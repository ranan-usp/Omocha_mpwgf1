magic
tech gf180mcuD
magscale 1 10
timestamp 1701760189
<< checkpaint >>
rect -2334 -2356 2334 2356
<< pwell >>
rect -334 -356 334 356
<< mvnmos >>
rect -70 -100 70 100
<< mvndiff >>
rect -158 87 -70 100
rect -158 -87 -145 87
rect -99 -87 -70 87
rect -158 -100 -70 -87
rect 70 87 158 100
rect 70 -87 99 87
rect 145 -87 158 87
rect 70 -100 158 -87
<< mvndiffc >>
rect -145 -87 -99 87
rect 99 -87 145 87
<< mvpsubdiff >>
rect -302 252 302 324
rect -302 -252 -230 252
rect 230 -252 302 252
rect -302 -265 302 -252
rect -302 -311 -186 -265
rect 186 -311 302 -265
rect -302 -324 302 -311
<< mvpsubdiffcont >>
rect -186 -311 186 -265
<< polysilicon >>
rect -70 179 70 192
rect -70 133 -57 179
rect 57 133 70 179
rect -70 100 70 133
rect -70 -183 70 -100
<< polycontact >>
rect -57 133 57 179
<< metal1 >>
rect -68 133 -57 179
rect 57 133 68 179
rect -145 87 -99 83
rect -145 -98 -99 -102
rect 99 87 145 83
rect 99 -98 145 -102
<< labels >>
flabel metal1 0 31 0 31 0 FreeSans 240 0 0 0 G
<< properties >>
string FIXED_BBOX -266 -288 266 288
<< end >>


