* NGSPICE file created from carray.ext - technology: gf180mcuD

.subckt carray n9 n0 n8 n7 n6 n5 n4 n3 n2 n1 ndum
C0 n8 cap_unit_9/out 0.420152p
C1 n2 ndum 0.041162f
C2 n9 cap_unit_9/out 0.846153p
C3 ndum n7 0.06073f
C4 n1 n5 0.134705f
C5 cap_unit_9/out n4 26.32268f
C6 ndum n3 0.025424f
C7 n6 cap_unit_9/out 0.105055p
C8 n2 n5 0.207999f
C9 n8 n1 0.278221f
C10 n5 n7 3.36878f
C11 n9 n1 0.342393f
C12 n2 n8 0.770114f
C13 n8 n7 50.178104f
C14 n2 n9 0.996568f
C15 n0 cap_unit_9/out 1.684219f
C16 n9 n7 29.51607f
C17 n1 n4 0.134826f
C18 n3 n5 0.346757f
C19 n6 n1 0.134562f
C20 n2 n4 0.213096f
C21 ndum n5 0.025424f
C22 n8 n3 1.46111f
C23 n2 n6 0.207877f
C24 n4 n7 1.70387f
C25 n3 n9 1.911225f
C26 n6 n7 34.326103f
C27 ndum n8 0.097254f
C28 ndum n9 0.127951f
C29 n0 n1 8.469265f
C30 n3 n4 25.8929f
C31 n2 n0 0.099202f
C32 n6 n3 0.336612f
C33 ndum n4 0.025424f
C34 n0 n7 0.06073f
C35 ndum n6 0.025424f
C36 n8 n5 5.60732f
C37 n9 n5 7.39935f
C38 cap_unit_9/out n1 3.365891f
C39 n3 n0 0.051666f
C40 n8 n9 87.10265f
C41 n2 cap_unit_9/out 6.640605f
C42 n5 n4 27.491999f
C43 cap_unit_9/out n7 0.210032p
C44 n6 n5 28.589401f
C45 n8 n4 2.84323f
C46 n8 n6 11.2161f
C47 n9 n4 3.740571f
C48 n3 cap_unit_9/out 13.201303f
C49 n6 n9 14.716781f
C50 n2 n1 16.597801f
C51 n0 n5 0.025424f
C52 ndum cap_unit_9/out 1.640173f
C53 n1 n7 0.205173f
C54 n6 n4 0.614078f
C55 n8 n0 0.097254f
C56 n2 n7 0.485242f
C57 n9 n0 0.184985f
C58 n3 n1 0.137399f
C59 cap_unit_9/out n5 52.565495f
C60 n2 n3 22.8406f
C61 ndum n1 8.161696f
C62 n0 n4 0.040502f
C63 n3 n7 0.891504f
C64 n6 n0 0.025424f
C65 n4 VSUBS 42.229664f
C66 ndum VSUBS 13.717415f
C67 n5 VSUBS 53.137516f
C68 n9 VSUBS 0.118402p
C69 cap_unit_9/out VSUBS 0.11849p
C70 n8 VSUBS 89.94086f
C71 n7 VSUBS 82.3075f
C72 n6 VSUBS 66.7443f
C73 n0 VSUBS 16.393326f
C74 n2 VSUBS 30.40069f
C75 n1 VSUBS 16.634346f
C76 n3 VSUBS 34.668854f
.ends

