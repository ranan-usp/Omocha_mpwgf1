magic
tech gf180mcuD
magscale 1 10
timestamp 1701965359
<< obsm1 >>
rect 216059 225784 408304 278832
<< metal2 >>
rect 11032 595560 11256 597000
rect 33096 595560 33320 597000
rect 55160 595560 55384 597000
rect 77224 595560 77448 597000
rect 99288 595560 99512 597000
rect 121352 595560 121576 597000
rect 143416 595560 143640 597000
rect 165480 595560 165704 597000
rect 187544 595560 187768 597000
rect 209608 595560 209832 597000
rect 231672 595560 231896 597000
rect 253736 595560 253960 597000
rect 275800 595560 276024 597000
rect 297864 595560 298088 597000
rect 319928 595560 320152 597000
rect 341992 595560 342216 597000
rect 364056 595560 364280 597000
rect 386120 595560 386344 597000
rect 408184 595560 408408 597000
rect 430248 595560 430472 597000
rect 452312 595560 452536 597000
rect 474376 595560 474600 597000
rect 496440 595560 496664 597000
rect 518504 595560 518728 597000
rect 540568 595560 540792 597000
rect 562632 595560 562856 597000
rect 584696 595560 584920 597000
rect 11368 -960 11592 480
rect 13272 -960 13496 480
rect 15176 -960 15400 480
rect 17080 -960 17304 480
rect 18984 -960 19208 480
rect 20888 -960 21112 480
rect 22792 -960 23016 480
rect 24696 -960 24920 480
rect 26600 -960 26824 480
rect 28504 -960 28728 480
rect 30408 -960 30632 480
rect 32312 -960 32536 480
rect 34216 -960 34440 480
rect 36120 -960 36344 480
rect 38024 -960 38248 480
rect 39928 -960 40152 480
rect 41832 -960 42056 480
rect 43736 -960 43960 480
rect 45640 -960 45864 480
rect 47544 -960 47768 480
rect 49448 -960 49672 480
rect 51352 -960 51576 480
rect 53256 -960 53480 480
rect 55160 -960 55384 480
rect 57064 -960 57288 480
rect 58968 -960 59192 480
rect 60872 -960 61096 480
rect 62776 -960 63000 480
rect 64680 -960 64904 480
rect 66584 -960 66808 480
rect 68488 -960 68712 480
rect 70392 -960 70616 480
rect 72296 -960 72520 480
rect 74200 -960 74424 480
rect 76104 -960 76328 480
rect 78008 -960 78232 480
rect 79912 -960 80136 480
rect 81816 -960 82040 480
rect 83720 -960 83944 480
rect 85624 -960 85848 480
rect 87528 -960 87752 480
rect 89432 -960 89656 480
rect 91336 -960 91560 480
rect 93240 -960 93464 480
rect 95144 -960 95368 480
rect 97048 -960 97272 480
rect 98952 -960 99176 480
rect 100856 -960 101080 480
rect 102760 -960 102984 480
rect 104664 -960 104888 480
rect 106568 -960 106792 480
rect 108472 -960 108696 480
rect 110376 -960 110600 480
rect 112280 -960 112504 480
rect 114184 -960 114408 480
rect 116088 -960 116312 480
rect 117992 -960 118216 480
rect 119896 -960 120120 480
rect 121800 -960 122024 480
rect 123704 -960 123928 480
rect 125608 -960 125832 480
rect 127512 -960 127736 480
rect 129416 -960 129640 480
rect 131320 -960 131544 480
rect 133224 -960 133448 480
rect 135128 -960 135352 480
rect 137032 -960 137256 480
rect 138936 -960 139160 480
rect 140840 -960 141064 480
rect 142744 -960 142968 480
rect 144648 -960 144872 480
rect 146552 -960 146776 480
rect 148456 -960 148680 480
rect 150360 -960 150584 480
rect 152264 -960 152488 480
rect 154168 -960 154392 480
rect 156072 -960 156296 480
rect 157976 -960 158200 480
rect 159880 -960 160104 480
rect 161784 -960 162008 480
rect 163688 -960 163912 480
rect 165592 -960 165816 480
rect 167496 -960 167720 480
rect 169400 -960 169624 480
rect 171304 -960 171528 480
rect 173208 -960 173432 480
rect 175112 -960 175336 480
rect 177016 -960 177240 480
rect 178920 -960 179144 480
rect 180824 -960 181048 480
rect 182728 -960 182952 480
rect 184632 -960 184856 480
rect 186536 -960 186760 480
rect 188440 -960 188664 480
rect 190344 -960 190568 480
rect 192248 -960 192472 480
rect 194152 -960 194376 480
rect 196056 -960 196280 480
rect 197960 -960 198184 480
rect 199864 -960 200088 480
rect 201768 -960 201992 480
rect 203672 -960 203896 480
rect 205576 -960 205800 480
rect 207480 -960 207704 480
rect 209384 -960 209608 480
rect 211288 -960 211512 480
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580664 -960 580888 480
rect 582568 -960 582792 480
rect 584472 -960 584696 480
<< obsm2 >>
rect 11340 540 574980 577440
rect 11652 392 13212 540
rect 13556 392 15116 540
rect 15460 392 17020 540
rect 17364 392 18924 540
rect 19268 392 20828 540
rect 21172 392 22732 540
rect 23076 392 24636 540
rect 24980 392 26540 540
rect 26884 392 28444 540
rect 28788 392 30348 540
rect 30692 392 32252 540
rect 32596 392 34156 540
rect 34500 392 36060 540
rect 36404 392 37964 540
rect 38308 392 39868 540
rect 40212 392 41772 540
rect 42116 392 43676 540
rect 44020 392 45580 540
rect 45924 392 47484 540
rect 47828 392 49388 540
rect 49732 392 51292 540
rect 51636 392 53196 540
rect 53540 392 55100 540
rect 55444 392 57004 540
rect 57348 392 58908 540
rect 59252 392 60812 540
rect 61156 392 62716 540
rect 63060 392 64620 540
rect 64964 392 66524 540
rect 66868 392 68428 540
rect 68772 392 70332 540
rect 70676 392 72236 540
rect 72580 392 74140 540
rect 74484 392 76044 540
rect 76388 392 77948 540
rect 78292 392 79852 540
rect 80196 392 81756 540
rect 82100 392 83660 540
rect 84004 392 85564 540
rect 85908 392 87468 540
rect 87812 392 89372 540
rect 89716 392 91276 540
rect 91620 392 93180 540
rect 93524 392 95084 540
rect 95428 392 96988 540
rect 97332 392 98892 540
rect 99236 392 100796 540
rect 101140 392 102700 540
rect 103044 392 104604 540
rect 104948 392 106508 540
rect 106852 392 108412 540
rect 108756 392 110316 540
rect 110660 392 112220 540
rect 112564 392 114124 540
rect 114468 392 116028 540
rect 116372 392 117932 540
rect 118276 392 119836 540
rect 120180 392 121740 540
rect 122084 392 123644 540
rect 123988 392 125548 540
rect 125892 392 127452 540
rect 127796 392 129356 540
rect 129700 392 131260 540
rect 131604 392 133164 540
rect 133508 392 135068 540
rect 135412 392 136972 540
rect 137316 392 138876 540
rect 139220 392 140780 540
rect 141124 392 142684 540
rect 143028 392 144588 540
rect 144932 392 146492 540
rect 146836 392 148396 540
rect 148740 392 150300 540
rect 150644 392 152204 540
rect 152548 392 154108 540
rect 154452 392 156012 540
rect 156356 392 157916 540
rect 158260 392 159820 540
rect 160164 392 161724 540
rect 162068 392 163628 540
rect 163972 392 165532 540
rect 165876 392 167436 540
rect 167780 392 169340 540
rect 169684 392 171244 540
rect 171588 392 173148 540
rect 173492 392 175052 540
rect 175396 392 176956 540
rect 177300 392 178860 540
rect 179204 392 180764 540
rect 181108 392 182668 540
rect 183012 392 184572 540
rect 184916 392 186476 540
rect 186820 392 188380 540
rect 188724 392 190284 540
rect 190628 392 192188 540
rect 192532 392 194092 540
rect 194436 392 195996 540
rect 196340 392 197900 540
rect 198244 392 199804 540
rect 200148 392 201708 540
rect 202052 392 203612 540
rect 203956 392 205516 540
rect 205860 392 207420 540
rect 207764 392 209324 540
rect 209668 392 211228 540
rect 211572 392 213132 540
rect 213476 392 215036 540
rect 215380 392 216940 540
rect 217284 392 218844 540
rect 219188 392 220748 540
rect 221092 392 222652 540
rect 222996 392 224556 540
rect 224900 392 226460 540
rect 226804 392 228364 540
rect 228708 392 230268 540
rect 230612 392 232172 540
rect 232516 392 234076 540
rect 234420 392 235980 540
rect 236324 392 237884 540
rect 238228 392 239788 540
rect 240132 392 241692 540
rect 242036 392 243596 540
rect 243940 392 245500 540
rect 245844 392 247404 540
rect 247748 392 249308 540
rect 249652 392 251212 540
rect 251556 392 253116 540
rect 253460 392 255020 540
rect 255364 392 256924 540
rect 257268 392 258828 540
rect 259172 392 260732 540
rect 261076 392 262636 540
rect 262980 392 264540 540
rect 264884 392 266444 540
rect 266788 392 268348 540
rect 268692 392 270252 540
rect 270596 392 272156 540
rect 272500 392 274060 540
rect 274404 392 275964 540
rect 276308 392 277868 540
rect 278212 392 279772 540
rect 280116 392 281676 540
rect 282020 392 283580 540
rect 283924 392 285484 540
rect 285828 392 287388 540
rect 287732 392 289292 540
rect 289636 392 291196 540
rect 291540 392 293100 540
rect 293444 392 295004 540
rect 295348 392 296908 540
rect 297252 392 298812 540
rect 299156 392 300716 540
rect 301060 392 302620 540
rect 302964 392 304524 540
rect 304868 392 306428 540
rect 306772 392 308332 540
rect 308676 392 310236 540
rect 310580 392 312140 540
rect 312484 392 314044 540
rect 314388 392 315948 540
rect 316292 392 317852 540
rect 318196 392 319756 540
rect 320100 392 321660 540
rect 322004 392 323564 540
rect 323908 392 325468 540
rect 325812 392 327372 540
rect 327716 392 329276 540
rect 329620 392 331180 540
rect 331524 392 333084 540
rect 333428 392 334988 540
rect 335332 392 336892 540
rect 337236 392 338796 540
rect 339140 392 340700 540
rect 341044 392 342604 540
rect 342948 392 344508 540
rect 344852 392 346412 540
rect 346756 392 348316 540
rect 348660 392 350220 540
rect 350564 392 352124 540
rect 352468 392 354028 540
rect 354372 392 355932 540
rect 356276 392 357836 540
rect 358180 392 359740 540
rect 360084 392 361644 540
rect 361988 392 363548 540
rect 363892 392 365452 540
rect 365796 392 367356 540
rect 367700 392 369260 540
rect 369604 392 371164 540
rect 371508 392 373068 540
rect 373412 392 374972 540
rect 375316 392 376876 540
rect 377220 392 378780 540
rect 379124 392 380684 540
rect 381028 392 382588 540
rect 382932 392 384492 540
rect 384836 392 386396 540
rect 386740 392 388300 540
rect 388644 392 390204 540
rect 390548 392 392108 540
rect 392452 392 394012 540
rect 394356 392 395916 540
rect 396260 392 397820 540
rect 398164 392 399724 540
rect 400068 392 401628 540
rect 401972 392 403532 540
rect 403876 392 405436 540
rect 405780 392 407340 540
rect 407684 392 409244 540
rect 409588 392 411148 540
rect 411492 392 413052 540
rect 413396 392 414956 540
rect 415300 392 416860 540
rect 417204 392 418764 540
rect 419108 392 420668 540
rect 421012 392 422572 540
rect 422916 392 424476 540
rect 424820 392 426380 540
rect 426724 392 428284 540
rect 428628 392 430188 540
rect 430532 392 432092 540
rect 432436 392 433996 540
rect 434340 392 435900 540
rect 436244 392 437804 540
rect 438148 392 439708 540
rect 440052 392 441612 540
rect 441956 392 443516 540
rect 443860 392 445420 540
rect 445764 392 447324 540
rect 447668 392 449228 540
rect 449572 392 451132 540
rect 451476 392 453036 540
rect 453380 392 454940 540
rect 455284 392 456844 540
rect 457188 392 458748 540
rect 459092 392 460652 540
rect 460996 392 462556 540
rect 462900 392 464460 540
rect 464804 392 466364 540
rect 466708 392 468268 540
rect 468612 392 470172 540
rect 470516 392 472076 540
rect 472420 392 473980 540
rect 474324 392 475884 540
rect 476228 392 477788 540
rect 478132 392 479692 540
rect 480036 392 481596 540
rect 481940 392 483500 540
rect 483844 392 485404 540
rect 485748 392 487308 540
rect 487652 392 489212 540
rect 489556 392 491116 540
rect 491460 392 493020 540
rect 493364 392 494924 540
rect 495268 392 496828 540
rect 497172 392 498732 540
rect 499076 392 500636 540
rect 500980 392 502540 540
rect 502884 392 504444 540
rect 504788 392 506348 540
rect 506692 392 508252 540
rect 508596 392 510156 540
rect 510500 392 512060 540
rect 512404 392 513964 540
rect 514308 392 515868 540
rect 516212 392 517772 540
rect 518116 392 519676 540
rect 520020 392 521580 540
rect 521924 392 523484 540
rect 523828 392 525388 540
rect 525732 392 527292 540
rect 527636 392 529196 540
rect 529540 392 531100 540
rect 531444 392 533004 540
rect 533348 392 534908 540
rect 535252 392 536812 540
rect 537156 392 538716 540
rect 539060 392 540620 540
rect 540964 392 542524 540
rect 542868 392 544428 540
rect 544772 392 546332 540
rect 546676 392 548236 540
rect 548580 392 550140 540
rect 550484 392 552044 540
rect 552388 392 553948 540
rect 554292 392 555852 540
rect 556196 392 557756 540
rect 558100 392 559660 540
rect 560004 392 561564 540
rect 561908 392 563468 540
rect 563812 392 565372 540
rect 565716 392 567276 540
rect 567620 392 569180 540
rect 569524 392 571084 540
rect 571428 392 572988 540
rect 573332 392 574892 540
<< metal3 >>
rect 595560 588616 597000 588840
rect -960 587160 480 587384
rect 595560 575400 597000 575624
rect -960 573048 480 573272
rect 595560 562184 597000 562408
rect -960 558936 480 559160
rect 595560 548968 597000 549192
rect -960 544824 480 545048
rect 595560 535752 597000 535976
rect -960 530712 480 530936
rect 595560 522536 597000 522760
rect -960 516600 480 516824
rect 595560 509320 597000 509544
rect -960 502488 480 502712
rect 595560 496104 597000 496328
rect -960 488376 480 488600
rect 595560 482888 597000 483112
rect -960 474264 480 474488
rect 595560 469672 597000 469896
rect -960 460152 480 460376
rect 595560 456456 597000 456680
rect -960 446040 480 446264
rect 595560 443240 597000 443464
rect -960 431928 480 432152
rect 595560 430024 597000 430248
rect -960 417816 480 418040
rect 595560 416808 597000 417032
rect -960 403704 480 403928
rect 595560 403592 597000 403816
rect 595560 390376 597000 390600
rect -960 389592 480 389816
rect 595560 377160 597000 377384
rect -960 375480 480 375704
rect 595560 363944 597000 364168
rect -960 361368 480 361592
rect 595560 350728 597000 350952
rect -960 347256 480 347480
rect 595560 337512 597000 337736
rect -960 333144 480 333368
rect 595560 324296 597000 324520
rect -960 319032 480 319256
rect 595560 311080 597000 311304
rect -960 304920 480 305144
rect 595560 297864 597000 298088
rect -960 290808 480 291032
rect 595560 284648 597000 284872
rect -960 276696 480 276920
rect 595560 271432 597000 271656
rect -960 262584 480 262808
rect 595560 258216 597000 258440
rect -960 248472 480 248696
rect 595560 245000 597000 245224
rect -960 234360 480 234584
rect 595560 231784 597000 232008
rect -960 220248 480 220472
rect 595560 218568 597000 218792
rect -960 206136 480 206360
rect 595560 205352 597000 205576
rect -960 192024 480 192248
rect 595560 192136 597000 192360
rect 595560 178920 597000 179144
rect -960 177912 480 178136
rect 595560 165704 597000 165928
rect -960 163800 480 164024
rect 595560 152488 597000 152712
rect -960 149688 480 149912
rect 595560 139272 597000 139496
rect -960 135576 480 135800
rect 595560 126056 597000 126280
rect -960 121464 480 121688
rect 595560 112840 597000 113064
rect -960 107352 480 107576
rect 595560 99624 597000 99848
rect -960 93240 480 93464
rect 595560 86408 597000 86632
rect -960 79128 480 79352
rect 595560 73192 597000 73416
rect -960 65016 480 65240
rect 595560 59976 597000 60200
rect -960 50904 480 51128
rect 595560 46760 597000 46984
rect -960 36792 480 37016
rect 595560 33544 597000 33768
rect -960 22680 480 22904
rect 595560 20328 597000 20552
rect -960 8568 480 8792
rect 595560 7112 597000 7336
<< obsm3 >>
rect 392 573332 574990 577440
rect 540 572988 574990 573332
rect 392 559220 574990 572988
rect 540 558876 574990 559220
rect 392 545108 574990 558876
rect 540 544764 574990 545108
rect 392 530996 574990 544764
rect 540 530652 574990 530996
rect 392 516884 574990 530652
rect 540 516540 574990 516884
rect 392 502772 574990 516540
rect 540 502428 574990 502772
rect 392 488660 574990 502428
rect 540 488316 574990 488660
rect 392 474548 574990 488316
rect 540 474204 574990 474548
rect 392 460436 574990 474204
rect 540 460092 574990 460436
rect 392 446324 574990 460092
rect 540 445980 574990 446324
rect 392 432212 574990 445980
rect 540 431868 574990 432212
rect 392 418100 574990 431868
rect 540 417756 574990 418100
rect 392 403988 574990 417756
rect 540 403644 574990 403988
rect 392 389876 574990 403644
rect 540 389532 574990 389876
rect 392 375764 574990 389532
rect 540 375420 574990 375764
rect 392 361652 574990 375420
rect 540 361308 574990 361652
rect 392 347540 574990 361308
rect 540 347196 574990 347540
rect 392 333428 574990 347196
rect 540 333084 574990 333428
rect 392 319316 574990 333084
rect 540 318972 574990 319316
rect 392 305204 574990 318972
rect 540 304860 574990 305204
rect 392 291092 574990 304860
rect 540 290748 574990 291092
rect 392 276980 574990 290748
rect 540 276636 574990 276980
rect 392 262868 574990 276636
rect 540 262524 574990 262868
rect 392 248756 574990 262524
rect 540 248412 574990 248756
rect 392 234644 574990 248412
rect 540 234300 574990 234644
rect 392 220532 574990 234300
rect 540 220188 574990 220532
rect 392 206420 574990 220188
rect 540 206076 574990 206420
rect 392 192308 574990 206076
rect 540 191964 574990 192308
rect 392 178196 574990 191964
rect 540 177852 574990 178196
rect 392 164084 574990 177852
rect 540 163740 574990 164084
rect 392 149972 574990 163740
rect 540 149628 574990 149972
rect 392 135860 574990 149628
rect 540 135516 574990 135860
rect 392 121748 574990 135516
rect 540 121404 574990 121748
rect 392 107636 574990 121404
rect 540 107292 574990 107636
rect 392 93524 574990 107292
rect 540 93180 574990 93524
rect 392 79412 574990 93180
rect 540 79068 574990 79412
rect 392 65300 574990 79068
rect 540 64956 574990 65300
rect 392 51188 574990 64956
rect 540 50844 574990 51188
rect 392 37076 574990 50844
rect 540 36732 574990 37076
rect 392 22964 574990 36732
rect 540 22620 574990 22964
rect 392 8852 574990 22620
rect 540 8508 574990 8852
rect 392 4172 574990 8508
<< metal4 >>
rect -1916 -1644 -1296 598268
rect -956 -684 -336 597308
rect 5418 -1644 6038 598268
rect 9138 -1644 9758 598268
rect 36138 550512 36758 598268
rect 39858 560472 40478 598268
rect 66858 551592 67478 598268
rect 70578 541632 71198 598268
rect 97578 573912 98198 598268
rect 101298 568272 101918 598268
rect 128298 577636 128918 598268
rect 132018 577636 132638 598268
rect 159018 563592 159638 598268
rect 162738 573432 163358 598268
rect 36138 -1644 36758 517448
rect 39858 -1644 40478 527288
rect 66858 -1644 67478 518408
rect 70578 -1644 71198 508448
rect 97578 -1644 98198 553328
rect 189738 549192 190358 598268
rect 101298 -1644 101918 547808
rect 193458 539352 194078 598268
rect 220458 572592 221078 598268
rect 224178 566952 224798 598268
rect 251178 577632 251798 598268
rect 254898 577632 255518 598268
rect 128298 -1644 128918 507368
rect 132018 -1644 132638 507368
rect 159018 487164 159638 519728
rect 162738 487164 163358 529328
rect 220458 487164 221078 546008
rect 224178 487164 224798 540488
rect 281898 487164 282518 598268
rect 285618 487164 286238 598268
rect 312618 487164 313238 598268
rect 316338 487164 316958 598268
rect 343338 487164 343958 598268
rect 347058 487164 347678 598268
rect 374058 487164 374678 598268
rect 377778 487164 378398 598268
rect 404778 487164 405398 598268
rect 408498 487164 409118 598268
rect 435498 487164 436118 598268
rect 439218 487164 439838 598268
rect 466218 487164 466838 598268
rect 469938 487164 470558 598268
rect 159018 -1644 159638 17452
rect 162738 -1644 163358 17452
rect 189738 -1644 190358 17452
rect 193458 -1644 194078 17452
rect 220458 -1644 221078 17452
rect 224178 -1644 224798 17452
rect 251178 -1644 251798 17452
rect 254898 -1644 255518 17452
rect 281898 -1644 282518 17452
rect 285618 -1644 286238 17452
rect 312618 -1644 313238 17452
rect 316338 -1644 316958 17452
rect 343338 -1644 343958 17452
rect 347058 -1644 347678 17452
rect 374058 -1644 374678 17452
rect 377778 -1644 378398 17452
rect 404778 -1644 405398 17452
rect 408498 -1644 409118 17452
rect 435498 -1644 436118 17452
rect 439218 -1644 439838 17452
rect 466218 -1644 466838 17452
rect 469938 -1644 470558 17452
rect 496938 -1644 497558 598268
rect 500658 -1644 501278 598268
rect 527658 -1644 528278 598268
rect 531378 -1644 531998 598268
rect 558378 -1644 558998 598268
rect 562098 -1644 562718 598268
rect 589098 -1644 589718 598268
rect 592818 -1644 593438 598268
rect 596400 -684 597020 597308
rect 597360 -1644 597980 598268
<< obsm4 >>
rect 4172 19568 5358 575940
rect 6098 19568 9078 575940
rect 9818 550452 36078 575940
rect 36818 560412 39798 575940
rect 40538 560412 66798 575940
rect 36818 551532 66798 560412
rect 67538 551532 70518 575940
rect 36818 550452 70518 551532
rect 9818 541572 70518 550452
rect 71258 573852 97518 575940
rect 98258 573852 101238 575940
rect 71258 568212 101238 573852
rect 101978 568212 158958 575940
rect 71258 563532 158958 568212
rect 159698 573372 162678 575940
rect 163418 573372 189678 575940
rect 159698 563532 189678 573372
rect 71258 553388 189678 563532
rect 71258 541572 97518 553388
rect 9818 527348 97518 541572
rect 9818 517508 39798 527348
rect 9818 19568 36078 517508
rect 36818 19568 39798 517508
rect 40538 518468 97518 527348
rect 40538 19568 66798 518468
rect 67538 508508 97518 518468
rect 67538 19568 70518 508508
rect 71258 19568 97518 508508
rect 98258 549132 189678 553388
rect 190418 549132 193398 575940
rect 98258 547868 193398 549132
rect 98258 19568 101238 547868
rect 101978 539292 193398 547868
rect 194138 572532 220398 575940
rect 221138 572532 224118 575940
rect 194138 566892 224118 572532
rect 224858 566892 281838 575940
rect 194138 546068 281838 566892
rect 194138 539292 220398 546068
rect 101978 529388 220398 539292
rect 101978 519788 162678 529388
rect 101978 507428 158958 519788
rect 101978 19568 128238 507428
rect 128978 19568 131958 507428
rect 132698 487104 158958 507428
rect 159698 487104 162678 519788
rect 163418 487104 220398 529388
rect 221138 540548 281838 546068
rect 221138 487104 224118 540548
rect 224858 487104 281838 540548
rect 282578 487104 285558 575940
rect 286298 487104 312558 575940
rect 313298 487104 316278 575940
rect 317018 487104 343278 575940
rect 344018 487104 346998 575940
rect 347738 487104 373998 575940
rect 374738 487104 377718 575940
rect 378458 487104 404718 575940
rect 405458 487104 408438 575940
rect 409178 487104 435438 575940
rect 436178 487104 439158 575940
rect 439898 487104 466158 575940
rect 466898 487104 469878 575940
rect 470618 487104 483960 575940
rect 132698 19568 483960 487104
<< metal5 >>
rect -1916 597648 597980 598268
rect -956 596688 597020 597308
rect -1916 586636 597980 587636
rect -1916 579636 597980 580636
rect -1916 568636 597980 569636
rect -1916 561636 597980 562636
rect -1916 550636 597980 551636
rect -1916 543636 597980 544636
rect -1916 532636 597980 533636
rect -1916 525636 597980 526636
rect -1916 514636 597980 515636
rect -1916 507636 597980 508636
rect -1916 496636 597980 497636
rect -1916 489636 597980 490636
rect -1916 478636 597980 479636
rect -1916 471636 597980 472636
rect -1916 460636 597980 461636
rect -1916 453636 597980 454636
rect -1916 442636 189012 443636
rect 442948 442636 597980 443636
rect -1916 435636 189012 436636
rect 442948 435636 597980 436636
rect -1916 424636 189012 425636
rect 442948 424636 597980 425636
rect -1916 417636 189012 418636
rect 442948 417636 597980 418636
rect -1916 406636 189012 407636
rect 442948 406636 597980 407636
rect -1916 399636 189012 400636
rect 442948 399636 597980 400636
rect -1916 388636 189012 389636
rect 442948 388636 597980 389636
rect -1916 381636 189012 382636
rect 442948 381636 597980 382636
rect -1916 370636 189012 371636
rect 442948 370636 597980 371636
rect -1916 363636 152116 364636
rect -1916 352636 152116 353636
rect -1916 345636 152116 346636
rect -1916 334636 152116 335636
rect -1916 327636 152116 328636
rect -1916 316636 152116 317636
rect -1916 309636 152116 310636
rect -1916 298636 152116 299636
rect -1916 291636 152116 292636
rect -1916 280636 152116 281636
rect -1916 273636 152116 274636
rect -1916 262636 152116 263636
rect -1916 255636 152116 256636
rect -1916 244636 152116 245636
rect -1916 237636 152116 238636
rect -1916 226636 152116 227636
rect -1916 219636 152116 220636
rect -1916 208636 152116 209636
rect -1916 201636 152116 202636
rect -1916 190636 152116 191636
rect -1916 183636 152116 184636
rect -1916 172636 152116 173636
rect -1916 165636 152116 166636
rect -1916 154636 152116 155636
rect -1916 147636 152116 148636
rect 479844 363636 597980 364636
rect 479844 352636 597980 353636
rect 479844 345636 597980 346636
rect 479844 334636 597980 335636
rect 479844 327636 597980 328636
rect 479844 316636 597980 317636
rect 479844 309636 597980 310636
rect 479844 298636 597980 299636
rect 479844 291636 597980 292636
rect 479844 280636 597980 281636
rect 479844 273636 597980 274636
rect 479844 262636 597980 263636
rect 479844 255636 597980 256636
rect 479844 244636 597980 245636
rect 479844 237636 597980 238636
rect 479844 226636 597980 227636
rect 479844 219636 597980 220636
rect 479844 208636 597980 209636
rect 479844 201636 597980 202636
rect 479844 190636 597980 191636
rect 479844 183636 597980 184636
rect 479844 172636 597980 173636
rect 479844 165636 597980 166636
rect 479844 154636 597980 155636
rect 479844 147636 597980 148636
rect -1916 136636 189012 137636
rect 442948 136636 597980 137636
rect -1916 129636 189012 130636
rect 442948 129636 597980 130636
rect -1916 118636 189012 119636
rect 442948 118636 597980 119636
rect -1916 111636 189012 112636
rect 442948 111636 597980 112636
rect -1916 100636 189012 101636
rect 442948 100636 597980 101636
rect -1916 93636 189012 94636
rect 442948 93636 597980 94636
rect -1916 82636 189012 83636
rect 442948 82636 597980 83636
rect -1916 75636 189012 76636
rect 442948 75636 597980 76636
rect -1916 64636 189012 65636
rect 442948 64636 597980 65636
rect -1916 57636 189012 58636
rect 442948 57636 597980 58636
rect -1916 46636 597980 47636
rect -1916 39636 597980 40636
rect -1916 28636 597980 29636
rect -1916 21636 597980 22636
rect -1916 10636 597980 11636
rect -1916 3636 597980 4636
rect -956 -684 597020 -64
rect -1916 -1644 597980 -1024
<< obsm5 >>
rect 154300 443736 477660 447548
rect 189112 442536 442848 443736
rect 154300 436736 477660 442536
rect 189112 435536 442848 436736
rect 154300 425736 477660 435536
rect 189112 424536 442848 425736
rect 154300 418736 477660 424536
rect 189112 417536 442848 418736
rect 154300 407736 477660 417536
rect 189112 406536 442848 407736
rect 154300 400736 477660 406536
rect 189112 399536 442848 400736
rect 154300 389736 477660 399536
rect 189112 388536 442848 389736
rect 154300 382736 477660 388536
rect 189112 381536 442848 382736
rect 154300 371736 477660 381536
rect 189112 370536 442848 371736
rect 154300 137736 477660 370536
rect 189112 136536 442848 137736
rect 154300 130736 477660 136536
rect 189112 129536 442848 130736
rect 154300 119736 477660 129536
rect 189112 118536 442848 119736
rect 154300 112736 477660 118536
rect 189112 111536 442848 112736
rect 154300 101736 477660 111536
rect 189112 100536 442848 101736
rect 154300 94736 477660 100536
rect 189112 93536 442848 94736
rect 154300 83736 477660 93536
rect 189112 82536 442848 83736
rect 154300 76736 477660 82536
rect 189112 75536 442848 76736
rect 154300 65736 477660 75536
rect 189112 64536 442848 65736
rect 154300 58736 477660 64536
rect 189112 57536 442848 58736
rect 154300 57068 477660 57536
<< labels >>
rlabel metal3 s 595560 7112 597000 7336 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 595560 403592 597000 403816 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 595560 443240 597000 443464 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 595560 482888 597000 483112 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 595560 522536 597000 522760 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 595560 562184 597000 562408 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 584696 595560 584920 597000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 518504 595560 518728 597000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 452312 595560 452536 597000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 386120 595560 386344 597000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 319928 595560 320152 597000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 595560 46760 597000 46984 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 253736 595560 253960 597000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 187544 595560 187768 597000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 121352 595560 121576 597000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 55160 595560 55384 597000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -960 587160 480 587384 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -960 544824 480 545048 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -960 502488 480 502712 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -960 460152 480 460376 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -960 417816 480 418040 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -960 375480 480 375704 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 595560 86408 597000 86632 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -960 333144 480 333368 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -960 290808 480 291032 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -960 248472 480 248696 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -960 206136 480 206360 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -960 163800 480 164024 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -960 121464 480 121688 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -960 79128 480 79352 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -960 36792 480 37016 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 595560 126056 597000 126280 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 595560 165704 597000 165928 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 595560 205352 597000 205576 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 595560 245000 597000 245224 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 595560 284648 597000 284872 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 595560 324296 597000 324520 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 595560 363944 597000 364168 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 595560 33544 597000 33768 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 595560 430024 597000 430248 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 595560 469672 597000 469896 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 595560 509320 597000 509544 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 595560 548968 597000 549192 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 595560 588616 597000 588840 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 540568 595560 540792 597000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 474376 595560 474600 597000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 408184 595560 408408 597000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 341992 595560 342216 597000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 275800 595560 276024 597000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 595560 73192 597000 73416 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 209608 595560 209832 597000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 143416 595560 143640 597000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 77224 595560 77448 597000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 11032 595560 11256 597000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -960 558936 480 559160 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -960 516600 480 516824 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -960 474264 480 474488 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -960 431928 480 432152 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -960 389592 480 389816 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -960 347256 480 347480 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 595560 112840 597000 113064 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -960 304920 480 305144 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -960 262584 480 262808 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -960 220248 480 220472 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -960 177912 480 178136 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -960 135576 480 135800 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -960 93240 480 93464 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -960 50904 480 51128 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -960 8568 480 8792 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 595560 152488 597000 152712 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 595560 192136 597000 192360 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 595560 231784 597000 232008 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 595560 271432 597000 271656 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 595560 311080 597000 311304 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 595560 350728 597000 350952 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 595560 390376 597000 390600 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 595560 20328 597000 20552 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 595560 416808 597000 417032 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 595560 456456 597000 456680 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 595560 496104 597000 496328 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 595560 535752 597000 535976 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 595560 575400 597000 575624 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 562632 595560 562856 597000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 496440 595560 496664 597000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 430248 595560 430472 597000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 364056 595560 364280 597000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 297864 595560 298088 597000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 595560 59976 597000 60200 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 231672 595560 231896 597000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 165480 595560 165704 597000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 99288 595560 99512 597000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 33096 595560 33320 597000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -960 573048 480 573272 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -960 530712 480 530936 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -960 488376 480 488600 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -960 446040 480 446264 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -960 403704 480 403928 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -960 361368 480 361592 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 595560 99624 597000 99848 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -960 319032 480 319256 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -960 276696 480 276920 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -960 234360 480 234584 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -960 192024 480 192248 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -960 149688 480 149912 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -960 107352 480 107576 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -960 65016 480 65240 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -960 22680 480 22904 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 595560 139272 597000 139496 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 595560 178920 597000 179144 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 595560 218568 597000 218792 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 595560 258216 597000 258440 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 595560 297864 597000 298088 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 595560 337512 597000 337736 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 595560 377160 597000 377384 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 213192 -960 213416 480 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 270312 -960 270536 480 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 276024 -960 276248 480 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 281736 -960 281960 480 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 287448 -960 287672 480 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 293160 -960 293384 480 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 298872 -960 299096 480 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 304584 -960 304808 480 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 310296 -960 310520 480 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 316008 -960 316232 480 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 321720 -960 321944 480 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 218904 -960 219128 480 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 327432 -960 327656 480 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 333144 -960 333368 480 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 338856 -960 339080 480 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 344568 -960 344792 480 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 350280 -960 350504 480 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 355992 -960 356216 480 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 361704 -960 361928 480 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 367416 -960 367640 480 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 373128 -960 373352 480 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 378840 -960 379064 480 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 224616 -960 224840 480 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 384552 -960 384776 480 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 390264 -960 390488 480 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 395976 -960 396200 480 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 401688 -960 401912 480 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 407400 -960 407624 480 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 413112 -960 413336 480 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 418824 -960 419048 480 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 424536 -960 424760 480 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 430248 -960 430472 480 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 435960 -960 436184 480 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 230328 -960 230552 480 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 441672 -960 441896 480 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 447384 -960 447608 480 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 453096 -960 453320 480 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 458808 -960 459032 480 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 464520 -960 464744 480 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 470232 -960 470456 480 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 475944 -960 476168 480 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 481656 -960 481880 480 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 487368 -960 487592 480 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 493080 -960 493304 480 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 236040 -960 236264 480 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 498792 -960 499016 480 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 504504 -960 504728 480 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 510216 -960 510440 480 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 515928 -960 516152 480 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 521640 -960 521864 480 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 527352 -960 527576 480 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 533064 -960 533288 480 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 538776 -960 539000 480 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 544488 -960 544712 480 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 550200 -960 550424 480 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 241752 -960 241976 480 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 555912 -960 556136 480 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 561624 -960 561848 480 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 567336 -960 567560 480 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 573048 -960 573272 480 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 247464 -960 247688 480 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 253176 -960 253400 480 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 258888 -960 259112 480 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 264600 -960 264824 480 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 215096 -960 215320 480 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 272216 -960 272440 480 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 277928 -960 278152 480 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 283640 -960 283864 480 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 289352 -960 289576 480 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 295064 -960 295288 480 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 300776 -960 301000 480 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 306488 -960 306712 480 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 312200 -960 312424 480 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 317912 -960 318136 480 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 323624 -960 323848 480 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 220808 -960 221032 480 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 329336 -960 329560 480 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 335048 -960 335272 480 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 340760 -960 340984 480 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 346472 -960 346696 480 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 352184 -960 352408 480 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 357896 -960 358120 480 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 363608 -960 363832 480 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 369320 -960 369544 480 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 375032 -960 375256 480 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 380744 -960 380968 480 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 226520 -960 226744 480 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 386456 -960 386680 480 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 392168 -960 392392 480 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 397880 -960 398104 480 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 403592 -960 403816 480 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 409304 -960 409528 480 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 415016 -960 415240 480 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 420728 -960 420952 480 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 426440 -960 426664 480 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 432152 -960 432376 480 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 437864 -960 438088 480 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 232232 -960 232456 480 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 443576 -960 443800 480 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 449288 -960 449512 480 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 455000 -960 455224 480 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 460712 -960 460936 480 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 466424 -960 466648 480 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 472136 -960 472360 480 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 477848 -960 478072 480 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 483560 -960 483784 480 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 489272 -960 489496 480 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 494984 -960 495208 480 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 237944 -960 238168 480 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 500696 -960 500920 480 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 506408 -960 506632 480 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 512120 -960 512344 480 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 517832 -960 518056 480 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 523544 -960 523768 480 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 529256 -960 529480 480 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 534968 -960 535192 480 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 540680 -960 540904 480 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 546392 -960 546616 480 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 552104 -960 552328 480 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 243656 -960 243880 480 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 557816 -960 558040 480 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 563528 -960 563752 480 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 569240 -960 569464 480 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 574952 -960 575176 480 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 249368 -960 249592 480 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 255080 -960 255304 480 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 260792 -960 261016 480 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 266504 -960 266728 480 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 217000 -960 217224 480 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 274120 -960 274344 480 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 279832 -960 280056 480 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 285544 -960 285768 480 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 291256 -960 291480 480 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 296968 -960 297192 480 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 302680 -960 302904 480 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 308392 -960 308616 480 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 314104 -960 314328 480 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 319816 -960 320040 480 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 325528 -960 325752 480 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 222712 -960 222936 480 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 331240 -960 331464 480 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 336952 -960 337176 480 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 342664 -960 342888 480 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 348376 -960 348600 480 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 354088 -960 354312 480 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 359800 -960 360024 480 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 365512 -960 365736 480 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 371224 -960 371448 480 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 376936 -960 377160 480 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 382648 -960 382872 480 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 228424 -960 228648 480 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 388360 -960 388584 480 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 394072 -960 394296 480 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 399784 -960 400008 480 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 405496 -960 405720 480 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 411208 -960 411432 480 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 416920 -960 417144 480 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 422632 -960 422856 480 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 428344 -960 428568 480 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 434056 -960 434280 480 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 439768 -960 439992 480 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 234136 -960 234360 480 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 445480 -960 445704 480 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 451192 -960 451416 480 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 456904 -960 457128 480 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 462616 -960 462840 480 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 468328 -960 468552 480 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 474040 -960 474264 480 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 479752 -960 479976 480 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 485464 -960 485688 480 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 491176 -960 491400 480 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 496888 -960 497112 480 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 239848 -960 240072 480 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 502600 -960 502824 480 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 508312 -960 508536 480 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 514024 -960 514248 480 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 519736 -960 519960 480 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 525448 -960 525672 480 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 531160 -960 531384 480 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 536872 -960 537096 480 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 542584 -960 542808 480 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 548296 -960 548520 480 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 554008 -960 554232 480 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 245560 -960 245784 480 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 559720 -960 559944 480 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 565432 -960 565656 480 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 571144 -960 571368 480 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 576856 -960 577080 480 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 251272 -960 251496 480 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 256984 -960 257208 480 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 262696 -960 262920 480 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 268408 -960 268632 480 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 578760 -960 578984 480 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 580664 -960 580888 480 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 582568 -960 582792 480 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 584472 -960 584696 480 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s -956 -684 -336 597308 4 vdd
port 311 nsew power bidirectional
rlabel metal5 s -956 -684 597020 -64 8 vdd
port 311 nsew power bidirectional
rlabel metal5 s -956 596688 597020 597308 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 596400 -684 597020 597308 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 5418 -1644 6038 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 36138 -1644 36758 517448 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 36138 550512 36758 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 66858 -1644 67478 518408 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 66858 551592 67478 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 97578 -1644 98198 553328 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 97578 573912 98198 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 128298 -1644 128918 507368 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 128298 577636 128918 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 159018 -1644 159638 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 159018 487164 159638 519728 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 159018 563592 159638 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 189738 -1644 190358 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 189738 549192 190358 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 220458 -1644 221078 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 220458 487164 221078 546008 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 220458 572592 221078 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 251178 -1644 251798 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 251178 577632 251798 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 281898 -1644 282518 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 281898 487164 282518 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 312618 -1644 313238 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 312618 487164 313238 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 343338 -1644 343958 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 343338 487164 343958 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 374058 -1644 374678 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 374058 487164 374678 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 404778 -1644 405398 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 404778 487164 405398 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 435498 -1644 436118 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 435498 487164 436118 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 466218 -1644 466838 17452 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 466218 487164 466838 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 496938 -1644 497558 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 527658 -1644 528278 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 558378 -1644 558998 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 589098 -1644 589718 598268 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 3636 597980 4636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 21636 597980 22636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 39636 597980 40636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 57636 189012 58636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 75636 189012 76636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 93636 189012 94636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 111636 189012 112636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 129636 189012 130636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 147636 152116 148636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 165636 152116 166636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 183636 152116 184636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 201636 152116 202636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 219636 152116 220636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 237636 152116 238636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 255636 152116 256636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 273636 152116 274636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 291636 152116 292636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 309636 152116 310636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 327636 152116 328636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 345636 152116 346636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 363636 152116 364636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 381636 189012 382636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 399636 189012 400636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 417636 189012 418636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 435636 189012 436636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 453636 597980 454636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 471636 597980 472636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 489636 597980 490636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 507636 597980 508636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 525636 597980 526636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 543636 597980 544636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 561636 597980 562636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1916 579636 597980 580636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 57636 597980 58636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 75636 597980 76636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 93636 597980 94636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 111636 597980 112636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 129636 597980 130636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 381636 597980 382636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 399636 597980 400636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 417636 597980 418636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 442948 435636 597980 436636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 147636 597980 148636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 165636 597980 166636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 183636 597980 184636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 201636 597980 202636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 219636 597980 220636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 237636 597980 238636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 255636 597980 256636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 273636 597980 274636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 291636 597980 292636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 309636 597980 310636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 327636 597980 328636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 345636 597980 346636 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 479844 363636 597980 364636 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s -1916 -1644 -1296 598268 4 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 -1644 597980 -1024 8 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 597648 597980 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 597360 -1644 597980 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 9138 -1644 9758 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 39858 -1644 40478 527288 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 39858 560472 40478 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 70578 -1644 71198 508448 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 70578 541632 71198 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 101298 -1644 101918 547808 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 101298 568272 101918 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 132018 -1644 132638 507368 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 132018 577636 132638 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 162738 -1644 163358 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 162738 487164 163358 529328 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 162738 573432 163358 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 193458 -1644 194078 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 193458 539352 194078 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 224178 -1644 224798 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 224178 487164 224798 540488 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 224178 566952 224798 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 254898 -1644 255518 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 254898 577632 255518 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 285618 -1644 286238 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 285618 487164 286238 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 316338 -1644 316958 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 316338 487164 316958 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 347058 -1644 347678 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 347058 487164 347678 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 377778 -1644 378398 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 377778 487164 378398 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 408498 -1644 409118 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 408498 487164 409118 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 439218 -1644 439838 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 439218 487164 439838 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 469938 -1644 470558 17452 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 469938 487164 470558 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 500658 -1644 501278 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 531378 -1644 531998 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 562098 -1644 562718 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 592818 -1644 593438 598268 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 10636 597980 11636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 28636 597980 29636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 46636 597980 47636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 64636 189012 65636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 82636 189012 83636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 100636 189012 101636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 118636 189012 119636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 136636 189012 137636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 154636 152116 155636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 172636 152116 173636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 190636 152116 191636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 208636 152116 209636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 226636 152116 227636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 244636 152116 245636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 262636 152116 263636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 280636 152116 281636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 298636 152116 299636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 316636 152116 317636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 334636 152116 335636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 352636 152116 353636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 370636 189012 371636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 388636 189012 389636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 406636 189012 407636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 424636 189012 425636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 442636 189012 443636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 460636 597980 461636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 478636 597980 479636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 496636 597980 497636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 514636 597980 515636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 532636 597980 533636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 550636 597980 551636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 568636 597980 569636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1916 586636 597980 587636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 64636 597980 65636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 82636 597980 83636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 100636 597980 101636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 118636 597980 119636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 136636 597980 137636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 370636 597980 371636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 388636 597980 389636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 406636 597980 407636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 424636 597980 425636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 442948 442636 597980 443636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 154636 597980 155636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 172636 597980 173636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 190636 597980 191636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 208636 597980 209636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 226636 597980 227636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 244636 597980 245636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 262636 597980 263636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 280636 597980 281636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 298636 597980 299636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 316636 597980 317636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 334636 597980 335636 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s 479844 352636 597980 353636 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 11368 -960 11592 480 8 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 13272 -960 13496 480 8 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 15176 -960 15400 480 8 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 22792 -960 23016 480 8 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 87528 -960 87752 480 8 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 93240 -960 93464 480 8 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 98952 -960 99176 480 8 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 104664 -960 104888 480 8 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 110376 -960 110600 480 8 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 116088 -960 116312 480 8 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 121800 -960 122024 480 8 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 127512 -960 127736 480 8 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 133224 -960 133448 480 8 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 138936 -960 139160 480 8 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 30408 -960 30632 480 8 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 144648 -960 144872 480 8 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 150360 -960 150584 480 8 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 156072 -960 156296 480 8 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 161784 -960 162008 480 8 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 167496 -960 167720 480 8 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 173208 -960 173432 480 8 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 178920 -960 179144 480 8 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 184632 -960 184856 480 8 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 190344 -960 190568 480 8 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 196056 -960 196280 480 8 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 38024 -960 38248 480 8 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 201768 -960 201992 480 8 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 207480 -960 207704 480 8 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 45640 -960 45864 480 8 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 53256 -960 53480 480 8 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 58968 -960 59192 480 8 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 64680 -960 64904 480 8 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 70392 -960 70616 480 8 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 76104 -960 76328 480 8 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 81816 -960 82040 480 8 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 17080 -960 17304 480 8 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 24696 -960 24920 480 8 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 89432 -960 89656 480 8 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 95144 -960 95368 480 8 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 100856 -960 101080 480 8 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 106568 -960 106792 480 8 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 112280 -960 112504 480 8 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 117992 -960 118216 480 8 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 123704 -960 123928 480 8 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 129416 -960 129640 480 8 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 135128 -960 135352 480 8 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 140840 -960 141064 480 8 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 32312 -960 32536 480 8 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 146552 -960 146776 480 8 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 152264 -960 152488 480 8 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 157976 -960 158200 480 8 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 163688 -960 163912 480 8 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 169400 -960 169624 480 8 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 175112 -960 175336 480 8 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 180824 -960 181048 480 8 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 186536 -960 186760 480 8 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 192248 -960 192472 480 8 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 197960 -960 198184 480 8 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 39928 -960 40152 480 8 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 203672 -960 203896 480 8 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 209384 -960 209608 480 8 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 47544 -960 47768 480 8 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 55160 -960 55384 480 8 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 60872 -960 61096 480 8 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 66584 -960 66808 480 8 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 72296 -960 72520 480 8 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 78008 -960 78232 480 8 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 83720 -960 83944 480 8 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 26600 -960 26824 480 8 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 91336 -960 91560 480 8 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 97048 -960 97272 480 8 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 102760 -960 102984 480 8 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 108472 -960 108696 480 8 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 114184 -960 114408 480 8 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 119896 -960 120120 480 8 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 125608 -960 125832 480 8 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 131320 -960 131544 480 8 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 137032 -960 137256 480 8 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 142744 -960 142968 480 8 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 34216 -960 34440 480 8 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 148456 -960 148680 480 8 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 154168 -960 154392 480 8 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 159880 -960 160104 480 8 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 165592 -960 165816 480 8 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 171304 -960 171528 480 8 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 177016 -960 177240 480 8 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 182728 -960 182952 480 8 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 188440 -960 188664 480 8 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 194152 -960 194376 480 8 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 199864 -960 200088 480 8 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 41832 -960 42056 480 8 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 205576 -960 205800 480 8 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 211288 -960 211512 480 8 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 49448 -960 49672 480 8 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 57064 -960 57288 480 8 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 62776 -960 63000 480 8 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 68488 -960 68712 480 8 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 74200 -960 74424 480 8 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 79912 -960 80136 480 8 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 85624 -960 85848 480 8 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 28504 -960 28728 480 8 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 36120 -960 36344 480 8 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 43736 -960 43960 480 8 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 51352 -960 51576 480 8 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 18984 -960 19208 480 8 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 20888 -960 21112 480 8 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 596040 596040
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 19900960
string GDS_FILE /home/oe23ranan/gf_analog/openlane/user_project_wrapper/runs/23_12_07_23_57/results/signoff/user_project_wrapper.magic.gds
string GDS_START 9713058
<< end >>

