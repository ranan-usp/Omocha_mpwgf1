* NGSPICE file created from dac.ext - technology: gf180mcuD

.subckt XM1_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 D S 0.038197f
C2 G S 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM4_bs G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# S 0.021189f
C1 D G 0.002389f
C2 D S 0.045397f
C3 S G 0.002389f
C4 D w_n319_n356# 0.019807f
C5 w_n319_n356# G 0.186402f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMs1_bs G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 D S 0.038197f
C2 G S 0.002868f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365275f
.ends

.subckt bs_cap I1_1_1_R0_BOT I1_1_1_R0_TOP VSUBS
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.339999u c_length=12.339999u
C0 I1_1_1_R0_BOT I1_1_1_R0_TOP 2.24198f
C1 I1_1_1_R0_TOP VSUBS 2.33555f
C2 I1_1_1_R0_BOT VSUBS 2.1391f
.ends

.subckt XM3_bs G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# S 0.021189f
C1 D G 0.002389f
C2 D S 0.045397f
C3 S G 0.002389f
C4 D w_n319_n356# 0.019807f
C5 w_n319_n356# G 0.186402f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XM1_bs_inv G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 D S 0.038197f
C2 G S 0.002868f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365365f
.ends

.subckt XM2_bs_inv G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# S 0.019807f
C1 D G 0.002389f
C2 D S 0.045397f
C3 S G 0.002389f
C4 D w_n319_n356# 0.019807f
C5 w_n319_n356# G 0.186609f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48751f
.ends

.subckt bs_inv inv_in inv_out vdd vss
XXM1_bs_inv_0 inv_in inv_out vss vss XM1_bs_inv
XXM2_bs_inv_0 inv_in inv_out vdd vdd vss XM2_bs_inv
C0 vdd inv_out 0.092565f
C1 inv_in inv_out 0.075645f
C2 inv_out vss 0.04895f
C3 inv_in vdd 0.07083f
C4 vdd vss 0.043239f
C5 inv_in vss 0.037258f
C6 vdd 0 1.650725f
C7 inv_out 0 0.392313f
C8 vss 0 0.277512f
C9 inv_in 0 0.605506f
.ends

.subckt XMs_bs G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D S 0.038197f
C2 D G 0.002868f
C3 D a_n302_n324# 0.061336f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361785f
.ends

.subckt XM2_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 D G 0.002868f
C2 S G 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XMs2_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 D G 0.002868f
C2 S G 0.002868f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.068446f
C5 G a_n302_n324# 0.365186f
.ends

.subckt bootstrapped_sw vg vs vdd en enb bs_in bs_out vbsl vss vbsh
XXM1_bs_0 vg vbsl vss vss bs_in XM1_bs
XXM4_bs_0 vg vdd vbsh vbsh vss XM4_bs
XXMs1_bs_0 vdd vs vss vg XMs1_bs
Xbs_cap_0 vbsl vbsh vss bs_cap
Xbs_cap_1 vbsl vbsh vss bs_cap
XXM3_bs_0 enb vg vbsh vbsh vss XM3_bs
Xbs_cap_2 vbsl vbsh vss bs_cap
Xbs_cap_4 vbsl vbsh vss bs_cap
Xbs_cap_3 vbsl vbsh vss bs_cap
Xbs_inv_0 en enb vdd vss bs_inv
XXMs_bs_0 vg bs_out vss bs_in XMs_bs
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 enb vss vss vss vs XMs2_bs
C0 vbsh bs_in 0.013047f
C1 vs enb 0.00173f
C2 vs vg 0.006382f
C3 vbsh vbsl 3.67197f
C4 vdd enb 0.426791f
C5 vg enb 0.693229f
C6 vg vdd 0.490821f
C7 vg bs_in 0.079028f
C8 vbsl enb 0.01529f
C9 vbsl vdd 0.002507f
C10 vbsl vg 0.040934f
C11 vbsl bs_in 0.272985f
C12 bs_out vbsh 0.119559f
C13 en enb 0.018916f
C14 en vdd 0.086628f
C15 en vg 0.002156f
C16 bs_out enb 0.001285f
C17 bs_out vdd 0.008497f
C18 bs_out vg 0.066304f
C19 vbsh enb 0.0922f
C20 bs_out vbsl 0.05557f
C21 vbsh vdd 0.205818f
C22 vbsh vg 0.287508f
C23 enb vss 1.704268f
C24 bs_out vss 0.895635f
C25 bs_in vss 0.378553f
C26 vg vss 1.570874f
C27 vdd vss 3.559775f
C28 en vss 0.896531f
C29 vbsh vss 12.08863f
C30 vbsl vss 10.320489f
C31 vs vss 0.04326f
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VDD I 0.074838f
C1 VDD VSS 0.029045f
C2 ZN I 0.58604f
C3 VSS ZN 0.180794f
C4 VDD VNW 0.082022f
C5 ZN VNW 0.023676f
C6 VSS I 0.091531f
C7 VDD ZN 0.271625f
C8 I VNW 0.285482f
C9 VSS VNW 0.006277f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu inv$1_1/I inv$1_8/I inv$1_7/ZN inv$1_1/ZN inv$1_3/I inv$1_5/I
+ inv$1_7/I inv$1_9/ZN inv$1_9/I inv$1_3/ZN inv$1_6/ZN vdd inv$1_0/ZN inv$1_0/I inv$1_4/ZN
+ inv$1_2/I inv$1_10/I inv$1_4/I inv$1_10/ZN inv$1_8/ZN vss inv$1_6/I inv$1_2/ZN inv$1_5/ZN
Xinv$1_10 vss inv$1_10/ZN inv$1_10/I vdd vdd inv$1_10/VPW vss inv$1
Xinv$1_0 vss inv$1_0/ZN inv$1_0/I vdd vdd inv$1_0/VPW vss inv$1
Xinv$1_1 vss inv$1_1/ZN inv$1_1/I vdd vdd inv$1_1/VPW vss inv$1
Xinv$1_2 vss inv$1_2/ZN inv$1_2/I vdd vdd inv$1_2/VPW vss inv$1
Xinv$1_3 vss inv$1_3/ZN inv$1_3/I vdd vdd inv$1_3/VPW vss inv$1
Xinv$1_4 vss inv$1_4/ZN inv$1_4/I vdd vdd inv$1_4/VPW vss inv$1
Xinv$1_5 vss inv$1_5/ZN inv$1_5/I vdd vdd inv$1_5/VPW vss inv$1
Xinv$1_6 vss inv$1_6/ZN inv$1_6/I vdd vdd inv$1_6/VPW vss inv$1
Xinv$1_7 vss inv$1_7/ZN inv$1_7/I vdd vdd inv$1_7/VPW vss inv$1
Xinv$1_8 vss inv$1_8/ZN inv$1_8/I vdd vdd inv$1_8/VPW vss inv$1
Xinv$1_9 vss inv$1_9/ZN inv$1_9/I vdd vdd inv$1_9/VPW vss inv$1
C0 inv$1_5/ZN vdd 0.159176f
C1 inv$1_9/ZN inv$1_10/I 0.002086f
C2 inv$1_10/ZN inv$1_9/I 0.028928f
C3 inv$1_7/I inv$1_6/I 0.084161f
C4 inv$1_10/I vss 0.166388f
C5 inv$1_1/ZN vdd 0.159176f
C6 inv$1_5/ZN inv$1_5/I 0.029333f
C7 inv$1_5/ZN inv$1_6/I 0.002086f
C8 inv$1_8/I inv$1_7/ZN 0.002086f
C9 inv$1_4/I vss 0.166388f
C10 inv$1_3/I inv$1_1/ZN 0.028928f
C11 inv$1_7/ZN vss 0.003326f
C12 inv$1_8/ZN inv$1_7/ZN 0.080571f
C13 inv$1_0/ZN inv$1_3/ZN 0.080571f
C14 inv$1_4/ZN vss 0.003326f
C15 inv$1_2/ZN inv$1_10/ZN 0.080571f
C16 inv$1_6/ZN inv$1_7/ZN 0.080571f
C17 inv$1_7/I inv$1_8/I 0.084161f
C18 inv$1_3/I vdd 0.019437f
C19 inv$1_7/I vss 0.166388f
C20 inv$1_8/ZN inv$1_7/I 0.028928f
C21 inv$1_5/I vdd 0.019437f
C22 inv$1_6/I vdd 0.019437f
C23 inv$1_2/I inv$1_10/I 0.084161f
C24 inv$1_5/ZN vss 0.003326f
C25 inv$1_7/I inv$1_6/ZN 0.002086f
C26 inv$1_0/I vdd 0.026972f
C27 inv$1_5/I inv$1_6/I 0.084161f
C28 inv$1_5/ZN inv$1_6/ZN 0.080571f
C29 inv$1_3/I inv$1_0/I 0.08416f
C30 inv$1_1/ZN vss 0.003326f
C31 inv$1_9/ZN vdd 0.159176f
C32 inv$1_8/I vdd 0.019437f
C33 inv$1_9/I inv$1_10/I 0.084161f
C34 vss vdd 0.009518f
C35 inv$1_8/ZN vdd 0.159176f
C36 inv$1_3/I vss 0.166388f
C37 inv$1_6/ZN vdd 0.159176f
C38 inv$1_5/I vss 0.166388f
C39 inv$1_6/I vss 0.166388f
C40 inv$1_10/ZN inv$1_10/I 0.029333f
C41 inv$1_2/ZN inv$1_10/I 0.028928f
C42 inv$1_0/I vss 0.170492f
C43 inv$1_5/I inv$1_6/ZN 0.028928f
C44 inv$1_6/I inv$1_6/ZN 0.029333f
C45 inv$1_9/ZN inv$1_8/I 0.028928f
C46 inv$1_2/I vdd 0.035575f
C47 inv$1_9/ZN vss 0.003326f
C48 inv$1_8/ZN inv$1_9/ZN 0.080571f
C49 inv$1_1/I inv$1_3/ZN 0.002086f
C50 inv$1_0/ZN vdd 0.184001f
C51 inv$1_8/I vss 0.166388f
C52 inv$1_8/ZN inv$1_8/I 0.029333f
C53 inv$1_8/ZN vss 0.003326f
C54 inv$1_3/I inv$1_0/ZN 0.002086f
C55 inv$1_6/ZN vss 0.003326f
C56 inv$1_0/ZN inv$1_0/I 0.029333f
C57 inv$1_9/I vdd 0.019437f
C58 inv$1_4/I inv$1_1/I 0.084161f
C59 inv$1_10/ZN vdd 0.159176f
C60 inv$1_2/I vss 0.164788f
C61 inv$1_1/I inv$1_4/ZN 0.028928f
C62 inv$1_2/ZN vdd 0.174722f
C63 inv$1_0/ZN vss 0.005399f
C64 inv$1_9/ZN inv$1_9/I 0.029333f
C65 inv$1_8/I inv$1_9/I 0.084161f
C66 inv$1_3/ZN inv$1_1/ZN 0.080571f
C67 inv$1_4/I inv$1_4/ZN 0.029333f
C68 inv$1_9/I vss 0.166388f
C69 inv$1_8/ZN inv$1_9/I 0.002086f
C70 inv$1_1/I inv$1_1/ZN 0.029333f
C71 inv$1_10/ZN inv$1_9/ZN 0.080571f
C72 inv$1_3/ZN vdd 0.159176f
C73 inv$1_7/I inv$1_7/ZN 0.029333f
C74 inv$1_10/ZN vss 0.003326f
C75 inv$1_5/ZN inv$1_4/I 0.028928f
C76 inv$1_3/I inv$1_3/ZN 0.029333f
C77 inv$1_2/ZN vss 0.005014f
C78 inv$1_1/I vdd 0.019437f
C79 inv$1_5/ZN inv$1_4/ZN 0.080571f
C80 inv$1_3/I inv$1_1/I 0.084161f
C81 inv$1_4/I inv$1_1/ZN 0.002086f
C82 inv$1_3/ZN inv$1_0/I 0.028928f
C83 inv$1_1/ZN inv$1_4/ZN 0.080571f
C84 inv$1_10/I vdd 0.019437f
C85 inv$1_4/I vdd 0.019437f
C86 inv$1_7/ZN vdd 0.159176f
C87 inv$1_10/ZN inv$1_2/I 0.002086f
C88 inv$1_4/ZN vdd 0.159176f
C89 inv$1_2/ZN inv$1_2/I 0.029333f
C90 inv$1_3/ZN vss 0.003326f
C91 inv$1_5/I inv$1_4/I 0.084161f
C92 inv$1_6/I inv$1_7/ZN 0.028928f
C93 inv$1_7/I vdd 0.019437f
C94 inv$1_5/I inv$1_4/ZN 0.002086f
C95 inv$1_1/I vss 0.166388f
C96 inv$1_9/ZN 0 0.131999f
C97 inv$1_9/I 0 0.64919f
C98 inv$1_8/ZN 0 0.131999f
C99 inv$1_8/I 0 0.64919f
C100 inv$1_7/ZN 0 0.131999f
C101 inv$1_7/I 0 0.64919f
C102 inv$1_6/ZN 0 0.131999f
C103 inv$1_6/I 0 0.64919f
C104 inv$1_5/ZN 0 0.131999f
C105 inv$1_5/I 0 0.64919f
C106 inv$1_4/ZN 0 0.131999f
C107 inv$1_4/I 0 0.64919f
C108 inv$1_3/ZN 0 0.131999f
C109 inv$1_3/I 0 0.64919f
C110 vss 0 3.02573f
C111 inv$1_2/ZN 0 0.206166f
C112 vdd 0 16.013325f
C113 inv$1_2/I 0 0.750024f
C114 inv$1_1/ZN 0 0.131999f
C115 inv$1_1/I 0 0.64919f
C116 inv$1_0/ZN 0 0.209411f
C117 inv$1_0/I 0 0.731246f
C118 inv$1_10/ZN 0 0.131999f
C119 inv$1_10/I 0 0.64919f
.ends

.subckt dac vdd vss dac_in dac_out dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9
+ ctl10 sample
Xbootstrapped_sw_0 bootstrapped_sw_0/vg bootstrapped_sw_0/vs vdd sample bootstrapped_sw_0/enb
+ dac_in dac_out bootstrapped_sw_0/vbsl vss bootstrapped_sw_0/vbsh bootstrapped_sw
Xinv_renketu_0 ctl2 ctl7 carray_0/n6 carray_0/n2 ctl1 ctl4 ctl6 carray_0/n8 ctl8 carray_0/n1
+ carray_0/n5 vdd carray_0/ndum dum carray_0/n3 ctl10 ctl9 ctl3 carray_0/n9 carray_0/n7
+ vss ctl5 carray_0/n0 carray_0/n4 inv_renketu
C0 carray_0/n4 carray_0/n8 2.84323f
C1 carray_0/n8 dac_out 0.420151p
C2 carray_0/n1 carray_0/n3 0.145048f
C3 carray_0/n9 carray_0/n4 3.740573f
C4 vdd carray_0/n1 0.002151f
C5 carray_0/n9 dac_out 0.846161p
C6 carray_0/n4 carray_0/n1 0.142475f
C7 carray_0/n9 carray_0/n8 87.43918f
C8 dac_out carray_0/n1 3.367623f
C9 ctl10 ctl9 0.104537f
C10 carray_0/n6 carray_0/n3 0.336612f
C11 carray_0/n8 carray_0/n1 0.28587f
C12 ctl5 ctl6 0.104537f
C13 vdd carray_0/n6 0.002151f
C14 carray_0/n9 carray_0/n1 0.350042f
C15 ctl9 ctl8 0.104537f
C16 ctl3 ctl4 0.104537f
C17 carray_0/ndum carray_0/n3 0.025424f
C18 carray_0/n4 carray_0/n6 0.614078f
C19 carray_0/n5 carray_0/n3 0.346757f
C20 carray_0/n0 carray_0/n3 0.051666f
C21 carray_0/ndum vdd 0.004405f
C22 vdd carray_0/n0 0.002151f
C23 carray_0/n5 vdd 0.002151f
C24 dac_out carray_0/n6 0.105055p
C25 ctl3 ctl2 0.104537f
C26 carray_0/n2 carray_0/n7 0.485355f
C27 carray_0/n8 carray_0/n6 11.2161f
C28 carray_0/ndum carray_0/n4 0.025424f
C29 carray_0/n0 carray_0/n4 0.040502f
C30 carray_0/n5 carray_0/n4 27.828503f
C31 carray_0/ndum dac_out 1.640173f
C32 carray_0/n0 dac_out 1.750611f
C33 carray_0/n5 dac_out 52.565514f
C34 carray_0/n9 carray_0/n6 14.716789f
C35 carray_0/ndum carray_0/n8 0.097254f
C36 carray_0/n0 carray_0/n8 0.097254f
C37 carray_0/n5 carray_0/n8 5.60732f
C38 carray_0/n1 carray_0/n6 0.142211f
C39 carray_0/ndum carray_0/n9 0.127951f
C40 carray_0/n9 carray_0/n0 0.521489f
C41 carray_0/n5 carray_0/n9 7.399346f
C42 carray_0/ndum carray_0/n1 8.498201f
C43 carray_0/n0 carray_0/n1 8.476914f
C44 carray_0/n5 carray_0/n1 0.142354f
C45 dac_out bootstrapped_sw_0/vbsh 0.254082f
C46 carray_0/ndum carray_0/n6 0.025424f
C47 carray_0/n0 carray_0/n6 0.025424f
C48 carray_0/n5 carray_0/n6 28.925901f
C49 carray_0/n2 carray_0/n3 23.177217f
C50 carray_0/n7 carray_0/n3 0.891504f
C51 vdd carray_0/n2 0.002151f
C52 vdd carray_0/n7 0.002151f
C53 ctl7 ctl6 0.104537f
C54 carray_0/n5 carray_0/ndum 0.025424f
C55 carray_0/n5 carray_0/n0 0.025424f
C56 carray_0/n4 carray_0/n2 0.213209f
C57 carray_0/n4 carray_0/n7 1.70387f
C58 carray_0/n2 dac_out 6.640605f
C59 dac_out carray_0/n7 0.210031p
C60 ctl5 ctl4 0.104537f
C61 carray_0/n8 carray_0/n2 0.770227f
C62 carray_0/n8 carray_0/n7 50.51461f
C63 carray_0/n9 carray_0/n2 0.996681f
C64 carray_0/n9 carray_0/n7 29.516087f
C65 sample carray_0/ndum 0.045492f
C66 carray_0/n2 carray_0/n1 16.941952f
C67 carray_0/n1 carray_0/n7 0.212822f
C68 ctl1 ctl2 0.104537f
C69 ctl1 dum 0.104537f
C70 carray_0/n2 carray_0/n6 0.20799f
C71 carray_0/n7 carray_0/n6 34.662605f
C72 vdd carray_0/n3 0.002151f
C73 carray_0/n4 carray_0/n3 26.229403f
C74 carray_0/ndum carray_0/n2 0.041162f
C75 carray_0/ndum carray_0/n7 0.06073f
C76 carray_0/n0 carray_0/n2 0.099314f
C77 carray_0/n5 carray_0/n2 0.208112f
C78 vdd carray_0/n4 0.002151f
C79 carray_0/n0 carray_0/n7 0.06073f
C80 carray_0/n5 carray_0/n7 3.36878f
C81 dac_out carray_0/n3 13.201303f
C82 carray_0/n8 carray_0/n3 1.46111f
C83 vdd carray_0/n8 0.002151f
C84 dac_out bootstrapped_sw_0/vbsl 0.193675f
C85 carray_0/n4 dac_out 26.32268f
C86 carray_0/n9 carray_0/n3 1.911224f
C87 ctl8 ctl7 0.104537f
C88 carray_0/n9 vdd 0.002151f
C89 ctl8 vss 0.916847f
C90 ctl7 vss 0.916847f
C91 ctl6 vss 0.916847f
C92 ctl5 vss 0.916847f
C93 ctl4 vss 0.916847f
C94 ctl3 vss 0.916847f
C95 ctl1 vss 0.916847f
C96 carray_0/n0 vss 17.633558f
C97 vdd vss 19.890364f
C98 ctl10 vss 1.146163f
C99 ctl2 vss 0.916847f
C100 carray_0/ndum vss 14.881693f
C101 dum vss 1.125528f
C102 ctl9 vss 0.916847f
C103 carray_0/n4 vss 39.983223f
C104 carray_0/n5 vss 48.006485f
C105 carray_0/n9 vss 14.963586f
C106 dac_out vss -0.683691p
C107 carray_0/n8 vss 40.580837f
C108 carray_0/n7 vss 56.915478f
C109 carray_0/n6 vss 53.64827f
C110 carray_0/n2 vss 30.783176f
C111 carray_0/n1 vss 17.779491f
C112 carray_0/n3 vss 34.26559f
C113 bootstrapped_sw_0/enb vss 1.50362f
C114 dac_in vss 0.363227f
C115 bootstrapped_sw_0/vg vss 1.495112f
C116 sample vss 21.11657f
C117 bootstrapped_sw_0/vbsh vss 12.07361f
C118 bootstrapped_sw_0/vbsl vss 10.152523f
C119 bootstrapped_sw_0/vs vss 0.054281f
.ends

