* NGSPICE file created from sarlogic.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW a_36_472# a_572_375# a_124_375#
+ a_484_472#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 a_36_472# a_484_472# 0.013276f
C1 a_124_375# VNW 0.180172f
C2 a_572_375# VDD 0.129266f
C3 VSS a_484_472# 0.148682f
C4 a_484_472# VNW 0.024396f
C5 a_36_472# VDD 0.093681f
C6 a_572_375# VSS 0.082563f
C7 VDD VSS 0.013184f
C8 a_124_375# a_484_472# 0.086742f
C9 a_572_375# VNW 0.18122f
C10 a_36_472# VSS 0.151218f
C11 VDD VNW 0.11314f
C12 a_124_375# a_572_375# 0.012222f
C13 a_36_472# VNW 0.025611f
C14 a_124_375# VDD 0.12673f
C15 VSS VNW 0.008822f
C16 a_124_375# a_36_472# 0.285629f
C17 a_572_375# a_484_472# 0.285629f
C18 a_124_375# VSS 0.136476f
C19 VDD a_484_472# 0.179463f
C20 VSS VPW 0.360066f
C21 VDD VPW 0.286281f
C22 VNW VPW 1.65967f
C23 a_484_472# VPW 0.345058f
C24 a_36_472# VPW 0.404746f
C25 a_572_375# VPW 0.232991f
C26 a_124_375# VPW 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VNW VPW
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 VNW I 0.027206f
C1 I VDD 0.017439f
C2 I VSS 0.031625f
C3 VNW VDD 0.048519f
C4 VNW VSS 0.007461f
C5 VDD VSS 0.009725f
C6 VSS VPW 0.12617f
C7 VDD VPW 0.087026f
C8 I VPW 0.139667f
C9 VNW VPW 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW a_224_472#
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 VNW A2 0.128798f
C1 a_224_472# VDD 0.013964f
C2 ZN VNW 0.019783f
C3 VDD VSS 0.023219f
C4 a_224_472# A2 0.008979f
C5 VNW A1 0.136915f
C6 a_224_472# ZN 0.023693f
C7 VDD A2 0.255318f
C8 VDD ZN 0.117921f
C9 VSS A2 0.043352f
C10 ZN VSS 0.08687f
C11 VDD A1 0.028041f
C12 ZN A2 0.378409f
C13 VSS A1 0.168633f
C14 A2 A1 0.037814f
C15 ZN A1 0.579732f
C16 VDD VNW 0.093678f
C17 VSS VNW 0.010571f
C18 VSS VPW 0.331491f
C19 ZN VPW 0.058886f
C20 VDD VPW 0.218051f
C21 A1 VPW 0.331856f
C22 A2 VPW 0.334514f
C23 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VNW VPW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_1456_156#
+ a_1288_156# a_2248_156# a_2560_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VPW nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 a_2248_156# RN 0.094336f
C1 a_36_151# a_448_472# 0.536965f
C2 a_2665_112# VNW 0.354715f
C3 a_2560_156# VDD 0.00217f
C4 a_36_151# RN 0.080102f
C5 a_2665_112# VSS 0.184997f
C6 a_448_472# CLK 0.002757f
C7 a_448_472# a_1308_423# 0.882105f
C8 a_1204_472# a_448_472# 0.008996f
C9 a_1308_423# RN 0.079294f
C10 a_796_472# D 0.082858f
C11 VNW VSS 0.010602f
C12 VDD D 0.009367f
C13 a_1000_472# VNW 0.241357f
C14 a_1000_472# VSS 0.04356f
C15 a_1204_472# RN 0.021039f
C16 a_2665_112# a_2248_156# 0.633318f
C17 a_2248_156# VNW 0.212431f
C18 a_2665_112# a_36_151# 0.019043f
C19 a_2248_156# VSS 0.030473f
C20 a_1000_472# a_2248_156# 0.001232f
C21 a_36_151# VNW 1.28833f
C22 a_448_472# a_1456_156# 0.00227f
C23 a_36_151# VSS 0.291264f
C24 a_2665_112# Q 0.109436f
C25 a_448_472# a_796_472# 0.401636f
C26 a_448_472# VDD 0.456269f
C27 a_36_151# a_1000_472# 0.08126f
C28 a_1308_423# VNW 0.149014f
C29 VNW CLK 0.137037f
C30 a_1308_423# VSS 0.013866f
C31 VNW Q 0.034443f
C32 CLK VSS 0.021952f
C33 VDD RN 0.034984f
C34 a_1204_472# VNW 0.016269f
C35 a_1000_472# a_1308_423# 0.934191f
C36 VSS Q 0.113401f
C37 a_36_151# a_2248_156# 0.042802f
C38 a_1000_472# a_1204_472# 0.66083f
C39 a_2248_156# a_1308_423# 0.056721f
C40 a_2560_156# a_448_472# 0.277491f
C41 a_2248_156# Q 0.014355f
C42 a_36_151# CLK 0.669598f
C43 a_36_151# a_1308_423# 0.05539f
C44 a_2560_156# RN 0.038779f
C45 a_2665_112# VDD 0.102046f
C46 a_448_472# D 0.328788f
C47 a_36_151# a_1204_472# 0.006996f
C48 a_796_472# VNW 0.010232f
C49 a_3041_156# RN 0.01068f
C50 VNW VDD 0.503557f
C51 a_1456_156# VSS 0.001901f
C52 a_796_472# VSS 0.05215f
C53 VDD VSS 0.01338f
C54 a_1000_472# VDD 0.119211f
C55 a_1204_472# a_1308_423# 0.026665f
C56 a_1000_472# a_796_472# 0.048436f
C57 a_2560_156# a_2665_112# 0.116059f
C58 a_2248_156# VDD 1.11667f
C59 a_1288_156# a_448_472# 0.002067f
C60 a_2560_156# VNW 0.020165f
C61 a_2665_112# a_3041_156# 0.001774f
C62 a_36_151# a_796_472# 0.011851f
C63 a_36_151# VDD 0.417088f
C64 a_2560_156# VSS 0.128503f
C65 a_448_472# RN 0.078731f
C66 a_1308_423# VDD 0.094185f
C67 CLK VDD 0.02303f
C68 VNW D 0.128231f
C69 VDD Q 0.149344f
C70 D VSS 0.064618f
C71 a_1204_472# VDD 0.282626f
C72 a_2560_156# a_2248_156# 0.119687f
C73 a_2560_156# a_36_151# 0.003674f
C74 a_2665_112# a_448_472# 0.020455f
C75 a_36_151# D 0.094113f
C76 a_1288_156# VSS 0.001702f
C77 a_2665_112# RN 0.336469f
C78 a_448_472# VNW 0.341284f
C79 a_448_472# VSS 1.20207f
C80 a_1000_472# a_448_472# 0.361958f
C81 VNW RN 0.329494f
C82 RN VSS 0.441968f
C83 a_1000_472# RN 0.0832f
C84 a_2248_156# a_448_472# 0.510371f
C85 Q VPW 0.114762f
C86 VSS VPW 1.26186f
C87 RN VPW 1.36673f
C88 D VPW 0.253406f
C89 VDD VPW 0.79945f
C90 CLK VPW 0.291241f
C91 VNW VPW 6.1377f
C92 a_2560_156# VPW 0.016968f
C93 a_2665_112# VPW 0.62251f
C94 a_2248_156# VPW 0.371662f
C95 a_1204_472# VPW 0.012971f
C96 a_1000_472# VPW 0.291735f
C97 a_796_472# VPW 0.023206f
C98 a_1308_423# VPW 0.279043f
C99 a_448_472# VPW 0.684413f
C100 a_36_151# VPW 1.43589f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VNW VPW a_36_68# a_244_472#
+ a_692_472#
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 VSS B2 0.025295f
C1 VSS A2 0.087422f
C2 a_244_472# B2 0.002003f
C3 VNW B1 0.125926f
C4 ZN VNW 0.010694f
C5 VSS B1 0.025138f
C6 VSS ZN 0.085273f
C7 A1 VNW 0.115376f
C8 VDD VNW 0.139306f
C9 a_244_472# B1 0.003598f
C10 a_36_68# VNW 0.040298f
C11 B2 B1 0.036483f
C12 A2 ZN 0.390894f
C13 VSS A1 0.084232f
C14 VSS VDD 0.011512f
C15 VSS a_36_68# 0.392965f
C16 VDD a_244_472# 0.00636f
C17 a_244_472# a_36_68# 0.027448f
C18 A2 A1 0.038725f
C19 a_36_68# B2 0.369561f
C20 VDD B2 0.246452f
C21 A2 a_36_68# 0.340509f
C22 A2 VDD 0.019572f
C23 ZN a_692_472# 0.011665f
C24 ZN B1 0.079f
C25 VDD a_692_472# 0.004194f
C26 A1 B1 0.163724f
C27 a_692_472# a_36_68# 0.015646f
C28 ZN A1 0.430191f
C29 a_36_68# B1 0.437534f
C30 VDD B1 0.014643f
C31 ZN a_36_68# 0.419486f
C32 ZN VDD 0.004634f
C33 VSS VNW 0.010714f
C34 A1 a_36_68# 0.160084f
C35 VDD A1 0.014671f
C36 VDD a_36_68# 0.787847f
C37 VNW B2 0.133721f
C38 A2 VNW 0.125671f
C39 VSS VPW 0.383233f
C40 ZN VPW 0.012598f
C41 VDD VPW 0.318857f
C42 A2 VPW 0.2826f
C43 A1 VPW 0.258579f
C44 B1 VPW 0.257485f
C45 B2 VPW 0.309037f
C46 VNW VPW 2.00777f
C47 a_36_68# VPW 0.150048f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW a_49_472#
+ a_665_69# a_257_69#
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
C0 VSS a_665_69# 0.003829f
C1 B1 a_257_69# 0.003901f
C2 VDD ZN 0.004108f
C3 A2 A1 0.392541f
C4 a_665_69# A2 0.006702f
C5 ZN a_49_472# 0.239204f
C6 VNW ZN 0.017894f
C7 a_665_69# A1 0.002008f
C8 VSS VDD 0.00787f
C9 VSS a_49_472# 0.02154f
C10 VSS VNW 0.011011f
C11 B2 VDD 0.026097f
C12 B2 a_49_472# 0.151151f
C13 B2 VNW 0.129409f
C14 A2 VDD 0.013575f
C15 VDD A1 0.013859f
C16 A2 a_49_472# 0.075759f
C17 VNW A2 0.131727f
C18 A1 a_49_472# 0.021757f
C19 VSS a_257_69# 0.00576f
C20 VNW A1 0.10965f
C21 B2 a_257_69# 0.003563f
C22 B1 ZN 0.367665f
C23 B1 VSS 0.095385f
C24 VDD a_49_472# 0.887006f
C25 VNW VDD 0.112326f
C26 VNW a_49_472# 0.026629f
C27 B1 B2 0.18297f
C28 B1 A1 0.041046f
C29 VSS ZN 0.071892f
C30 B1 VDD 0.017923f
C31 B2 ZN 0.001886f
C32 B1 a_49_472# 0.069833f
C33 B1 VNW 0.109456f
C34 A2 ZN 0.102518f
C35 VSS B2 0.06757f
C36 ZN A1 0.447732f
C37 a_665_69# ZN 0.001059f
C38 VSS A2 0.150463f
C39 VSS A1 0.087393f
C40 VSS VPW 0.39457f
C41 ZN VPW 0.021794f
C42 VDD VPW 0.243433f
C43 A2 VPW 0.322629f
C44 A1 VPW 0.250967f
C45 B1 VPW 0.261124f
C46 B2 VPW 0.322244f
C47 VNW VPW 1.83372f
C48 a_49_472# VPW 0.054843f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VNW VPW a_36_160#
X0 Z a_36_160# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VPW nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 a_36_160# I 0.545454f
C1 a_36_160# VNW 0.170864f
C2 I VNW 0.2276f
C3 VDD Z 0.128274f
C4 VSS VDD 0.009574f
C5 a_36_160# VDD 0.2736f
C6 I VDD 0.02612f
C7 VDD VNW 0.087464f
C8 VSS Z 0.146199f
C9 a_36_160# Z 0.281838f
C10 I Z 0.041707f
C11 VSS a_36_160# 0.074156f
C12 Z VNW 0.030347f
C13 VSS I 0.12329f
C14 VSS VNW 0.009324f
C15 VSS VPW 0.28275f
C16 Z VPW 0.10469f
C17 VDD VPW 0.178615f
C18 I VPW 0.323491f
C19 VNW VPW 1.31158f
C20 a_36_160# VPW 0.386641f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD I 0.157124f
C1 ZN VSS 0.077008f
C2 VDD ZN 0.098026f
C3 ZN I 0.47009f
C4 VNW VSS 0.011085f
C5 VNW VDD 0.076212f
C6 VNW I 0.135368f
C7 VNW ZN 0.031181f
C8 VDD VSS 0.025441f
C9 VSS I 0.058937f
C10 VSS VPW 0.242183f
C11 ZN VPW 0.095505f
C12 VDD VPW 0.182097f
C13 I VPW 0.355642f
C14 VNW VPW 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 ZN VSS 0.115297f
C1 VDD I 0.041847f
C2 VDD ZN 0.137375f
C3 ZN I 0.262199f
C4 VNW VSS 0.011339f
C5 VNW VDD 0.076257f
C6 VNW I 0.137757f
C7 VNW ZN 0.022202f
C8 VDD VSS 0.025626f
C9 VSS I 0.0533f
C10 VSS VPW 0.2316f
C11 ZN VPW 0.113404f
C12 VDD VPW 0.181139f
C13 I VPW 0.341982f
C14 VNW VPW 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW a_36_472# a_124_375#
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 a_124_375# VNW 0.179924f
C1 VDD VSS 0.006592f
C2 a_124_375# VDD 0.126034f
C3 VNW VDD 0.061035f
C4 a_36_472# VSS 0.150876f
C5 a_36_472# a_124_375# 0.285629f
C6 a_36_472# VNW 0.025989f
C7 a_36_472# VDD 0.093681f
C8 a_124_375# VSS 0.082879f
C9 VNW VSS 0.004411f
C10 VSS VPW 0.218985f
C11 VDD VPW 0.182777f
C12 VNW VPW 0.96348f
C13 a_36_472# VPW 0.417394f
C14 a_124_375# VPW 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VNW VPW a_224_472#
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 a_224_472# I 0.796069f
C1 a_224_472# VNW 1.14633f
C2 VDD Z 0.819024f
C3 I VNW 0.55539f
C4 VSS VDD 0.031131f
C5 a_224_472# VDD 0.74621f
C6 I VDD 0.1311f
C7 VDD VNW 0.305516f
C8 VSS Z 0.70427f
C9 a_224_472# Z 2.29481f
C10 I Z 0.001907f
C11 VSS a_224_472# 0.659695f
C12 Z VNW 0.038011f
C13 VSS I 0.158668f
C14 VSS VNW 0.01282f
C15 VSS VPW 0.910368f
C16 Z VPW 0.18914f
C17 VDD VPW 0.724491f
C18 I VPW 1.16773f
C19 VNW VPW 4.79254f
C20 a_224_472# VPW 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW a_36_472# a_244_68#
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
C0 B VDD 0.071777f
C1 a_36_472# VNW 0.013943f
C2 a_36_472# VDD 0.581285f
C3 A2 A1 0.047589f
C4 VDD VNW 0.11216f
C5 ZN A1 0.245346f
C6 B ZN 0.00761f
C7 a_36_472# A2 0.10395f
C8 a_244_68# VSS 0.00255f
C9 a_36_472# ZN 0.088503f
C10 VNW A2 0.128282f
C11 ZN VNW 0.014655f
C12 VDD A2 0.015143f
C13 VDD ZN 0.003129f
C14 VSS A1 0.021732f
C15 ZN A2 0.248411f
C16 B VSS 0.080416f
C17 a_36_472# VSS 0.004325f
C18 VNW VSS 0.009145f
C19 VDD VSS 0.01275f
C20 B A1 0.157699f
C21 a_36_472# A1 0.104556f
C22 a_244_68# ZN 0.008784f
C23 A2 VSS 0.069479f
C24 VNW A1 0.122087f
C25 B a_36_472# 0.01027f
C26 VDD A1 0.0167f
C27 ZN VSS 0.304078f
C28 B VNW 0.137038f
C29 VSS VPW 0.361309f
C30 VDD VPW 0.259458f
C31 ZN VPW 0.040013f
C32 B VPW 0.378232f
C33 A1 VPW 0.264815f
C34 A2 VPW 0.3189f
C35 VNW VPW 1.65967f
C36 a_36_472# VPW 0.031137f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW a_36_113#
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 a_36_113# VNW 0.160792f
C1 Z I 0.031362f
C2 VSS I 0.070302f
C3 a_36_113# VDD 0.278283f
C4 a_36_113# Z 0.191876f
C5 VNW VDD 0.088196f
C6 a_36_113# VSS 0.11114f
C7 VNW Z 0.030118f
C8 VNW VSS 0.009307f
C9 a_36_113# I 0.476912f
C10 Z VDD 0.085355f
C11 VSS VDD 0.009561f
C12 VNW I 0.152645f
C13 VSS Z 0.136942f
C14 I VDD 0.028968f
C15 VSS VPW 0.283681f
C16 Z VPW 0.117185f
C17 VDD VPW 0.180237f
C18 I VPW 0.336876f
C19 VNW VPW 1.31158f
C20 a_36_113# VPW 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW a_1916_375# a_1380_472#
+ a_3260_375# a_36_472# a_932_472# a_2812_375# a_2276_472# a_1828_472# a_3172_472#
+ a_572_375# a_2724_472# a_124_375# a_1468_375# a_1020_375# a_484_472# a_2364_375#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 VDD a_1916_375# 0.129962f
C1 VSS a_932_472# 0.142721f
C2 a_2364_375# a_2276_472# 0.285629f
C3 VSS a_1020_375# 0.131736f
C4 VDD a_572_375# 0.129962f
C5 a_2364_375# a_2724_472# 0.087174f
C6 a_2812_375# a_2724_472# 0.285629f
C7 a_3172_472# VSS 0.139489f
C8 VNW a_2276_472# 0.024018f
C9 VNW a_2724_472# 0.024018f
C10 a_1380_472# a_932_472# 0.013276f
C11 a_484_472# VNW 0.024018f
C12 a_1020_375# a_1380_472# 0.087174f
C13 a_1020_375# a_932_472# 0.285629f
C14 a_2276_472# a_2724_472# 0.013276f
C15 VDD a_2364_375# 0.129962f
C16 VDD a_2812_375# 0.129962f
C17 VNW a_1468_375# 0.181468f
C18 VSS a_1828_472# 0.142721f
C19 a_124_375# a_572_375# 0.013103f
C20 VSS a_1916_375# 0.131736f
C21 VSS a_572_375# 0.131736f
C22 VNW VDD 0.425768f
C23 VDD a_2276_472# 0.179463f
C24 a_1380_472# a_1828_472# 0.013276f
C25 VDD a_2724_472# 0.179463f
C26 a_2812_375# a_3260_375# 0.013103f
C27 a_484_472# VDD 0.179463f
C28 a_572_375# a_932_472# 0.087174f
C29 a_1020_375# a_572_375# 0.013103f
C30 VSS a_2364_375# 0.131736f
C31 VSS a_2812_375# 0.131736f
C32 VDD a_1468_375# 0.129962f
C33 VNW a_3260_375# 0.18122f
C34 a_124_375# VNW 0.180172f
C35 VNW VSS 0.035286f
C36 VSS a_2276_472# 0.142721f
C37 a_484_472# a_124_375# 0.087174f
C38 VSS a_2724_472# 0.142721f
C39 a_1828_472# a_1916_375# 0.285629f
C40 a_36_472# VNW 0.025611f
C41 a_484_472# VSS 0.142721f
C42 a_3172_472# a_2812_375# 0.087174f
C43 VNW a_1380_472# 0.024018f
C44 VSS a_1468_375# 0.131736f
C45 VNW a_932_472# 0.024018f
C46 VDD a_3260_375# 0.129266f
C47 a_484_472# a_36_472# 0.013276f
C48 VNW a_1020_375# 0.181468f
C49 a_3172_472# VNW 0.024396f
C50 a_124_375# VDD 0.12673f
C51 VDD VSS 0.052737f
C52 a_484_472# a_932_472# 0.013276f
C53 a_3172_472# a_2724_472# 0.013276f
C54 a_1380_472# a_1468_375# 0.285629f
C55 a_2364_375# a_1916_375# 0.013103f
C56 a_36_472# VDD 0.093681f
C57 a_1020_375# a_1468_375# 0.013103f
C58 VDD a_1380_472# 0.179463f
C59 VNW a_1828_472# 0.024018f
C60 VSS a_3260_375# 0.081304f
C61 VDD a_932_472# 0.179463f
C62 VNW a_1916_375# 0.181468f
C63 VDD a_1020_375# 0.129962f
C64 VNW a_572_375# 0.181468f
C65 a_1828_472# a_2276_472# 0.013276f
C66 a_2276_472# a_1916_375# 0.087174f
C67 a_3172_472# VDD 0.179463f
C68 a_124_375# VSS 0.131736f
C69 a_484_472# a_572_375# 0.285629f
C70 a_2812_375# a_2364_375# 0.013103f
C71 a_1828_472# a_1468_375# 0.087174f
C72 a_124_375# a_36_472# 0.285629f
C73 a_1468_375# a_1916_375# 0.013103f
C74 a_36_472# VSS 0.142026f
C75 VNW a_2364_375# 0.181468f
C76 VNW a_2812_375# 0.181468f
C77 VDD a_1828_472# 0.179463f
C78 a_3172_472# a_3260_375# 0.285629f
C79 VSS a_1380_472# 0.142721f
C80 VSS VPW 1.20585f
C81 VDD VPW 0.907304f
C82 VNW VPW 5.83682f
C83 a_3172_472# VPW 0.345058f
C84 a_2724_472# VPW 0.33241f
C85 a_2276_472# VPW 0.33241f
C86 a_1828_472# VPW 0.33241f
C87 a_1380_472# VPW 0.33241f
C88 a_932_472# VPW 0.33241f
C89 a_484_472# VPW 0.33241f
C90 a_36_472# VPW 0.404746f
C91 a_3260_375# VPW 0.233093f
C92 a_2812_375# VPW 0.17167f
C93 a_2364_375# VPW 0.17167f
C94 a_1916_375# VPW 0.17167f
C95 a_1468_375# VPW 0.17167f
C96 a_1020_375# VPW 0.17167f
C97 a_572_375# VPW 0.17167f
C98 a_124_375# VPW 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_455_68# a_271_68#
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 ZN a_271_68# 0.001916f
C1 ZN a_455_68# 0.002926f
C2 VSS a_271_68# 0.006038f
C3 VSS a_455_68# 0.006909f
C4 VNW A2 0.121191f
C5 A2 ZN 0.078589f
C6 A1 VDD 0.022021f
C7 A2 VSS 0.104901f
C8 VNW A1 0.12917f
C9 A3 A2 0.117566f
C10 A2 a_271_68# 0.004027f
C11 A2 a_455_68# 0.005127f
C12 A1 ZN 0.384588f
C13 A1 VSS 0.084906f
C14 A1 a_455_68# 0.004981f
C15 VNW VDD 0.112537f
C16 A2 A1 0.133044f
C17 ZN VDD 0.33173f
C18 VSS VDD 0.008734f
C19 VNW ZN 0.034322f
C20 VNW VSS 0.008577f
C21 A3 VDD 0.079999f
C22 VNW A3 0.148237f
C23 VSS ZN 0.064021f
C24 A3 ZN 0.008403f
C25 A2 VDD 0.023177f
C26 A3 VSS 0.07804f
C27 VSS VPW 0.307914f
C28 ZN VPW 0.133449f
C29 VDD VPW 0.241872f
C30 A1 VPW 0.287469f
C31 A2 VPW 0.25736f
C32 A3 VPW 0.326833f
C33 VNW VPW 1.48562f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW a_245_68#
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
C0 A1 a_245_68# 0.008831f
C1 A2 ZN 0.038658f
C2 A2 VDD 0.039698f
C3 a_245_68# VSS 0.002295f
C4 ZN VDD 0.240333f
C5 A1 VSS 0.131667f
C6 A1 VNW 0.119756f
C7 VSS VNW 0.006174f
C8 A1 A2 0.226398f
C9 A1 ZN 0.351362f
C10 A2 VSS 0.051087f
C11 A1 VDD 0.027485f
C12 ZN VSS 0.098328f
C13 VSS VDD 0.017706f
C14 A2 VNW 0.125396f
C15 ZN VNW 0.02653f
C16 VNW VDD 0.084263f
C17 VSS VPW 0.238729f
C18 ZN VPW 0.105772f
C19 VDD VPW 0.243067f
C20 A1 VPW 0.290957f
C21 A2 VPW 0.314823f
C22 VNW VPW 1.13753f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW a_255_603# a_67_603#
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VSS Z 0.158265f
C1 A2 a_255_603# 0.001961f
C2 VSS a_67_603# 0.250493f
C3 Z a_67_603# 0.181586f
C4 A2 A1 0.062395f
C5 VNW A1 0.220003f
C6 A2 VDD 0.147628f
C7 VNW VDD 0.11771f
C8 A2 VSS 0.025748f
C9 VNW VSS 0.010039f
C10 a_255_603# VDD 0.005359f
C11 A2 Z 0.027598f
C12 VNW Z 0.033884f
C13 A2 a_67_603# 0.505374f
C14 VNW a_67_603# 0.157241f
C15 VDD A1 0.01431f
C16 a_255_603# a_67_603# 0.007617f
C17 VSS A1 0.050738f
C18 VDD VSS 0.008648f
C19 A1 a_67_603# 0.540888f
C20 A2 VNW 0.216313f
C21 VDD Z 0.196046f
C22 VDD a_67_603# 0.307039f
C23 VSS VPW 0.359722f
C24 Z VPW 0.102754f
C25 VDD VPW 0.233025f
C26 A2 VPW 0.313441f
C27 A1 VPW 0.39469f
C28 VNW VPW 1.65967f
C29 a_67_603# VPW 0.345683f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VNW VPW a_36_68# a_1612_497#
+ a_2124_68# a_244_497# a_2960_68# a_3368_68# a_2552_68# a_1164_497# a_716_497#
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
C0 ZN C 0.514613f
C1 B VDD 0.100578f
C2 A2 a_36_68# 0.108262f
C3 VSS a_2960_68# 0.002422f
C4 A2 VDD 0.15752f
C5 VSS a_3368_68# 0.004815f
C6 a_1164_497# VDD 0.008664f
C7 VSS a_2552_68# 0.002422f
C8 a_2124_68# a_36_68# 0.012118f
C9 ZN VSS 0.006216f
C10 VDD a_36_68# 0.021485f
C11 ZN a_244_497# 0.009475f
C12 A2 A1 1.73987f
C13 B C 1.73339f
C14 ZN VNW 0.056895f
C15 a_1612_497# ZN 0.024559f
C16 A1 a_36_68# 0.065645f
C17 VDD A1 0.078657f
C18 B VSS 0.072527f
C19 C a_36_68# 0.105844f
C20 VDD C 0.095093f
C21 VSS A2 0.060501f
C22 A2 a_244_497# 0.01347f
C23 B VNW 0.600992f
C24 VNW A2 0.590323f
C25 B a_2960_68# 0.002626f
C26 VSS a_2124_68# 0.004133f
C27 VSS a_36_68# 3.64719f
C28 VSS VDD 0.005699f
C29 a_1612_497# A2 0.010709f
C30 VDD a_244_497# 0.020528f
C31 ZN a_716_497# 0.027752f
C32 B a_2552_68# 0.002588f
C33 VNW a_36_68# 0.004654f
C34 VNW VDD 0.366897f
C35 B ZN 0.426118f
C36 ZN A2 1.2828f
C37 a_2960_68# a_36_68# 0.009506f
C38 a_36_68# a_3368_68# 0.007478f
C39 a_1612_497# VDD 0.009792f
C40 VSS A1 0.060963f
C41 a_1164_497# ZN 0.021094f
C42 VSS C 0.092809f
C43 a_2552_68# a_36_68# 0.009506f
C44 ZN a_36_68# 1.98502f
C45 VNW A1 0.51833f
C46 ZN VDD 2.06829f
C47 A2 a_716_497# 0.00653f
C48 VNW C 0.636287f
C49 B A2 0.037299f
C50 a_1164_497# A2 0.009095f
C51 VDD a_716_497# 0.008599f
C52 ZN A1 1.37575f
C53 VSS VNW 0.004483f
C54 B a_36_68# 1.37417f
C55 VSS VPW 1.08055f
C56 ZN VPW 0.051826f
C57 VDD VPW 0.846798f
C58 C VPW 1.06351f
C59 B VPW 1.11555f
C60 A1 VPW 1.1956f
C61 A2 VPW 1.16629f
C62 VNW VPW 5.892971f
C63 a_36_68# VPW 0.063181f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW a_36_160#
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
C0 I Z 0.016176f
C1 I VNW 0.1633f
C2 I VDD 0.028233f
C3 Z VNW 0.021185f
C4 I VSS 0.178818f
C5 Z VDD 0.161733f
C6 I a_36_160# 0.564508f
C7 VSS Z 0.111496f
C8 VDD VNW 0.111398f
C9 a_36_160# Z 0.426617f
C10 VSS VNW 0.00834f
C11 VSS VDD 0.01316f
C12 a_36_160# VNW 0.302514f
C13 a_36_160# VDD 0.31851f
C14 VSS a_36_160# 0.114407f
C15 VSS VPW 0.397291f
C16 Z VPW 0.097163f
C17 VDD VPW 0.238155f
C18 I VPW 0.333888f
C19 VNW VPW 1.65967f
C20 a_36_160# VPW 0.696445f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW a_1380_472# a_36_472#
+ a_932_472# a_572_375# a_124_375# a_1468_375# a_1020_375# a_484_472#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_572_375# VDD 0.129962f
C1 a_572_375# a_484_472# 0.285629f
C2 VNW a_932_472# 0.024018f
C3 a_1468_375# a_1380_472# 0.285629f
C4 VSS VDD 0.026369f
C5 VNW a_124_375# 0.180172f
C6 a_484_472# VSS 0.148077f
C7 a_484_472# VDD 0.179463f
C8 a_1468_375# a_1020_375# 0.012552f
C9 a_1380_472# VSS 0.144845f
C10 a_1380_472# VDD 0.179463f
C11 a_572_375# a_1020_375# 0.012552f
C12 VSS a_1020_375# 0.134699f
C13 a_1020_375# VDD 0.129962f
C14 a_36_472# VSS 0.147381f
C15 a_36_472# VDD 0.093681f
C16 a_484_472# a_36_472# 0.013276f
C17 a_932_472# a_572_375# 0.086905f
C18 a_1380_472# a_1020_375# 0.086905f
C19 a_124_375# a_572_375# 0.012552f
C20 a_932_472# VSS 0.148077f
C21 a_932_472# VDD 0.179463f
C22 VNW a_1468_375# 0.18122f
C23 a_932_472# a_484_472# 0.013276f
C24 VNW a_572_375# 0.181468f
C25 a_1380_472# a_932_472# 0.013276f
C26 a_124_375# VSS 0.134699f
C27 a_124_375# VDD 0.12673f
C28 a_124_375# a_484_472# 0.086905f
C29 VNW VSS 0.017643f
C30 VNW VDD 0.217349f
C31 VNW a_484_472# 0.024018f
C32 a_932_472# a_1020_375# 0.285629f
C33 VNW a_1380_472# 0.024396f
C34 a_124_375# a_36_472# 0.285629f
C35 VNW a_1020_375# 0.181468f
C36 VNW a_36_472# 0.025611f
C37 a_1468_375# VSS 0.082091f
C38 a_572_375# VSS 0.134699f
C39 a_1468_375# VDD 0.129266f
C40 VSS VPW 0.642184f
C41 VDD VPW 0.493288f
C42 VNW VPW 3.05206f
C43 a_1380_472# VPW 0.345058f
C44 a_932_472# VPW 0.33241f
C45 a_484_472# VPW 0.33241f
C46 a_36_472# VPW 0.404746f
C47 a_1468_375# VPW 0.233029f
C48 a_1020_375# VPW 0.171606f
C49 a_572_375# VPW 0.171606f
C50 a_124_375# VPW 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW a_36_68#
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 a_36_68# I 0.731677f
C1 a_36_68# VNW 0.296832f
C2 I VNW 0.133333f
C3 Z VSS 0.133443f
C4 Z VDD 0.172592f
C5 VDD VSS 0.014283f
C6 a_36_68# Z 0.432914f
C7 a_36_68# VSS 0.156367f
C8 I Z 0.018906f
C9 I VSS 0.128735f
C10 Z VNW 0.023138f
C11 VNW VSS 0.009972f
C12 a_36_68# VDD 0.271105f
C13 I VDD 0.029139f
C14 VDD VNW 0.114912f
C15 VSS VPW 0.338876f
C16 Z VPW 0.103236f
C17 VDD VPW 0.234026f
C18 I VPW 0.298844f
C19 VNW VPW 1.65967f
C20 a_36_68# VPW 0.69549f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW a_848_380# a_1084_68#
+ a_124_24# a_1152_472# a_692_472#
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
C0 Z I1 0.027341f
C1 Z VNW 0.020389f
C2 VNW I0 0.103064f
C3 a_124_24# a_1152_472# 0.00128f
C4 a_124_24# a_692_472# 0.033243f
C5 a_124_24# I1 0.564972f
C6 S a_1084_68# 0.001644f
C7 a_124_24# VNW 0.277682f
C8 a_848_380# S 0.754833f
C9 I1 a_692_472# 0.001219f
C10 Z VDD 0.20273f
C11 I0 VDD 0.028914f
C12 VNW I1 0.127749f
C13 Z VSS 0.129676f
C14 I0 VSS 0.124513f
C15 a_124_24# VDD 0.309232f
C16 a_124_24# VSS 0.501844f
C17 a_1152_472# VDD 0.00645f
C18 VDD a_692_472# 0.009663f
C19 I1 VDD 0.227359f
C20 I1 VSS 0.026996f
C21 VNW VDD 0.182986f
C22 VNW VSS 0.009598f
C23 S I0 0.533789f
C24 I0 a_1084_68# 0.00492f
C25 a_124_24# S 0.245829f
C26 a_848_380# I0 0.082224f
C27 VSS VDD 0.028952f
C28 a_124_24# a_1084_68# 0.002839f
C29 S a_692_472# 0.002582f
C30 a_848_380# a_124_24# 0.302602f
C31 S I1 0.042269f
C32 VNW S 0.253706f
C33 a_848_380# a_1152_472# 0.007362f
C34 a_124_24# a_692_68# 0.006853f
C35 a_848_380# a_692_472# 0.003985f
C36 a_848_380# I1 0.013444f
C37 a_848_380# VNW 0.174516f
C38 S VDD 0.056165f
C39 S VSS 0.081531f
C40 a_848_380# VDD 0.319708f
C41 VSS a_1084_68# 0.009508f
C42 a_848_380# VSS 0.130064f
C43 Z a_124_24# 0.219295f
C44 a_124_24# I0 0.004772f
C45 VSS a_692_68# 0.001982f
C46 VSS VPW 0.565512f
C47 Z VPW 0.047467f
C48 VDD VPW 0.424967f
C49 I0 VPW 0.267152f
C50 S VPW 0.549493f
C51 I1 VPW 0.247562f
C52 VNW VPW 2.87801f
C53 a_848_380# VPW 0.40208f
C54 a_124_24# VPW 0.591898f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW a_36_68# a_244_472#
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 VSS B 0.198567f
C1 A2 VDD 0.017122f
C2 ZN a_244_472# 0.014146f
C3 ZN VDD 0.006004f
C4 VSS a_36_68# 0.117681f
C5 A2 VNW 0.122386f
C6 A2 A1 0.038725f
C7 VDD a_244_472# 0.004051f
C8 ZN VNW 0.011308f
C9 ZN A1 0.496662f
C10 VDD VNW 0.117098f
C11 VDD A1 0.014914f
C12 A2 a_36_68# 0.489122f
C13 VSS A2 0.083821f
C14 ZN a_36_68# 0.56857f
C15 A1 VNW 0.117811f
C16 VDD B 0.07579f
C17 VSS ZN 0.088946f
C18 a_36_68# a_244_472# 0.013419f
C19 VDD a_36_68# 0.753239f
C20 B VNW 0.163023f
C21 VSS VDD 0.004855f
C22 B A1 0.034707f
C23 a_36_68# VNW 0.038286f
C24 a_36_68# A1 0.292244f
C25 VSS VNW 0.0064f
C26 VSS A1 0.090903f
C27 A2 ZN 0.400775f
C28 B a_36_68# 0.389329f
C29 VSS VPW 0.342662f
C30 ZN VPW 0.011384f
C31 VDD VPW 0.256635f
C32 B VPW 0.339176f
C33 A1 VPW 0.256004f
C34 A2 VPW 0.28395f
C35 VNW VPW 1.65967f
C36 a_36_68# VPW 0.112263f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW a_224_552#
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
C0 a_224_552# I 0.421587f
C1 a_224_552# VNW 0.5926f
C2 I VNW 0.376531f
C3 Z VSS 0.275062f
C4 Z VDD 0.356369f
C5 VDD VSS 0.030201f
C6 a_224_552# Z 1.17071f
C7 a_224_552# VSS 0.331404f
C8 I Z 0.002319f
C9 Z VNW 0.027266f
C10 I VSS 0.061715f
C11 VNW VSS 0.009226f
C12 a_224_552# VDD 0.347549f
C13 I VDD 0.069894f
C14 VDD VNW 0.176912f
C15 VSS VPW 0.628617f
C16 Z VPW 0.102362f
C17 VDD VPW 0.415149f
C18 I VPW 0.471574f
C19 VNW VPW 2.70396f
C20 a_224_552# VPW 1.31114f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW a_234_472# a_672_472#
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 a_234_472# ZN 0.003154f
C1 VSS VNW 0.010681f
C2 A1 VDD 0.037494f
C3 ZN VNW 0.03148f
C4 a_672_472# VDD 0.005379f
C5 ZN VSS 0.460527f
C6 A1 A2 0.636124f
C7 A2 VDD 0.13595f
C8 a_672_472# A2 0.0147f
C9 a_234_472# VDD 0.0121f
C10 VNW A1 0.25895f
C11 VNW VDD 0.137685f
C12 VSS A1 0.052992f
C13 a_234_472# A2 0.018681f
C14 VSS VDD 0.023993f
C15 ZN A1 0.274601f
C16 ZN VDD 0.517479f
C17 VNW A2 0.275679f
C18 a_672_472# ZN 0.023475f
C19 VSS A2 0.07211f
C20 ZN A2 0.509001f
C21 VSS VPW 0.451405f
C22 ZN VPW 0.138491f
C23 VDD VPW 0.322159f
C24 A1 VPW 0.557317f
C25 A2 VPW 0.617688f
C26 VNW VPW 2.00777f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_448_472# a_244_472#
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
C0 A3 a_244_472# 0.019089f
C1 VSS A1 0.025677f
C2 A3 VDD 0.201466f
C3 ZN a_244_472# 0.001803f
C4 ZN VDD 0.116419f
C5 A3 VNW 0.136756f
C6 VDD a_244_472# 0.006513f
C7 A3 A2 0.416588f
C8 ZN VNW 0.040402f
C9 ZN A2 0.096665f
C10 a_244_472# A2 0.003952f
C11 VDD VNW 0.11801f
C12 VDD A2 0.09496f
C13 ZN A1 0.499849f
C14 VSS A3 0.058214f
C15 ZN a_448_472# 0.006209f
C16 A2 VNW 0.116878f
C17 VDD A1 0.095023f
C18 VSS ZN 0.283414f
C19 VDD a_448_472# 0.013539f
C20 A1 VNW 0.127941f
C21 VSS VDD 0.01583f
C22 A1 A2 0.145555f
C23 a_448_472# A2 0.012315f
C24 VSS VNW 0.008407f
C25 VSS A2 0.027728f
C26 A3 ZN 0.035547f
C27 A1 a_448_472# 0.012619f
C28 VSS VPW 0.367618f
C29 ZN VPW 0.134331f
C30 VDD VPW 0.264623f
C31 A1 VPW 0.311038f
C32 A2 VPW 0.285534f
C33 A3 VPW 0.334053f
C34 VNW VPW 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VNW VPW a_36_68# a_1732_68#
+ a_244_68# a_1100_68# a_1528_68# a_672_68#
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
C0 ZN A2 1.77619f
C1 A1 A2 0.077487f
C2 ZN VNW 0.095885f
C3 VNW A1 0.700258f
C4 a_36_68# a_1100_68# 0.012396f
C5 a_36_68# a_672_68# 0.012389f
C6 a_36_68# A2 0.223434f
C7 a_36_68# VNW 0.007741f
C8 ZN VDD 1.57207f
C9 A1 VDD 0.115489f
C10 ZN VSS 0.00864f
C11 VNW A2 0.630933f
C12 A1 VSS 0.065524f
C13 a_36_68# VDD 0.029088f
C14 a_36_68# VSS 2.77545f
C15 A2 VDD 0.124271f
C16 VSS a_1100_68# 0.003125f
C17 VSS a_672_68# 0.003125f
C18 A2 VSS 0.070822f
C19 VNW VDD 0.292073f
C20 VNW VSS 0.003704f
C21 ZN A3 0.150755f
C22 A3 A1 0.001696f
C23 ZN a_1732_68# 0.002613f
C24 a_36_68# A3 1.03106f
C25 VSS VDD 0.004708f
C26 A3 a_1100_68# 0.003385f
C27 a_36_68# a_1732_68# 0.011094f
C28 A3 a_672_68# 0.003442f
C29 a_244_68# a_36_68# 0.009768f
C30 A3 A2 1.65768f
C31 VNW A3 0.599629f
C32 a_36_68# a_1528_68# 0.012072f
C33 A3 VDD 0.107959f
C34 A3 VSS 0.09506f
C35 ZN A1 1.266f
C36 VSS a_1732_68# 0.002237f
C37 a_244_68# VSS 0.006268f
C38 ZN a_36_68# 0.885472f
C39 a_36_68# A1 0.118844f
C40 VSS a_1528_68# 0.003775f
C41 VSS VPW 0.861061f
C42 ZN VPW 0.103891f
C43 VDD VPW 0.701563f
C44 A1 VPW 1.27704f
C45 A3 VPW 1.11693f
C46 A2 VPW 1.08692f
C47 VNW VPW 4.73584f
C48 a_36_68# VPW 0.061249f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW a_36_159#
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
C0 A1 a_36_159# 0.377122f
C1 VSS a_36_159# 0.244357f
C2 VSS Z 0.102819f
C3 A1 VNW 0.206765f
C4 A1 A2 0.061431f
C5 Z a_36_159# 0.215269f
C6 VSS VNW 0.007925f
C7 VSS A2 0.011099f
C8 a_36_159# VNW 0.162496f
C9 A1 VDD 0.04397f
C10 a_36_159# A2 0.472781f
C11 Z VNW 0.032842f
C12 Z A2 0.020174f
C13 VSS VDD 0.014131f
C14 VDD a_36_159# 0.130189f
C15 VSS a_244_159# 0.001449f
C16 A2 VNW 0.20463f
C17 Z VDD 0.158212f
C18 a_244_159# a_36_159# 0.003343f
C19 VDD VNW 0.125609f
C20 VDD A2 0.184025f
C21 A1 VSS 0.010276f
C22 VSS VPW 0.35312f
C23 Z VPW 0.096476f
C24 VDD VPW 0.251252f
C25 A2 VPW 0.262264f
C26 A1 VPW 0.321274f
C27 VNW VPW 1.65967f
C28 a_36_159# VPW 0.374116f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VNW VPW a_2590_472#
+ a_170_472# a_1602_69# a_786_69# a_3126_472# a_1194_69# a_3662_472# a_2034_472# a_358_69#
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VPW nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VPW nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VPW nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
C0 a_170_472# VDD 2.96356f
C1 ZN VSS 1.77446f
C2 a_170_472# a_3126_472# 0.01307f
C3 VDD a_3126_472# 0.00779f
C4 ZN A2 1.83822f
C5 a_170_472# a_2590_472# 0.013379f
C6 VDD a_2590_472# 0.007681f
C7 ZN B 0.231932f
C8 A1 VSS 0.087217f
C9 VSS VNW 0.012025f
C10 A1 A2 1.72617f
C11 VNW A2 0.513788f
C12 A1 B 0.001644f
C13 VNW B 0.617219f
C14 a_170_472# VSS 0.00801f
C15 VDD VSS 0.016824f
C16 ZN C 1.79111f
C17 a_170_472# A2 0.109943f
C18 VDD A2 0.052548f
C19 a_170_472# B 2.12702f
C20 VSS a_1602_69# 0.005669f
C21 VDD B 0.110239f
C22 B a_3126_472# 0.007345f
C23 VSS a_1194_69# 0.005069f
C24 A1 C 0.001754f
C25 B a_2590_472# 0.007345f
C26 C VNW 0.61926f
C27 ZN a_358_69# 0.011344f
C28 ZN a_786_69# 0.008749f
C29 a_170_472# C 0.075372f
C30 VDD C 0.089678f
C31 VSS A2 0.104058f
C32 A1 a_358_69# 0.001641f
C33 VSS B 0.119454f
C34 A1 a_786_69# 0.001203f
C35 B A2 0.05388f
C36 a_2034_472# a_170_472# 0.020753f
C37 a_2034_472# VDD 0.008673f
C38 VSS C 0.088883f
C39 a_170_472# a_3662_472# 0.013628f
C40 VDD a_3662_472# 0.007223f
C41 C B 1.34577f
C42 A1 ZN 1.40746f
C43 ZN VNW 0.045695f
C44 VSS a_358_69# 0.005318f
C45 VSS a_786_69# 0.003966f
C46 a_170_472# ZN 0.818521f
C47 ZN VDD 0.008843f
C48 A1 VNW 0.480244f
C49 a_2034_472# B 0.008709f
C50 ZN a_1602_69# 0.008113f
C51 A1 a_170_472# 0.0698f
C52 ZN a_1194_69# 0.00847f
C53 A1 VDD 0.051939f
C54 a_170_472# VNW 0.018375f
C55 B a_3662_472# 0.007338f
C56 VDD VNW 0.393677f
C57 VSS VPW 1.33264f
C58 VDD VPW 0.809429f
C59 ZN VPW 0.171181f
C60 C VPW 1.26656f
C61 B VPW 1.19887f
C62 A1 VPW 1.12703f
C63 A2 VPW 1.09165f
C64 VNW VPW 6.53302f
C65 a_170_472# VPW 0.077257f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW a_1792_472# a_224_472#
+ a_1568_472# a_36_472# a_1120_472# a_672_472#
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
C0 VNW A2 0.539636f
C1 a_1120_472# VDD 0.011157f
C2 VSS VNW 0.009996f
C3 a_1568_472# a_36_472# 0.025433f
C4 A3 A2 1.6562f
C5 VDD ZN 0.005367f
C6 VSS A3 0.10353f
C7 a_224_472# a_36_472# 0.01823f
C8 VSS A2 0.128956f
C9 VNW a_36_472# 0.031928f
C10 VDD A1 0.054887f
C11 A1 ZN 1.56829f
C12 a_1792_472# a_36_472# 0.022081f
C13 A3 a_36_472# 0.100976f
C14 a_36_472# A2 0.993181f
C15 a_672_472# A2 0.002647f
C16 VSS a_36_472# 0.020716f
C17 a_1568_472# VDD 0.005385f
C18 a_1568_472# A1 0.002055f
C19 a_224_472# VDD 0.010911f
C20 a_1120_472# A2 0.002647f
C21 VNW VDD 0.286001f
C22 VNW ZN 0.046016f
C23 a_672_472# a_36_472# 0.01823f
C24 a_1792_472# VDD 0.002998f
C25 VNW A1 0.520086f
C26 a_1792_472# ZN 0.004144f
C27 A3 VDD 0.09322f
C28 VDD A2 0.082489f
C29 A3 ZN 1.42151f
C30 A2 ZN 0.250963f
C31 a_1792_472# A1 0.006624f
C32 VSS VDD 0.012739f
C33 a_1120_472# a_36_472# 0.01951f
C34 VSS ZN 2.18568f
C35 A3 A1 0.008795f
C36 A1 A2 0.085569f
C37 VSS A1 0.115774f
C38 a_36_472# VDD 1.90933f
C39 a_36_472# ZN 0.362263f
C40 a_672_472# VDD 0.01105f
C41 a_1568_472# A2 0.004974f
C42 a_36_472# A1 0.174868f
C43 VNW A3 0.478769f
C44 a_224_472# A2 0.002647f
C45 VSS VPW 0.918064f
C46 ZN VPW 0.159858f
C47 VDD VPW 0.61695f
C48 A1 VPW 1.35739f
C49 A3 VPW 1.33073f
C50 A2 VPW 1.29013f
C51 VNW VPW 4.79254f
C52 a_36_472# VPW 0.137725f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW a_468_472# a_244_472#
+ a_1130_472# a_906_472#
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 VDD VNW 0.178574f
C1 VNW A2 0.241313f
C2 A3 a_1130_472# 0.016495f
C3 VDD A1 0.038139f
C4 A2 A1 0.570018f
C5 A3 a_906_472# 0.017829f
C6 VDD ZN 0.579119f
C7 A2 ZN 0.694728f
C8 ZN a_468_472# 0.015602f
C9 VDD VSS 0.009106f
C10 ZN a_244_472# 0.019831f
C11 VSS A2 0.043139f
C12 VNW A1 0.254404f
C13 VNW ZN 0.031771f
C14 VDD A3 0.178286f
C15 A3 A2 0.624599f
C16 VDD a_1130_472# 0.011629f
C17 ZN A1 0.084783f
C18 VNW VSS 0.007164f
C19 VDD a_906_472# 0.011614f
C20 A3 a_468_472# 0.010018f
C21 A3 a_244_472# 0.010666f
C22 VNW A3 0.28584f
C23 VSS A1 0.044587f
C24 VSS ZN 1.3936f
C25 A3 A1 0.292395f
C26 A3 ZN 1.03634f
C27 VDD A2 0.038421f
C28 ZN a_1130_472# 0.001342f
C29 ZN a_906_472# 0.002855f
C30 VSS A3 0.0525f
C31 VDD a_468_472# 0.00502f
C32 VDD a_244_472# 0.00632f
C33 VSS VPW 0.509614f
C34 ZN VPW 0.172636f
C35 VDD VPW 0.441158f
C36 A1 VPW 0.622214f
C37 A2 VPW 0.627317f
C38 A3 VPW 0.692739f
C39 VNW VPW 2.70396f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VNW VPW a_1492_488#
+ a_244_68# a_1044_488# a_636_68# a_36_488#
X0 VSS B ZN VPW nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VPW nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
C0 a_244_68# VSS 0.004878f
C1 a_36_488# ZN 0.459425f
C2 a_36_488# VDD 1.67897f
C3 ZN VDD 0.004894f
C4 A2 B 0.036672f
C5 VSS B 0.089442f
C6 A2 A1 0.652956f
C7 a_36_488# C 0.041645f
C8 VSS A1 0.090485f
C9 ZN C 0.191881f
C10 VSS A2 0.077665f
C11 C VDD 0.040747f
C12 B a_1492_488# 0.007233f
C13 VNW a_36_488# 0.010653f
C14 VNW ZN 0.028815f
C15 VNW VDD 0.191798f
C16 VSS a_636_68# 0.002222f
C17 a_36_488# a_1044_488# 0.018358f
C18 VNW C 0.268332f
C19 a_244_68# ZN 0.001328f
C20 a_1044_488# VDD 0.004195f
C21 a_36_488# B 0.80489f
C22 a_36_488# A1 0.031215f
C23 B ZN 0.413891f
C24 ZN A1 0.372797f
C25 B VDD 0.04259f
C26 A2 a_36_488# 0.076279f
C27 VSS a_36_488# 0.005331f
C28 A1 VDD 0.026261f
C29 A2 ZN 0.752866f
C30 VSS ZN 0.708286f
C31 A2 VDD 0.02614f
C32 B C 0.560408f
C33 VSS VDD 0.009527f
C34 a_36_488# a_1492_488# 0.017313f
C35 VSS C 0.05406f
C36 a_1492_488# VDD 0.00909f
C37 a_636_68# ZN 0.00593f
C38 VNW B 0.298561f
C39 VNW A1 0.25321f
C40 VNW A2 0.280457f
C41 VNW VSS 0.008434f
C42 a_244_68# A1 0.003444f
C43 a_1044_488# B 0.012375f
C44 VSS VPW 0.653933f
C45 VDD VPW 0.406726f
C46 ZN VPW 0.089692f
C47 C VPW 0.626227f
C48 B VPW 0.654892f
C49 A1 VPW 0.552174f
C50 A2 VPW 0.559992f
C51 VNW VPW 3.2261f
C52 a_36_488# VPW 0.101145f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VNW VPW a_244_524# a_2215_68#
+ a_56_524# a_718_524# a_728_93# a_1936_472# a_1336_472#
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
C0 A2 a_718_524# 0.107911f
C1 A1 VNW 0.293766f
C2 A3 a_1336_472# 0.490376f
C3 Z a_728_93# 0.402606f
C4 A3 a_1936_472# 0.018144f
C5 VDD A1 0.018915f
C6 a_1336_472# Z 0.021039f
C7 A3 VSS 0.056027f
C8 a_1936_472# Z 0.337902f
C9 A2 a_244_524# 0.004824f
C10 a_56_524# a_728_93# 0.016741f
C11 Z VSS 0.277351f
C12 A3 VNW 0.268193f
C13 a_1336_472# a_728_93# 0.62718f
C14 a_1936_472# a_728_93# 0.105997f
C15 A3 VDD 0.028848f
C16 A2 A1 0.321942f
C17 VSS a_56_524# 0.214447f
C18 Z VNW 0.028011f
C19 VSS a_728_93# 0.709567f
C20 a_1936_472# a_1336_472# 0.004622f
C21 VDD Z 0.01058f
C22 a_1336_472# VSS 0.326133f
C23 a_56_524# VNW 0.188846f
C24 VNW a_728_93# 0.346549f
C25 VDD a_56_524# 0.049641f
C26 A1 a_718_524# 0.026418f
C27 VDD a_728_93# 0.575073f
C28 a_1336_472# VNW 0.144065f
C29 a_1936_472# VNW 0.004015f
C30 a_1336_472# VDD 0.033982f
C31 a_1936_472# VDD 0.595117f
C32 VSS VNW 0.007756f
C33 VDD VSS 0.013872f
C34 A2 a_56_524# 0.908796f
C35 a_2215_68# Z 0.008507f
C36 A2 a_728_93# 0.416172f
C37 VDD VNW 0.360391f
C38 a_1336_472# A2 0.001757f
C39 A2 VSS 0.047538f
C40 a_56_524# a_718_524# 0.009198f
C41 a_718_524# a_728_93# 0.329834f
C42 a_728_93# a_1524_472# 0.007139f
C43 A2 VNW 0.369075f
C44 a_2215_68# VSS 0.004309f
C45 a_1336_472# a_1524_472# 0.001046f
C46 A2 VDD 0.208821f
C47 A1 a_56_524# 0.569057f
C48 VNW a_718_524# 0.020055f
C49 A1 a_728_93# 0.12992f
C50 VDD a_718_524# 0.554575f
C51 a_952_93# a_728_93# 0.00421f
C52 A3 Z 0.259021f
C53 A1 VSS 0.139902f
C54 VDD a_244_524# 0.004322f
C55 A3 a_728_93# 0.720358f
C56 VSS VPW 0.861752f
C57 Z VPW 0.085787f
C58 A1 VPW 0.602985f
C59 A2 VPW 0.640744f
C60 VDD VPW 0.543474f
C61 A3 VPW 0.593976f
C62 VNW VPW 4.270391f
C63 a_1936_472# VPW 0.009918f
C64 a_718_524# VPW 0.005143f
C65 a_56_524# VPW 0.41096f
C66 a_728_93# VPW 0.654825f
C67 a_1336_472# VPW 0.316639f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VNW VPW a_652_68# a_244_68#
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
C0 A1 VSS 0.115936f
C1 ZN VDD 0.409997f
C2 A1 VDD 0.050088f
C3 ZN a_244_68# 0.001926f
C4 VNW A2 0.277885f
C5 VDD VSS 0.020712f
C6 A1 a_244_68# 0.004867f
C7 VSS a_244_68# 0.006834f
C8 VNW ZN 0.033841f
C9 VNW A1 0.232646f
C10 VNW VSS 0.008805f
C11 VNW VDD 0.123338f
C12 ZN A2 0.891023f
C13 A2 A1 0.708017f
C14 A2 VSS 0.057292f
C15 a_652_68# ZN 0.008436f
C16 ZN A1 0.363066f
C17 A2 VDD 0.070487f
C18 a_652_68# VSS 0.003855f
C19 ZN VSS 0.2597f
C20 VSS VPW 0.385688f
C21 ZN VPW 0.120217f
C22 VDD VPW 0.305683f
C23 A1 VPW 0.522064f
C24 A2 VPW 0.568932f
C25 VNW VPW 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VNW VPW a_36_68# a_1612_497#
+ a_692_497# a_1388_497# a_960_497#
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
C0 VSS B 0.047409f
C1 A2 a_1388_497# 0.008156f
C2 VDD a_692_497# 0.00542f
C3 A2 a_1612_497# 0.006056f
C4 VDD B 0.119783f
C5 A3 A1 0.206693f
C6 a_36_68# VSS 2.0408f
C7 a_36_68# VDD 0.001802f
C8 A2 a_960_497# 0.003506f
C9 VSS ZN 0.006088f
C10 VDD ZN 1.08837f
C11 a_36_68# B 0.184521f
C12 A2 A1 0.703324f
C13 VSS A3 0.03178f
C14 ZN a_692_497# 0.018589f
C15 ZN B 0.244028f
C16 A3 VDD 0.555327f
C17 VNW A1 0.279057f
C18 a_36_68# ZN 1.49222f
C19 A3 a_692_497# 0.019827f
C20 A3 B 0.036798f
C21 A1 a_1612_497# 0.003158f
C22 A2 VSS 0.030287f
C23 A2 VDD 0.030601f
C24 a_36_68# A3 0.036843f
C25 A3 ZN 1.02771f
C26 VNW VSS 0.008187f
C27 A2 a_692_497# 0.001398f
C28 VNW VDD 0.248379f
C29 VDD a_1388_497# 0.005409f
C30 VDD a_1612_497# 0.009412f
C31 a_36_68# A2 0.032025f
C32 VNW B 0.309147f
C33 A2 ZN 0.152712f
C34 VDD a_960_497# 0.003264f
C35 a_36_68# VNW 0.001442f
C36 VNW ZN 0.025446f
C37 VSS A1 0.032188f
C38 A2 A3 1.11591f
C39 A1 VDD 0.091309f
C40 ZN a_1388_497# 0.001168f
C41 VNW A3 0.297068f
C42 ZN a_960_497# 0.012124f
C43 A3 a_1388_497# 0.02079f
C44 A3 a_1612_497# 0.030605f
C45 a_36_68# A1 0.158235f
C46 VSS VDD 0.010407f
C47 A1 ZN 0.619225f
C48 A3 a_960_497# 0.014254f
C49 A2 VNW 0.281901f
C50 VSS VPW 0.663038f
C51 ZN VPW 0.080495f
C52 VDD VPW 0.512998f
C53 A1 VPW 0.643779f
C54 A2 VPW 0.561227f
C55 A3 VPW 0.573818f
C56 B VPW 0.585725f
C57 VNW VPW 3.48825f
C58 a_36_68# VPW 0.048026f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VNW VPW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_2248_156#
+ a_2560_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VPW nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 VSS a_2665_112# 0.21484f
C1 a_36_151# RN 0.080119f
C2 a_448_472# a_1456_156# 0.00227f
C3 a_2248_156# VSS 0.030372f
C4 a_36_151# a_1308_423# 0.05539f
C5 a_1000_472# VSS 0.04356f
C6 VDD a_2560_156# 0.00302f
C7 VNW a_36_151# 1.28833f
C8 a_448_472# a_1288_156# 0.002067f
C9 a_1204_472# a_1000_472# 0.66083f
C10 VDD a_2665_112# 0.152571f
C11 a_2560_156# a_2665_112# 0.116229f
C12 a_796_472# a_1000_472# 0.048436f
C13 a_448_472# RN 0.078731f
C14 a_2248_156# VDD 1.12036f
C15 a_2248_156# a_2560_156# 0.119687f
C16 a_2248_156# a_2665_112# 0.63615f
C17 a_448_472# a_1308_423# 0.882105f
C18 a_36_151# VSS 0.291264f
C19 a_1000_472# VDD 0.119211f
C20 a_1204_472# a_36_151# 0.006996f
C21 VNW a_448_472# 0.341284f
C22 a_36_151# a_796_472# 0.011851f
C23 a_2248_156# a_1000_472# 0.001232f
C24 RN a_3041_156# 0.014924f
C25 VNW D 0.128231f
C26 a_36_151# VDD 0.417101f
C27 a_36_151# a_2560_156# 0.003674f
C28 VNW CLK 0.137037f
C29 a_448_472# VSS 1.20207f
C30 a_36_151# a_2665_112# 0.019033f
C31 VNW Q 0.026596f
C32 a_448_472# a_1204_472# 0.008996f
C33 a_2248_156# a_36_151# 0.042802f
C34 a_448_472# a_796_472# 0.401636f
C35 D VSS 0.064618f
C36 CLK VSS 0.021952f
C37 a_36_151# a_1000_472# 0.08126f
C38 Q VSS 0.170514f
C39 a_448_472# VDD 0.456269f
C40 a_796_472# D 0.082858f
C41 a_1308_423# RN 0.079294f
C42 a_448_472# a_2560_156# 0.277491f
C43 VSS a_1456_156# 0.001901f
C44 a_448_472# a_2665_112# 0.020455f
C45 VSS a_3041_156# 0.004935f
C46 VNW RN 0.304626f
C47 D VDD 0.009367f
C48 a_2248_156# a_448_472# 0.510371f
C49 CLK VDD 0.02303f
C50 VNW a_1308_423# 0.149014f
C51 VSS a_1288_156# 0.001702f
C52 Q VDD 0.260055f
C53 a_448_472# a_1000_472# 0.361958f
C54 Q a_2665_112# 0.263315f
C55 RN VSS 0.436942f
C56 a_1204_472# RN 0.021039f
C57 a_2665_112# a_3041_156# 0.001841f
C58 a_2248_156# Q 0.013765f
C59 a_1308_423# VSS 0.013866f
C60 a_1204_472# a_1308_423# 0.026665f
C61 a_448_472# a_36_151# 0.536965f
C62 VNW VSS 0.012596f
C63 VNW a_1204_472# 0.016269f
C64 RN VDD 0.035003f
C65 RN a_2560_156# 0.038779f
C66 VNW a_796_472# 0.010232f
C67 RN a_2665_112# 0.322698f
C68 a_36_151# D 0.094113f
C69 a_1308_423# VDD 0.094185f
C70 CLK a_36_151# 0.669598f
C71 a_2248_156# RN 0.080362f
C72 VNW VDD 0.546785f
C73 VNW a_2560_156# 0.019282f
C74 VNW a_2665_112# 0.486803f
C75 a_2248_156# a_1308_423# 0.056721f
C76 a_796_472# VSS 0.05215f
C77 a_1000_472# RN 0.0832f
C78 VNW a_2248_156# 0.181292f
C79 a_1308_423# a_1000_472# 0.934191f
C80 a_448_472# D 0.328788f
C81 VSS VDD 0.02167f
C82 a_448_472# CLK 0.002757f
C83 VSS a_2560_156# 0.128503f
C84 a_1204_472# VDD 0.282626f
C85 VNW a_1000_472# 0.241357f
C86 Q VPW 0.061347f
C87 VSS VPW 1.33519f
C88 RN VPW 1.37098f
C89 D VPW 0.253406f
C90 VDD VPW 0.859994f
C91 CLK VPW 0.291241f
C92 VNW VPW 6.48579f
C93 a_2560_156# VPW 0.016968f
C94 a_2665_112# VPW 0.91969f
C95 a_2248_156# VPW 0.30886f
C96 a_1204_472# VPW 0.012971f
C97 a_1000_472# VPW 0.291735f
C98 a_796_472# VPW 0.023206f
C99 a_1308_423# VPW 0.279043f
C100 a_448_472# VPW 0.684413f
C101 a_36_151# VPW 1.43587f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW a_438_68#
+ a_244_68# a_1254_68# a_1060_68# a_632_68# a_1458_68#
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
C0 A4 A2 0.762551f
C1 A3 A4 0.297972f
C2 VNW A4 0.388525f
C3 a_1060_68# VSS 0.001868f
C4 a_438_68# VSS 0.00542f
C5 A1 A2 0.516286f
C6 A3 a_632_68# 0.0083f
C7 VDD VSS 0.004026f
C8 A3 A1 0.831807f
C9 a_1060_68# ZN 0.007219f
C10 VNW A1 0.345207f
C11 A3 A2 0.40854f
C12 VNW A2 0.317841f
C13 VDD ZN 1.39778f
C14 VNW A3 0.300046f
C15 ZN VSS 0.89636f
C16 a_1254_68# VSS 0.002331f
C17 a_1254_68# ZN 0.008913f
C18 a_244_68# VSS 0.007139f
C19 A4 VDD 0.047422f
C20 a_1458_68# VSS 0.002548f
C21 A4 VSS 0.056757f
C22 a_1458_68# ZN 0.01082f
C23 A4 ZN 1.94271f
C24 A1 VDD 0.044019f
C25 A3 a_1060_68# 0.004303f
C26 a_632_68# VSS 0.005832f
C27 VDD A2 0.041932f
C28 A1 VSS 0.037456f
C29 A3 a_438_68# 0.007312f
C30 A2 VSS 0.036637f
C31 A3 VDD 0.040467f
C32 VNW VDD 0.1769f
C33 a_632_68# ZN 0.001673f
C34 A3 VSS 0.248503f
C35 A1 ZN 0.071728f
C36 VNW VSS 0.006403f
C37 ZN A2 0.068627f
C38 A3 ZN 0.881941f
C39 VNW ZN 0.062752f
C40 A3 a_1254_68# 0.004873f
C41 a_244_68# A3 0.007f
C42 A4 A1 0.451294f
C43 VSS VPW 0.597574f
C44 VDD VPW 0.397078f
C45 ZN VPW 0.12583f
C46 A1 VPW 0.558392f
C47 A2 VPW 0.513744f
C48 A3 VPW 0.547819f
C49 A4 VPW 0.580825f
C50 VNW VPW 3.05206f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
C0 VDD I 0.164681f
C1 VNW VDD 0.103267f
C2 VNW I 0.283715f
C3 VSS ZN 0.15979f
C4 VDD VSS 0.022662f
C5 VSS I 0.071429f
C6 VNW VSS 0.01054f
C7 VDD ZN 0.24022f
C8 ZN I 0.614595f
C9 VNW ZN 0.025997f
C10 VSS VPW 0.345063f
C11 ZN VPW 0.094435f
C12 VDD VPW 0.235951f
C13 I VPW 0.642286f
C14 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VNW VPW a_468_472#
+ a_224_472# a_244_68# a_916_472#
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
C0 B1 VDD 0.015317f
C1 VSS a_224_472# 0.00124f
C2 VDD VNW 0.158216f
C3 B2 a_244_68# 0.29062f
C4 A1 A2 0.038953f
C5 B1 VNW 0.116377f
C6 VDD A3 0.236688f
C7 a_244_68# a_916_472# 0.018012f
C8 VNW A3 0.13805f
C9 a_468_472# a_244_68# 0.022611f
C10 VSS B2 0.072128f
C11 VSS a_244_68# 0.329999f
C12 a_224_472# A2 0.014544f
C13 VDD ZN 0.006472f
C14 B1 ZN 0.457921f
C15 ZN VNW 0.012941f
C16 A1 VDD 0.015114f
C17 A2 a_244_68# 0.356992f
C18 A1 B1 0.13457f
C19 A1 VNW 0.125824f
C20 a_468_472# A2 0.002382f
C21 VSS A2 0.030842f
C22 a_224_472# VDD 0.016257f
C23 A1 ZN 0.164807f
C24 a_224_472# A3 0.012212f
C25 VDD B2 0.018546f
C26 VDD a_244_68# 0.520053f
C27 B1 B2 0.038725f
C28 B1 a_244_68# 0.212448f
C29 VDD a_916_472# 0.004169f
C30 B2 VNW 0.125762f
C31 a_244_68# VNW 0.043485f
C32 a_468_472# VDD 0.005594f
C33 VSS VDD 0.027141f
C34 a_244_68# A3 0.010697f
C35 VSS B1 0.072063f
C36 VSS VNW 0.013582f
C37 VSS A3 0.046517f
C38 ZN B2 0.371232f
C39 ZN a_244_68# 0.2576f
C40 ZN a_916_472# 0.008827f
C41 A2 VDD 0.071137f
C42 VSS ZN 0.069913f
C43 A2 VNW 0.121626f
C44 A1 a_244_68# 0.480797f
C45 A2 A3 0.129823f
C46 A1 a_468_472# 0.001494f
C47 A1 VSS 0.029231f
C48 a_224_472# a_244_68# 0.004752f
C49 VSS VPW 0.474343f
C50 ZN VPW 0.00986f
C51 VDD VPW 0.363224f
C52 B2 VPW 0.282623f
C53 B1 VPW 0.257203f
C54 A1 VPW 0.255736f
C55 A2 VPW 0.254473f
C56 A3 VPW 0.308666f
C57 VNW VPW 2.35586f
C58 a_244_68# VPW 0.138666f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_244_567# a_718_527#
+ a_2172_497# a_56_567# a_1948_68# a_728_93# a_1296_93#
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
C0 a_1948_68# VNW 0.002346f
C1 a_56_567# a_718_527# 0.00772f
C2 VSS A3 0.047056f
C3 VSS VNW 0.009921f
C4 a_1296_93# ZN 0.029802f
C5 a_718_527# A2 0.141128f
C6 a_728_93# a_1296_93# 0.624643f
C7 a_56_567# A2 0.174541f
C8 A1 a_718_527# 0.023145f
C9 a_56_567# A1 0.368741f
C10 A3 VNW 0.298581f
C11 a_952_93# VSS 0.003841f
C12 A1 A2 0.757944f
C13 a_718_527# VDD 0.618394f
C14 a_56_567# VDD 0.056918f
C15 a_1948_68# a_1296_93# 0.005923f
C16 A2 VDD 0.210416f
C17 A1 VDD 0.022573f
C18 a_1296_93# VSS 0.379749f
C19 a_728_93# a_718_527# 0.21558f
C20 a_1296_93# A3 0.356198f
C21 a_728_93# a_56_567# 0.070648f
C22 a_1296_93# VNW 0.155715f
C23 a_2172_497# VDD 0.010751f
C24 a_728_93# A2 0.516752f
C25 a_728_93# A1 0.281966f
C26 ZN VDD 0.47211f
C27 a_728_93# VDD 0.78216f
C28 ZN a_2172_497# 0.03345f
C29 a_728_93# a_2172_497# 0.010602f
C30 a_56_567# VSS 0.400197f
C31 a_56_567# a_244_567# 0.00105f
C32 VSS A2 0.051212f
C33 a_718_527# VNW 0.020227f
C34 VSS a_1504_93# 0.003902f
C35 A1 VSS 0.0538f
C36 a_56_567# VNW 0.187311f
C37 a_1948_68# VDD 0.001604f
C38 a_728_93# ZN 0.663929f
C39 a_244_567# A2 0.004089f
C40 A2 VNW 0.388997f
C41 A1 VNW 0.342048f
C42 VSS VDD 0.011823f
C43 a_244_567# VDD 0.006111f
C44 A3 VDD 0.022483f
C45 a_1948_68# ZN 0.381585f
C46 VDD VNW 0.370487f
C47 a_728_93# a_1948_68# 0.02618f
C48 ZN VSS 0.004739f
C49 a_728_93# VSS 0.328386f
C50 ZN A3 0.033406f
C51 a_1296_93# A2 0.002759f
C52 a_728_93# A3 0.721889f
C53 ZN VNW 0.032895f
C54 a_1296_93# a_1504_93# 0.003723f
C55 a_728_93# VNW 0.385878f
C56 a_1948_68# VSS 0.719859f
C57 a_728_93# a_952_93# 0.003723f
C58 a_1296_93# VDD 0.030892f
C59 a_1948_68# A3 0.069927f
C60 VSS VPW 0.875791f
C61 ZN VPW 0.08517f
C62 A1 VPW 0.604039f
C63 A2 VPW 0.633287f
C64 VDD VPW 0.584594f
C65 A3 VPW 0.573218f
C66 VNW VPW 4.42794f
C67 a_1948_68# VPW 0.022025f
C68 a_718_527# VPW 0.001795f
C69 a_56_567# VPW 0.424713f
C70 a_728_93# VPW 0.65929f
C71 a_1296_93# VPW 0.317801f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VNW VPW a_36_68# a_244_497#
+ a_1657_68# a_1229_68# a_716_497#
X0 a_1229_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
C0 VNW B 0.311256f
C1 C VSS 0.04168f
C2 A1 VSS 0.031008f
C3 A2 VNW 0.30827f
C4 ZN VNW 0.042076f
C5 A2 B 0.037237f
C6 a_1229_68# VSS 0.002856f
C7 A2 a_716_497# 0.010693f
C8 ZN B 0.3603f
C9 C a_36_68# 0.055076f
C10 ZN a_716_497# 0.025301f
C11 a_1657_68# VSS 0.002208f
C12 A1 a_36_68# 0.039393f
C13 A2 a_244_497# 0.020646f
C14 ZN a_244_497# 0.006285f
C15 C VDD 0.056662f
C16 a_1229_68# a_36_68# 0.011792f
C17 A1 VDD 0.033883f
C18 ZN A2 1.02528f
C19 a_36_68# VSS 2.1107f
C20 a_1657_68# a_36_68# 0.009002f
C21 VDD VSS 0.007619f
C22 VDD a_36_68# 0.019083f
C23 VNW C 0.309331f
C24 A1 VNW 0.269127f
C25 C B 0.698524f
C26 VNW VSS 0.005994f
C27 B a_1229_68# 0.003462f
C28 a_1657_68# B 0.002626f
C29 B VSS 0.032629f
C30 ZN C 0.501479f
C31 A2 A1 0.722847f
C32 ZN A1 0.622246f
C33 VNW a_36_68# 0.00468f
C34 B a_36_68# 0.587375f
C35 A2 VSS 0.030494f
C36 VNW VDD 0.219901f
C37 ZN VSS 0.004788f
C38 VDD B 0.089771f
C39 VDD a_716_497# 0.008883f
C40 A2 a_36_68# 0.091399f
C41 VDD a_244_497# 0.016799f
C42 ZN a_36_68# 0.528658f
C43 A2 VDD 0.147417f
C44 ZN VDD 0.761655f
C45 VSS VPW 0.620026f
C46 ZN VPW 0.062404f
C47 VDD VPW 0.531064f
C48 C VPW 0.529789f
C49 B VPW 0.589191f
C50 A1 VPW 0.58772f
C51 A2 VPW 0.613706f
C52 VNW VPW 3.34705f
C53 a_36_68# VPW 0.052951f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW a_428_148# a_36_148#
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
C0 A2 VDD 0.022493f
C1 a_36_148# a_428_148# 0.007047f
C2 A3 A2 0.340591f
C3 VNW A2 0.189332f
C4 a_36_148# A1 0.205722f
C5 Z VDD 0.164783f
C6 A3 Z 0.001054f
C7 VNW Z 0.033257f
C8 a_36_148# VSS 0.798993f
C9 A3 VDD 0.022574f
C10 VNW VDD 0.134134f
C11 VNW A3 0.213241f
C12 VSS A1 0.00434f
C13 a_36_148# A2 0.141951f
C14 A2 A1 0.307806f
C15 a_36_148# a_244_148# 0.004781f
C16 a_36_148# Z 0.156534f
C17 a_36_148# VDD 0.556761f
C18 A2 VSS 0.004456f
C19 A3 a_428_148# 0.001335f
C20 a_244_148# A1 0.002081f
C21 A3 a_36_148# 0.477475f
C22 VNW a_36_148# 0.194548f
C23 VDD A1 0.021719f
C24 Z VSS 0.093779f
C25 VNW A1 0.214361f
C26 VSS VDD 0.012823f
C27 A3 VSS 0.005273f
C28 VNW VSS 0.007319f
C29 VSS VPW 0.415001f
C30 Z VPW 0.095371f
C31 VDD VPW 0.277732f
C32 A3 VPW 0.275015f
C33 A2 VPW 0.257076f
C34 A1 VPW 0.330738f
C35 VNW VPW 2.00777f
C36 a_36_148# VPW 0.388358f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW a_1044_68# a_452_68#
+ a_276_68# a_860_68#
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 A1 ZN 0.430404f
C1 VNW ZN 0.034063f
C2 A1 VNW 0.280755f
C3 ZN a_1044_68# 0.001223f
C4 ZN VSS 0.476547f
C5 A1 VSS 0.050488f
C6 VNW VSS 0.007349f
C7 A3 ZN 1.24554f
C8 A1 A3 0.037905f
C9 VSS a_1044_68# 0.00861f
C10 VNW A3 0.347673f
C11 A2 ZN 0.082264f
C12 A1 A2 0.708241f
C13 A3 VSS 0.074424f
C14 A2 VNW 0.279783f
C15 ZN VDD 0.550625f
C16 ZN a_860_68# 0.001808f
C17 A1 VDD 0.041745f
C18 ZN a_452_68# 0.007752f
C19 A2 a_1044_68# 0.006328f
C20 A1 a_452_68# 0.001247f
C21 a_276_68# ZN 0.007178f
C22 VNW VDD 0.172362f
C23 A2 VSS 0.130985f
C24 A2 A3 1.13496f
C25 VSS VDD 0.009236f
C26 VSS a_860_68# 0.005864f
C27 VSS a_452_68# 0.003244f
C28 a_276_68# VSS 0.003438f
C29 A3 VDD 0.099291f
C30 A2 VDD 0.041181f
C31 A2 a_860_68# 0.003842f
C32 VSS VPW 0.511432f
C33 ZN VPW 0.112753f
C34 VDD VPW 0.407724f
C35 A1 VPW 0.540441f
C36 A2 VPW 0.524145f
C37 A3 VPW 0.582222f
C38 VNW VPW 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW a_692_473#
+ a_254_473# a_66_473# a_2700_473# a_1660_473# a_3220_473# a_1212_473# a_2180_473#
+ a_3740_473# a_1920_473#
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VPW nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
C0 a_66_473# a_3740_473# 0.028219f
C1 A1 VDD 0.055928f
C2 a_66_473# A2 0.182327f
C3 a_3220_473# a_66_473# 0.021354f
C4 a_1920_473# a_66_473# 0.023791f
C5 A1 VNW 0.553741f
C6 VDD a_1212_473# 0.014305f
C7 A2 VSS 0.076134f
C8 a_254_473# VDD 0.012952f
C9 A4 A3 1.96796f
C10 A2 a_3740_473# 0.010293f
C11 VDD A3 0.086829f
C12 A4 VDD 0.110338f
C13 VDD a_2180_473# 0.00368f
C14 A3 VNW 0.567739f
C15 A1 ZN 1.60655f
C16 A4 VNW 0.513548f
C17 VDD VNW 0.394018f
C18 a_1660_473# A3 0.0054f
C19 VDD a_1660_473# 0.008572f
C20 a_66_473# A1 0.077909f
C21 ZN A3 0.417545f
C22 a_2700_473# VDD 0.003457f
C23 A4 ZN 1.44735f
C24 ZN a_2180_473# 0.018904f
C25 VDD ZN 0.007051f
C26 A1 VSS 0.093176f
C27 a_66_473# a_1212_473# 0.018664f
C28 a_254_473# a_66_473# 0.016207f
C29 ZN VNW 0.038639f
C30 a_66_473# A3 1.66251f
C31 a_66_473# A4 0.100571f
C32 a_66_473# a_2180_473# 0.020817f
C33 A2 A1 2.13585f
C34 ZN a_1660_473# 0.00216f
C35 a_66_473# VDD 3.19476f
C36 a_66_473# VNW 0.040351f
C37 VSS A3 0.078892f
C38 A4 VSS 0.099821f
C39 a_2700_473# ZN 0.019492f
C40 VDD VSS 0.009708f
C41 a_66_473# a_1660_473# 0.035002f
C42 VDD a_692_473# 0.017923f
C43 A2 A3 0.0303f
C44 VDD a_3740_473# 0.003118f
C45 VSS VNW 0.006947f
C46 a_66_473# a_2700_473# 0.021497f
C47 A2 VDD 0.054912f
C48 a_3220_473# VDD 0.003326f
C49 a_1920_473# VDD 0.004058f
C50 a_66_473# ZN 0.956309f
C51 A2 VNW 0.584134f
C52 ZN VSS 4.39577f
C53 ZN a_3740_473# 0.004594f
C54 A2 ZN 2.14591f
C55 a_3220_473# ZN 0.019778f
C56 a_1920_473# ZN 0.017667f
C57 a_66_473# VSS 0.01197f
C58 a_66_473# a_692_473# 0.022803f
C59 VSS VPW 1.3434f
C60 ZN VPW 0.240026f
C61 VDD VPW 0.844436f
C62 A1 VPW 1.40024f
C63 A2 VPW 1.30271f
C64 A4 VPW 1.33565f
C65 A3 VPW 1.29175f
C66 VNW VPW 6.70706f
C67 a_66_473# VPW 0.11665f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VNW VPW a_49_472# a_1133_69#
+ a_741_69#
X0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VPW nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VPW nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
C0 ZN A2 0.800412f
C1 a_49_472# VSS 0.01207f
C2 a_741_69# VSS 0.002035f
C3 VNW a_49_472# 0.012852f
C4 VNW VSS 0.0086f
C5 a_49_472# A1 0.03417f
C6 ZN a_1133_69# 0.001193f
C7 A1 VSS 0.129775f
C8 VNW A1 0.241301f
C9 VDD a_49_472# 1.09818f
C10 VDD VSS 0.009099f
C11 VNW VDD 0.151549f
C12 VDD A1 0.028601f
C13 B a_49_472# 0.234399f
C14 B VSS 0.061328f
C15 VNW B 0.260678f
C16 B VDD 0.045174f
C17 A2 a_49_472# 0.086717f
C18 a_741_69# A2 0.001142f
C19 A2 VSS 0.047574f
C20 VNW A2 0.272677f
C21 A2 A1 0.809974f
C22 ZN a_49_472# 0.475008f
C23 a_1133_69# VSS 0.00441f
C24 ZN a_741_69# 0.006341f
C25 ZN VSS 0.784804f
C26 A2 VDD 0.029358f
C27 ZN VNW 0.025755f
C28 a_1133_69# A1 0.003427f
C29 ZN A1 0.182845f
C30 ZN VDD 0.008463f
C31 B A2 0.029994f
C32 ZN B 0.20884f
C33 VSS VPW 0.510011f
C34 ZN VPW 0.070911f
C35 VDD VPW 0.327438f
C36 A1 VPW 0.556927f
C37 A2 VPW 0.56333f
C38 B VPW 0.662515f
C39 VNW VPW 2.52991f
C40 a_49_472# VPW 0.098072f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 ZN VSS 0.179304f
C1 VNW VSS 0.010163f
C2 VNW ZN 0.027829f
C3 VDD I 0.074838f
C4 VSS I 0.091531f
C5 ZN I 0.58604f
C6 VNW I 0.285482f
C7 VDD VSS 0.023187f
C8 ZN VDD 0.266247f
C9 VNW VDD 0.097124f
C10 VSS VPW 0.308828f
C11 ZN VPW 0.100523f
C12 VDD VPW 0.240805f
C13 I VPW 0.610668f
C14 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VNW VPW a_448_472#
+ a_36_151# a_1293_527# a_3081_151# a_1284_156# a_1040_527# a_1353_112# a_836_156#
+ a_1697_156# a_2449_156# a_3129_107# a_2225_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VPW nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VPW nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VPW nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VPW nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VPW nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VPW nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
C0 SETN VDD 0.127822f
C1 VDD a_1353_112# 0.016257f
C2 VDD a_2449_156# 0.208631f
C3 VNW a_2225_156# 0.209033f
C4 VNW D 0.1615f
C5 SETN a_2225_156# 0.070597f
C6 a_2225_156# a_1353_112# 0.152869f
C7 VNW SETN 0.811046f
C8 VNW a_1353_112# 0.219511f
C9 a_2449_156# a_2225_156# 0.569174f
C10 VDD a_36_151# 1.41468f
C11 VNW a_2449_156# 0.043816f
C12 VSS CLK 0.021941f
C13 a_448_472# a_1697_156# 0.007618f
C14 VSS a_3129_107# 0.136769f
C15 a_448_472# CLK 0.001313f
C16 a_2225_156# a_3081_151# 0.004129f
C17 SETN a_1353_112# 0.072983f
C18 a_1040_527# VDD 0.039677f
C19 SETN a_2449_156# 0.302222f
C20 a_2225_156# a_36_151# 0.153684f
C21 a_836_156# VSS 0.050008f
C22 a_448_472# VSS 1.07431f
C23 VNW a_36_151# 0.909435f
C24 a_448_472# a_836_156# 0.427756f
C25 a_2449_156# a_3081_151# 0.001203f
C26 a_36_151# D 0.092705f
C27 SETN a_36_151# 0.077775f
C28 a_36_151# a_1353_112# 0.840879f
C29 VNW a_1040_527# 0.223863f
C30 a_2449_156# a_36_151# 0.005967f
C31 SETN a_1040_527# 0.063241f
C32 a_1040_527# a_1353_112# 0.387423f
C33 Q a_3129_107# 0.179468f
C34 VSS Q 0.131272f
C35 VDD CLK 0.022091f
C36 VDD a_3129_107# 0.351307f
C37 a_1040_527# a_36_151# 0.206392f
C38 VSS VDD 0.013814f
C39 a_448_472# VDD 0.624585f
C40 a_2225_156# a_3129_107# 0.514036f
C41 VNW CLK 0.136589f
C42 VNW a_3129_107# 0.323464f
C43 a_1697_156# a_1353_112# 0.002752f
C44 VSS a_2225_156# 1.18908f
C45 a_448_472# a_2225_156# 0.153996f
C46 VNW VSS 0.009462f
C47 SETN a_3129_107# 0.089288f
C48 a_836_156# VNW 0.01368f
C49 a_448_472# VNW 0.400964f
C50 a_2449_156# a_3129_107# 0.00955f
C51 VSS D 0.067877f
C52 a_836_156# D 0.108102f
C53 a_448_472# D 0.400104f
C54 SETN VSS 0.008083f
C55 VSS a_1353_112# 0.027348f
C56 a_448_472# SETN 0.083903f
C57 a_448_472# a_1353_112# 0.317251f
C58 a_448_472# a_2449_156# 0.056679f
C59 a_36_151# CLK 0.700974f
C60 VDD Q 0.282179f
C61 a_36_151# a_1293_527# 0.008379f
C62 VSS a_36_151# 0.286331f
C63 a_836_156# a_36_151# 0.015697f
C64 a_448_472# a_36_151# 0.473132f
C65 a_1040_527# a_1293_527# 0.00215f
C66 VNW Q 0.031621f
C67 a_1040_527# VSS 0.060221f
C68 a_836_156# a_1040_527# 0.068207f
C69 a_448_472# a_1040_527# 0.869605f
C70 VDD a_2225_156# 0.073415f
C71 VSS a_1284_156# 0.003637f
C72 VNW VDD 0.539099f
C73 a_448_472# a_1284_156# 0.002691f
C74 VDD D 0.004944f
C75 Q VPW 0.105566f
C76 VSS VPW 1.35707f
C77 SETN VPW 0.710246f
C78 D VPW 0.247102f
C79 VDD VPW 0.833181f
C80 CLK VPW 0.290467f
C81 VNW VPW 6.44257f
C82 a_2449_156# VPW 0.049992f
C83 a_2225_156# VPW 0.434082f
C84 a_3129_107# VPW 0.58406f
C85 a_836_156# VPW 0.019766f
C86 a_1040_527# VPW 0.302082f
C87 a_1353_112# VPW 0.286513f
C88 a_448_472# VPW 1.21246f
C89 a_36_151# VPW 1.31409f
.ends

.subckt sarlogic cal clk clkc comp ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5]
+ ctln[6] ctln[7] ctln[8] ctln[9] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5]
+ ctlp[6] ctlp[7] ctlp[8] ctlp[9] en result[0] result[1] result[2] result[3] result[4]
+ result[5] result[6] result[7] result[8] result[9] rstn sample trim[0] trim[1] trim[2]
+ trim[3] trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] valid vdd vss _000_
+ _001_ _002_ _003_ _004_ _005_ _006_ _007_ _008_ _009_ _010_ _011_ _012_ _013_ _014_
+ _015_ _016_ _017_ _018_ _019_ _020_ _021_ _022_ _023_ _024_ _025_ _026_ _027_ _028_
+ _029_ _030_ _031_ _032_ _033_ _034_ _035_ _036_ _037_ _038_ _039_ _040_ _041_ _042_
+ _043_ _044_ _045_ _046_ _047_ _048_ _049_ _050_ _051_ _052_ _053_ _054_ _055_ _056_
+ _057_ _058_ _059_ _060_ _061_ _062_ _063_ _064_ _065_ _066_ _067_ _068_ _069_ _070_
+ _071_ _072_ _073_ _074_ _075_ _076_ _077_ _078_ _079_ _080_ _081_ _082_ _083_ _084_
+ _085_ _086_ _087_ _088_ _089_ _090_ _091_ _092_ _093_ _094_ _095_ _096_ _097_ _098_
+ _099_ _100_ _101_ _102_ _103_ _104_ _105_ _106_ _107_ _108_ _109_ _110_ _111_ _112_
+ _113_ _114_ _115_ _116_ _117_ _118_ _119_ _120_ _121_ _122_ _123_ _124_ _125_ _126_
+ _127_ _128_ _129_ _130_ _131_ _132_ _133_ _134_ _135_ _136_ _137_ _138_ _139_ _140_
+ _141_ _142_ _143_ _144_ _145_ _146_ _147_ _148_ _149_ _150_ _151_ _152_ _153_ _154_
+ _155_ _156_ _157_ _158_ _159_ _160_ _161_ _162_ _163_ _164_ _165_ _166_ _167_ _168_
+ _169_ _170_ _171_ _172_ _173_ _174_ _175_ _176_ _177_ _178_ _179_ _180_ _181_ _182_
+ _183_ _184_ _185_ _186_ _187_ _188_ cal_count\[0\] cal_count\[1\] cal_count\[2\]
+ cal_count\[3\] cal_itt\[0\] cal_itt\[1\] cal_itt\[2\] cal_itt\[3\] calibrate en_co_clk
+ mask\[0\] mask\[1\] mask\[2\] mask\[3\] mask\[4\] mask\[5\] mask\[6\] mask\[7\]
+ mask\[8\] mask\[9\] net1 net10 net11 net12 net13 net14 net15 net16 net17 net18 net19
+ net2 net20 net21 net22 net23 net24 net25 net26 net27 net28 net29 net3 net30 net31
+ net32 net33 net34 net35 net36 net37 net38 net39 net4 net40 net41 net42 net43 net44
+ net45 net46 net47 net48 net49 net5 net50 net51 net52 net53 net54 net55 net56 net57
+ net58 net59 net6 net60 net61 net62 net63 net64 net65 net66 net67 net68 net69 net7
+ net70 net71 net72 net73 net74 net75 net76 net77 net78 net79 net8 net80 net81 net82
+ net9 state\[0\] state\[1\] state\[2\] trim_mask\[0\] trim_mask\[1\] trim_mask\[2\]
+ trim_mask\[3\] trim_mask\[4\] trim_val\[0\] trim_val\[1\] trim_val\[2\] trim_val\[3\]
+ trim_val\[4\]
XFILLER_0_17_200 vdd vss vdd vss FILLER_0_17_200/a_36_472# FILLER_0_17_200/a_572_375#
+ FILLER_0_17_200/a_124_375# FILLER_0_17_200/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_294_ vdd vss _008_ _104_ _106_ vdd vss _294_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_432_ _021_ mask\[3\] net63 vss net80 vdd vdd vss _432_/a_2665_112# _432_/a_448_472#
+ _432_/a_796_472# _432_/a_36_151# _432_/a_1204_472# _432_/a_3041_156# _432_/a_1000_472#
+ _432_/a_1308_423# _432_/a_1456_156# _432_/a_1288_156# _432_/a_2248_156# _432_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ vdd vss _363_/a_36_68# _363_/a_244_472#
+ _363_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ vdd vss _346_/a_49_472# _346_/a_665_69#
+ _346_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd vdd vss _415_/a_2665_112# _415_/a_448_472#
+ _415_/a_796_472# _415_/a_36_151# _415_/a_1204_472# _415_/a_3041_156# _415_/a_1000_472#
+ _415_/a_1308_423# _415_/a_1456_156# _415_/a_1288_156# _415_/a_2248_156# _415_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd vdd vss _277_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss vdd vss FILLER_0_19_125/a_36_472# FILLER_0_19_125/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss vdd vss FILLER_0_15_150/a_36_472# FILLER_0_15_150/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss vdd vss FILLER_0_21_142/a_36_472# FILLER_0_21_142/a_572_375#
+ FILLER_0_21_142/a_124_375# FILLER_0_21_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss vdd vss FILLER_0_16_73/a_36_472# FILLER_0_16_73/a_572_375#
+ FILLER_0_16_73/a_124_375# FILLER_0_16_73/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss vdd vss output20/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss vdd vss output31/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss vdd vss output42/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 ctln[0] net7 vdd vss vdd vss output7/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss vdd vss FILLER_0_5_117/a_36_472# FILLER_0_5_117/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss vdd vss FILLER_0_5_128/a_36_472# FILLER_0_5_128/a_572_375#
+ FILLER_0_5_128/a_124_375# FILLER_0_5_128/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_293_ net31 vdd vss _106_ mask\[4\] _105_ vdd vss _293_/a_36_472# _293_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_431_ _020_ mask\[2\] net53 vss net70 vdd vdd vss _431_/a_2665_112# _431_/a_448_472#
+ _431_/a_796_472# _431_/a_36_151# _431_/a_1204_472# _431_/a_3041_156# _431_/a_1000_472#
+ _431_/a_1308_423# _431_/a_1456_156# _431_/a_1288_156# _431_/a_2248_156# _431_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_362_ vdd vss trim_mask\[1\] _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_345_ vss _144_ _132_ vdd vdd vss _345_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ vss _093_ _092_ vdd vdd vss _276_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd vdd vss _414_/a_2665_112# _414_/a_448_472#
+ _414_/a_796_472# _414_/a_36_151# _414_/a_1204_472# _414_/a_3041_156# _414_/a_1000_472#
+ _414_/a_1308_423# _414_/a_1456_156# _414_/a_1288_156# _414_/a_2248_156# _414_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd vdd vss _328_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss vdd vss FILLER_0_9_28/a_1916_375# FILLER_0_9_28/a_1380_472#
+ FILLER_0_9_28/a_3260_375# FILLER_0_9_28/a_36_472# FILLER_0_9_28/a_932_472# FILLER_0_9_28/a_2812_375#
+ FILLER_0_9_28/a_2276_472# FILLER_0_9_28/a_1828_472# FILLER_0_9_28/a_3172_472# FILLER_0_9_28/a_572_375#
+ FILLER_0_9_28/a_2724_472# FILLER_0_9_28/a_124_375# FILLER_0_9_28/a_1468_375# FILLER_0_9_28/a_1020_375#
+ FILLER_0_9_28/a_484_472# FILLER_0_9_28/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_204 vdd vss vdd vss FILLER_0_3_204/a_36_472# FILLER_0_3_204/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _078_ vdd vss _080_ _073_ _076_ vdd vss _259_/a_455_68# _259_/a_271_68# gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd vss vdd vss FILLER_0_16_107/a_36_472# FILLER_0_16_107/a_572_375#
+ FILLER_0_16_107/a_124_375# FILLER_0_16_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss vdd vss output21/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss vdd vss output43/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss vdd vss output32/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss vdd vss output10/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss vdd vss output8/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ vss _105_ _098_ vdd vdd vss _292_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_430_ _019_ mask\[1\] net63 vss net80 vdd vdd vss _430_/a_2665_112# _430_/a_448_472#
+ _430_/a_796_472# _430_/a_36_151# _430_/a_1204_472# _430_/a_3041_156# _430_/a_1000_472#
+ _430_/a_1308_423# _430_/a_1456_156# _430_/a_1288_156# _430_/a_2248_156# _430_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_361_ vdd vss _154_ _086_ _119_ vdd vss _361_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss vdd vss FILLER_0_7_72/a_1916_375# FILLER_0_7_72/a_1380_472#
+ FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472# FILLER_0_7_72/a_932_472# FILLER_0_7_72/a_2812_375#
+ FILLER_0_7_72/a_2276_472# FILLER_0_7_72/a_1828_472# FILLER_0_7_72/a_3172_472# FILLER_0_7_72/a_572_375#
+ FILLER_0_7_72/a_2724_472# FILLER_0_7_72/a_124_375# FILLER_0_7_72/a_1468_375# FILLER_0_7_72/a_1020_375#
+ FILLER_0_7_72/a_484_472# FILLER_0_7_72/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ vdd vss _275_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__191__I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd vdd vss _413_/a_2665_112# _413_/a_448_472#
+ _413_/a_796_472# _413_/a_36_151# _413_/a_1204_472# _413_/a_3041_156# _413_/a_1000_472#
+ _413_/a_1308_423# _413_/a_1456_156# _413_/a_1288_156# _413_/a_2248_156# _413_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_96 vdd vss vdd vss FILLER_0_24_96/a_36_472# FILLER_0_24_96/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss vdd vss FILLER_0_24_63/a_36_472# FILLER_0_24_63/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ vdd vss _043_ net27 mask\[0\] vdd vss _189_/a_255_603# _189_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_327_ _131_ vdd vss _016_ _127_ _130_ vdd vss _327_/a_36_472# _327_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ vss _079_ _078_ vdd vdd vss _258_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss vdd vss FILLER_0_18_171/a_36_472# FILLER_0_18_171/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss vdd vss FILLER_0_24_130/a_36_472# FILLER_0_24_130/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss vdd vss FILLER_0_21_133/a_36_472# FILLER_0_21_133/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss vdd vss FILLER_0_8_138/a_36_472# FILLER_0_8_138/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss vdd vss FILLER_0_8_127/a_36_472# FILLER_0_8_127/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 ctlp[5] net22 vdd vss vdd vss output22/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 result[6] net33 vdd vss vdd vss output33/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss vdd vss output44/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss vdd vss output11/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss vdd vss output9/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd vdd vss _291_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss vdd vss FILLER_0_4_152/a_36_472# FILLER_0_4_152/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss vdd vss FILLER_0_4_185/a_36_472# FILLER_0_4_185/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd vdd vss _360_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss vdd vss FILLER_0_13_65/a_36_472# FILLER_0_13_65/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ vdd vss _343_/a_49_472# _343_/a_665_69#
+ _343_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ vdd vss _274_/a_36_68# _274_/a_1612_497#
+ _274_/a_2124_68# _274_/a_244_497# _274_/a_2960_68# _274_/a_3368_68# _274_/a_2552_68#
+ _274_/a_1164_497# _274_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd vdd vss _412_/a_2665_112# _412_/a_448_472#
+ _412_/a_796_472# _412_/a_36_151# _412_/a_1204_472# _412_/a_3041_156# _412_/a_1000_472#
+ _412_/a_1308_423# _412_/a_1456_156# _412_/a_1288_156# _412_/a_2248_156# _412_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__292__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ vdd vss _326_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ vdd vss _257_/a_36_472# _257_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__301__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss vdd vss FILLER_0_15_142/a_36_472# FILLER_0_15_142/a_572_375#
+ FILLER_0_15_142/a_124_375# FILLER_0_15_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 ctlp[6] net23 vdd vss vdd vss output23/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss vdd vss output45/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss vdd vss output34/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss vdd vss output12/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss vdd vss FILLER_0_5_109/a_36_472# FILLER_0_5_109/a_572_375#
+ FILLER_0_5_109/a_124_375# FILLER_0_5_109/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss vdd vss FILLER_0_17_226/a_36_472# FILLER_0_17_226/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss vdd vss FILLER_0_4_197/a_1380_472# FILLER_0_4_197/a_36_472#
+ FILLER_0_4_197/a_932_472# FILLER_0_4_197/a_572_375# FILLER_0_4_197/a_124_375# FILLER_0_4_197/a_1468_375#
+ FILLER_0_4_197/a_1020_375# FILLER_0_4_197/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ vdd vss _290_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss vdd vss FILLER_0_9_223/a_36_472# FILLER_0_9_223/a_572_375#
+ FILLER_0_9_223/a_124_375# FILLER_0_9_223/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_273_ vss _090_ state\[0\] vdd vdd vss _273_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd vdd vss _411_/a_2665_112# _411_/a_448_472#
+ _411_/a_796_472# _411_/a_36_151# _411_/a_1204_472# _411_/a_3041_156# _411_/a_1000_472#
+ _411_/a_1308_423# _411_/a_1456_156# _411_/a_1288_156# _411_/a_2248_156# _411_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout80 vss net80 net81 vdd vdd vss fanout80/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_325_ vdd vss _130_ _118_ _129_ vdd vss _325_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd vss vdd vss FILLER_0_10_78/a_1380_472# FILLER_0_10_78/a_36_472#
+ FILLER_0_10_78/a_932_472# FILLER_0_10_78/a_572_375# FILLER_0_10_78/a_124_375# FILLER_0_10_78/a_1468_375#
+ FILLER_0_10_78/a_1020_375# FILLER_0_10_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ vdd vss _256_/a_36_68# _256_/a_1612_497#
+ _256_/a_2124_68# _256_/a_244_497# _256_/a_2960_68# _256_/a_3368_68# _256_/a_2552_68#
+ _256_/a_1164_497# _256_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ vdd vss _308_/a_848_380# _308_/a_1084_68#
+ _308_/a_124_24# _308_/a_1152_472# _308_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss vdd vss FILLER_0_1_98/a_36_472# FILLER_0_1_98/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ vdd vss _239_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss vdd vss FILLER_0_12_124/a_36_472# FILLER_0_12_124/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss vdd vss FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 ctlp[7] net24 vdd vss vdd vss output24/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss vdd vss output35/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss vdd vss output46/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss vdd vss FILLER_0_18_2/a_1916_375# FILLER_0_18_2/a_1380_472#
+ FILLER_0_18_2/a_3260_375# FILLER_0_18_2/a_36_472# FILLER_0_18_2/a_932_472# FILLER_0_18_2/a_2812_375#
+ FILLER_0_18_2/a_2276_472# FILLER_0_18_2/a_1828_472# FILLER_0_18_2/a_3172_472# FILLER_0_18_2/a_572_375#
+ FILLER_0_18_2/a_2724_472# FILLER_0_18_2/a_124_375# FILLER_0_18_2/a_1468_375# FILLER_0_18_2/a_1020_375#
+ FILLER_0_18_2/a_484_472# FILLER_0_18_2/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 ctln[6] net13 vdd vss vdd vss output13/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss vdd vss FILLER_0_7_162/a_36_472# FILLER_0_7_162/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss vdd vss FILLER_0_7_195/a_36_472# FILLER_0_7_195/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ vdd vss _341_/a_49_472# _341_/a_665_69#
+ _341_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss vdd vss _410_/a_36_68# _410_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ vdd vss _272_/a_36_472# _272_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd vdd vss fanout70/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ _076_ vss vdd _057_ vdd vss _255_/a_224_552# gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_324_ vdd vss _129_ calibrate _062_ vdd vss _324_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output40_I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 vss net81 net82 vdd vdd vss fanout81/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_55 vdd vss vdd vss FILLER_0_19_55/a_36_472# FILLER_0_19_55/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_307_ vdd vss _114_ _113_ _096_ vdd vss _307_/a_234_472# _307_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] vdd vss _238_/a_255_603# _238_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss vdd vss FILLER_0_21_125/a_36_472# FILLER_0_21_125/a_572_375#
+ FILLER_0_21_125/a_124_375# FILLER_0_21_125/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss vdd vss FILLER_0_16_89/a_1380_472# FILLER_0_16_89/a_36_472#
+ FILLER_0_16_89/a_932_472# FILLER_0_16_89/a_572_375# FILLER_0_16_89/a_124_375# FILLER_0_16_89/a_1468_375#
+ FILLER_0_16_89/a_1020_375# FILLER_0_16_89/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss vdd vss FILLER_0_12_136/a_1380_472# FILLER_0_12_136/a_36_472#
+ FILLER_0_12_136/a_932_472# FILLER_0_12_136/a_572_375# FILLER_0_12_136/a_124_375#
+ FILLER_0_12_136/a_1468_375# FILLER_0_12_136/a_1020_375# FILLER_0_12_136/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 ctlp[8] net25 vdd vss vdd vss output25/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss vdd vss output47/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 result[9] net36 vdd vss vdd vss output36/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss vdd vss output14/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss vdd vss FILLER_0_4_144/a_36_472# FILLER_0_4_144/a_572_375#
+ FILLER_0_4_144/a_124_375# FILLER_0_4_144/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss vdd vss FILLER_0_4_177/a_36_472# FILLER_0_4_177/a_572_375#
+ FILLER_0_4_177/a_124_375# FILLER_0_4_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd vdd vss _340_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss vdd vss FILLER_0_10_256/a_36_472# FILLER_0_10_256/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__200__I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_99 vdd vss vdd vss FILLER_0_4_99/a_36_472# FILLER_0_4_99/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss vdd vss FILLER_0_6_239/a_36_472# FILLER_0_6_239/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout71 vss net71 net73 vdd vdd vss fanout71/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 net60 vss vdd net61 vdd vss fanout60/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_323_ vss _015_ _128_ vdd vdd vss _323_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd vdd vss fanout82/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ vdd vss _254_/a_448_472# _254_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_237_ vdd vss net40 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_306_ vss _113_ _057_ vdd vdd vss _306_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_57 vdd vss vdd vss FILLER_0_16_57/a_1380_472# FILLER_0_16_57/a_36_472#
+ FILLER_0_16_57/a_932_472# FILLER_0_16_57/a_572_375# FILLER_0_16_57/a_124_375# FILLER_0_16_57/a_1468_375#
+ FILLER_0_16_57/a_1020_375# FILLER_0_16_57/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss vdd vss output26/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss vdd vss output15/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss vdd vss output37/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss vdd vss output48/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss vdd vss FILLER_0_17_218/a_36_472# FILLER_0_17_218/a_572_375#
+ FILLER_0_17_218/a_124_375# FILLER_0_17_218/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss vdd vss FILLER_0_4_123/a_36_472# FILLER_0_4_123/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ vdd vss _270_/a_36_472# _270_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ vdd vss _399_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ vdd vss _322_/a_848_380# _322_/a_1084_68# _322_/a_124_24#
+ _322_/a_1152_472# _322_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd vdd vss fanout61/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd vdd vss fanout72/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd vss vdd vss FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net50 vss vdd net52 vdd vss fanout50/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] vdd vss _253_/a_36_68#
+ _253_/a_1732_68# _253_/a_244_68# _253_/a_1100_68# _253_/a_1528_68# _253_/a_672_68#
+ gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_305_ vdd vss _112_ net1 _081_ vdd vss _305_/a_36_159# gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ net40 vss vdd _064_ vdd vss _236_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss vdd vss FILLER_0_20_193/a_36_472# FILLER_0_20_193/a_572_375#
+ FILLER_0_20_193/a_124_375# FILLER_0_20_193/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd vdd vss _219_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss vdd vss output27/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss vdd vss output16/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss vdd vss output38/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss vdd vss FILLER_0_16_241/a_36_472# FILLER_0_16_241/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd vdd vss _398_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vss vdd vss FILLER_0_10_247/a_36_472# FILLER_0_10_247/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_214 vdd vss vdd vss FILLER_0_10_214/a_36_472# FILLER_0_10_214/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_91 vdd vss vdd vss FILLER_0_14_91/a_36_472# FILLER_0_14_91/a_572_375#
+ FILLER_0_14_91/a_124_375# FILLER_0_14_91/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__209__I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss vdd vss FILLER_0_19_47/a_36_472# FILLER_0_19_47/a_572_375#
+ FILLER_0_19_47/a_124_375# FILLER_0_19_47/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd vdd vss fanout73/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 net62 vss vdd net64 vdd vss fanout62/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vss net51 net52 vdd vdd vss fanout51/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ vdd vss _321_/a_2590_472# _321_/a_170_472#
+ _321_/a_1602_69# _321_/a_786_69# _321_/a_3126_472# _321_/a_1194_69# _321_/a_3662_472#
+ _321_/a_2034_472# _321_/a_358_69# gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_252_ vdd vss cal_itt\[0\] _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_100 vdd vss vdd vss FILLER_0_18_100/a_36_472# FILLER_0_18_100/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss vdd vss FILLER_0_18_177/a_1916_375# FILLER_0_18_177/a_1380_472#
+ FILLER_0_18_177/a_3260_375# FILLER_0_18_177/a_36_472# FILLER_0_18_177/a_932_472#
+ FILLER_0_18_177/a_2812_375# FILLER_0_18_177/a_2276_472# FILLER_0_18_177/a_1828_472#
+ FILLER_0_18_177/a_3172_472# FILLER_0_18_177/a_572_375# FILLER_0_18_177/a_2724_472#
+ FILLER_0_18_177/a_124_375# FILLER_0_18_177/a_1468_375# FILLER_0_18_177/a_1020_375#
+ FILLER_0_18_177/a_484_472# FILLER_0_18_177/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ vdd vss _304_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] vdd vss _235_/a_255_603# _235_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss vdd vss FILLER_0_16_37/a_36_472# FILLER_0_16_37/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss vdd vss output17/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss vdd vss output28/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss vdd vss output39/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss vdd vss FILLER_0_13_212/a_1380_472# FILLER_0_13_212/a_36_472#
+ FILLER_0_13_212/a_932_472# FILLER_0_13_212/a_572_375# FILLER_0_13_212/a_124_375#
+ FILLER_0_13_212/a_1468_375# FILLER_0_13_212/a_1020_375# FILLER_0_13_212/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ vdd vss _397_/a_36_472# _397_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss vdd vss FILLER_0_14_81/a_36_472# FILLER_0_14_81/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout63 net63 vss vdd net64 vdd vss fanout63/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ vdd vss _320_/a_1792_472# _320_/a_224_472#
+ _320_/a_1568_472# _320_/a_36_472# _320_/a_1120_472# _320_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_28 vdd vss vdd vss FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 vss net74 net82 vdd vdd vss fanout74/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net52 vss vdd net57 vdd vss fanout52/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ vdd vss _251_/a_468_472# _251_/a_244_472# _251_/a_1130_472#
+ _251_/a_906_472# gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_449_ _038_ en_co_clk net55 vss net72 vdd vdd vss _449_/a_2665_112# _449_/a_448_472#
+ _449_/a_796_472# _449_/a_36_151# _449_/a_1204_472# _449_/a_3041_156# _449_/a_1000_472#
+ _449_/a_1308_423# _449_/a_1456_156# _449_/a_1288_156# _449_/a_2248_156# _449_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ vdd vss _303_/a_36_472# _303_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_217_ vss net26 _052_ vdd vdd vss _217_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_181 vdd vss vdd vss FILLER_0_14_181/a_36_472# FILLER_0_14_181/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 ctlp[1] net18 vdd vss vdd vss output18/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss vdd vss output29/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ vdd vss _396_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout53 net53 vss vdd net56 vdd vss fanout53/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_250_ vss _072_ _071_ vdd vdd vss _250_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 vss net75 net76 vdd vdd vss fanout75/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd vdd vss fanout64/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd vdd vss _448_/a_2665_112# _448_/a_448_472#
+ _448_/a_796_472# _448_/a_36_151# _448_/a_1204_472# _448_/a_3041_156# _448_/a_1000_472#
+ _448_/a_1308_423# _448_/a_1456_156# _448_/a_1288_156# _448_/a_2248_156# _448_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ vdd vss _379_/a_36_472# _379_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_302_ vdd vss _012_ _093_ _110_ vdd vss _302_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss vdd vss FILLER_0_21_28/a_1916_375# FILLER_0_21_28/a_1380_472#
+ FILLER_0_21_28/a_3260_375# FILLER_0_21_28/a_36_472# FILLER_0_21_28/a_932_472# FILLER_0_21_28/a_2812_375#
+ FILLER_0_21_28/a_2276_472# FILLER_0_21_28/a_1828_472# FILLER_0_21_28/a_3172_472#
+ FILLER_0_21_28/a_572_375# FILLER_0_21_28/a_2724_472# FILLER_0_21_28/a_124_375# FILLER_0_21_28/a_1468_375#
+ FILLER_0_21_28/a_1020_375# FILLER_0_21_28/a_484_472# FILLER_0_21_28/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__216__A2 vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ vss net39 _063_ vdd vdd vss _233_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss vdd vss FILLER_0_15_116/a_36_472# FILLER_0_15_116/a_572_375#
+ FILLER_0_15_116/a_124_375# FILLER_0_15_116/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_216_ vdd vss _052_ mask\[9\] net36 vdd vss _216_/a_255_603# _216_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_146 vdd vss vdd vss FILLER_0_7_146/a_36_472# FILLER_0_7_146/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 ctlp[2] net19 vdd vss vdd vss output19/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss vdd vss FILLER_0_7_59/a_36_472# FILLER_0_7_59/a_572_375# FILLER_0_7_59/a_124_375#
+ FILLER_0_7_59/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss vdd vss FILLER_0_16_255/a_36_472# FILLER_0_16_255/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss vdd vss FILLER_0_0_130/a_36_472# FILLER_0_0_130/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss vdd vss FILLER_0_8_263/a_36_472# FILLER_0_8_263/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss vdd vss FILLER_0_14_50/a_36_472# FILLER_0_14_50/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ vdd vss _395_/a_1492_488# _395_/a_244_68#
+ _395_/a_1044_488# _395_/a_636_68# _395_/a_36_488# gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss vdd vss FILLER_0_4_49/a_36_472# FILLER_0_4_49/a_572_375# FILLER_0_4_49/a_124_375#
+ FILLER_0_4_49/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 vdd vss fanout54/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd vdd vss fanout76/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd vdd vss fanout65/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss vdd vss FILLER_0_19_28/a_36_472# FILLER_0_19_28/a_572_375#
+ FILLER_0_19_28/a_124_375# FILLER_0_19_28/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd vdd vss _447_/a_2665_112# _447_/a_448_472#
+ _447_/a_796_472# _447_/a_36_151# _447_/a_1204_472# _447_/a_3041_156# _447_/a_1000_472#
+ _447_/a_1308_423# _447_/a_1456_156# _447_/a_1288_156# _447_/a_2248_156# _447_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_2 vdd vss vdd vss FILLER_0_3_2/a_36_472# FILLER_0_3_2/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ vdd vss _033_ _160_ _165_ vdd vss _378_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ vdd vss _301_/a_36_472# _301_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] vdd vss _232_/a_255_603# _232_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss vdd vss FILLER_0_11_142/a_36_472# FILLER_0_11_142/a_572_375#
+ FILLER_0_11_142/a_124_375# FILLER_0_11_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss vdd vss FILLER_0_2_93/a_36_472# FILLER_0_2_93/a_572_375# FILLER_0_2_93/a_124_375#
+ FILLER_0_2_93/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss vdd vss FILLER_0_17_72/a_1916_375# FILLER_0_17_72/a_1380_472#
+ FILLER_0_17_72/a_3260_375# FILLER_0_17_72/a_36_472# FILLER_0_17_72/a_932_472# FILLER_0_17_72/a_2812_375#
+ FILLER_0_17_72/a_2276_472# FILLER_0_17_72/a_1828_472# FILLER_0_17_72/a_3172_472#
+ FILLER_0_17_72/a_572_375# FILLER_0_17_72/a_2724_472# FILLER_0_17_72/a_124_375# FILLER_0_17_72/a_1468_375#
+ FILLER_0_17_72/a_1020_375# FILLER_0_17_72/a_484_472# FILLER_0_17_72/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss vdd vss FILLER_0_3_172/a_1916_375# FILLER_0_3_172/a_1380_472#
+ FILLER_0_3_172/a_3260_375# FILLER_0_3_172/a_36_472# FILLER_0_3_172/a_932_472# FILLER_0_3_172/a_2812_375#
+ FILLER_0_3_172/a_2276_472# FILLER_0_3_172/a_1828_472# FILLER_0_3_172/a_3172_472#
+ FILLER_0_3_172/a_572_375# FILLER_0_3_172/a_2724_472# FILLER_0_3_172/a_124_375# FILLER_0_3_172/a_1468_375#
+ FILLER_0_3_172/a_1020_375# FILLER_0_3_172/a_484_472# FILLER_0_3_172/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] vdd vss _394_/a_244_524# _394_/a_2215_68#
+ _394_/a_56_524# _394_/a_718_524# _394_/a_728_93# _394_/a_1936_472# _394_/a_1336_472#
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 vdd vss fanout55/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss vdd vss FILLER_0_5_212/a_36_472# FILLER_0_5_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd vdd vss fanout77/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd vdd vss _446_/a_2665_112# _446_/a_448_472#
+ _446_/a_796_472# _446_/a_36_151# _446_/a_1204_472# _446_/a_3041_156# _446_/a_1000_472#
+ _446_/a_1308_423# _446_/a_1456_156# _446_/a_1288_156# _446_/a_2248_156# _446_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout66 vss net66 net68 vdd vdd vss fanout66/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ vdd vss _377_/a_36_472# _377_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd vss _011_ _104_ _109_ vdd vss _300_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ vdd vss _231_/a_652_68# _231_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd vdd vss _429_/a_2665_112# _429_/a_448_472#
+ _429_/a_796_472# _429_/a_36_151# _429_/a_1204_472# _429_/a_3041_156# _429_/a_1000_472#
+ _429_/a_1308_423# _429_/a_1456_156# _429_/a_1288_156# _429_/a_2248_156# _429_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd vdd vss input1/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd vdd vss _214_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss vdd vss FILLER_0_7_104/a_1380_472# FILLER_0_7_104/a_36_472#
+ FILLER_0_7_104/a_932_472# FILLER_0_7_104/a_572_375# FILLER_0_7_104/a_124_375# FILLER_0_7_104/a_1468_375#
+ FILLER_0_7_104/a_1020_375# FILLER_0_7_104/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss vdd vss FILLER_0_4_107/a_1380_472# FILLER_0_4_107/a_36_472#
+ FILLER_0_4_107/a_932_472# FILLER_0_4_107/a_572_375# FILLER_0_4_107/a_124_375# FILLER_0_4_107/a_1468_375#
+ FILLER_0_4_107/a_1020_375# FILLER_0_4_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss vdd vss FILLER_0_24_290/a_36_472# FILLER_0_24_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss vdd vss FILLER_0_15_290/a_36_472# FILLER_0_15_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss vdd vss FILLER_0_0_198/a_36_472# FILLER_0_0_198/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd vdd vss fanout78/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd vdd vss fanout56/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd vdd vss fanout67/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd vdd vss _445_/a_2665_112# _445_/a_448_472#
+ _445_/a_796_472# _445_/a_36_151# _445_/a_1204_472# _445_/a_3041_156# _445_/a_1000_472#
+ _445_/a_1308_423# _445_/a_1456_156# _445_/a_1288_156# _445_/a_2248_156# _445_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vss _164_ _163_ vdd vdd vss _376_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd vss _062_ _060_ _061_ vdd vss _230_/a_652_68# _230_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vss vdd vss FILLER_0_5_72/a_1380_472# FILLER_0_5_72/a_36_472# FILLER_0_5_72/a_932_472#
+ FILLER_0_5_72/a_572_375# FILLER_0_5_72/a_124_375# FILLER_0_5_72/a_1468_375# FILLER_0_5_72/a_1020_375#
+ FILLER_0_5_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ _017_ state\[2\] net53 vss net70 vdd vdd vss _428_/a_2665_112# _428_/a_448_472#
+ _428_/a_796_472# _428_/a_36_151# _428_/a_1204_472# _428_/a_3041_156# _428_/a_1000_472#
+ _428_/a_1308_423# _428_/a_1456_156# _428_/a_1288_156# _428_/a_2248_156# _428_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd vss vdd vss FILLER_0_11_64/a_36_472# FILLER_0_11_64/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ vdd vss _359_/a_1492_488# _359_/a_244_68#
+ _359_/a_1044_488# _359_/a_636_68# _359_/a_36_488# gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vss net2 clk vdd vdd vss input2/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output22_I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 vdd vss _213_/a_255_603# _213_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_177 vdd vss vdd vss FILLER_0_20_177/a_1380_472# FILLER_0_20_177/a_36_472#
+ FILLER_0_20_177/a_932_472# FILLER_0_20_177/a_572_375# FILLER_0_20_177/a_124_375#
+ FILLER_0_20_177/a_1468_375# FILLER_0_20_177/a_1020_375# FILLER_0_20_177/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_206 vdd vss vdd vss FILLER_0_13_206/a_36_472# FILLER_0_13_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss vdd vss FILLER_0_13_228/a_36_472# FILLER_0_13_228/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss vdd vss _392_/a_36_68# _392_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__282__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 vss net79 net81 vdd vdd vss fanout79/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_2 vdd vss vdd vss FILLER_0_12_2/a_36_472# FILLER_0_12_2/a_572_375# FILLER_0_12_2/a_124_375#
+ FILLER_0_12_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout68 vss net68 net69 vdd vdd vss fanout68/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 vss net57 net65 vdd vdd vss fanout57/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd vdd vss _444_/a_2665_112# _444_/a_448_472#
+ _444_/a_796_472# _444_/a_36_151# _444_/a_1204_472# _444_/a_3041_156# _444_/a_1000_472#
+ _444_/a_1308_423# _444_/a_1456_156# _444_/a_1288_156# _444_/a_2248_156# _444_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] vdd vss _375_/a_36_68# _375_/a_1612_497#
+ _375_/a_692_497# _375_/a_1388_497# _375_/a_960_497# gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__277__I vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd vss vdd vss FILLER_0_18_139/a_1380_472# FILLER_0_18_139/a_36_472#
+ FILLER_0_18_139/a_932_472# FILLER_0_18_139/a_572_375# FILLER_0_18_139/a_124_375#
+ FILLER_0_18_139/a_1468_375# FILLER_0_18_139/a_1020_375# FILLER_0_18_139/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_161 vdd vss vdd vss FILLER_0_17_161/a_36_472# FILLER_0_17_161/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ _016_ state\[1\] net53 vdd vss net70 vdd vss _427_/a_2665_112# _427_/a_448_472#
+ _427_/a_796_472# _427_/a_36_151# _427_/a_1204_472# _427_/a_3041_156# _427_/a_1000_472#
+ _427_/a_1308_423# _427_/a_2248_156# _427_/a_2560_156# gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_358_ vdd vss _053_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ vdd vss _289_/a_36_472# _289_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd vdd vss input3/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss vdd vss FILLER_0_22_86/a_1380_472# FILLER_0_22_86/a_36_472#
+ FILLER_0_22_86/a_932_472# FILLER_0_22_86/a_572_375# FILLER_0_22_86/a_124_375# FILLER_0_22_86/a_1468_375#
+ FILLER_0_22_86/a_1020_375# FILLER_0_22_86/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss vdd vss FILLER_0_11_101/a_36_472# FILLER_0_11_101/a_572_375#
+ FILLER_0_11_101/a_124_375# FILLER_0_11_101/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss vdd vss FILLER_0_17_64/a_36_472# FILLER_0_17_64/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss vdd vss FILLER_0_3_142/a_36_472# FILLER_0_3_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ vdd vss _391_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 vss net69 net74 vdd vdd vss fanout69/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net58 vss vdd net59 vdd vss fanout58/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_374_ vdd _061_ _056_ _162_ calibrate vss vdd vss _374_/a_36_68# _374_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd vdd vss _443_/a_2665_112# _443_/a_448_472#
+ _443_/a_796_472# _443_/a_36_151# _443_/a_1204_472# _443_/a_3041_156# _443_/a_1000_472#
+ _443_/a_1308_423# _443_/a_1456_156# _443_/a_1288_156# _443_/a_2248_156# _443_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_107 vdd vss vdd vss FILLER_0_18_107/a_1916_375# FILLER_0_18_107/a_1380_472#
+ FILLER_0_18_107/a_3260_375# FILLER_0_18_107/a_36_472# FILLER_0_18_107/a_932_472#
+ FILLER_0_18_107/a_2812_375# FILLER_0_18_107/a_2276_472# FILLER_0_18_107/a_1828_472#
+ FILLER_0_18_107/a_3172_472# FILLER_0_18_107/a_572_375# FILLER_0_18_107/a_2724_472#
+ FILLER_0_18_107/a_124_375# FILLER_0_18_107/a_1468_375# FILLER_0_18_107/a_1020_375#
+ FILLER_0_18_107/a_484_472# FILLER_0_18_107/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ vdd vss _288_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ _015_ state\[0\] net64 vss net81 vdd vdd vss _426_/a_2665_112# _426_/a_448_472#
+ _426_/a_796_472# _426_/a_36_151# _426_/a_1204_472# _426_/a_3041_156# _426_/a_1000_472#
+ _426_/a_1308_423# _426_/a_1456_156# _426_/a_1288_156# _426_/a_2248_156# _426_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 vss net4 en vdd vdd vss input4/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_211_ vss net24 _050_ vdd vdd vss _211_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ vdd vss _409_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd vss vdd vss FILLER_0_11_135/a_36_472# FILLER_0_11_135/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vss vdd vss FILLER_0_11_124/a_36_472# FILLER_0_11_124/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss vdd vss FILLER_0_15_282/a_36_472# FILLER_0_15_282/a_572_375#
+ FILLER_0_15_282/a_124_375# FILLER_0_15_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ vdd vss _390_/a_36_68# _390_/a_244_472#
+ _390_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss vdd vss FILLER_0_14_99/a_36_472# FILLER_0_14_99/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 vdd vss fanout59/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ vdd vss _373_/a_438_68# _373_/a_244_68#
+ _373_/a_1254_68# _373_/a_1060_68# _373_/a_632_68# _373_/a_1458_68# gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd vdd vss _442_/a_2665_112# _442_/a_448_472#
+ _442_/a_796_472# _442_/a_36_151# _442_/a_1204_472# _442_/a_3041_156# _442_/a_1000_472#
+ _442_/a_1308_423# _442_/a_1456_156# _442_/a_1288_156# _442_/a_2248_156# _442_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ vdd vss _356_/a_36_472# _356_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ vdd vss _287_/a_36_472# _287_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss vdd vss FILLER_0_11_78/a_36_472# FILLER_0_11_78/a_572_375#
+ FILLER_0_11_78/a_124_375# FILLER_0_11_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd vdd vss input5/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd vdd vss _425_/a_2665_112# _425_/a_448_472#
+ _425_/a_796_472# _425_/a_36_151# _425_/a_1204_472# _425_/a_3041_156# _425_/a_1000_472#
+ _425_/a_1308_423# _425_/a_1456_156# _425_/a_1288_156# _425_/a_2248_156# _425_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 vdd vss _210_/a_255_603# _210_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss vdd vss FILLER_0_20_169/a_36_472# FILLER_0_20_169/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] vdd vss _408_/a_244_524# _408_/a_2215_68#
+ _408_/a_56_524# _408_/a_718_524# _408_/a_728_93# _408_/a_1936_472# _408_/a_1336_472#
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd vdd vss _339_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss vdd vss FILLER_0_21_286/a_36_472# FILLER_0_21_286/a_572_375#
+ FILLER_0_21_286/a_124_375# FILLER_0_21_286/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss vdd vss FILLER_0_12_220/a_1380_472# FILLER_0_12_220/a_36_472#
+ FILLER_0_12_220/a_932_472# FILLER_0_12_220/a_572_375# FILLER_0_12_220/a_124_375#
+ FILLER_0_12_220/a_1468_375# FILLER_0_12_220/a_1020_375# FILLER_0_12_220/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss vdd vss FILLER_0_8_247/a_1380_472# FILLER_0_8_247/a_36_472#
+ FILLER_0_8_247/a_932_472# FILLER_0_8_247/a_572_375# FILLER_0_8_247/a_124_375# FILLER_0_8_247/a_1468_375#
+ FILLER_0_8_247/a_1020_375# FILLER_0_8_247/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 net49 vss vdd net50 vdd vss fanout49/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_206 vdd vss vdd vss FILLER_0_5_206/a_36_472# FILLER_0_5_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd vdd vss _441_/a_2665_112# _441_/a_448_472#
+ _441_/a_796_472# _441_/a_36_151# _441_/a_1204_472# _441_/a_3041_156# _441_/a_1000_472#
+ _441_/a_1308_423# _441_/a_1456_156# _441_/a_1288_156# _441_/a_2248_156# _441_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ vdd vss _372_/a_2590_472# _372_/a_170_472#
+ _372_/a_1602_69# _372_/a_786_69# _372_/a_3126_472# _372_/a_1194_69# _372_/a_3662_472#
+ _372_/a_2034_472# _372_/a_358_69# gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__303__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vss vdd vss FILLER_0_17_142/a_36_472# FILLER_0_17_142/a_572_375#
+ FILLER_0_17_142/a_124_375# FILLER_0_17_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_54 vdd vss vdd vss FILLER_0_5_54/a_1380_472# FILLER_0_5_54/a_36_472# FILLER_0_5_54/a_932_472#
+ FILLER_0_5_54/a_572_375# FILLER_0_5_54/a_124_375# FILLER_0_5_54/a_1468_375# FILLER_0_5_54/a_1020_375#
+ FILLER_0_5_54/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_355_ vdd vss _149_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd vdd vss _424_/a_2665_112# _424_/a_448_472#
+ _424_/a_796_472# _424_/a_36_151# _424_/a_1204_472# _424_/a_3041_156# _424_/a_1000_472#
+ _424_/a_1308_423# _424_/a_1456_156# _424_/a_1288_156# _424_/a_2248_156# _424_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ vdd vss _005_ _094_ _101_ vdd vss _286_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_123 vdd vss vdd vss FILLER_0_14_123/a_36_472# FILLER_0_14_123/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ vdd vss _407_/a_36_472# _407_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ vdd vss _269_/a_36_472# _269_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss vdd vss FILLER_0_17_56/a_36_472# FILLER_0_17_56/a_572_375#
+ FILLER_0_17_56/a_124_375# FILLER_0_17_56/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vss _032_ _159_ vdd vdd vss _371_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd vdd vss _440_/a_2665_112# _440_/a_448_472#
+ _440_/a_796_472# _440_/a_36_151# _440_/a_1204_472# _440_/a_3041_156# _440_/a_1000_472#
+ _440_/a_1308_423# _440_/a_1456_156# _440_/a_1288_156# _440_/a_2248_156# _440_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd vss vdd vss FILLER_0_5_88/a_36_472# FILLER_0_5_88/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ _012_ net35 net55 vss net72 vdd vdd vss _423_/a_2665_112# _423_/a_448_472#
+ _423_/a_796_472# _423_/a_36_151# _423_/a_1204_472# _423_/a_3041_156# _423_/a_1000_472#
+ _423_/a_1308_423# _423_/a_1456_156# _423_/a_1288_156# _423_/a_2248_156# _423_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ vdd vss _354_/a_49_472# _354_/a_665_69#
+ _354_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_285_ net28 vdd vss _101_ mask\[1\] _099_ vdd vss _285_/a_36_472# _285_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_199_ net20 vss vdd _046_ vdd vss _199_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ vdd vss _337_/a_49_472# _337_/a_665_69#
+ _337_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] vdd vss _406_/a_36_159# gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ vdd vss _268_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss vdd vss FILLER_0_24_274/a_1380_472# FILLER_0_24_274/a_36_472#
+ FILLER_0_24_274/a_932_472# FILLER_0_24_274/a_572_375# FILLER_0_24_274/a_124_375#
+ FILLER_0_24_274/a_1468_375# FILLER_0_24_274/a_1020_375# FILLER_0_24_274/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ vdd vss _370_/a_848_380# _370_/a_1084_68#
+ _370_/a_124_24# _370_/a_1152_472# _370_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss vdd vss FILLER_0_1_266/a_36_472# FILLER_0_1_266/a_572_375#
+ FILLER_0_1_266/a_124_375# FILLER_0_1_266/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_422_ _011_ net34 net61 vss net78 vdd vdd vss _422_/a_2665_112# _422_/a_448_472#
+ _422_/a_796_472# _422_/a_36_151# _422_/a_1204_472# _422_/a_3041_156# _422_/a_1000_472#
+ _422_/a_1308_423# _422_/a_1456_156# _422_/a_1288_156# _422_/a_2248_156# _422_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_353_ vdd vss _148_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss vdd vss FILLER_0_17_133/a_36_472# FILLER_0_17_133/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output36_I vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_284_ vdd vss _004_ _094_ _100_ vdd vss _284_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_198_ vdd vss _046_ mask\[3\] net30 vdd vss _198_/a_255_603# _198_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_336_ vdd vss _138_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] vdd vss _405_/a_255_603# _405_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] vdd vss _267_/a_1792_472# _267_/a_224_472#
+ _267_/a_1568_472# _267_/a_36_472# _267_/a_1120_472# _267_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss vdd vss FILLER_0_6_177/a_36_472# FILLER_0_6_177/a_572_375#
+ FILLER_0_6_177/a_124_375# FILLER_0_6_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ vdd vss _319_/a_234_472# _319_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss vdd vss FILLER_0_8_239/a_36_472# FILLER_0_8_239/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss vdd vss FILLER_0_1_212/a_36_472# FILLER_0_1_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd vdd vss _421_/a_2665_112# _421_/a_448_472#
+ _421_/a_796_472# _421_/a_36_151# _421_/a_1204_472# _421_/a_3041_156# _421_/a_1000_472#
+ _421_/a_1308_423# _421_/a_1456_156# _421_/a_1288_156# _421_/a_2248_156# _421_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ vdd vss _352_/a_49_472# _352_/a_665_69#
+ _352_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ vdd vss _283_/a_36_472# _283_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vdd vss vdd vss FILLER_0_9_142/a_36_472# FILLER_0_9_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vss vdd vss FILLER_0_20_107/a_36_472# FILLER_0_20_107/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ vdd vss _404_/a_36_472# _404_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ vdd vss _335_/a_49_472# _335_/a_665_69#
+ _335_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_266_ vdd vss _055_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_197_ vdd vss net19 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd vss _124_ _115_ _118_ vdd vss _318_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd vss vdd vss FILLER_0_8_24/a_36_472# FILLER_0_8_24/a_572_375# FILLER_0_8_24/a_124_375#
+ FILLER_0_8_24/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss vdd vss FILLER_0_8_2/a_36_472# FILLER_0_8_2/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd vdd vss _420_/a_2665_112# _420_/a_448_472#
+ _420_/a_796_472# _420_/a_36_151# _420_/a_1204_472# _420_/a_3041_156# _420_/a_1000_472#
+ _420_/a_1308_423# _420_/a_1456_156# _420_/a_1288_156# _420_/a_2248_156# _420_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd vdd vss _282_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_334_ vss _137_ _132_ vdd vdd vss _334_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_403_ vdd vss _183_ cal_count\[2\] _176_ vdd vss _403_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vss vdd vss FILLER_0_6_90/a_36_472# FILLER_0_6_90/a_572_375# FILLER_0_6_90/a_124_375#
+ FILLER_0_6_90/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net19 vss vdd _045_ vdd vss _196_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ vdd vss _265_/a_468_472# _265_/a_224_472#
+ _265_/a_244_68# _265_/a_916_472# gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd vss vdd vss FILLER_0_17_38/a_36_472# FILLER_0_17_38/a_572_375#
+ FILLER_0_17_38/a_124_375# FILLER_0_17_38/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_248_ vss _070_ _069_ vdd vdd vss _248_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__409__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd vdd vss _317_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss vdd vss FILLER_0_2_171/a_36_472# FILLER_0_2_171/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss vdd vss FILLER_0_12_236/a_36_472# FILLER_0_12_236/a_572_375#
+ FILLER_0_12_236/a_124_375# FILLER_0_12_236/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ vdd vss _350_/a_49_472# _350_/a_665_69#
+ _350_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ vdd vss _281_/a_234_472# _281_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd vdd vss _333_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 vdd vss _195_/a_255_603# _195_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] vdd vss _402_/a_244_567# _402_/a_718_527#
+ _402_/a_2172_497# _402_/a_56_567# _402_/a_1948_68# _402_/a_728_93# _402_/a_1296_93#
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss vdd vss FILLER_0_11_109/a_36_472# FILLER_0_11_109/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] vdd vss _264_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss vdd vss FILLER_0_12_50/a_36_472# FILLER_0_12_50/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ vdd vss _247_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate vdd vss _316_/a_848_380# _316_/a_1084_68#
+ _316_/a_124_24# _316_/a_1152_472# _316_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_60 vdd vss vdd vss FILLER_0_23_60/a_36_472# FILLER_0_23_60/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vss vdd vss FILLER_0_15_212/a_1380_472# FILLER_0_15_212/a_36_472#
+ FILLER_0_15_212/a_932_472# FILLER_0_15_212/a_572_375# FILLER_0_15_212/a_124_375#
+ FILLER_0_15_212/a_1468_375# FILLER_0_15_212/a_1020_375# FILLER_0_15_212/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vss vdd vss FILLER_0_8_37/a_36_472# FILLER_0_8_37/a_572_375# FILLER_0_8_37/a_124_375#
+ FILLER_0_8_37/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss vdd vss FILLER_0_17_104/a_1380_472# FILLER_0_17_104/a_36_472#
+ FILLER_0_17_104/a_932_472# FILLER_0_17_104/a_572_375# FILLER_0_17_104/a_124_375#
+ FILLER_0_17_104/a_1468_375# FILLER_0_17_104/a_1020_375# FILLER_0_17_104/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_72 vdd vss vdd vss FILLER_0_15_72/a_36_472# FILLER_0_15_72/a_572_375#
+ FILLER_0_15_72/a_124_375# FILLER_0_15_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd vss vdd vss FILLER_0_1_204/a_36_472# FILLER_0_1_204/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ vdd vss _280_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss vdd vss FILLER_0_14_107/a_1380_472# FILLER_0_14_107/a_36_472#
+ FILLER_0_14_107/a_932_472# FILLER_0_14_107/a_572_375# FILLER_0_14_107/a_124_375#
+ FILLER_0_14_107/a_1468_375# FILLER_0_14_107/a_1020_375# FILLER_0_14_107/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ vdd _180_ _179_ _181_ _174_ vss vdd vss _401_/a_36_68# _401_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_332_ _126_ vdd vss _017_ _127_ _135_ vdd vss _332_/a_36_472# _332_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_194_ vss net8 net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ vdd vss _263_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss vdd vss FILLER_0_5_181/a_36_472# FILLER_0_5_181/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_246_ vss _068_ _055_ vdd vdd vss _246_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss vdd vss _315_/a_36_68# _315_/a_244_497#
+ _315_/a_1657_68# _315_/a_1229_68# _315_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_290 vdd vss vdd vss FILLER_0_23_290/a_36_472# FILLER_0_23_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss vdd vss FILLER_0_15_235/a_36_472# FILLER_0_15_235/a_572_375#
+ FILLER_0_15_235/a_124_375# FILLER_0_15_235/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ vdd vss _229_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss vdd vss FILLER_0_18_61/a_36_472# FILLER_0_18_61/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss vdd vss FILLER_0_11_282/a_36_472# FILLER_0_11_282/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss vdd vss FILLER_0_4_213/a_36_472# FILLER_0_4_213/a_572_375#
+ FILLER_0_4_213/a_124_375# FILLER_0_4_213/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ vdd vss _180_ cal_count\[1\] _178_ vdd vss _400_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_193_ net18 vss vdd _044_ vdd vss _193_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_331_ _134_ vdd vss _135_ _086_ _132_ vdd vss _331_/a_448_472# _331_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ vdd vss _121_ _085_ _069_ vdd vss _314_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_245_ vdd vss net6 _067_ net67 vdd vss _245_/a_234_472# _245_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_206 vdd vss vdd vss FILLER_0_21_206/a_36_472# FILLER_0_21_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd vdd vss _228_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss vdd vss FILLER_0_7_233/a_36_472# FILLER_0_7_233/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss vdd vss FILLER_0_9_60/a_36_472# FILLER_0_9_60/a_572_375# FILLER_0_9_60/a_124_375#
+ FILLER_0_9_60/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vss vdd vss FILLER_0_13_142/a_1380_472# FILLER_0_13_142/a_36_472#
+ FILLER_0_13_142/a_932_472# FILLER_0_13_142/a_572_375# FILLER_0_13_142/a_124_375#
+ FILLER_0_13_142/a_1468_375# FILLER_0_13_142/a_1020_375# FILLER_0_13_142/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ vdd vss _044_ mask\[1\] net28 vdd vss _192_/a_255_603# _192_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_261_ vss _081_ _059_ vdd vdd vss _261_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_330_ vdd vss _134_ _133_ _062_ vdd vss _330_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss vdd vss FILLER_0_12_20/a_36_472# FILLER_0_12_20/a_572_375#
+ FILLER_0_12_20/a_124_375# FILLER_0_12_20/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss vdd vss FILLER_0_5_172/a_36_472# FILLER_0_5_172/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ vdd vss en_co_clk _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__190__I vss _043_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_313_ vdd vss _120_ _059_ _119_ vdd vss _313_/a_255_603# _313_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__257__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd vdd vss _227_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss vdd vss FILLER_0_20_31/a_36_472# FILLER_0_20_31/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss vdd vss FILLER_0_9_72/a_1380_472# FILLER_0_9_72/a_36_472# FILLER_0_9_72/a_932_472#
+ FILLER_0_9_72/a_572_375# FILLER_0_9_72/a_124_375# FILLER_0_9_72/a_1468_375# FILLER_0_9_72/a_1020_375#
+ FILLER_0_9_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss vdd vss FILLER_0_0_96/a_36_472# FILLER_0_0_96/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss vdd vss _260_/a_36_68# _260_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ vdd vss _389_/a_428_148# _389_/a_36_148# gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ vdd vss _312_/a_234_472# _312_/a_672_472#
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd vss net47 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd vss vdd vss FILLER_0_23_282/a_36_472# FILLER_0_23_282/a_572_375#
+ FILLER_0_23_282/a_124_375# FILLER_0_23_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss vdd vss FILLER_0_15_205/a_36_472# FILLER_0_15_205/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss vdd vss FILLER_0_2_165/a_36_472# FILLER_0_2_165/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss vdd vss FILLER_0_18_53/a_36_472# FILLER_0_18_53/a_572_375#
+ FILLER_0_18_53/a_124_375# FILLER_0_18_53/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ vdd vss _226_/a_1044_68# _226_/a_452_68# _226_/a_276_68#
+ _226_/a_860_68# gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_98 vdd vss vdd vss FILLER_0_20_98/a_36_472# FILLER_0_20_98/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_87 vdd vss vdd vss FILLER_0_20_87/a_36_472# FILLER_0_20_87/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss vdd vss FILLER_0_19_171/a_1380_472# FILLER_0_19_171/a_36_472#
+ FILLER_0_19_171/a_932_472# FILLER_0_19_171/a_572_375# FILLER_0_19_171/a_124_375#
+ FILLER_0_19_171/a_1468_375# FILLER_0_19_171/a_1020_375# FILLER_0_19_171/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss vdd vss FILLER_0_15_10/a_36_472# FILLER_0_15_10/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss vdd vss FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_572_375# FILLER_0_15_2/a_124_375#
+ FILLER_0_15_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss vdd vss FILLER_0_22_177/a_1380_472# FILLER_0_22_177/a_36_472#
+ FILLER_0_22_177/a_932_472# FILLER_0_22_177/a_572_375# FILLER_0_22_177/a_124_375#
+ FILLER_0_22_177/a_1468_375# FILLER_0_22_177/a_1020_375# FILLER_0_22_177/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss vdd vss FILLER_0_13_100/a_36_472# FILLER_0_13_100/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss vdd vss FILLER_0_9_105/a_36_472# FILLER_0_9_105/a_572_375#
+ FILLER_0_9_105/a_124_375# FILLER_0_9_105/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ vdd vss _190_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ vdd vss _311_/a_692_473# _311_/a_254_473#
+ _311_/a_66_473# _311_/a_2700_473# _311_/a_1660_473# _311_/a_3220_473# _311_/a_1212_473#
+ _311_/a_2180_473# _311_/a_3740_473# _311_/a_1920_473# gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_242_ net47 vss vdd _066_ vdd vss _242_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_228 vdd vss vdd vss FILLER_0_15_228/a_36_472# FILLER_0_15_228/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss vdd vss FILLER_0_2_111/a_1380_472# FILLER_0_2_111/a_36_472#
+ FILLER_0_2_111/a_932_472# FILLER_0_2_111/a_572_375# FILLER_0_2_111/a_124_375# FILLER_0_2_111/a_1468_375#
+ FILLER_0_2_111/a_1020_375# FILLER_0_2_111/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss vdd vss FILLER_0_2_177/a_36_472# FILLER_0_2_177/a_572_375#
+ FILLER_0_2_177/a_124_375# FILLER_0_2_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd vdd vss _225_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss vdd vss FILLER_0_18_76/a_36_472# FILLER_0_18_76/a_572_375#
+ FILLER_0_18_76/a_124_375# FILLER_0_18_76/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ vdd vss _208_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd vdd vss _387_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_310_ _090_ vdd vss _117_ _060_ _113_ vdd vss _310_/a_49_472# _310_/a_1133_69# _310_/a_741_69#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_164 vdd vss vdd vss FILLER_0_5_164/a_36_472# FILLER_0_5_164/a_572_375#
+ FILLER_0_5_164/a_124_375# FILLER_0_5_164/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd vss vdd vss FILLER_0_23_88/a_36_472# FILLER_0_23_88/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss vdd vss FILLER_0_23_44/a_1380_472# FILLER_0_23_44/a_36_472#
+ FILLER_0_23_44/a_932_472# FILLER_0_23_44/a_572_375# FILLER_0_23_44/a_124_375# FILLER_0_23_44/a_1468_375#
+ FILLER_0_23_44/a_1020_375# FILLER_0_23_44/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] vdd vss _241_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd vdd vss _439_/a_2665_112# _439_/a_448_472#
+ _439_/a_796_472# _439_/a_36_151# _439_/a_1204_472# _439_/a_3041_156# _439_/a_1000_472#
+ _439_/a_1308_423# _439_/a_1456_156# _439_/a_1288_156# _439_/a_2248_156# _439_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd vss vdd vss FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss vdd vss FILLER_0_3_54/a_36_472# FILLER_0_3_54/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd vss _049_ mask\[6\] net33 vdd vss _207_/a_255_603# _207_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss vdd vss FILLER_0_19_195/a_36_472# FILLER_0_19_195/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss vdd vss FILLER_0_0_232/a_36_472# FILLER_0_0_232/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss vdd vss FILLER_0_16_154/a_1380_472# FILLER_0_16_154/a_36_472#
+ FILLER_0_16_154/a_932_472# FILLER_0_16_154/a_572_375# FILLER_0_16_154/a_124_375#
+ FILLER_0_16_154/a_1468_375# FILLER_0_16_154/a_1020_375# FILLER_0_16_154/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss vdd vss FILLER_0_20_2/a_36_472# FILLER_0_20_2/a_572_375# FILLER_0_20_2/a_124_375#
+ FILLER_0_20_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ vdd vss _386_/a_848_380# _386_/a_1084_68#
+ _386_/a_124_24# _386_/a_1152_472# _386_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss vdd vss FILLER_0_5_198/a_36_472# FILLER_0_5_198/a_572_375#
+ FILLER_0_5_198/a_124_375# FILLER_0_5_198/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_240_ vdd vss net41 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_282 vdd vss vdd vss FILLER_0_17_282/a_36_472# FILLER_0_17_282/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_274 vdd vss vdd vss FILLER_0_23_274/a_36_472# FILLER_0_23_274/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd vdd vss _438_/a_2665_112# _438_/a_448_472#
+ _438_/a_796_472# _438_/a_36_151# _438_/a_1204_472# _438_/a_3041_156# _438_/a_1000_472#
+ _438_/a_1308_423# _438_/a_1456_156# _438_/a_1288_156# _438_/a_2248_156# _438_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ vdd vss _369_/a_36_68# _369_/a_244_472#
+ _369_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss vdd vss FILLER_0_14_263/a_36_472# FILLER_0_14_263/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] vdd vss _223_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss vdd vss FILLER_0_9_290/a_36_472# FILLER_0_9_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss vdd vss FILLER_0_0_266/a_36_472# FILLER_0_0_266/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss vdd vss _385_/a_36_68# _385_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ vdd vss _299_/a_36_472# _299_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd vdd vss _437_/a_2665_112# _437_/a_448_472#
+ _437_/a_796_472# _437_/a_36_151# _437_/a_1204_472# _437_/a_3041_156# _437_/a_1000_472#
+ _437_/a_1308_423# _437_/a_1456_156# _437_/a_1288_156# _437_/a_2248_156# _437_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_78 vdd vss vdd vss FILLER_0_3_78/a_36_472# FILLER_0_3_78/a_572_375# FILLER_0_3_78/a_124_375#
+ FILLER_0_3_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_368_ vdd vss trim_mask\[4\] _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_222_ vdd vss net38 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ vdd vss _205_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss vdd vss FILLER_0_19_142/a_36_472# FILLER_0_19_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd vdd vss _453_/a_2665_112# _453_/a_448_472#
+ _453_/a_796_472# _453_/a_36_151# _453_/a_1204_472# _453_/a_3041_156# _453_/a_1000_472#
+ _453_/a_1308_423# _453_/a_1456_156# _453_/a_1288_156# _453_/a_2248_156# _453_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ vdd vss _384_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss vdd vss FILLER_0_10_107/a_36_472# FILLER_0_10_107/a_572_375#
+ FILLER_0_10_107/a_124_375# FILLER_0_10_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ vdd vss _298_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd vdd vss _436_/a_2665_112# _436_/a_448_472#
+ _436_/a_796_472# _436_/a_36_151# _436_/a_1204_472# _436_/a_3041_156# _436_/a_1000_472#
+ _436_/a_1308_423# _436_/a_1456_156# _436_/a_1288_156# _436_/a_2248_156# _436_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ vdd vss _367_/a_36_68# _367_/a_244_472#
+ _367_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss vdd vss FILLER_0_13_80/a_36_472# FILLER_0_13_80/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss vdd vss FILLER_0_1_192/a_36_472# FILLER_0_1_192/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd vss vdd vss FILLER_0_9_270/a_36_472# FILLER_0_9_270/a_572_375#
+ FILLER_0_9_270/a_124_375# FILLER_0_9_270/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vss net38 _054_ vdd vdd vss _221_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ _008_ net31 net60 vss net77 vdd vdd vss _419_/a_2665_112# _419_/a_448_472#
+ _419_/a_796_472# _419_/a_36_151# _419_/a_1204_472# _419_/a_3041_156# _419_/a_1000_472#
+ _419_/a_1308_423# _419_/a_1456_156# _419_/a_1288_156# _419_/a_2248_156# _419_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 vdd vss _204_/a_255_603# _204_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss vdd vss FILLER_0_20_15/a_1380_472# FILLER_0_20_15/a_36_472#
+ FILLER_0_20_15/a_932_472# FILLER_0_20_15/a_572_375# FILLER_0_20_15/a_124_375# FILLER_0_20_15/a_1468_375#
+ FILLER_0_20_15/a_1020_375# FILLER_0_20_15/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss vdd vss FILLER_0_19_187/a_36_472# FILLER_0_19_187/a_572_375#
+ FILLER_0_19_187/a_124_375# FILLER_0_19_187/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss vdd vss FILLER_0_3_221/a_1380_472# FILLER_0_3_221/a_36_472#
+ FILLER_0_3_221/a_932_472# FILLER_0_3_221/a_572_375# FILLER_0_3_221/a_124_375# FILLER_0_3_221/a_1468_375#
+ FILLER_0_3_221/a_1020_375# FILLER_0_3_221/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss vdd vss FILLER_0_15_59/a_36_472# FILLER_0_15_59/a_572_375#
+ FILLER_0_15_59/a_124_375# FILLER_0_15_59/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd vss vdd vss FILLER_0_6_79/a_36_472# FILLER_0_6_79/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 vdd vss _452_/a_448_472# _452_/a_36_151#
+ _452_/a_1293_527# _452_/a_3081_151# _452_/a_1284_156# _452_/a_1040_527# _452_/a_1353_112#
+ _452_/a_836_156# _452_/a_1697_156# _452_/a_2449_156# _452_/a_3129_107# _452_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ vdd vss _383_/a_36_472# _383_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ vdd vss _297_/a_36_472# _297_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd vdd vss _435_/a_2665_112# _435_/a_448_472#
+ _435_/a_796_472# _435_/a_36_151# _435_/a_1204_472# _435_/a_3041_156# _435_/a_1000_472#
+ _435_/a_1308_423# _435_/a_1456_156# _435_/a_1288_156# _435_/a_2248_156# _435_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A2 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ vdd vss trim_mask\[3\] _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_127 vdd vss vdd vss FILLER_0_2_127/a_36_472# FILLER_0_2_127/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vss vdd vss FILLER_0_18_37/a_1380_472# FILLER_0_18_37/a_36_472#
+ FILLER_0_18_37/a_932_472# FILLER_0_18_37/a_572_375# FILLER_0_18_37/a_124_375# FILLER_0_18_37/a_1468_375#
+ FILLER_0_18_37/a_1020_375# FILLER_0_18_37/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vss vdd vss FILLER_0_9_282/a_36_472# FILLER_0_9_282/a_572_375#
+ FILLER_0_9_282/a_124_375# FILLER_0_9_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd vss _054_ trim_val\[0\] _053_ vdd vss _220_/a_255_603# _220_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_349_ vdd vss _146_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _007_ net30 net60 vss net77 vdd vdd vss _418_/a_2665_112# _418_/a_448_472#
+ _418_/a_796_472# _418_/a_36_151# _418_/a_1204_472# _418_/a_3041_156# _418_/a_1000_472#
+ _418_/a_1308_423# _418_/a_1456_156# _418_/a_1288_156# _418_/a_2248_156# _418_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output21_I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss vdd vss FILLER_0_19_155/a_36_472# FILLER_0_19_155/a_572_375#
+ FILLER_0_19_155/a_124_375# FILLER_0_19_155/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss vdd vss FILLER_0_19_111/a_36_472# FILLER_0_19_111/a_572_375#
+ FILLER_0_19_111/a_124_375# FILLER_0_19_111/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss vdd vss FILLER_0_22_128/a_1916_375# FILLER_0_22_128/a_1380_472#
+ FILLER_0_22_128/a_3260_375# FILLER_0_22_128/a_36_472# FILLER_0_22_128/a_932_472#
+ FILLER_0_22_128/a_2812_375# FILLER_0_22_128/a_2276_472# FILLER_0_22_128/a_1828_472#
+ FILLER_0_22_128/a_3172_472# FILLER_0_22_128/a_572_375# FILLER_0_22_128/a_2724_472#
+ FILLER_0_22_128/a_124_375# FILLER_0_22_128/a_1468_375# FILLER_0_22_128/a_1020_375#
+ FILLER_0_22_128/a_484_472# FILLER_0_22_128/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss vdd vss FILLER_0_15_180/a_36_472# FILLER_0_15_180/a_572_375#
+ FILLER_0_15_180/a_124_375# FILLER_0_15_180/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss vdd vss FILLER_0_21_150/a_36_472# FILLER_0_21_150/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss vdd vss FILLER_0_6_47/a_1916_375# FILLER_0_6_47/a_1380_472#
+ FILLER_0_6_47/a_3260_375# FILLER_0_6_47/a_36_472# FILLER_0_6_47/a_932_472# FILLER_0_6_47/a_2812_375#
+ FILLER_0_6_47/a_2276_472# FILLER_0_6_47/a_1828_472# FILLER_0_6_47/a_3172_472# FILLER_0_6_47/a_572_375#
+ FILLER_0_6_47/a_2724_472# FILLER_0_6_47/a_124_375# FILLER_0_6_47/a_1468_375# FILLER_0_6_47/a_1020_375#
+ FILLER_0_6_47/a_484_472# FILLER_0_6_47/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 vdd vss _451_/a_448_472# _451_/a_36_151#
+ _451_/a_1293_527# _451_/a_3081_151# _451_/a_1284_156# _451_/a_1040_527# _451_/a_1353_112#
+ _451_/a_836_156# _451_/a_1697_156# _451_/a_2449_156# _451_/a_3129_107# _451_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_28 vdd vss vdd vss FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd vss _035_ _160_ _167_ vdd vss _382_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss vdd vss FILLER_0_18_209/a_36_472# FILLER_0_18_209/a_572_375#
+ FILLER_0_18_209/a_124_375# FILLER_0_18_209/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss vdd vss FILLER_0_5_136/a_36_472# FILLER_0_5_136/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ vdd vss _296_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd vdd vss _434_/a_2665_112# _434_/a_448_472#
+ _434_/a_796_472# _434_/a_36_151# _434_/a_1204_472# _434_/a_3041_156# _434_/a_1000_472#
+ _434_/a_1308_423# _434_/a_1456_156# _434_/a_1288_156# _434_/a_2248_156# _434_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ vdd vss _365_/a_36_68# _365_/a_244_472#
+ _365_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ vdd vss _348_/a_49_472# _348_/a_665_69#
+ _348_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd vdd vss _417_/a_2665_112# _417_/a_448_472#
+ _417_/a_796_472# _417_/a_36_151# _417_/a_1204_472# _417_/a_3041_156# _417_/a_1000_472#
+ _417_/a_1308_423# _417_/a_1456_156# _417_/a_1288_156# _417_/a_2248_156# _417_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_279_ vdd vss _096_ _090_ state\[1\] vdd vss _279_/a_652_68# _279_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_231 vdd vss vdd vss FILLER_0_6_231/a_36_472# FILLER_0_6_231/a_572_375#
+ FILLER_0_6_231/a_124_375# FILLER_0_6_231/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ vdd vss _202_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output14_I vss net14 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd vss vdd vss FILLER_0_4_91/a_36_472# FILLER_0_4_91/a_572_375# FILLER_0_4_91/a_124_375#
+ FILLER_0_4_91/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_94 vdd vss vdd vss FILLER_0_10_94/a_36_472# FILLER_0_10_94/a_572_375#
+ FILLER_0_10_94/a_124_375# FILLER_0_10_94/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss vdd vss FILLER_0_3_212/a_36_472# FILLER_0_3_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss vdd vss FILLER_0_19_134/a_36_472# FILLER_0_19_134/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss vdd vss FILLER_0_16_115/a_36_472# FILLER_0_16_115/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss vdd vss FILLER_0_22_107/a_36_472# FILLER_0_22_107/a_572_375#
+ FILLER_0_22_107/a_124_375# FILLER_0_22_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss vdd vss FILLER_0_21_60/a_36_472# FILLER_0_21_60/a_572_375#
+ FILLER_0_21_60/a_124_375# FILLER_0_21_60/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss vdd vss FILLER_0_6_37/a_36_472# FILLER_0_6_37/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd vss vdd vss FILLER_0_8_156/a_36_472# FILLER_0_8_156/a_572_375#
+ FILLER_0_8_156/a_124_375# FILLER_0_8_156/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I vss rstn vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__243__I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 vdd vss _450_/a_448_472# _450_/a_36_151#
+ _450_/a_1293_527# _450_/a_3081_151# _450_/a_1284_156# _450_/a_1040_527# _450_/a_1353_112#
+ _450_/a_836_156# _450_/a_1697_156# _450_/a_2449_156# _450_/a_3129_107# _450_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xoutput40 trim[2] net40 vdd vss vdd vss output40/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ vdd vss _381_/a_36_472# _381_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_148 vdd vss vdd vss FILLER_0_5_148/a_36_472# FILLER_0_5_148/a_572_375#
+ FILLER_0_5_148/a_124_375# FILLER_0_5_148/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd vdd vss _433_/a_2665_112# _433_/a_448_472#
+ _433_/a_796_472# _433_/a_36_151# _433_/a_1204_472# _433_/a_3041_156# _433_/a_1000_472#
+ _433_/a_1308_423# _433_/a_1456_156# _433_/a_1288_156# _433_/a_2248_156# _433_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ vdd vss _295_/a_36_472# _295_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss vdd vss FILLER_0_14_235/a_36_472# FILLER_0_14_235/a_572_375#
+ FILLER_0_14_235/a_124_375# FILLER_0_14_235/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss vdd vss FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_572_375#
+ FILLER_0_13_72/a_124_375# FILLER_0_13_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_347_ vdd vss _145_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 vdd vss _278_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_290 vdd vss vdd vss FILLER_0_13_290/a_36_472# FILLER_0_13_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ _005_ net28 net62 vss net79 vdd vdd vss _416_/a_2665_112# _416_/a_448_472#
+ _416_/a_796_472# _416_/a_36_151# _416_/a_1204_472# _416_/a_3041_156# _416_/a_1000_472#
+ _416_/a_1308_423# _416_/a_1456_156# _416_/a_1288_156# _416_/a_2248_156# _416_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_201_ vdd vss _047_ mask\[4\] net31 vdd vss _201_/a_255_603# _201_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 result[3] net30 vdd vss vdd vss output30/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_196 vdd vss vdd vss FILLER_0_12_196/a_36_472# FILLER_0_12_196/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 clkc net6 vdd vss vdd vss output6/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss vdd vss output41/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ vdd vss _380_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
C0 FILLER_0_3_172/a_36_472# FILLER_0_5_172/a_124_375# 0.0027f
C1 net52 trim_val\[3\] 0.082691f
C2 net82 FILLER_0_4_213/a_124_375# 0.00123f
C3 _056_ _070_ 0.045548f
C4 FILLER_0_17_72/a_3172_472# vss 0.001338f
C5 FILLER_0_11_124/a_36_472# _120_ 0.014712f
C6 _443_/a_36_151# net69 0.069715f
C7 FILLER_0_9_142/a_124_375# calibrate 0.001505f
C8 net61 _009_ 0.042703f
C9 fanout61/a_36_113# net79 0.001865f
C10 output35/a_224_472# FILLER_0_22_177/a_1380_472# 0.002486f
C11 fanout80/a_36_113# _136_ 0.006151f
C12 net50 trim_mask\[0\] 0.002835f
C13 _126_ _085_ 0.02154f
C14 _144_ _346_/a_49_472# 0.036821f
C15 _323_/a_36_113# net64 0.06154f
C16 net38 _039_ 0.059899f
C17 net16 net40 0.039189f
C18 vss output6/a_224_472# 0.004205f
C19 net52 FILLER_0_0_130/a_124_375# 0.004055f
C20 _105_ net78 0.004705f
C21 _105_ net60 0.042726f
C22 net16 trim_mask\[2\] 0.002527f
C23 _126_ _018_ 0.001243f
C24 net79 net22 0.042486f
C25 _141_ net56 0.012364f
C26 net16 _447_/a_1308_423# 0.001178f
C27 ctln[9] _447_/a_36_151# 0.010503f
C28 net57 FILLER_0_13_100/a_124_375# 0.012636f
C29 net61 fanout78/a_36_113# 0.056484f
C30 fanout60/a_36_160# net61 0.001167f
C31 FILLER_0_4_197/a_572_375# vdd 0.002455f
C32 net17 net51 0.026974f
C33 _015_ FILLER_0_8_247/a_932_472# 0.005458f
C34 net81 net79 0.178225f
C35 en net64 0.01789f
C36 _048_ _047_ 0.007849f
C37 _343_/a_257_69# mask\[4\] 0.001786f
C38 FILLER_0_16_107/a_36_472# net14 0.004691f
C39 net18 net30 0.09055f
C40 net58 net18 0.091503f
C41 _024_ vdd 0.091532f
C42 _424_/a_36_151# vdd 0.125156f
C43 net60 _010_ 0.108311f
C44 _098_ _434_/a_2665_112# 0.013854f
C45 _441_/a_796_472# vss 0.001231f
C46 _066_ _386_/a_848_380# 0.00416f
C47 _079_ _080_ 0.022852f
C48 output20/a_224_472# mask\[7\] 0.024731f
C49 _133_ _058_ 0.092697f
C50 state\[2\] _427_/a_2665_112# 0.007007f
C51 _425_/a_2665_112# net18 0.003301f
C52 FILLER_0_23_290/a_124_375# FILLER_0_23_282/a_572_375# 0.012001f
C53 net55 _452_/a_36_151# 0.042427f
C54 net57 net70 0.012088f
C55 _015_ _426_/a_796_472# 0.007696f
C56 FILLER_0_13_206/a_36_472# vdd 0.011681f
C57 _009_ _108_ 1.645945f
C58 FILLER_0_13_206/a_124_375# vss 0.051723f
C59 _193_/a_36_160# FILLER_0_13_290/a_124_375# 0.005732f
C60 _447_/a_448_472# vdd 0.014537f
C61 _447_/a_36_151# vss 0.001541f
C62 FILLER_0_18_2/a_2812_375# vdd 0.021655f
C63 _068_ _315_/a_244_497# 0.004768f
C64 _115_ FILLER_0_9_105/a_36_472# 0.004013f
C65 net57 net47 0.279638f
C66 _440_/a_2665_112# vss 0.008703f
C67 result[2] output30/a_224_472# 0.045862f
C68 _439_/a_1308_423# vss 0.009355f
C69 net80 _434_/a_1204_472# 0.003997f
C70 mask\[5\] net21 0.212814f
C71 _091_ FILLER_0_13_212/a_484_472# 0.04953f
C72 _412_/a_1308_423# net58 0.037719f
C73 fanout56/a_36_113# vss 0.03072f
C74 _411_/a_36_151# vdd 0.077963f
C75 FILLER_0_2_93/a_36_472# _441_/a_2665_112# 0.007491f
C76 FILLER_0_8_107/a_36_472# net14 0.001596f
C77 _098_ mask\[2\] 0.06158f
C78 _098_ _437_/a_796_472# 0.0049f
C79 net20 FILLER_0_3_221/a_1380_472# 0.008749f
C80 _053_ _152_ 0.032961f
C81 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_36_472# 0.003468f
C82 FILLER_0_7_72/a_36_472# _439_/a_36_151# 0.013806f
C83 FILLER_0_7_104/a_1468_375# _129_ 0.001165f
C84 FILLER_0_7_104/a_36_472# _131_ 0.002019f
C85 net36 _438_/a_1000_472# 0.072117f
C86 net27 FILLER_0_11_282/a_36_472# 0.001526f
C87 _386_/a_848_380# net37 0.006086f
C88 net56 _433_/a_2665_112# 0.003434f
C89 FILLER_0_15_180/a_124_375# vdd 0.016985f
C90 net63 _434_/a_2665_112# 0.120476f
C91 _021_ _091_ 0.016024f
C92 net15 _441_/a_448_472# 0.049213f
C93 trim[1] vss 0.085436f
C94 _155_ FILLER_0_7_104/a_124_375# 0.007925f
C95 net35 _207_/a_67_603# 0.005045f
C96 net67 _221_/a_36_160# 0.008581f
C97 mask\[5\] FILLER_0_20_177/a_484_472# 0.016114f
C98 mask\[9\] net14 0.090939f
C99 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_36_472# 0.002296f
C100 _126_ _320_/a_224_472# 0.003754f
C101 net17 _381_/a_36_472# 0.002796f
C102 _077_ _251_/a_906_472# 0.001076f
C103 _004_ fanout79/a_36_160# 0.048599f
C104 net35 _435_/a_36_151# 0.038368f
C105 en vss 0.466499f
C106 _259_/a_455_68# _076_ 0.002372f
C107 FILLER_0_16_73/a_484_472# _040_ 0.004877f
C108 _028_ FILLER_0_6_79/a_124_375# 0.015932f
C109 FILLER_0_14_99/a_36_472# _043_ 0.001242f
C110 net15 _440_/a_1204_472# 0.01349f
C111 net65 net75 0.135447f
C112 FILLER_0_21_142/a_36_472# FILLER_0_22_128/a_1468_375# 0.001543f
C113 _088_ _083_ 0.007169f
C114 net32 output33/a_224_472# 0.018183f
C115 net15 _439_/a_36_151# 0.068183f
C116 FILLER_0_3_78/a_36_472# _168_ 0.063262f
C117 _161_ _228_/a_36_68# 0.055774f
C118 _311_/a_254_473# vdd 0.001207f
C119 _292_/a_36_160# net22 0.001864f
C120 _452_/a_1353_112# net40 0.003745f
C121 _053_ trim_val\[0\] 0.446477f
C122 mask\[5\] FILLER_0_18_177/a_124_375# 0.002726f
C123 net34 net80 0.041846f
C124 net63 mask\[2\] 0.553545f
C125 _232_/a_67_603# net66 0.001758f
C126 FILLER_0_7_146/a_36_472# _076_ 0.001843f
C127 FILLER_0_7_146/a_124_375# _068_ 0.033245f
C128 FILLER_0_22_86/a_1380_472# net14 0.039176f
C129 result[4] _418_/a_36_151# 0.005556f
C130 output31/a_224_472# net19 0.072666f
C131 net36 FILLER_0_15_212/a_572_375# 0.004606f
C132 _435_/a_1308_423# vdd 0.012856f
C133 FILLER_0_19_111/a_36_472# net14 0.00143f
C134 _448_/a_2665_112# net59 0.005948f
C135 _176_ _267_/a_36_472# 0.001681f
C136 _085_ _267_/a_224_472# 0.002907f
C137 net31 _419_/a_2665_112# 0.004446f
C138 _176_ FILLER_0_15_59/a_572_375# 0.007169f
C139 _144_ _098_ 1.252524f
C140 _031_ _160_ 0.004547f
C141 _408_/a_1336_472# _184_ 0.003286f
C142 _427_/a_1000_472# vss 0.012657f
C143 _374_/a_36_68# vdd 0.075685f
C144 FILLER_0_21_133/a_36_472# net54 0.02286f
C145 FILLER_0_7_72/a_2276_472# vdd 0.004035f
C146 _392_/a_36_68# FILLER_0_12_50/a_36_472# 0.002811f
C147 FILLER_0_15_235/a_124_375# net62 0.001315f
C148 FILLER_0_15_282/a_124_375# net18 0.048284f
C149 ctln[3] net58 0.00479f
C150 FILLER_0_9_223/a_124_375# _128_ 0.004252f
C151 net65 fanout65/a_36_113# 0.019148f
C152 FILLER_0_9_28/a_2364_375# vdd 0.004562f
C153 FILLER_0_8_24/a_124_375# _054_ 0.008177f
C154 vss FILLER_0_21_60/a_572_375# 0.021222f
C155 vdd FILLER_0_21_60/a_36_472# 0.08419f
C156 _161_ calibrate 0.044443f
C157 FILLER_0_8_127/a_124_375# vss 0.019066f
C158 FILLER_0_8_127/a_36_472# vdd 0.069117f
C159 mask\[5\] FILLER_0_19_171/a_1380_472# 0.007596f
C160 _451_/a_448_472# _040_ 0.026819f
C161 _281_/a_672_472# vdd 0.001069f
C162 FILLER_0_7_162/a_124_375# vdd 0.011809f
C163 _427_/a_1000_472# net74 0.009646f
C164 FILLER_0_21_28/a_1380_472# net17 0.001709f
C165 _331_/a_448_472# vdd 0.001343f
C166 net27 FILLER_0_8_263/a_124_375# 0.016669f
C167 net44 _450_/a_836_156# 0.006278f
C168 net62 net30 0.339141f
C169 FILLER_0_13_290/a_36_472# _416_/a_36_151# 0.001723f
C170 FILLER_0_22_177/a_484_472# net33 0.013149f
C171 _398_/a_36_113# _043_ 0.005985f
C172 net68 _453_/a_448_472# 0.01245f
C173 FILLER_0_8_127/a_124_375# net74 0.026604f
C174 FILLER_0_13_212/a_572_375# vdd 0.001551f
C175 FILLER_0_13_212/a_124_375# vss 0.007116f
C176 _053_ _070_ 2.345795f
C177 FILLER_0_17_72/a_1020_375# _131_ 0.005847f
C178 _439_/a_36_151# net51 0.00711f
C179 vdd _145_ 0.082579f
C180 _016_ FILLER_0_12_136/a_1020_375# 0.001659f
C181 _127_ _395_/a_36_488# 0.00519f
C182 _140_ mask\[7\] 0.064343f
C183 _111_ _110_ 0.00195f
C184 FILLER_0_5_72/a_1468_375# net47 0.005049f
C185 output21/a_224_472# net22 0.022576f
C186 _140_ _148_ 0.011699f
C187 _162_ _061_ 0.001665f
C188 FILLER_0_2_177/a_36_472# net22 0.002517f
C189 output24/a_224_472# _025_ 0.010601f
C190 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_484_472# 0.026657f
C191 _337_/a_49_472# vdd 0.028131f
C192 _277_/a_36_160# _102_ 0.061995f
C193 _428_/a_36_151# _095_ 0.006658f
C194 FILLER_0_9_223/a_124_375# state\[0\] 0.002912f
C195 _401_/a_36_68# _179_ 0.007074f
C196 _360_/a_36_160# _152_ 0.040508f
C197 cal_itt\[3\] net22 0.134309f
C198 _407_/a_36_472# vdd 0.095308f
C199 trim[4] net47 0.009333f
C200 _274_/a_36_68# FILLER_0_12_220/a_932_472# 0.001237f
C201 net35 net14 0.040959f
C202 mask\[7\] FILLER_0_22_128/a_124_375# 0.01319f
C203 _057_ _311_/a_254_473# 0.002364f
C204 FILLER_0_20_193/a_36_472# net21 0.001099f
C205 _065_ ctln[8] 0.193903f
C206 _325_/a_224_472# _118_ 0.004845f
C207 ctln[1] net8 0.678616f
C208 output39/a_224_472# _444_/a_36_151# 0.062717f
C209 FILLER_0_7_59/a_484_472# vdd 0.00824f
C210 FILLER_0_7_59/a_36_472# vss 0.004006f
C211 FILLER_0_17_200/a_124_375# net21 0.048656f
C212 _132_ net53 0.035348f
C213 _412_/a_36_151# net81 0.014094f
C214 net80 FILLER_0_22_177/a_124_375# 0.013214f
C215 net35 FILLER_0_22_128/a_3260_375# 0.012732f
C216 FILLER_0_1_204/a_36_472# vss 0.002247f
C217 net36 _451_/a_36_151# 0.02414f
C218 _114_ FILLER_0_12_136/a_484_472# 0.003953f
C219 _144_ FILLER_0_22_128/a_3172_472# 0.001287f
C220 _395_/a_36_488# _071_ 0.00276f
C221 _437_/a_2665_112# FILLER_0_22_107/a_572_375# 0.001597f
C222 net68 FILLER_0_6_47/a_1020_375# 0.029857f
C223 FILLER_0_12_20/a_572_375# net17 0.041149f
C224 fanout72/a_36_113# _174_ 0.026207f
C225 _013_ _424_/a_1308_423# 0.007751f
C226 net58 _425_/a_2560_156# 0.004835f
C227 FILLER_0_9_72/a_1020_375# _439_/a_36_151# 0.059049f
C228 _255_/a_224_552# _056_ 0.033615f
C229 output19/a_224_472# _422_/a_2665_112# 0.024396f
C230 net20 _294_/a_224_472# 0.008053f
C231 input1/a_36_113# input2/a_36_113# 0.029417f
C232 trim_mask\[1\] FILLER_0_6_47/a_1916_375# 0.007169f
C233 _365_/a_36_68# net14 0.017522f
C234 FILLER_0_3_142/a_124_375# vdd 0.00167f
C235 _274_/a_36_68# _091_ 0.025773f
C236 net63 FILLER_0_22_177/a_1020_375# 0.003419f
C237 net38 clkc 0.088241f
C238 FILLER_0_0_96/a_124_375# net14 0.077876f
C239 _080_ vss 0.012982f
C240 trimb[1] cal_count\[2\] 0.003178f
C241 net57 state\[1\] 0.154183f
C242 FILLER_0_22_128/a_36_472# vss 0.001309f
C243 FILLER_0_22_128/a_484_472# vdd 0.002467f
C244 FILLER_0_16_89/a_124_375# _451_/a_448_472# 0.001597f
C245 net72 FILLER_0_17_64/a_36_472# 0.001145f
C246 _033_ _166_ 0.004448f
C247 FILLER_0_7_72/a_3260_375# net14 0.025344f
C248 _444_/a_1308_423# vdd 0.005677f
C249 FILLER_0_21_28/a_1916_375# _423_/a_36_151# 0.001597f
C250 net73 _334_/a_36_160# 0.003275f
C251 trim_val\[0\] _164_ 0.133785f
C252 _077_ FILLER_0_8_239/a_124_375# 0.001772f
C253 _127_ calibrate 0.004656f
C254 fanout49/a_36_160# FILLER_0_5_88/a_124_375# 0.001154f
C255 net52 _376_/a_36_160# 0.00267f
C256 net54 _438_/a_2248_156# 0.014423f
C257 fanout77/a_36_113# _419_/a_36_151# 0.002361f
C258 _075_ _081_ 0.001195f
C259 FILLER_0_15_282/a_124_375# net62 0.012711f
C260 FILLER_0_7_59/a_124_375# net15 0.004662f
C261 _128_ net4 0.039671f
C262 FILLER_0_7_146/a_124_375# vdd 0.034288f
C263 net41 _186_ 0.054661f
C264 net26 FILLER_0_23_44/a_124_375# 0.007775f
C265 _073_ FILLER_0_3_221/a_1380_472# 0.045839f
C266 net20 FILLER_0_15_228/a_124_375# 0.047331f
C267 net65 _413_/a_1000_472# 0.02866f
C268 en_co_clk fanout55/a_36_160# 0.041263f
C269 _052_ FILLER_0_19_28/a_484_472# 0.003325f
C270 net22 FILLER_0_18_209/a_124_375# 0.012909f
C271 fanout56/a_36_113# _097_ 0.062226f
C272 net27 FILLER_0_9_270/a_484_472# 0.023461f
C273 FILLER_0_10_78/a_1020_375# vss 0.002352f
C274 FILLER_0_10_78/a_1468_375# vdd 0.001778f
C275 _408_/a_718_524# _043_ 0.003719f
C276 net38 _064_ 0.02996f
C277 FILLER_0_19_28/a_124_375# net17 0.007234f
C278 _288_/a_224_472# net19 0.002252f
C279 _104_ _420_/a_2665_112# 0.053555f
C280 _413_/a_448_472# net21 0.052657f
C281 net23 FILLER_0_8_156/a_36_472# 0.004939f
C282 FILLER_0_16_107/a_484_472# net36 0.003765f
C283 _149_ _148_ 0.001124f
C284 _306_/a_36_68# _113_ 0.010109f
C285 FILLER_0_18_2/a_932_472# net38 0.020589f
C286 FILLER_0_8_2/a_36_472# net40 0.002477f
C287 output34/a_224_472# output18/a_224_472# 0.002121f
C288 net63 FILLER_0_18_177/a_2364_375# 0.009893f
C289 FILLER_0_5_54/a_36_472# net47 0.00679f
C290 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_36_472# 0.009654f
C291 net29 _005_ 0.020239f
C292 FILLER_0_19_55/a_36_472# FILLER_0_18_53/a_124_375# 0.001684f
C293 FILLER_0_9_72/a_932_472# vss 0.007033f
C294 FILLER_0_9_72/a_1380_472# vdd 0.007659f
C295 _028_ vss 0.410396f
C296 FILLER_0_12_124/a_124_375# _131_ 0.07304f
C297 net82 FILLER_0_3_172/a_36_472# 0.007612f
C298 _432_/a_36_151# _143_ 0.001486f
C299 _360_/a_36_160# _070_ 0.012463f
C300 net4 FILLER_0_12_236/a_124_375# 0.001558f
C301 _404_/a_36_472# vdd 0.034854f
C302 cal_itt\[3\] _076_ 0.002726f
C303 _414_/a_1308_423# net21 0.06986f
C304 _328_/a_36_113# vss 0.044028f
C305 net58 FILLER_0_8_247/a_1380_472# 0.0597f
C306 _185_ cal_count\[2\] 0.205002f
C307 _033_ trim_mask\[1\] 0.001251f
C308 _173_ _042_ 0.002294f
C309 FILLER_0_2_111/a_1468_375# _160_ 0.001026f
C310 fanout62/a_36_160# result[1] 0.036633f
C311 _094_ _418_/a_448_472# 0.042782f
C312 FILLER_0_17_72/a_1468_375# _150_ 0.001076f
C313 _137_ FILLER_0_16_154/a_484_472# 0.00631f
C314 _028_ FILLER_0_7_72/a_2812_375# 0.003873f
C315 _414_/a_2665_112# _075_ 0.050503f
C316 FILLER_0_9_28/a_124_375# net42 0.007403f
C317 output35/a_224_472# result[8] 0.016867f
C318 mask\[4\] FILLER_0_20_177/a_36_472# 0.001215f
C319 fanout52/a_36_160# vdd 0.026513f
C320 _114_ FILLER_0_12_124/a_124_375# 0.006974f
C321 net73 net36 0.073334f
C322 state\[0\] net4 0.13193f
C323 _119_ FILLER_0_8_127/a_124_375# 0.013315f
C324 mask\[9\] FILLER_0_20_87/a_36_472# 0.00596f
C325 fanout82/a_36_113# vss 0.023533f
C326 FILLER_0_16_89/a_1380_472# _136_ 0.009079f
C327 _328_/a_36_113# net74 0.002214f
C328 _132_ FILLER_0_11_109/a_36_472# 0.005748f
C329 net24 vdd 0.223761f
C330 _091_ _069_ 0.741596f
C331 _432_/a_36_151# _136_ 0.004543f
C332 _308_/a_848_380# vss 0.043591f
C333 _098_ FILLER_0_15_212/a_1380_472# 0.009972f
C334 FILLER_0_12_136/a_484_472# _126_ 0.014541f
C335 net52 trim_mask\[4\] 0.034276f
C336 _176_ _118_ 0.392531f
C337 _053_ FILLER_0_7_72/a_1020_375# 0.014569f
C338 _086_ net76 0.049988f
C339 _122_ FILLER_0_8_156/a_124_375# 0.032617f
C340 _024_ _147_ 0.006801f
C341 FILLER_0_20_15/a_572_375# vdd 0.003301f
C342 net15 FILLER_0_9_72/a_36_472# 0.006905f
C343 _141_ vss 0.308762f
C344 net82 cal_itt\[1\] 0.396149f
C345 fanout51/a_36_113# FILLER_0_9_72/a_36_472# 0.001391f
C346 _105_ output33/a_224_472# 0.099107f
C347 FILLER_0_17_72/a_1380_472# net36 0.021039f
C348 net52 FILLER_0_11_78/a_36_472# 0.005678f
C349 _099_ vdd 0.326559f
C350 _132_ FILLER_0_14_107/a_36_472# 0.002187f
C351 trim_mask\[2\] FILLER_0_3_78/a_124_375# 0.010185f
C352 _372_/a_2590_472# _059_ 0.002974f
C353 _392_/a_36_68# _039_ 0.001522f
C354 _008_ ctlp[1] 0.002566f
C355 FILLER_0_3_221/a_36_472# FILLER_0_3_212/a_36_472# 0.001963f
C356 FILLER_0_5_136/a_36_472# vss 0.007658f
C357 _281_/a_234_472# _097_ 0.004169f
C358 _257_/a_36_472# _068_ 0.002986f
C359 _127_ _125_ 0.053419f
C360 _077_ _449_/a_36_151# 0.002475f
C361 _422_/a_36_151# _109_ 0.036674f
C362 FILLER_0_21_28/a_3172_472# vss 0.001574f
C363 FILLER_0_6_90/a_36_472# vss 0.001409f
C364 FILLER_0_6_90/a_484_472# vdd 0.003146f
C365 valid net82 0.060784f
C366 _428_/a_36_151# vss 0.00285f
C367 _428_/a_448_472# vdd 0.034564f
C368 FILLER_0_15_142/a_124_375# net53 0.033224f
C369 FILLER_0_16_89/a_932_472# FILLER_0_17_72/a_2812_375# 0.001723f
C370 mask\[4\] FILLER_0_19_171/a_932_472# 0.004669f
C371 net66 net17 0.023639f
C372 ctln[2] FILLER_0_1_266/a_124_375# 0.047145f
C373 _430_/a_36_151# FILLER_0_17_200/a_36_472# 0.001723f
C374 _320_/a_1120_472# _090_ 0.001215f
C375 trimb[0] trimb[2] 0.00878f
C376 cal_itt\[2\] net82 0.663246f
C377 net74 FILLER_0_5_136/a_36_472# 0.003704f
C378 fanout68/a_36_113# FILLER_0_3_54/a_124_375# 0.015816f
C379 FILLER_0_7_72/a_2364_375# FILLER_0_6_90/a_484_472# 0.001684f
C380 _163_ FILLER_0_5_148/a_484_472# 0.002734f
C381 net37 FILLER_0_6_231/a_124_375# 0.001989f
C382 FILLER_0_8_263/a_36_472# net64 0.00399f
C383 _445_/a_1308_423# net17 0.002172f
C384 net81 _425_/a_2248_156# 0.058229f
C385 FILLER_0_15_116/a_36_472# net70 0.051129f
C386 _428_/a_36_151# net74 0.020444f
C387 fanout50/a_36_160# vss 0.009871f
C388 cal vss 0.424638f
C389 net57 _385_/a_36_68# 0.03315f
C390 output48/a_224_472# _425_/a_448_472# 0.001155f
C391 vdd _202_/a_36_160# 0.06338f
C392 _443_/a_448_472# vdd 0.007773f
C393 _443_/a_36_151# vss 0.019802f
C394 net48 _123_ 0.153061f
C395 _422_/a_36_151# _421_/a_2248_156# 0.001189f
C396 _432_/a_448_472# _091_ 0.050539f
C397 _074_ _265_/a_224_472# 0.001223f
C398 net55 _423_/a_36_151# 0.001124f
C399 _165_ FILLER_0_6_37/a_124_375# 0.002884f
C400 FILLER_0_7_72/a_1468_375# net52 0.003576f
C401 FILLER_0_7_72/a_572_375# net50 0.012932f
C402 _096_ net57 0.05086f
C403 net82 FILLER_0_2_171/a_124_375# 0.003818f
C404 vss _433_/a_2665_112# 0.035903f
C405 net75 _079_ 0.071974f
C406 output23/a_224_472# vdd 0.033718f
C407 _449_/a_2248_156# _176_ 0.013753f
C408 ctlp[5] vdd 0.293399f
C409 _091_ FILLER_0_18_209/a_484_472# 0.001212f
C410 FILLER_0_13_228/a_124_375# net4 0.002641f
C411 FILLER_0_16_255/a_36_472# net36 0.034335f
C412 FILLER_0_20_177/a_1468_375# _434_/a_2248_156# 0.001221f
C413 net52 FILLER_0_2_93/a_484_472# 0.009006f
C414 net50 FILLER_0_2_93/a_572_375# 0.00275f
C415 _088_ FILLER_0_3_212/a_36_472# 0.005583f
C416 net74 _443_/a_36_151# 0.003682f
C417 _059_ _242_/a_36_160# 0.001942f
C418 net79 FILLER_0_13_290/a_36_472# 0.038324f
C419 _449_/a_36_151# _453_/a_36_151# 0.007757f
C420 FILLER_0_12_124/a_124_375# _126_ 0.02249f
C421 net52 _448_/a_2248_156# 0.002555f
C422 cal_count\[3\] net14 0.028995f
C423 _067_ net17 0.17227f
C424 net55 _424_/a_1000_472# 0.001357f
C425 _020_ net73 0.057454f
C426 _065_ vdd 0.646511f
C427 _269_/a_36_472# _080_ 0.003981f
C428 _083_ _260_/a_36_68# 0.047191f
C429 net16 FILLER_0_18_37/a_124_375# 0.017482f
C430 _321_/a_1194_69# vss 0.0011f
C431 FILLER_0_2_177/a_572_375# vdd 0.022268f
C432 FILLER_0_2_177/a_124_375# vss 0.00252f
C433 _417_/a_2665_112# net62 0.006083f
C434 _058_ FILLER_0_8_156/a_484_472# 0.013955f
C435 _310_/a_49_472# _060_ 0.001122f
C436 FILLER_0_17_218/a_572_375# vss 0.078608f
C437 FILLER_0_17_218/a_36_472# vdd 0.084913f
C438 _139_ FILLER_0_15_180/a_572_375# 0.022254f
C439 FILLER_0_5_88/a_124_375# vdd 0.020896f
C440 net71 FILLER_0_22_107/a_572_375# 0.006403f
C441 FILLER_0_18_2/a_932_472# net55 0.012117f
C442 _154_ net14 0.02512f
C443 result[8] mask\[7\] 0.110637f
C444 FILLER_0_8_263/a_36_472# vss 0.001089f
C445 _072_ _070_ 2.141346f
C446 _418_/a_36_151# _417_/a_36_151# 0.005373f
C447 output11/a_224_472# _411_/a_36_151# 0.095813f
C448 _426_/a_2665_112# FILLER_0_8_239/a_124_375# 0.010736f
C449 FILLER_0_24_63/a_124_375# vss 0.03143f
C450 FILLER_0_24_63/a_36_472# vdd 0.055524f
C451 mask\[5\] FILLER_0_19_187/a_484_472# 0.007596f
C452 FILLER_0_20_31/a_36_472# vss 0.004923f
C453 _383_/a_36_472# vss 0.002794f
C454 _074_ _317_/a_36_113# 0.003383f
C455 FILLER_0_7_72/a_1916_375# FILLER_0_5_88/a_36_472# 0.0027f
C456 net16 FILLER_0_10_28/a_124_375# 0.002225f
C457 net54 FILLER_0_21_150/a_124_375# 0.007123f
C458 _433_/a_36_151# _145_ 0.004437f
C459 FILLER_0_5_128/a_484_472# FILLER_0_5_136/a_36_472# 0.013276f
C460 mask\[3\] _102_ 0.142836f
C461 FILLER_0_21_286/a_572_375# vdd 0.03062f
C462 FILLER_0_21_286/a_124_375# vss 0.005049f
C463 net79 FILLER_0_12_236/a_124_375# 0.010367f
C464 _045_ net62 0.029263f
C465 FILLER_0_4_144/a_572_375# net47 0.011686f
C466 clk rstn 0.541051f
C467 sample net18 0.103617f
C468 FILLER_0_10_78/a_572_375# cal_count\[3\] 0.002314f
C469 FILLER_0_5_198/a_572_375# net37 0.009149f
C470 _132_ _127_ 0.112364f
C471 _091_ FILLER_0_19_171/a_1020_375# 0.005708f
C472 net81 _426_/a_1308_423# 0.002332f
C473 _132_ FILLER_0_16_115/a_36_472# 0.015199f
C474 _413_/a_36_151# FILLER_0_3_172/a_1916_375# 0.059049f
C475 cal_count\[2\] _402_/a_1296_93# 0.022009f
C476 net44 FILLER_0_12_2/a_124_375# 0.01836f
C477 _137_ mask\[2\] 0.440828f
C478 _101_ _196_/a_36_160# 0.009836f
C479 _134_ FILLER_0_9_105/a_124_375# 0.005919f
C480 cal_count\[3\] FILLER_0_9_72/a_484_472# 0.004129f
C481 _448_/a_448_472# _037_ 0.044085f
C482 output20/a_224_472# ctlp[2] 0.085373f
C483 FILLER_0_4_123/a_36_472# _153_ 0.001419f
C484 _053_ _363_/a_244_472# 0.001236f
C485 fanout53/a_36_160# _136_ 0.001471f
C486 _069_ _161_ 0.017831f
C487 _077_ FILLER_0_9_60/a_572_375# 0.018665f
C488 FILLER_0_4_197/a_1020_375# net82 0.00123f
C489 _412_/a_2665_112# output37/a_224_472# 0.002025f
C490 _323_/a_36_113# FILLER_0_10_247/a_36_472# 0.00136f
C491 _012_ FILLER_0_23_44/a_484_472# 0.001572f
C492 _053_ FILLER_0_6_47/a_1828_472# 0.006408f
C493 _436_/a_2248_156# net35 0.014499f
C494 _441_/a_448_472# net66 0.023761f
C495 result[7] _419_/a_448_472# 0.021809f
C496 output34/a_224_472# _419_/a_2248_156# 0.022045f
C497 FILLER_0_16_89/a_1468_375# vss 0.048986f
C498 FILLER_0_16_89/a_36_472# vdd 0.040085f
C499 _081_ net22 0.103561f
C500 _257_/a_36_472# vdd -0.001779f
C501 net44 vdd 0.897202f
C502 net41 _452_/a_448_472# 0.052165f
C503 _417_/a_2560_156# net30 0.049334f
C504 net80 _146_ 0.021227f
C505 vdd _107_ 0.038236f
C506 _171_ vdd 0.038202f
C507 _430_/a_2248_156# _091_ 0.053571f
C508 _412_/a_2665_112# net5 0.042084f
C509 _181_ _401_/a_36_68# 0.010647f
C510 FILLER_0_21_142/a_572_375# net54 0.043619f
C511 FILLER_0_19_134/a_124_375# _145_ 0.023167f
C512 FILLER_0_15_142/a_36_472# fanout73/a_36_113# 0.009544f
C513 output35/a_224_472# _098_ 0.003653f
C514 _018_ mask\[1\] 0.001206f
C515 net49 _440_/a_1308_423# 0.022006f
C516 net25 net15 0.013745f
C517 output7/a_224_472# ctln[9] 0.001987f
C518 net19 net8 0.056454f
C519 ctln[5] ctln[6] 0.017291f
C520 ctln[1] FILLER_0_3_221/a_1020_375# 0.001554f
C521 output8/a_224_472# FILLER_0_3_221/a_1380_472# 0.001699f
C522 output32/a_224_472# _418_/a_36_151# 0.07368f
C523 _245_/a_234_472# net6 0.001301f
C524 net20 _078_ 0.105266f
C525 net15 net36 0.265646f
C526 net32 _419_/a_1308_423# 0.00191f
C527 _436_/a_2665_112# vss 0.007905f
C528 result[5] _419_/a_36_151# 0.006539f
C529 mask\[3\] _198_/a_67_603# 0.024102f
C530 net48 _305_/a_36_159# 0.059079f
C531 _415_/a_1204_472# net27 0.006198f
C532 FILLER_0_22_128/a_484_472# _433_/a_36_151# 0.001653f
C533 FILLER_0_4_197/a_1380_472# net59 0.022002f
C534 trimb[1] FILLER_0_20_2/a_124_375# 0.003431f
C535 output42/a_224_472# FILLER_0_8_2/a_124_375# 0.030009f
C536 calibrate net23 0.032259f
C537 vss _034_ 0.008249f
C538 _430_/a_2560_156# mask\[2\] 0.010268f
C539 _427_/a_36_151# FILLER_0_14_123/a_124_375# 0.023595f
C540 net21 net11 0.10869f
C541 _033_ _054_ 0.003394f
C542 net75 net64 0.037337f
C543 _270_/a_36_472# net22 0.002857f
C544 input3/a_36_113# net3 0.015124f
C545 output39/a_224_472# net49 0.039256f
C546 _011_ _299_/a_36_472# 0.004407f
C547 FILLER_0_17_104/a_124_375# vdd 0.030663f
C548 net55 FILLER_0_17_56/a_124_375# 0.014472f
C549 net72 FILLER_0_17_56/a_484_472# 0.003359f
C550 output7/a_224_472# vss 0.00746f
C551 FILLER_0_12_220/a_36_472# _248_/a_36_68# 0.006596f
C552 FILLER_0_5_54/a_572_375# FILLER_0_6_47/a_1380_472# 0.001597f
C553 _085_ vss 0.132721f
C554 _176_ vdd 0.874707f
C555 FILLER_0_16_73/a_572_375# FILLER_0_17_72/a_572_375# 0.026339f
C556 FILLER_0_16_73/a_36_472# FILLER_0_17_72/a_124_375# 0.001723f
C557 FILLER_0_5_164/a_572_375# vdd 0.0042f
C558 _414_/a_2665_112# net22 0.004067f
C559 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_572_375# 0.086635f
C560 output15/a_224_472# ctln[8] 0.079231f
C561 net20 net10 0.02842f
C562 _306_/a_36_68# vdd 0.044152f
C563 net63 output35/a_224_472# 0.148302f
C564 _341_/a_665_69# _141_ 0.001064f
C565 net82 net59 0.102279f
C566 trim[1] _445_/a_36_151# 0.008362f
C567 net39 _445_/a_1308_423# 0.008252f
C568 _220_/a_67_603# vdd 0.020078f
C569 _008_ _418_/a_2248_156# 0.047066f
C570 _335_/a_49_472# vdd 0.085394f
C571 FILLER_0_11_101/a_36_472# _070_ 0.033113f
C572 net52 FILLER_0_6_47/a_2276_472# 0.003298f
C573 net82 net4 1.982825f
C574 net38 FILLER_0_20_15/a_484_472# 0.003376f
C575 _018_ vss 0.022336f
C576 FILLER_0_13_228/a_124_375# net79 0.008554f
C577 ctlp[1] _421_/a_2665_112# 0.008695f
C578 _251_/a_906_472# vss 0.0016f
C579 fanout65/a_36_113# net64 0.002858f
C580 state\[2\] FILLER_0_13_142/a_1020_375# 0.007311f
C581 net53 FILLER_0_13_142/a_36_472# 0.059367f
C582 _442_/a_2665_112# vss 0.001727f
C583 _442_/a_2560_156# vdd 0.006195f
C584 net15 _160_ 0.046497f
C585 _425_/a_36_151# _316_/a_848_380# 0.035903f
C586 result[7] _420_/a_2665_112# 0.039448f
C587 _446_/a_2665_112# net17 0.00149f
C588 _036_ vdd 0.364747f
C589 _131_ _451_/a_3129_107# 0.001608f
C590 _144_ FILLER_0_19_125/a_36_472# 0.153815f
C591 net56 mask\[2\] 0.090254f
C592 net15 _423_/a_2560_156# 0.007083f
C593 net54 FILLER_0_19_142/a_124_375# 0.056556f
C594 _445_/a_2665_112# vdd 0.055628f
C595 result[9] net30 0.231442f
C596 FILLER_0_13_212/a_36_472# _429_/a_1308_423# 0.009119f
C597 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1380_472# 0.013276f
C598 _127_ _069_ 0.048146f
C599 _056_ _228_/a_36_68# 0.043669f
C600 FILLER_0_5_117/a_36_472# _153_ 0.028773f
C601 _076_ _081_ 0.010091f
C602 _133_ _152_ 0.124374f
C603 net52 _066_ 0.022601f
C604 vss output30/a_224_472# 0.030732f
C605 net75 vss 0.662689f
C606 mask\[4\] _201_/a_67_603# 0.029139f
C607 FILLER_0_6_90/a_124_375# _163_ 0.013948f
C608 net81 _005_ 0.003646f
C609 _091_ _090_ 0.117348f
C610 fanout61/a_36_113# ctlp[1] 0.019606f
C611 mask\[5\] FILLER_0_19_155/a_572_375# 0.007026f
C612 net73 FILLER_0_18_107/a_1916_375# 0.014643f
C613 FILLER_0_7_104/a_1380_472# _133_ 0.004838f
C614 trim_val\[3\] FILLER_0_2_93/a_36_472# 0.015653f
C615 FILLER_0_14_181/a_124_375# vdd 0.040138f
C616 _077_ _453_/a_2560_156# 0.001286f
C617 _430_/a_448_472# vss 0.003371f
C618 _430_/a_1308_423# vdd 0.00218f
C619 _425_/a_1204_472# vdd 0.015969f
C620 net64 FILLER_0_8_247/a_1468_375# 0.002559f
C621 _013_ _216_/a_67_603# 0.006454f
C622 mask\[7\] _435_/a_2560_156# 0.011544f
C623 _106_ _092_ 0.140596f
C624 net15 _030_ 0.355335f
C625 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_484_472# 0.026657f
C626 output36/a_224_472# _196_/a_36_160# 0.001309f
C627 _104_ vss 0.564464f
C628 FILLER_0_4_177/a_36_472# _386_/a_848_380# 0.007646f
C629 _061_ _055_ 0.853642f
C630 net65 FILLER_0_1_266/a_484_472# 0.004635f
C631 _122_ FILLER_0_6_231/a_124_375# 0.013183f
C632 _070_ FILLER_0_10_94/a_484_472# 0.003573f
C633 FILLER_0_8_24/a_572_375# net17 0.007101f
C634 output44/a_224_472# net38 0.106923f
C635 _056_ calibrate 0.00931f
C636 _426_/a_36_151# net64 0.022056f
C637 _094_ _006_ 0.090405f
C638 _091_ net22 0.031921f
C639 _420_/a_448_472# vdd 0.010071f
C640 _420_/a_36_151# vss 0.043027f
C641 net34 _422_/a_2248_156# 0.005617f
C642 _185_ _402_/a_56_567# 0.107713f
C643 fanout65/a_36_113# vss 0.053899f
C644 net26 net17 0.132516f
C645 trimb[2] net43 0.011999f
C646 _320_/a_672_472# vdd 0.008437f
C647 _098_ FILLER_0_15_180/a_572_375# 0.01526f
C648 _436_/a_2665_112# FILLER_0_22_128/a_1020_375# 0.029834f
C649 _091_ net81 0.03653f
C650 _057_ _176_ 0.001304f
C651 _415_/a_796_472# _004_ 0.005395f
C652 _013_ FILLER_0_18_37/a_572_375# 0.003828f
C653 net19 _419_/a_36_151# 0.009613f
C654 _057_ _306_/a_36_68# 0.019072f
C655 FILLER_0_21_125/a_572_375# vdd -0.013698f
C656 FILLER_0_10_78/a_1020_375# _389_/a_36_148# 0.001335f
C657 _093_ _099_ 0.001725f
C658 _003_ _087_ 0.054908f
C659 _089_ _079_ 0.126206f
C660 FILLER_0_18_139/a_484_472# FILLER_0_19_142/a_124_375# 0.001723f
C661 _449_/a_1308_423# _038_ 0.021006f
C662 FILLER_0_13_142/a_124_375# vdd 0.02675f
C663 net45 vdd 0.087369f
C664 FILLER_0_16_57/a_1468_375# _176_ 0.006445f
C665 FILLER_0_18_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001684f
C666 _410_/a_36_68# _173_ 0.009636f
C667 _339_/a_36_160# FILLER_0_19_171/a_36_472# 0.195478f
C668 _413_/a_36_151# FILLER_0_1_192/a_36_472# 0.046516f
C669 _183_ vdd 0.109252f
C670 _434_/a_2248_156# mask\[6\] 0.022666f
C671 mask\[4\] FILLER_0_19_187/a_36_472# 0.004669f
C672 _449_/a_36_151# _095_ 0.003412f
C673 result[9] _421_/a_1204_472# 0.014964f
C674 FILLER_0_17_72/a_2812_375# _136_ 0.017702f
C675 net61 FILLER_0_21_286/a_484_472# 0.001829f
C676 net16 _178_ 0.30147f
C677 fanout68/a_36_113# trim_mask\[2\] 0.003509f
C678 _082_ vdd 0.191411f
C679 net79 _416_/a_1204_472# 0.006493f
C680 net57 _374_/a_36_68# 0.001052f
C681 FILLER_0_8_247/a_1468_375# vss 0.054783f
C682 FILLER_0_8_247/a_36_472# vdd 0.112197f
C683 trim_mask\[4\] _152_ 0.224909f
C684 fanout77/a_36_113# vdd 0.032109f
C685 vss FILLER_0_6_37/a_124_375# 0.030885f
C686 vdd FILLER_0_6_37/a_36_472# 0.138008f
C687 _058_ _122_ 0.040376f
C688 net23 FILLER_0_22_128/a_2276_472# 0.011079f
C689 net63 mask\[7\] 0.069252f
C690 _070_ _133_ 0.436976f
C691 net20 net36 0.03843f
C692 FILLER_0_4_123/a_124_375# _160_ 0.038272f
C693 result[9] FILLER_0_15_282/a_124_375# 0.001233f
C694 net68 _042_ 0.037716f
C695 FILLER_0_10_214/a_36_472# _069_ 0.085701f
C696 FILLER_0_7_162/a_124_375# net57 0.033245f
C697 _426_/a_36_151# vss 0.003014f
C698 _426_/a_448_472# vdd 0.042167f
C699 cal_itt\[0\] net8 0.026229f
C700 _095_ FILLER_0_13_100/a_36_472# 0.003036f
C701 net82 FILLER_0_3_142/a_36_472# 0.0172f
C702 _430_/a_36_151# FILLER_0_18_177/a_2276_472# 0.001793f
C703 FILLER_0_16_37/a_124_375# cal_count\[2\] 0.008393f
C704 _446_/a_796_472# net40 0.001504f
C705 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_572_375# 0.086635f
C706 _074_ _375_/a_36_68# 0.003157f
C707 net80 _435_/a_448_472# 0.005274f
C708 ctlp[5] _147_ 0.001406f
C709 _064_ _446_/a_36_151# 0.006723f
C710 _235_/a_67_603# _446_/a_2665_112# 0.017036f
C711 _122_ FILLER_0_5_198/a_572_375# 0.001352f
C712 _187_ net51 0.04894f
C713 net20 ctln[4] 0.00225f
C714 _210_/a_255_603# vss 0.001246f
C715 _073_ _078_ 0.098575f
C716 _173_ _120_ 0.004205f
C717 net65 FILLER_0_3_172/a_36_472# 0.014671f
C718 _448_/a_448_472# FILLER_0_3_172/a_572_375# 0.00123f
C719 _448_/a_36_151# FILLER_0_3_172/a_1020_375# 0.001512f
C720 net17 FILLER_0_23_44/a_124_375# 0.007634f
C721 _436_/a_36_151# net24 0.075327f
C722 _013_ FILLER_0_18_61/a_124_375# 0.016976f
C723 FILLER_0_16_154/a_932_472# vdd 0.00549f
C724 FILLER_0_16_154/a_484_472# vss 0.003464f
C725 FILLER_0_3_172/a_2364_375# net21 0.004803f
C726 _412_/a_1204_472# cal_itt\[1\] 0.001547f
C727 FILLER_0_8_239/a_124_375# vss 0.017196f
C728 FILLER_0_8_239/a_36_472# vdd 0.079402f
C729 FILLER_0_11_101/a_484_472# FILLER_0_11_109/a_36_472# 0.013276f
C730 net69 FILLER_0_3_54/a_124_375# 0.004245f
C731 _141_ FILLER_0_17_142/a_572_375# 0.029028f
C732 _265_/a_244_68# vdd 0.022571f
C733 _061_ _058_ 0.02828f
C734 FILLER_0_12_136/a_1380_472# _076_ 0.001809f
C735 net19 _420_/a_2248_156# 0.058662f
C736 _076_ FILLER_0_9_142/a_124_375# 0.001774f
C737 FILLER_0_10_78/a_932_472# _439_/a_2665_112# 0.001182f
C738 net32 mask\[6\] 0.003248f
C739 _405_/a_67_603# net40 0.015326f
C740 _112_ vdd 0.086153f
C741 _415_/a_2248_156# net64 0.051575f
C742 FILLER_0_21_125/a_36_472# _140_ 0.101284f
C743 _093_ FILLER_0_17_218/a_36_472# 0.006994f
C744 fanout81/a_36_160# vss 0.02458f
C745 FILLER_0_7_104/a_36_472# vss 0.002797f
C746 FILLER_0_7_104/a_484_472# vdd 0.021325f
C747 output13/a_224_472# net23 0.00255f
C748 fanout64/a_36_160# vdd 0.010802f
C749 net81 FILLER_0_10_256/a_124_375# 0.026113f
C750 _120_ net14 0.024442f
C751 _436_/a_1000_472# _050_ 0.02064f
C752 output15/a_224_472# vdd 0.025731f
C753 FILLER_0_18_107/a_3260_375# vdd 0.004983f
C754 FILLER_0_18_107/a_2812_375# vss 0.002392f
C755 net65 cal_itt\[1\] 0.049124f
C756 _413_/a_1204_472# vdd 0.001027f
C757 _161_ _090_ 0.207838f
C758 result[1] FILLER_0_11_282/a_36_472# 0.01775f
C759 _346_/a_665_69# _141_ 0.002048f
C760 state\[1\] FILLER_0_13_142/a_1380_472# 0.006475f
C761 FILLER_0_14_107/a_124_375# _451_/a_36_151# 0.059049f
C762 vdd FILLER_0_10_94/a_124_375# 0.020076f
C763 _163_ _160_ 0.120564f
C764 _448_/a_1000_472# net22 0.011389f
C765 FILLER_0_16_89/a_124_375# _040_ 0.006315f
C766 mask\[8\] _354_/a_49_472# 0.105272f
C767 ctln[1] vdd 0.825166f
C768 FILLER_0_21_28/a_1468_375# _012_ 0.00351f
C769 _443_/a_2665_112# FILLER_0_2_165/a_124_375# 0.006271f
C770 _421_/a_2560_156# net19 0.006572f
C771 net57 FILLER_0_3_142/a_124_375# 0.003738f
C772 output44/a_224_472# net55 0.011586f
C773 FILLER_0_20_15/a_1380_472# net40 0.014911f
C774 output21/a_224_472# result[8] 0.149245f
C775 _053_ _439_/a_2665_112# 0.006037f
C776 FILLER_0_24_274/a_932_472# vss 0.001001f
C777 net65 valid 0.074257f
C778 _414_/a_2248_156# vdd 0.00901f
C779 ctln[2] net76 0.001008f
C780 FILLER_0_5_117/a_124_375# _160_ 0.008534f
C781 net45 output17/a_224_472# 0.01994f
C782 FILLER_0_4_49/a_484_472# _160_ 0.001336f
C783 FILLER_0_10_78/a_572_375# _120_ 0.006134f
C784 net65 cal_itt\[2\] 0.514538f
C785 net2 _082_ 0.034094f
C786 FILLER_0_5_164/a_484_472# net37 0.013857f
C787 FILLER_0_19_47/a_36_472# net26 0.050805f
C788 _008_ _199_/a_36_160# 0.002015f
C789 _025_ FILLER_0_22_107/a_484_472# 0.00892f
C790 _057_ _310_/a_741_69# 0.001002f
C791 _134_ FILLER_0_10_107/a_36_472# 0.006746f
C792 _093_ FILLER_0_16_89/a_36_472# 0.001338f
C793 _002_ net21 0.056631f
C794 output28/a_224_472# net18 0.015144f
C795 _053_ calibrate 0.081635f
C796 _415_/a_2665_112# vdd 0.017004f
C797 _415_/a_2248_156# vss 0.00818f
C798 net34 _023_ 0.00872f
C799 _162_ _118_ 0.005444f
C800 _120_ FILLER_0_9_72/a_484_472# 0.001645f
C801 _420_/a_2248_156# _009_ 0.00681f
C802 _016_ _427_/a_796_472# 0.001666f
C803 net67 net15 0.109181f
C804 FILLER_0_22_177/a_572_375# mask\[6\] 0.002657f
C805 _414_/a_36_151# net76 0.037157f
C806 _450_/a_1353_112# _039_ 0.019843f
C807 mask\[4\] FILLER_0_19_155/a_124_375# 0.043876f
C808 net52 net13 0.018118f
C809 _015_ calibrate 0.105287f
C810 _379_/a_244_68# _160_ 0.001202f
C811 net65 FILLER_0_2_171/a_124_375# 0.023202f
C812 FILLER_0_18_177/a_3260_375# net22 0.049279f
C813 net18 _416_/a_796_472# 0.007144f
C814 FILLER_0_8_138/a_36_472# _313_/a_67_603# 0.005759f
C815 _443_/a_1204_472# net23 0.026261f
C816 _449_/a_448_472# vdd 0.007757f
C817 _449_/a_36_151# vss 0.014774f
C818 _094_ _007_ 0.170362f
C819 _106_ FILLER_0_17_226/a_36_472# 0.050907f
C820 net50 _441_/a_2665_112# 0.056602f
C821 FILLER_0_13_65/a_36_472# _449_/a_36_151# 0.001723f
C822 net64 mask\[2\] 0.046428f
C823 _440_/a_1308_423# net47 0.009738f
C824 FILLER_0_12_220/a_484_472# vdd 0.002383f
C825 FILLER_0_12_220/a_36_472# vss 0.023702f
C826 _301_/a_36_472# FILLER_0_22_86/a_36_472# 0.010679f
C827 FILLER_0_4_49/a_36_472# net49 0.010951f
C828 FILLER_0_13_212/a_1380_472# net79 0.006824f
C829 FILLER_0_5_128/a_124_375# _152_ 0.017496f
C830 FILLER_0_5_128/a_572_375# _081_ 0.023853f
C831 FILLER_0_9_28/a_572_375# _054_ 0.002983f
C832 FILLER_0_21_125/a_36_472# _149_ 0.008849f
C833 net55 FILLER_0_18_37/a_1468_375# 0.009059f
C834 FILLER_0_4_107/a_932_472# _160_ 0.014254f
C835 mask\[2\] mask\[1\] 0.059794f
C836 net35 _434_/a_2248_156# 0.026885f
C837 FILLER_0_17_72/a_1020_375# vss 0.005441f
C838 FILLER_0_17_72/a_1468_375# vdd 0.003316f
C839 FILLER_0_8_37/a_484_472# vss 0.001267f
C840 _069_ _429_/a_448_472# 0.035108f
C841 FILLER_0_4_49/a_36_472# net68 0.00894f
C842 FILLER_0_11_142/a_36_472# FILLER_0_13_142/a_124_375# 0.0027f
C843 net58 net37 0.15273f
C844 net78 _420_/a_448_472# 0.001091f
C845 FILLER_0_21_142/a_36_472# FILLER_0_21_133/a_124_375# 0.007947f
C846 _093_ FILLER_0_17_104/a_124_375# 0.01418f
C847 net82 _443_/a_1308_423# 0.006706f
C848 _089_ vss 0.018272f
C849 net50 _439_/a_2248_156# 0.007461f
C850 _003_ vdd 0.032367f
C851 _321_/a_170_472# _176_ 0.059301f
C852 _449_/a_36_151# net74 0.032989f
C853 result[2] _416_/a_36_151# 0.010509f
C854 trimb[1] FILLER_0_18_2/a_1916_375# 0.001855f
C855 _095_ FILLER_0_14_107/a_1020_375# 0.014156f
C856 net57 fanout52/a_36_160# 0.122432f
C857 FILLER_0_8_127/a_36_472# _129_ 0.060819f
C858 _425_/a_2665_112# net37 0.008519f
C859 FILLER_0_22_86/a_124_375# vdd 0.024158f
C860 mask\[4\] FILLER_0_18_177/a_2724_472# 0.014625f
C861 FILLER_0_13_100/a_36_472# vss 0.003094f
C862 net38 _450_/a_1040_527# 0.027925f
C863 _116_ FILLER_0_12_196/a_124_375# 0.005332f
C864 result[9] _417_/a_2665_112# 0.060365f
C865 _131_ _332_/a_36_472# 0.006825f
C866 _010_ _420_/a_2560_156# 0.070902f
C867 net65 FILLER_0_2_165/a_124_375# 0.001177f
C868 _069_ net23 0.418375f
C869 _434_/a_2560_156# vdd 0.002922f
C870 _434_/a_2665_112# vss 0.00127f
C871 fanout73/a_36_113# _095_ 0.003989f
C872 clk net59 0.052607f
C873 _435_/a_36_151# _434_/a_1308_423# 0.001518f
C874 FILLER_0_18_107/a_572_375# net14 0.00258f
C875 FILLER_0_12_136/a_932_472# vdd 0.005266f
C876 FILLER_0_12_136/a_484_472# vss 0.007054f
C877 _422_/a_796_472# _009_ 0.001178f
C878 ctlp[1] FILLER_0_23_282/a_484_472# 0.007608f
C879 _417_/a_1000_472# vss 0.001822f
C880 output13/a_224_472# trim_val\[4\] 0.001014f
C881 net49 FILLER_0_3_78/a_484_472# 0.048729f
C882 _031_ FILLER_0_2_111/a_1380_472# 0.01562f
C883 net20 result[6] 0.026511f
C884 result[8] ctlp[2] 0.068359f
C885 _077_ FILLER_0_9_223/a_124_375# 0.008762f
C886 net25 _423_/a_2248_156# 0.005535f
C887 _092_ FILLER_0_18_209/a_572_375# 0.00609f
C888 _065_ _447_/a_2560_156# 0.012523f
C889 net74 FILLER_0_13_100/a_36_472# 0.003924f
C890 net36 FILLER_0_18_76/a_36_472# 0.001728f
C891 FILLER_0_12_136/a_572_375# _427_/a_1308_423# 0.001238f
C892 net13 _387_/a_36_113# 0.00189f
C893 net67 net51 0.010753f
C894 _114_ _332_/a_36_472# 0.021351f
C895 en_co_clk _172_ 0.025699f
C896 FILLER_0_15_142/a_124_375# net23 0.002212f
C897 _443_/a_2665_112# net59 0.0434f
C898 _161_ _076_ 0.042123f
C899 _017_ vdd 0.26981f
C900 FILLER_0_17_72/a_124_375# net15 0.006492f
C901 _411_/a_1308_423# net8 0.0176f
C902 net82 FILLER_0_2_177/a_36_472# 0.001777f
C903 cal_count\[2\] _452_/a_2225_156# 0.003086f
C904 net60 _421_/a_796_472# 0.002046f
C905 fanout77/a_36_113# net78 0.019286f
C906 mask\[2\] vss 0.536426f
C907 _437_/a_1000_472# vdd 0.001777f
C908 _441_/a_2560_156# _164_ 0.049213f
C909 ctln[1] net2 0.126801f
C910 net47 _365_/a_36_68# 0.020511f
C911 FILLER_0_8_138/a_36_472# _058_ 0.005325f
C912 net57 _428_/a_448_472# 0.032029f
C913 net61 _422_/a_36_151# 0.003736f
C914 _292_/a_36_160# _098_ 0.048643f
C915 _412_/a_36_151# net82 0.064296f
C916 FILLER_0_4_213/a_124_375# vss 0.006145f
C917 FILLER_0_4_213/a_572_375# vdd 0.026692f
C918 calibrate net18 0.014127f
C919 _308_/a_848_380# FILLER_0_9_105/a_124_375# 0.005599f
C920 _431_/a_2248_156# FILLER_0_15_142/a_572_375# 0.001374f
C921 net80 _141_ 0.077957f
C922 FILLER_0_22_177/a_124_375# _023_ 0.001195f
C923 FILLER_0_17_200/a_124_375# mask\[3\] 0.01841f
C924 output16/a_224_472# net16 0.054603f
C925 net47 FILLER_0_5_148/a_124_375# 0.008947f
C926 ctlp[4] mask\[7\] 0.080163f
C927 FILLER_0_1_192/a_124_375# net11 0.003537f
C928 _032_ vdd 0.174834f
C929 _250_/a_36_68# vdd 0.014409f
C930 result[7] vss 0.49466f
C931 _086_ FILLER_0_7_104/a_1468_375# 0.065371f
C932 FILLER_0_10_37/a_124_375# net51 0.006198f
C933 _273_/a_36_68# _090_ 0.034955f
C934 FILLER_0_23_44/a_36_472# vss 0.002194f
C935 FILLER_0_23_44/a_484_472# vdd 0.003276f
C936 output28/a_224_472# net62 0.206137f
C937 _144_ mask\[8\] 0.131592f
C938 FILLER_0_21_125/a_572_375# _433_/a_36_151# 0.059049f
C939 _141_ FILLER_0_18_139/a_1468_375# 0.005239f
C940 net53 FILLER_0_14_107/a_1380_472# 0.059367f
C941 net57 _443_/a_448_472# 0.001956f
C942 _302_/a_224_472# _012_ 0.002675f
C943 fanout63/a_36_160# _098_ 0.003627f
C944 _067_ FILLER_0_12_20/a_484_472# 0.011046f
C945 mask\[3\] FILLER_0_16_154/a_1020_375# 0.001996f
C946 _412_/a_1204_472# net59 0.001824f
C947 net72 FILLER_0_15_59/a_484_472# 0.008749f
C948 result[5] vdd 0.142481f
C949 _077_ FILLER_0_11_64/a_124_375# 0.013507f
C950 net48 _074_ 1.192591f
C951 _412_/a_2665_112# en 0.015256f
C952 mask\[5\] output19/a_224_472# 0.092961f
C953 _258_/a_36_160# net76 0.015203f
C954 _144_ vss 0.411237f
C955 net65 _411_/a_448_472# 0.006279f
C956 FILLER_0_7_104/a_1468_375# _154_ 0.003683f
C957 sample fanout59/a_36_160# 0.001854f
C958 output8/a_224_472# _078_ 0.001267f
C959 _430_/a_448_472# _019_ 0.019666f
C960 _422_/a_36_151# _108_ 0.062205f
C961 _091_ FILLER_0_18_177/a_932_472# 0.002113f
C962 FILLER_0_12_124/a_124_375# vss 0.012672f
C963 FILLER_0_12_124/a_36_472# vdd 0.040515f
C964 _370_/a_848_380# FILLER_0_5_136/a_124_375# 0.014613f
C965 _077_ _439_/a_1000_472# 0.030609f
C966 _091_ _140_ 0.006511f
C967 FILLER_0_9_60/a_36_472# vdd 0.08419f
C968 FILLER_0_9_60/a_572_375# vss 0.022532f
C969 _069_ _056_ 0.035189f
C970 net69 _369_/a_244_472# 0.002456f
C971 FILLER_0_10_214/a_36_472# _090_ 0.011963f
C972 FILLER_0_15_290/a_36_472# vss 0.010015f
C973 FILLER_0_22_86/a_484_472# FILLER_0_23_88/a_124_375# 0.001684f
C974 FILLER_0_3_172/a_932_472# net22 0.012284f
C975 _291_/a_36_160# mask\[4\] 0.00591f
C976 net65 net59 0.790496f
C977 _105_ mask\[6\] 0.029716f
C978 net66 _160_ 0.097885f
C979 _074_ FILLER_0_6_177/a_124_375# 0.003608f
C980 net63 fanout63/a_36_160# 0.011149f
C981 mask\[5\] FILLER_0_20_169/a_124_375# 0.011078f
C982 _343_/a_257_69# _141_ 0.001515f
C983 FILLER_0_12_124/a_124_375# net74 0.049113f
C984 _424_/a_1308_423# _012_ 0.007041f
C985 ctln[0] trim[2] 0.011834f
C986 net65 net4 0.614946f
C987 FILLER_0_7_72/a_124_375# vdd 0.01526f
C988 _126_ _332_/a_36_472# 0.009299f
C989 _127_ _076_ 0.137964f
C990 ctln[3] _411_/a_1000_472# 0.00283f
C991 cal_itt\[1\] FILLER_0_3_221/a_1468_375# 0.020427f
C992 _445_/a_36_151# _034_ 0.005488f
C993 trim_mask\[1\] _166_ 0.124855f
C994 net35 FILLER_0_22_177/a_572_375# 0.007797f
C995 net20 _317_/a_36_113# 0.00189f
C996 FILLER_0_11_109/a_124_375# vdd 0.079069f
C997 net20 FILLER_0_24_274/a_36_472# 0.009746f
C998 net54 net36 0.005827f
C999 _163_ _156_ 0.001616f
C1000 FILLER_0_10_214/a_36_472# net22 0.001634f
C1001 cal_count\[3\] _408_/a_1936_472# 0.007046f
C1002 FILLER_0_2_93/a_124_375# vdd 0.008901f
C1003 _077_ net4 0.656292f
C1004 FILLER_0_10_78/a_124_375# _115_ 0.001718f
C1005 _069_ FILLER_0_13_212/a_36_472# 0.047013f
C1006 cal_count\[2\] _182_ 0.044348f
C1007 FILLER_0_11_135/a_124_375# vdd 0.042201f
C1008 _399_/a_224_472# net16 0.003817f
C1009 FILLER_0_17_282/a_36_472# vss 0.007765f
C1010 _448_/a_796_472# vdd 0.002153f
C1011 FILLER_0_11_64/a_124_375# _453_/a_36_151# 0.005577f
C1012 ctln[7] ctln[8] 0.004643f
C1013 net38 _035_ 0.02987f
C1014 net75 _416_/a_2665_112# 0.001785f
C1015 _072_ _395_/a_36_488# 0.024944f
C1016 _088_ FILLER_0_3_172/a_3260_375# 0.002239f
C1017 FILLER_0_14_235/a_572_375# net62 0.017549f
C1018 FILLER_0_14_107/a_1468_375# vdd 0.007687f
C1019 _057_ _250_/a_36_68# 0.014333f
C1020 ctlp[1] FILLER_0_24_290/a_36_472# 0.037615f
C1021 _431_/a_1204_472# _137_ 0.005886f
C1022 net75 FILLER_0_10_247/a_36_472# 0.001184f
C1023 FILLER_0_22_177/a_1468_375# vdd -0.007187f
C1024 net66 _030_ 0.087608f
C1025 net41 _041_ 0.076779f
C1026 net69 _441_/a_1204_472# 0.014374f
C1027 trim_mask\[2\] net69 0.051795f
C1028 output31/a_224_472# net30 0.149277f
C1029 FILLER_0_3_172/a_124_375# FILLER_0_2_171/a_124_375# 0.026339f
C1030 _151_ net14 0.009212f
C1031 FILLER_0_5_109/a_572_375# vdd 0.024724f
C1032 cal_itt\[2\] FILLER_0_3_221/a_1468_375# 0.016021f
C1033 fanout73/a_36_113# vss 0.01873f
C1034 FILLER_0_16_37/a_36_472# _402_/a_728_93# 0.0108f
C1035 _321_/a_358_69# _121_ 0.00135f
C1036 _162_ vdd 0.073371f
C1037 _091_ _128_ 0.003717f
C1038 net71 _437_/a_2248_156# 0.025557f
C1039 net63 FILLER_0_17_218/a_484_472# 0.002672f
C1040 net41 _181_ 0.043679f
C1041 _445_/a_448_472# net49 0.00122f
C1042 _075_ _056_ 0.001957f
C1043 FILLER_0_7_72/a_2724_472# _077_ 0.004635f
C1044 _122_ FILLER_0_5_164/a_484_472# 0.002997f
C1045 _267_/a_36_472# _055_ 0.035376f
C1046 net34 FILLER_0_22_128/a_1916_375# 0.04185f
C1047 _128_ FILLER_0_9_142/a_124_375# 0.004439f
C1048 _430_/a_36_151# _432_/a_2665_112# 0.030053f
C1049 FILLER_0_9_28/a_2812_375# _077_ 0.006629f
C1050 _072_ _228_/a_36_68# 0.005788f
C1051 output9/a_224_472# net18 0.114757f
C1052 _327_/a_36_472# _428_/a_2248_156# 0.001757f
C1053 _273_/a_36_68# _076_ 0.001503f
C1054 net31 _104_ 0.102776f
C1055 _137_ FILLER_0_15_180/a_572_375# 0.028083f
C1056 net20 FILLER_0_12_220/a_1020_375# 0.047331f
C1057 _253_/a_244_68# _073_ 0.002878f
C1058 net52 FILLER_0_5_72/a_572_375# 0.024148f
C1059 _246_/a_36_68# _090_ 0.001712f
C1060 FILLER_0_22_128/a_36_472# _022_ 0.001541f
C1061 net76 net21 0.041873f
C1062 state\[0\] FILLER_0_12_220/a_932_472# 0.001003f
C1063 fanout73/a_36_113# net74 0.04136f
C1064 FILLER_0_15_235/a_572_375# FILLER_0_14_235/a_572_375# 0.05841f
C1065 _000_ net82 0.032846f
C1066 _079_ cal_itt\[1\] 0.012324f
C1067 FILLER_0_12_136/a_1380_472# FILLER_0_11_142/a_572_375# 0.001543f
C1068 _124_ _134_ 0.002508f
C1069 vss rstn 0.149553f
C1070 _205_/a_36_160# vdd 0.016131f
C1071 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_124_375# 0.007947f
C1072 FILLER_0_12_136/a_36_472# cal_count\[3\] 0.006102f
C1073 result[9] _418_/a_2665_112# 0.053489f
C1074 FILLER_0_18_177/a_2812_375# vdd 0.003766f
C1075 FILLER_0_21_206/a_124_375# _434_/a_2665_112# 0.002259f
C1076 _132_ _428_/a_1000_472# 0.027767f
C1077 _339_/a_36_160# vss 0.027338f
C1078 _372_/a_786_69# _163_ 0.001179f
C1079 _428_/a_1308_423# _131_ 0.037599f
C1080 net19 vdd 2.167778f
C1081 _093_ FILLER_0_18_107/a_3260_375# 0.008393f
C1082 _043_ net14 0.037706f
C1083 _418_/a_1000_472# vss 0.001193f
C1084 _411_/a_2560_156# net75 0.007047f
C1085 _076_ FILLER_0_8_156/a_572_375# 0.010751f
C1086 output9/a_224_472# _412_/a_1308_423# 0.001352f
C1087 net26 FILLER_0_21_28/a_2276_472# 0.001561f
C1088 _136_ _451_/a_1697_156# 0.001053f
C1089 ctln[5] FILLER_0_1_192/a_124_375# 0.001391f
C1090 _070_ net37 0.036662f
C1091 _072_ calibrate 0.539702f
C1092 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_124_375# 0.012001f
C1093 FILLER_0_23_88/a_124_375# vdd 0.03583f
C1094 FILLER_0_17_200/a_484_472# net21 0.017997f
C1095 _453_/a_2560_156# vss 0.00337f
C1096 _026_ _437_/a_796_472# 0.008884f
C1097 _149_ _437_/a_1204_472# 0.024276f
C1098 net41 _446_/a_1308_423# 0.056251f
C1099 cal_count\[3\] net47 0.043032f
C1100 net28 _426_/a_448_472# 0.00154f
C1101 net57 _176_ 0.192223f
C1102 _091_ state\[0\] 0.012343f
C1103 net75 _123_ 0.173358f
C1104 FILLER_0_9_223/a_36_472# _090_ 0.001057f
C1105 FILLER_0_18_107/a_3260_375# FILLER_0_19_134/a_124_375# 0.026339f
C1106 _439_/a_36_151# FILLER_0_6_47/a_2364_375# 0.002807f
C1107 net57 _306_/a_36_68# 0.042596f
C1108 cal_itt\[2\] _079_ 0.017071f
C1109 _126_ net79 0.085443f
C1110 _432_/a_36_151# _021_ 0.033849f
C1111 FILLER_0_15_212/a_1380_472# mask\[1\] 0.041503f
C1112 mask\[0\] FILLER_0_13_206/a_124_375# 0.005989f
C1113 _187_ _067_ 0.035532f
C1114 FILLER_0_13_142/a_36_472# net23 0.003007f
C1115 input2/a_36_113# vdd 0.096633f
C1116 _425_/a_2560_156# calibrate 0.010842f
C1117 net68 _120_ 0.001304f
C1118 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_124_375# 0.012001f
C1119 net47 _154_ 0.055128f
C1120 _053_ net50 0.711279f
C1121 result[2] net79 0.077934f
C1122 _103_ mask\[2\] 0.002168f
C1123 FILLER_0_13_212/a_484_472# net62 0.059367f
C1124 FILLER_0_1_266/a_484_472# vss 0.001113f
C1125 FILLER_0_1_204/a_124_375# net21 0.008041f
C1126 net18 FILLER_0_9_282/a_36_472# 0.041571f
C1127 _449_/a_2248_156# fanout55/a_36_160# 0.027388f
C1128 mask\[5\] FILLER_0_20_193/a_36_472# 0.013533f
C1129 FILLER_0_3_54/a_36_472# vdd 0.00827f
C1130 FILLER_0_9_28/a_2724_472# net68 0.010755f
C1131 net15 _453_/a_2248_156# 0.044493f
C1132 result[7] _103_ 0.298427f
C1133 FILLER_0_17_38/a_484_472# _182_ 0.00527f
C1134 _095_ FILLER_0_13_72/a_572_375# 0.003559f
C1135 net20 net34 0.003775f
C1136 net47 _169_ 0.528536f
C1137 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_124_375# 0.003732f
C1138 output44/a_224_472# FILLER_0_20_15/a_36_472# 0.0323f
C1139 _397_/a_36_472# _131_ 0.012338f
C1140 _325_/a_224_472# _129_ 0.003137f
C1141 FILLER_0_12_2/a_36_472# net67 0.013281f
C1142 output12/a_224_472# net59 0.015069f
C1143 vdd FILLER_0_16_115/a_124_375# 0.020393f
C1144 ctln[1] output11/a_224_472# 0.004299f
C1145 output10/a_224_472# ctln[2] 0.024524f
C1146 FILLER_0_6_47/a_932_472# vdd 0.003435f
C1147 net72 _052_ 0.138281f
C1148 net55 _217_/a_36_160# 0.001311f
C1149 FILLER_0_15_212/a_1380_472# vss 0.007595f
C1150 _429_/a_448_472# net22 0.054866f
C1151 _093_ FILLER_0_17_72/a_1468_375# 0.005785f
C1152 _337_/a_257_69# _137_ 0.001822f
C1153 _415_/a_2665_112# FILLER_0_9_290/a_124_375# 0.001597f
C1154 result[5] net78 0.020038f
C1155 result[5] net60 0.16275f
C1156 FILLER_0_19_47/a_572_375# FILLER_0_18_53/a_36_472# 0.001684f
C1157 _009_ vdd 0.693198f
C1158 FILLER_0_8_127/a_36_472# _322_/a_124_24# 0.00171f
C1159 FILLER_0_4_49/a_36_472# net47 0.002964f
C1160 FILLER_0_14_181/a_36_472# _098_ 0.004669f
C1161 _425_/a_36_151# FILLER_0_8_247/a_572_375# 0.001597f
C1162 net81 _429_/a_448_472# 0.018517f
C1163 _111_ vdd 0.3227f
C1164 _008_ _046_ 0.067769f
C1165 FILLER_0_4_197/a_36_472# net22 0.003404f
C1166 FILLER_0_4_197/a_1380_472# _081_ 0.001345f
C1167 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_124_375# 0.012001f
C1168 output38/a_224_472# output39/a_224_472# 0.002978f
C1169 FILLER_0_8_247/a_1380_472# calibrate 0.008605f
C1170 _178_ net3 0.257606f
C1171 net35 _051_ 0.019252f
C1172 _077_ FILLER_0_10_78/a_36_472# 0.002486f
C1173 output47/a_224_472# net3 0.002186f
C1174 trimb[4] input3/a_36_113# 0.001221f
C1175 _091_ FILLER_0_13_228/a_124_375# 0.001657f
C1176 _422_/a_1000_472# mask\[7\] 0.039617f
C1177 net52 _443_/a_2248_156# 0.045316f
C1178 FILLER_0_3_172/a_124_375# net59 0.001045f
C1179 trim[4] net44 0.188184f
C1180 net55 _038_ 0.05656f
C1181 en_co_clk _136_ 0.034892f
C1182 cal_count\[2\] FILLER_0_15_2/a_36_472# 0.037661f
C1183 _430_/a_448_472# net80 0.00896f
C1184 _426_/a_1000_472# calibrate 0.002865f
C1185 net4 _248_/a_36_68# 0.054512f
C1186 _162_ FILLER_0_5_172/a_36_472# 0.001501f
C1187 fanout78/a_36_113# vdd 0.061637f
C1188 fanout60/a_36_160# vdd 0.090968f
C1189 _446_/a_2665_112# _160_ 0.013745f
C1190 _379_/a_36_472# net47 0.016584f
C1191 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_124_375# 0.012267f
C1192 _055_ _113_ 0.153988f
C1193 _023_ _146_ 0.006636f
C1194 FILLER_0_16_241/a_36_472# FILLER_0_15_235/a_572_375# 0.001543f
C1195 _128_ _161_ 0.027657f
C1196 _102_ _419_/a_2248_156# 0.001679f
C1197 net2 net19 0.031976f
C1198 _453_/a_2248_156# net51 0.05329f
C1199 _363_/a_36_68# FILLER_0_5_109/a_36_472# 0.001024f
C1200 _426_/a_2665_112# net4 0.011288f
C1201 _402_/a_2172_497# cal_count\[1\] 0.008211f
C1202 net57 FILLER_0_13_142/a_124_375# 0.011369f
C1203 _421_/a_2665_112# net33 0.007127f
C1204 _415_/a_1204_472# result[1] 0.004051f
C1205 FILLER_0_16_89/a_484_472# _131_ 0.01075f
C1206 _177_ _040_ 0.061289f
C1207 _430_/a_796_472# net63 0.002914f
C1208 FILLER_0_4_107/a_484_472# net47 0.001975f
C1209 output24/a_224_472# net71 0.001495f
C1210 FILLER_0_21_125/a_36_472# _098_ 0.002923f
C1211 FILLER_0_18_171/a_124_375# FILLER_0_19_171/a_124_375# 0.05841f
C1212 net47 _278_/a_36_160# 0.001838f
C1213 FILLER_0_4_197/a_572_375# _088_ 0.013597f
C1214 FILLER_0_5_181/a_36_472# vss 0.001068f
C1215 FILLER_0_12_20/a_124_375# net47 0.047331f
C1216 _052_ _424_/a_36_151# 0.010844f
C1217 net4 _060_ 0.327437f
C1218 FILLER_0_21_28/a_1468_375# vdd -0.008892f
C1219 _304_/a_224_472# net15 0.001451f
C1220 FILLER_0_3_172/a_36_472# vss 0.001848f
C1221 FILLER_0_3_172/a_484_472# vdd 0.007258f
C1222 _386_/a_124_24# vss 0.009702f
C1223 _386_/a_848_380# vdd 0.054849f
C1224 valid net64 0.022969f
C1225 FILLER_0_9_223/a_36_472# _076_ 0.00146f
C1226 _053_ _075_ 0.634359f
C1227 vdd FILLER_0_8_156/a_124_375# 0.005213f
C1228 net4 FILLER_0_3_221/a_1468_375# 0.006974f
C1229 net75 _305_/a_36_159# 0.049563f
C1230 FILLER_0_8_239/a_124_375# _123_ 0.001286f
C1231 _091_ _139_ 0.05535f
C1232 _235_/a_67_603# net17 0.018056f
C1233 result[8] ctlp[1] 0.049662f
C1234 ctln[7] vdd 0.359832f
C1235 FILLER_0_18_100/a_124_375# vss 0.025563f
C1236 FILLER_0_18_100/a_36_472# vdd 0.012574f
C1237 input2/a_36_113# net2 0.015844f
C1238 _413_/a_2248_156# net82 0.009308f
C1239 net81 FILLER_0_14_235/a_124_375# 0.01391f
C1240 FILLER_0_18_2/a_1468_375# net17 0.004803f
C1241 net12 net59 0.001028f
C1242 _446_/a_2248_156# net49 0.006196f
C1243 net15 _168_ 0.04897f
C1244 _144_ _433_/a_448_472# 0.075144f
C1245 fanout49/a_36_160# _441_/a_2248_156# 0.027388f
C1246 net52 _170_ 0.378738f
C1247 FILLER_0_10_214/a_124_375# vdd 0.018944f
C1248 _005_ _416_/a_1204_472# 0.014873f
C1249 net50 _164_ 0.080818f
C1250 FILLER_0_19_195/a_36_472# _434_/a_2248_156# 0.001731f
C1251 FILLER_0_14_81/a_124_375# _451_/a_3129_107# 0.009542f
C1252 FILLER_0_7_59/a_572_375# FILLER_0_6_47/a_1916_375# 0.05841f
C1253 _118_ _055_ 0.042556f
C1254 _056_ _090_ 0.177189f
C1255 _132_ FILLER_0_17_104/a_1468_375# 0.051996f
C1256 net1 _265_/a_224_472# 0.005504f
C1257 _019_ mask\[2\] 0.155325f
C1258 _261_/a_36_160# FILLER_0_5_136/a_124_375# 0.003477f
C1259 net76 FILLER_0_3_172/a_1468_375# 0.039469f
C1260 net36 _195_/a_67_603# 0.034361f
C1261 _131_ FILLER_0_17_104/a_572_375# 0.003214f
C1262 _451_/a_2225_156# vdd 0.012404f
C1263 _451_/a_3129_107# vss 0.01f
C1264 ctln[1] _411_/a_2665_112# 0.004748f
C1265 FILLER_0_5_72/a_1380_472# trim_mask\[1\] 0.01221f
C1266 fanout58/a_36_160# vdd 0.101571f
C1267 _086_ state\[1\] 0.043298f
C1268 _176_ _129_ 0.036112f
C1269 cal_itt\[1\] vss 0.327626f
C1270 cal_itt\[0\] vdd 0.438996f
C1271 net33 net22 0.066751f
C1272 output21/a_224_472# ctlp[4] 0.052556f
C1273 _095_ net40 0.674445f
C1274 _059_ _163_ 0.038651f
C1275 _413_/a_3041_156# net59 0.001022f
C1276 net39 net17 0.099429f
C1277 fanout55/a_36_160# vdd 0.016488f
C1278 output18/a_224_472# output19/a_224_472# 0.00124f
C1279 net57 FILLER_0_16_154/a_932_472# 0.003453f
C1280 _425_/a_36_151# _317_/a_36_113# 0.002361f
C1281 _076_ net23 0.105196f
C1282 cal_count\[3\] state\[1\] 0.236393f
C1283 _079_ net59 0.102335f
C1284 FILLER_0_7_233/a_36_472# vss 0.005354f
C1285 net38 _452_/a_1353_112# 0.005918f
C1286 _014_ _122_ 0.001529f
C1287 _056_ net22 0.075673f
C1288 _008_ net18 0.113775f
C1289 _401_/a_36_68# vdd 0.003745f
C1290 _193_/a_36_160# vdd 0.092266f
C1291 net67 _067_ 0.151887f
C1292 _431_/a_796_472# net73 0.002306f
C1293 valid vss 0.308766f
C1294 mask\[3\] FILLER_0_18_177/a_1020_375# 0.002924f
C1295 FILLER_0_16_57/a_1468_375# _111_ 0.001371f
C1296 _098_ FILLER_0_16_154/a_1380_472# 0.00417f
C1297 _118_ _313_/a_67_603# 0.001793f
C1298 FILLER_0_12_28/a_36_472# _039_ 0.007926f
C1299 _079_ net4 0.023763f
C1300 net16 _233_/a_36_160# 0.01152f
C1301 output29/a_224_472# result[2] 0.058798f
C1302 _103_ _418_/a_1000_472# 0.006239f
C1303 _415_/a_36_151# net75 0.024047f
C1304 net41 FILLER_0_18_37/a_36_472# 0.007459f
C1305 _091_ _429_/a_1000_472# 0.029742f
C1306 net78 net19 0.507249f
C1307 net60 net19 0.102311f
C1308 cal_itt\[2\] vss 0.249871f
C1309 cal_count\[1\] _451_/a_3129_107# 0.028519f
C1310 mask\[5\] output18/a_224_472# 0.00133f
C1311 mask\[4\] net54 0.009909f
C1312 vdd FILLER_0_13_72/a_36_472# 0.108152f
C1313 vss FILLER_0_13_72/a_572_375# 0.061657f
C1314 trim_val\[4\] net22 0.144267f
C1315 _127_ _128_ 0.257374f
C1316 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_36_472# 0.012267f
C1317 _387_/a_36_113# _170_ 0.017801f
C1318 _340_/a_36_160# FILLER_0_20_169/a_124_375# 0.005494f
C1319 mask\[5\] _340_/a_36_160# 0.031249f
C1320 net58 FILLER_0_9_282/a_484_472# 0.091905f
C1321 FILLER_0_16_89/a_124_375# _177_ 0.008257f
C1322 output31/a_224_472# _417_/a_2665_112# 0.011048f
C1323 _164_ trim_mask\[3\] 0.016366f
C1324 _432_/a_1000_472# _091_ 0.026097f
C1325 net65 FILLER_0_1_212/a_124_375# 0.005253f
C1326 FILLER_0_8_127/a_124_375# _124_ 0.022175f
C1327 FILLER_0_13_212/a_36_472# net22 0.002402f
C1328 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_124_375# 0.012001f
C1329 FILLER_0_6_177/a_36_472# vss 0.001617f
C1330 FILLER_0_6_177/a_484_472# vdd 0.007991f
C1331 _321_/a_170_472# FILLER_0_11_135/a_124_375# 0.001153f
C1332 output48/a_224_472# net76 0.069862f
C1333 _068_ _055_ 0.443477f
C1334 FILLER_0_2_171/a_124_375# vss 0.049142f
C1335 net65 FILLER_0_2_177/a_36_472# 0.016652f
C1336 FILLER_0_2_171/a_36_472# vdd 0.029996f
C1337 net74 FILLER_0_13_72/a_572_375# 0.012891f
C1338 net55 FILLER_0_11_78/a_484_472# 0.038269f
C1339 output13/a_224_472# FILLER_0_0_130/a_124_375# 0.00363f
C1340 _242_/a_36_160# FILLER_0_5_164/a_124_375# 0.005705f
C1341 _114_ trim_mask\[0\] 0.021887f
C1342 _133_ calibrate 0.0188f
C1343 _070_ _122_ 0.153373f
C1344 net64 _416_/a_36_151# 0.013586f
C1345 fanout80/a_36_113# net81 0.097873f
C1346 net65 _412_/a_36_151# 0.015454f
C1347 vdd _047_ 0.175913f
C1348 net16 net55 0.035875f
C1349 FILLER_0_7_104/a_36_472# FILLER_0_9_105/a_124_375# 0.001188f
C1350 output35/a_224_472# vss 0.01667f
C1351 FILLER_0_4_144/a_36_472# _443_/a_36_151# 0.00271f
C1352 FILLER_0_4_123/a_36_472# _159_ 0.004956f
C1353 _274_/a_36_68# _072_ 0.001647f
C1354 FILLER_0_5_109/a_484_472# FILLER_0_4_107/a_572_375# 0.001684f
C1355 FILLER_0_4_197/a_1380_472# FILLER_0_4_213/a_36_472# 0.013277f
C1356 _033_ _444_/a_36_151# 0.014843f
C1357 _077_ cal_itt\[3\] 0.009816f
C1358 _068_ _311_/a_1212_473# 0.002835f
C1359 net79 _248_/a_36_68# 0.018243f
C1360 _104_ FILLER_0_23_274/a_124_375# 0.002159f
C1361 net31 result[7] 0.231528f
C1362 _427_/a_2248_156# _095_ 0.022479f
C1363 net68 FILLER_0_5_54/a_932_472# 0.013043f
C1364 _058_ _118_ 0.001451f
C1365 _324_/a_224_472# net74 0.001704f
C1366 _068_ _313_/a_67_603# 0.012208f
C1367 _273_/a_36_68# _128_ 0.005719f
C1368 net15 FILLER_0_23_60/a_124_375# 0.038706f
C1369 ctlp[3] _107_ 0.132316f
C1370 FILLER_0_2_165/a_36_472# vdd -0.003333f
C1371 FILLER_0_2_165/a_124_375# vss 0.008386f
C1372 FILLER_0_9_223/a_572_375# vdd 0.007158f
C1373 FILLER_0_9_223/a_124_375# vss 0.009569f
C1374 _445_/a_448_472# net47 0.005429f
C1375 _118_ _315_/a_36_68# 0.005792f
C1376 FILLER_0_14_123/a_36_472# _043_ 0.001782f
C1377 _420_/a_36_151# FILLER_0_23_274/a_124_375# 0.059049f
C1378 _451_/a_448_472# net14 0.04399f
C1379 _216_/a_67_603# _012_ 0.001014f
C1380 _369_/a_692_472# vdd 0.003899f
C1381 _076_ FILLER_0_6_231/a_572_375# 0.001647f
C1382 _069_ net62 0.010033f
C1383 net50 trim_val\[3\] 0.111824f
C1384 net82 FILLER_0_4_213/a_36_472# 0.003042f
C1385 _056_ _076_ 0.938912f
C1386 _061_ _070_ 0.02813f
C1387 net79 _060_ 0.019511f
C1388 _443_/a_1308_423# net69 0.004128f
C1389 _032_ _442_/a_36_151# 0.005632f
C1390 _443_/a_36_151# _031_ 0.014344f
C1391 fanout71/a_36_113# FILLER_0_20_107/a_124_375# 0.002853f
C1392 net78 _009_ 0.02395f
C1393 net60 _009_ 0.006086f
C1394 trim_mask\[2\] FILLER_0_4_91/a_484_472# 0.0022f
C1395 _093_ FILLER_0_18_177/a_2812_375# 0.001989f
C1396 net2 fanout58/a_36_160# 0.010424f
C1397 net29 net62 0.082455f
C1398 _086_ FILLER_0_5_181/a_124_375# 0.006872f
C1399 _415_/a_36_151# _426_/a_36_151# 0.002121f
C1400 _062_ net14 0.003317f
C1401 vss _416_/a_36_151# 0.044403f
C1402 output27/a_224_472# FILLER_0_9_282/a_572_375# 0.029138f
C1403 _429_/a_36_151# vdd 0.076815f
C1404 _114_ FILLER_0_13_142/a_572_375# 0.00191f
C1405 net35 _024_ 0.001335f
C1406 vdd net6 0.134918f
C1407 _079_ FILLER_0_5_198/a_124_375# 0.013896f
C1408 _095_ FILLER_0_13_80/a_124_375# 0.001989f
C1409 _128_ FILLER_0_10_214/a_36_472# 0.00186f
C1410 _398_/a_36_113# cal_count\[2\] 0.004895f
C1411 _178_ _405_/a_67_603# 0.02427f
C1412 net16 _447_/a_1000_472# 0.003207f
C1413 output16/a_224_472# _447_/a_2665_112# 0.005471f
C1414 fanout78/a_36_113# net78 0.004202f
C1415 fanout60/a_36_160# net60 0.019034f
C1416 net64 net59 0.005832f
C1417 FILLER_0_4_197/a_1020_375# vss 0.001981f
C1418 FILLER_0_4_197/a_1468_375# vdd 0.019672f
C1419 FILLER_0_18_171/a_124_375# _143_ 0.005331f
C1420 _273_/a_36_68# state\[0\] 0.012187f
C1421 mask\[1\] FILLER_0_15_180/a_572_375# 0.011186f
C1422 net4 net64 0.060449f
C1423 FILLER_0_22_86/a_572_375# _098_ 0.001139f
C1424 net18 result[3] 0.237732f
C1425 net58 net8 0.175026f
C1426 _449_/a_2665_112# FILLER_0_13_80/a_124_375# 0.010688f
C1427 vss net40 0.898805f
C1428 _424_/a_448_472# vss 0.002076f
C1429 _424_/a_1308_423# vdd 0.002386f
C1430 ctlp[1] _098_ 0.0012f
C1431 _072_ _069_ 0.265737f
C1432 net54 _437_/a_448_472# 0.004418f
C1433 _441_/a_2248_156# vdd -0.003818f
C1434 trim_val\[2\] vdd 0.160419f
C1435 _441_/a_1204_472# vss 0.011996f
C1436 trim_mask\[2\] vss 0.182675f
C1437 FILLER_0_11_64/a_124_375# vss 0.021069f
C1438 FILLER_0_11_64/a_36_472# vdd 0.015144f
C1439 _091_ _098_ 1.501073f
C1440 _444_/a_2665_112# trim_val\[0\] 0.007249f
C1441 _133_ _125_ 0.014858f
C1442 _068_ _058_ 0.092852f
C1443 _096_ cal_count\[3\] 0.016393f
C1444 net55 _452_/a_1353_112# 0.030679f
C1445 net57 _017_ 0.045694f
C1446 _015_ _426_/a_1204_472# 0.008883f
C1447 _447_/a_796_472# vdd 0.001959f
C1448 FILLER_0_22_128/a_2364_375# FILLER_0_21_150/a_36_472# 0.001543f
C1449 ctlp[0] net17 0.006778f
C1450 FILLER_0_18_2/a_3260_375# vss 0.026159f
C1451 FILLER_0_18_2/a_36_472# vdd 0.104532f
C1452 _068_ _315_/a_36_68# 0.003516f
C1453 _114_ FILLER_0_11_101/a_124_375# 0.013348f
C1454 trim_val\[3\] trim_mask\[3\] 0.48462f
C1455 _274_/a_244_497# net27 0.010334f
C1456 _431_/a_2248_156# vdd 0.00968f
C1457 _101_ _094_ 0.304499f
C1458 net76 FILLER_0_1_192/a_124_375# 0.00275f
C1459 _083_ _001_ 0.002625f
C1460 FILLER_0_18_177/a_1916_375# FILLER_0_19_195/a_36_472# 0.001684f
C1461 mask\[8\] mask\[7\] 0.021731f
C1462 _126_ FILLER_0_14_181/a_36_472# 0.008653f
C1463 _430_/a_1204_472# _069_ 0.001629f
C1464 _446_/a_36_151# _035_ 0.012914f
C1465 _439_/a_1000_472# vss 0.032923f
C1466 net34 net54 0.003682f
C1467 input3/a_36_113# vss 0.043862f
C1468 _091_ FILLER_0_13_212/a_1380_472# 0.003507f
C1469 _412_/a_1000_472# net58 0.030238f
C1470 mask\[8\] _148_ 0.356546f
C1471 _017_ _135_ 0.094281f
C1472 _443_/a_36_151# _371_/a_36_113# 0.001252f
C1473 _411_/a_448_472# vss 0.009447f
C1474 _176_ FILLER_0_10_107/a_572_375# 0.012296f
C1475 _098_ _437_/a_1204_472# 0.005729f
C1476 _053_ net22 0.039386f
C1477 _093_ FILLER_0_16_115/a_124_375# 0.003988f
C1478 _232_/a_67_603# _160_ 0.001684f
C1479 FILLER_0_7_104/a_932_472# _131_ 0.011713f
C1480 FILLER_0_21_125/a_124_375# _022_ 0.007023f
C1481 _402_/a_1948_68# _179_ 0.005403f
C1482 net57 _250_/a_36_68# 0.001141f
C1483 _055_ vdd 0.406945f
C1484 FILLER_0_4_152/a_124_375# net23 0.039975f
C1485 net17 net42 0.056318f
C1486 mask\[7\] vss 0.85153f
C1487 FILLER_0_15_180/a_572_375# vss 0.010974f
C1488 FILLER_0_15_180/a_36_472# vdd 0.017678f
C1489 net28 net19 0.115252f
C1490 _132_ FILLER_0_18_107/a_932_472# 0.001369f
C1491 net15 _441_/a_796_472# 0.021664f
C1492 net63 _091_ 0.767908f
C1493 net59 vss 1.191297f
C1494 mask\[5\] FILLER_0_20_177/a_1380_472# 0.016114f
C1495 FILLER_0_16_57/a_1020_375# net55 0.003303f
C1496 FILLER_0_16_57/a_484_472# net72 0.017841f
C1497 _148_ vss 0.025751f
C1498 _432_/a_448_472# FILLER_0_19_171/a_572_375# 0.00184f
C1499 net80 mask\[2\] 0.048734f
C1500 _190_/a_36_160# _450_/a_36_151# 0.002486f
C1501 _447_/a_36_151# net15 0.001598f
C1502 _093_ _111_ 0.555171f
C1503 net4 vss 0.774455f
C1504 _155_ _156_ 0.037229f
C1505 _128_ _246_/a_36_68# 0.01024f
C1506 _320_/a_36_472# _043_ 0.019162f
C1507 net65 _000_ 0.093773f
C1508 _086_ FILLER_0_6_177/a_572_375# 0.012909f
C1509 net81 _015_ 0.002818f
C1510 FILLER_0_15_10/a_124_375# vdd 0.021578f
C1511 FILLER_0_21_142/a_484_472# FILLER_0_22_128/a_1916_375# 0.001543f
C1512 net19 _416_/a_2248_156# 0.024466f
C1513 _311_/a_1212_473# vdd 0.001387f
C1514 _452_/a_836_156# net40 0.023204f
C1515 _428_/a_36_151# _451_/a_36_151# 0.003608f
C1516 _075_ _072_ 0.024301f
C1517 _077_ trim_mask\[0\] 0.090587f
C1518 net20 net48 0.035427f
C1519 net65 _425_/a_2248_156# 0.003451f
C1520 mask\[5\] FILLER_0_18_177/a_1020_375# 0.001604f
C1521 _313_/a_67_603# vdd -0.002183f
C1522 _254_/a_244_472# _074_ 0.002716f
C1523 _114_ FILLER_0_10_94/a_572_375# 0.008375f
C1524 output31/a_224_472# _418_/a_2665_112# 0.008243f
C1525 net36 FILLER_0_15_212/a_1468_375# 0.005276f
C1526 _430_/a_36_151# net21 0.019114f
C1527 net51 output6/a_224_472# 0.006462f
C1528 _435_/a_1000_472# vdd 0.032539f
C1529 _301_/a_36_472# _098_ 0.010091f
C1530 _119_ _324_/a_224_472# 0.00368f
C1531 output27/a_224_472# net18 0.058296f
C1532 _176_ FILLER_0_15_59/a_484_472# 0.007596f
C1533 _140_ net23 0.06742f
C1534 FILLER_0_18_171/a_36_472# _091_ 0.00395f
C1535 _370_/a_848_380# net47 0.004223f
C1536 vdd FILLER_0_6_231/a_124_375# 0.024542f
C1537 net16 _392_/a_36_68# 0.002191f
C1538 _427_/a_2248_156# vss 0.018484f
C1539 _427_/a_2665_112# vdd 0.033395f
C1540 FILLER_0_7_72/a_3172_472# vdd 0.003913f
C1541 _102_ _006_ 0.006115f
C1542 FILLER_0_15_282/a_36_472# net18 0.036858f
C1543 FILLER_0_4_177/a_124_375# net22 0.006125f
C1544 FILLER_0_9_223/a_36_472# _128_ 0.00702f
C1545 _164_ _382_/a_224_472# 0.011658f
C1546 FILLER_0_9_28/a_3260_375# vdd 0.017581f
C1547 FILLER_0_8_24/a_36_472# _054_ 0.007348f
C1548 vss FILLER_0_21_60/a_484_472# 0.004134f
C1549 _276_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C1550 fanout61/a_36_113# net18 0.001668f
C1551 _451_/a_1040_527# _040_ 0.007154f
C1552 FILLER_0_7_162/a_36_472# vss 0.006392f
C1553 _093_ FILLER_0_18_100/a_36_472# 0.077197f
C1554 _320_/a_36_472# net21 0.025762f
C1555 net52 FILLER_0_2_111/a_124_375# 0.00483f
C1556 _126_ FILLER_0_11_101/a_124_375# 0.011403f
C1557 net62 result[3] 0.451989f
C1558 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_124_375# 0.003732f
C1559 FILLER_0_8_138/a_36_472# _070_ 0.001342f
C1560 FILLER_0_8_37/a_124_375# _054_ 0.014206f
C1561 FILLER_0_22_177/a_1380_472# net33 0.016037f
C1562 net68 _453_/a_796_472# 0.001516f
C1563 FILLER_0_1_98/a_36_472# vdd 0.009937f
C1564 net72 cal_count\[3\] 0.059493f
C1565 _411_/a_2665_112# net19 0.00934f
C1566 FILLER_0_13_212/a_1468_375# vdd -0.013698f
C1567 FILLER_0_13_212/a_1020_375# vss 0.041631f
C1568 ctln[8] net52 0.005231f
C1569 net1 net5 0.266194f
C1570 _053_ _076_ 0.108358f
C1571 FILLER_0_6_177/a_124_375# _163_ 0.025831f
C1572 FILLER_0_20_107/a_124_375# net71 0.03452f
C1573 net32 _094_ 0.027571f
C1574 FILLER_0_17_72/a_1916_375# _131_ 0.006589f
C1575 net74 _332_/a_36_472# 0.003752f
C1576 FILLER_0_11_109/a_124_375# _135_ 0.009057f
C1577 _016_ FILLER_0_12_136/a_36_472# 0.016227f
C1578 _057_ _055_ 0.290639f
C1579 ctlp[2] _420_/a_2665_112# 0.01544f
C1580 FILLER_0_13_80/a_36_472# vdd 0.087291f
C1581 FILLER_0_13_80/a_124_375# vss 0.042254f
C1582 FILLER_0_5_72/a_484_472# net47 0.00169f
C1583 net81 net18 0.102876f
C1584 output40/a_224_472# output41/a_224_472# 0.292611f
C1585 _058_ vdd 0.511536f
C1586 net15 FILLER_0_21_60/a_572_375# 0.03167f
C1587 _448_/a_2665_112# trim_val\[4\] 0.004707f
C1588 _128_ net23 0.041791f
C1589 output36/a_224_472# _094_ 0.001477f
C1590 FILLER_0_24_130/a_36_472# output23/a_224_472# 0.001994f
C1591 net79 net64 0.049663f
C1592 _428_/a_1308_423# _095_ 0.001504f
C1593 FILLER_0_9_223/a_36_472# state\[0\] 0.002846f
C1594 net74 FILLER_0_13_80/a_124_375# 0.012889f
C1595 result[7] FILLER_0_24_274/a_124_375# 0.006125f
C1596 FILLER_0_14_91/a_36_472# _067_ 0.004194f
C1597 _272_/a_36_472# _089_ 0.003862f
C1598 _408_/a_56_524# net47 0.040511f
C1599 net79 mask\[1\] 0.029512f
C1600 mask\[7\] FILLER_0_22_128/a_1020_375# 0.035799f
C1601 _057_ _311_/a_1212_473# 0.004869f
C1602 net46 vss 0.110452f
C1603 _140_ net33 0.026401f
C1604 net24 FILLER_0_22_86/a_1380_472# 0.003096f
C1605 FILLER_0_5_198/a_572_375# vdd 0.005402f
C1606 _189_/a_67_603# FILLER_0_12_236/a_124_375# 0.00221f
C1607 _095_ FILLER_0_15_72/a_124_375# 0.001474f
C1608 net55 FILLER_0_21_28/a_3260_375# 0.006399f
C1609 net72 FILLER_0_21_28/a_932_472# 0.015756f
C1610 _412_/a_1308_423# net81 0.006961f
C1611 FILLER_0_11_142/a_572_375# net23 0.010863f
C1612 net80 FILLER_0_22_177/a_1020_375# 0.00258f
C1613 net53 _131_ 0.059223f
C1614 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_36_472# 0.086635f
C1615 net35 FILLER_0_22_128/a_484_472# 0.004578f
C1616 FILLER_0_15_150/a_124_375# mask\[2\] 0.002588f
C1617 _239_/a_36_160# net17 0.014703f
C1618 _126_ FILLER_0_10_94/a_572_375# 0.027249f
C1619 FILLER_0_8_24/a_124_375# net47 0.025599f
C1620 net36 _451_/a_1353_112# 0.01266f
C1621 _114_ FILLER_0_12_136/a_1380_472# 0.003953f
C1622 _437_/a_2665_112# FILLER_0_22_107/a_484_472# 0.007376f
C1623 net68 FILLER_0_6_47/a_1916_375# 0.00799f
C1624 mask\[0\] _018_ 0.328328f
C1625 _120_ _453_/a_2665_112# 0.002925f
C1626 FILLER_0_12_20/a_484_472# net17 0.05005f
C1627 _013_ _424_/a_1000_472# 0.037585f
C1628 FILLER_0_9_72/a_36_472# _439_/a_36_151# 0.001723f
C1629 output33/a_224_472# net19 0.12997f
C1630 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1380_472# 0.013276f
C1631 FILLER_0_3_142/a_36_472# vss 0.012379f
C1632 _094_ FILLER_0_17_282/a_124_375# 0.001151f
C1633 _114_ net53 0.001275f
C1634 fanout57/a_36_113# net22 0.024465f
C1635 _074_ _251_/a_906_472# 0.002887f
C1636 _106_ vdd 0.232973f
C1637 cal_itt\[3\] _079_ 0.015743f
C1638 FILLER_0_22_128/a_1380_472# vdd 0.005746f
C1639 FILLER_0_22_128/a_932_472# vss 0.003452f
C1640 net55 FILLER_0_17_64/a_124_375# 0.020021f
C1641 _444_/a_1000_472# vdd 0.004148f
C1642 _341_/a_49_472# net23 0.031763f
C1643 FILLER_0_16_73/a_572_375# _176_ 0.006454f
C1644 net50 _376_/a_36_160# 0.018407f
C1645 FILLER_0_9_28/a_1916_375# net51 0.001008f
C1646 FILLER_0_9_28/a_2364_375# _042_ 0.001216f
C1647 _035_ _164_ 0.056332f
C1648 _132_ fanout71/a_36_113# 0.055078f
C1649 FILLER_0_3_142/a_36_472# net74 0.001098f
C1650 FILLER_0_15_282/a_36_472# net62 0.013655f
C1651 _452_/a_36_151# _041_ 0.013289f
C1652 net79 vss 0.770834f
C1653 _150_ _136_ 0.039815f
C1654 FILLER_0_7_146/a_36_472# vss 0.029149f
C1655 _394_/a_1336_472# FILLER_0_13_72/a_124_375# 0.001597f
C1656 net26 FILLER_0_23_44/a_1020_375# 0.001646f
C1657 net75 _074_ 1.343862f
C1658 net80 _339_/a_36_160# 0.016897f
C1659 result[7] FILLER_0_23_274/a_124_375# 0.017938f
C1660 _233_/a_36_160# _063_ 0.002771f
C1661 net65 _413_/a_2248_156# 0.036792f
C1662 fanout61/a_36_113# net62 0.031315f
C1663 net22 FILLER_0_18_209/a_36_472# 0.018061f
C1664 vss trim[3] 0.235724f
C1665 _269_/a_36_472# net59 0.011985f
C1666 FILLER_0_10_78/a_36_472# vss 0.008832f
C1667 FILLER_0_10_78/a_484_472# vdd 0.004673f
C1668 trim[0] _064_ 0.014422f
C1669 _326_/a_36_160# _115_ 0.051266f
C1670 FILLER_0_19_28/a_36_472# net17 0.009277f
C1671 _428_/a_2665_112# net53 0.002379f
C1672 FILLER_0_21_28/a_484_472# net40 0.022617f
C1673 mask\[8\] FILLER_0_22_107/a_124_375# 0.015331f
C1674 _274_/a_716_497# net64 0.007904f
C1675 _327_/a_36_472# vdd 0.00142f
C1676 FILLER_0_17_200/a_484_472# FILLER_0_18_177/a_3172_472# 0.026657f
C1677 net4 _269_/a_36_472# 0.033296f
C1678 output42/a_224_472# vdd 0.04917f
C1679 FILLER_0_18_2/a_1828_472# net38 0.006713f
C1680 net20 _323_/a_36_113# 0.002161f
C1681 _033_ net49 0.003904f
C1682 FILLER_0_5_54/a_932_472# net47 0.006386f
C1683 _057_ _058_ 0.098076f
C1684 result[2] _005_ 0.060821f
C1685 FILLER_0_19_55/a_124_375# FILLER_0_18_53/a_484_472# 0.001684f
C1686 net82 FILLER_0_3_172/a_932_472# 0.007986f
C1687 FILLER_0_10_107/a_124_375# FILLER_0_10_94/a_572_375# 0.003228f
C1688 _128_ _056_ 0.026612f
C1689 net4 FILLER_0_12_236/a_36_472# 0.016315f
C1690 net38 net3 0.103189f
C1691 _150_ _356_/a_36_472# 0.007271f
C1692 ctln[7] _442_/a_36_151# 0.007057f
C1693 net75 FILLER_0_6_239/a_36_472# 0.009325f
C1694 FILLER_0_9_282/a_124_375# vdd 0.01273f
C1695 FILLER_0_12_220/a_1468_375# _043_ 0.002509f
C1696 vdd _167_ 0.012869f
C1697 net35 net24 0.01339f
C1698 FILLER_0_4_144/a_124_375# _081_ 0.004558f
C1699 _414_/a_1000_472# net21 0.042244f
C1700 _093_ _302_/a_224_472# 0.011376f
C1701 _185_ _184_ 0.047803f
C1702 vss FILLER_0_22_107/a_124_375# 0.002881f
C1703 vdd FILLER_0_22_107/a_572_375# 0.005745f
C1704 _094_ _418_/a_796_472# 0.005889f
C1705 FILLER_0_17_72/a_2364_375# _150_ 0.001083f
C1706 _086_ _374_/a_36_68# 0.009872f
C1707 _137_ FILLER_0_16_154/a_1380_472# 0.005667f
C1708 _028_ FILLER_0_7_72/a_36_472# 0.020625f
C1709 _414_/a_2665_112# _077_ 0.001675f
C1710 net81 net62 0.245647f
C1711 ctln[1] input5/a_36_113# 0.01908f
C1712 _253_/a_1100_68# _074_ 0.001563f
C1713 net43 FILLER_0_20_15/a_484_472# 0.001534f
C1714 fanout63/a_36_160# net64 0.016132f
C1715 net77 _007_ 0.002591f
C1716 _072_ _090_ 0.091468f
C1717 FILLER_0_15_282/a_572_375# result[3] 0.038939f
C1718 net52 _440_/a_36_151# 0.01571f
C1719 FILLER_0_13_100/a_124_375# _043_ 0.010818f
C1720 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_36_472# 0.016748f
C1721 fanout63/a_36_160# mask\[1\] 0.009907f
C1722 _119_ FILLER_0_7_162/a_36_472# 0.005739f
C1723 net38 _245_/a_672_472# 0.006341f
C1724 FILLER_0_12_136/a_1380_472# _126_ 0.014722f
C1725 _086_ _331_/a_448_472# 0.004356f
C1726 _189_/a_67_603# FILLER_0_13_228/a_124_375# 0.00744f
C1727 _053_ FILLER_0_7_72/a_1916_375# 0.013335f
C1728 _122_ FILLER_0_8_156/a_36_472# 0.047846f
C1729 _104_ _422_/a_2248_156# 0.041703f
C1730 mask\[4\] FILLER_0_18_177/a_572_375# 0.015941f
C1731 FILLER_0_20_15/a_1468_375# vdd 0.009742f
C1732 net50 FILLER_0_4_91/a_124_375# 0.022557f
C1733 _129_ FILLER_0_11_135/a_124_375# 0.009882f
C1734 _000_ FILLER_0_3_221/a_1468_375# 0.054354f
C1735 calibrate net37 0.101109f
C1736 _028_ net15 0.223301f
C1737 net57 _280_/a_224_472# 0.001032f
C1738 _069_ state\[2\] 0.023375f
C1739 FILLER_0_17_72/a_2276_472# net36 0.004399f
C1740 _130_ net53 0.00399f
C1741 _421_/a_2665_112# _109_ 0.002029f
C1742 _132_ FILLER_0_14_107/a_932_472# 0.014911f
C1743 FILLER_0_0_232/a_124_375# vdd 0.012494f
C1744 _441_/a_2248_156# FILLER_0_3_78/a_572_375# 0.001068f
C1745 output13/a_224_472# _448_/a_2248_156# 0.009013f
C1746 _423_/a_2248_156# FILLER_0_23_60/a_124_375# 0.001901f
C1747 _013_ FILLER_0_17_56/a_124_375# 0.001047f
C1748 trim_mask\[2\] FILLER_0_3_78/a_36_472# 0.005209f
C1749 _392_/a_244_472# cal_count\[0\] 0.003287f
C1750 _114_ FILLER_0_11_109/a_36_472# 0.023029f
C1751 _292_/a_36_160# vss 0.009517f
C1752 _072_ net22 0.147672f
C1753 net70 _043_ 0.045182f
C1754 _256_/a_716_497# net4 0.001936f
C1755 net81 FILLER_0_15_235/a_572_375# 0.009675f
C1756 _411_/a_2665_112# cal_itt\[0\] 0.010667f
C1757 _043_ net47 0.043824f
C1758 net32 output34/a_224_472# 0.027498f
C1759 _428_/a_796_472# vdd 0.003502f
C1760 net69 FILLER_0_2_127/a_124_375# 0.08337f
C1761 FILLER_0_15_142/a_36_472# net53 0.080484f
C1762 FILLER_0_16_89/a_1380_472# FILLER_0_17_72/a_3260_375# 0.001723f
C1763 ctln[2] FILLER_0_1_266/a_36_472# 0.052489f
C1764 _430_/a_1204_472# net22 0.028536f
C1765 _114_ FILLER_0_14_107/a_36_472# 0.00191f
C1766 _214_/a_36_160# vdd 0.010812f
C1767 output44/a_224_472# net43 0.001041f
C1768 net57 _386_/a_848_380# 0.041622f
C1769 FILLER_0_7_72/a_1828_472# _163_ 0.002095f
C1770 _185_ net47 0.185634f
C1771 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_36_472# 0.001723f
C1772 fanout76/a_36_160# vdd 0.108854f
C1773 _144_ _022_ 0.139742f
C1774 _369_/a_36_68# _158_ 0.042315f
C1775 net37 FILLER_0_6_231/a_36_472# 0.002982f
C1776 net57 FILLER_0_8_156/a_124_375# 0.001628f
C1777 FILLER_0_15_72/a_572_375# vdd 0.003801f
C1778 fanout63/a_36_160# vss 0.008974f
C1779 FILLER_0_15_72/a_124_375# vss 0.048711f
C1780 FILLER_0_12_2/a_36_472# output6/a_224_472# 0.00108f
C1781 net81 _425_/a_2560_156# 0.022037f
C1782 _428_/a_1308_423# net74 0.0098f
C1783 net21 _434_/a_2248_156# 0.001467f
C1784 FILLER_0_15_116/a_572_375# net53 0.012526f
C1785 net52 vdd 1.32956f
C1786 _114_ _161_ 0.024297f
C1787 _181_ _402_/a_1948_68# 0.001223f
C1788 _123_ FILLER_0_7_233/a_36_472# 0.002812f
C1789 net48 _425_/a_36_151# 0.020568f
C1790 _141_ FILLER_0_19_155/a_124_375# 0.029562f
C1791 _443_/a_1308_423# vss 0.031091f
C1792 _446_/a_2665_112# trim_val\[1\] 0.001275f
C1793 FILLER_0_7_162/a_124_375# _169_ 0.00336f
C1794 trim_val\[4\] _386_/a_1084_68# 0.002659f
C1795 FILLER_0_7_72/a_1468_375# net50 0.020186f
C1796 _000_ _079_ 0.032884f
C1797 mask\[3\] FILLER_0_17_200/a_484_472# 0.014805f
C1798 _028_ net51 0.002321f
C1799 net36 FILLER_0_15_228/a_124_375# 0.00167f
C1800 net27 _426_/a_448_472# 0.023676f
C1801 output22/a_224_472# _435_/a_448_472# 0.010723f
C1802 _431_/a_448_472# net36 0.010914f
C1803 _070_ _267_/a_36_472# 0.002617f
C1804 net50 FILLER_0_2_93/a_484_472# 0.002377f
C1805 _261_/a_36_160# net47 0.010976f
C1806 net48 net1 0.006424f
C1807 FILLER_0_3_204/a_124_375# FILLER_0_4_197/a_932_472# 0.001597f
C1808 FILLER_0_1_212/a_36_472# vdd 0.10765f
C1809 FILLER_0_1_212/a_124_375# vss 0.011796f
C1810 net16 _164_ 0.015161f
C1811 _216_/a_67_603# vdd 0.030831f
C1812 ctlp[7] net24 0.078667f
C1813 FILLER_0_15_72/a_124_375# cal_count\[1\] 0.00816f
C1814 net55 _424_/a_2248_156# 0.057967f
C1815 FILLER_0_6_239/a_124_375# FILLER_0_8_239/a_36_472# 0.001512f
C1816 net41 vdd 1.983262f
C1817 output21/a_224_472# vss 0.082781f
C1818 net16 FILLER_0_18_37/a_1020_375# 0.005406f
C1819 net57 fanout55/a_36_160# 0.017476f
C1820 FILLER_0_18_2/a_124_375# net44 0.051228f
C1821 _397_/a_36_472# vss 0.003673f
C1822 fanout50/a_36_160# net15 0.029852f
C1823 result[9] net29 0.001272f
C1824 FILLER_0_2_177/a_484_472# vdd 0.008489f
C1825 _132_ net71 0.099427f
C1826 FILLER_0_17_218/a_484_472# vss 0.035317f
C1827 net20 FILLER_0_1_204/a_36_472# 0.001278f
C1828 _139_ FILLER_0_15_180/a_484_472# 0.004763f
C1829 output47/a_224_472# trimb[4] 0.044883f
C1830 FILLER_0_5_88/a_36_472# vss 0.005793f
C1831 net71 FILLER_0_22_107/a_484_472# 0.00689f
C1832 FILLER_0_18_2/a_1828_472# net55 0.011802f
C1833 _153_ net14 0.260217f
C1834 FILLER_0_5_206/a_36_472# net59 0.060133f
C1835 output29/a_224_472# vss 0.013148f
C1836 ctlp[1] _419_/a_448_472# 0.020153f
C1837 cal_itt\[3\] vss 0.15522f
C1838 FILLER_0_14_181/a_36_472# _095_ 0.071989f
C1839 _412_/a_448_472# vdd 0.011f
C1840 _412_/a_36_151# vss 0.003515f
C1841 _072_ _076_ 0.068172f
C1842 _418_/a_1308_423# _417_/a_36_151# 0.001518f
C1843 _387_/a_36_113# vdd 0.041853f
C1844 _008_ result[9] 0.048497f
C1845 net46 FILLER_0_21_28/a_484_472# 0.001795f
C1846 _126_ FILLER_0_11_109/a_36_472# 0.00136f
C1847 _091_ _137_ 0.486022f
C1848 _406_/a_36_159# vdd 0.020825f
C1849 _433_/a_1308_423# _145_ 0.026613f
C1850 _414_/a_1204_472# _074_ 0.003142f
C1851 FILLER_0_18_37/a_124_375# vss 0.002958f
C1852 FILLER_0_18_37/a_572_375# vdd 0.02259f
C1853 FILLER_0_21_286/a_36_472# vss 0.004123f
C1854 FILLER_0_21_286/a_484_472# vdd 0.007903f
C1855 output45/a_224_472# net17 0.092967f
C1856 net79 FILLER_0_12_236/a_36_472# 0.009225f
C1857 net20 _080_ 0.093195f
C1858 FILLER_0_4_144/a_484_472# net47 0.008338f
C1859 _126_ FILLER_0_11_135/a_36_472# 0.002321f
C1860 FILLER_0_5_198/a_484_472# net37 0.009858f
C1861 FILLER_0_14_81/a_36_472# _394_/a_1936_472# 0.010394f
C1862 _346_/a_49_472# net23 0.022558f
C1863 _127_ _131_ 0.470047f
C1864 _091_ FILLER_0_19_171/a_36_472# 0.029168f
C1865 output44/a_224_472# _452_/a_448_472# 0.004683f
C1866 _050_ net14 0.001835f
C1867 net53 _137_ 0.008376f
C1868 _077_ FILLER_0_12_50/a_124_375# 0.008485f
C1869 result[8] net33 0.474056f
C1870 _413_/a_36_151# FILLER_0_3_172/a_2812_375# 0.059049f
C1871 _157_ _160_ 0.010231f
C1872 _131_ FILLER_0_16_115/a_36_472# 0.008241f
C1873 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_36_472# 0.086635f
C1874 cal_count\[2\] _402_/a_56_567# 0.07745f
C1875 _134_ FILLER_0_9_105/a_36_472# 0.004375f
C1876 FILLER_0_10_28/a_124_375# vss 0.013087f
C1877 FILLER_0_10_28/a_36_472# vdd 0.092132f
C1878 _448_/a_796_472# _037_ 0.009263f
C1879 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_124_375# 0.004426f
C1880 trim[0] _446_/a_448_472# 0.007307f
C1881 _053_ _363_/a_36_68# 0.021227f
C1882 _114_ _127_ 0.006414f
C1883 _077_ FILLER_0_9_60/a_484_472# 0.024249f
C1884 _012_ FILLER_0_23_44/a_1380_472# 0.001572f
C1885 _053_ FILLER_0_6_47/a_2724_472# 0.001777f
C1886 _436_/a_2560_156# net35 0.003198f
C1887 _441_/a_448_472# _030_ 0.038429f
C1888 _441_/a_36_151# net49 0.010951f
C1889 net82 net23 0.18994f
C1890 FILLER_0_16_89/a_932_472# vdd 0.002218f
C1891 FILLER_0_16_89/a_484_472# vss -0.001894f
C1892 _308_/a_124_24# FILLER_0_9_72/a_1468_375# 0.007188f
C1893 FILLER_0_18_2/a_2724_472# net40 0.011079f
C1894 _335_/a_257_69# mask\[1\] 0.001543f
C1895 ctlp[6] output24/a_224_472# 0.004288f
C1896 net68 _441_/a_36_151# 0.031891f
C1897 fanout76/a_36_160# net2 0.023033f
C1898 _172_ vdd 0.008764f
C1899 _430_/a_2560_156# _091_ 0.047345f
C1900 _445_/a_36_151# net40 0.007227f
C1901 FILLER_0_21_142/a_484_472# net54 0.038728f
C1902 FILLER_0_18_209/a_124_375# vss 0.004598f
C1903 FILLER_0_18_209/a_572_375# vdd 0.021356f
C1904 _040_ net14 0.069672f
C1905 net49 _440_/a_1000_472# 0.020434f
C1906 net9 net8 0.027272f
C1907 output36/a_224_472# FILLER_0_14_263/a_124_375# 0.029138f
C1908 _030_ _157_ 0.011014f
C1909 fanout74/a_36_113# net82 0.018392f
C1910 _067_ output6/a_224_472# 0.001611f
C1911 net68 _440_/a_1000_472# 0.002604f
C1912 _431_/a_448_472# _020_ 0.05255f
C1913 net57 FILLER_0_2_165/a_36_472# 0.001562f
C1914 _415_/a_2665_112# net27 0.030051f
C1915 ctlp[2] vss 0.131085f
C1916 fanout80/a_36_113# _139_ 0.009968f
C1917 _127_ _428_/a_2665_112# 0.001162f
C1918 FILLER_0_22_128/a_1380_472# _433_/a_36_151# 0.001973f
C1919 output23/a_224_472# FILLER_0_22_128/a_1468_375# 0.00242f
C1920 trimb[1] FILLER_0_20_2/a_36_472# 0.003628f
C1921 net72 _403_/a_224_472# 0.002276f
C1922 _440_/a_2248_156# trim_mask\[1\] 0.004408f
C1923 FILLER_0_11_109/a_36_472# FILLER_0_10_107/a_124_375# 0.001684f
C1924 output26/a_224_472# net26 0.047008f
C1925 FILLER_0_18_61/a_124_375# vdd 0.022663f
C1926 _028_ _163_ 0.199021f
C1927 _114_ _071_ 0.040513f
C1928 _178_ _095_ 0.839141f
C1929 trim[1] net66 0.007756f
C1930 _079_ _081_ 1.441057f
C1931 FILLER_0_17_104/a_1020_375# vdd 0.012531f
C1932 _174_ _179_ 0.003183f
C1933 net55 FILLER_0_17_56/a_36_472# 0.019193f
C1934 net7 vdd 0.321735f
C1935 FILLER_0_14_91/a_484_472# _043_ 0.00134f
C1936 FILLER_0_5_54/a_36_472# FILLER_0_6_47/a_932_472# 0.026657f
C1937 FILLER_0_5_54/a_1020_375# FILLER_0_6_47/a_1828_472# 0.001597f
C1938 output47/a_224_472# _095_ 0.012266f
C1939 state\[1\] _043_ 0.1587f
C1940 FILLER_0_16_73/a_484_472# FILLER_0_17_72/a_572_375# 0.001723f
C1941 FILLER_0_5_164/a_36_472# vss 0.001809f
C1942 FILLER_0_5_164/a_484_472# vdd 0.005235f
C1943 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_484_472# 0.013276f
C1944 FILLER_0_14_181/a_36_472# mask\[1\] 0.006352f
C1945 _106_ _093_ 0.045972f
C1946 _413_/a_448_472# _002_ 0.044695f
C1947 net39 _445_/a_1000_472# 0.007782f
C1948 _429_/a_36_151# FILLER_0_15_205/a_36_472# 0.001723f
C1949 _077_ _161_ 0.023053f
C1950 _010_ FILLER_0_23_274/a_36_472# 0.008718f
C1951 _008_ _418_/a_2560_156# 0.006651f
C1952 net47 _450_/a_2449_156# 0.004488f
C1953 net29 _287_/a_244_68# 0.001262f
C1954 net52 FILLER_0_6_47/a_3172_472# 0.047876f
C1955 FILLER_0_5_206/a_124_375# FILLER_0_5_198/a_572_375# 0.012001f
C1956 _070_ _113_ 0.01052f
C1957 _274_/a_1612_497# state\[0\] 0.001071f
C1958 comp input3/a_36_113# 0.022213f
C1959 FILLER_0_4_49/a_124_375# _167_ 0.009437f
C1960 FILLER_0_12_220/a_932_472# _060_ 0.002471f
C1961 _412_/a_448_472# net2 0.033994f
C1962 net18 FILLER_0_13_290/a_36_472# 0.079901f
C1963 FILLER_0_19_171/a_124_375# vdd -0.009473f
C1964 net67 net17 0.04175f
C1965 FILLER_0_21_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001723f
C1966 _427_/a_3041_156# net23 0.001305f
C1967 _377_/a_36_472# net67 0.005639f
C1968 state\[2\] FILLER_0_13_142/a_36_472# 0.022678f
C1969 net56 net53 0.053535f
C1970 net53 FILLER_0_13_142/a_932_472# 0.059367f
C1971 _303_/a_36_472# FILLER_0_20_87/a_36_472# 0.005725f
C1972 FILLER_0_18_107/a_2812_375# FILLER_0_17_133/a_36_472# 0.001543f
C1973 _091_ _248_/a_36_68# 0.071763f
C1974 net3 FILLER_0_15_10/a_36_472# 0.002825f
C1975 FILLER_0_15_235/a_124_375# vdd -0.006807f
C1976 _270_/a_36_472# _079_ 0.036715f
C1977 calibrate _122_ 0.074949f
C1978 FILLER_0_18_177/a_1916_375# net21 0.004339f
C1979 _098_ net23 0.036637f
C1980 FILLER_0_8_107/a_36_472# FILLER_0_7_104/a_484_472# 0.026657f
C1981 _163_ FILLER_0_5_136/a_36_472# 0.007779f
C1982 trim_mask\[0\] vss 0.014228f
C1983 _127_ _126_ 0.398279f
C1984 _068_ _152_ 0.006744f
C1985 _130_ _127_ 0.195571f
C1986 _414_/a_36_151# FILLER_0_6_177/a_572_375# 0.073306f
C1987 state\[1\] net21 0.210202f
C1988 _105_ output34/a_224_472# 0.007506f
C1989 vdd net30 0.636147f
C1990 _000_ vss 0.205593f
C1991 net58 vdd 0.929215f
C1992 FILLER_0_6_90/a_36_472# _163_ 0.016147f
C1993 _091_ _060_ 0.085764f
C1994 output20/a_224_472# _109_ 0.003452f
C1995 FILLER_0_2_93/a_572_375# net69 0.015032f
C1996 mask\[5\] FILLER_0_19_155/a_484_472# 0.043011f
C1997 net73 FILLER_0_18_107/a_2812_375# 0.018753f
C1998 _086_ _325_/a_224_472# 0.003155f
C1999 FILLER_0_7_72/a_2812_375# trim_mask\[0\] 0.005302f
C2000 FILLER_0_16_107/a_124_375# _136_ 0.00661f
C2001 FILLER_0_14_181/a_36_472# vss 0.002955f
C2002 _242_/a_36_160# _386_/a_124_24# 0.031797f
C2003 _425_/a_2665_112# vdd 0.012933f
C2004 _033_ net47 0.056436f
C2005 _069_ FILLER_0_11_142/a_124_375# 0.030279f
C2006 _070_ _118_ 0.302298f
C2007 net41 cal_count\[0\] 0.001014f
C2008 _119_ cal_itt\[3\] 0.010152f
C2009 net1 en 0.068102f
C2010 net82 trim_val\[4\] 0.511271f
C2011 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_932_472# 0.026657f
C2012 FILLER_0_20_98/a_124_375# vdd 0.0135f
C2013 net57 _055_ 0.008619f
C2014 _122_ FILLER_0_6_231/a_36_472# 0.015997f
C2015 FILLER_0_8_24/a_484_472# net17 0.010321f
C2016 _021_ _432_/a_796_472# 0.001666f
C2017 _115_ _134_ 0.051655f
C2018 _426_/a_1308_423# net64 0.021119f
C2019 _432_/a_2665_112# _337_/a_49_472# 0.001051f
C2020 _098_ FILLER_0_14_235/a_124_375# 0.001228f
C2021 _420_/a_1308_423# vss 0.001461f
C2022 input2/a_36_113# input5/a_36_113# 0.01088f
C2023 vss _450_/a_36_151# 0.02803f
C2024 vdd _450_/a_448_472# 0.011591f
C2025 _185_ _402_/a_718_527# 0.001973f
C2026 ctlp[3] _009_ 0.018168f
C2027 _126_ _071_ 0.090032f
C2028 net70 _451_/a_448_472# 0.043107f
C2029 fanout70/a_36_113# _136_ 0.002788f
C2030 _098_ FILLER_0_15_180/a_484_472# 0.014511f
C2031 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_124_375# 0.001597f
C2032 _415_/a_1204_472# _004_ 0.002391f
C2033 _013_ FILLER_0_18_37/a_1468_375# 0.017213f
C2034 output20/a_224_472# _422_/a_448_472# 0.009204f
C2035 net19 _419_/a_1308_423# 0.056469f
C2036 mask\[3\] FILLER_0_17_218/a_124_375# 0.016168f
C2037 _073_ _080_ 0.455535f
C2038 FILLER_0_21_125/a_36_472# vss 0.00143f
C2039 FILLER_0_21_125/a_484_472# vdd 0.002728f
C2040 _449_/a_1000_472# _038_ 0.021492f
C2041 FILLER_0_16_57/a_484_472# _176_ 0.013507f
C2042 FILLER_0_13_142/a_1020_375# vdd 0.018221f
C2043 trimb[2] vdd 0.084666f
C2044 FILLER_0_13_142/a_572_375# vss 0.04084f
C2045 _232_/a_67_603# trim_val\[1\] 0.009588f
C2046 net16 _378_/a_224_472# 0.001007f
C2047 FILLER_0_18_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001684f
C2048 _004_ _101_ 0.001514f
C2049 FILLER_0_9_142/a_36_472# _118_ 0.01533f
C2050 net80 mask\[7\] 0.020051f
C2051 net38 _190_/a_36_160# 0.062343f
C2052 _434_/a_2560_156# mask\[6\] 0.010913f
C2053 _008_ net61 0.004059f
C2054 ctlp[8] _051_ 0.010337f
C2055 net79 _416_/a_2665_112# 0.035115f
C2056 net57 _427_/a_2665_112# 0.016685f
C2057 FILLER_0_8_247/a_484_472# vss -0.001894f
C2058 FILLER_0_8_247/a_932_472# vdd 0.008645f
C2059 _421_/a_1204_472# vdd 0.002198f
C2060 trim_mask\[4\] net22 0.027368f
C2061 FILLER_0_7_59/a_572_375# trim_mask\[1\] 0.001548f
C2062 _331_/a_448_472# _120_ 0.001496f
C2063 net74 FILLER_0_13_142/a_572_375# 0.001412f
C2064 net23 FILLER_0_22_128/a_3172_472# 0.015058f
C2065 _133_ _076_ 0.11688f
C2066 _070_ _068_ 1.019801f
C2067 _258_/a_36_160# FILLER_0_7_233/a_124_375# 0.001633f
C2068 net34 _350_/a_49_472# 0.008001f
C2069 _422_/a_36_151# vdd 0.177717f
C2070 net55 _131_ 0.314732f
C2071 FILLER_0_13_290/a_36_472# net62 0.003157f
C2072 result[9] FILLER_0_15_282/a_36_472# 0.003213f
C2073 ctln[5] net11 0.004569f
C2074 cal_count\[3\] _171_ 0.00961f
C2075 net52 FILLER_0_2_101/a_36_472# 0.00749f
C2076 _426_/a_796_472# vdd 0.007178f
C2077 _084_ net8 0.001821f
C2078 trim_mask\[1\] net14 0.024935f
C2079 _096_ _043_ 0.842762f
C2080 _430_/a_36_151# FILLER_0_18_177/a_3172_472# 0.001512f
C2081 FILLER_0_15_282/a_124_375# vdd 0.011964f
C2082 _446_/a_1204_472# net40 0.026414f
C2083 trim[4] net6 0.002404f
C2084 _436_/a_36_151# FILLER_0_22_107/a_572_375# 0.059049f
C2085 _178_ vss 0.150839f
C2086 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_484_472# 0.013276f
C2087 FILLER_0_11_101/a_572_375# vdd 0.023482f
C2088 _064_ _446_/a_1308_423# 0.001728f
C2089 _157_ _156_ 0.005264f
C2090 _122_ FILLER_0_5_198/a_484_472# 0.002999f
C2091 output47/a_224_472# vss 0.002843f
C2092 _091_ _095_ 0.005006f
C2093 net10 ctln[4] 0.1323f
C2094 _088_ FILLER_0_4_213/a_572_375# 0.022684f
C2095 FILLER_0_17_104/a_1380_472# FILLER_0_16_115/a_124_375# 0.001723f
C2096 _305_/a_36_159# net59 0.007898f
C2097 net63 net33 0.048496f
C2098 net67 _439_/a_36_151# 0.136402f
C2099 _438_/a_36_151# net71 0.053065f
C2100 _332_/a_244_68# _135_ 0.001325f
C2101 net65 FILLER_0_3_172/a_932_472# 0.002604f
C2102 _086_ _176_ 0.837546f
C2103 output11/a_224_472# FILLER_0_0_232/a_124_375# 0.00515f
C2104 net58 net2 0.070564f
C2105 _315_/a_244_497# _120_ 0.006419f
C2106 _412_/a_2248_156# fanout58/a_36_160# 0.005856f
C2107 FILLER_0_16_154/a_1380_472# vss 0.003609f
C2108 net53 _095_ 0.431214f
C2109 _412_/a_2665_112# cal_itt\[1\] 0.015571f
C2110 FILLER_0_3_172/a_3260_375# net21 0.049606f
C2111 fanout80/a_36_113# _098_ 0.011559f
C2112 net19 _196_/a_36_160# 0.027835f
C2113 _141_ FILLER_0_17_142/a_484_472# 0.004527f
C2114 _408_/a_728_93# net40 0.084147f
C2115 net19 _420_/a_2560_156# 0.010978f
C2116 net57 _058_ 0.028536f
C2117 _176_ cal_count\[3\] 0.067683f
C2118 _152_ vdd 0.354509f
C2119 _081_ vss 0.733408f
C2120 _068_ FILLER_0_9_142/a_36_472# 0.009073f
C2121 _221_/a_36_160# net40 0.002952f
C2122 net57 _315_/a_36_68# 0.0036f
C2123 _306_/a_36_68# cal_count\[3\] 0.007663f
C2124 net39 net67 0.049482f
C2125 _077_ FILLER_0_8_156/a_572_375# 0.007238f
C2126 _372_/a_170_472# net23 0.025555f
C2127 _178_ cal_count\[1\] 0.470244f
C2128 _415_/a_2560_156# net64 0.066438f
C2129 _075_ net37 0.001054f
C2130 FILLER_0_7_104/a_1380_472# vdd 0.011752f
C2131 output13/a_224_472# net13 0.058196f
C2132 _072_ _128_ 0.072191f
C2133 FILLER_0_14_99/a_36_472# net14 0.036527f
C2134 FILLER_0_17_56/a_124_375# _041_ 0.001489f
C2135 FILLER_0_3_78/a_124_375# _164_ 0.023555f
C2136 net74 _081_ 0.093806f
C2137 _318_/a_224_472# vdd 0.001873f
C2138 _436_/a_2248_156# _050_ 0.023725f
C2139 _043_ FILLER_0_13_72/a_124_375# 0.013517f
C2140 _038_ FILLER_0_11_78/a_36_472# 0.001782f
C2141 FILLER_0_18_107/a_484_472# vdd 0.035309f
C2142 FILLER_0_18_107/a_36_472# vss 0.003245f
C2143 FILLER_0_2_127/a_36_472# vdd 0.08468f
C2144 FILLER_0_2_127/a_124_375# vss 0.008566f
C2145 net64 _005_ 0.006192f
C2146 FILLER_0_19_195/a_36_472# _202_/a_36_160# 0.002647f
C2147 _114_ net23 0.029535f
C2148 _413_/a_2248_156# vss 0.004157f
C2149 _413_/a_2665_112# vdd 0.02286f
C2150 _161_ _060_ 0.042838f
C2151 vss FILLER_0_10_94/a_572_375# 0.013232f
C2152 vdd FILLER_0_10_94/a_36_472# 0.086035f
C2153 _143_ vdd 0.074199f
C2154 _448_/a_2248_156# net22 0.07925f
C2155 net54 FILLER_0_22_128/a_36_472# 0.020739f
C2156 FILLER_0_18_139/a_36_472# _145_ 0.002415f
C2157 _005_ mask\[1\] 0.246517f
C2158 FILLER_0_16_89/a_1020_375# _040_ 0.004252f
C2159 _348_/a_49_472# vdd 0.038046f
C2160 _417_/a_448_472# _006_ 0.068545f
C2161 FILLER_0_16_37/a_124_375# net47 0.002638f
C2162 output15/a_224_472# FILLER_0_0_96/a_124_375# 0.00515f
C2163 trim_val\[0\] vdd 0.056059f
C2164 trim_mask\[4\] _076_ 0.001824f
C2165 FILLER_0_21_28/a_2364_375# _012_ 0.017669f
C2166 _421_/a_448_472# net77 0.003958f
C2167 _292_/a_36_160# net31 0.010041f
C2168 net16 _186_ 0.225785f
C2169 _014_ vdd 0.035382f
C2170 _010_ _419_/a_1000_472# 0.001598f
C2171 net69 _367_/a_244_472# 0.001708f
C2172 _442_/a_2248_156# _153_ 0.0011f
C2173 net74 FILLER_0_2_127/a_124_375# 0.001389f
C2174 net27 net19 0.036883f
C2175 _414_/a_2665_112# vss 0.010021f
C2176 net68 fanout67/a_36_160# 0.02648f
C2177 FILLER_0_5_164/a_124_375# _163_ 0.048663f
C2178 _063_ _164_ 0.326812f
C2179 _144_ net73 0.003657f
C2180 trimb[2] output17/a_224_472# 0.008375f
C2181 output45/a_224_472# ctlp[0] 0.007867f
C2182 FILLER_0_8_138/a_36_472# calibrate 0.047835f
C2183 _413_/a_448_472# net76 0.029504f
C2184 _136_ vdd 1.020301f
C2185 _092_ _069_ 0.040267f
C2186 fanout72/a_36_113# _095_ 0.001842f
C2187 _149_ FILLER_0_20_98/a_36_472# 0.067283f
C2188 _093_ FILLER_0_16_89/a_932_472# 0.002018f
C2189 _091_ net64 0.079488f
C2190 state\[0\] _072_ 0.030642f
C2191 net72 FILLER_0_17_38/a_572_375# 0.010272f
C2192 fanout82/a_36_113# _425_/a_36_151# 0.030783f
C2193 _415_/a_2560_156# vss 0.001286f
C2194 net36 FILLER_0_20_87/a_124_375# 0.005853f
C2195 net20 net75 0.092951f
C2196 net60 net30 0.001168f
C2197 ctln[3] FILLER_0_0_266/a_36_472# 0.012298f
C2198 _091_ mask\[1\] 0.064614f
C2199 _120_ FILLER_0_9_72/a_1380_472# 0.001723f
C2200 _420_/a_2560_156# _009_ 0.001487f
C2201 FILLER_0_22_177/a_1468_375# mask\[6\] 0.002149f
C2202 _093_ FILLER_0_18_209/a_572_375# 0.064723f
C2203 net72 _043_ 0.05655f
C2204 mask\[4\] FILLER_0_19_155/a_36_472# 0.047448f
C2205 _450_/a_836_156# _039_ 0.019042f
C2206 _430_/a_36_151# mask\[3\] 0.005848f
C2207 net22 _048_ 0.268142f
C2208 _431_/a_36_151# net70 0.031018f
C2209 trim_mask\[1\] FILLER_0_6_90/a_572_375# 0.001263f
C2210 _005_ vss 0.01812f
C2211 _104_ _291_/a_36_160# 0.006129f
C2212 net18 _416_/a_1204_472# 0.027218f
C2213 _070_ vdd 1.546772f
C2214 _021_ FILLER_0_18_171/a_124_375# 0.004621f
C2215 _449_/a_1308_423# vss 0.027539f
C2216 net20 _104_ 0.482229f
C2217 _356_/a_36_472# vdd 0.016338f
C2218 _440_/a_1000_472# net47 0.011283f
C2219 FILLER_0_12_220/a_932_472# vss 0.003677f
C2220 FILLER_0_12_220/a_1380_472# vdd 0.002025f
C2221 net35 FILLER_0_22_86/a_124_375# 0.01209f
C2222 mask\[8\] FILLER_0_22_86/a_572_375# 0.013048f
C2223 FILLER_0_15_150/a_124_375# _427_/a_2248_156# 0.001221f
C2224 net52 _442_/a_36_151# 0.029373f
C2225 FILLER_0_5_128/a_36_472# _152_ 0.013822f
C2226 FILLER_0_5_128/a_484_472# _081_ 0.00169f
C2227 FILLER_0_9_28/a_1468_375# _054_ 0.005381f
C2228 _093_ FILLER_0_18_61/a_124_375# 0.031062f
C2229 net55 FILLER_0_18_37/a_484_472# 0.006153f
C2230 net50 _447_/a_2248_156# 0.007602f
C2231 _114_ _311_/a_1660_473# 0.003304f
C2232 _077_ _246_/a_36_68# 0.006077f
C2233 net32 _011_ 0.072502f
C2234 FILLER_0_17_72/a_2364_375# vdd 0.002455f
C2235 FILLER_0_17_72/a_1916_375# vss 0.001345f
C2236 FILLER_0_11_142/a_484_472# FILLER_0_13_142/a_572_375# 0.0027f
C2237 _174_ _181_ 0.079407f
C2238 _069_ _429_/a_796_472# 0.003099f
C2239 FILLER_0_16_89/a_572_375# net36 0.003629f
C2240 _093_ FILLER_0_17_104/a_1020_375# 0.01418f
C2241 net82 _443_/a_1000_472# 0.008161f
C2242 net50 _439_/a_2560_156# 0.006321f
C2243 _321_/a_2590_472# _176_ 0.001932f
C2244 _069_ _395_/a_1044_488# 0.002244f
C2245 output29/a_224_472# _416_/a_2665_112# 0.011048f
C2246 _095_ FILLER_0_14_107/a_36_472# 0.011439f
C2247 _105_ _204_/a_255_603# 0.002146f
C2248 _293_/a_36_472# _105_ 0.004667f
C2249 _255_/a_224_552# _118_ 0.002405f
C2250 state\[1\] _062_ 0.001179f
C2251 FILLER_0_7_72/a_1916_375# _376_/a_36_160# 0.001925f
C2252 net44 FILLER_0_15_2/a_124_375# 0.017852f
C2253 FILLER_0_22_86/a_1020_375# vdd 0.008761f
C2254 net38 _450_/a_1293_527# 0.001307f
C2255 _114_ _056_ 0.034246f
C2256 FILLER_0_12_2/a_572_375# net44 0.041552f
C2257 _033_ FILLER_0_6_47/a_36_472# 0.001185f
C2258 ctlp[1] vss 0.32843f
C2259 _126_ net23 0.030487f
C2260 _140_ _348_/a_257_69# 0.001089f
C2261 FILLER_0_7_59/a_124_375# net67 0.036499f
C2262 _091_ vss 0.56693f
C2263 _020_ _334_/a_36_160# 0.028435f
C2264 net79 _100_ 0.170973f
C2265 _422_/a_1204_472# _009_ 0.009783f
C2266 _417_/a_2665_112# vdd 0.03015f
C2267 net73 fanout73/a_36_113# 0.02062f
C2268 FILLER_0_12_136/a_1380_472# vss 0.031524f
C2269 _449_/a_36_151# net15 0.020788f
C2270 _074_ FILLER_0_5_181/a_36_472# 0.002385f
C2271 FILLER_0_9_142/a_36_472# vdd 0.107619f
C2272 FILLER_0_9_142/a_124_375# vss 0.006851f
C2273 _050_ _208_/a_36_160# 0.001038f
C2274 _295_/a_244_68# _107_ 0.00123f
C2275 _077_ FILLER_0_9_223/a_36_472# 0.005511f
C2276 _092_ FILLER_0_18_209/a_484_472# 0.006303f
C2277 output31/a_224_472# _008_ 0.051074f
C2278 net53 vss 0.426484f
C2279 _411_/a_1000_472# net8 0.007241f
C2280 FILLER_0_13_206/a_36_472# _043_ 0.011439f
C2281 _105_ _422_/a_2665_112# 0.011125f
C2282 net20 _421_/a_1308_423# 0.012036f
C2283 net61 _421_/a_2665_112# 0.001339f
C2284 net78 _421_/a_1204_472# 0.006482f
C2285 net60 _421_/a_1204_472# 0.021679f
C2286 output8/a_224_472# _080_ 0.001971f
C2287 _045_ vdd 0.246567f
C2288 _437_/a_2248_156# vdd 0.054674f
C2289 _129_ _058_ 0.050726f
C2290 _373_/a_1060_68# _090_ 0.002234f
C2291 cal net1 0.336092f
C2292 _029_ FILLER_0_5_88/a_36_472# 0.007596f
C2293 net57 _428_/a_796_472# 0.003017f
C2294 net61 _422_/a_1308_423# 0.002171f
C2295 net60 _422_/a_36_151# 0.008119f
C2296 net78 _422_/a_36_151# 0.023285f
C2297 FILLER_0_4_213/a_484_472# vdd 0.007084f
C2298 FILLER_0_4_213/a_36_472# vss 0.003969f
C2299 _308_/a_848_380# FILLER_0_9_105/a_36_472# 0.15783f
C2300 _093_ net30 0.001859f
C2301 net53 net74 0.164124f
C2302 _390_/a_36_68# net14 0.010844f
C2303 _448_/a_36_151# FILLER_0_1_192/a_36_472# 0.008172f
C2304 _431_/a_2248_156# FILLER_0_15_142/a_484_472# 0.016128f
C2305 output16/a_224_472# ctln[9] 0.08624f
C2306 net47 FILLER_0_5_148/a_36_472# 0.004409f
C2307 _144_ _352_/a_257_69# 0.001662f
C2308 _192_/a_67_603# vdd 0.027014f
C2309 _028_ FILLER_0_7_104/a_124_375# 0.008248f
C2310 _069_ _122_ 0.002164f
C2311 FILLER_0_4_197/a_572_375# net21 0.041173f
C2312 _273_/a_36_68# _060_ 0.010339f
C2313 _301_/a_36_472# mask\[8\] 0.016751f
C2314 _074_ cal_itt\[1\] 0.120296f
C2315 output20/a_224_472# result[9] 0.001884f
C2316 net54 _433_/a_2665_112# 0.047439f
C2317 net57 net52 0.016136f
C2318 net61 fanout61/a_36_113# 0.023179f
C2319 _043_ FILLER_0_15_180/a_124_375# 0.003099f
C2320 _255_/a_224_552# _068_ 0.002412f
C2321 _057_ _070_ 0.033401f
C2322 FILLER_0_21_125/a_484_472# _433_/a_36_151# 0.001723f
C2323 FILLER_0_5_128/a_572_375# _133_ 0.00134f
C2324 FILLER_0_5_128/a_36_472# _070_ 0.036f
C2325 FILLER_0_11_78/a_124_375# vss 0.006233f
C2326 FILLER_0_11_78/a_572_375# vdd -0.006646f
C2327 _077_ net23 0.0245f
C2328 _432_/a_36_151# FILLER_0_17_161/a_124_375# 0.035117f
C2329 _020_ net36 0.001995f
C2330 trimb[4] net38 0.124219f
C2331 _412_/a_2665_112# net59 0.055415f
C2332 _162_ _312_/a_234_472# 0.003812f
C2333 net67 net42 0.101108f
C2334 fanout57/a_36_113# net82 0.017696f
C2335 _074_ FILLER_0_7_233/a_36_472# 0.001341f
C2336 net20 FILLER_0_8_239/a_124_375# 0.004302f
C2337 _444_/a_36_151# _054_ 0.011342f
C2338 net58 FILLER_0_9_290/a_124_375# 0.001157f
C2339 output16/a_224_472# vss 0.009875f
C2340 FILLER_0_13_206/a_36_472# net21 0.00171f
C2341 _050_ _210_/a_67_603# 0.006444f
C2342 ctlp[4] net33 0.001734f
C2343 _301_/a_36_472# vss 0.003975f
C2344 FILLER_0_12_50/a_36_472# vdd 0.012805f
C2345 FILLER_0_12_50/a_124_375# vss 0.004123f
C2346 _415_/a_36_151# net79 0.001156f
C2347 _321_/a_1602_69# _120_ 0.00262f
C2348 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_36_472# 0.086635f
C2349 trim_val\[4\] _443_/a_2665_112# 0.018733f
C2350 _325_/a_224_472# _120_ 0.00233f
C2351 _094_ _099_ 0.193065f
C2352 _423_/a_36_151# _012_ 0.021631f
C2353 _013_ _217_/a_36_160# 0.001614f
C2354 _028_ FILLER_0_5_72/a_932_472# 0.003042f
C2355 _430_/a_796_472# _019_ 0.006511f
C2356 cal_itt\[2\] _074_ 0.082824f
C2357 _422_/a_1308_423# _108_ 0.019345f
C2358 fanout66/a_36_113# _441_/a_36_151# 0.032681f
C2359 FILLER_0_9_60/a_484_472# vss 0.005321f
C2360 _077_ _439_/a_2248_156# 0.038814f
C2361 _069_ _061_ 0.024151f
C2362 net69 _369_/a_36_68# 0.008024f
C2363 _031_ _369_/a_244_472# 0.002741f
C2364 FILLER_0_4_152/a_124_375# trim_mask\[4\] 0.01182f
C2365 FILLER_0_10_214/a_36_472# _060_ 0.001378f
C2366 fanout72/a_36_113# vss 0.053396f
C2367 FILLER_0_7_72/a_3172_472# _219_/a_36_160# 0.035111f
C2368 FILLER_0_13_65/a_36_472# fanout72/a_36_113# 0.193651f
C2369 output42/a_224_472# trim[4] 0.017153f
C2370 FILLER_0_3_172/a_1828_472# net22 0.009883f
C2371 FILLER_0_4_144/a_124_375# net23 0.011315f
C2372 FILLER_0_10_256/a_124_375# vss 0.006036f
C2373 FILLER_0_10_256/a_36_472# vdd 0.025204f
C2374 _030_ _160_ 0.063581f
C2375 net66 _034_ 0.139638f
C2376 net49 _166_ 0.007445f
C2377 _074_ FILLER_0_6_177/a_36_472# 0.045576f
C2378 FILLER_0_23_282/a_572_375# vdd -0.013698f
C2379 FILLER_0_23_282/a_124_375# vss 0.005048f
C2380 _430_/a_2248_156# _092_ 0.003124f
C2381 net22 net37 0.03068f
C2382 output26/a_224_472# net17 0.004277f
C2383 _424_/a_1000_472# _012_ 0.00675f
C2384 FILLER_0_7_72/a_1020_375# vdd 0.004039f
C2385 FILLER_0_7_72/a_572_375# vss 0.006884f
C2386 fanout72/a_36_113# net74 0.02894f
C2387 _075_ _122_ 0.030339f
C2388 ctln[3] _411_/a_2248_156# 0.001208f
C2389 _445_/a_1308_423# _034_ 0.002494f
C2390 _137_ net23 0.031218f
C2391 net35 FILLER_0_22_177/a_1468_375# 0.048182f
C2392 FILLER_0_22_86/a_36_472# net71 0.005766f
C2393 net81 net37 0.18149f
C2394 FILLER_0_11_109/a_36_472# vss 0.003131f
C2395 _285_/a_36_472# mask\[1\] 0.036335f
C2396 FILLER_0_2_93/a_572_375# vss 0.055237f
C2397 _002_ FILLER_0_3_172/a_2364_375# 0.016984f
C2398 _052_ FILLER_0_21_28/a_1468_375# 0.001757f
C2399 FILLER_0_10_78/a_1020_375# _115_ 0.064761f
C2400 _311_/a_254_473# net21 0.003733f
C2401 net75 _073_ 0.34505f
C2402 FILLER_0_11_135/a_36_472# vss 0.006739f
C2403 FILLER_0_21_28/a_124_375# net17 0.005751f
C2404 _345_/a_36_160# _145_ 0.001141f
C2405 output35/a_224_472# _204_/a_67_603# 0.012678f
C2406 _437_/a_36_151# net14 0.014361f
C2407 FILLER_0_16_255/a_124_375# net19 0.008033f
C2408 _448_/a_1204_472# vdd 0.002228f
C2409 trim[0] _035_ 0.171633f
C2410 net15 FILLER_0_9_60/a_572_375# 0.047331f
C2411 _077_ _311_/a_1660_473# 0.001653f
C2412 FILLER_0_13_212/a_572_375# _043_ 0.01418f
C2413 net69 net23 0.064573f
C2414 _072_ _395_/a_1492_488# 0.003088f
C2415 _155_ _028_ 0.049284f
C2416 FILLER_0_14_235/a_484_472# net62 0.017862f
C2417 FILLER_0_14_107/a_484_472# vdd 0.030114f
C2418 FILLER_0_14_107/a_36_472# vss 0.003706f
C2419 _431_/a_2665_112# _137_ 0.010924f
C2420 sample vdd 0.154389f
C2421 FILLER_0_22_177/a_36_472# vss 0.002984f
C2422 FILLER_0_22_177/a_484_472# vdd 0.006974f
C2423 _115_ FILLER_0_9_72/a_932_472# 0.001837f
C2424 _449_/a_448_472# cal_count\[3\] 0.007511f
C2425 _053_ _372_/a_170_472# 0.05895f
C2426 _219_/a_36_160# _058_ 0.014194f
C2427 _053_ _131_ 0.086215f
C2428 net69 _441_/a_2665_112# 0.014995f
C2429 _111_ mask\[9\] 0.127919f
C2430 _120_ _171_ 0.414533f
C2431 _063_ _378_/a_224_472# 0.002323f
C2432 _439_/a_36_151# _453_/a_2248_156# 0.001082f
C2433 FILLER_0_5_109/a_484_472# vdd 0.007355f
C2434 cal_itt\[2\] FILLER_0_3_221/a_484_472# 0.016997f
C2435 _161_ vss 0.134214f
C2436 net71 _437_/a_2560_156# 0.037081f
C2437 fanout74/a_36_113# net69 0.006779f
C2438 net49 trim_mask\[1\] 0.003402f
C2439 _077_ _056_ 1.777574f
C2440 _447_/a_2665_112# trim_val\[3\] 0.002721f
C2441 net50 _444_/a_2665_112# 0.023342f
C2442 net38 _095_ 0.032393f
C2443 _429_/a_36_151# FILLER_0_15_212/a_124_375# 0.059049f
C2444 FILLER_0_0_130/a_36_472# net13 0.002757f
C2445 net34 FILLER_0_22_128/a_2812_375# 0.005158f
C2446 fanout73/a_36_113# _427_/a_36_151# 0.032681f
C2447 net65 trim_val\[4\] 0.015549f
C2448 _436_/a_2665_112# net54 0.042428f
C2449 _452_/a_36_151# vdd 0.109842f
C2450 net68 trim_mask\[1\] 0.054055f
C2451 result[8] _422_/a_448_472# 0.002989f
C2452 output9/a_224_472# net8 0.020421f
C2453 _016_ _428_/a_448_472# 0.00347f
C2454 _101_ _283_/a_36_472# 0.002471f
C2455 _008_ FILLER_0_17_226/a_36_472# 0.001842f
C2456 _137_ FILLER_0_15_180/a_484_472# 0.046411f
C2457 _041_ FILLER_0_18_37/a_1468_375# 0.001032f
C2458 FILLER_0_4_123/a_36_472# net47 0.012399f
C2459 _432_/a_36_151# _098_ 0.00957f
C2460 _308_/a_1084_68# _114_ 0.00178f
C2461 _308_/a_848_380# _115_ 0.00763f
C2462 net35 FILLER_0_23_88/a_124_375# 0.009071f
C2463 _407_/a_36_472# _185_ 0.009281f
C2464 net32 _102_ 0.038622f
C2465 FILLER_0_16_73/a_124_375# net55 0.007695f
C2466 FILLER_0_12_136/a_932_472# cal_count\[3\] 0.007247f
C2467 _077_ _392_/a_36_68# 0.055912f
C2468 FILLER_0_18_177/a_3260_375# vss 0.055219f
C2469 FILLER_0_18_177/a_36_472# vdd 0.110153f
C2470 _176_ _120_ 0.169846f
C2471 _428_/a_1000_472# _131_ 0.035998f
C2472 net9 vdd 0.190349f
C2473 _093_ FILLER_0_18_107/a_484_472# 0.008683f
C2474 _091_ _097_ 0.036863f
C2475 _255_/a_224_552# vdd 0.082462f
C2476 output24/a_224_472# vdd 0.08781f
C2477 _418_/a_2665_112# vdd 0.028061f
C2478 _411_/a_2665_112# net58 0.018133f
C2479 _076_ FILLER_0_8_156/a_484_472# 0.008487f
C2480 _105_ _011_ 0.003998f
C2481 FILLER_0_9_60/a_572_375# net51 0.002279f
C2482 _017_ cal_count\[3\] 0.003939f
C2483 _076_ net37 0.072179f
C2484 _450_/a_2225_156# net40 0.04513f
C2485 _143_ _093_ 0.003295f
C2486 FILLER_0_18_100/a_36_472# mask\[9\] 0.005719f
C2487 FILLER_0_23_88/a_36_472# vss 0.003481f
C2488 FILLER_0_5_206/a_36_472# _081_ 0.014328f
C2489 net75 _425_/a_36_151# 0.02868f
C2490 _149_ _437_/a_2665_112# 0.020763f
C2491 _026_ _437_/a_1204_472# 0.022954f
C2492 net41 _446_/a_1000_472# 0.01097f
C2493 _095_ _451_/a_2449_156# 0.001843f
C2494 FILLER_0_16_57/a_124_375# vdd 0.008567f
C2495 _440_/a_36_151# FILLER_0_6_47/a_1828_472# 0.001512f
C2496 trimb[4] net55 0.01379f
C2497 _086_ _250_/a_36_68# 0.001132f
C2498 FILLER_0_12_28/a_124_375# vdd 0.040988f
C2499 _287_/a_36_472# vdd 0.072871f
C2500 _432_/a_36_151# net63 0.001392f
C2501 net56 net23 0.930833f
C2502 FILLER_0_13_142/a_932_472# net23 0.020589f
C2503 net47 _153_ 0.755476f
C2504 _250_/a_36_68# cal_count\[3\] 0.004136f
C2505 _441_/a_448_472# _168_ 0.033059f
C2506 _092_ net22 0.010937f
C2507 _093_ _136_ 0.226819f
C2508 FILLER_0_13_212/a_1380_472# net62 0.059367f
C2509 net20 mask\[2\] 0.050364f
C2510 net75 net1 0.098901f
C2511 net41 _408_/a_1336_472# 0.063099f
C2512 FILLER_0_1_204/a_124_375# net11 0.01048f
C2513 FILLER_0_5_72/a_1020_375# _164_ 0.018398f
C2514 _327_/a_244_68# _130_ 0.00117f
C2515 fanout71/a_36_113# _149_ 0.001315f
C2516 _431_/a_2665_112# net56 0.048214f
C2517 FILLER_0_3_204/a_36_472# net22 0.036788f
C2518 _098_ FILLER_0_19_171/a_572_375# 0.001946f
C2519 net15 _453_/a_2560_156# 0.049334f
C2520 _095_ FILLER_0_13_72/a_484_472# 0.027852f
C2521 _098_ FILLER_0_15_235/a_572_375# 0.001343f
C2522 net20 result[7] 0.134149f
C2523 _127_ vss 0.343764f
C2524 output44/a_224_472# FILLER_0_20_15/a_932_472# 0.0323f
C2525 _432_/a_36_151# FILLER_0_18_171/a_36_472# 0.059367f
C2526 FILLER_0_12_50/a_36_472# cal_count\[0\] 0.001857f
C2527 net16 _013_ 0.060401f
C2528 _413_/a_2665_112# output11/a_224_472# 0.001492f
C2529 _074_ net59 0.030221f
C2530 output34/a_224_472# _099_ 0.001498f
C2531 net76 FILLER_0_5_212/a_124_375# 0.004635f
C2532 _093_ _356_/a_36_472# 0.009235f
C2533 _363_/a_244_472# vdd 0.002075f
C2534 vss FILLER_0_16_115/a_36_472# 0.003243f
C2535 _074_ net4 0.088616f
C2536 FILLER_0_6_47/a_1828_472# vdd 0.002735f
C2537 FILLER_0_6_47/a_1380_472# vss 0.001431f
C2538 _085_ _121_ 0.027373f
C2539 output20/a_224_472# net61 0.177946f
C2540 _429_/a_796_472# net22 0.020124f
C2541 FILLER_0_12_124/a_36_472# cal_count\[3\] 0.004109f
C2542 _093_ FILLER_0_17_72/a_2364_375# 0.010888f
C2543 _402_/a_1948_68# vdd 0.001429f
C2544 FILLER_0_5_117/a_36_472# net47 0.005919f
C2545 _127_ net74 0.0588f
C2546 vdd _039_ 0.219985f
C2547 _228_/a_36_68# _113_ 0.021898f
C2548 output13/a_224_472# _170_ 0.024999f
C2549 output42/a_224_472# _236_/a_36_160# 0.001892f
C2550 net81 _429_/a_796_472# 0.002847f
C2551 net70 _040_ 0.018254f
C2552 _156_ _160_ 0.299745f
C2553 FILLER_0_4_197/a_932_472# net22 0.0473f
C2554 fanout67/a_36_160# FILLER_0_9_60/a_124_375# 0.02985f
C2555 _098_ FILLER_0_20_98/a_36_472# 0.0127f
C2556 _418_/a_448_472# _007_ 0.050316f
C2557 net82 FILLER_0_3_221/a_124_375# 0.015932f
C2558 _255_/a_224_552# _057_ 0.024333f
C2559 _077_ FILLER_0_10_78/a_932_472# 0.002503f
C2560 _132_ FILLER_0_15_116/a_124_375# 0.047331f
C2561 FILLER_0_21_125/a_124_375# net54 0.008377f
C2562 _086_ FILLER_0_11_135/a_124_375# 0.008238f
C2563 _422_/a_2248_156# mask\[7\] 0.015008f
C2564 _449_/a_36_151# _394_/a_728_93# 0.002727f
C2565 net52 _443_/a_2560_156# 0.020855f
C2566 _426_/a_36_151# _425_/a_36_151# 0.006252f
C2567 net67 _160_ 0.003659f
C2568 _071_ vss 0.126519f
C2569 net65 FILLER_0_9_282/a_572_375# 0.001388f
C2570 en_co_clk _038_ 0.014475f
C2571 _426_/a_2248_156# calibrate 0.004597f
C2572 cal_count\[3\] FILLER_0_11_109/a_124_375# 0.004618f
C2573 _430_/a_36_151# FILLER_0_17_200/a_124_375# 0.059049f
C2574 net17 output6/a_224_472# 0.047757f
C2575 ctlp[9] vdd 0.17413f
C2576 FILLER_0_14_91/a_572_375# net14 0.005527f
C2577 _446_/a_2665_112# _034_ 0.002484f
C2578 _273_/a_36_68# vss 0.095582f
C2579 _136_ FILLER_0_17_142/a_124_375# 0.001315f
C2580 clk net18 0.003519f
C2581 output46/a_224_472# FILLER_0_20_2/a_124_375# 0.030009f
C2582 net55 _095_ 0.055644f
C2583 cal_count\[3\] FILLER_0_11_135/a_124_375# 0.004365f
C2584 _174_ FILLER_0_15_59/a_572_375# 0.007123f
C2585 net2 net9 0.001033f
C2586 _453_/a_2560_156# net51 0.013556f
C2587 net57 FILLER_0_13_142/a_1020_375# 0.009442f
C2588 _402_/a_2172_497# _180_ 0.001094f
C2589 FILLER_0_7_162/a_36_472# _074_ 0.003809f
C2590 _415_/a_2665_112# result[1] 0.010555f
C2591 _428_/a_448_472# _043_ 0.063478f
C2592 _140_ net71 0.005182f
C2593 net38 vss 0.633752f
C2594 FILLER_0_16_89/a_1380_472# _131_ 0.004201f
C2595 _086_ _162_ 0.107276f
C2596 _433_/a_1288_156# _022_ 0.001147f
C2597 output20/a_224_472# _108_ 0.022243f
C2598 mask\[3\] _282_/a_36_160# 0.005823f
C2599 _143_ FILLER_0_17_161/a_36_472# 0.00363f
C2600 _430_/a_1204_472# net63 0.013728f
C2601 FILLER_0_4_107/a_1380_472# net47 0.008874f
C2602 _030_ _156_ 0.153053f
C2603 FILLER_0_3_221/a_484_472# net59 0.001655f
C2604 FILLER_0_12_20/a_36_472# net47 0.020589f
C2605 FILLER_0_4_197/a_36_472# _079_ 0.002448f
C2606 FILLER_0_4_197/a_1468_375# _088_ 0.012367f
C2607 _052_ _424_/a_1308_423# 0.008633f
C2608 FILLER_0_21_28/a_2364_375# vdd -0.011393f
C2609 _403_/a_224_472# _183_ 0.007508f
C2610 ctln[5] net76 0.001707f
C2611 FILLER_0_3_172/a_1380_472# vdd 0.043045f
C2612 _442_/a_36_151# FILLER_0_2_127/a_36_472# 0.012873f
C2613 _449_/a_2665_112# net55 0.057694f
C2614 _053_ _077_ 0.123663f
C2615 net4 FILLER_0_3_221/a_484_472# 0.043027f
C2616 vss FILLER_0_8_156/a_572_375# 0.007969f
C2617 vdd FILLER_0_8_156/a_36_472# 0.002891f
C2618 _438_/a_2665_112# net14 0.026903f
C2619 _091_ _019_ 0.031681f
C2620 result[6] _421_/a_36_151# 0.032036f
C2621 _413_/a_2560_156# net82 0.00101f
C2622 _122_ net22 0.024638f
C2623 net55 FILLER_0_17_72/a_484_472# 0.019636f
C2624 net81 FILLER_0_14_235/a_36_472# 0.002571f
C2625 _447_/a_36_151# net17 0.001448f
C2626 _081_ _123_ 0.007811f
C2627 FILLER_0_18_2/a_2364_375# net17 0.048345f
C2628 _144_ _433_/a_796_472# 0.008448f
C2629 FILLER_0_4_152/a_124_375# _066_ 0.003354f
C2630 ctln[7] FILLER_0_0_96/a_124_375# 0.025944f
C2631 FILLER_0_16_37/a_124_375# net72 0.013591f
C2632 net52 _037_ 0.103749f
C2633 FILLER_0_5_109/a_572_375# _154_ 0.014669f
C2634 FILLER_0_20_87/a_36_472# _437_/a_36_151# 0.001723f
C2635 FILLER_0_5_72/a_1380_472# net49 0.002057f
C2636 FILLER_0_10_214/a_36_472# vss 0.008006f
C2637 _005_ _416_/a_2665_112# 0.014205f
C2638 _036_ _446_/a_2248_156# 0.001763f
C2639 _443_/a_1204_472# _170_ 0.002808f
C2640 _056_ _060_ 0.085489f
C2641 _061_ _090_ 0.00832f
C2642 _132_ FILLER_0_17_104/a_484_472# 0.002737f
C2643 net1 _265_/a_916_472# 0.002088f
C2644 net48 _316_/a_848_380# 0.026413f
C2645 _131_ FILLER_0_17_104/a_1468_375# 0.006022f
C2646 net16 _179_ 0.007397f
C2647 trim_val\[4\] FILLER_0_3_172/a_124_375# 0.002076f
C2648 _095_ net23 0.053365f
C2649 output8/a_224_472# net75 0.044765f
C2650 _395_/a_244_68# _070_ 0.001481f
C2651 FILLER_0_9_72/a_36_472# _453_/a_2248_156# 0.013656f
C2652 _084_ vdd 0.134578f
C2653 result[2] net18 0.086474f
C2654 net22 _435_/a_2665_112# 0.004214f
C2655 FILLER_0_5_109/a_124_375# _163_ 0.002658f
C2656 _061_ net22 0.123662f
C2657 net68 _054_ 0.08092f
C2658 _431_/a_1204_472# net73 0.026905f
C2659 mask\[3\] FILLER_0_18_177/a_1916_375# 0.003052f
C2660 FILLER_0_12_28/a_124_375# cal_count\[0\] 0.001414f
C2661 net53 FILLER_0_17_142/a_572_375# 0.023771f
C2662 net21 _202_/a_36_160# 0.09166f
C2663 FILLER_0_4_107/a_124_375# vdd 0.036972f
C2664 _103_ _418_/a_2248_156# 0.012186f
C2665 _091_ _429_/a_2248_156# 0.006148f
C2666 FILLER_0_5_212/a_36_472# _078_ 0.002235f
C2667 _374_/a_36_68# _062_ 0.004248f
C2668 net60 _418_/a_2665_112# 0.042307f
C2669 net28 _045_ 0.05144f
C2670 fanout77/a_36_113# _094_ 0.002244f
C2671 _149_ net71 0.827628f
C2672 net31 ctlp[1] 0.050993f
C2673 vss FILLER_0_13_72/a_484_472# 0.008682f
C2674 _436_/a_36_151# _437_/a_2248_156# 0.001837f
C2675 mask\[5\] _434_/a_2248_156# 0.003462f
C2676 trimb[1] net44 0.089379f
C2677 _387_/a_36_113# _037_ 0.003577f
C2678 net31 _091_ 0.001465f
C2679 net65 net18 0.879399f
C2680 net68 FILLER_0_8_37/a_124_375# 0.004818f
C2681 FILLER_0_8_127/a_36_472# _062_ 0.01783f
C2682 net47 _166_ 0.034342f
C2683 _010_ net77 0.009534f
C2684 _432_/a_2248_156# _091_ 0.007123f
C2685 mask\[0\] net79 0.243338f
C2686 FILLER_0_7_162/a_124_375# _062_ 0.010242f
C2687 _132_ FILLER_0_19_125/a_124_375# 0.009167f
C2688 trim_mask\[4\] _158_ 0.022724f
C2689 _233_/a_36_160# vss 0.01649f
C2690 net28 _192_/a_67_603# 0.119061f
C2691 _079_ FILLER_0_6_231/a_572_375# 0.002768f
C2692 _199_/a_36_160# vss 0.004608f
C2693 net74 FILLER_0_13_72/a_484_472# 0.007142f
C2694 _246_/a_36_68# vss 0.024639f
C2695 _114_ _072_ 0.078148f
C2696 _401_/a_244_472# _180_ 0.001689f
C2697 result[8] result[9] 0.242998f
C2698 _242_/a_36_160# FILLER_0_5_164/a_36_472# 0.193804f
C2699 _028_ FILLER_0_6_47/a_2364_375# 0.016593f
C2700 _127_ FILLER_0_11_142/a_484_472# 0.001177f
C2701 _095_ FILLER_0_15_10/a_36_472# 0.00335f
C2702 net54 _354_/a_49_472# 0.002169f
C2703 _068_ calibrate 0.110297f
C2704 _076_ _122_ 0.097035f
C2705 _002_ net76 0.213703f
C2706 net65 _412_/a_1308_423# 0.024499f
C2707 FILLER_0_7_104/a_484_472# FILLER_0_9_105/a_572_375# 0.001188f
C2708 _449_/a_36_151# _067_ 0.031377f
C2709 _189_/a_67_603# net64 0.064691f
C2710 result[8] FILLER_0_23_282/a_36_472# 0.001908f
C2711 net15 FILLER_0_13_72/a_572_375# 0.003021f
C2712 net57 _136_ 0.168299f
C2713 _033_ _444_/a_1308_423# 0.002877f
C2714 net32 output19/a_224_472# 0.101682f
C2715 _053_ FILLER_0_6_47/a_572_375# 0.008213f
C2716 mask\[4\] FILLER_0_20_193/a_484_472# 0.001215f
C2717 _394_/a_1936_472# _175_ 0.017848f
C2718 _068_ _311_/a_1920_473# 0.001498f
C2719 _427_/a_2560_156# _095_ 0.009888f
C2720 _039_ cal_count\[0\] 0.219667f
C2721 _417_/a_36_151# output30/a_224_472# 0.004902f
C2722 _370_/a_124_24# _081_ 0.015048f
C2723 FILLER_0_14_81/a_124_375# net55 0.038949f
C2724 _125_ _118_ 0.239695f
C2725 output38/a_224_472# output41/a_224_472# 0.00607f
C2726 _235_/a_67_603# _447_/a_36_151# 0.038675f
C2727 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3260_375# 0.086905f
C2728 FILLER_0_0_198/a_124_375# vdd 0.04491f
C2729 _305_/a_36_159# _081_ 0.039192f
C2730 cal_count\[3\] _373_/a_244_68# 0.002341f
C2731 net55 vss 0.947665f
C2732 FILLER_0_9_223/a_36_472# vss 0.019592f
C2733 FILLER_0_9_223/a_484_472# vdd 0.004285f
C2734 trim_mask\[1\] net47 0.306848f
C2735 _451_/a_1040_527# net14 0.029964f
C2736 FILLER_0_3_204/a_124_375# vdd 0.023302f
C2737 mask\[4\] FILLER_0_18_139/a_1380_472# 0.003851f
C2738 sample FILLER_0_9_290/a_124_375# 0.00195f
C2739 net20 FILLER_0_15_212/a_1380_472# 0.001449f
C2740 _369_/a_36_68# vss 0.002343f
C2741 fanout57/a_36_113# net65 0.035361f
C2742 output28/a_224_472# vdd 0.044767f
C2743 net17 _452_/a_1697_156# 0.001184f
C2744 _061_ _076_ 0.024289f
C2745 net18 _419_/a_448_472# 0.037373f
C2746 net57 _070_ 0.202843f
C2747 FILLER_0_10_256/a_36_472# net28 0.00136f
C2748 _443_/a_1000_472# net69 0.008276f
C2749 net32 mask\[5\] 0.304094f
C2750 FILLER_0_12_2/a_124_375# clkc 0.003601f
C2751 FILLER_0_5_172/a_124_375# net37 0.014083f
C2752 result[2] net62 0.311075f
C2753 net82 trim_mask\[4\] 0.21475f
C2754 net55 net74 0.048927f
C2755 FILLER_0_14_99/a_124_375# FILLER_0_13_100/a_36_472# 0.001597f
C2756 vss _416_/a_1308_423# 0.001962f
C2757 _176_ _043_ 0.04106f
C2758 output27/a_224_472# FILLER_0_9_282/a_484_472# 0.001711f
C2759 net27 FILLER_0_9_282/a_124_375# 0.003572f
C2760 _069_ _267_/a_36_472# 0.003607f
C2761 _429_/a_448_472# vss 0.035246f
C2762 net64 FILLER_0_14_235/a_124_375# 0.046554f
C2763 _119_ FILLER_0_8_156/a_572_375# 0.01739f
C2764 _114_ FILLER_0_13_142/a_1468_375# 0.001931f
C2765 _423_/a_36_151# vdd 0.088377f
C2766 vdd clkc 0.190259f
C2767 _306_/a_36_68# _043_ 0.001086f
C2768 _088_ FILLER_0_5_198/a_572_375# 0.001374f
C2769 _079_ FILLER_0_5_198/a_36_472# 0.012251f
C2770 _335_/a_49_472# _043_ 0.00367f
C2771 _395_/a_36_488# vdd 0.066813f
C2772 result[4] FILLER_0_15_290/a_36_472# 0.001422f
C2773 state\[1\] FILLER_0_12_196/a_36_472# 0.030132f
C2774 _189_/a_67_603# vss 0.004088f
C2775 net55 cal_count\[1\] 0.204733f
C2776 _292_/a_36_160# _204_/a_67_603# 0.003478f
C2777 FILLER_0_4_197/a_484_472# vdd 0.002749f
C2778 ctln[1] ctln[2] 0.047127f
C2779 _053_ _165_ 0.123461f
C2780 FILLER_0_8_107/a_36_472# _058_ 0.015262f
C2781 _432_/a_1308_423# vdd 0.029938f
C2782 mask\[1\] FILLER_0_15_180/a_484_472# 0.003594f
C2783 _008_ _419_/a_36_151# 0.014476f
C2784 net23 vss 1.922425f
C2785 FILLER_0_20_107/a_124_375# vdd 0.04384f
C2786 _343_/a_49_472# _143_ 0.00918f
C2787 FILLER_0_7_146/a_124_375# _062_ 0.028312f
C2788 vss trim[2] 0.026644f
C2789 _238_/a_67_603# trim_mask\[2\] 0.003021f
C2790 result[8] _048_ 0.006006f
C2791 FILLER_0_23_290/a_36_472# vdd 0.089567f
C2792 FILLER_0_23_290/a_124_375# vss 0.033011f
C2793 _424_/a_1000_472# vdd 0.002952f
C2794 _176_ _175_ 0.054439f
C2795 _150_ _438_/a_36_151# 0.032532f
C2796 _441_/a_2665_112# vss 0.005169f
C2797 _444_/a_448_472# net17 0.022222f
C2798 _072_ _126_ 0.012566f
C2799 FILLER_0_22_128/a_2812_375# _146_ 0.001336f
C2800 _064_ vdd 0.874293f
C2801 _059_ _160_ 0.037235f
C2802 net55 _452_/a_836_156# 0.010887f
C2803 net69 _164_ 0.040362f
C2804 _015_ _426_/a_2665_112# 0.018623f
C2805 _228_/a_36_68# vdd 0.036391f
C2806 _447_/a_1204_472# vdd 0.001085f
C2807 FILLER_0_18_2/a_932_472# vdd 0.002342f
C2808 FILLER_0_18_2/a_484_472# vss 0.001228f
C2809 net74 net23 0.0064f
C2810 _114_ FILLER_0_11_101/a_36_472# 0.00501f
C2811 fanout74/a_36_113# vss 0.048756f
C2812 net39 trim[1] 0.115976f
C2813 _005_ _100_ 0.004305f
C2814 result[4] FILLER_0_17_282/a_36_472# 0.017375f
C2815 _431_/a_2665_112# vss 0.033886f
C2816 _148_ _352_/a_257_69# 0.001417f
C2817 _446_/a_1308_423# _035_ 0.002639f
C2818 FILLER_0_9_28/a_124_375# net40 0.047331f
C2819 _439_/a_2248_156# vss 0.003954f
C2820 _439_/a_2665_112# vdd 0.015979f
C2821 _127_ _321_/a_2034_472# 0.003159f
C2822 FILLER_0_20_193/a_572_375# _434_/a_2665_112# 0.002362f
C2823 _372_/a_2034_472# _152_ 0.00171f
C2824 _129_ _152_ 0.041257f
C2825 _412_/a_2248_156# net58 0.010702f
C2826 _091_ net80 0.23053f
C2827 FILLER_0_14_181/a_124_375# _043_ 0.008393f
C2828 mask\[8\] _025_ 0.036686f
C2829 _411_/a_796_472# vss 0.00159f
C2830 _176_ FILLER_0_10_107/a_484_472# 0.009571f
C2831 _386_/a_848_380# _169_ 0.001355f
C2832 _386_/a_124_24# _163_ 0.001234f
C2833 _098_ _437_/a_2665_112# 0.003567f
C2834 vdd FILLER_0_14_235/a_572_375# 0.006167f
C2835 vss FILLER_0_14_235/a_124_375# 0.002686f
C2836 fanout74/a_36_113# net74 0.007425f
C2837 FILLER_0_24_96/a_36_472# output25/a_224_472# 0.010475f
C2838 FILLER_0_21_125/a_36_472# _022_ 0.002295f
C2839 _432_/a_36_151# _137_ 0.051293f
C2840 result[6] net34 0.072393f
C2841 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_124_375# 0.001597f
C2842 net41 _450_/a_3129_107# 0.059083f
C2843 result[1] net19 0.084617f
C2844 net63 _434_/a_3041_156# 0.001449f
C2845 FILLER_0_15_180/a_484_472# vss 0.001207f
C2846 calibrate vdd 0.857987f
C2847 _132_ FILLER_0_18_107/a_1828_472# 0.045833f
C2848 net15 _441_/a_1204_472# 0.005939f
C2849 trim_mask\[2\] net15 0.026132f
C2850 _155_ FILLER_0_7_104/a_36_472# 0.005042f
C2851 FILLER_0_11_64/a_124_375# net15 0.047331f
C2852 _436_/a_36_151# output24/a_224_472# 0.053592f
C2853 fanout51/a_36_113# FILLER_0_11_64/a_124_375# 0.002335f
C2854 _025_ vss 0.016676f
C2855 _164_ FILLER_0_6_47/a_572_375# 0.010099f
C2856 _144_ net54 0.095482f
C2857 net67 FILLER_0_8_24/a_484_472# 0.001065f
C2858 FILLER_0_17_72/a_2724_472# net14 0.007133f
C2859 _086_ FILLER_0_6_177/a_484_472# 0.017841f
C2860 result[8] FILLER_0_24_290/a_124_375# 0.00562f
C2861 FILLER_0_15_10/a_36_472# vss 0.002605f
C2862 fanout71/a_36_113# _098_ 0.012725f
C2863 _132_ FILLER_0_16_107/a_124_375# 0.003315f
C2864 net20 FILLER_0_7_233/a_36_472# 0.035074f
C2865 net15 _439_/a_1000_472# 0.001798f
C2866 cal_itt\[3\] _074_ 0.584958f
C2867 _311_/a_1920_473# vdd 0.007492f
C2868 _077_ _072_ 0.178678f
C2869 FILLER_0_2_101/a_124_375# _367_/a_36_68# 0.001176f
C2870 FILLER_0_9_28/a_932_472# net16 0.017841f
C2871 net33 vss 0.674927f
C2872 mask\[5\] FILLER_0_18_177/a_1916_375# 0.002014f
C2873 fanout80/a_36_113# mask\[1\] 0.020046f
C2874 _053_ _079_ 0.007118f
C2875 _114_ FILLER_0_10_94/a_484_472# 0.011954f
C2876 _137_ FILLER_0_17_104/a_1468_375# 0.002679f
C2877 mask\[2\] FILLER_0_16_154/a_572_375# 0.026605f
C2878 FILLER_0_13_142/a_124_375# _043_ 0.009328f
C2879 FILLER_0_18_2/a_1828_472# _452_/a_448_472# 0.005748f
C2880 net36 FILLER_0_15_212/a_484_472# 0.007742f
C2881 _430_/a_1308_423# net21 0.008506f
C2882 _435_/a_2248_156# vdd 0.00571f
C2883 net20 cal_itt\[2\] 0.715447f
C2884 _053_ FILLER_0_6_79/a_124_375# 0.003818f
C2885 _081_ _242_/a_36_160# 0.025059f
C2886 vss FILLER_0_6_231/a_572_375# 0.057794f
C2887 vdd FILLER_0_6_231/a_36_472# 0.014642f
C2888 net20 _298_/a_224_472# 0.001861f
C2889 net17 FILLER_0_20_15/a_124_375# 0.005919f
C2890 _427_/a_2560_156# vss 0.003576f
C2891 _056_ vss 0.193804f
C2892 _414_/a_448_472# _089_ 0.003905f
C2893 _414_/a_36_151# _003_ 0.021191f
C2894 _434_/a_36_151# _348_/a_49_472# 0.017459f
C2895 FILLER_0_4_177/a_36_472# net22 0.006506f
C2896 FILLER_0_21_133/a_124_375# FILLER_0_21_125/a_572_375# 0.012001f
C2897 trim_val\[1\] _160_ 0.024279f
C2898 FILLER_0_9_28/a_36_472# vss -0.001119f
C2899 FILLER_0_9_28/a_484_472# vdd 0.010868f
C2900 FILLER_0_11_109/a_124_375# _120_ 0.016902f
C2901 _141_ FILLER_0_21_150/a_124_375# 0.02192f
C2902 cal_count\[2\] _184_ 0.033241f
C2903 _018_ _138_ 0.008093f
C2904 FILLER_0_14_263/a_36_472# output30/a_224_472# 0.002002f
C2905 FILLER_0_11_135/a_124_375# _120_ 0.017316f
C2906 _057_ _228_/a_36_68# 0.002062f
C2907 net51 net40 0.060626f
C2908 _443_/a_2248_156# net22 0.001984f
C2909 FILLER_0_10_37/a_36_472# FILLER_0_8_37/a_124_375# 0.001512f
C2910 _053_ FILLER_0_8_107/a_124_375# 0.002386f
C2911 FILLER_0_17_56/a_124_375# vdd 0.008529f
C2912 trim_val\[4\] vss 0.192567f
C2913 FILLER_0_11_64/a_124_375# net51 0.027848f
C2914 net52 FILLER_0_2_111/a_1020_375# 0.00245f
C2915 _126_ FILLER_0_11_101/a_36_472# 0.062336f
C2916 _372_/a_170_472# _133_ 0.031518f
C2917 _069_ _113_ 0.027402f
C2918 _131_ _133_ 0.20118f
C2919 _129_ _070_ 0.056776f
C2920 FILLER_0_8_138/a_36_472# _076_ 0.016628f
C2921 _392_/a_36_68# vss 0.002019f
C2922 fanout62/a_36_160# FILLER_0_11_282/a_36_472# 0.005262f
C2923 net72 _182_ 0.044895f
C2924 FILLER_0_8_37/a_36_472# _054_ 0.015053f
C2925 net16 _041_ 0.029736f
C2926 ctlp[3] _422_/a_36_151# 0.002627f
C2927 result[2] FILLER_0_15_282/a_572_375# 0.0011f
C2928 _165_ _164_ 0.351097f
C2929 result[8] net61 0.001106f
C2930 _072_ _267_/a_224_472# 0.004269f
C2931 FILLER_0_13_212/a_36_472# vss 0.005259f
C2932 ctln[8] net50 0.0032f
C2933 FILLER_0_6_177/a_36_472# _163_ 0.025039f
C2934 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_36_472# 0.026657f
C2935 fanout80/a_36_113# vss 0.003526f
C2936 result[5] _094_ 0.065897f
C2937 FILLER_0_17_72/a_2812_375# _131_ 0.006589f
C2938 net16 _181_ 0.48682f
C2939 net42 output6/a_224_472# 0.009273f
C2940 _292_/a_36_160# _201_/a_67_603# 0.003917f
C2941 FILLER_0_1_98/a_36_472# FILLER_0_0_96/a_124_375# 0.001684f
C2942 FILLER_0_5_72/a_1380_472# net47 0.003924f
C2943 FILLER_0_4_177/a_572_375# _087_ 0.006527f
C2944 FILLER_0_4_99/a_36_472# _153_ 0.066147f
C2945 FILLER_0_17_226/a_124_375# vdd 0.026497f
C2946 _057_ calibrate 0.002047f
C2947 mask\[4\] net34 0.001774f
C2948 FILLER_0_21_28/a_124_375# FILLER_0_19_28/a_36_472# 0.001512f
C2949 _125_ vdd 0.218505f
C2950 net15 FILLER_0_21_60/a_484_472# 0.001552f
C2951 _021_ vdd 0.022473f
C2952 fanout57/a_36_113# FILLER_0_3_172/a_124_375# 0.006548f
C2953 net52 FILLER_0_6_79/a_36_472# 0.012286f
C2954 net66 FILLER_0_3_54/a_124_375# 0.038548f
C2955 net50 fanout49/a_36_160# 0.059373f
C2956 _428_/a_1000_472# _095_ 0.001101f
C2957 FILLER_0_5_72/a_124_375# _440_/a_36_151# 0.059049f
C2958 _105_ output19/a_224_472# 0.107668f
C2959 _274_/a_2960_68# _070_ 0.001963f
C2960 result[7] FILLER_0_24_274/a_1020_375# 0.006125f
C2961 FILLER_0_7_72/a_3260_375# _058_ 0.00258f
C2962 _119_ net23 0.0245f
C2963 FILLER_0_21_150/a_124_375# _433_/a_2665_112# 0.029834f
C2964 mask\[7\] FILLER_0_22_128/a_1916_375# 0.007718f
C2965 _069_ _118_ 0.010986f
C2966 trimb[3] vss 0.161605f
C2967 _140_ _049_ 0.003069f
C2968 _052_ _216_/a_67_603# 0.006658f
C2969 FILLER_0_16_241/a_124_375# vss 0.04897f
C2970 FILLER_0_16_241/a_36_472# vdd 0.012388f
C2971 FILLER_0_15_150/a_124_375# net53 0.041074f
C2972 net2 calibrate 0.003482f
C2973 net47 _054_ 0.171966f
C2974 net39 _444_/a_448_472# 0.002089f
C2975 _168_ _160_ 0.03261f
C2976 _422_/a_2665_112# _107_ 0.005055f
C2977 FILLER_0_5_212/a_124_375# FILLER_0_3_212/a_36_472# 0.001512f
C2978 net41 _052_ 0.001927f
C2979 _412_/a_1000_472# net81 0.012828f
C2980 net16 _444_/a_2665_112# 0.011295f
C2981 cal_count\[2\] net47 0.274891f
C2982 net40 _381_/a_36_472# 0.020876f
C2983 FILLER_0_11_142/a_484_472# net23 0.006988f
C2984 net35 FILLER_0_22_128/a_1380_472# 0.016004f
C2985 net80 FILLER_0_22_177/a_36_472# 0.018848f
C2986 FILLER_0_14_91/a_484_472# FILLER_0_14_99/a_36_472# 0.013276f
C2987 net36 _451_/a_836_156# 0.007104f
C2988 FILLER_0_2_111/a_124_375# trim_mask\[3\] 0.004993f
C2989 trim_mask\[2\] _381_/a_36_472# 0.034251f
C2990 FILLER_0_8_24/a_36_472# net47 0.097212f
C2991 result[8] _108_ 0.007884f
C2992 output9/a_224_472# vdd 0.102412f
C2993 _105_ mask\[5\] 0.706158f
C2994 _013_ _424_/a_2248_156# 0.001828f
C2995 FILLER_0_9_72/a_932_472# _439_/a_36_151# 0.001723f
C2996 net64 FILLER_0_9_282/a_572_375# 0.002322f
C2997 _028_ _439_/a_36_151# 0.009268f
C2998 FILLER_0_11_64/a_36_472# cal_count\[3\] 0.0081f
C2999 ctlp[2] _422_/a_2248_156# 0.001328f
C3000 trim_mask\[1\] FILLER_0_6_47/a_36_472# 0.004319f
C3001 _098_ _048_ 0.092201f
C3002 _174_ vdd 0.18623f
C3003 _274_/a_3368_68# _091_ 0.001328f
C3004 _114_ state\[2\] 0.528838f
C3005 result[6] _419_/a_2665_112# 0.001225f
C3006 _207_/a_67_603# FILLER_0_22_128/a_3260_375# 0.00744f
C3007 net63 FILLER_0_22_177/a_932_472# 0.060639f
C3008 fanout53/a_36_160# _137_ 0.001852f
C3009 _248_/a_36_68# net62 0.002178f
C3010 _122_ FILLER_0_5_172/a_124_375# 0.001352f
C3011 FILLER_0_22_128/a_1828_472# vss 0.009137f
C3012 FILLER_0_22_128/a_2276_472# vdd 0.00565f
C3013 FILLER_0_16_89/a_36_472# _451_/a_448_472# 0.011974f
C3014 _052_ FILLER_0_18_37/a_572_375# 0.00706f
C3015 _444_/a_2248_156# vdd 0.041347f
C3016 _341_/a_665_69# net23 0.001508f
C3017 FILLER_0_16_73/a_484_472# _176_ 0.010681f
C3018 _128_ _122_ 0.019207f
C3019 _086_ _055_ 0.113385f
C3020 _446_/a_448_472# vdd 0.006805f
C3021 _030_ _168_ 0.015729f
C3022 FILLER_0_21_142/a_572_375# _433_/a_2665_112# 0.001092f
C3023 FILLER_0_21_142/a_124_375# _433_/a_2560_156# 0.001178f
C3024 FILLER_0_20_193/a_36_472# FILLER_0_18_177/a_1916_375# 0.0027f
C3025 FILLER_0_6_79/a_124_375# _164_ 0.061565f
C3026 FILLER_0_5_72/a_124_375# vdd -0.005497f
C3027 _394_/a_1336_472# FILLER_0_13_72/a_36_472# 0.008136f
C3028 _394_/a_728_93# FILLER_0_13_72/a_572_375# 0.001064f
C3029 _036_ _384_/a_224_472# 0.001921f
C3030 net82 _066_ 0.029681f
C3031 net26 FILLER_0_23_44/a_36_472# 0.013977f
C3032 _000_ _074_ 0.003542f
C3033 _015_ net64 1.212892f
C3034 _009_ _296_/a_224_472# 0.001278f
C3035 _016_ FILLER_0_12_124/a_36_472# 0.002661f
C3036 net65 _413_/a_2560_156# 0.011101f
C3037 cal_count\[3\] _055_ 0.039546f
C3038 FILLER_0_10_78/a_932_472# vss 0.002987f
C3039 net25 FILLER_0_23_60/a_124_375# 0.004431f
C3040 mask\[0\] FILLER_0_14_181/a_36_472# 0.001234f
C3041 _428_/a_2665_112# state\[2\] 0.001746f
C3042 FILLER_0_21_28/a_1828_472# _424_/a_36_151# 0.001723f
C3043 _413_/a_1204_472# net21 0.011236f
C3044 net35 FILLER_0_22_107/a_572_375# 0.010438f
C3045 mask\[8\] FILLER_0_22_107/a_36_472# 0.017159f
C3046 _216_/a_67_603# mask\[9\] 0.003086f
C3047 _098_ net71 1.076897f
C3048 _073_ cal_itt\[1\] 0.058541f
C3049 _069_ _068_ 0.003779f
C3050 net63 FILLER_0_18_177/a_484_472# 0.061539f
C3051 net20 _411_/a_448_472# 0.002167f
C3052 _267_/a_36_472# _090_ 0.001109f
C3053 fanout82/a_36_113# _316_/a_848_380# 0.001292f
C3054 net38 _445_/a_36_151# 0.112205f
C3055 _415_/a_36_151# FILLER_0_10_256/a_124_375# 0.035117f
C3056 FILLER_0_17_104/a_124_375# _451_/a_448_472# 0.001718f
C3057 FILLER_0_17_104/a_572_375# _451_/a_36_151# 0.001619f
C3058 _077_ FILLER_0_10_94/a_484_472# 0.001548f
C3059 _119_ _313_/a_255_603# 0.001151f
C3060 _195_/a_67_603# mask\[2\] 0.003161f
C3061 net82 FILLER_0_3_172/a_1828_472# 0.004472f
C3062 _079_ fanout75/a_36_113# 0.059598f
C3063 FILLER_0_15_116/a_36_472# _136_ 0.003818f
C3064 _128_ _061_ 0.76584f
C3065 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_572_375# 0.007947f
C3066 _072_ _248_/a_36_68# 0.001683f
C3067 _176_ _451_/a_448_472# 0.007191f
C3068 output14/a_224_472# _442_/a_2665_112# 0.009771f
C3069 FILLER_0_9_282/a_36_472# vdd 0.106034f
C3070 FILLER_0_9_282/a_572_375# vss 0.058599f
C3071 FILLER_0_4_107/a_36_472# _369_/a_36_68# 0.001709f
C3072 FILLER_0_4_144/a_36_472# _081_ 0.003547f
C3073 _414_/a_2248_156# net21 0.00415f
C3074 _132_ vdd 0.960634f
C3075 _277_/a_36_160# _099_ 0.001628f
C3076 _094_ net19 0.06304f
C3077 FILLER_0_5_54/a_572_375# _440_/a_36_151# 0.026916f
C3078 FILLER_0_8_138/a_124_375# vdd 0.024547f
C3079 vdd FILLER_0_22_107/a_484_472# 0.035591f
C3080 vss FILLER_0_22_107/a_36_472# 0.001514f
C3081 _094_ _418_/a_1204_472# 0.009231f
C3082 net20 net59 0.045227f
C3083 net82 net37 0.037195f
C3084 _046_ vss 0.088886f
C3085 _119_ _056_ 0.008929f
C3086 _028_ FILLER_0_7_72/a_932_472# 0.001777f
C3087 net58 net27 0.190417f
C3088 output13/a_224_472# vdd 0.045929f
C3089 FILLER_0_21_206/a_124_375# net33 0.001579f
C3090 _053_ vss 0.85895f
C3091 net20 net4 0.650415f
C3092 FILLER_0_7_195/a_124_375# cal_itt\[3\] 0.034632f
C3093 cal_itt\[2\] _073_ 0.202415f
C3094 net27 _425_/a_2665_112# 0.001323f
C3095 _072_ _060_ 0.080908f
C3096 _052_ FILLER_0_18_61/a_124_375# 0.006877f
C3097 net52 _440_/a_1308_423# 0.047012f
C3098 FILLER_0_15_282/a_484_472# result[3] 0.026996f
C3099 _321_/a_170_472# _395_/a_36_488# 0.007047f
C3100 FILLER_0_12_20/a_124_375# net6 0.003726f
C3101 ctln[2] net19 0.073057f
C3102 net17 _034_ 0.020793f
C3103 net72 _394_/a_56_524# 0.066156f
C3104 _053_ FILLER_0_7_72/a_2812_375# 0.016329f
C3105 _015_ vss 0.090048f
C3106 FILLER_0_23_282/a_124_375# FILLER_0_23_274/a_124_375# 0.003732f
C3107 _104_ _422_/a_2560_156# 0.003223f
C3108 mask\[4\] FILLER_0_18_177/a_1468_375# 0.01587f
C3109 _053_ net74 0.09773f
C3110 net50 FILLER_0_4_91/a_36_472# 0.058499f
C3111 net72 FILLER_0_19_28/a_572_375# 0.010026f
C3112 output7/a_224_472# net17 0.001164f
C3113 _443_/a_2665_112# trim_mask\[4\] 0.013708f
C3114 net76 _083_ 0.002446f
C3115 _256_/a_244_497# calibrate 0.002421f
C3116 _140_ FILLER_0_22_128/a_2724_472# 0.004196f
C3117 _432_/a_1308_423# _093_ 0.016365f
C3118 FILLER_0_15_290/a_36_472# _417_/a_36_151# 0.027236f
C3119 _126_ state\[2\] 0.030985f
C3120 net35 _214_/a_36_160# 0.0116f
C3121 FILLER_0_0_232/a_36_472# vss 0.007185f
C3122 fanout53/a_36_160# net56 0.196684f
C3123 _013_ FILLER_0_17_56/a_36_472# 0.002659f
C3124 _065_ _441_/a_36_151# 0.00701f
C3125 net48 _251_/a_244_472# 0.001259f
C3126 net64 net18 1.557441f
C3127 _017_ _043_ 0.02569f
C3128 output11/a_224_472# FILLER_0_0_198/a_124_375# 0.00363f
C3129 _256_/a_1612_497# net4 0.002497f
C3130 net81 FILLER_0_15_235/a_484_472# 0.0047f
C3131 output9/a_224_472# net2 0.003405f
C3132 _075_ _068_ 0.006297f
C3133 _077_ _133_ 0.003921f
C3134 FILLER_0_12_20/a_572_375# net40 0.007477f
C3135 _422_/a_1000_472# _109_ 0.003473f
C3136 _239_/a_36_160# _447_/a_36_151# 0.137659f
C3137 _070_ FILLER_0_10_107/a_572_375# 0.003959f
C3138 output32/a_224_472# result[7] 0.063135f
C3139 _428_/a_1204_472# vdd 0.001231f
C3140 _031_ FILLER_0_2_127/a_124_375# 0.013811f
C3141 _086_ _058_ 0.054155f
C3142 FILLER_0_5_54/a_572_375# vdd 0.004086f
C3143 net31 _199_/a_36_160# 0.007888f
C3144 _183_ FILLER_0_18_53/a_124_375# 0.001032f
C3145 output22/a_224_472# mask\[7\] 0.05527f
C3146 _086_ _315_/a_36_68# 0.003329f
C3147 FILLER_0_4_177/a_572_375# vdd 0.001622f
C3148 FILLER_0_4_177/a_124_375# vss 0.002462f
C3149 net57 FILLER_0_8_156/a_36_472# 0.001544f
C3150 FILLER_0_17_282/a_36_472# _417_/a_36_151# 0.001723f
C3151 FILLER_0_15_72/a_484_472# vdd 0.002283f
C3152 FILLER_0_15_72/a_36_472# vss 0.038986f
C3153 _415_/a_448_472# net19 0.03569f
C3154 FILLER_0_12_2/a_572_375# net6 0.058881f
C3155 output28/a_224_472# net28 0.048681f
C3156 _445_/a_2248_156# net17 0.06175f
C3157 _428_/a_1000_472# net74 0.00735f
C3158 FILLER_0_15_116/a_484_472# net53 0.002804f
C3159 net50 vdd 0.661261f
C3160 net20 FILLER_0_13_212/a_1020_375# 0.003962f
C3161 FILLER_0_4_99/a_124_375# _160_ 0.005563f
C3162 _440_/a_448_472# _164_ 0.0036f
C3163 FILLER_0_22_177/a_36_472# _434_/a_448_472# 0.012285f
C3164 _141_ FILLER_0_19_155/a_36_472# 0.05777f
C3165 net55 FILLER_0_18_76/a_124_375# 0.001706f
C3166 _443_/a_1000_472# vss 0.031435f
C3167 net1 cal_itt\[1\] 0.229522f
C3168 output44/a_224_472# vdd 0.043902f
C3169 _033_ FILLER_0_6_37/a_36_472# 0.017695f
C3170 FILLER_0_19_28/a_124_375# net40 0.047489f
C3171 FILLER_0_7_72/a_2364_375# net50 0.017301f
C3172 vss _433_/a_3041_156# 0.001287f
C3173 output28/a_224_472# _416_/a_2248_156# 0.023576f
C3174 result[1] _416_/a_448_472# 0.008784f
C3175 _074_ _081_ 0.070546f
C3176 _378_/a_224_472# _165_ 0.00481f
C3177 net27 _426_/a_796_472# 0.001678f
C3178 _444_/a_448_472# net42 0.002526f
C3179 net18 vss 1.110302f
C3180 _176_ FILLER_0_17_72/a_1828_472# 0.001028f
C3181 valid net1 0.00347f
C3182 FILLER_0_16_57/a_572_375# _131_ 0.015859f
C3183 _067_ FILLER_0_13_72/a_572_375# 0.001874f
C3184 fanout78/a_36_113# _094_ 0.01312f
C3185 fanout56/a_36_113# net36 0.021321f
C3186 net19 FILLER_0_23_274/a_36_472# 0.075097f
C3187 FILLER_0_17_64/a_124_375# FILLER_0_17_56/a_572_375# 0.012001f
C3188 _174_ cal_count\[0\] 0.009645f
C3189 FILLER_0_15_72/a_36_472# cal_count\[1\] 0.006408f
C3190 net55 _424_/a_2560_156# 0.003707f
C3191 net15 FILLER_0_15_72/a_124_375# 0.006566f
C3192 _078_ _080_ 0.030094f
C3193 net16 FILLER_0_18_37/a_36_472# 0.001132f
C3194 _001_ _082_ 0.46787f
C3195 FILLER_0_18_2/a_1020_375# net44 0.009108f
C3196 _069_ vdd 0.985405f
C3197 result[9] result[2] 0.001669f
C3198 _308_/a_124_24# net14 0.005016f
C3199 _090_ _113_ 0.263235f
C3200 FILLER_0_18_2/a_2724_472# net55 0.007511f
C3201 _360_/a_36_160# vss 0.028817f
C3202 net34 FILLER_0_22_177/a_124_375# 0.006974f
C3203 net29 vdd 0.611195f
C3204 _371_/a_36_113# FILLER_0_2_127/a_124_375# 0.002437f
C3205 ctlp[1] _419_/a_796_472# 0.001178f
C3206 FILLER_0_10_78/a_124_375# FILLER_0_9_72/a_932_472# 0.001543f
C3207 _432_/a_36_151# mask\[1\] 0.003001f
C3208 _232_/a_255_603# net47 0.001241f
C3209 FILLER_0_3_204/a_36_472# net82 0.008268f
C3210 output25/a_224_472# vdd 0.03413f
C3211 FILLER_0_15_142/a_124_375# vdd -0.003809f
C3212 trim_mask\[3\] vdd 0.233305f
C3213 _164_ vss 0.597051f
C3214 _431_/a_2665_112# FILLER_0_17_142/a_572_375# 0.001092f
C3215 _431_/a_2560_156# FILLER_0_17_142/a_124_375# 0.001178f
C3216 output48/a_224_472# _082_ 0.002393f
C3217 _433_/a_1000_472# _145_ 0.004227f
C3218 _414_/a_2665_112# _074_ 0.004912f
C3219 FILLER_0_18_37/a_1468_375# vdd 0.021186f
C3220 _008_ vdd 0.284571f
C3221 _259_/a_455_68# net20 0.001427f
C3222 _360_/a_36_160# net74 0.001912f
C3223 FILLER_0_10_78/a_484_472# cal_count\[3\] 0.001112f
C3224 _102_ _099_ 0.151018f
C3225 _322_/a_124_24# _070_ 0.033355f
C3226 _091_ FILLER_0_19_171/a_932_472# 0.002509f
C3227 _440_/a_2665_112# _160_ 0.008418f
C3228 FILLER_0_6_90/a_572_375# net14 0.031929f
C3229 net64 net62 0.078454f
C3230 _227_/a_36_160# FILLER_0_8_156/a_124_375# 0.005398f
C3231 _116_ FILLER_0_13_206/a_124_375# 0.003926f
C3232 net20 net79 0.046876f
C3233 mask\[9\] FILLER_0_20_98/a_124_375# 0.003444f
C3234 _404_/a_36_472# _182_ 0.036415f
C3235 cal_count\[2\] _402_/a_718_527# 0.004645f
C3236 _411_/a_448_472# _073_ 0.004279f
C3237 mask\[1\] net62 0.227329f
C3238 fanout57/a_36_113# vss 0.046378f
C3239 _448_/a_2665_112# _170_ 0.002715f
C3240 _448_/a_1204_472# _037_ 0.008883f
C3241 FILLER_0_4_144/a_124_375# trim_mask\[4\] 0.014395f
C3242 result[8] _435_/a_2665_112# 0.001855f
C3243 _265_/a_244_68# _001_ 0.008874f
C3244 _053_ _119_ 0.038651f
C3245 _118_ _090_ 0.005469f
C3246 FILLER_0_4_197/a_932_472# net82 0.001826f
C3247 output34/a_224_472# net19 0.001308f
C3248 net66 net40 0.124825f
C3249 _436_/a_448_472# _025_ 0.044246f
C3250 _441_/a_796_472# _030_ 0.024278f
C3251 net34 _419_/a_2665_112# 0.001468f
C3252 result[7] _419_/a_1204_472# 0.018181f
C3253 FILLER_0_16_89/a_1380_472# vss 0.005351f
C3254 trim_mask\[2\] net66 0.036211f
C3255 FILLER_0_4_152/a_124_375# _170_ 0.029927f
C3256 _013_ _131_ 0.001178f
C3257 fanout53/a_36_160# _095_ 0.007436f
C3258 net39 _034_ 0.004367f
C3259 _075_ vdd 0.190898f
C3260 _321_/a_170_472# _125_ 0.008492f
C3261 FILLER_0_17_226/a_124_375# _093_ 0.001604f
C3262 _073_ net59 0.028673f
C3263 _112_ _001_ 0.002527f
C3264 _432_/a_448_472# vdd 0.035246f
C3265 _432_/a_36_151# vss 0.003647f
C3266 _036_ _441_/a_36_151# 0.005754f
C3267 _021_ _093_ 0.049589f
C3268 _445_/a_1308_423# net40 0.046345f
C3269 _073_ net4 0.076114f
C3270 _009_ FILLER_0_23_274/a_36_472# 0.005531f
C3271 FILLER_0_18_209/a_484_472# vdd 0.00367f
C3272 FILLER_0_18_209/a_36_472# vss 0.005442f
C3273 net49 _440_/a_2248_156# 0.025137f
C3274 _414_/a_1288_156# cal_itt\[3\] 0.001354f
C3275 net64 FILLER_0_15_235/a_572_375# 0.007219f
C3276 FILLER_0_20_177/a_124_375# vdd 0.001964f
C3277 ctln[3] vss 0.133697f
C3278 _322_/a_848_380# FILLER_0_9_142/a_124_375# 0.001721f
C3279 _103_ _046_ 0.010317f
C3280 net32 _419_/a_2248_156# 0.034827f
C3281 _104_ _294_/a_224_472# 0.003008f
C3282 trim_mask\[4\] net69 0.185121f
C3283 _431_/a_796_472# _020_ 0.012284f
C3284 _442_/a_2665_112# _157_ 0.001587f
C3285 net38 _221_/a_36_160# 0.029767f
C3286 _091_ FILLER_0_15_212/a_572_375# 0.022582f
C3287 FILLER_0_15_235/a_572_375# mask\[1\] 0.013718f
C3288 output48/a_224_472# _112_ 0.027383f
C3289 fanout80/a_36_113# _019_ 0.003644f
C3290 FILLER_0_11_109/a_124_375# FILLER_0_10_107/a_484_472# 0.001684f
C3291 output23/a_224_472# FILLER_0_22_128/a_2364_375# 0.002439f
C3292 _057_ _069_ 0.053765f
C3293 _198_/a_67_603# _099_ 0.0109f
C3294 FILLER_0_18_61/a_36_472# vss 0.00605f
C3295 output8/a_224_472# cal_itt\[1\] 0.003894f
C3296 _028_ FILLER_0_6_90/a_124_375# 0.012573f
C3297 FILLER_0_16_255/a_124_375# net30 0.001055f
C3298 vss net62 1.17087f
C3299 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_124_375# 0.012001f
C3300 _116_ _311_/a_66_473# 0.001527f
C3301 _091_ mask\[0\] 0.04171f
C3302 _087_ net22 0.028009f
C3303 FILLER_0_17_104/a_1468_375# vss 0.001786f
C3304 FILLER_0_17_104/a_36_472# vdd 0.095484f
C3305 result[9] _419_/a_448_472# 0.015767f
C3306 ctln[0] vdd 0.051631f
C3307 FILLER_0_5_54/a_484_472# FILLER_0_6_47/a_1380_472# 0.026657f
C3308 FILLER_0_5_54/a_1468_375# FILLER_0_6_47/a_2276_472# 0.001597f
C3309 _105_ output18/a_224_472# 0.105478f
C3310 _067_ net40 0.040115f
C3311 _110_ _098_ 0.09704f
C3312 net31 net33 0.002465f
C3313 net82 _122_ 0.001375f
C3314 _426_/a_2248_156# _076_ 0.015189f
C3315 _402_/a_56_567# net47 0.026503f
C3316 _196_/a_36_160# _045_ 0.036714f
C3317 _413_/a_796_472# _002_ 0.009261f
C3318 net39 _445_/a_2248_156# 0.003571f
C3319 output37/a_224_472# net5 0.072504f
C3320 net52 FILLER_0_9_72/a_572_375# 0.022582f
C3321 FILLER_0_15_59/a_124_375# vdd 0.017243f
C3322 FILLER_0_21_286/a_572_375# net77 0.044323f
C3323 net20 _274_/a_716_497# 0.001321f
C3324 mask\[3\] _099_ 0.10534f
C3325 net48 _317_/a_36_113# 0.018494f
C3326 ctln[6] ctln[7] 0.00499f
C3327 net57 _395_/a_36_488# 0.026081f
C3328 net24 _050_ 0.049889f
C3329 net75 _316_/a_848_380# 0.044673f
C3330 FILLER_0_4_49/a_36_472# _167_ 0.063278f
C3331 output8/a_224_472# cal_itt\[2\] 0.05561f
C3332 net44 _452_/a_2225_156# 0.044858f
C3333 _283_/a_36_472# _099_ 0.004667f
C3334 net63 _092_ 0.008819f
C3335 _412_/a_796_472# net2 0.00566f
C3336 FILLER_0_11_64/a_36_472# _120_ 0.011673f
C3337 FILLER_0_21_142/a_36_472# _210_/a_67_603# 0.001547f
C3338 FILLER_0_19_171/a_1020_375# vdd 0.025918f
C3339 FILLER_0_20_87/a_36_472# net14 0.001471f
C3340 _348_/a_49_472# mask\[6\] 0.005525f
C3341 net52 cal_count\[3\] 0.348542f
C3342 state\[2\] FILLER_0_13_142/a_932_472# 0.004118f
C3343 _159_ net47 0.01358f
C3344 _205_/a_36_160# net21 0.020847f
C3345 FILLER_0_15_235/a_572_375# vss 0.002683f
C3346 FILLER_0_15_235/a_36_472# vdd 0.019127f
C3347 trim_val\[3\] vss 0.249446f
C3348 _132_ _433_/a_36_151# 0.024768f
C3349 FILLER_0_18_177/a_2812_375# net21 0.048071f
C3350 _438_/a_36_151# vdd 0.111691f
C3351 _063_ _444_/a_2665_112# 0.001996f
C3352 _432_/a_796_472# _098_ 0.038458f
C3353 _072_ vss 0.439154f
C3354 net52 _154_ 0.001512f
C3355 _068_ net22 0.088209f
C3356 FILLER_0_20_107/a_36_472# _098_ 0.011046f
C3357 FILLER_0_10_28/a_124_375# net51 0.00979f
C3358 result[2] FILLER_0_13_290/a_124_375# 0.015011f
C3359 net20 fanout63/a_36_160# 0.084165f
C3360 ctln[4] FILLER_0_1_204/a_36_472# 0.006408f
C3361 fanout69/a_36_113# net69 0.040451f
C3362 _414_/a_36_151# FILLER_0_6_177/a_484_472# 0.006095f
C3363 vdd result[3] 0.181788f
C3364 FILLER_0_9_28/a_1468_375# net68 0.013121f
C3365 FILLER_0_2_93/a_484_472# net69 0.0127f
C3366 _443_/a_2665_112# _066_ 0.001654f
C3367 net73 FILLER_0_18_107/a_36_472# 0.002425f
C3368 FILLER_0_0_130/a_36_472# vdd 0.050082f
C3369 FILLER_0_0_130/a_124_375# vss 0.018073f
C3370 mask\[5\] _145_ 0.012075f
C3371 FILLER_0_16_89/a_1020_375# net14 0.029702f
C3372 FILLER_0_24_96/a_124_375# vdd 0.029269f
C3373 _131_ _179_ 0.034602f
C3374 FILLER_0_16_107/a_36_472# _136_ 0.011469f
C3375 net1 net59 0.920133f
C3376 _430_/a_2248_156# vdd 0.008989f
C3377 net54 mask\[7\] 0.262465f
C3378 _132_ _093_ 0.105039f
C3379 net64 FILLER_0_8_247/a_1380_472# 0.001021f
C3380 _076_ _118_ 0.06281f
C3381 _136_ FILLER_0_17_133/a_124_375# 0.001315f
C3382 FILLER_0_4_99/a_124_375# _156_ 0.081915f
C3383 net41 cal_count\[3\] 0.028902f
C3384 net1 net4 0.03357f
C3385 _230_/a_244_68# net21 0.00165f
C3386 FILLER_0_20_98/a_36_472# vss 0.00206f
C3387 net54 _148_ 0.098648f
C3388 FILLER_0_18_107/a_484_472# mask\[9\] 0.001955f
C3389 result[9] _420_/a_2665_112# 0.037019f
C3390 FILLER_0_19_47/a_572_375# _183_ 0.001186f
C3391 net19 FILLER_0_14_263/a_124_375# 0.032085f
C3392 _123_ FILLER_0_6_231/a_572_375# 0.00487f
C3393 _311_/a_66_473# _117_ 0.001055f
C3394 _103_ net18 0.11279f
C3395 net57 calibrate 0.037299f
C3396 FILLER_0_18_139/a_1468_375# net23 0.04546f
C3397 _426_/a_1000_472# net64 0.008796f
C3398 _189_/a_67_603# _100_ 0.002818f
C3399 _132_ FILLER_0_19_134/a_124_375# 0.00141f
C3400 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_124_375# 0.026339f
C3401 _420_/a_1000_472# vss 0.002146f
C3402 net20 FILLER_0_1_212/a_124_375# 0.084041f
C3403 vdd _450_/a_1040_527# 0.005529f
C3404 output23/a_224_472# _050_ 0.014495f
C3405 net53 _451_/a_36_151# 0.030715f
C3406 net70 _451_/a_1040_527# 0.002679f
C3407 _109_ vss 0.023215f
C3408 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_572_375# 0.086635f
C3409 FILLER_0_8_247/a_36_472# _316_/a_124_24# 0.001386f
C3410 _313_/a_67_603# _120_ 0.005873f
C3411 _291_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C3412 _186_ _095_ 0.042856f
C3413 net19 _419_/a_1000_472# 0.012949f
C3414 mask\[3\] FILLER_0_17_218/a_36_472# 0.015535f
C3415 _376_/a_36_160# FILLER_0_6_79/a_124_375# 0.004736f
C3416 _449_/a_2248_156# _038_ 0.016483f
C3417 FILLER_0_16_57/a_1380_472# _176_ 0.01346f
C3418 FILLER_0_13_142/a_36_472# vdd 0.104785f
C3419 _136_ mask\[9\] 0.015204f
C3420 fanout53/a_36_160# vss 0.006674f
C3421 FILLER_0_13_142/a_1468_375# vss 0.00614f
C3422 FILLER_0_18_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001684f
C3423 net41 FILLER_0_21_28/a_932_472# 0.014034f
C3424 net67 output6/a_224_472# 0.070024f
C3425 _382_/a_224_472# vdd 0.001663f
C3426 FILLER_0_8_107/a_124_375# _133_ 0.048874f
C3427 FILLER_0_8_107/a_36_472# _070_ 0.001287f
C3428 _008_ net78 0.032202f
C3429 _008_ net60 0.314106f
C3430 FILLER_0_7_59/a_572_375# net68 0.005738f
C3431 _069_ _314_/a_224_472# 0.003461f
C3432 _430_/a_36_151# FILLER_0_17_200/a_484_472# 0.001723f
C3433 FILLER_0_8_247/a_1380_472# vss 0.001338f
C3434 FILLER_0_5_88/a_36_472# _163_ 0.006541f
C3435 _421_/a_2665_112# vdd 0.029293f
C3436 net72 cal_count\[2\] 0.073818f
C3437 net49 net14 0.00344f
C3438 cal_itt\[3\] _163_ 0.021146f
C3439 trimb[0] vss 0.097724f
C3440 _442_/a_2248_156# net14 0.025334f
C3441 _067_ FILLER_0_13_80/a_124_375# 0.001857f
C3442 ctln[5] _448_/a_448_472# 0.010887f
C3443 net52 FILLER_0_3_78/a_484_472# 0.003143f
C3444 output27/a_224_472# vdd 0.070751f
C3445 _076_ _068_ 0.35956f
C3446 net32 _297_/a_36_472# 0.001843f
C3447 _422_/a_1308_423# vdd 0.004083f
C3448 result[4] net79 0.048452f
C3449 FILLER_0_10_256/a_36_472# net27 0.008331f
C3450 cal_count\[3\] _172_ 0.03048f
C3451 net80 net33 0.037227f
C3452 _356_/a_36_472# mask\[9\] 0.047632f
C3453 _426_/a_1204_472# vdd 0.003412f
C3454 _415_/a_36_151# _416_/a_1308_423# 0.00119f
C3455 _444_/a_36_151# net49 0.007102f
C3456 ctlp[4] _108_ 0.002002f
C3457 _132_ _436_/a_36_151# 0.00162f
C3458 _326_/a_36_160# _134_ 0.003299f
C3459 FILLER_0_15_282/a_572_375# vss 0.058168f
C3460 FILLER_0_15_282/a_36_472# vdd 0.10628f
C3461 _432_/a_36_151# _097_ 0.003144f
C3462 _446_/a_2665_112# net40 0.027712f
C3463 trim[4] clkc 0.005f
C3464 _436_/a_36_151# FILLER_0_22_107/a_484_472# 0.001723f
C3465 _074_ _161_ 0.191658f
C3466 FILLER_0_11_101/a_484_472# vdd 0.009482f
C3467 FILLER_0_11_101/a_36_472# vss 0.001641f
C3468 _090_ vdd 0.751973f
C3469 fanout61/a_36_113# vdd 0.108255f
C3470 _088_ FILLER_0_4_213/a_484_472# 0.018066f
C3471 _112_ _316_/a_124_24# 0.032665f
C3472 FILLER_0_3_221/a_124_375# vss 0.034009f
C3473 _058_ _120_ 0.008566f
C3474 FILLER_0_4_49/a_572_375# _164_ 0.005532f
C3475 net34 _146_ 0.004718f
C3476 net66 trim[3] 0.00567f
C3477 _315_/a_36_68# _120_ 0.00572f
C3478 net17 FILLER_0_23_44/a_36_472# 0.071244f
C3479 _144_ _350_/a_49_472# 0.033348f
C3480 net63 _435_/a_2665_112# 0.039512f
C3481 output8/a_224_472# _411_/a_448_472# 0.010723f
C3482 state\[2\] _095_ 0.001426f
C3483 fanout55/a_36_160# _043_ 0.019538f
C3484 _176_ _182_ 0.008217f
C3485 net73 net53 0.094507f
C3486 net65 net37 0.008382f
C3487 _420_/a_448_472# net77 0.001276f
C3488 _413_/a_36_151# net59 0.02781f
C3489 _021_ net57 0.00736f
C3490 net31 _046_ 0.008368f
C3491 _321_/a_170_472# _069_ 0.025551f
C3492 net22 vdd 1.920713f
C3493 net20 ctlp[2] 0.254928f
C3494 FILLER_0_15_150/a_124_375# net23 0.03361f
C3495 _093_ _069_ 0.008325f
C3496 _077_ FILLER_0_8_156/a_484_472# 0.006446f
C3497 output8/a_224_472# net59 0.00398f
C3498 _414_/a_36_151# _055_ 0.001987f
C3499 _178_ _180_ 0.004668f
C3500 _077_ net37 0.003374f
C3501 FILLER_0_8_24/a_572_375# net40 0.038492f
C3502 net81 vdd 1.658963f
C3503 fanout80/a_36_113# net80 0.004615f
C3504 FILLER_0_3_78/a_36_472# _164_ 0.022063f
C3505 _125_ _135_ 0.001926f
C3506 _015_ FILLER_0_10_247/a_36_472# 0.007508f
C3507 FILLER_0_17_56/a_36_472# _041_ 0.004881f
C3508 _313_/a_67_603# _227_/a_36_160# 0.032438f
C3509 output8/a_224_472# net4 0.015359f
C3510 _081_ FILLER_0_5_148/a_572_375# 0.01425f
C3511 _436_/a_2560_156# _050_ 0.01099f
C3512 _043_ FILLER_0_13_72/a_36_472# 0.017766f
C3513 net26 net40 0.001136f
C3514 net26 _424_/a_448_472# 0.063966f
C3515 FILLER_0_2_101/a_36_472# trim_mask\[3\] 0.013363f
C3516 FILLER_0_18_107/a_1380_472# vdd 0.009462f
C3517 fanout67/a_36_160# _220_/a_67_603# 0.005474f
C3518 _119_ _072_ 0.189217f
C3519 _413_/a_2560_156# vss 0.001097f
C3520 _217_/a_36_160# vdd 0.092586f
C3521 _406_/a_36_159# _278_/a_36_160# 0.001331f
C3522 net61 _419_/a_448_472# 0.024246f
C3523 _208_/a_36_160# FILLER_0_22_128/a_3260_375# 0.001948f
C3524 _049_ FILLER_0_22_128/a_3172_472# 0.01125f
C3525 _008_ _093_ 0.252609f
C3526 vss FILLER_0_10_94/a_484_472# 0.001244f
C3527 FILLER_0_14_107/a_36_472# _451_/a_36_151# 0.001723f
C3528 _448_/a_2560_156# net22 0.00766f
C3529 net54 FILLER_0_22_128/a_932_472# 0.014735f
C3530 _322_/a_848_380# _127_ 0.018892f
C3531 FILLER_0_16_89/a_36_472# _040_ 0.015634f
C3532 _417_/a_796_472# _006_ 0.014427f
C3533 _058_ FILLER_0_9_105/a_572_375# 0.003832f
C3534 output43/a_224_472# output46/a_224_472# 0.292611f
C3535 output47/a_224_472# _452_/a_3129_107# 0.018181f
C3536 FILLER_0_21_28/a_3260_375# _012_ 0.016427f
C3537 fanout77/a_36_113# net77 0.031558f
C3538 _035_ vdd 0.215473f
C3539 net69 _367_/a_36_68# 0.008893f
C3540 net63 FILLER_0_17_226/a_36_472# 0.001822f
C3541 FILLER_0_5_164/a_36_472# _163_ 0.001777f
C3542 _422_/a_2665_112# net19 0.006987f
C3543 FILLER_0_18_171/a_124_375# _098_ 0.032114f
C3544 _372_/a_170_472# _122_ 0.018399f
C3545 _129_ calibrate 0.04134f
C3546 FILLER_0_10_78/a_484_472# _120_ 0.004669f
C3547 _294_/a_224_472# mask\[2\] 0.001715f
C3548 _038_ vdd 0.043998f
C3549 _057_ _090_ 0.112325f
C3550 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001597f
C3551 net55 FILLER_0_17_38/a_124_375# 0.003236f
C3552 net72 FILLER_0_17_38/a_484_472# 0.00547f
C3553 net23 _242_/a_36_160# 0.007466f
C3554 _432_/a_448_472# _093_ 0.048289f
C3555 FILLER_0_16_255/a_124_375# _417_/a_2665_112# 0.003856f
C3556 _162_ _062_ 0.033583f
C3557 _186_ vss 0.0718f
C3558 net10 net75 0.073869f
C3559 net20 _000_ 0.159624f
C3560 net60 result[3] 0.001124f
C3561 net4 FILLER_0_12_220/a_124_375# 0.016485f
C3562 FILLER_0_22_177/a_484_472# mask\[6\] 0.006573f
C3563 FILLER_0_22_177/a_124_375# _146_ 0.001864f
C3564 mask\[5\] _202_/a_36_160# 0.00164f
C3565 _093_ FILLER_0_18_209/a_484_472# 0.014737f
C3566 _450_/a_3129_107# _039_ 0.012762f
C3567 _176_ _040_ 0.272465f
C3568 trim_mask\[1\] FILLER_0_6_90/a_484_472# 0.014443f
C3569 _058_ _227_/a_36_160# 0.008511f
C3570 net19 _001_ 0.018424f
C3571 net54 FILLER_0_22_107/a_124_375# 0.003502f
C3572 _133_ vss 0.18326f
C3573 _076_ vdd 0.806117f
C3574 _449_/a_1000_472# vss 0.029565f
C3575 FILLER_0_18_100/a_124_375# _438_/a_2248_156# 0.001068f
C3576 net28 net29 0.178557f
C3577 _440_/a_2248_156# net47 0.017063f
C3578 _057_ net22 0.163773f
C3579 mask\[8\] FILLER_0_22_86/a_1468_375# 0.015339f
C3580 net35 FILLER_0_22_86/a_1020_375# 0.010202f
C3581 net52 _442_/a_1308_423# 0.017208f
C3582 net55 FILLER_0_18_37/a_1380_472# 0.007432f
C3583 _114_ _311_/a_2180_473# 0.00515f
C3584 _132_ net57 0.029479f
C3585 net32 _006_ 0.0012f
C3586 net31 net18 0.114197f
C3587 FILLER_0_17_72/a_3260_375# vdd 0.007427f
C3588 _376_/a_36_160# vss 0.03081f
C3589 net21 _047_ 0.048701f
C3590 _069_ _429_/a_1204_472# 0.025254f
C3591 _075_ FILLER_0_5_206/a_124_375# 0.001024f
C3592 fanout59/a_36_160# net64 0.006298f
C3593 _183_ _182_ 0.002134f
C3594 _093_ FILLER_0_17_104/a_36_472# 0.014431f
C3595 output48/a_224_472# net19 0.054227f
C3596 net74 _133_ 0.696379f
C3597 _429_/a_36_151# _043_ 0.002771f
C3598 _321_/a_3662_472# _176_ 0.002006f
C3599 _186_ cal_count\[1\] 0.003341f
C3600 trimb[1] FILLER_0_18_2/a_36_472# 0.010728f
C3601 _095_ FILLER_0_14_107/a_932_472# 0.014431f
C3602 _128_ _426_/a_2248_156# 0.019019f
C3603 net44 FILLER_0_15_2/a_36_472# 0.007808f
C3604 FILLER_0_22_86/a_36_472# vdd -0.001506f
C3605 FILLER_0_22_86/a_1468_375# vss 0.013146f
C3606 _132_ _135_ 0.345161f
C3607 _090_ _279_/a_244_68# 0.001986f
C3608 _192_/a_255_603# mask\[1\] 0.001059f
C3609 net33 _434_/a_448_472# 0.003049f
C3610 FILLER_0_9_28/a_2276_472# _053_ 0.002243f
C3611 output36/a_224_472# _006_ 0.022685f
C3612 _114_ _061_ 0.123371f
C3613 FILLER_0_12_2/a_484_472# net44 0.046864f
C3614 FILLER_0_24_63/a_36_472# _423_/a_2665_112# 0.001873f
C3615 _131_ FILLER_0_17_56/a_572_375# 0.006224f
C3616 FILLER_0_7_59/a_36_472# net67 0.021549f
C3617 _128_ _113_ 0.002117f
C3618 FILLER_0_24_130/a_36_472# output24/a_224_472# 0.023414f
C3619 FILLER_0_3_204/a_36_472# net65 0.001777f
C3620 net81 net2 1.204674f
C3621 _422_/a_2665_112# _009_ 0.061508f
C3622 mask\[8\] _437_/a_2665_112# 0.007907f
C3623 _449_/a_1308_423# net15 0.015651f
C3624 FILLER_0_13_212/a_1020_375# FILLER_0_12_220/a_124_375# 0.05841f
C3625 net41 FILLER_0_18_2/a_3172_472# 0.00982f
C3626 state\[2\] vss 0.185787f
C3627 input1/a_36_113# clk 0.001121f
C3628 _411_/a_2248_156# net8 0.06032f
C3629 net41 _445_/a_448_472# 0.002211f
C3630 FILLER_0_11_101/a_572_375# cal_count\[3\] 0.002017f
C3631 _093_ _438_/a_36_151# 0.088469f
C3632 net20 _421_/a_1000_472# 0.012469f
C3633 net60 _421_/a_2665_112# 0.044114f
C3634 _219_/a_36_160# _439_/a_2665_112# 0.002537f
C3635 _437_/a_2665_112# vss 0.002056f
C3636 _437_/a_2560_156# vdd 0.0026f
C3637 _444_/a_448_472# net67 0.046278f
C3638 _129_ _125_ 0.069221f
C3639 net53 _427_/a_36_151# 0.13192f
C3640 output19/a_224_472# _107_ 0.005034f
C3641 _131_ _041_ 0.035642f
C3642 net57 _428_/a_1204_472# 0.015233f
C3643 trim_mask\[1\] FILLER_0_5_88/a_124_375# 0.072632f
C3644 net61 _422_/a_1000_472# 0.001947f
C3645 _429_/a_36_151# net21 0.054289f
C3646 net82 _170_ 0.080348f
C3647 FILLER_0_7_195/a_124_375# _161_ 0.005368f
C3648 FILLER_0_17_282/a_124_375# _006_ 0.004694f
C3649 FILLER_0_9_60/a_572_375# _439_/a_36_151# 0.001107f
C3650 net52 _120_ 0.023363f
C3651 _004_ net19 0.112289f
C3652 state\[2\] net74 0.024462f
C3653 fanout59/a_36_160# vss 0.010949f
C3654 state\[0\] _426_/a_2248_156# 0.001198f
C3655 FILLER_0_22_177/a_36_472# _023_ 0.007019f
C3656 _029_ _164_ 0.031781f
C3657 trim_mask\[4\] vss 0.641217f
C3658 _128_ _118_ 0.58787f
C3659 _127_ _124_ 0.035569f
C3660 FILLER_0_16_89/a_124_375# _176_ 0.002781f
C3661 _028_ FILLER_0_7_104/a_1020_375# 0.004954f
C3662 _086_ FILLER_0_7_104/a_1380_472# 0.034829f
C3663 net34 _435_/a_448_472# 0.013341f
C3664 _105_ _297_/a_36_472# 0.03208f
C3665 fanout61/a_36_113# net78 0.009579f
C3666 vdd FILLER_0_4_91/a_572_375# 0.019853f
C3667 _236_/a_36_160# _064_ 0.039922f
C3668 _043_ FILLER_0_15_180/a_36_472# 0.001219f
C3669 _057_ _076_ 0.041986f
C3670 _086_ _318_/a_224_472# 0.007024f
C3671 mask\[5\] _107_ 0.01249f
C3672 fanout71/a_36_113# vss 0.007654f
C3673 _141_ FILLER_0_18_139/a_1380_472# 0.016119f
C3674 _402_/a_1296_93# _401_/a_36_68# 0.001523f
C3675 _087_ FILLER_0_5_172/a_124_375# 0.003043f
C3676 FILLER_0_5_128/a_484_472# _133_ 0.037369f
C3677 FILLER_0_11_78/a_484_472# vdd 0.001756f
C3678 FILLER_0_11_78/a_36_472# vss 0.00471f
C3679 output20/a_224_472# vdd 0.09529f
C3680 _160_ _034_ 0.00905f
C3681 mask\[3\] FILLER_0_16_154/a_932_472# 0.002604f
C3682 net74 trim_mask\[4\] 0.548293f
C3683 _444_/a_1308_423# _054_ 0.005457f
C3684 net81 FILLER_0_12_236/a_572_375# 0.021025f
C3685 net16 vdd 2.255325f
C3686 FILLER_0_12_20/a_124_375# _450_/a_448_472# 0.001597f
C3687 _416_/a_2665_112# net62 0.037195f
C3688 net20 _081_ 0.024512f
C3689 net43 vss 0.132286f
C3690 _429_/a_2248_156# net62 0.012262f
C3691 FILLER_0_16_107/a_484_472# FILLER_0_16_115/a_36_472# 0.013276f
C3692 FILLER_0_21_133/a_36_472# mask\[7\] 0.003404f
C3693 _444_/a_1308_423# FILLER_0_8_24/a_36_472# 0.009119f
C3694 FILLER_0_7_104/a_1380_472# _154_ 0.002799f
C3695 _423_/a_1308_423# _012_ 0.01389f
C3696 _422_/a_1000_472# _108_ 0.027806f
C3697 _430_/a_448_472# net36 0.011598f
C3698 _412_/a_36_151# net1 0.020184f
C3699 result[9] vss 0.348416f
C3700 FILLER_0_4_185/a_124_375# FILLER_0_4_177/a_572_375# 0.012001f
C3701 _077_ _439_/a_2560_156# 0.012523f
C3702 _327_/a_36_472# _016_ 0.04536f
C3703 net79 _286_/a_224_472# 0.001276f
C3704 _031_ _369_/a_36_68# 0.050502f
C3705 net57 _069_ 0.026933f
C3706 _116_ _085_ 0.049304f
C3707 ctln[4] net75 0.00718f
C3708 FILLER_0_13_100/a_124_375# net14 0.041373f
C3709 FILLER_0_3_172/a_2724_472# net22 0.012284f
C3710 net79 FILLER_0_12_220/a_124_375# 0.010895f
C3711 _427_/a_2665_112# _043_ 0.002612f
C3712 _081_ _163_ 0.427672f
C3713 _055_ net21 0.025995f
C3714 FILLER_0_4_144/a_36_472# net23 0.016933f
C3715 net20 _413_/a_2248_156# 0.002515f
C3716 FILLER_0_23_282/a_36_472# vss 0.003317f
C3717 _430_/a_2560_156# _092_ 0.001333f
C3718 fanout51/a_36_113# FILLER_0_11_78/a_124_375# 0.005683f
C3719 mask\[4\] _141_ 0.948091f
C3720 _424_/a_2248_156# _012_ 0.009377f
C3721 FILLER_0_7_72/a_1468_375# vss 0.003253f
C3722 FILLER_0_7_72/a_1916_375# vdd 0.015888f
C3723 output16/a_224_472# net15 0.013768f
C3724 _077_ _122_ 0.144611f
C3725 output42/a_224_472# FILLER_0_8_24/a_124_375# 0.001168f
C3726 cal_count\[3\] _136_ 0.00703f
C3727 _128_ _068_ 0.863174f
C3728 net58 result[1] 0.004614f
C3729 _445_/a_1000_472# _034_ 0.007034f
C3730 _445_/a_2665_112# _166_ 0.002292f
C3731 net35 FILLER_0_22_177/a_484_472# 0.00632f
C3732 fanout69/a_36_113# vss 0.002239f
C3733 cal_itt\[1\] FILLER_0_3_221/a_1380_472# 0.004939f
C3734 _062_ FILLER_0_8_156/a_124_375# 0.008116f
C3735 FILLER_0_22_86/a_932_472# net71 0.005789f
C3736 net70 net14 0.106631f
C3737 result[6] FILLER_0_21_286/a_124_375# 0.019179f
C3738 output37/a_224_472# en 0.003788f
C3739 FILLER_0_2_93/a_484_472# vss 0.003689f
C3740 _002_ FILLER_0_3_172/a_3260_375# 0.001683f
C3741 _052_ FILLER_0_21_28/a_2364_375# 0.002388f
C3742 _119_ _133_ 0.038875f
C3743 _086_ _070_ 0.123033f
C3744 FILLER_0_10_78/a_36_472# _115_ 0.002611f
C3745 _000_ _073_ 0.222349f
C3746 net47 net14 0.033547f
C3747 FILLER_0_21_28/a_1020_375# net17 0.001134f
C3748 _437_/a_1308_423# net14 0.085815f
C3749 _448_/a_2248_156# vss 0.003807f
C3750 _448_/a_2665_112# vdd 0.005876f
C3751 _001_ cal_itt\[0\] 0.004843f
C3752 net15 FILLER_0_9_60/a_484_472# 0.020589f
C3753 FILLER_0_13_212/a_1468_375# _043_ 0.01418f
C3754 net69 net13 0.005834f
C3755 en net5 0.892091f
C3756 FILLER_0_8_138/a_124_375# _129_ 0.006506f
C3757 fanout72/a_36_113# net15 0.010284f
C3758 net79 _417_/a_36_151# 0.082646f
C3759 _079_ FILLER_0_3_172/a_1828_472# 0.001638f
C3760 FILLER_0_11_142/a_36_472# _076_ 0.003047f
C3761 fanout69/a_36_113# net74 0.034782f
C3762 net19 _044_ 0.138869f
C3763 FILLER_0_14_107/a_1380_472# vdd 0.002511f
C3764 cal_count\[3\] _070_ 0.059233f
C3765 FILLER_0_22_177/a_932_472# vss -0.001894f
C3766 FILLER_0_22_177/a_1380_472# vdd 0.007188f
C3767 _444_/a_36_151# net47 0.016691f
C3768 FILLER_0_4_152/a_124_375# vdd -0.001403f
C3769 _043_ FILLER_0_13_80/a_36_472# 0.016194f
C3770 FILLER_0_22_177/a_572_375# _435_/a_36_151# 0.059049f
C3771 _053_ _372_/a_2590_472# 0.001932f
C3772 _079_ net37 0.408392f
C3773 _120_ _172_ 0.010275f
C3774 net68 net49 0.607379f
C3775 cal_itt\[2\] FILLER_0_3_221/a_1380_472# 0.015024f
C3776 output27/a_224_472# FILLER_0_9_290/a_124_375# 0.02894f
C3777 _447_/a_2248_156# net69 0.001126f
C3778 output12/a_224_472# FILLER_0_0_198/a_36_472# 0.023414f
C3779 _077_ _061_ 0.031458f
C3780 _106_ output34/a_224_472# 0.01606f
C3781 _429_/a_36_151# FILLER_0_15_212/a_1020_375# 0.035849f
C3782 _267_/a_1568_472# _055_ 0.001681f
C3783 result[5] net77 0.142532f
C3784 _452_/a_1353_112# vdd 0.008539f
C3785 _448_/a_448_472# net76 0.003937f
C3786 _093_ net22 0.041918f
C3787 FILLER_0_4_49/a_124_375# _035_ 0.00215f
C3788 mask\[4\] _433_/a_2665_112# 0.005353f
C3789 net20 FILLER_0_12_220/a_932_472# 0.007397f
C3790 net52 FILLER_0_5_72/a_484_472# 0.050714f
C3791 net50 FILLER_0_5_72/a_1468_375# 0.001777f
C3792 _445_/a_2665_112# trim_mask\[1\] 0.00183f
C3793 mask\[0\] _429_/a_448_472# 0.061449f
C3794 FILLER_0_0_130/a_36_472# _442_/a_36_151# 0.001723f
C3795 _011_ _009_ 0.035129f
C3796 _276_/a_36_160# _092_ 0.06772f
C3797 _415_/a_2248_156# FILLER_0_11_282/a_124_375# 0.001221f
C3798 FILLER_0_16_73/a_36_472# net55 0.002576f
C3799 _048_ vss 0.056146f
C3800 FILLER_0_18_177/a_484_472# vss -0.001894f
C3801 FILLER_0_18_177/a_932_472# vdd 0.029926f
C3802 _189_/a_67_603# mask\[0\] 0.043158f
C3803 _140_ vdd 0.598538f
C3804 _070_ _169_ 0.006335f
C3805 FILLER_0_20_177/a_572_375# _098_ 0.015373f
C3806 _428_/a_2248_156# _131_ 0.005621f
C3807 _093_ FILLER_0_18_107/a_1380_472# 0.001782f
C3808 _398_/a_36_113# net44 0.011803f
C3809 _432_/a_36_151# net80 0.035794f
C3810 FILLER_0_5_128/a_572_375# vdd 0.008326f
C3811 _144_ FILLER_0_22_128/a_2812_375# 0.001601f
C3812 FILLER_0_9_60/a_484_472# net51 0.061362f
C3813 net27 output28/a_224_472# 0.011692f
C3814 net20 ctlp[1] 0.024556f
C3815 mask\[8\] net71 0.424276f
C3816 _431_/a_36_151# FILLER_0_16_115/a_124_375# 0.035117f
C3817 FILLER_0_5_206/a_124_375# net22 0.019537f
C3818 net20 _091_ 0.0557f
C3819 net75 _425_/a_1308_423# 0.034219f
C3820 _058_ net21 0.004383f
C3821 net41 _446_/a_2248_156# 0.016492f
C3822 _053_ FILLER_0_5_54/a_484_472# 0.001135f
C3823 FILLER_0_16_57/a_572_375# vss 0.00372f
C3824 FILLER_0_16_57/a_1020_375# vdd 0.004428f
C3825 _440_/a_36_151# FILLER_0_6_47/a_2724_472# 0.001653f
C3826 FILLER_0_6_37/a_124_375# _160_ 0.04948f
C3827 FILLER_0_3_2/a_36_472# _446_/a_36_151# 0.004032f
C3828 _439_/a_1308_423# FILLER_0_6_47/a_3260_375# 0.001224f
C3829 FILLER_0_12_28/a_36_472# vss 0.003004f
C3830 _114_ _428_/a_2248_156# 0.004516f
C3831 _012_ _098_ 0.002778f
C3832 FILLER_0_22_128/a_124_375# vdd 0.013058f
C3833 FILLER_0_5_128/a_124_375# net74 0.013683f
C3834 FILLER_0_22_86/a_1468_375# _211_/a_36_160# 0.010334f
C3835 ctln[6] net52 0.1064f
C3836 _415_/a_36_151# net18 0.015992f
C3837 _072_ _311_/a_3740_473# 0.005483f
C3838 FILLER_0_5_198/a_572_375# net21 0.023563f
C3839 _414_/a_448_472# cal_itt\[3\] 0.109704f
C3840 net71 vss 0.335256f
C3841 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_124_375# 0.009654f
C3842 fanout74/a_36_113# _371_/a_36_113# 0.01088f
C3843 net63 FILLER_0_20_177/a_572_375# 0.00281f
C3844 FILLER_0_17_56/a_572_375# FILLER_0_15_59/a_36_472# 0.001188f
C3845 _099_ _195_/a_255_603# 0.002146f
C3846 mask\[0\] FILLER_0_14_235/a_124_375# 0.009674f
C3847 cal_count\[3\] FILLER_0_11_78/a_572_375# 0.010243f
C3848 net47 FILLER_0_5_136/a_124_375# 0.010674f
C3849 FILLER_0_24_290/a_36_472# vdd 0.089567f
C3850 FILLER_0_24_290/a_124_375# vss 0.034103f
C3851 FILLER_0_5_172/a_124_375# vdd 0.028449f
C3852 vdd FILLER_0_13_290/a_36_472# 0.027484f
C3853 vss FILLER_0_13_290/a_124_375# 0.031844f
C3854 _426_/a_36_151# FILLER_0_9_270/a_36_472# 0.008172f
C3855 net16 cal_count\[0\] 0.152321f
C3856 _098_ FILLER_0_15_235/a_484_472# 0.004898f
C3857 FILLER_0_18_2/a_572_375# net38 0.007477f
C3858 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_36_472# 0.009654f
C3859 _128_ vdd 0.217501f
C3860 _098_ _438_/a_448_472# 0.008962f
C3861 cal_count\[3\] FILLER_0_12_50/a_36_472# 0.063276f
C3862 net81 net28 0.034606f
C3863 _073_ _081_ 0.046537f
C3864 _100_ net62 0.006742f
C3865 _363_/a_36_68# vdd 0.04306f
C3866 net75 _263_/a_224_472# 0.004396f
C3867 FILLER_0_6_47/a_2724_472# vdd 0.002467f
C3868 FILLER_0_6_47/a_2276_472# vss 0.004086f
C3869 output20/a_224_472# net78 0.001495f
C3870 _429_/a_1204_472# net22 0.001899f
C3871 net75 FILLER_0_8_247/a_572_375# 0.003962f
C3872 _093_ FILLER_0_17_72/a_3260_375# 0.011936f
C3873 FILLER_0_11_142/a_124_375# vss 0.008766f
C3874 FILLER_0_11_142/a_572_375# vdd 0.014107f
C3875 _149_ vdd 0.379674f
C3876 _104_ result[6] 0.096535f
C3877 output13/a_224_472# _037_ 0.019694f
C3878 ctln[6] _387_/a_36_113# 0.007687f
C3879 _425_/a_36_151# FILLER_0_8_247/a_484_472# 0.059367f
C3880 net81 _429_/a_1204_472# 0.005046f
C3881 _013_ vss 0.163674f
C3882 net27 FILLER_0_14_235/a_572_375# 0.006429f
C3883 FILLER_0_3_204/a_124_375# _088_ 0.00269f
C3884 net63 FILLER_0_19_171/a_1468_375# 0.006671f
C3885 net81 FILLER_0_10_247/a_124_375# 0.044906f
C3886 FILLER_0_12_236/a_124_375# vdd 0.005169f
C3887 output24/a_224_472# ctlp[7] 0.060657f
C3888 net33 _204_/a_67_603# 0.022193f
C3889 _418_/a_796_472# _007_ 0.012286f
C3890 net82 FILLER_0_3_221/a_1020_375# 0.010208f
C3891 result[6] _420_/a_36_151# 0.011901f
C3892 _132_ FILLER_0_15_116/a_36_472# 0.020589f
C3893 result[9] _103_ 0.034463f
C3894 FILLER_0_21_125/a_36_472# net54 0.016672f
C3895 _074_ FILLER_0_6_231/a_572_375# 0.009029f
C3896 net27 calibrate 0.017426f
C3897 mask\[0\] _056_ 0.001878f
C3898 _422_/a_2560_156# mask\[7\] 0.010664f
C3899 _390_/a_36_68# _171_ 0.001252f
C3900 FILLER_0_3_172/a_1916_375# net59 0.001221f
C3901 _074_ _056_ 0.002397f
C3902 _426_/a_36_151# _425_/a_1308_423# 0.001518f
C3903 _367_/a_36_68# vss 0.001589f
C3904 _066_ vss 0.08113f
C3905 net56 fanout54/a_36_160# 0.044466f
C3906 _341_/a_49_472# vdd 0.026636f
C3907 net61 vss 0.254538f
C3908 _102_ net19 0.011979f
C3909 state\[0\] vdd 0.120171f
C3910 net44 _054_ 0.003562f
C3911 _253_/a_36_68# _082_ 0.013108f
C3912 _126_ _428_/a_2248_156# 0.001131f
C3913 en_co_clk _095_ 0.003753f
C3914 FILLER_0_17_72/a_1020_375# net36 0.001777f
C3915 net15 FILLER_0_6_47/a_1380_472# 0.00464f
C3916 _130_ _428_/a_2248_156# 0.006602f
C3917 net44 cal_count\[2\] 0.191151f
C3918 net7 _446_/a_2248_156# 0.001166f
C3919 net57 FILLER_0_13_142/a_36_472# 0.011199f
C3920 _428_/a_796_472# _043_ 0.007935f
C3921 trim[0] vss 0.132654f
C3922 _322_/a_124_24# _125_ 0.01165f
C3923 FILLER_0_8_138/a_36_472# _077_ 0.005953f
C3924 _094_ net30 0.188507f
C3925 _430_/a_2665_112# net63 0.075661f
C3926 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_572_375# 0.086635f
C3927 FILLER_0_4_197/a_484_472# _088_ 0.014756f
C3928 _052_ _424_/a_1000_472# 0.007574f
C3929 FILLER_0_21_28/a_3260_375# vdd -0.001166f
C3930 FILLER_0_3_172/a_2276_472# vdd 0.00806f
C3931 net79 _418_/a_36_151# 0.059124f
C3932 FILLER_0_8_2/a_124_375# vss 0.003001f
C3933 FILLER_0_8_2/a_36_472# vdd 0.104141f
C3934 _449_/a_2665_112# en_co_clk 0.002966f
C3935 net17 net40 1.095167f
C3936 FILLER_0_13_212/a_36_472# mask\[0\] 0.001366f
C3937 fanout80/a_36_113# mask\[0\] 0.002212f
C3938 net4 FILLER_0_3_221/a_1380_472# 0.003953f
C3939 vss FILLER_0_8_156/a_484_472# 0.004078f
C3940 ctln[8] _447_/a_2665_112# 0.001271f
C3941 fanout82/a_36_113# output37/a_224_472# 0.023409f
C3942 trim_mask\[2\] net17 0.084388f
C3943 _117_ _310_/a_49_472# 0.018229f
C3944 _193_/a_36_160# _044_ 0.025719f
C3945 output33/a_224_472# _421_/a_2665_112# 0.010726f
C3946 result[6] _421_/a_1308_423# 0.023269f
C3947 net79 _138_ 0.024731f
C3948 net37 vss 0.666835f
C3949 _415_/a_36_151# net62 0.00514f
C3950 _176_ _390_/a_36_68# 0.005007f
C3951 FILLER_0_11_101/a_572_375# _120_ 0.006382f
C3952 _447_/a_1308_423# net17 0.002531f
C3953 net55 FILLER_0_17_72/a_1380_472# 0.021108f
C3954 _112_ _425_/a_448_472# 0.002335f
C3955 ctln[2] net58 0.025352f
C3956 _144_ _433_/a_1204_472# 0.009472f
C3957 fanout58/a_36_160# input4/a_36_68# 0.059453f
C3958 mask\[7\] _350_/a_49_472# 0.035293f
C3959 _057_ _128_ 0.036548f
C3960 _432_/a_2665_112# _136_ 0.002691f
C3961 FILLER_0_5_109/a_572_375# _153_ 0.03228f
C3962 FILLER_0_5_109/a_484_472# _154_ 0.039428f
C3963 _062_ _055_ 0.29425f
C3964 FILLER_0_17_64/a_124_375# vdd 0.027957f
C3965 _443_/a_2665_112# _170_ 0.019855f
C3966 _061_ _060_ 0.066418f
C3967 net76 FILLER_0_5_181/a_124_375# 0.031324f
C3968 _108_ vss 0.160825f
C3969 _132_ FILLER_0_17_104/a_1380_472# 0.02114f
C3970 _086_ _255_/a_224_552# 0.073601f
C3971 _131_ FILLER_0_17_104/a_484_472# 0.003483f
C3972 _176_ cal_count\[2\] 0.005783f
C3973 _059_ FILLER_0_5_136/a_36_472# 0.001755f
C3974 net36 mask\[2\] 0.871463f
C3975 _426_/a_36_151# FILLER_0_8_247/a_572_375# 0.059049f
C3976 output8/a_224_472# _000_ 0.182377f
C3977 _054_ _220_/a_67_603# 0.004333f
C3978 net1 _081_ 0.111227f
C3979 FILLER_0_8_37/a_484_472# _160_ 0.001767f
C3980 net56 FILLER_0_18_139/a_124_375# 0.00281f
C3981 _175_ FILLER_0_15_72/a_572_375# 0.04785f
C3982 _428_/a_36_151# FILLER_0_14_107/a_124_375# 0.001597f
C3983 net75 _317_/a_36_113# 0.030797f
C3984 _009_ net77 0.001183f
C3985 FILLER_0_21_206/a_124_375# _048_ 0.018458f
C3986 _098_ _113_ 0.001472f
C3987 FILLER_0_20_177/a_124_375# _434_/a_36_151# 0.059049f
C3988 _412_/a_2665_112# net18 0.001321f
C3989 _104_ mask\[4\] 0.001621f
C3990 net41 _043_ 0.03188f
C3991 FILLER_0_5_109/a_36_472# _163_ 0.00319f
C3992 FILLER_0_10_37/a_36_472# net68 0.005405f
C3993 _079_ _122_ 0.003853f
C3994 FILLER_0_0_266/a_124_375# vss 0.007654f
C3995 FILLER_0_0_266/a_36_472# vdd 0.05043f
C3996 _161_ _163_ 0.024512f
C3997 _042_ _039_ 0.003075f
C3998 net38 _452_/a_3129_107# 0.005269f
C3999 net57 net22 0.003595f
C4000 _179_ vss 0.089947f
C4001 FILLER_0_3_78/a_124_375# vdd 0.002419f
C4002 mask\[9\] FILLER_0_20_107/a_124_375# 0.004716f
C4003 _431_/a_2665_112# net73 0.001495f
C4004 FILLER_0_15_205/a_36_472# net22 0.037011f
C4005 FILLER_0_13_228/a_124_375# vdd -0.007362f
C4006 net53 FILLER_0_17_142/a_484_472# 0.001286f
C4007 cal_count\[3\] FILLER_0_12_28/a_124_375# 0.013328f
C4008 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_124_375# 0.001597f
C4009 FILLER_0_2_101/a_124_375# vdd 0.044073f
C4010 net41 _185_ 0.029318f
C4011 FILLER_0_4_107/a_1020_375# vdd 0.025121f
C4012 _114_ _267_/a_36_472# 0.011923f
C4013 net54 FILLER_0_18_107/a_36_472# 0.002116f
C4014 _103_ _418_/a_2560_156# 0.002179f
C4015 net70 FILLER_0_14_123/a_36_472# 0.009456f
C4016 _091_ _429_/a_2560_156# 0.001502f
C4017 net20 _418_/a_2248_156# 0.003507f
C4018 fanout78/a_36_113# net77 0.036366f
C4019 FILLER_0_5_117/a_36_472# FILLER_0_5_109/a_572_375# 0.086635f
C4020 net81 FILLER_0_15_205/a_36_472# 0.081574f
C4021 _026_ net71 0.406369f
C4022 cal net5 0.039735f
C4023 _293_/a_36_472# _106_ 0.04279f
C4024 net65 net8 0.203388f
C4025 FILLER_0_16_89/a_36_472# _177_ 0.048163f
C4026 net68 FILLER_0_8_37/a_36_472# 0.001088f
C4027 _435_/a_2248_156# mask\[6\] 0.001778f
C4028 result[4] _417_/a_2248_156# 0.001436f
C4029 _063_ vdd 0.201806f
C4030 _406_/a_36_159# _185_ 0.001573f
C4031 _079_ FILLER_0_6_231/a_484_472# 0.008159f
C4032 _448_/a_36_151# FILLER_0_2_177/a_124_375# 0.001597f
C4033 FILLER_0_4_185/a_124_375# net22 0.004776f
C4034 _179_ cal_count\[1\] 0.088667f
C4035 _028_ FILLER_0_6_47/a_3260_375# 0.013006f
C4036 _115_ trim_mask\[0\] 0.008966f
C4037 FILLER_0_9_28/a_2724_472# trim_val\[0\] 0.001183f
C4038 _139_ vdd 0.085044f
C4039 net65 _412_/a_1000_472# 0.00929f
C4040 result[8] vdd 0.590386f
C4041 net67 FILLER_0_6_37/a_124_375# 0.002918f
C4042 FILLER_0_7_195/a_36_472# _055_ 0.03271f
C4043 _449_/a_1308_423# _067_ 0.021042f
C4044 net15 FILLER_0_13_72/a_484_472# 0.002925f
C4045 _033_ _444_/a_1000_472# 0.00692f
C4046 _165_ _444_/a_2665_112# 0.044447f
C4047 _110_ mask\[8\] 0.05045f
C4048 _235_/a_67_603# net40 0.001273f
C4049 _053_ FILLER_0_6_47/a_1468_375# 0.008103f
C4050 net49 net47 0.53353f
C4051 _068_ _311_/a_2700_473# 0.001846f
C4052 _211_/a_36_160# net71 0.035804f
C4053 net76 FILLER_0_6_177/a_572_375# 0.073022f
C4054 _058_ _062_ 1.676625f
C4055 _140_ _433_/a_36_151# 0.020943f
C4056 _092_ vss 0.346097f
C4057 _235_/a_67_603# trim_mask\[2\] 0.022726f
C4058 _417_/a_1308_423# output30/a_224_472# 0.001434f
C4059 _370_/a_692_472# _081_ 0.00129f
C4060 _370_/a_848_380# _152_ 0.031499f
C4061 cal_count\[3\] _039_ 0.004827f
C4062 _177_ _176_ 0.226424f
C4063 net68 net47 0.063835f
C4064 _426_/a_36_151# _317_/a_36_113# 0.001082f
C4065 _070_ _120_ 0.838223f
C4066 FILLER_0_0_198/a_36_472# vss 0.00344f
C4067 cal_count\[3\] _373_/a_632_68# 0.004529f
C4068 en_co_clk vss 0.014954f
C4069 FILLER_0_15_150/a_124_375# fanout53/a_36_160# 0.004079f
C4070 FILLER_0_3_204/a_36_472# vss 0.003572f
C4071 _053_ _074_ 0.503728f
C4072 _140_ _147_ 0.08953f
C4073 _158_ vdd 0.131365f
C4074 cal_count\[2\] _183_ 0.034303f
C4075 _110_ vss 0.131865f
C4076 output29/a_224_472# FILLER_0_14_263/a_36_472# 0.0323f
C4077 net18 _419_/a_796_472# 0.006586f
C4078 trim_mask\[2\] _157_ 0.002951f
C4079 FILLER_0_1_192/a_36_472# net59 0.082738f
C4080 net57 _076_ 0.028356f
C4081 cal FILLER_0_1_266/a_572_375# 0.001707f
C4082 FILLER_0_19_47/a_36_472# _424_/a_448_472# 0.004782f
C4083 en_co_clk net74 0.039096f
C4084 fanout73/a_36_113# net36 0.01199f
C4085 net46 net17 0.791341f
C4086 net39 net40 0.279259f
C4087 _256_/a_244_497# _128_ 0.002372f
C4088 vss _416_/a_1000_472# 0.001784f
C4089 net27 FILLER_0_9_282/a_36_472# 0.002962f
C4090 result[0] FILLER_0_9_282/a_124_375# 0.00283f
C4091 net33 _023_ 0.015172f
C4092 net64 FILLER_0_14_235/a_36_472# 0.067888f
C4093 _119_ FILLER_0_8_156/a_484_472# 0.00979f
C4094 _423_/a_1308_423# vdd 0.00335f
C4095 _423_/a_448_472# vss 0.002481f
C4096 _064_ output39/a_224_472# 0.107406f
C4097 output34/a_224_472# net30 0.002189f
C4098 _414_/a_448_472# _081_ 0.024533f
C4099 net55 net15 1.200864f
C4100 output31/a_224_472# vss -0.003316f
C4101 _136_ FILLER_0_16_154/a_124_375# 0.00252f
C4102 FILLER_0_9_142/a_36_472# _120_ 0.035902f
C4103 _346_/a_49_472# vdd -0.002208f
C4104 fanout51/a_36_113# net55 0.010147f
C4105 _095_ _041_ 0.002104f
C4106 FILLER_0_4_197/a_1380_472# vdd 0.00581f
C4107 _432_/a_1000_472# vdd 0.010431f
C4108 net53 FILLER_0_14_99/a_124_375# 0.00494f
C4109 FILLER_0_17_161/a_124_375# vdd 0.014253f
C4110 net13 vss 0.071697f
C4111 _070_ FILLER_0_9_105/a_572_375# 0.017191f
C4112 FILLER_0_18_177/a_1380_472# _139_ 0.00195f
C4113 _104_ net34 0.293336f
C4114 FILLER_0_22_86/a_484_472# _098_ 0.003294f
C4115 FILLER_0_20_107/a_36_472# vss 0.004557f
C4116 _238_/a_67_603# _441_/a_2665_112# 0.015187f
C4117 _095_ _181_ 0.008117f
C4118 _424_/a_2248_156# vdd -0.005751f
C4119 _024_ _435_/a_36_151# 0.10993f
C4120 _098_ FILLER_0_19_111/a_124_375# 0.001331f
C4121 _027_ _438_/a_36_151# 0.010763f
C4122 _150_ _438_/a_1308_423# 0.001472f
C4123 _427_/a_36_151# net23 0.006844f
C4124 net69 _170_ 0.006468f
C4125 net55 _452_/a_3129_107# 0.006395f
C4126 _447_/a_2665_112# vdd 0.022038f
C4127 _447_/a_2248_156# vss 0.003961f
C4128 FILLER_0_18_2/a_1380_472# vss -0.001894f
C4129 FILLER_0_18_2/a_1828_472# vdd 0.001953f
C4130 net23 FILLER_0_5_148/a_572_375# 0.039975f
C4131 _274_/a_36_68# net27 0.027359f
C4132 net82 vdd 1.014512f
C4133 _114_ _113_ 0.201729f
C4134 _446_/a_1000_472# _035_ 0.00349f
C4135 FILLER_0_14_50/a_124_375# _179_ 0.021823f
C4136 FILLER_0_4_197/a_572_375# net76 0.006026f
C4137 _439_/a_2560_156# vss 0.001309f
C4138 net3 vdd 0.118499f
C4139 net17 trim[3] 0.001664f
C4140 _412_/a_2560_156# net58 0.005111f
C4141 fanout50/a_36_160# _168_ 0.033707f
C4142 net52 _384_/a_224_472# 0.001238f
C4143 _411_/a_1204_472# vss 0.001746f
C4144 _411_/a_2248_156# vdd 0.006283f
C4145 vdd FILLER_0_14_235/a_484_472# 0.010228f
C4146 vss FILLER_0_14_235/a_36_472# 0.001602f
C4147 FILLER_0_12_50/a_124_375# _067_ 0.011869f
C4148 FILLER_0_11_78/a_572_375# _120_ 0.01683f
C4149 _069_ FILLER_0_15_212/a_124_375# 0.039975f
C4150 _182_ _401_/a_36_68# 0.088487f
C4151 result[6] result[7] 0.119475f
C4152 net41 _402_/a_1296_93# 0.001707f
C4153 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_572_375# 0.001597f
C4154 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_36_472# 0.026657f
C4155 _070_ _227_/a_36_160# 0.00254f
C4156 net23 FILLER_0_19_155/a_124_375# 0.001347f
C4157 _131_ _118_ 0.001685f
C4158 _122_ vss 0.750387f
C4159 _436_/a_36_151# _140_ 0.031519f
C4160 _132_ FILLER_0_18_107/a_2724_472# 0.002229f
C4161 FILLER_0_4_99/a_36_472# net14 0.022408f
C4162 net55 net51 0.007067f
C4163 _436_/a_1308_423# output24/a_224_472# 0.005632f
C4164 fanout72/a_36_113# _067_ 0.005796f
C4165 output19/a_224_472# net19 0.030721f
C4166 FILLER_0_16_57/a_932_472# net55 0.00179f
C4167 net29 _196_/a_36_160# 0.073294f
C4168 FILLER_0_12_50/a_36_472# _120_ 0.005447f
C4169 FILLER_0_12_20/a_124_375# _039_ 0.004669f
C4170 _390_/a_244_472# _136_ 0.001777f
C4171 FILLER_0_13_212/a_124_375# FILLER_0_13_206/a_124_375# 0.005439f
C4172 net35 _435_/a_2248_156# 0.001854f
C4173 net44 FILLER_0_20_2/a_124_375# 0.001564f
C4174 _320_/a_1568_472# _043_ 0.00177f
C4175 _308_/a_848_380# _134_ 0.001299f
C4176 _132_ FILLER_0_16_107/a_36_472# 0.001538f
C4177 _114_ _118_ 0.074399f
C4178 FILLER_0_16_107/a_124_375# _131_ 0.016011f
C4179 input1/a_36_113# vss 0.05331f
C4180 fanout66/a_36_113# net49 0.001044f
C4181 FILLER_0_20_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001543f
C4182 mask\[5\] _205_/a_36_160# 0.003775f
C4183 FILLER_0_4_107/a_124_375# _154_ 0.00183f
C4184 FILLER_0_9_28/a_1828_472# net16 0.001946f
C4185 FILLER_0_19_142/a_36_472# _145_ 0.010377f
C4186 _049_ vss 0.026036f
C4187 net68 fanout66/a_36_113# 0.01746f
C4188 _115_ FILLER_0_10_94/a_572_375# 0.00887f
C4189 _408_/a_728_93# _186_ 0.003815f
C4190 FILLER_0_20_169/a_36_472# _339_/a_36_160# 0.001448f
C4191 fanout54/a_36_160# vss 0.061573f
C4192 _072_ _375_/a_692_497# 0.001113f
C4193 mask\[2\] FILLER_0_16_154/a_1468_375# 0.014254f
C4194 FILLER_0_13_142/a_1020_375# _043_ 0.005672f
C4195 net32 _421_/a_448_472# 0.022214f
C4196 FILLER_0_18_2/a_3172_472# _452_/a_36_151# 0.059367f
C4197 FILLER_0_18_2/a_2724_472# _452_/a_448_472# 0.008967f
C4198 net36 FILLER_0_15_212/a_1380_472# 0.006416f
C4199 _430_/a_1000_472# net21 0.053061f
C4200 FILLER_0_15_150/a_36_472# _136_ 0.002967f
C4201 FILLER_0_14_91/a_572_375# _176_ 0.002444f
C4202 _435_/a_2560_156# vdd 0.001372f
C4203 _435_/a_2665_112# vss 0.002665f
C4204 _436_/a_448_472# net71 0.005274f
C4205 net34 _210_/a_255_603# 0.002153f
C4206 _094_ _045_ 0.102437f
C4207 vss FILLER_0_6_231/a_484_472# 0.005629f
C4208 net17 FILLER_0_20_15/a_1020_375# 0.039975f
C4209 _061_ vss 0.046487f
C4210 _141_ _146_ 0.020044f
C4211 FILLER_0_24_63/a_124_375# output26/a_224_472# 0.00515f
C4212 FILLER_0_15_142/a_572_375# net56 0.001809f
C4213 _414_/a_796_472# _089_ 0.001426f
C4214 FILLER_0_15_205/a_124_375# vdd 0.015886f
C4215 FILLER_0_18_76/a_124_375# net71 0.008427f
C4216 trim_val\[1\] _034_ 0.001535f
C4217 net41 _033_ 0.033812f
C4218 FILLER_0_9_28/a_1380_472# vdd 0.01306f
C4219 _291_/a_36_160# _199_/a_36_160# 0.005575f
C4220 _428_/a_2665_112# _118_ 0.001007f
C4221 fanout70/a_36_113# _131_ 0.003364f
C4222 FILLER_0_14_263/a_124_375# net30 0.016642f
C4223 ctlp[1] FILLER_0_24_274/a_1020_375# 0.004803f
C4224 _451_/a_2225_156# _040_ 0.015815f
C4225 _098_ vdd 2.272938f
C4226 FILLER_0_12_2/a_572_375# _039_ 0.005407f
C4227 _286_/a_224_472# _005_ 0.001254f
C4228 net20 _199_/a_36_160# 0.05178f
C4229 trim_mask\[4\] _370_/a_124_24# 0.015021f
C4230 FILLER_0_3_54/a_124_375# _160_ 0.004602f
C4231 FILLER_0_17_56/a_572_375# vss 0.05884f
C4232 FILLER_0_17_56/a_36_472# vdd 0.040007f
C4233 output37/a_224_472# fanout65/a_36_113# 0.013171f
C4234 net23 FILLER_0_22_128/a_1916_375# 0.004205f
C4235 net52 FILLER_0_2_111/a_36_472# 0.0659f
C4236 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_36_472# 0.009654f
C4237 _372_/a_2034_472# _076_ 0.007461f
C4238 _372_/a_170_472# _068_ 0.037034f
C4239 _126_ _113_ 0.547055f
C4240 FILLER_0_21_28/a_572_375# FILLER_0_20_31/a_124_375# 0.026339f
C4241 _129_ _076_ 0.043637f
C4242 _132_ mask\[9\] 0.203851f
C4243 FILLER_0_13_212/a_932_472# vss 0.022933f
C4244 fanout65/a_36_113# net5 0.027955f
C4245 FILLER_0_17_72/a_36_472# _131_ 0.002672f
C4246 output19/a_224_472# _009_ 0.003174f
C4247 net82 net2 0.451147f
C4248 _425_/a_448_472# net19 0.034226f
C4249 _114_ _068_ 1.097353f
C4250 FILLER_0_4_177/a_484_472# _087_ 0.005486f
C4251 FILLER_0_4_152/a_124_375# net57 0.001947f
C4252 FILLER_0_17_226/a_36_472# vss 0.007552f
C4253 net38 FILLER_0_15_2/a_572_375# 0.007477f
C4254 FILLER_0_14_181/a_36_472# _138_ 0.002748f
C4255 FILLER_0_21_28/a_572_375# FILLER_0_19_28/a_484_472# 0.001512f
C4256 FILLER_0_6_239/a_36_472# fanout75/a_36_113# 0.00191f
C4257 FILLER_0_18_139/a_124_375# vss 0.006869f
C4258 FILLER_0_18_139/a_572_375# vdd 0.004039f
C4259 _086_ _395_/a_36_488# 0.00825f
C4260 _041_ vss 0.012963f
C4261 FILLER_0_5_206/a_36_472# net37 0.009858f
C4262 net63 vdd 1.002883f
C4263 net50 FILLER_0_6_79/a_36_472# 0.001614f
C4264 FILLER_0_24_130/a_124_375# ctlp[6] 0.021926f
C4265 _412_/a_448_472# _001_ 0.01124f
C4266 mask\[0\] net62 0.552008f
C4267 FILLER_0_11_109/a_124_375# FILLER_0_9_105/a_484_472# 0.0027f
C4268 result[7] FILLER_0_24_274/a_36_472# 0.006454f
C4269 _091_ FILLER_0_12_220/a_124_375# 0.006907f
C4270 _181_ vss 0.003673f
C4271 FILLER_0_0_130/a_124_375# _031_ 0.001861f
C4272 net42 net40 0.007686f
C4273 _037_ net22 0.079675f
C4274 mask\[7\] FILLER_0_22_128/a_2812_375# 0.001476f
C4275 mask\[5\] _009_ 0.001095f
C4276 _126_ _118_ 0.215385f
C4277 _130_ _118_ 0.053869f
C4278 _144_ FILLER_0_18_107/a_1916_375# 0.003148f
C4279 _253_/a_36_68# net19 0.019615f
C4280 FILLER_0_10_78/a_36_472# _439_/a_36_151# 0.00271f
C4281 _079_ net8 0.001928f
C4282 net80 FILLER_0_22_177/a_932_472# 0.002472f
C4283 net35 FILLER_0_22_128/a_2276_472# 0.014483f
C4284 net65 FILLER_0_3_221/a_1020_375# 0.001641f
C4285 _320_/a_36_472# state\[1\] 0.013058f
C4286 fanout68/a_36_113# vdd 0.012621f
C4287 _144_ mask\[4\] 0.268823f
C4288 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3172_472# 0.013276f
C4289 _053_ _312_/a_672_472# 0.001065f
C4290 net36 _451_/a_3129_107# 0.013154f
C4291 net20 _429_/a_448_472# 0.002244f
C4292 net68 FILLER_0_6_47/a_36_472# 0.001248f
C4293 _115_ FILLER_0_9_142/a_124_375# 0.010167f
C4294 FILLER_0_18_171/a_124_375# vss 0.048769f
C4295 FILLER_0_18_171/a_36_472# vdd 0.010704f
C4296 net64 FILLER_0_9_282/a_484_472# 0.005717f
C4297 trim_mask\[1\] FILLER_0_6_47/a_932_472# 0.007542f
C4298 output31/a_224_472# _103_ 0.006731f
C4299 net20 _189_/a_67_603# 0.011939f
C4300 _396_/a_224_472# _095_ 0.001351f
C4301 net67 FILLER_0_9_60/a_572_375# 0.011073f
C4302 net31 net61 0.053131f
C4303 cal_count\[3\] _228_/a_36_68# 0.01871f
C4304 FILLER_0_22_128/a_3172_472# vdd 0.003395f
C4305 FILLER_0_22_128/a_2724_472# vss 0.005195f
C4306 _108_ _295_/a_36_472# 0.014558f
C4307 _052_ FILLER_0_18_37/a_1468_375# 0.001585f
C4308 FILLER_0_7_72/a_2276_472# net14 0.004375f
C4309 result[9] FILLER_0_24_274/a_124_375# 0.008195f
C4310 _176_ FILLER_0_18_53/a_36_472# 0.001868f
C4311 _341_/a_49_472# FILLER_0_17_161/a_36_472# 0.079018f
C4312 _444_/a_2665_112# vss 0.002271f
C4313 _444_/a_2560_156# vdd 0.025035f
C4314 _181_ cal_count\[1\] 0.186904f
C4315 net70 FILLER_0_13_100/a_124_375# 0.017886f
C4316 _152_ _261_/a_36_160# 0.001102f
C4317 FILLER_0_9_28/a_36_472# net51 0.002082f
C4318 net16 _408_/a_1336_472# 0.022364f
C4319 _410_/a_36_68# _039_ 0.016062f
C4320 _072_ _074_ 2.017168f
C4321 FILLER_0_22_86/a_124_375# _437_/a_36_151# 0.001597f
C4322 _119_ _122_ 0.155432f
C4323 _086_ calibrate 0.041755f
C4324 FILLER_0_20_193/a_484_472# FILLER_0_18_177/a_2364_375# 0.0027f
C4325 _132_ _142_ 0.006253f
C4326 FILLER_0_5_72/a_1020_375# vdd 0.009501f
C4327 FILLER_0_5_72/a_572_375# vss 0.006023f
C4328 _452_/a_836_156# _041_ 0.001052f
C4329 _136_ _043_ 0.040107f
C4330 _394_/a_728_93# FILLER_0_13_72/a_484_472# 0.018997f
C4331 net26 FILLER_0_23_44/a_932_472# 0.001889f
C4332 _177_ FILLER_0_17_72/a_1468_375# 0.026469f
C4333 FILLER_0_12_236/a_572_375# FILLER_0_14_235/a_484_472# 0.001026f
C4334 net23 _163_ 0.034799f
C4335 _078_ net59 0.168928f
C4336 output38/a_224_472# net49 0.002434f
C4337 net38 net66 0.040578f
C4338 FILLER_0_21_28/a_2724_472# _424_/a_36_151# 0.001723f
C4339 FILLER_0_10_28/a_124_375# net17 0.00917f
C4340 net35 FILLER_0_22_107/a_484_472# 0.008026f
C4341 _413_/a_2665_112# net21 0.002828f
C4342 net4 _078_ 0.487587f
C4343 _126_ _068_ 0.01065f
C4344 net63 FILLER_0_18_177/a_1380_472# 0.070445f
C4345 FILLER_0_15_142/a_572_375# _095_ 0.003935f
C4346 net10 _411_/a_448_472# 0.010544f
C4347 _137_ _113_ 0.030279f
C4348 net38 _445_/a_1308_423# 0.006454f
C4349 trim[0] _445_/a_36_151# 0.008302f
C4350 net82 FILLER_0_3_172/a_2724_472# 0.007912f
C4351 trim_val\[1\] FILLER_0_6_37/a_124_375# 0.007292f
C4352 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_484_472# 0.001963f
C4353 _405_/a_67_603# vdd 0.034681f
C4354 FILLER_0_9_282/a_484_472# vss 0.00561f
C4355 net57 _128_ 0.040656f
C4356 _009_ _299_/a_36_472# 0.006927f
C4357 net41 FILLER_0_16_37/a_124_375# 0.008195f
C4358 _372_/a_170_472# vdd 0.031606f
C4359 FILLER_0_5_54/a_1468_375# _440_/a_36_151# 0.059049f
C4360 FILLER_0_8_138/a_36_472# vss 0.008189f
C4361 _094_ _418_/a_2665_112# 0.035668f
C4362 _131_ vdd 1.344823f
C4363 FILLER_0_15_116/a_124_375# _095_ 0.002659f
C4364 net52 _441_/a_36_151# 0.013755f
C4365 _028_ FILLER_0_7_72/a_1828_472# 0.001777f
C4366 _119_ _061_ 0.132725f
C4367 _120_ _039_ 0.148356f
C4368 net72 FILLER_0_20_31/a_124_375# 0.011347f
C4369 net58 result[0] 0.443436f
C4370 FILLER_0_12_124/a_36_472# FILLER_0_11_124/a_36_472# 0.05841f
C4371 fanout70/a_36_113# FILLER_0_15_116/a_572_375# 0.003553f
C4372 FILLER_0_5_128/a_124_375# _370_/a_124_24# 0.023285f
C4373 result[9] FILLER_0_23_274/a_124_375# 0.003102f
C4374 fanout63/a_36_160# FILLER_0_15_228/a_124_375# 0.001177f
C4375 FILLER_0_20_177/a_124_375# mask\[6\] 0.001158f
C4376 _136_ net21 0.022198f
C4377 output22/a_224_472# net23 0.008048f
C4378 net52 _440_/a_1000_472# 0.013793f
C4379 _287_/a_36_472# _094_ 0.029751f
C4380 FILLER_0_12_20/a_36_472# net6 0.007073f
C4381 _114_ vdd 1.30767f
C4382 ctln[2] net9 0.022757f
C4383 calibrate _169_ 0.001883f
C4384 output44/a_224_472# FILLER_0_18_2/a_124_375# 0.001168f
C4385 net38 _067_ 0.062447f
C4386 net72 _394_/a_718_524# 0.001558f
C4387 net55 _394_/a_728_93# 0.0026f
C4388 _053_ FILLER_0_7_72/a_36_472# 0.01287f
C4389 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_124_375# 0.009654f
C4390 FILLER_0_20_15/a_1380_472# vdd 0.007068f
C4391 mask\[4\] FILLER_0_18_177/a_2364_375# 0.01602f
C4392 net72 FILLER_0_19_28/a_484_472# 0.004312f
C4393 net55 FILLER_0_19_28/a_124_375# 0.002644f
C4394 _000_ FILLER_0_3_221/a_1380_472# 0.025567f
C4395 _123_ net37 0.002942f
C4396 mask\[4\] _339_/a_36_160# 0.003234f
C4397 _165_ FILLER_0_6_47/a_124_375# 0.014312f
C4398 _432_/a_1000_472# _093_ 0.007509f
C4399 _093_ FILLER_0_17_161/a_124_375# 0.002431f
C4400 _070_ net21 0.03068f
C4401 _239_/a_36_160# net40 0.010925f
C4402 net20 FILLER_0_6_231/a_572_375# 0.01215f
C4403 net69 FILLER_0_2_111/a_124_375# 0.010762f
C4404 FILLER_0_9_28/a_3260_375# fanout67/a_36_160# 0.001925f
C4405 net48 _251_/a_906_472# 0.001362f
C4406 _077_ _068_ 0.601166f
C4407 FILLER_0_12_20/a_484_472# net40 0.003391f
C4408 _178_ _402_/a_728_93# 0.050963f
C4409 _070_ FILLER_0_10_107/a_484_472# 0.007421f
C4410 _053_ net15 0.041871f
C4411 _127_ _121_ 0.023125f
C4412 en_co_clk _389_/a_36_148# 0.001249f
C4413 _428_/a_2665_112# vdd 0.004735f
C4414 cal en 0.482495f
C4415 _120_ FILLER_0_8_156/a_36_472# 0.005842f
C4416 _086_ _125_ 0.490983f
C4417 FILLER_0_5_54/a_1020_375# vss 0.003196f
C4418 FILLER_0_5_54/a_1468_375# vdd 0.014683f
C4419 _424_/a_36_151# FILLER_0_20_31/a_124_375# 0.012574f
C4420 _183_ FILLER_0_18_53/a_36_472# 0.007412f
C4421 FILLER_0_14_50/a_124_375# _181_ 0.00402f
C4422 _155_ FILLER_0_5_109/a_36_472# 0.001872f
C4423 _144_ net34 0.029247f
C4424 clk vdd 0.053789f
C4425 net29 FILLER_0_16_255/a_124_375# 0.085055f
C4426 FILLER_0_1_98/a_36_472# _153_ 0.001463f
C4427 net57 _386_/a_1084_68# 0.005716f
C4428 net58 output48/a_224_472# 0.065357f
C4429 net75 net48 0.10167f
C4430 _096_ _320_/a_36_472# 0.052438f
C4431 FILLER_0_4_177/a_36_472# vss 0.001806f
C4432 FILLER_0_4_177/a_484_472# vdd 0.010663f
C4433 _412_/a_2665_112# fanout59/a_36_160# 0.016426f
C4434 net73 FILLER_0_17_104/a_1468_375# 0.002342f
C4435 output28/a_224_472# result[1] 0.054333f
C4436 _415_/a_796_472# net19 0.001468f
C4437 FILLER_0_12_2/a_484_472# net6 0.005586f
C4438 _445_/a_2560_156# net17 0.010829f
C4439 _428_/a_2248_156# net74 0.072805f
C4440 _421_/a_448_472# _010_ 0.039422f
C4441 net69 fanout49/a_36_160# 0.005942f
C4442 ctln[1] FILLER_0_1_266/a_124_375# 0.002958f
C4443 _103_ _288_/a_224_472# 0.002992f
C4444 net55 FILLER_0_18_76/a_36_472# 0.003695f
C4445 _443_/a_2248_156# vss 0.008696f
C4446 _443_/a_2665_112# vdd 0.011824f
C4447 FILLER_0_19_125/a_124_375# FILLER_0_18_107/a_2276_472# 0.001684f
C4448 _369_/a_244_472# _160_ 0.00146f
C4449 trim_val\[4\] _163_ 0.03439f
C4450 net55 _423_/a_2248_156# 0.001188f
C4451 _253_/a_36_68# cal_itt\[0\] 0.001495f
C4452 FILLER_0_19_28/a_36_472# net40 0.020968f
C4453 net31 _092_ 0.04309f
C4454 FILLER_0_7_72/a_484_472# net52 0.049487f
C4455 output27/a_224_472# net27 0.046353f
C4456 net81 FILLER_0_15_212/a_124_375# 0.005049f
C4457 ctlp[6] vss 0.115894f
C4458 FILLER_0_14_50/a_36_472# _174_ 0.015387f
C4459 net70 FILLER_0_14_107/a_572_375# 0.018214f
C4460 _071_ _121_ 0.007734f
C4461 ctlp[5] _435_/a_36_151# 0.003815f
C4462 ctlp[3] output20/a_224_472# 0.023589f
C4463 net8 vss 0.171128f
C4464 FILLER_0_16_57/a_1468_375# _131_ 0.015859f
C4465 output25/a_224_472# net35 0.016177f
C4466 output46/a_224_472# FILLER_0_20_15/a_572_375# 0.00135f
C4467 _426_/a_2248_156# _060_ 0.00106f
C4468 _114_ _057_ 0.30288f
C4469 ctlp[4] vdd 0.278868f
C4470 net15 FILLER_0_15_72/a_36_472# 0.007185f
C4471 _174_ cal_count\[3\] 0.053844f
C4472 net16 FILLER_0_18_37/a_932_472# 0.008749f
C4473 net20 FILLER_0_16_241/a_124_375# 0.002327f
C4474 _098_ _433_/a_36_151# 0.023263f
C4475 _126_ vdd 0.682779f
C4476 net17 _450_/a_36_151# 0.006157f
C4477 _130_ vdd 0.046379f
C4478 cal_itt\[2\] _253_/a_244_68# 0.001073f
C4479 _004_ net58 0.00116f
C4480 net24 net14 0.172253f
C4481 _091_ FILLER_0_18_177/a_572_375# 0.004285f
C4482 _113_ _060_ 0.01991f
C4483 _190_/a_36_160# vdd 0.031799f
C4484 _140_ _434_/a_36_151# 0.025956f
C4485 _150_ vss 0.016993f
C4486 FILLER_0_5_206/a_36_472# _122_ 0.003017f
C4487 net34 FILLER_0_22_177/a_1020_375# 0.006974f
C4488 net36 FILLER_0_15_180/a_572_375# 0.002531f
C4489 result[2] vdd 0.18482f
C4490 _442_/a_36_151# _158_ 0.001257f
C4491 _256_/a_36_68# _058_ 0.001402f
C4492 FILLER_0_10_78/a_572_375# FILLER_0_9_72/a_1380_472# 0.001543f
C4493 ctlp[1] _419_/a_1204_472# 0.007338f
C4494 mask\[9\] _438_/a_36_151# 0.060632f
C4495 _170_ vss 0.280383f
C4496 FILLER_0_3_172/a_572_375# net22 0.013048f
C4497 FILLER_0_9_28/a_572_375# net41 0.025588f
C4498 FILLER_0_19_55/a_124_375# net55 0.005311f
C4499 net40 _160_ 0.152292f
C4500 FILLER_0_15_142/a_572_375# vss 0.095176f
C4501 FILLER_0_15_142/a_36_472# vdd 0.106034f
C4502 _056_ FILLER_0_12_196/a_124_375# 0.027077f
C4503 output31/a_224_472# net31 0.002146f
C4504 trim_val\[2\] _166_ 0.014514f
C4505 trim_mask\[2\] _160_ 0.367302f
C4506 _433_/a_2248_156# _145_ 0.009108f
C4507 _106_ mask\[3\] 0.249479f
C4508 FILLER_0_18_37/a_36_472# vss 0.003026f
C4509 FILLER_0_18_37/a_484_472# vdd 0.008381f
C4510 _093_ _098_ 0.556613f
C4511 net81 net27 1.118985f
C4512 FILLER_0_0_96/a_124_375# trim_mask\[3\] 0.006277f
C4513 FILLER_0_7_195/a_124_375# _072_ 0.012244f
C4514 ctln[4] net59 0.10527f
C4515 _322_/a_692_472# _070_ 0.002328f
C4516 output10/a_224_472# _411_/a_36_151# 0.001362f
C4517 _305_/a_36_159# net37 0.015682f
C4518 _128_ _129_ 0.029628f
C4519 _216_/a_255_603# net15 0.002146f
C4520 net76 FILLER_0_2_177/a_572_375# 0.053951f
C4521 FILLER_0_14_91/a_124_375# net53 0.065572f
C4522 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_124_375# 0.012222f
C4523 FILLER_0_15_116/a_572_375# vdd 0.017636f
C4524 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_572_375# 0.086635f
C4525 FILLER_0_6_90/a_484_472# net14 0.014785f
C4526 FILLER_0_15_142/a_572_375# net74 0.001652f
C4527 _227_/a_36_160# FILLER_0_8_156/a_36_472# 0.006647f
C4528 _132_ _086_ 0.014693f
C4529 _381_/a_244_68# _167_ 0.001153f
C4530 FILLER_0_10_78/a_1468_375# _308_/a_124_24# 0.001565f
C4531 _119_ FILLER_0_8_138/a_36_472# 0.003894f
C4532 FILLER_0_13_212/a_1380_472# FILLER_0_13_228/a_36_472# 0.013277f
C4533 FILLER_0_14_107/a_484_472# _043_ 0.001641f
C4534 net65 vdd 1.430654f
C4535 _448_/a_2665_112# _037_ 0.042225f
C4536 FILLER_0_23_88/a_124_375# _437_/a_36_151# 0.002709f
C4537 FILLER_0_4_144/a_36_472# trim_mask\[4\] 0.017557f
C4538 FILLER_0_9_223/a_572_375# _223_/a_36_160# 0.001177f
C4539 net55 _067_ 0.053438f
C4540 _427_/a_2248_156# net36 0.004462f
C4541 _115_ _127_ 0.042389f
C4542 _118_ _060_ 0.002868f
C4543 _132_ cal_count\[3\] 0.193553f
C4544 _030_ net40 0.002509f
C4545 _436_/a_796_472# _025_ 0.026852f
C4546 net15 _164_ 0.026132f
C4547 trim_mask\[2\] _030_ 1.467465f
C4548 result[7] _419_/a_2665_112# 0.002471f
C4549 _308_/a_124_24# FILLER_0_9_72/a_1380_472# 0.003595f
C4550 _077_ vdd 1.61568f
C4551 _178_ net17 0.115251f
C4552 net2 clk 0.046099f
C4553 _093_ FILLER_0_18_139/a_572_375# 0.008393f
C4554 FILLER_0_10_107/a_124_375# vdd 0.045066f
C4555 output47/a_224_472# net17 0.081437f
C4556 net63 _093_ 0.109689f
C4557 _445_/a_1000_472# net40 0.015508f
C4558 FILLER_0_12_136/a_572_375# _127_ 0.00116f
C4559 _447_/a_448_472# net68 0.012962f
C4560 net49 _440_/a_2560_156# 0.011378f
C4561 _064_ _445_/a_448_472# 0.080931f
C4562 FILLER_0_7_72/a_2364_375# _077_ 0.002969f
C4563 net79 FILLER_0_11_282/a_124_375# 0.002239f
C4564 _152_ _062_ 0.097086f
C4565 net64 FILLER_0_15_235/a_484_472# 0.005893f
C4566 result[5] _418_/a_448_472# 0.007308f
C4567 output32/a_224_472# _418_/a_2248_156# 0.024448f
C4568 FILLER_0_20_177/a_1020_375# vdd 0.005483f
C4569 net32 _419_/a_2560_156# 0.029586f
C4570 trim_mask\[4\] _031_ 0.001262f
C4571 net20 _046_ 0.194455f
C4572 _431_/a_1204_472# _020_ 0.002176f
C4573 _091_ FILLER_0_15_212/a_1468_375# 0.002531f
C4574 FILLER_0_15_235/a_484_472# mask\[1\] 0.014415f
C4575 trim[4] FILLER_0_8_2/a_36_472# 0.019134f
C4576 _116_ net4 0.00603f
C4577 _057_ _126_ 0.022413f
C4578 _028_ FILLER_0_6_90/a_36_472# 0.013106f
C4579 net22 mask\[6\] 0.612004f
C4580 _065_ net14 0.005438f
C4581 _088_ net22 0.17798f
C4582 FILLER_0_4_144/a_124_375# vdd 0.005512f
C4583 FILLER_0_17_104/a_932_472# vdd 0.020019f
C4584 _274_/a_36_68# FILLER_0_12_236/a_484_472# 0.001237f
C4585 _012_ vss 0.454371f
C4586 _328_/a_36_113# _428_/a_36_151# 0.030244f
C4587 FILLER_0_5_54/a_932_472# FILLER_0_6_47/a_1828_472# 0.026657f
C4588 _044_ net30 0.005104f
C4589 _050_ FILLER_0_22_107/a_572_375# 0.001825f
C4590 _095_ _113_ 0.004037f
C4591 net20 _015_ 0.005917f
C4592 ctlp[7] output25/a_224_472# 0.002088f
C4593 mask\[2\] FILLER_0_15_212/a_484_472# 0.001641f
C4594 net26 FILLER_0_21_28/a_1916_375# 0.008721f
C4595 _419_/a_448_472# vdd 0.022174f
C4596 _419_/a_36_151# vss -0.00139f
C4597 _136_ _451_/a_448_472# 0.047841f
C4598 _251_/a_244_472# net4 0.005273f
C4599 _277_/a_36_160# net30 0.014059f
C4600 _430_/a_2665_112# mask\[1\] 0.004574f
C4601 _413_/a_1204_472# _002_ 0.003057f
C4602 net39 _445_/a_2560_156# 0.003401f
C4603 _317_/a_36_113# FILLER_0_7_233/a_36_472# 0.003531f
C4604 net52 FILLER_0_9_72/a_1468_375# 0.003576f
C4605 _053_ _163_ 0.763235f
C4606 _267_/a_36_472# vss 0.001495f
C4607 _137_ vdd 0.945976f
C4608 FILLER_0_15_59/a_572_375# vss 0.018573f
C4609 FILLER_0_15_59/a_36_472# vdd 0.031071f
C4610 FILLER_0_21_286/a_484_472# net77 0.02147f
C4611 _217_/a_36_160# _052_ 0.016695f
C4612 _453_/a_36_151# vdd 0.164654f
C4613 net20 _274_/a_1612_497# 0.002057f
C4614 net54 net23 0.084191f
C4615 _414_/a_2560_156# _075_ 0.026328f
C4616 _320_/a_36_472# FILLER_0_13_206/a_36_472# 0.038251f
C4617 _131_ FILLER_0_17_64/a_36_472# 0.002638f
C4618 FILLER_0_19_171/a_36_472# vdd 0.004762f
C4619 FILLER_0_19_171/a_1468_375# vss 0.054352f
C4620 _238_/a_67_603# trim_val\[3\] 0.024283f
C4621 net69 vdd 1.102677f
C4622 net41 output41/a_224_472# 0.008587f
C4623 _272_/a_36_472# net37 0.002669f
C4624 FILLER_0_15_235/a_484_472# vss 0.003614f
C4625 _178_ FILLER_0_16_37/a_36_472# 0.007425f
C4626 _087_ _079_ 0.251042f
C4627 output45/a_224_472# net40 0.001284f
C4628 _242_/a_36_160# _066_ 0.044262f
C4629 net59 FILLER_0_3_212/a_124_375# 0.057221f
C4630 FILLER_0_24_96/a_124_375# net35 0.001886f
C4631 FILLER_0_17_282/a_36_472# _418_/a_1308_423# 0.001295f
C4632 _122_ _123_ 0.242965f
C4633 _438_/a_448_472# vss 0.00615f
C4634 _055_ _223_/a_36_160# 0.012271f
C4635 output46/a_224_472# net44 0.003804f
C4636 FILLER_0_4_152/a_124_375# FILLER_0_4_144/a_572_375# 0.012001f
C4637 _011_ _422_/a_36_151# 0.015698f
C4638 net4 FILLER_0_3_212/a_124_375# 0.001739f
C4639 FILLER_0_17_72/a_2364_375# _451_/a_448_472# 0.001512f
C4640 net5 rstn 0.101356f
C4641 _360_/a_36_160# FILLER_0_4_123/a_124_375# 0.013555f
C4642 net57 net82 0.91473f
C4643 _077_ _057_ 0.584179f
C4644 cal_count\[2\] _401_/a_36_68# 0.008136f
C4645 trim_mask\[4\] _371_/a_36_113# 0.007529f
C4646 _032_ _159_ 0.053405f
C4647 _415_/a_2665_112# fanout62/a_36_160# 0.016426f
C4648 cal_count\[1\] FILLER_0_15_59/a_572_375# 0.008797f
C4649 FILLER_0_9_28/a_2364_375# net68 0.019969f
C4650 _086_ _069_ 0.580351f
C4651 net73 FILLER_0_18_107/a_932_472# 0.016711f
C4652 FILLER_0_19_125/a_36_472# vdd 0.003414f
C4653 FILLER_0_19_125/a_124_375# vss 0.001974f
C4654 net16 _450_/a_3129_107# 0.064714f
C4655 net65 net2 0.035908f
C4656 _070_ _062_ 0.06973f
C4657 FILLER_0_24_96/a_36_472# vss 0.003218f
C4658 _430_/a_2665_112# vss 0.031646f
C4659 _432_/a_796_472# net80 0.007731f
C4660 calibrate _120_ 0.001106f
C4661 _171_ net14 0.020479f
C4662 output26/a_224_472# FILLER_0_23_44/a_36_472# 0.026108f
C4663 _126_ FILLER_0_11_142/a_36_472# 0.001428f
C4664 _141_ _433_/a_2665_112# 0.013144f
C4665 _093_ _131_ 0.254316f
C4666 _069_ cal_count\[3\] 0.012382f
C4667 _242_/a_36_160# net37 0.02401f
C4668 FILLER_0_4_177/a_124_375# _163_ 0.004052f
C4669 net47 _385_/a_36_68# 0.011168f
C4670 net54 _025_ 0.00573f
C4671 net32 _105_ 2.08459f
C4672 FILLER_0_6_47/a_572_375# vdd 0.003158f
C4673 _043_ _039_ 0.001161f
C4674 trim_val\[3\] net15 0.068273f
C4675 _123_ FILLER_0_6_231/a_484_472# 0.001396f
C4676 cal_itt\[3\] _078_ 0.024443f
C4677 _164_ _381_/a_36_472# 0.007224f
C4678 net20 net18 0.025322f
C4679 _426_/a_2248_156# net64 0.01109f
C4680 _420_/a_2665_112# vdd 0.024431f
C4681 _420_/a_2248_156# vss -0.001f
C4682 net10 FILLER_0_1_212/a_124_375# 0.002314f
C4683 _121_ net23 0.078786f
C4684 FILLER_0_7_72/a_124_375# FILLER_0_6_47/a_2812_375# 0.026339f
C4685 net53 _451_/a_1353_112# 0.028324f
C4686 _263_/a_224_472# net59 0.002558f
C4687 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_484_472# 0.013276f
C4688 _013_ FILLER_0_18_37/a_1380_472# 0.01384f
C4689 net19 _419_/a_2248_156# 0.012726f
C4690 FILLER_0_17_104/a_124_375# net14 0.010099f
C4691 _061_ _311_/a_3740_473# 0.006728f
C4692 mask\[1\] _113_ 0.032744f
C4693 output12/a_224_472# vdd 0.106635f
C4694 fanout70/a_36_113# _095_ 0.003087f
C4695 _431_/a_2248_156# FILLER_0_18_139/a_932_472# 0.001148f
C4696 _176_ net14 0.031922f
C4697 _449_/a_2560_156# _038_ 0.010532f
C4698 trim[0] FILLER_0_3_2/a_36_472# 0.017429f
C4699 net56 vdd 0.277166f
C4700 FILLER_0_13_142/a_484_472# vss 0.024835f
C4701 _392_/a_36_68# _067_ 0.020085f
C4702 FILLER_0_16_57/a_484_472# FILLER_0_15_59/a_124_375# 0.001543f
C4703 _413_/a_36_151# FILLER_0_4_197/a_36_472# 0.001512f
C4704 FILLER_0_17_72/a_1828_472# _136_ 0.004161f
C4705 FILLER_0_7_59/a_484_472# net68 0.002785f
C4706 _213_/a_67_603# vdd 0.014901f
C4707 FILLER_0_1_266/a_572_375# rstn 0.00328f
C4708 fanout69/a_36_113# _371_/a_36_113# 0.259508f
C4709 FILLER_0_16_73/a_124_375# vdd 0.008987f
C4710 FILLER_0_18_107/a_124_375# FILLER_0_20_107/a_36_472# 0.00108f
C4711 _360_/a_36_160# _163_ 0.008593f
C4712 _177_ _451_/a_2225_156# 0.031347f
C4713 _248_/a_36_68# vdd 0.038887f
C4714 _430_/a_36_151# _337_/a_49_472# 0.023882f
C4715 net74 FILLER_0_13_142/a_484_472# 0.001771f
C4716 trim_mask\[2\] _156_ 0.018332f
C4717 _077_ cal_count\[0\] 0.018501f
C4718 FILLER_0_3_172/a_124_375# vdd 0.010886f
C4719 _116_ net79 0.081785f
C4720 _276_/a_36_160# vdd 0.010213f
C4721 ctln[5] _448_/a_796_472# 0.001484f
C4722 FILLER_0_1_266/a_124_375# net19 0.007016f
C4723 _422_/a_1000_472# vdd 0.005284f
C4724 _163_ _164_ 0.021311f
C4725 _165_ vdd 0.168803f
C4726 net7 output41/a_224_472# 0.019483f
C4727 net57 _098_ 0.062604f
C4728 trim_mask\[4\] FILLER_0_2_111/a_1468_375# 0.001226f
C4729 _177_ fanout55/a_36_160# 0.002687f
C4730 _426_/a_2248_156# vss 0.002303f
C4731 _426_/a_2665_112# vdd 0.008893f
C4732 net67 net40 0.886781f
C4733 _098_ FILLER_0_15_205/a_36_472# 0.010528f
C4734 _265_/a_224_472# net59 0.001052f
C4735 FILLER_0_10_78/a_572_375# _176_ 0.005927f
C4736 net26 net55 0.002901f
C4737 FILLER_0_5_117/a_124_375# _360_/a_36_160# 0.004736f
C4738 FILLER_0_15_282/a_484_472# vss 0.005507f
C4739 _446_/a_36_151# net66 0.034846f
C4740 _060_ vdd 0.349556f
C4741 FILLER_0_24_96/a_124_375# ctlp[7] 0.004486f
C4742 _113_ vss 0.147905f
C4743 _064_ _446_/a_2248_156# 0.04774f
C4744 trimb[4] vdd 0.081023f
C4745 net20 fanout75/a_36_113# 0.001027f
C4746 _112_ _316_/a_692_472# 0.001614f
C4747 net35 net22 0.001381f
C4748 fanout50/a_36_160# _383_/a_36_472# 0.096296f
C4749 FILLER_0_3_221/a_1020_375# vss 0.003948f
C4750 FILLER_0_3_221/a_1468_375# vdd 0.008815f
C4751 _125_ _120_ 0.006198f
C4752 _102_ net30 0.043037f
C4753 FILLER_0_4_49/a_484_472# _164_ 0.003258f
C4754 _236_/a_36_160# FILLER_0_8_2/a_36_472# 0.01395f
C4755 net65 FILLER_0_3_172/a_2724_472# 0.001777f
C4756 FILLER_0_5_72/a_572_375# _029_ 0.010208f
C4757 fanout63/a_36_160# net36 0.004435f
C4758 ctln[8] ctln[9] 0.003265f
C4759 _413_/a_1308_423# net59 0.018948f
C4760 sample result[0] 0.081581f
C4761 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1468_375# 0.086635f
C4762 _321_/a_170_472# _126_ 0.018831f
C4763 net12 vdd 0.082923f
C4764 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_124_375# 0.003732f
C4765 net16 _052_ 0.022236f
C4766 _431_/a_36_151# _136_ 0.03371f
C4767 _130_ _321_/a_170_472# 0.001018f
C4768 net63 FILLER_0_15_205/a_36_472# 0.047903f
C4769 _048_ _204_/a_67_603# 0.004547f
C4770 _372_/a_3662_472# net23 0.002864f
C4771 FILLER_0_2_111/a_572_375# vdd 0.012666f
C4772 FILLER_0_8_24/a_484_472# net40 0.004383f
C4773 net20 net62 0.058892f
C4774 output45/a_224_472# net46 0.005906f
C4775 net34 output35/a_224_472# 0.0731f
C4776 _330_/a_224_472# vdd 0.001701f
C4777 FILLER_0_4_99/a_36_472# net47 0.003903f
C4778 _144_ _146_ 0.333799f
C4779 _004_ _192_/a_67_603# 0.020219f
C4780 FILLER_0_18_2/a_36_472# cal_count\[2\] 0.001929f
C4781 _081_ FILLER_0_5_148/a_484_472# 0.016132f
C4782 _118_ vss 0.217218f
C4783 net26 _424_/a_796_472# 0.006496f
C4784 _057_ net56 0.002158f
C4785 _174_ _120_ 0.002521f
C4786 FILLER_0_18_107/a_2276_472# vdd 0.004405f
C4787 ctln[8] vss 0.351742f
C4788 _115_ net23 0.018953f
C4789 net78 _419_/a_448_472# 0.0122f
C4790 net60 _419_/a_448_472# 0.05959f
C4791 net61 _419_/a_796_472# 0.00438f
C4792 fanout69/a_36_113# FILLER_0_2_111/a_1468_375# 0.015816f
C4793 FILLER_0_24_130/a_124_375# vdd 0.027763f
C4794 _341_/a_257_69# _137_ 0.004351f
C4795 _322_/a_124_24# _128_ 0.02077f
C4796 net54 FILLER_0_22_128/a_1828_472# 0.009504f
C4797 net73 fanout71/a_36_113# 0.004833f
C4798 FILLER_0_16_89/a_932_472# _040_ 0.00702f
C4799 _417_/a_1204_472# _006_ 0.014354f
C4800 _058_ FILLER_0_9_105/a_484_472# 0.00148f
C4801 _087_ vss 0.09895f
C4802 _079_ vdd 0.476075f
C4803 net74 _118_ 0.060991f
C4804 _112_ net76 0.011948f
C4805 FILLER_0_16_107/a_572_375# vdd 0.019922f
C4806 FILLER_0_16_107/a_124_375# vss 0.002683f
C4807 _397_/a_36_472# net36 0.010045f
C4808 _198_/a_67_603# net30 0.017304f
C4809 net41 FILLER_0_19_28/a_572_375# 0.040551f
C4810 FILLER_0_6_79/a_124_375# vdd 0.015119f
C4811 FILLER_0_12_136/a_572_375# net23 0.00281f
C4812 fanout49/a_36_160# vss 0.025717f
C4813 FILLER_0_16_73/a_124_375# FILLER_0_16_57/a_1468_375# 0.012222f
C4814 net5 cal_itt\[1\] 0.057623f
C4815 _115_ _439_/a_2248_156# 0.003553f
C4816 ctln[4] FILLER_0_1_212/a_124_375# 0.008197f
C4817 FILLER_0_10_78/a_1380_472# _120_ 0.003228f
C4818 output37/a_224_472# valid 0.039402f
C4819 _315_/a_1229_68# _121_ 0.003401f
C4820 _414_/a_2560_156# net22 0.00603f
C4821 _057_ _060_ 0.033334f
C4822 net55 FILLER_0_17_38/a_36_472# 0.010728f
C4823 cal_count\[2\] FILLER_0_15_10/a_124_375# 0.017594f
C4824 ctlp[3] result[8] 0.278543f
C4825 FILLER_0_18_171/a_124_375# net80 0.024341f
C4826 _095_ vdd 1.051346f
C4827 FILLER_0_13_65/a_124_375# _095_ 0.002035f
C4828 mask\[3\] net30 0.451388f
C4829 net10 _000_ 0.001954f
C4830 valid net5 0.044555f
C4831 net4 FILLER_0_12_220/a_1020_375# 0.020782f
C4832 FILLER_0_8_107/a_124_375# vdd 0.049132f
C4833 _004_ FILLER_0_10_256/a_36_472# 0.00402f
C4834 net66 FILLER_0_5_54/a_124_375# 0.002093f
C4835 _096_ state\[1\] 0.083332f
C4836 FILLER_0_7_104/a_572_375# _058_ 0.006125f
C4837 FILLER_0_22_177/a_1380_472# mask\[6\] 0.006573f
C4838 FILLER_0_17_64/a_124_375# FILLER_0_15_59/a_484_472# 0.001188f
C4839 _450_/a_2449_156# _039_ 0.013285f
C4840 _132_ _120_ 0.034714f
C4841 fanout71/a_36_113# FILLER_0_19_111/a_484_472# 0.007864f
C4842 _431_/a_448_472# net53 0.002087f
C4843 net18 _416_/a_1288_156# 0.001147f
C4844 FILLER_0_8_138/a_124_375# _120_ 0.12254f
C4845 _072_ _163_ 0.016226f
C4846 net54 FILLER_0_22_107/a_36_472# 0.043792f
C4847 _068_ vss 0.547532f
C4848 FILLER_0_5_54/a_1020_375# _029_ 0.024737f
C4849 _449_/a_2248_156# vss 0.008071f
C4850 _449_/a_2665_112# vdd 0.012848f
C4851 _440_/a_2560_156# net47 0.003888f
C4852 net35 FILLER_0_22_86/a_36_472# 0.00797f
C4853 mask\[8\] FILLER_0_22_86/a_484_472# 0.012439f
C4854 fanout70/a_36_113# net74 0.002663f
C4855 net52 _442_/a_1000_472# 0.016308f
C4856 _114_ _311_/a_3220_473# 0.003283f
C4857 result[4] net18 0.048179f
C4858 FILLER_0_17_72/a_36_472# vss 0.036865f
C4859 net57 _131_ 0.030577f
C4860 FILLER_0_16_89/a_484_472# net36 0.003595f
C4861 net60 _420_/a_2665_112# 0.038894f
C4862 net78 _420_/a_2665_112# 0.039469f
C4863 net52 trim_mask\[1\] 0.04149f
C4864 _093_ FILLER_0_17_104/a_932_472# 0.014431f
C4865 _255_/a_224_552# _062_ 0.009032f
C4866 result[2] _416_/a_2248_156# 0.001396f
C4867 _449_/a_2248_156# net74 0.004565f
C4868 _186_ _180_ 0.003034f
C4869 trimb[1] FILLER_0_18_2/a_932_472# 0.011513f
C4870 net65 output11/a_224_472# 0.001529f
C4871 _083_ _082_ 0.018442f
C4872 output9/a_224_472# ctln[2] 0.080206f
C4873 FILLER_0_22_86/a_932_472# vdd 0.001826f
C4874 _122_ _242_/a_36_160# 0.005377f
C4875 _113_ _279_/a_652_68# 0.001425f
C4876 _192_/a_67_603# _044_ 0.002571f
C4877 net38 _450_/a_1284_156# 0.001291f
C4878 _131_ _135_ 0.068855f
C4879 _131_ FILLER_0_17_56/a_484_472# 0.002672f
C4880 cal_itt\[3\] _116_ 0.001364f
C4881 _093_ _137_ 0.201779f
C4882 _114_ net57 0.22998f
C4883 _140_ mask\[6\] 0.605898f
C4884 FILLER_0_19_111/a_572_375# vdd -0.008314f
C4885 _432_/a_2560_156# _136_ 0.001178f
C4886 FILLER_0_19_187/a_124_375# vdd 0.030349f
C4887 output15/a_224_472# net14 0.003312f
C4888 FILLER_0_0_198/a_124_375# net21 0.004256f
C4889 _065_ net49 0.001576f
C4890 _086_ _090_ 0.065807f
C4891 _449_/a_1000_472# net15 0.056791f
C4892 net69 FILLER_0_3_78/a_572_375# 0.002984f
C4893 net14 FILLER_0_10_94/a_124_375# 0.007086f
C4894 FILLER_0_3_204/a_124_375# net21 0.010054f
C4895 net27 FILLER_0_12_236/a_124_375# 0.044776f
C4896 FILLER_0_13_212/a_1468_375# FILLER_0_12_220/a_572_375# 0.05841f
C4897 net34 mask\[7\] 0.901671f
C4898 FILLER_0_19_125/a_36_472# _433_/a_36_151# 0.059367f
C4899 _065_ net68 0.194392f
C4900 net69 FILLER_0_2_101/a_36_472# 0.00845f
C4901 _114_ _135_ 0.018715f
C4902 _003_ net76 0.080782f
C4903 FILLER_0_19_55/a_36_472# _216_/a_67_603# 0.00254f
C4904 _411_/a_2560_156# net8 0.013106f
C4905 _408_/a_728_93# _181_ 0.018292f
C4906 FILLER_0_4_123/a_36_472# _152_ 0.003937f
C4907 _074_ net37 0.064705f
C4908 FILLER_0_11_101/a_484_472# cal_count\[3\] 0.00702f
C4909 _093_ _438_/a_1308_423# 0.001057f
C4910 _176_ _394_/a_718_524# 0.00141f
C4911 cal_count\[3\] _090_ 0.243462f
C4912 net60 _421_/a_1288_156# 0.001147f
C4913 _098_ _434_/a_36_151# 0.019342f
C4914 net66 _164_ 0.093385f
C4915 _444_/a_796_472# net67 0.006859f
C4916 net53 _427_/a_1308_423# 0.007426f
C4917 FILLER_0_12_236/a_572_375# _060_ 0.001597f
C4918 net57 _428_/a_2665_112# 0.027291f
C4919 _407_/a_36_472# _184_ 0.004667f
C4920 net61 _422_/a_2248_156# 0.027973f
C4921 _086_ net22 0.00117f
C4922 _231_/a_652_68# _062_ 0.001555f
C4923 _057_ _095_ 0.001346f
C4924 _083_ _265_/a_244_68# 0.004022f
C4925 net64 vdd 1.155692f
C4926 _440_/a_448_472# vdd 0.007263f
C4927 _440_/a_36_151# vss 0.016458f
C4928 mask\[1\] vdd 0.741266f
C4929 _078_ _081_ 0.445443f
C4930 _028_ FILLER_0_7_104/a_36_472# 0.006408f
C4931 net75 FILLER_0_8_263/a_36_472# 0.020293f
C4932 net34 _435_/a_796_472# 0.002288f
C4933 FILLER_0_4_197/a_484_472# net21 0.046864f
C4934 FILLER_0_6_239/a_36_472# net37 0.004187f
C4935 output23/a_224_472# _208_/a_36_160# 0.014541f
C4936 vdd FILLER_0_4_91/a_484_472# 0.007304f
C4937 _112_ _083_ 0.003571f
C4938 FILLER_0_7_162/a_124_375# net47 0.030995f
C4939 _119_ _118_ 0.001596f
C4940 mask\[9\] _140_ 0.00126f
C4941 net1 net18 0.047886f
C4942 FILLER_0_21_206/a_36_472# net22 0.012952f
C4943 net63 _434_/a_36_151# 0.005153f
C4944 _053_ FILLER_0_7_104/a_124_375# 0.012564f
C4945 _152_ _153_ 0.002954f
C4946 _444_/a_1000_472# _054_ 0.002998f
C4947 net81 FILLER_0_12_236/a_484_472# 0.001419f
C4948 ctln[9] vdd 0.221231f
C4949 _228_/a_36_68# net21 0.055313f
C4950 FILLER_0_12_20/a_36_472# _450_/a_448_472# 0.058631f
C4951 FILLER_0_17_142/a_124_375# _137_ 0.006974f
C4952 mask\[8\] vdd 0.423606f
C4953 net73 net71 0.033964f
C4954 _429_/a_2560_156# net62 0.002164f
C4955 _069_ _120_ 0.030804f
C4956 FILLER_0_12_2/a_124_375# vss 0.002871f
C4957 _423_/a_1000_472# _012_ 0.013415f
C4958 _422_/a_2248_156# _108_ 0.019477f
C4959 _430_/a_796_472# net36 0.00117f
C4960 _412_/a_1308_423# net1 0.022273f
C4961 FILLER_0_18_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001684f
C4962 result[4] net62 0.050684f
C4963 FILLER_0_14_81/a_124_375# vdd 0.023163f
C4964 FILLER_0_21_286/a_124_375# _420_/a_36_151# 0.001597f
C4965 net57 _126_ 0.021705f
C4966 _093_ net56 0.040124f
C4967 FILLER_0_22_86/a_124_375# net14 0.003962f
C4968 net19 _006_ 0.090449f
C4969 ctln[4] _000_ 0.002823f
C4970 net79 FILLER_0_12_220/a_1020_375# 0.010818f
C4971 vdd vss 15.42941f
C4972 FILLER_0_13_65/a_36_472# vdd 0.005885f
C4973 FILLER_0_13_65/a_124_375# vss 0.030194f
C4974 _448_/a_36_151# net59 0.062656f
C4975 output42/a_224_472# _054_ 0.013225f
C4976 _053_ _414_/a_448_472# 0.065053f
C4977 fanout67/a_36_160# trim_val\[0\] 0.003096f
C4978 calibrate net21 0.036773f
C4979 fanout51/a_36_113# FILLER_0_11_78/a_36_472# 0.193759f
C4980 _143_ mask\[3\] 0.023322f
C4981 mask\[7\] FILLER_0_22_177/a_124_375# 0.001315f
C4982 _424_/a_2560_156# _012_ 0.002513f
C4983 _106_ output18/a_224_472# 0.005393f
C4984 FILLER_0_7_72/a_2812_375# vdd 0.02125f
C4985 output37/a_224_472# net59 0.001014f
C4986 cal_count\[3\] _038_ 0.682941f
C4987 _126_ _135_ 0.011447f
C4988 output23/a_224_472# _210_/a_67_603# 0.021084f
C4989 _432_/a_1204_472# _137_ 0.006554f
C4990 FILLER_0_17_161/a_36_472# _137_ 0.013985f
C4991 FILLER_0_18_76/a_572_375# _438_/a_36_151# 0.059049f
C4992 net35 FILLER_0_22_177/a_1380_472# 0.01447f
C4993 _276_/a_36_160# _093_ 0.019339f
C4994 net74 vdd 1.451847f
C4995 FILLER_0_13_65/a_124_375# net74 0.020091f
C4996 _017_ net14 0.014743f
C4997 _095_ cal_count\[0\] 0.005211f
C4998 result[6] FILLER_0_21_286/a_36_472# 0.015369f
C4999 mask\[5\] FILLER_0_19_171/a_124_375# 0.002206f
C5000 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1468_375# 0.086635f
C5001 net38 net17 1.634286f
C5002 net71 FILLER_0_19_111/a_484_472# 0.004544f
C5003 _052_ FILLER_0_21_28/a_3260_375# 0.002388f
C5004 _119_ _068_ 0.040944f
C5005 _086_ _076_ 0.79237f
C5006 net5 net59 0.923076f
C5007 FILLER_0_10_78/a_932_472# _115_ 0.013773f
C5008 fanout75/a_36_113# net1 0.011428f
C5009 FILLER_0_11_64/a_124_375# _453_/a_2248_156# 0.001901f
C5010 _437_/a_1000_472# net14 0.028506f
C5011 FILLER_0_13_212/a_484_472# _043_ 0.011439f
C5012 _129_ _372_/a_170_472# 0.001985f
C5013 net4 net5 0.104296f
C5014 net68 _220_/a_67_603# 0.030878f
C5015 _131_ _129_ 0.017222f
C5016 _088_ FILLER_0_3_172/a_2276_472# 0.024532f
C5017 _435_/a_2248_156# net21 0.012406f
C5018 FILLER_0_17_38/a_124_375# _041_ 0.009172f
C5019 cal_count\[1\] vdd 0.516859f
C5020 mask\[9\] _149_ 0.040342f
C5021 _444_/a_1308_423# net47 0.040252f
C5022 FILLER_0_4_152/a_36_472# vss 0.009467f
C5023 FILLER_0_22_177/a_1468_375# _435_/a_36_151# 0.059049f
C5024 _053_ _372_/a_3662_472# 0.002006f
C5025 output13/a_224_472# ctln[6] 0.080817f
C5026 _442_/a_36_151# net69 0.048683f
C5027 _036_ net49 0.005235f
C5028 _447_/a_2560_156# net69 0.001774f
C5029 _445_/a_2665_112# net49 0.03968f
C5030 _053_ _155_ 0.122798f
C5031 net58 FILLER_0_9_270/a_572_375# 0.006256f
C5032 _077_ net57 0.025864f
C5033 net68 _036_ 0.168017f
C5034 _429_/a_36_151# FILLER_0_15_212/a_36_472# 0.001723f
C5035 result[5] _007_ 0.0249f
C5036 net35 _140_ 0.12583f
C5037 _452_/a_836_156# vdd 0.002533f
C5038 FILLER_0_4_107/a_1380_472# _152_ 0.001297f
C5039 _101_ _099_ 0.198807f
C5040 net52 FILLER_0_5_72/a_1380_472# 0.001523f
C5041 net29 _094_ 0.313846f
C5042 net48 FILLER_0_7_233/a_36_472# 0.01015f
C5043 _450_/a_1697_156# net6 0.00236f
C5044 net56 FILLER_0_17_142/a_124_375# 0.004803f
C5045 _041_ FILLER_0_18_37/a_1380_472# 0.003776f
C5046 mask\[0\] _429_/a_796_472# 0.007281f
C5047 net16 _042_ 0.012486f
C5048 _308_/a_1084_68# _115_ 0.001451f
C5049 net55 FILLER_0_18_53/a_572_375# 0.015895f
C5050 result[6] ctlp[2] 0.001324f
C5051 FILLER_0_18_177/a_1828_472# vdd 0.004845f
C5052 FILLER_0_18_177/a_1380_472# vss -0.001894f
C5053 _008_ _094_ 0.234346f
C5054 _132_ _428_/a_1456_156# 0.001009f
C5055 output47/a_224_472# FILLER_0_15_2/a_484_472# 0.038484f
C5056 net72 FILLER_0_21_28/a_572_375# 0.005742f
C5057 _133_ _163_ 0.034905f
C5058 FILLER_0_20_177/a_1468_375# _098_ 0.012889f
C5059 _428_/a_2560_156# _131_ 0.002853f
C5060 _093_ FILLER_0_18_107/a_2276_472# 0.001996f
C5061 net35 FILLER_0_22_128/a_124_375# 0.010439f
C5062 _057_ vss 0.169369f
C5063 _379_/a_36_472# _035_ 0.002226f
C5064 FILLER_0_4_123/a_124_375# trim_mask\[4\] 0.004312f
C5065 FILLER_0_5_212/a_36_472# net59 0.058827f
C5066 _136_ _040_ 0.788826f
C5067 _174_ _043_ 0.964645f
C5068 FILLER_0_7_72/a_124_375# FILLER_0_7_59/a_572_375# 0.003228f
C5069 _256_/a_36_68# _070_ 0.019259f
C5070 _256_/a_1164_497# _076_ 0.001871f
C5071 _376_/a_36_160# _163_ 0.006811f
C5072 mask\[4\] FILLER_0_17_218/a_484_472# 0.001232f
C5073 net58 _425_/a_448_472# 0.002474f
C5074 net75 _425_/a_1000_472# 0.038919f
C5075 FILLER_0_10_78/a_124_375# FILLER_0_11_78/a_124_375# 0.05841f
C5076 net41 _446_/a_2560_156# 0.005695f
C5077 _053_ FILLER_0_5_54/a_1380_472# 0.00114f
C5078 FILLER_0_16_57/a_1468_375# vss 0.062643f
C5079 FILLER_0_16_57/a_36_472# vdd 0.088011f
C5080 FILLER_0_16_107/a_572_375# _093_ 0.002827f
C5081 net50 FILLER_0_8_24/a_124_375# 0.001597f
C5082 net57 _137_ 0.006142f
C5083 FILLER_0_22_128/a_572_375# vss 0.00243f
C5084 FILLER_0_22_128/a_1020_375# vdd 0.002503f
C5085 FILLER_0_5_128/a_36_472# net74 0.01163f
C5086 net2 vss 0.213737f
C5087 _415_/a_1308_423# net18 0.010051f
C5088 _428_/a_36_151# FILLER_0_13_100/a_36_472# 0.004032f
C5089 net64 FILLER_0_12_236/a_572_375# 0.005704f
C5090 FILLER_0_5_198/a_484_472# net21 0.051161f
C5091 _414_/a_796_472# cal_itt\[3\] 0.019699f
C5092 net76 net19 0.02061f
C5093 _233_/a_36_160# net17 0.003831f
C5094 output17/a_224_472# vss 0.009426f
C5095 _441_/a_1204_472# _168_ 0.009437f
C5096 trim_mask\[2\] _168_ 0.00704f
C5097 net16 FILLER_0_14_50/a_36_472# 0.001377f
C5098 _141_ mask\[2\] 0.084094f
C5099 FILLER_0_2_93/a_124_375# net14 0.007439f
C5100 net63 FILLER_0_20_177/a_1468_375# 0.018435f
C5101 FILLER_0_5_72/a_932_472# _164_ 0.011079f
C5102 _000_ _253_/a_244_68# 0.001243f
C5103 net75 _253_/a_1100_68# 0.001047f
C5104 mask\[0\] FILLER_0_14_235/a_36_472# 0.287093f
C5105 net41 _054_ 0.035503f
C5106 FILLER_0_19_47/a_124_375# _013_ 0.023766f
C5107 cal_count\[3\] FILLER_0_11_78/a_484_472# 0.011737f
C5108 _098_ FILLER_0_19_171/a_484_472# 0.010731f
C5109 _079_ FILLER_0_5_206/a_124_375# 0.009128f
C5110 _367_/a_244_472# _157_ 0.002529f
C5111 net41 cal_count\[2\] 0.079279f
C5112 _428_/a_448_472# net70 0.007116f
C5113 FILLER_0_5_172/a_36_472# vss 0.003406f
C5114 _085_ _310_/a_49_472# 0.001093f
C5115 result[8] mask\[6\] 0.111221f
C5116 FILLER_0_21_28/a_124_375# net40 0.060428f
C5117 _279_/a_652_68# vdd 0.001562f
C5118 _132_ _345_/a_36_160# 0.078243f
C5119 fanout80/a_36_113# _138_ 0.002489f
C5120 FILLER_0_16_57/a_572_375# net15 0.013085f
C5121 net16 cal_count\[3\] 0.082821f
C5122 FILLER_0_18_2/a_1468_375# net38 0.016983f
C5123 _074_ _122_ 0.300373f
C5124 FILLER_0_9_60/a_484_472# FILLER_0_9_72/a_36_472# 0.002296f
C5125 trimb[1] FILLER_0_20_15/a_484_472# 0.001292f
C5126 _126_ _129_ 0.039006f
C5127 _413_/a_2248_156# ctln[4] 0.001253f
C5128 _067_ _450_/a_1353_112# 0.007106f
C5129 _188_ FILLER_0_12_50/a_36_472# 0.006464f
C5130 _130_ _129_ 0.021732f
C5131 FILLER_0_14_50/a_124_375# vdd 0.026996f
C5132 _064_ _033_ 0.001986f
C5133 _132_ _043_ 0.038747f
C5134 net54 FILLER_0_20_98/a_36_472# 0.059367f
C5135 _081_ _160_ 0.00816f
C5136 FILLER_0_9_72/a_124_375# vdd -0.003896f
C5137 net82 FILLER_0_3_172/a_572_375# 0.010972f
C5138 _119_ vdd 0.38257f
C5139 _214_/a_36_160# _437_/a_36_151# 0.001542f
C5140 _142_ _341_/a_49_472# 0.011026f
C5141 FILLER_0_6_47/a_3172_472# vss 0.014726f
C5142 net75 FILLER_0_8_247/a_1468_375# 0.047331f
C5143 FILLER_0_15_150/a_124_375# FILLER_0_15_142/a_572_375# 0.012001f
C5144 _093_ FILLER_0_17_72/a_484_472# 0.008637f
C5145 _406_/a_36_159# cal_count\[2\] 0.028829f
C5146 net55 net17 0.056153f
C5147 _269_/a_36_472# vdd 0.03432f
C5148 mask\[4\] FILLER_0_18_209/a_124_375# 0.020811f
C5149 trim_mask\[4\] _163_ 0.003686f
C5150 FILLER_0_7_146/a_36_472# _059_ 0.073041f
C5151 FILLER_0_11_142/a_36_472# vss 0.008744f
C5152 FILLER_0_11_142/a_484_472# vdd 0.006641f
C5153 vss cal_count\[0\] 0.160743f
C5154 _026_ vdd 0.15542f
C5155 _425_/a_448_472# FILLER_0_8_247/a_932_472# 0.012285f
C5156 net81 _429_/a_2665_112# 0.012675f
C5157 FILLER_0_6_239/a_36_472# _122_ 0.01785f
C5158 net18 _417_/a_36_151# 0.020548f
C5159 net27 FILLER_0_14_235/a_484_472# 0.010072f
C5160 _144_ _141_ 0.095441f
C5161 FILLER_0_15_212/a_124_375# FILLER_0_15_205/a_124_375# 0.004426f
C5162 FILLER_0_12_236/a_572_375# vss 0.025768f
C5163 FILLER_0_12_236/a_36_472# vdd 0.086431f
C5164 output10/a_224_472# ctln[1] 0.083631f
C5165 net38 net39 0.066083f
C5166 net75 _426_/a_36_151# 0.070626f
C5167 FILLER_0_10_37/a_124_375# FILLER_0_10_28/a_124_375# 0.003228f
C5168 FILLER_0_21_206/a_124_375# vdd 0.038521f
C5169 FILLER_0_16_89/a_124_375# _136_ 0.011795f
C5170 net82 FILLER_0_3_221/a_36_472# 0.015923f
C5171 result[6] _420_/a_1308_423# 0.008756f
C5172 _097_ vdd 0.191424f
C5173 _104_ _421_/a_1308_423# 0.001621f
C5174 _093_ FILLER_0_19_111/a_572_375# 0.002743f
C5175 FILLER_0_18_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001597f
C5176 FILLER_0_4_49/a_572_375# _440_/a_36_151# 0.073306f
C5177 _074_ FILLER_0_6_231/a_484_472# 0.004409f
C5178 result[0] calibrate 0.00287f
C5179 net20 result[9] 1.593573f
C5180 _098_ FILLER_0_15_212/a_124_375# 0.008125f
C5181 _390_/a_36_68# _172_ 0.033476f
C5182 _074_ _061_ 0.007152f
C5183 _350_/a_49_472# net23 0.002397f
C5184 _103_ vdd 0.590261f
C5185 net60 vss 0.382678f
C5186 net78 vss 0.167812f
C5187 _072_ _121_ 0.041039f
C5188 FILLER_0_23_88/a_124_375# net14 0.002894f
C5189 FILLER_0_17_72/a_1916_375# net36 0.015395f
C5190 net15 FILLER_0_6_47/a_2276_472# 0.049487f
C5191 output44/a_224_472# trimb[1] 0.046391f
C5192 mask\[5\] _143_ 0.032539f
C5193 net57 FILLER_0_13_142/a_932_472# 0.01158f
C5194 net57 net56 0.054294f
C5195 mask\[5\] _348_/a_49_472# 0.025962f
C5196 _004_ output28/a_224_472# 0.024204f
C5197 FILLER_0_12_124/a_124_375# _428_/a_36_151# 0.058722f
C5198 _343_/a_49_472# _137_ 0.001419f
C5199 net51 FILLER_0_12_28/a_36_472# 0.005661f
C5200 net25 FILLER_0_22_86/a_572_375# 0.002444f
C5201 net75 _265_/a_916_472# 0.001686f
C5202 _077_ _129_ 0.08682f
C5203 _422_/a_36_151# _299_/a_36_472# 0.004432f
C5204 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_484_472# 0.013277f
C5205 FILLER_0_4_197/a_1380_472# _088_ 0.017451f
C5206 _131_ FILLER_0_10_107/a_572_375# 0.007252f
C5207 FILLER_0_21_28/a_484_472# vdd 0.011209f
C5208 _052_ _424_/a_2248_156# 0.005116f
C5209 output15/a_224_472# net49 0.005626f
C5210 _211_/a_36_160# vdd 0.030216f
C5211 _287_/a_36_472# _102_ 0.028733f
C5212 _013_ net15 0.152142f
C5213 FILLER_0_3_172/a_3172_472# vdd 0.003804f
C5214 FILLER_0_5_88/a_124_375# net47 0.005083f
C5215 _099_ _282_/a_36_160# 0.005808f
C5216 _314_/a_224_472# vss 0.001399f
C5217 net23 FILLER_0_21_150/a_124_375# 0.045928f
C5218 _242_/a_36_160# _170_ 0.001933f
C5219 _117_ _310_/a_1133_69# 0.002654f
C5220 result[6] _421_/a_1000_472# 0.024206f
C5221 _091_ net36 0.067629f
C5222 _084_ _316_/a_124_24# 0.001501f
C5223 net63 FILLER_0_15_212/a_124_375# 0.001597f
C5224 _256_/a_244_497# vss 0.001274f
C5225 FILLER_0_11_101/a_484_472# _120_ 0.011393f
C5226 mask\[8\] _433_/a_36_151# 0.001402f
C5227 _144_ _433_/a_2665_112# 0.030413f
C5228 en cal_itt\[1\] 0.028447f
C5229 output32/a_224_472# net18 0.022521f
C5230 FILLER_0_5_109/a_484_472# _153_ 0.071582f
C5231 _088_ net82 0.160444f
C5232 net16 _379_/a_36_472# 0.01109f
C5233 trim_val\[0\] trim_mask\[1\] 0.003033f
C5234 FILLER_0_17_64/a_36_472# vss 0.006428f
C5235 net53 net36 3.423337f
C5236 FILLER_0_4_49/a_572_375# vdd 0.005972f
C5237 _443_/a_2665_112# _037_ 0.004052f
C5238 calibrate _062_ 2.032477f
C5239 output48/a_224_472# calibrate 0.003223f
C5240 net76 FILLER_0_3_172/a_484_472# 0.002542f
C5241 _131_ FILLER_0_17_104/a_1380_472# 0.004125f
C5242 net48 net59 0.015963f
C5243 _426_/a_36_151# FILLER_0_8_247/a_1468_375# 0.059049f
C5244 _413_/a_2248_156# FILLER_0_3_212/a_124_375# 0.030666f
C5245 vss _433_/a_36_151# 0.00618f
C5246 vdd _433_/a_448_472# 0.003821f
C5247 net56 FILLER_0_18_139/a_1020_375# 0.018398f
C5248 _175_ FILLER_0_15_72/a_484_472# 0.020589f
C5249 valid en 0.026142f
C5250 net48 net4 0.099614f
C5251 _093_ mask\[8\] 0.004026f
C5252 FILLER_0_20_177/a_1020_375# _434_/a_36_151# 0.059049f
C5253 _425_/a_448_472# _014_ 0.013561f
C5254 _069_ _043_ 0.04044f
C5255 _147_ vss 0.006333f
C5256 _118_ _311_/a_3740_473# 0.001244f
C5257 FILLER_0_21_142/a_572_375# net23 0.007884f
C5258 net38 _452_/a_2449_156# 0.058386f
C5259 FILLER_0_3_78/a_572_375# vss 0.04008f
C5260 FILLER_0_3_78/a_36_472# vdd 0.082597f
C5261 net72 _424_/a_36_151# 0.09381f
C5262 _431_/a_1288_156# net73 0.001033f
C5263 output39/a_224_472# _063_ 0.001019f
C5264 net39 _233_/a_36_160# 0.017979f
C5265 mask\[3\] FILLER_0_18_177/a_36_472# 0.005668f
C5266 _321_/a_170_472# vss 0.024882f
C5267 ctlp[4] ctlp[3] 0.027598f
C5268 FILLER_0_13_228/a_36_472# vss 0.006491f
C5269 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_572_375# 0.001597f
C5270 _141_ _339_/a_36_160# 0.011118f
C5271 FILLER_0_2_101/a_36_472# vss 0.004743f
C5272 FILLER_0_4_107/a_36_472# vdd 0.119007f
C5273 FILLER_0_4_107/a_1468_375# vss 0.055184f
C5274 _093_ vss 2.002012f
C5275 _114_ _267_/a_672_472# 0.001566f
C5276 _417_/a_36_151# net62 0.044051f
C5277 net53 FILLER_0_14_123/a_124_375# 0.003138f
C5278 input5/a_36_113# clk 0.01086f
C5279 net67 _450_/a_36_151# 0.067819f
C5280 fanout78/a_36_113# _007_ 0.003126f
C5281 FILLER_0_5_117/a_36_472# FILLER_0_5_109/a_484_472# 0.013276f
C5282 FILLER_0_18_2/a_1468_375# net55 0.007169f
C5283 _301_/a_36_472# net25 0.003165f
C5284 output25/a_224_472# ctlp[8] 0.018544f
C5285 net46 FILLER_0_21_28/a_124_375# 0.011995f
C5286 _091_ FILLER_0_20_169/a_36_472# 0.007537f
C5287 _086_ FILLER_0_5_172/a_124_375# 0.007355f
C5288 _321_/a_170_472# net74 0.020269f
C5289 result[4] _417_/a_2560_156# 0.001076f
C5290 vdd FILLER_0_19_134/a_36_472# 0.092128f
C5291 vss FILLER_0_19_134/a_124_375# 0.021427f
C5292 result[8] net35 0.001362f
C5293 _086_ _128_ 0.085571f
C5294 _195_/a_67_603# net62 0.002422f
C5295 output24/a_224_472# _050_ 0.061723f
C5296 net28 mask\[1\] 0.572459f
C5297 _369_/a_36_68# _157_ 0.068266f
C5298 _186_ _067_ 0.001907f
C5299 FILLER_0_5_128/a_124_375# _163_ 0.009765f
C5300 FILLER_0_19_171/a_36_472# _434_/a_36_151# 0.00271f
C5301 _363_/a_36_68# _086_ 0.007567f
C5302 FILLER_0_9_28/a_36_472# net17 0.012954f
C5303 net34 ctlp[2] 0.953441f
C5304 _448_/a_36_151# FILLER_0_2_177/a_36_472# 0.04556f
C5305 FILLER_0_9_290/a_124_375# vss 0.033914f
C5306 FILLER_0_9_290/a_36_472# vdd 0.094552f
C5307 ctln[6] FILLER_0_0_130/a_36_472# 0.023355f
C5308 _136_ FILLER_0_14_99/a_36_472# 0.01535f
C5309 _179_ _180_ 0.018662f
C5310 net32 _107_ 0.003155f
C5311 FILLER_0_5_206/a_36_472# vdd 0.090007f
C5312 FILLER_0_5_206/a_124_375# vss 0.050652f
C5313 _069_ net21 0.032615f
C5314 _038_ _120_ 0.00117f
C5315 _019_ vdd 0.015401f
C5316 FILLER_0_21_142/a_484_472# mask\[7\] 0.001603f
C5317 _098_ mask\[6\] 0.297837f
C5318 net65 _412_/a_2248_156# 0.039861f
C5319 _077_ _219_/a_36_160# 0.01438f
C5320 FILLER_0_10_247/a_124_375# net64 0.001597f
C5321 _086_ FILLER_0_11_142/a_572_375# 0.011726f
C5322 FILLER_0_17_200/a_36_472# net63 0.005648f
C5323 ctln[7] net14 0.197449f
C5324 FILLER_0_18_100/a_36_472# net14 0.046864f
C5325 _449_/a_1000_472# _067_ 0.021759f
C5326 _402_/a_1948_68# _182_ 0.016049f
C5327 FILLER_0_7_195/a_36_472# calibrate 0.010951f
C5328 _033_ _444_/a_2248_156# 0.011578f
C5329 _081_ _265_/a_224_472# 0.008598f
C5330 _412_/a_36_151# output37/a_224_472# 0.006358f
C5331 _053_ FILLER_0_6_47/a_2364_375# 0.007053f
C5332 _068_ _311_/a_3740_473# 0.001409f
C5333 _436_/a_36_151# mask\[8\] 0.032521f
C5334 net76 FILLER_0_6_177/a_484_472# 0.016333f
C5335 _125_ _062_ 0.061735f
C5336 FILLER_0_19_195/a_124_375# vdd 0.03587f
C5337 output11/a_224_472# vss 0.083244f
C5338 _235_/a_255_603# trim_val\[2\] 0.002471f
C5339 FILLER_0_11_142/a_572_375# cal_count\[3\] 0.014082f
C5340 _417_/a_448_472# net30 0.042386f
C5341 _370_/a_1152_472# _152_ 0.001423f
C5342 _188_ _039_ 0.002071f
C5343 FILLER_0_18_2/a_2364_375# net40 0.002024f
C5344 net57 _095_ 0.07431f
C5345 _363_/a_36_68# _154_ 0.149319f
C5346 vdd _295_/a_36_472# 0.0083f
C5347 cal_itt\[3\] _375_/a_36_68# 0.005168f
C5348 _076_ _120_ 0.736844f
C5349 trim_mask\[2\] _447_/a_36_151# 0.022881f
C5350 _389_/a_36_148# vdd 0.039639f
C5351 net81 _094_ 0.004737f
C5352 cal_count\[3\] _373_/a_1254_68# 0.001391f
C5353 _445_/a_2665_112# net47 0.041188f
C5354 FILLER_0_4_185/a_36_472# _087_ 0.008805f
C5355 net18 _418_/a_36_151# 0.017941f
C5356 FILLER_0_17_142/a_124_375# vss 0.008753f
C5357 FILLER_0_17_142/a_572_375# vdd 0.012885f
C5358 output8/a_224_472# FILLER_0_3_221/a_124_375# 0.03228f
C5359 net28 vss 0.185012f
C5360 net38 net42 0.012245f
C5361 net63 mask\[6\] 0.146994f
C5362 _436_/a_448_472# vdd 0.038494f
C5363 FILLER_0_4_197/a_124_375# net59 0.001026f
C5364 _232_/a_67_603# _164_ 0.076123f
C5365 _440_/a_36_151# _029_ 0.00874f
C5366 ctln[2] net81 0.003762f
C5367 vdd _380_/a_224_472# 0.001733f
C5368 _430_/a_448_472# mask\[2\] 0.045973f
C5369 FILLER_0_18_76/a_124_375# vdd 0.019258f
C5370 FILLER_0_16_73/a_572_375# _131_ 0.011479f
C5371 vdd _416_/a_2665_112# 0.027256f
C5372 net54 FILLER_0_22_86/a_1468_375# 0.001597f
C5373 trimb[3] net17 0.005798f
C5374 trim[1] net40 0.043114f
C5375 mask\[9\] _098_ 0.256513f
C5376 _429_/a_2248_156# vdd -0.006752f
C5377 _429_/a_1204_472# vss 0.002428f
C5378 _075_ net21 0.012335f
C5379 _423_/a_1000_472# vdd 0.001833f
C5380 result[4] result[9] 0.101112f
C5381 FILLER_0_10_247/a_124_375# vss 0.006235f
C5382 FILLER_0_10_247/a_36_472# vdd 0.111658f
C5383 FILLER_0_20_98/a_124_375# _437_/a_36_151# 0.059049f
C5384 _104_ mask\[2\] 0.002737f
C5385 FILLER_0_8_263/a_124_375# net19 0.039576f
C5386 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_124_375# 0.001597f
C5387 _414_/a_796_472# _081_ 0.003538f
C5388 _414_/a_36_151# net22 0.014398f
C5389 FILLER_0_19_28/a_572_375# _452_/a_36_151# 0.0027f
C5390 net60 _103_ 0.066266f
C5391 net31 vdd 0.542738f
C5392 _136_ FILLER_0_16_154/a_1020_375# 0.004387f
C5393 net20 net61 0.014444f
C5394 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_36_472# 0.086635f
C5395 result[6] ctlp[1] 0.677825f
C5396 _285_/a_36_472# net36 0.003032f
C5397 FILLER_0_13_206/a_124_375# net4 0.031251f
C5398 FILLER_0_19_125/a_124_375# _022_ 0.055527f
C5399 _432_/a_2248_156# vdd 0.02369f
C5400 _008_ _419_/a_1000_472# 0.003267f
C5401 FILLER_0_17_161/a_36_472# vss 0.003343f
C5402 cal_itt\[2\] _080_ 0.062471f
C5403 net52 FILLER_0_6_47/a_2812_375# 0.018463f
C5404 _070_ FILLER_0_9_105/a_484_472# 0.020248f
C5405 _110_ net15 0.016359f
C5406 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1468_375# 0.086635f
C5407 _104_ result[7] 0.475003f
C5408 _424_/a_2665_112# vss 0.013462f
C5409 _024_ _435_/a_1308_423# 0.002661f
C5410 _098_ FILLER_0_19_111/a_36_472# 0.003915f
C5411 _150_ _438_/a_1000_472# 0.003452f
C5412 _066_ _163_ 0.006401f
C5413 _444_/a_1204_472# net17 0.021952f
C5414 ctlp[1] _421_/a_36_151# 0.010453f
C5415 net54 _437_/a_2665_112# 0.061157f
C5416 _427_/a_1308_423# net23 0.004863f
C5417 _442_/a_448_472# vdd 0.006758f
C5418 _442_/a_36_151# vss 0.021278f
C5419 net1 fanout59/a_36_160# 0.002325f
C5420 _323_/a_36_113# net4 0.005657f
C5421 net25 FILLER_0_23_88/a_36_472# 0.192699f
C5422 FILLER_0_4_177/a_36_472# _074_ 0.002603f
C5423 net55 _452_/a_2449_156# 0.015878f
C5424 result[7] _420_/a_36_151# 0.006868f
C5425 _446_/a_36_151# net17 0.006518f
C5426 _132_ _451_/a_448_472# 0.001197f
C5427 _447_/a_2560_156# vss 0.00126f
C5428 FILLER_0_18_2/a_2724_472# vdd 0.004348f
C5429 FILLER_0_18_2/a_2276_472# vss 0.001865f
C5430 net23 FILLER_0_5_148/a_484_472# 0.047258f
C5431 _316_/a_124_24# calibrate 0.016936f
C5432 _415_/a_448_472# net81 0.004045f
C5433 net15 _423_/a_448_472# 0.004833f
C5434 _431_/a_3041_156# vss 0.001312f
C5435 net20 net37 0.039674f
C5436 _445_/a_36_151# vdd 0.052935f
C5437 _029_ vdd 0.223076f
C5438 FILLER_0_4_197/a_1468_375# net76 0.007667f
C5439 _322_/a_124_24# _126_ 0.019609f
C5440 _029_ _365_/a_244_472# 0.001956f
C5441 FILLER_0_15_290/a_36_472# output30/a_224_472# 0.001711f
C5442 _412_/a_1456_156# net58 0.001045f
C5443 en net59 0.490893f
C5444 _411_/a_2665_112# vss 0.00238f
C5445 _411_/a_2560_156# vdd 0.001315f
C5446 FILLER_0_2_93/a_572_375# _030_ 0.001718f
C5447 comp FILLER_0_12_2/a_124_375# 0.007468f
C5448 FILLER_0_15_282/a_572_375# _417_/a_36_151# 0.001597f
C5449 ctln[6] net22 0.014307f
C5450 fanout71/a_36_113# net54 0.001194f
C5451 net47 FILLER_0_6_37/a_36_472# 0.001161f
C5452 _119_ FILLER_0_4_107/a_1468_375# 0.001695f
C5453 _116_ _161_ 0.008003f
C5454 en net4 0.125535f
C5455 FILLER_0_11_78/a_484_472# _120_ 0.016839f
C5456 net20 _108_ 0.125627f
C5457 _077_ _453_/a_448_472# 0.057515f
C5458 net41 _402_/a_56_567# 0.021641f
C5459 _074_ net8 0.001023f
C5460 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_484_472# 0.026657f
C5461 mask\[1\] FILLER_0_15_205/a_36_472# 0.006921f
C5462 _163_ net37 0.079552f
C5463 _076_ _227_/a_36_160# 0.004997f
C5464 net23 FILLER_0_19_155/a_36_472# 0.019429f
C5465 FILLER_0_14_263/a_36_472# net62 0.019591f
C5466 _123_ vdd 0.214703f
C5467 output10/a_224_472# net19 0.037774f
C5468 mask\[7\] _435_/a_448_472# 0.064472f
C5469 net16 _120_ 0.009918f
C5470 comp vdd 0.108153f
C5471 net63 FILLER_0_19_187/a_572_375# 0.049706f
C5472 trim_val\[0\] _054_ 0.010002f
C5473 _056_ _226_/a_1044_68# 0.002852f
C5474 FILLER_0_12_20/a_36_472# _039_ 0.007881f
C5475 _091_ FILLER_0_16_154/a_1468_375# 0.003056f
C5476 output34/a_224_472# _421_/a_2665_112# 0.00151f
C5477 result[7] _421_/a_1308_423# 0.022204f
C5478 _447_/a_2248_156# net15 0.01843f
C5479 _390_/a_244_472# _038_ 0.001278f
C5480 _390_/a_36_68# _136_ 0.032598f
C5481 net44 FILLER_0_20_2/a_36_472# 0.037627f
C5482 net50 _033_ 0.003088f
C5483 _144_ FILLER_0_21_125/a_124_375# 0.009117f
C5484 _418_/a_36_151# net62 0.029844f
C5485 _406_/a_36_159# _402_/a_56_567# 0.001025f
C5486 FILLER_0_16_107/a_36_472# _131_ 0.008817f
C5487 FILLER_0_20_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001543f
C5488 FILLER_0_2_101/a_124_375# _154_ 0.003932f
C5489 FILLER_0_4_107/a_124_375# _153_ 0.073219f
C5490 FILLER_0_4_107/a_1020_375# _154_ 0.013746f
C5491 _053_ _377_/a_36_472# 0.023504f
C5492 mask\[5\] FILLER_0_18_177/a_36_472# 0.001063f
C5493 _093_ _103_ 0.124026f
C5494 _036_ fanout66/a_36_113# 0.014556f
C5495 net36 FILLER_0_16_115/a_36_472# 0.003805f
C5496 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_124_375# 0.026339f
C5497 _115_ FILLER_0_10_94/a_484_472# 0.015061f
C5498 _408_/a_1336_472# _095_ 0.011305f
C5499 _072_ _375_/a_1388_497# 0.001138f
C5500 mask\[2\] FILLER_0_16_154/a_484_472# 0.028444f
C5501 FILLER_0_13_142/a_36_472# _043_ 0.011974f
C5502 output12/a_224_472# _037_ 0.00827f
C5503 FILLER_0_18_2/a_2724_472# _452_/a_1040_527# 0.001138f
C5504 FILLER_0_18_2/a_932_472# _452_/a_2225_156# 0.001256f
C5505 FILLER_0_14_91/a_484_472# _176_ 0.003624f
C5506 net35 _098_ 0.017288f
C5507 _176_ state\[1\] 0.001641f
C5508 output37/a_224_472# _425_/a_2248_156# 0.00114f
C5509 output28/a_224_472# fanout79/a_36_160# 0.022393f
C5510 _272_/a_36_472# _087_ 0.048282f
C5511 _390_/a_36_68# _070_ 0.047478f
C5512 _306_/a_36_68# state\[1\] 0.028553f
C5513 net17 FILLER_0_20_15/a_36_472# 0.004375f
C5514 FILLER_0_15_142/a_484_472# net56 0.003214f
C5515 output33/a_224_472# vss 0.05089f
C5516 net57 vss 0.818311f
C5517 _414_/a_1000_472# _003_ 0.002053f
C5518 _143_ _340_/a_36_160# 0.001064f
C5519 cal cal_itt\[1\] 0.036277f
C5520 mask\[4\] _091_ 0.071954f
C5521 FILLER_0_15_205/a_36_472# vss 0.003239f
C5522 _340_/a_36_160# _348_/a_49_472# 0.001528f
C5523 FILLER_0_9_28/a_1828_472# vss 0.001663f
C5524 FILLER_0_9_28/a_2276_472# vdd 0.003276f
C5525 result[8] FILLER_0_21_206/a_36_472# 0.001292f
C5526 FILLER_0_12_2/a_484_472# _039_ 0.003082f
C5527 net72 _404_/a_36_472# 0.019911f
C5528 _135_ vss 0.097337f
C5529 FILLER_0_17_56/a_484_472# vss 0.006298f
C5530 FILLER_0_18_53/a_124_375# FILLER_0_18_37/a_1468_375# 0.012222f
C5531 net57 net74 2.360287f
C5532 net23 FILLER_0_22_128/a_2812_375# 0.050811f
C5533 net52 FILLER_0_2_111/a_932_472# 0.061249f
C5534 _372_/a_358_69# _070_ 0.001293f
C5535 cal valid 0.06045f
C5536 _444_/a_448_472# net40 0.055844f
C5537 _043_ _090_ 0.001578f
C5538 net63 net35 0.126544f
C5539 _161_ _117_ 0.25528f
C5540 fanout54/a_36_160# FILLER_0_19_155/a_124_375# 0.005705f
C5541 net80 vdd 1.045288f
C5542 FILLER_0_17_72/a_932_472# _131_ 0.002672f
C5543 _092_ _291_/a_36_160# 0.03297f
C5544 FILLER_0_9_105/a_124_375# vdd 0.029831f
C5545 net74 _135_ 0.002261f
C5546 _105_ _107_ 0.020727f
C5547 FILLER_0_4_185/a_124_375# vss 0.024832f
C5548 FILLER_0_4_185/a_36_472# vdd 0.122463f
C5549 net20 _092_ 0.001458f
C5550 FILLER_0_15_212/a_1468_375# net62 0.001106f
C5551 net38 FILLER_0_15_2/a_484_472# 0.003391f
C5552 FILLER_0_13_206/a_124_375# net79 0.009649f
C5553 FILLER_0_18_139/a_1020_375# vss 0.032606f
C5554 FILLER_0_18_139/a_1468_375# vdd 0.015542f
C5555 FILLER_0_1_204/a_36_472# net59 0.067975f
C5556 net65 FILLER_0_3_172/a_572_375# 0.008318f
C5557 _086_ _395_/a_1492_488# 0.001769f
C5558 _158_ _154_ 0.008872f
C5559 _043_ net22 0.041447f
C5560 net49 FILLER_0_3_54/a_36_472# 0.00186f
C5561 FILLER_0_5_72/a_36_472# _440_/a_36_151# 0.001723f
C5562 net15 FILLER_0_17_56/a_572_375# 0.007386f
C5563 result[7] FILLER_0_24_274/a_932_472# 0.006454f
C5564 _091_ FILLER_0_12_220/a_1020_375# 0.001598f
C5565 _069_ _062_ 0.029863f
C5566 _100_ vdd 0.212037f
C5567 net68 FILLER_0_3_54/a_36_472# 0.049455f
C5568 _037_ net12 0.007817f
C5569 output9/a_224_472# input4/a_36_68# 0.009732f
C5570 _370_/a_124_24# vdd 0.018613f
C5571 mask\[7\] FILLER_0_22_128/a_36_472# 0.013408f
C5572 _080_ net59 0.038227f
C5573 _305_/a_36_159# vdd 0.017293f
C5574 _067_ FILLER_0_12_28/a_36_472# 0.0127f
C5575 _148_ FILLER_0_22_128/a_36_472# 0.010386f
C5576 net35 FILLER_0_22_128/a_3172_472# 0.014415f
C5577 FILLER_0_15_116/a_124_375# _451_/a_36_151# 0.006111f
C5578 _090_ net21 0.038093f
C5579 _412_/a_36_151# net48 0.001091f
C5580 net4 _080_ 0.076128f
C5581 net36 _451_/a_2449_156# 0.016229f
C5582 FILLER_0_2_111/a_36_472# trim_mask\[3\] 0.007915f
C5583 ctlp[4] mask\[6\] 0.003054f
C5584 net16 _446_/a_2248_156# 0.010032f
C5585 _379_/a_36_472# _063_ 0.071695f
C5586 _116_ _071_ 0.017991f
C5587 net68 FILLER_0_6_47/a_932_472# 0.014935f
C5588 _436_/a_36_151# _211_/a_36_160# 0.068534f
C5589 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_572_375# 0.086635f
C5590 net38 _160_ 0.00247f
C5591 FILLER_0_18_107/a_124_375# vdd 0.030961f
C5592 _028_ _439_/a_1000_472# 0.003267f
C5593 trim_mask\[1\] FILLER_0_6_47/a_1828_472# 0.007542f
C5594 _093_ FILLER_0_19_134/a_36_472# 0.002415f
C5595 _180_ _041_ 0.00244f
C5596 _132_ _431_/a_36_151# 0.051016f
C5597 output31/a_224_472# net20 0.004424f
C5598 net67 FILLER_0_9_60/a_484_472# 0.001345f
C5599 net31 net60 0.012623f
C5600 result[4] net61 0.023257f
C5601 _343_/a_49_472# vss 0.002581f
C5602 FILLER_0_16_89/a_1380_472# _451_/a_1353_112# 0.010457f
C5603 _052_ FILLER_0_18_37/a_484_472# 0.003861f
C5604 net17 _164_ 0.007595f
C5605 FILLER_0_7_72/a_3172_472# net14 0.046751f
C5606 result[9] FILLER_0_24_274/a_1020_375# 0.001657f
C5607 net76 FILLER_0_5_198/a_572_375# 0.006974f
C5608 _377_/a_36_472# _164_ 0.03259f
C5609 _181_ _180_ 0.216908f
C5610 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_124_375# 0.005439f
C5611 _017_ FILLER_0_13_100/a_124_375# 0.001274f
C5612 FILLER_0_21_28/a_1828_472# _423_/a_36_151# 0.059367f
C5613 net22 net21 1.937266f
C5614 _144_ _354_/a_49_472# 0.03742f
C5615 _073_ net37 0.013152f
C5616 _421_/a_448_472# net19 0.058446f
C5617 _081_ _059_ 0.04053f
C5618 net54 net71 0.536043f
C5619 FILLER_0_19_55/a_124_375# _013_ 0.009611f
C5620 FILLER_0_24_274/a_124_375# vdd 0.012632f
C5621 FILLER_0_11_282/a_36_472# _416_/a_448_472# 0.011962f
C5622 FILLER_0_12_136/a_572_375# state\[2\] 0.001955f
C5623 FILLER_0_12_136/a_1468_375# net53 0.002709f
C5624 FILLER_0_5_72/a_36_472# vdd 0.107678f
C5625 FILLER_0_5_72/a_1468_375# vss 0.057097f
C5626 net81 net21 0.185411f
C5627 FILLER_0_8_107/a_124_375# _219_/a_36_160# 0.002515f
C5628 output10/a_224_472# cal_itt\[0\] 0.008003f
C5629 trim[0] net66 0.376153f
C5630 net70 _017_ 0.015488f
C5631 FILLER_0_1_98/a_36_472# net14 0.023583f
C5632 _128_ _120_ 0.053476f
C5633 trim[4] vss 0.033925f
C5634 _086_ _311_/a_2700_473# 0.00176f
C5635 _415_/a_36_151# vdd 0.115639f
C5636 net34 ctlp[1] 0.127025f
C5637 _408_/a_1336_472# vss 0.001022f
C5638 _408_/a_728_93# vdd 0.024163f
C5639 net63 FILLER_0_18_177/a_2276_472# 0.012025f
C5640 FILLER_0_15_142/a_484_472# _095_ 0.001509f
C5641 _096_ _306_/a_36_68# 0.016266f
C5642 _221_/a_36_160# vdd 0.073414f
C5643 _096_ _335_/a_49_472# 0.00151f
C5644 ctln[7] _442_/a_2248_156# 0.006094f
C5645 _093_ FILLER_0_17_142/a_572_375# 0.009547f
C5646 FILLER_0_15_150/a_124_375# vdd 0.026143f
C5647 _058_ net14 0.40635f
C5648 net20 _122_ 0.046817f
C5649 _129_ vss 0.141494f
C5650 FILLER_0_11_142/a_572_375# _120_ 0.009014f
C5651 FILLER_0_17_72/a_1380_472# _150_ 0.014154f
C5652 FILLER_0_15_116/a_36_472# _095_ 0.001098f
C5653 net50 _441_/a_36_151# 0.060777f
C5654 net52 _441_/a_1308_423# 0.059264f
C5655 _028_ FILLER_0_7_72/a_2724_472# 0.001777f
C5656 FILLER_0_9_28/a_36_472# net42 0.038355f
C5657 _119_ net57 0.30462f
C5658 fanout70/a_36_113# FILLER_0_15_116/a_484_472# 0.002001f
C5659 FILLER_0_13_212/a_124_375# net79 0.007396f
C5660 _093_ FILLER_0_18_76/a_124_375# 0.061549f
C5661 _429_/a_2248_156# FILLER_0_13_228/a_36_472# 0.035805f
C5662 net52 _440_/a_2248_156# 0.028463f
C5663 ctlp[5] _024_ 0.022549f
C5664 FILLER_0_23_274/a_124_375# vdd 0.014998f
C5665 output14/a_224_472# FILLER_0_0_130/a_124_375# 0.00515f
C5666 _272_/a_36_472# vdd 0.058326f
C5667 net52 _439_/a_448_472# 0.042072f
C5668 _129_ net74 0.476969f
C5669 _122_ _163_ 0.156898f
C5670 output44/a_224_472# FILLER_0_18_2/a_1020_375# 0.032639f
C5671 _053_ FILLER_0_7_72/a_932_472# 0.01339f
C5672 net55 net36 0.273956f
C5673 _425_/a_36_151# net37 0.003145f
C5674 net31 _093_ 0.274432f
C5675 mask\[4\] FILLER_0_18_177/a_3260_375# 0.013881f
C5676 _077_ FILLER_0_8_107/a_36_472# 0.007552f
C5677 net55 FILLER_0_19_28/a_36_472# 0.001572f
C5678 _010_ _420_/a_448_472# 0.027802f
C5679 net57 _097_ 0.100409f
C5680 _256_/a_36_68# calibrate 0.02084f
C5681 FILLER_0_7_72/a_2724_472# _308_/a_848_380# 0.001797f
C5682 _321_/a_358_69# net23 0.001718f
C5683 _432_/a_2248_156# _093_ 0.012955f
C5684 _434_/a_36_151# vss 0.006401f
C5685 _434_/a_448_472# vdd 0.020387f
C5686 FILLER_0_5_212/a_36_472# _081_ 0.01062f
C5687 _096_ FILLER_0_14_181/a_124_375# 0.002455f
C5688 _076_ net21 0.031683f
C5689 net41 output40/a_224_472# 0.018977f
C5690 net20 FILLER_0_6_231/a_484_472# 0.017025f
C5691 trimb[3] ctlp[0] 0.384753f
C5692 net69 FILLER_0_2_111/a_1020_375# 0.018655f
C5693 _031_ FILLER_0_2_111/a_124_375# 0.05482f
C5694 cal net59 0.297816f
C5695 net58 _264_/a_224_472# 0.001803f
C5696 net75 cal_itt\[1\] 0.704169f
C5697 _065_ _447_/a_448_472# 0.049072f
C5698 net1 net37 0.00519f
C5699 cal net4 0.026084f
C5700 FILLER_0_5_54/a_484_472# vdd 0.003166f
C5701 FILLER_0_5_54/a_36_472# vss 0.001756f
C5702 cal_count\[2\] _452_/a_36_151# 0.006982f
C5703 _242_/a_36_160# vdd 0.007995f
C5704 FILLER_0_20_31/a_36_472# net40 0.045181f
C5705 FILLER_0_17_133/a_124_375# _137_ 0.009198f
C5706 mask\[0\] _113_ 0.01678f
C5707 _441_/a_448_472# _164_ 0.016938f
C5708 FILLER_0_10_28/a_124_375# output6/a_224_472# 0.002633f
C5709 _071_ _225_/a_36_160# 0.002808f
C5710 _428_/a_2248_156# _427_/a_36_151# 0.035837f
C5711 net75 valid 0.002077f
C5712 _096_ _320_/a_672_472# 0.0082f
C5713 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_124_375# 0.001597f
C5714 net3 _278_/a_36_160# 0.014154f
C5715 FILLER_0_14_91/a_572_375# _136_ 0.049763f
C5716 _432_/a_2665_112# _139_ 0.004089f
C5717 FILLER_0_18_2/a_3260_375# FILLER_0_20_31/a_36_472# 0.001338f
C5718 _428_/a_2560_156# net74 0.002759f
C5719 net29 _044_ 0.01495f
C5720 net36 net23 0.028202f
C5721 _421_/a_796_472# _010_ 0.037434f
C5722 net20 FILLER_0_13_212/a_932_472# 0.003007f
C5723 cal_itt\[2\] net75 0.143064f
C5724 ctln[1] FILLER_0_1_266/a_36_472# 0.002068f
C5725 _443_/a_2560_156# vss 0.002467f
C5726 _322_/a_848_380# _118_ 0.047787f
C5727 net20 _288_/a_224_472# 0.003019f
C5728 _291_/a_36_160# FILLER_0_17_226/a_36_472# 0.035111f
C5729 net16 FILLER_0_17_38/a_572_375# 0.018281f
C5730 _428_/a_36_151# _332_/a_36_472# 0.004432f
C5731 _369_/a_36_68# _160_ 0.015312f
C5732 net55 _423_/a_2560_156# 0.002265f
C5733 _253_/a_36_68# _084_ 0.029805f
C5734 output27/a_224_472# result[0] 0.031252f
C5735 FILLER_0_7_72/a_1380_472# net52 0.003507f
C5736 FILLER_0_7_72/a_484_472# net50 0.059395f
C5737 net81 FILLER_0_15_212/a_1020_375# 0.006974f
C5738 _100_ FILLER_0_12_236/a_572_375# 0.015109f
C5739 vdd _022_ 0.082842f
C5740 FILLER_0_17_226/a_124_375# mask\[3\] 0.010642f
C5741 FILLER_0_2_177/a_124_375# net59 0.005212f
C5742 net28 _416_/a_2665_112# 0.008877f
C5743 _408_/a_718_524# FILLER_0_12_28/a_124_375# 0.001192f
C5744 net72 _176_ 0.059793f
C5745 FILLER_0_9_28/a_572_375# net50 0.002807f
C5746 _017_ FILLER_0_14_107/a_572_375# 0.003679f
C5747 net70 FILLER_0_14_107/a_1468_375# 0.007955f
C5748 output32/a_224_472# result[9] 0.047198f
C5749 _021_ mask\[3\] 0.036781f
C5750 net16 _043_ 0.049385f
C5751 _053_ FILLER_0_7_59/a_124_375# 0.015298f
C5752 output42/a_224_472# _444_/a_36_151# 0.002701f
C5753 _431_/a_2665_112# net36 0.001523f
C5754 net15 FILLER_0_5_54/a_1020_375# 0.015944f
C5755 FILLER_0_19_47/a_36_472# FILLER_0_18_37/a_1020_375# 0.001684f
C5756 net76 fanout76/a_36_160# 0.004503f
C5757 _104_ _298_/a_224_472# 0.001731f
C5758 _159_ _152_ 0.035925f
C5759 valid fanout65/a_36_113# 0.001646f
C5760 net27 _060_ 0.045136f
C5761 FILLER_0_16_57/a_484_472# _131_ 0.008223f
C5762 FILLER_0_17_38/a_124_375# vdd 0.01443f
C5763 FILLER_0_5_109/a_572_375# net47 0.011047f
C5764 net16 _185_ 0.086347f
C5765 mask\[3\] FILLER_0_16_241/a_36_472# 0.00209f
C5766 _162_ net47 0.004104f
C5767 _219_/a_36_160# vss 0.00157f
C5768 _098_ _433_/a_1308_423# 0.010653f
C5769 FILLER_0_3_2/a_124_375# vss 0.007235f
C5770 FILLER_0_3_2/a_36_472# vdd 0.106665f
C5771 FILLER_0_12_2/a_572_375# net3 0.001872f
C5772 _027_ vss 0.011873f
C5773 net34 FILLER_0_22_177/a_36_472# 0.003953f
C5774 net36 FILLER_0_15_180/a_484_472# 0.00702f
C5775 ctlp[1] _419_/a_2665_112# 0.009197f
C5776 mask\[9\] _438_/a_1308_423# 0.044336f
C5777 net23 _160_ 0.030085f
C5778 _412_/a_2248_156# vss 0.005692f
C5779 _412_/a_2665_112# vdd 0.014403f
C5780 _087_ _074_ 0.004231f
C5781 FILLER_0_19_125/a_124_375# net73 0.005414f
C5782 _037_ vss 0.051886f
C5783 FILLER_0_3_172/a_1468_375# net22 0.012895f
C5784 net40 _034_ 0.04333f
C5785 ctlp[3] vss 0.037106f
C5786 FILLER_0_15_142/a_484_472# vss 0.029611f
C5787 FILLER_0_17_72/a_1828_472# _438_/a_36_151# 0.001221f
C5788 output31/a_224_472# result[4] 0.049147f
C5789 _433_/a_2560_156# _145_ 0.007651f
C5790 FILLER_0_18_37/a_1380_472# vdd 0.004422f
C5791 output7/a_224_472# net40 0.009154f
C5792 net7 output40/a_224_472# 0.006944f
C5793 FILLER_0_15_142/a_572_375# _427_/a_36_151# 0.059049f
C5794 _322_/a_848_380# _068_ 0.009682f
C5795 _186_ _402_/a_728_93# 0.002381f
C5796 FILLER_0_14_91/a_36_472# net53 0.005849f
C5797 FILLER_0_15_228/a_124_375# net62 0.001408f
C5798 net76 FILLER_0_2_177/a_484_472# 0.012872f
C5799 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_36_472# 0.086743f
C5800 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_484_472# 0.013277f
C5801 net80 _147_ 0.022618f
C5802 FILLER_0_15_116/a_484_472# vdd 0.006111f
C5803 _408_/a_728_93# cal_count\[0\] 0.007633f
C5804 _413_/a_36_151# FILLER_0_3_172/a_1828_472# 0.001723f
C5805 _119_ _129_ 0.055585f
C5806 _086_ _131_ 0.886615f
C5807 net38 net67 1.762405f
C5808 cal_count\[2\] _402_/a_1948_68# 0.010022f
C5809 _412_/a_448_472# net76 0.026446f
C5810 FILLER_0_14_107/a_1380_472# _043_ 0.001641f
C5811 trimb[0] net17 0.006176f
C5812 _062_ _090_ 0.010805f
C5813 en_co_clk _067_ 0.272082f
C5814 _436_/a_2665_112# mask\[7\] 0.004274f
C5815 net80 _093_ 0.818824f
C5816 _416_/a_36_151# output30/a_224_472# 0.012025f
C5817 FILLER_0_9_223/a_484_472# _223_/a_36_160# 0.004695f
C5818 cal_count\[3\] _405_/a_67_603# 0.011131f
C5819 _436_/a_1204_472# _025_ 0.01349f
C5820 _131_ cal_count\[3\] 0.035391f
C5821 net52 net14 0.072003f
C5822 trim_val\[2\] net49 0.00301f
C5823 _441_/a_2248_156# net49 0.048164f
C5824 _073_ _122_ 0.002157f
C5825 _006_ net30 0.284414f
C5826 _095_ FILLER_0_13_142/a_1380_472# 0.001782f
C5827 _053_ _359_/a_36_488# 0.015831f
C5828 _053_ _078_ 0.137388f
C5829 _074_ _068_ 0.011897f
C5830 _086_ _114_ 1.371271f
C5831 _250_/a_36_68# state\[1\] 0.103037f
C5832 _093_ FILLER_0_18_139/a_1468_375# 0.004939f
C5833 trim_val\[3\] _441_/a_448_472# 0.00469f
C5834 FILLER_0_10_107/a_36_472# vdd 0.117291f
C5835 FILLER_0_10_107/a_572_375# vss 0.017711f
C5836 trim_val\[2\] net68 0.010894f
C5837 fanout81/a_36_160# cal_itt\[1\] 0.069457f
C5838 net81 _001_ 0.012492f
C5839 _445_/a_2248_156# net40 0.004545f
C5840 _013_ net26 0.174966f
C5841 input5/a_36_113# vss 0.005833f
C5842 FILLER_0_3_142/a_36_472# _443_/a_36_151# 0.001723f
C5843 _447_/a_796_472# net68 0.001593f
C5844 _447_/a_448_472# _036_ 0.015378f
C5845 _064_ _445_/a_796_472# 0.00673f
C5846 _131_ _154_ 0.019221f
C5847 net48 _081_ 0.137029f
C5848 _142_ _137_ 1.401722f
C5849 _114_ cal_count\[3\] 0.081644f
C5850 net32 net19 0.65591f
C5851 result[5] _418_/a_796_472# 0.001983f
C5852 FILLER_0_20_177/a_1468_375# vss 0.053913f
C5853 FILLER_0_20_177/a_36_472# vdd 0.114932f
C5854 _091_ FILLER_0_15_212/a_484_472# 0.049391f
C5855 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_124_375# 0.009654f
C5856 net72 _183_ 0.093818f
C5857 fanout80/a_36_113# net36 0.007625f
C5858 FILLER_0_7_104/a_932_472# _134_ 0.004249f
C5859 ctln[2] FILLER_0_0_266/a_36_472# 0.049163f
C5860 net81 output48/a_224_472# 0.040059f
C5861 _450_/a_36_151# output6/a_224_472# 0.134892f
C5862 FILLER_0_16_107/a_124_375# _451_/a_36_151# 0.001597f
C5863 net38 FILLER_0_8_24/a_484_472# 0.001223f
C5864 net70 FILLER_0_16_115/a_124_375# 0.025173f
C5865 FILLER_0_10_78/a_572_375# net52 0.003311f
C5866 output36/a_224_472# net19 0.106928f
C5867 FILLER_0_4_144/a_36_472# vdd 0.004289f
C5868 FILLER_0_4_144/a_572_375# vss 0.072463f
C5869 FILLER_0_17_104/a_1380_472# vss 0.001141f
C5870 _118_ _124_ 0.652002f
C5871 result[9] _419_/a_1204_472# 0.019627f
C5872 FILLER_0_5_54/a_1380_472# FILLER_0_6_47/a_2276_472# 0.026657f
C5873 _044_ result[3] 0.00251f
C5874 _093_ FILLER_0_18_107/a_124_375# 0.008393f
C5875 _081_ FILLER_0_6_177/a_124_375# 0.005524f
C5876 _411_/a_448_472# net75 0.072712f
C5877 mask\[2\] FILLER_0_15_212/a_1380_472# 0.001225f
C5878 net26 FILLER_0_21_28/a_2812_375# 0.001905f
C5879 _136_ _451_/a_1040_527# 0.00497f
C5880 net41 _444_/a_36_151# 0.013142f
C5881 _053_ FILLER_0_6_90/a_124_375# 0.003061f
C5882 net52 FILLER_0_9_72/a_484_472# 0.049391f
C5883 _343_/a_257_69# _093_ 0.001043f
C5884 FILLER_0_12_136/a_1468_375# _071_ 0.002023f
C5885 FILLER_0_15_59/a_484_472# vss 0.007866f
C5886 _008_ net77 0.029049f
C5887 _106_ FILLER_0_17_218/a_124_375# 0.004655f
C5888 _116_ _056_ 0.30649f
C5889 FILLER_0_21_133/a_124_375# _140_ 0.018383f
C5890 net29 _102_ 0.056837f
C5891 _453_/a_448_472# vss 0.00396f
C5892 _453_/a_1308_423# vdd 0.002896f
C5893 net10 FILLER_0_0_232/a_36_472# 0.016287f
C5894 _363_/a_36_68# _151_ 0.020916f
C5895 _003_ FILLER_0_5_181/a_124_375# 0.009929f
C5896 net54 FILLER_0_20_107/a_36_472# 0.050184f
C5897 FILLER_0_16_241/a_124_375# net36 0.004069f
C5898 net75 _316_/a_1084_68# 0.001531f
C5899 _375_/a_36_68# _161_ 0.028567f
C5900 net31 output33/a_224_472# 0.005087f
C5901 _429_/a_2665_112# _098_ 0.003225f
C5902 _002_ _270_/a_244_68# 0.001153f
C5903 net63 FILLER_0_19_195/a_36_472# 0.030832f
C5904 net75 net59 0.06935f
C5905 FILLER_0_15_212/a_124_375# mask\[1\] 0.007876f
C5906 FILLER_0_19_171/a_484_472# vss 0.001913f
C5907 FILLER_0_19_171/a_932_472# vdd 0.011399f
C5908 _196_/a_36_160# mask\[1\] 0.003254f
C5909 FILLER_0_14_181/a_124_375# FILLER_0_15_180/a_124_375# 0.026339f
C5910 _031_ vdd 0.327674f
C5911 _425_/a_36_151# _122_ 0.063131f
C5912 _425_/a_448_472# calibrate 0.105581f
C5913 _008_ _102_ 0.027578f
C5914 net75 net4 0.031823f
C5915 FILLER_0_9_28/a_2364_375# _220_/a_67_603# 0.002082f
C5916 _132_ _040_ 0.023821f
C5917 _079_ _088_ 0.012529f
C5918 _438_/a_796_472# vss 0.001171f
C5919 result[6] FILLER_0_23_290/a_124_375# 0.001492f
C5920 _289_/a_36_472# mask\[2\] 0.006392f
C5921 _004_ net81 0.993594f
C5922 _104_ mask\[7\] 0.069172f
C5923 net15 _012_ 0.043755f
C5924 _233_/a_36_160# net67 0.001315f
C5925 _394_/a_56_524# _174_ 0.015122f
C5926 _011_ _422_/a_1308_423# 0.001997f
C5927 net50 fanout67/a_36_160# 0.007195f
C5928 FILLER_0_17_72/a_1020_375# _451_/a_3129_107# 0.001202f
C5929 _320_/a_36_472# _055_ 0.001393f
C5930 cal_count\[1\] FILLER_0_15_59/a_484_472# 0.006408f
C5931 FILLER_0_15_282/a_124_375# _006_ 0.002249f
C5932 net16 _402_/a_1296_93# 0.053493f
C5933 FILLER_0_9_28/a_3260_375# net68 0.009969f
C5934 _086_ _126_ 0.063495f
C5935 net15 FILLER_0_15_59/a_572_375# 0.033245f
C5936 net32 _009_ 0.003756f
C5937 net73 FILLER_0_18_107/a_1828_472# 0.01544f
C5938 _086_ _130_ 0.008816f
C5939 _245_/a_234_472# _067_ 0.005071f
C5940 _333_/a_36_160# FILLER_0_15_180/a_36_472# 0.016014f
C5941 FILLER_0_16_89/a_932_472# net14 0.014714f
C5942 _076_ _062_ 0.978627f
C5943 _186_ net17 0.001172f
C5944 _432_/a_1204_472# net80 0.009362f
C5945 net47 _386_/a_848_380# 0.003045f
C5946 _322_/a_848_380# vdd 0.067623f
C5947 _322_/a_124_24# vss 0.003731f
C5948 _077_ _042_ 0.045685f
C5949 net80 FILLER_0_17_161/a_36_472# 0.003342f
C5950 output26/a_224_472# FILLER_0_23_44/a_932_472# 0.0323f
C5951 result[8] FILLER_0_24_274/a_572_375# 0.00726f
C5952 FILLER_0_21_125/a_124_375# mask\[7\] 0.00145f
C5953 _126_ cal_count\[3\] 0.418508f
C5954 FILLER_0_4_177/a_36_472# _163_ 0.002787f
C5955 _142_ net56 0.028797f
C5956 FILLER_0_1_98/a_124_375# _442_/a_2665_112# 0.003045f
C5957 _130_ cal_count\[3\] 0.037708f
C5958 _021_ mask\[5\] 0.001088f
C5959 net27 net64 1.364577f
C5960 FILLER_0_6_47/a_1468_375# vdd -0.014642f
C5961 FILLER_0_15_212/a_124_375# vss 0.005813f
C5962 FILLER_0_15_212/a_572_375# vdd -0.014642f
C5963 _369_/a_36_68# _156_ 0.001359f
C5964 FILLER_0_10_247/a_124_375# _100_ 0.001804f
C5965 FILLER_0_3_204/a_36_472# _413_/a_36_151# 0.001723f
C5966 _449_/a_36_151# FILLER_0_13_72/a_572_375# 0.035849f
C5967 input1/a_36_113# net1 0.003795f
C5968 _432_/a_2665_112# net63 0.067487f
C5969 FILLER_0_18_139/a_1380_472# net23 0.013087f
C5970 _322_/a_124_24# net74 0.05722f
C5971 _426_/a_2560_156# net64 0.00801f
C5972 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_36_472# 0.001723f
C5973 net58 net76 0.700034f
C5974 vdd _450_/a_2225_156# 0.020301f
C5975 _187_ _392_/a_36_68# 0.058263f
C5976 FILLER_0_7_72/a_572_375# FILLER_0_6_47/a_3260_375# 0.026339f
C5977 net53 _451_/a_836_156# 0.006521f
C5978 _008_ _198_/a_67_603# 0.012332f
C5979 mask\[0\] vdd 0.181371f
C5980 FILLER_0_8_247/a_124_375# calibrate 0.008393f
C5981 _074_ vdd 1.221102f
C5982 mask\[3\] _069_ 0.025564f
C5983 fanout54/a_36_160# net54 0.018583f
C5984 net35 _213_/a_67_603# 0.012955f
C5985 mask\[8\] _213_/a_255_603# 0.002776f
C5986 result[5] _010_ 0.00244f
C5987 net19 _419_/a_2560_156# 0.003213f
C5988 FILLER_0_17_104/a_1020_375# net14 0.002226f
C5989 _231_/a_244_68# _059_ 0.004384f
C5990 _056_ _117_ 0.065147f
C5991 _128_ net21 0.03068f
C5992 _204_/a_67_603# vdd 0.039556f
C5993 FILLER_0_10_78/a_1468_375# _171_ 0.034647f
C5994 _431_/a_2665_112# FILLER_0_18_139/a_1380_472# 0.001008f
C5995 _371_/a_36_113# vdd 0.007666f
C5996 _127_ _059_ 0.002878f
C5997 _057_ _267_/a_1120_472# 0.001833f
C5998 fanout70/a_36_113# net73 0.21211f
C5999 result[6] net33 0.363421f
C6000 FILLER_0_13_142/a_1380_472# vss 0.004953f
C6001 net16 _033_ 0.042852f
C6002 FILLER_0_20_31/a_124_375# FILLER_0_20_15/a_1468_375# 0.012001f
C6003 net18 FILLER_0_11_282/a_124_375# 0.042342f
C6004 fanout66/a_36_113# FILLER_0_3_54/a_36_472# 0.001645f
C6005 _077_ FILLER_0_9_72/a_572_375# 0.008103f
C6006 FILLER_0_9_28/a_1380_472# _120_ 0.00154f
C6007 FILLER_0_16_57/a_932_472# FILLER_0_15_59/a_572_375# 0.001543f
C6008 net82 _370_/a_848_380# 0.014538f
C6009 _086_ _077_ 0.058673f
C6010 FILLER_0_17_72/a_2724_472# _136_ 0.03065f
C6011 _453_/a_36_151# _042_ 0.035846f
C6012 _008_ mask\[3\] 0.799138f
C6013 FILLER_0_6_239/a_124_375# vss 0.017355f
C6014 FILLER_0_6_239/a_36_472# vdd 0.092399f
C6015 _210_/a_255_603# mask\[7\] 0.001329f
C6016 FILLER_0_16_73/a_572_375# vss 0.030752f
C6017 FILLER_0_16_73/a_36_472# vdd 0.08735f
C6018 _415_/a_36_151# net28 0.001195f
C6019 _433_/a_36_151# _022_ 0.017789f
C6020 result[8] FILLER_0_23_274/a_36_472# 0.001908f
C6021 mask\[4\] net23 0.111873f
C6022 ctlp[5] output23/a_224_472# 0.005152f
C6023 ctln[5] _448_/a_1204_472# 0.005186f
C6024 FILLER_0_3_172/a_1020_375# vdd 0.009809f
C6025 FILLER_0_1_266/a_36_472# net19 0.07227f
C6026 _077_ cal_count\[3\] 0.176576f
C6027 net27 vss 0.534444f
C6028 _422_/a_2248_156# vdd 0.005833f
C6029 ctln[2] net82 0.005498f
C6030 _449_/a_448_472# net72 0.01383f
C6031 ctln[0] output41/a_224_472# 0.001583f
C6032 output7/a_224_472# trim[3] 0.103375f
C6033 _122_ _121_ 0.034975f
C6034 _415_/a_2248_156# _416_/a_36_151# 0.001495f
C6035 fanout60/a_36_160# FILLER_0_17_282/a_124_375# 0.005489f
C6036 FILLER_0_10_78/a_1468_375# _176_ 0.013408f
C6037 _402_/a_56_567# _452_/a_36_151# 0.001915f
C6038 net55 FILLER_0_17_72/a_124_375# 0.019544f
C6039 net79 _018_ 0.069992f
C6040 _446_/a_1308_423# net66 0.005976f
C6041 _064_ _446_/a_2560_156# 0.029586f
C6042 net73 FILLER_0_19_111/a_124_375# 0.005778f
C6043 FILLER_0_3_221/a_36_472# vss 0.046345f
C6044 FILLER_0_3_221/a_484_472# vdd 0.002974f
C6045 _432_/a_448_472# mask\[3\] 0.005831f
C6046 net80 net57 0.002913f
C6047 result[7] _298_/a_224_472# 0.007724f
C6048 net54 FILLER_0_18_139/a_124_375# 0.002807f
C6049 _275_/a_224_472# _091_ 0.003461f
C6050 _000_ _080_ 0.002867f
C6051 ctln[4] FILLER_0_0_232/a_36_472# 0.012298f
C6052 _053_ _160_ 0.0539f
C6053 FILLER_0_20_193/a_124_375# _098_ 0.009717f
C6054 _451_/a_36_151# vdd 0.088651f
C6055 ctln[1] _411_/a_36_151# 0.018351f
C6056 FILLER_0_5_72/a_124_375# trim_mask\[1\] 0.010758f
C6057 FILLER_0_5_72/a_1468_375# _029_ 0.007876f
C6058 FILLER_0_3_172/a_2276_472# net21 0.003603f
C6059 fanout81/a_36_160# net4 0.002848f
C6060 _086_ _267_/a_224_472# 0.004041f
C6061 FILLER_0_20_98/a_124_375# net14 0.05242f
C6062 mask\[9\] FILLER_0_19_111/a_572_375# 0.027695f
C6063 ctln[3] net10 0.873575f
C6064 net26 _423_/a_448_472# 0.011612f
C6065 _413_/a_1000_472# net59 0.018099f
C6066 net34 _199_/a_36_160# 0.026709f
C6067 FILLER_0_17_200/a_36_472# vss 0.001182f
C6068 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_36_472# 0.009654f
C6069 _431_/a_1308_423# _136_ 0.027758f
C6070 net79 output30/a_224_472# 0.078502f
C6071 _105_ _205_/a_36_160# 0.001167f
C6072 output10/a_224_472# FILLER_0_0_232/a_124_375# 0.00363f
C6073 _057_ _074_ 0.013823f
C6074 FILLER_0_13_228/a_124_375# _043_ 0.133079f
C6075 FILLER_0_2_111/a_1468_375# vdd 0.011806f
C6076 net17 net43 0.144179f
C6077 net49 _167_ 0.031111f
C6078 cal_count\[3\] _453_/a_36_151# 0.023915f
C6079 output45/a_224_472# trimb[3] 0.076387f
C6080 _105_ net19 0.049611f
C6081 net41 FILLER_0_20_31/a_124_375# 0.049106f
C6082 _124_ vdd 0.040228f
C6083 net68 _167_ 0.001302f
C6084 net26 _424_/a_1204_472# 0.00194f
C6085 FILLER_0_18_107/a_2724_472# vss 0.003148f
C6086 FILLER_0_18_107/a_3172_472# vdd 0.004296f
C6087 net61 _418_/a_36_151# 0.042401f
C6088 net20 _419_/a_36_151# 0.001225f
C6089 _052_ vss 0.077815f
C6090 net78 _419_/a_796_472# 0.00376f
C6091 net61 _419_/a_1204_472# 0.012025f
C6092 net60 _419_/a_796_472# 0.003097f
C6093 net63 FILLER_0_20_193/a_124_375# 0.075841f
C6094 FILLER_0_24_130/a_36_472# vss 0.001687f
C6095 mask\[6\] vss 0.348967f
C6096 _417_/a_2665_112# _006_ 0.023025f
C6097 ctln[8] FILLER_0_0_96/a_36_472# 0.012298f
C6098 FILLER_0_11_109/a_36_472# _134_ 0.007739f
C6099 output31/a_224_472# _417_/a_36_151# 0.07368f
C6100 _088_ vss 0.326434f
C6101 FILLER_0_21_28/a_1380_472# _012_ 0.004453f
C6102 _010_ net19 0.408364f
C6103 FILLER_0_16_107/a_484_472# vdd 0.02929f
C6104 _119_ _322_/a_124_24# 0.020461f
C6105 net69 _154_ 0.05211f
C6106 net41 FILLER_0_19_28/a_484_472# 0.047447f
C6107 FILLER_0_6_79/a_36_472# vss 0.008693f
C6108 FILLER_0_12_136/a_1468_375# net23 0.021046f
C6109 net47 net6 0.23883f
C6110 FILLER_0_17_133/a_36_472# vdd 0.097394f
C6111 FILLER_0_17_133/a_124_375# vss 0.015434f
C6112 _076_ _226_/a_860_68# 0.001752f
C6113 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1468_375# 0.086742f
C6114 _308_/a_848_380# trim_mask\[0\] 0.035693f
C6115 _045_ _006_ 0.00216f
C6116 _372_/a_3662_472# _122_ 0.002653f
C6117 _074_ FILLER_0_5_172/a_36_472# 0.016713f
C6118 FILLER_0_14_81/a_36_472# _095_ 0.014706f
C6119 vdd _201_/a_67_603# 0.031337f
C6120 ctln[8] net15 0.205163f
C6121 net38 FILLER_0_20_2/a_572_375# 0.004413f
C6122 fanout61/a_36_113# net77 0.052643f
C6123 mask\[8\] mask\[9\] 0.078756f
C6124 net4 FILLER_0_12_220/a_36_472# 0.019348f
C6125 FILLER_0_8_107/a_36_472# vss 0.006371f
C6126 FILLER_0_18_107/a_3260_375# _145_ 0.00346f
C6127 net73 vdd 0.44835f
C6128 _423_/a_36_151# FILLER_0_23_44/a_572_375# 0.059049f
C6129 _091_ _323_/a_36_113# 0.001651f
C6130 _091_ fanout56/a_36_113# 0.001254f
C6131 _115_ _122_ 0.004082f
C6132 FILLER_0_22_177/a_36_472# _146_ 0.002f
C6133 _343_/a_49_472# net80 0.001646f
C6134 net16 FILLER_0_16_37/a_124_375# 0.033245f
C6135 _073_ net8 0.206839f
C6136 _430_/a_2248_156# mask\[3\] 0.004211f
C6137 _430_/a_2665_112# net20 0.005397f
C6138 _334_/a_36_160# FILLER_0_17_104/a_1468_375# 0.027706f
C6139 FILLER_0_18_177/a_3172_472# net22 0.037136f
C6140 _131_ _120_ 0.191602f
C6141 FILLER_0_5_54/a_572_375# trim_mask\[1\] 0.011664f
C6142 net34 net23 0.058486f
C6143 _449_/a_2560_156# vss 0.002544f
C6144 result[1] result[2] 0.072492f
C6145 net52 net49 0.092082f
C6146 mask\[9\] vss 0.649041f
C6147 mask\[8\] FILLER_0_22_86/a_1380_472# 0.012151f
C6148 net35 FILLER_0_22_86/a_932_472# 0.007806f
C6149 _105_ _009_ 0.01731f
C6150 net52 _442_/a_2248_156# 0.022954f
C6151 FILLER_0_9_28/a_484_472# _054_ 0.002831f
C6152 _139_ net21 0.004991f
C6153 net17 _452_/a_448_472# 0.043154f
C6154 _404_/a_36_472# _183_ 0.002637f
C6155 FILLER_0_17_72/a_1380_472# vdd 0.001762f
C6156 FILLER_0_17_72/a_932_472# vss 0.002754f
C6157 output32/a_224_472# output31/a_224_472# 0.00289f
C6158 _027_ FILLER_0_18_76/a_124_375# 0.001285f
C6159 FILLER_0_16_89/a_1380_472# net36 0.001657f
C6160 _360_/a_36_160# _160_ 0.052885f
C6161 net20 _420_/a_2248_156# 0.003737f
C6162 result[8] net21 0.166555f
C6163 FILLER_0_7_195/a_124_375# vdd 0.007788f
C6164 _131_ _403_/a_224_472# 0.003274f
C6165 _076_ FILLER_0_5_148/a_36_472# 0.011563f
C6166 net50 trim_mask\[1\] 0.502622f
C6167 _114_ _120_ 0.334426f
C6168 _164_ _160_ 1.863027f
C6169 _081_ _080_ 0.003905f
C6170 output25/a_224_472# _423_/a_2665_112# 0.001396f
C6171 _010_ _009_ 0.030637f
C6172 FILLER_0_24_130/a_124_375# ctlp[7] 0.002726f
C6173 _023_ vdd 0.062542f
C6174 FILLER_0_19_111/a_484_472# vdd 0.009246f
C6175 _013_ FILLER_0_18_53/a_572_375# 0.015534f
C6176 FILLER_0_19_187/a_572_375# vss 0.055266f
C6177 FILLER_0_19_187/a_36_472# vdd 0.09884f
C6178 FILLER_0_18_107/a_484_472# net14 0.002472f
C6179 FILLER_0_0_198/a_124_375# net11 0.071885f
C6180 output16/a_224_472# _447_/a_36_151# 0.200384f
C6181 net41 net49 0.392356f
C6182 FILLER_0_4_213/a_124_375# net59 0.039014f
C6183 _449_/a_2248_156# net15 0.001705f
C6184 net69 FILLER_0_3_78/a_484_472# 0.002068f
C6185 net14 FILLER_0_10_94/a_36_472# 0.003391f
C6186 _104_ fanout63/a_36_160# 0.007014f
C6187 net27 FILLER_0_12_236/a_36_472# 0.005414f
C6188 _065_ _036_ 0.031728f
C6189 net41 net68 0.009755f
C6190 _015_ FILLER_0_8_247/a_572_375# 0.00706f
C6191 net36 net62 0.034265f
C6192 _131_ FILLER_0_9_105/a_572_375# 0.031928f
C6193 net81 fanout79/a_36_160# 0.057526f
C6194 FILLER_0_17_72/a_36_472# net15 0.006905f
C6195 net17 FILLER_0_12_28/a_36_472# 0.012286f
C6196 ctln[3] ctln[4] 0.073214f
C6197 _093_ _438_/a_1000_472# 0.001556f
C6198 _176_ _394_/a_1936_472# 0.001255f
C6199 _078_ FILLER_0_3_221/a_124_375# 0.002694f
C6200 cal_count\[3\] _060_ 0.007037f
C6201 _098_ _434_/a_1308_423# 0.007057f
C6202 _079_ _260_/a_36_68# 0.043596f
C6203 _030_ _164_ 0.036025f
C6204 net53 _427_/a_1000_472# 0.008132f
C6205 FILLER_0_12_236/a_484_472# _060_ 0.002678f
C6206 net61 _422_/a_2560_156# 0.010748f
C6207 FILLER_0_18_2/a_124_375# vss 0.003207f
C6208 net3 _043_ 0.004313f
C6209 net20 _426_/a_2248_156# 0.007902f
C6210 FILLER_0_16_255/a_36_472# vdd 0.044615f
C6211 _136_ net14 0.417108f
C6212 _440_/a_1308_423# vss 0.028595f
C6213 FILLER_0_4_185/a_124_375# _272_/a_36_472# 0.001781f
C6214 _128_ _062_ 0.025708f
C6215 net34 net33 0.509436f
C6216 mask\[8\] _352_/a_49_472# 0.002573f
C6217 output29/a_224_472# output30/a_224_472# 0.005147f
C6218 _359_/a_1044_488# _152_ 0.001339f
C6219 _144_ mask\[7\] 0.111088f
C6220 _028_ FILLER_0_7_104/a_932_472# 0.003084f
C6221 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_124_375# 0.012221f
C6222 net80 _434_/a_36_151# 0.067037f
C6223 FILLER_0_16_89/a_36_472# _176_ 0.012173f
C6224 _091_ FILLER_0_13_212/a_124_375# 0.025558f
C6225 _412_/a_36_151# net75 0.060039f
C6226 net58 FILLER_0_8_263/a_124_375# 0.001876f
C6227 net34 _435_/a_1204_472# 0.004285f
C6228 mask\[8\] net35 2.631701f
C6229 output21/a_224_472# _104_ 0.002459f
C6230 net3 _185_ 0.004236f
C6231 _176_ _171_ 0.049997f
C6232 ctlp[6] net54 0.00409f
C6233 _144_ _148_ 0.038002f
C6234 net20 FILLER_0_3_221/a_1020_375# 0.025371f
C6235 FILLER_0_21_142/a_124_375# _140_ 0.016087f
C6236 net36 FILLER_0_15_235/a_572_375# 0.083299f
C6237 net1 net8 0.00497f
C6238 _035_ output41/a_224_472# 0.002168f
C6239 _059_ net23 0.265909f
C6240 FILLER_0_19_47/a_124_375# vdd 0.025971f
C6241 _402_/a_728_93# _179_ 0.011717f
C6242 _142_ vss 0.121933f
C6243 FILLER_0_14_91/a_124_375# en_co_clk 0.006788f
C6244 _174_ cal_count\[2\] 0.004821f
C6245 net63 _434_/a_1308_423# 0.003686f
C6246 _070_ net14 0.536953f
C6247 _132_ FILLER_0_18_107/a_1468_375# 0.089207f
C6248 _053_ FILLER_0_7_104/a_1020_375# 0.002671f
C6249 net55 _453_/a_2248_156# 0.001546f
C6250 _089_ FILLER_0_5_198/a_124_375# 0.001517f
C6251 _444_/a_2248_156# _054_ 0.002637f
C6252 mask\[5\] FILLER_0_20_177/a_124_375# 0.013531f
C6253 _356_/a_36_472# net14 0.001801f
C6254 FILLER_0_10_214/a_36_472# _247_/a_36_160# 0.004828f
C6255 FILLER_0_20_177/a_124_375# FILLER_0_20_169/a_124_375# 0.003732f
C6256 mask\[0\] FILLER_0_13_228/a_36_472# 0.002986f
C6257 net35 vss 0.434438f
C6258 FILLER_0_17_142/a_36_472# _137_ 0.003953f
C6259 mask\[3\] net22 0.036607f
C6260 net82 net21 0.037271f
C6261 _126_ _120_ 0.055349f
C6262 _130_ _120_ 0.014675f
C6263 result[6] net18 0.026875f
C6264 _423_/a_2248_156# _012_ 0.011646f
C6265 net15 _440_/a_36_151# 0.016061f
C6266 _088_ _269_/a_36_472# 0.004438f
C6267 _422_/a_2560_156# _108_ 0.008253f
C6268 net54 _150_ 0.001162f
C6269 _412_/a_1000_472# net1 0.027748f
C6270 FILLER_0_18_177/a_1828_472# FILLER_0_19_187/a_572_375# 0.001684f
C6271 _152_ FILLER_0_5_136/a_124_375# 0.039558f
C6272 _081_ FILLER_0_5_136/a_36_472# 0.0028f
C6273 FILLER_0_9_28/a_572_375# net16 0.042681f
C6274 FILLER_0_14_81/a_36_472# vss 0.007047f
C6275 FILLER_0_21_286/a_36_472# _420_/a_36_151# 0.059367f
C6276 _238_/a_67_603# vdd 0.004498f
C6277 _053_ net67 0.672744f
C6278 _077_ _410_/a_36_68# 0.020334f
C6279 net81 _283_/a_36_472# 0.032292f
C6280 FILLER_0_21_206/a_124_375# mask\[6\] 0.008881f
C6281 FILLER_0_22_86/a_1020_375# net14 0.047331f
C6282 _308_/a_124_24# FILLER_0_10_94/a_36_472# 0.001811f
C6283 _421_/a_36_151# net18 0.00659f
C6284 net79 FILLER_0_12_220/a_36_472# 0.005464f
C6285 FILLER_0_14_50/a_36_472# _095_ 0.013704f
C6286 FILLER_0_18_2/a_1468_375# _452_/a_448_472# 0.001597f
C6287 _365_/a_36_68# vss 0.029516f
C6288 _448_/a_1308_423# net59 0.014899f
C6289 _053_ _414_/a_796_472# 0.008213f
C6290 trim[4] _221_/a_36_160# 0.002685f
C6291 _345_/a_36_160# _098_ 0.002041f
C6292 _427_/a_36_151# vdd 0.107344f
C6293 FILLER_0_0_96/a_124_375# vss 0.008342f
C6294 FILLER_0_0_96/a_36_472# vdd 0.047982f
C6295 _256_/a_36_68# net22 0.019035f
C6296 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_124_375# 0.012222f
C6297 FILLER_0_7_72/a_36_472# vdd 0.106377f
C6298 FILLER_0_7_72/a_3260_375# vss 0.053035f
C6299 _016_ _131_ 0.017461f
C6300 _098_ _043_ 0.032706f
C6301 FILLER_0_18_76/a_484_472# _438_/a_36_151# 0.001723f
C6302 _287_/a_36_472# _006_ 0.00121f
C6303 output10/a_224_472# net58 0.025878f
C6304 vdd FILLER_0_5_148/a_572_375# -0.009701f
C6305 vss FILLER_0_5_148/a_124_375# 0.018465f
C6306 FILLER_0_9_28/a_124_375# vdd -0.004893f
C6307 net7 net68 0.032489f
C6308 cal_count\[3\] _095_ 0.06065f
C6309 mask\[5\] FILLER_0_19_171/a_1020_375# 0.007169f
C6310 ctln[2] clk 0.004558f
C6311 _443_/a_36_151# _081_ 0.001923f
C6312 FILLER_0_14_81/a_36_472# cal_count\[1\] 0.034486f
C6313 _437_/a_2248_156# net14 0.023718f
C6314 _264_/a_224_472# _084_ 0.007508f
C6315 _016_ _114_ 0.041462f
C6316 FILLER_0_13_212/a_1380_472# _043_ 0.014431f
C6317 fanout53/a_36_160# net36 0.028652f
C6318 _359_/a_36_488# _133_ 0.04287f
C6319 _072_ _116_ 0.283323f
C6320 _088_ FILLER_0_3_172/a_3172_472# 0.004381f
C6321 FILLER_0_22_177/a_124_375# net33 0.013581f
C6322 _087_ _163_ 0.004829f
C6323 FILLER_0_21_133/a_124_375# _098_ 0.006462f
C6324 net15 vdd 2.073988f
C6325 _104_ ctlp[2] 1.420577f
C6326 FILLER_0_17_38/a_36_472# _041_ 0.003805f
C6327 _180_ vdd 0.176915f
C6328 FILLER_0_13_65/a_124_375# net15 0.048002f
C6329 _077_ _120_ 0.205715f
C6330 _449_/a_2665_112# cal_count\[3\] 0.001422f
C6331 mask\[9\] _026_ 0.002924f
C6332 _444_/a_1000_472# net47 0.036015f
C6333 fanout51/a_36_113# vdd 0.013496f
C6334 _113_ FILLER_0_12_196/a_124_375# 0.001597f
C6335 _161_ _311_/a_66_473# 0.021817f
C6336 _090_ FILLER_0_12_196/a_36_472# 0.002321f
C6337 FILLER_0_22_177/a_484_472# _435_/a_36_151# 0.001723f
C6338 _120_ FILLER_0_10_107/a_124_375# 0.001834f
C6339 FILLER_0_19_155/a_124_375# vdd 0.019233f
C6340 _063_ _033_ 0.250192f
C6341 _442_/a_36_151# _031_ 0.013852f
C6342 net59 rstn 0.039664f
C6343 FILLER_0_3_172/a_36_472# FILLER_0_2_171/a_124_375# 0.001723f
C6344 _443_/a_36_151# FILLER_0_2_127/a_124_375# 0.073306f
C6345 net27 FILLER_0_9_290/a_36_472# 0.006729f
C6346 _410_/a_36_68# _453_/a_36_151# 0.002326f
C6347 _327_/a_36_472# FILLER_0_12_136/a_36_472# 0.096379f
C6348 ctln[5] FILLER_0_0_198/a_124_375# 0.002726f
C6349 _140_ _352_/a_665_69# 0.001363f
C6350 FILLER_0_15_205/a_124_375# net21 0.002912f
C6351 valid cal_itt\[1\] 0.011576f
C6352 _308_/a_124_24# _070_ 0.001465f
C6353 FILLER_0_3_142/a_124_375# _032_ 0.001153f
C6354 net58 FILLER_0_9_270/a_484_472# 0.061043f
C6355 _429_/a_36_151# FILLER_0_15_212/a_932_472# 0.001723f
C6356 state\[1\] _055_ 0.067603f
C6357 _414_/a_2560_156# vss 0.001078f
C6358 net34 FILLER_0_22_128/a_1828_472# 0.005158f
C6359 _098_ net21 0.133694f
C6360 _452_/a_3129_107# vdd 0.016611f
C6361 _162_ _374_/a_36_68# 0.005729f
C6362 FILLER_0_9_28/a_2724_472# _077_ 0.006001f
C6363 FILLER_0_3_54/a_124_375# net40 0.005766f
C6364 cal_itt\[2\] cal_itt\[1\] 0.057194f
C6365 _016_ _428_/a_2665_112# 0.050481f
C6366 net50 FILLER_0_5_72/a_1380_472# 0.002431f
C6367 trim_mask\[2\] FILLER_0_3_54/a_124_375# 0.015198f
C6368 net56 FILLER_0_17_142/a_36_472# 0.003603f
C6369 mask\[0\] _429_/a_1204_472# 0.005396f
C6370 output42/a_224_472# net47 0.083794f
C6371 _070_ FILLER_0_5_136/a_124_375# 0.001083f
C6372 net55 FILLER_0_18_53/a_484_472# 0.012319f
C6373 _321_/a_3126_472# _118_ 0.002754f
C6374 FILLER_0_18_177/a_2724_472# vdd 0.002749f
C6375 _065_ output15/a_224_472# 0.037721f
C6376 output8/a_224_472# net8 0.034396f
C6377 trimb[4] FILLER_0_15_2/a_124_375# 0.003305f
C6378 net72 FILLER_0_21_28/a_1468_375# 0.001823f
C6379 _412_/a_36_151# fanout81/a_36_160# 0.001725f
C6380 _068_ _163_ 0.04926f
C6381 FILLER_0_20_177/a_484_472# _098_ 0.009817f
C6382 net35 FILLER_0_22_128/a_1020_375# 0.010202f
C6383 _093_ FILLER_0_18_107/a_3172_472# 0.008787f
C6384 _044_ FILLER_0_13_290/a_36_472# 0.001194f
C6385 ctlp[7] vss 0.036681f
C6386 net47 _167_ 0.003019f
C6387 net75 _000_ 0.096899f
C6388 result[6] net62 0.005382f
C6389 _114_ FILLER_0_12_136/a_124_375# 0.006974f
C6390 net50 _054_ 0.131493f
C6391 _256_/a_36_68# _076_ 0.079206f
C6392 _256_/a_1612_497# _068_ 0.002759f
C6393 _376_/a_36_160# FILLER_0_6_90/a_124_375# 0.005705f
C6394 _120_ _453_/a_36_151# 0.001848f
C6395 _091_ _141_ 0.010074f
C6396 _042_ vss 0.008272f
C6397 net51 vdd 0.692054f
C6398 FILLER_0_10_78/a_572_375# FILLER_0_11_78/a_572_375# 0.05841f
C6399 ctlp[0] net43 0.003786f
C6400 FILLER_0_16_57/a_932_472# vdd 0.005518f
C6401 FILLER_0_16_57/a_484_472# vss 0.004107f
C6402 net63 net21 0.278824f
C6403 _176_ _183_ 0.024038f
C6404 net50 FILLER_0_8_24/a_36_472# 0.015187f
C6405 FILLER_0_18_107/a_3172_472# FILLER_0_19_134/a_124_375# 0.001723f
C6406 _427_/a_2665_112# state\[1\] 0.021573f
C6407 net73 _433_/a_36_151# 0.004541f
C6408 net57 _267_/a_1120_472# 0.002885f
C6409 net38 output6/a_224_472# 0.060017f
C6410 _260_/a_36_68# vss 0.030324f
C6411 FILLER_0_22_128/a_1468_375# vss 0.006619f
C6412 _093_ FILLER_0_17_133/a_36_472# 0.010432f
C6413 _432_/a_36_151# FILLER_0_16_154/a_1468_375# 0.001107f
C6414 net67 _164_ 0.030648f
C6415 _415_/a_1000_472# net18 0.006558f
C6416 FILLER_0_17_72/a_124_375# FILLER_0_15_72/a_36_472# 0.001512f
C6417 _414_/a_1204_472# cal_itt\[3\] 0.052432f
C6418 net64 FILLER_0_12_236/a_484_472# 0.010321f
C6419 _442_/a_36_151# _371_/a_36_113# 0.001089f
C6420 FILLER_0_9_28/a_2724_472# _453_/a_36_151# 0.013806f
C6421 net27 FILLER_0_10_247/a_36_472# 0.016681f
C6422 FILLER_0_15_290/a_36_472# net79 0.04083f
C6423 FILLER_0_2_93/a_36_472# net14 0.005108f
C6424 _016_ _126_ 0.051451f
C6425 FILLER_0_12_136/a_124_375# _428_/a_2665_112# 0.029834f
C6426 net63 FILLER_0_20_177/a_484_472# 0.002172f
C6427 net65 ctln[2] 0.113266f
C6428 _016_ _130_ 0.114514f
C6429 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2812_375# 0.001597f
C6430 net75 _253_/a_1732_68# 0.001047f
C6431 FILLER_0_17_133/a_36_472# FILLER_0_19_134/a_124_375# 0.001188f
C6432 _073_ FILLER_0_3_221/a_1020_375# 0.002563f
C6433 _140_ FILLER_0_19_155/a_572_375# 0.040109f
C6434 _217_/a_36_160# FILLER_0_19_28/a_572_375# 0.058908f
C6435 _095_ _278_/a_36_160# 0.030448f
C6436 _095_ FILLER_0_12_20/a_124_375# 0.001588f
C6437 FILLER_0_19_47/a_36_472# _013_ 0.03573f
C6438 output27/a_224_472# FILLER_0_9_270/a_572_375# 0.00135f
C6439 net73 _093_ 0.350073f
C6440 _408_/a_56_524# _190_/a_36_160# 0.004025f
C6441 _098_ FILLER_0_19_171/a_1380_472# 0.001764f
C6442 net16 _182_ 0.05291f
C6443 _367_/a_36_68# _157_ 0.013352f
C6444 _428_/a_448_472# _017_ 0.056f
C6445 _428_/a_36_151# net53 0.001124f
C6446 net41 _184_ 0.065857f
C6447 FILLER_0_21_28/a_1468_375# _424_/a_36_151# 0.059049f
C6448 FILLER_0_4_123/a_124_375# vdd 0.027816f
C6449 _077_ _227_/a_36_160# 0.012587f
C6450 FILLER_0_16_57/a_484_472# cal_count\[1\] 0.001664f
C6451 FILLER_0_16_57/a_1468_375# net15 0.012909f
C6452 _153_ FILLER_0_4_91/a_572_375# 0.001735f
C6453 net72 _401_/a_36_68# 0.006818f
C6454 FILLER_0_18_2/a_2364_375# net38 0.001683f
C6455 net63 FILLER_0_18_177/a_124_375# 0.001937f
C6456 FILLER_0_14_50/a_36_472# vss 0.002954f
C6457 FILLER_0_9_72/a_1020_375# vdd -0.014642f
C6458 FILLER_0_9_72/a_572_375# vss 0.007993f
C6459 _131_ _043_ 0.047425f
C6460 net82 FILLER_0_3_172/a_1468_375# 0.010439f
C6461 _086_ vss 0.615299f
C6462 _397_/a_36_472# FILLER_0_17_72/a_1020_375# 0.001781f
C6463 vdd _381_/a_36_472# 0.014305f
C6464 fanout75/a_36_113# _317_/a_36_113# 0.001442f
C6465 FILLER_0_4_144/a_124_375# _370_/a_848_380# 0.005599f
C6466 net75 FILLER_0_8_247/a_484_472# 0.003007f
C6467 _185_ _405_/a_67_603# 0.060789f
C6468 _093_ FILLER_0_17_72/a_1380_472# 0.008517f
C6469 mask\[4\] FILLER_0_18_209/a_36_472# 0.018888f
C6470 fanout63/a_36_160# mask\[2\] 0.026642f
C6471 net52 net47 0.039912f
C6472 _267_/a_36_472# _121_ 0.041237f
C6473 _394_/a_1336_472# _095_ 0.031869f
C6474 _137_ FILLER_0_16_154/a_124_375# 0.007998f
C6475 _028_ FILLER_0_7_72/a_572_375# 0.003837f
C6476 _173_ FILLER_0_12_28/a_124_375# 0.009218f
C6477 cal_count\[3\] vss 1.35143f
C6478 mask\[5\] net22 0.04021f
C6479 _147_ _023_ 0.004036f
C6480 FILLER_0_6_239/a_124_375# _123_ 0.044771f
C6481 net18 _417_/a_1308_423# 0.015651f
C6482 _114_ _043_ 0.071339f
C6483 _086_ net74 0.058077f
C6484 net63 FILLER_0_19_171/a_1380_472# 0.003014f
C6485 FILLER_0_12_236/a_484_472# vss 0.002739f
C6486 net75 _426_/a_1308_423# 0.002552f
C6487 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_36_472# 0.001963f
C6488 FILLER_0_21_206/a_36_472# vss 0.004971f
C6489 FILLER_0_16_89/a_1020_375# _136_ 0.019549f
C6490 net82 FILLER_0_3_221/a_932_472# 0.004092f
C6491 _089_ cal_itt\[3\] 0.049851f
C6492 result[6] _420_/a_1000_472# 0.007761f
C6493 FILLER_0_2_171/a_124_375# FILLER_0_2_165/a_124_375# 0.003598f
C6494 _328_/a_36_113# FILLER_0_11_109/a_36_472# 0.0161f
C6495 _093_ FILLER_0_19_111/a_484_472# 0.001009f
C6496 FILLER_0_18_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001597f
C6497 FILLER_0_4_49/a_484_472# _440_/a_36_151# 0.006095f
C6498 FILLER_0_12_136/a_124_375# _126_ 0.013041f
C6499 _098_ FILLER_0_15_212/a_1020_375# 0.00918f
C6500 _175_ _131_ 0.050098f
C6501 _291_/a_36_160# vdd 0.010802f
C6502 _154_ vss 0.200253f
C6503 _350_/a_665_69# net23 0.001468f
C6504 _130_ FILLER_0_12_136/a_124_375# 0.010514f
C6505 net57 _074_ 0.026184f
C6506 net39 FILLER_0_8_2/a_124_375# 0.008405f
C6507 FILLER_0_14_50/a_36_472# cal_count\[1\] 0.030015f
C6508 net74 cal_count\[3\] 0.040777f
C6509 _091_ FILLER_0_17_218/a_572_375# 0.001927f
C6510 net35 _211_/a_36_160# 0.009886f
C6511 net20 vdd 2.14128f
C6512 _443_/a_448_472# _032_ 0.036717f
C6513 _035_ _166_ 0.034749f
C6514 net82 _001_ 0.044461f
C6515 _316_/a_848_380# net37 0.01216f
C6516 _176_ FILLER_0_10_94/a_124_375# 0.009888f
C6517 _140_ FILLER_0_22_128/a_2364_375# 0.003037f
C6518 output33/a_224_472# _204_/a_67_603# 0.00401f
C6519 _096_ _055_ 0.047639f
C6520 _441_/a_36_151# FILLER_0_3_78/a_124_375# 0.035849f
C6521 ctlp[1] FILLER_0_21_286/a_124_375# 0.025059f
C6522 net41 net47 0.19549f
C6523 FILLER_0_3_221/a_124_375# FILLER_0_3_212/a_124_375# 0.002036f
C6524 net74 _154_ 0.002976f
C6525 _428_/a_2665_112# _043_ 0.021483f
C6526 net73 FILLER_0_17_142/a_124_375# 0.003021f
C6527 FILLER_0_21_28/a_1380_472# vdd 0.007073f
C6528 _052_ _424_/a_2560_156# 0.003401f
C6529 net23 _146_ 0.034955f
C6530 net75 _081_ 0.060976f
C6531 output48/a_224_472# net82 0.048965f
C6532 _053_ _059_ 0.042128f
C6533 _169_ vss 0.037006f
C6534 _163_ vdd 0.418075f
C6535 mask\[4\] FILLER_0_19_171/a_572_375# 0.006277f
C6536 trim_val\[4\] _241_/a_224_472# 0.003005f
C6537 _114_ net21 0.022033f
C6538 result[6] _421_/a_2248_156# 0.031832f
C6539 output43/a_224_472# trimb[2] 0.005445f
C6540 trimb[0] output45/a_224_472# 0.003753f
C6541 net63 FILLER_0_15_212/a_1020_375# 0.001012f
C6542 cal_itt\[1\] net59 0.227495f
C6543 _406_/a_36_159# net47 0.034933f
C6544 FILLER_0_13_142/a_1468_375# _225_/a_36_160# 0.027706f
C6545 FILLER_0_18_2/a_1380_472# net17 0.003603f
C6546 FILLER_0_4_107/a_572_375# _157_ 0.001032f
C6547 _112_ _425_/a_1204_472# 0.001132f
C6548 _173_ _039_ 0.0326f
C6549 result[8] _011_ 0.001294f
C6550 net68 trim_val\[0\] 0.052045f
C6551 net4 cal_itt\[1\] 0.048147f
C6552 FILLER_0_5_117/a_124_375# vdd 0.035079f
C6553 net81 _425_/a_448_472# 0.056225f
C6554 _181_ _402_/a_728_93# 0.064373f
C6555 _428_/a_36_151# FILLER_0_11_109/a_36_472# 0.001221f
C6556 _133_ _160_ 0.043549f
C6557 FILLER_0_4_49/a_36_472# vss 0.001931f
C6558 FILLER_0_4_49/a_484_472# vdd 0.003356f
C6559 net37 FILLER_0_5_148/a_484_472# 0.001212f
C6560 FILLER_0_19_195/a_124_375# FILLER_0_19_187/a_572_375# 0.012001f
C6561 mask\[9\] FILLER_0_18_76/a_124_375# 0.004592f
C6562 net76 FILLER_0_3_172/a_1380_472# 0.015215f
C6563 valid net59 0.577796f
C6564 _426_/a_36_151# FILLER_0_8_247/a_484_472# 0.001723f
C6565 net4 FILLER_0_7_233/a_36_472# 0.036721f
C6566 vss _433_/a_1308_423# 0.002695f
C6567 net56 FILLER_0_18_139/a_36_472# 0.002172f
C6568 FILLER_0_10_28/a_36_472# net47 0.002783f
C6569 output22/a_224_472# vdd 0.111234f
C6570 _428_/a_36_151# FILLER_0_14_107/a_36_472# 0.02628f
C6571 net26 _012_ 0.066032f
C6572 cal_itt\[2\] net59 0.014956f
C6573 FILLER_0_20_177/a_36_472# _434_/a_36_151# 0.001723f
C6574 FILLER_0_20_177/a_1468_375# _434_/a_448_472# 0.008952f
C6575 _350_/a_49_472# _049_ 0.025442f
C6576 cal_itt\[2\] net4 0.333682f
C6577 _126_ _043_ 0.128227f
C6578 net51 cal_count\[0\] 0.030963f
C6579 FILLER_0_21_142/a_484_472# net23 0.005353f
C6580 FILLER_0_3_78/a_484_472# vss 0.005811f
C6581 _190_/a_36_160# _043_ 0.06415f
C6582 _269_/a_36_472# _260_/a_36_68# 0.002875f
C6583 _265_/a_244_68# _082_ 0.031951f
C6584 mask\[3\] FILLER_0_18_177/a_932_472# 0.005654f
C6585 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_36_472# 0.002296f
C6586 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_36_472# 0.026657f
C6587 _187_ _186_ 0.032149f
C6588 FILLER_0_4_107/a_932_472# vdd 0.00987f
C6589 net15 FILLER_0_17_64/a_36_472# 0.015524f
C6590 _417_/a_1308_423# net62 0.006676f
C6591 _430_/a_36_151# _136_ 0.02044f
C6592 FILLER_0_2_171/a_124_375# net59 0.006603f
C6593 net67 _450_/a_1353_112# 0.025358f
C6594 FILLER_0_12_20/a_572_375# vdd 0.013384f
C6595 net24 FILLER_0_23_88/a_124_375# 0.020193f
C6596 FILLER_0_18_2/a_2364_375# net55 0.005899f
C6597 net48 _056_ 0.001581f
C6598 ctln[6] net69 0.003695f
C6599 _367_/a_692_472# net14 0.00423f
C6600 vdd FILLER_0_12_196/a_124_375# 0.015159f
C6601 net33 _146_ 0.306187f
C6602 output35/a_224_472# mask\[7\] 0.004608f
C6603 net27 _100_ 0.006783f
C6604 _105_ _106_ 0.038327f
C6605 _053_ FILLER_0_5_212/a_36_472# 0.007052f
C6606 result[1] net64 0.048458f
C6607 net70 FILLER_0_17_104/a_1020_375# 0.001894f
C6608 _050_ _140_ 0.001f
C6609 _053_ trim_val\[1\] 0.00385f
C6610 ctlp[7] _211_/a_36_160# 0.003488f
C6611 output37/a_224_472# net18 0.046654f
C6612 FILLER_0_17_200/a_124_375# net22 0.003602f
C6613 FILLER_0_5_128/a_36_472# _163_ 0.009857f
C6614 FILLER_0_19_171/a_932_472# _434_/a_36_151# 0.00271f
C6615 _136_ _333_/a_36_160# 0.00842f
C6616 _322_/a_848_380# _129_ 0.048486f
C6617 _119_ _086_ 0.419383f
C6618 ctlp[4] net21 0.04068f
C6619 _429_/a_36_151# FILLER_0_13_206/a_36_472# 0.059367f
C6620 _394_/a_728_93# vdd 0.006211f
C6621 _394_/a_1336_472# vss 0.040135f
C6622 _126_ net21 0.024842f
C6623 _142_ FILLER_0_17_142/a_572_375# 0.012321f
C6624 _429_/a_2665_112# net64 0.013014f
C6625 trim_mask\[4\] _160_ 0.244284f
C6626 net5 net18 0.015361f
C6627 FILLER_0_2_165/a_124_375# net59 0.00999f
C6628 net38 _444_/a_448_472# 0.031117f
C6629 FILLER_0_14_50/a_124_375# cal_count\[3\] 0.002524f
C6630 FILLER_0_21_125/a_36_472# _354_/a_49_472# 0.063744f
C6631 _093_ net15 0.145303f
C6632 _086_ FILLER_0_11_142/a_484_472# 0.008338f
C6633 FILLER_0_19_28/a_124_375# vdd 0.028695f
C6634 _076_ _223_/a_36_160# 0.001756f
C6635 FILLER_0_18_177/a_2812_375# _202_/a_36_160# 0.026361f
C6636 _429_/a_2665_112# mask\[1\] 0.001022f
C6637 FILLER_0_4_91/a_124_375# _160_ 0.009765f
C6638 _050_ FILLER_0_22_128/a_124_375# 0.002607f
C6639 _449_/a_2248_156# _067_ 0.040648f
C6640 FILLER_0_15_2/a_572_375# vdd 0.017581f
C6641 _093_ FILLER_0_19_155/a_124_375# 0.001864f
C6642 FILLER_0_15_2/a_124_375# vss 0.002713f
C6643 FILLER_0_9_223/a_124_375# net4 0.061757f
C6644 net31 FILLER_0_16_255/a_124_375# 0.029277f
C6645 _378_/a_224_472# net67 0.00211f
C6646 FILLER_0_12_2/a_572_375# vss 0.017629f
C6647 FILLER_0_12_2/a_36_472# vdd 0.104425f
C6648 trim_mask\[2\] net40 0.401672f
C6649 _081_ _265_/a_916_472# 0.002264f
C6650 _012_ FILLER_0_23_44/a_124_375# 0.002474f
C6651 _053_ FILLER_0_6_47/a_3260_375# 0.002746f
C6652 _436_/a_448_472# net35 0.012374f
C6653 FILLER_0_19_195/a_36_472# vss 0.005146f
C6654 net52 _453_/a_2665_112# 0.073881f
C6655 _417_/a_448_472# result[3] 0.003109f
C6656 FILLER_0_11_142/a_484_472# cal_count\[3\] 0.014314f
C6657 net80 mask\[6\] 0.080689f
C6658 FILLER_0_18_2/a_3260_375# net40 0.035372f
C6659 net16 _166_ 0.146913f
C6660 _363_/a_36_68# _153_ 0.008003f
C6661 _119_ _154_ 0.01697f
C6662 _447_/a_2665_112# _441_/a_36_151# 0.028591f
C6663 FILLER_0_13_80/a_124_375# FILLER_0_13_72/a_572_375# 0.012001f
C6664 _430_/a_448_472# _091_ 0.065306f
C6665 trim_val\[1\] FILLER_0_5_54/a_124_375# 0.001814f
C6666 _438_/a_36_151# _437_/a_36_151# 0.002668f
C6667 _118_ _121_ 0.02882f
C6668 net66 _440_/a_36_151# 0.041433f
C6669 FILLER_0_7_104/a_1468_375# _152_ 0.009263f
C6670 _104_ ctlp[1] 0.076863f
C6671 FILLER_0_15_150/a_36_472# net56 0.011741f
C6672 _394_/a_1336_472# cal_count\[1\] 0.018116f
C6673 net18 _418_/a_1308_423# 0.015651f
C6674 FILLER_0_17_142/a_36_472# vss 0.008239f
C6675 FILLER_0_17_142/a_484_472# vdd 0.004902f
C6676 ctln[5] output13/a_224_472# 0.023159f
C6677 output8/a_224_472# FILLER_0_3_221/a_1020_375# 0.03228f
C6678 result[1] vss 0.311464f
C6679 net17 _041_ 0.002779f
C6680 FILLER_0_5_172/a_36_472# _163_ 0.006934f
C6681 net18 _419_/a_2665_112# 0.0371f
C6682 _436_/a_796_472# vdd 0.005009f
C6683 output32/a_224_472# _419_/a_36_151# 0.129117f
C6684 net65 net21 0.04444f
C6685 _415_/a_36_151# net27 0.019856f
C6686 _127_ _428_/a_36_151# 0.030717f
C6687 ctlp[1] _420_/a_36_151# 0.067975f
C6688 _093_ FILLER_0_18_177/a_2724_472# 0.003036f
C6689 FILLER_0_4_197/a_1020_375# net59 0.008989f
C6690 _073_ vdd 0.258125f
C6691 net55 FILLER_0_21_60/a_572_375# 0.041903f
C6692 _430_/a_796_472# mask\[2\] 0.006305f
C6693 FILLER_0_18_76/a_36_472# vdd 0.014249f
C6694 FILLER_0_18_76/a_572_375# vss 0.007413f
C6695 FILLER_0_16_73/a_484_472# _131_ 0.007761f
C6696 _256_/a_36_68# _128_ 0.001702f
C6697 FILLER_0_21_142/a_124_375# _098_ 0.006558f
C6698 _429_/a_2665_112# vss 0.012165f
C6699 _077_ net21 0.032627f
C6700 _423_/a_2248_156# vdd 0.013707f
C6701 _432_/a_2560_156# _139_ 0.002737f
C6702 _137_ _043_ 0.007284f
C6703 FILLER_0_8_107/a_36_472# FILLER_0_9_105/a_124_375# 0.001684f
C6704 _414_/a_1308_423# net22 0.011978f
C6705 _341_/a_49_472# mask\[3\] 0.00631f
C6706 net20 net78 1.100401f
C6707 result[4] vdd 0.205815f
C6708 _136_ FILLER_0_16_154/a_36_472# 0.00615f
C6709 fanout69/a_36_113# _160_ 0.005933f
C6710 net20 net60 0.033919f
C6711 output39/a_224_472# _445_/a_36_151# 0.11862f
C6712 _078_ net37 0.459092f
C6713 FILLER_0_12_20/a_484_472# FILLER_0_12_28/a_36_472# 0.013277f
C6714 FILLER_0_1_266/a_572_375# net18 0.080358f
C6715 _008_ _418_/a_448_472# 0.052899f
C6716 net47 _450_/a_448_472# 0.012172f
C6717 _432_/a_2665_112# vss 0.002577f
C6718 net16 trim_mask\[1\] 0.007065f
C6719 FILLER_0_12_136/a_932_472# FILLER_0_13_142/a_124_375# 0.001684f
C6720 FILLER_0_9_270/a_124_375# vdd 0.013312f
C6721 net38 FILLER_0_20_15/a_124_375# 0.012947f
C6722 _053_ _385_/a_244_472# 0.00134f
C6723 net32 net30 0.004658f
C6724 _024_ _435_/a_1000_472# 0.002902f
C6725 _027_ _438_/a_1000_472# 0.010911f
C6726 net66 vdd 0.646189f
C6727 ctlp[1] _421_/a_1308_423# 0.002417f
C6728 _427_/a_1000_472# net23 0.003046f
C6729 _446_/a_1308_423# net17 0.033125f
C6730 FILLER_0_22_128/a_2724_472# FILLER_0_21_150/a_124_375# 0.001543f
C6731 _316_/a_848_380# _122_ 0.002234f
C6732 _316_/a_692_472# calibrate 0.006232f
C6733 _068_ _121_ 0.008802f
C6734 _345_/a_36_160# FILLER_0_19_125/a_36_472# 0.006647f
C6735 _415_/a_796_472# net81 0.002008f
C6736 net34 _109_ 0.001298f
C6737 _083_ _084_ 0.016693f
C6738 _445_/a_1308_423# vdd 0.001478f
C6739 _148_ mask\[7\] 0.010238f
C6740 fanout54/a_36_160# FILLER_0_19_142/a_124_375# 0.005489f
C6741 FILLER_0_18_177/a_2276_472# FILLER_0_19_195/a_124_375# 0.001684f
C6742 output36/a_224_472# net30 0.083671f
C6743 _414_/a_36_151# _079_ 0.037562f
C6744 net20 _256_/a_244_497# 0.005033f
C6745 trim_val\[1\] _164_ 0.100504f
C6746 FILLER_0_4_123/a_124_375# FILLER_0_4_107/a_1468_375# 0.012001f
C6747 FILLER_0_4_197/a_484_472# net76 0.003719f
C6748 FILLER_0_19_55/a_124_375# vdd 0.035786f
C6749 _029_ _365_/a_36_68# 0.013994f
C6750 _410_/a_36_68# vss 0.02717f
C6751 FILLER_0_20_87/a_124_375# net71 0.003629f
C6752 net74 _442_/a_1308_423# 0.001618f
C6753 net4 net59 0.102012f
C6754 _214_/a_36_160# _051_ 0.207388f
C6755 FILLER_0_2_93/a_36_472# net49 0.001451f
C6756 FILLER_0_15_282/a_484_472# _417_/a_36_151# 0.059367f
C6757 FILLER_0_15_282/a_36_472# _417_/a_448_472# 0.011962f
C6758 _086_ _321_/a_2034_472# 0.001815f
C6759 net75 FILLER_0_10_256/a_124_375# 0.027258f
C6760 FILLER_0_7_104/a_1020_375# _133_ 0.008772f
C6761 _085_ _161_ 0.008926f
C6762 state\[2\] _225_/a_36_160# 0.037565f
C6763 _069_ FILLER_0_15_212/a_36_472# 0.046864f
C6764 _372_/a_170_472# _062_ 0.014919f
C6765 _131_ _062_ 0.120189f
C6766 net36 net71 0.148833f
C6767 _425_/a_36_151# vdd 0.078723f
C6768 _077_ _453_/a_796_472# 0.003409f
C6769 net41 _402_/a_718_527# 0.019628f
C6770 net15 _424_/a_2665_112# 0.046592f
C6771 _129_ _124_ 0.010499f
C6772 output10/a_224_472# net9 0.003212f
C6773 _089_ _081_ 0.002206f
C6774 mask\[7\] _435_/a_796_472# 0.009587f
C6775 net63 FILLER_0_19_187/a_484_472# 0.020823f
C6776 _053_ net48 0.003159f
C6777 FILLER_0_18_107/a_124_375# mask\[9\] 0.006029f
C6778 _447_/a_2560_156# net15 0.001586f
C6779 result[7] _421_/a_1000_472# 0.015328f
C6780 _067_ vdd 0.853589f
C6781 _390_/a_36_68# _038_ 0.019355f
C6782 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_124_375# 0.016748f
C6783 FILLER_0_13_65/a_124_375# _067_ 0.001283f
C6784 _114_ _062_ 0.028432f
C6785 FILLER_0_11_124/a_124_375# _118_ 0.030768f
C6786 FILLER_0_17_282/a_124_375# net30 0.001288f
C6787 _144_ FILLER_0_21_125/a_36_472# 0.008287f
C6788 FILLER_0_5_128/a_124_375# _160_ 0.001157f
C6789 _115_ _118_ 1.045555f
C6790 output45/a_224_472# net43 0.024629f
C6791 FILLER_0_20_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001543f
C6792 net1 vdd 0.63891f
C6793 _420_/a_36_151# FILLER_0_23_282/a_124_375# 0.059049f
C6794 _291_/a_36_160# _093_ 0.017281f
C6795 FILLER_0_14_99/a_124_375# vdd 0.040312f
C6796 net20 FILLER_0_13_228/a_36_472# 0.020589f
C6797 _016_ _095_ 0.034744f
C6798 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_36_472# 0.001723f
C6799 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_572_375# 0.026339f
C6800 _120_ vss 0.42505f
C6801 _408_/a_56_524# _095_ 0.01643f
C6802 mask\[5\] _140_ 0.103728f
C6803 net54 vdd 0.877573f
C6804 FILLER_0_20_169/a_124_375# _140_ 0.01799f
C6805 net20 _093_ 0.398457f
C6806 mask\[2\] FILLER_0_16_154/a_1380_472# 0.017868f
C6807 _056_ _311_/a_66_473# 0.026074f
C6808 FILLER_0_13_142/a_932_472# _043_ 0.011974f
C6809 _053_ FILLER_0_6_177/a_124_375# 0.009352f
C6810 result[6] result[9] 0.026511f
C6811 net41 output38/a_224_472# 0.017358f
C6812 _089_ _270_/a_36_472# 0.00437f
C6813 net46 net40 0.254778f
C6814 net17 FILLER_0_20_15/a_932_472# 0.047256f
C6815 _152_ net47 0.242864f
C6816 FILLER_0_15_150/a_36_472# _095_ 0.001526f
C6817 _168_ _164_ 0.092012f
C6818 net41 FILLER_0_21_28/a_572_375# 0.054443f
C6819 _013_ net36 0.032392f
C6820 net74 _120_ 0.027885f
C6821 _434_/a_448_472# mask\[6\] 0.060756f
C6822 fanout68/a_36_113# _441_/a_36_151# 0.138322f
C6823 net80 net35 0.028982f
C6824 net79 _416_/a_36_151# 0.062626f
C6825 ctlp[1] FILLER_0_24_274/a_932_472# 0.003603f
C6826 _094_ mask\[1\] 0.49634f
C6827 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1468_375# 0.086742f
C6828 _009_ _107_ 0.027726f
C6829 output36/a_224_472# FILLER_0_15_282/a_124_375# 0.002977f
C6830 _307_/a_234_472# _126_ 0.00204f
C6831 ctlp[3] _422_/a_2248_156# 0.001888f
C6832 cal_count\[3\] _389_/a_36_148# 0.024777f
C6833 FILLER_0_5_117/a_36_472# FILLER_0_4_107/a_1020_375# 0.001684f
C6834 _444_/a_796_472# net40 0.005776f
C6835 FILLER_0_20_193/a_572_375# vdd 0.029393f
C6836 _064_ _444_/a_36_151# 0.001296f
C6837 fanout54/a_36_160# FILLER_0_19_155/a_36_472# 0.193804f
C6838 FILLER_0_10_256/a_124_375# _426_/a_36_151# 0.001597f
C6839 FILLER_0_16_73/a_124_375# _175_ 0.005727f
C6840 _439_/a_2665_112# net14 0.004943f
C6841 FILLER_0_17_72/a_1828_472# _131_ 0.004882f
C6842 FILLER_0_9_105/a_36_472# vdd 0.009746f
C6843 FILLER_0_9_105/a_572_375# vss 0.020145f
C6844 _410_/a_244_472# _042_ 0.003902f
C6845 _127_ _085_ 0.00179f
C6846 FILLER_0_5_198/a_124_375# net59 0.00174f
C6847 _115_ _068_ 0.889978f
C6848 net20 output11/a_224_472# 0.036556f
C6849 net70 _136_ 0.032219f
C6850 net40 trim[3] 0.084824f
C6851 FILLER_0_18_139/a_36_472# vss 0.007877f
C6852 FILLER_0_18_139/a_484_472# vdd 0.003106f
C6853 _258_/a_36_160# _079_ 0.026618f
C6854 net65 result[0] 0.011634f
C6855 FILLER_0_16_154/a_572_375# vdd 0.004706f
C6856 FILLER_0_16_154/a_124_375# vss 0.004317f
C6857 _412_/a_36_151# cal_itt\[1\] 0.025078f
C6858 _121_ vdd 0.106437f
C6859 net15 FILLER_0_17_56/a_484_472# 0.001758f
C6860 _374_/a_36_68# _058_ 0.010442f
C6861 _091_ FILLER_0_12_220/a_36_472# 0.003655f
C6862 net19 _420_/a_448_472# 0.05745f
C6863 _094_ vss 0.24519f
C6864 _036_ FILLER_0_3_54/a_36_472# 0.002156f
C6865 net2 _425_/a_36_151# 0.012359f
C6866 _370_/a_848_380# vss 0.051599f
C6867 mask\[7\] FILLER_0_22_128/a_932_472# 0.017448f
C6868 _367_/a_36_68# _160_ 0.013113f
C6869 FILLER_0_8_127/a_36_472# _058_ 0.003283f
C6870 net55 FILLER_0_21_28/a_3172_472# 0.06297f
C6871 _202_/a_36_160# _047_ 0.02265f
C6872 _415_/a_448_472# net64 0.02484f
C6873 FILLER_0_15_116/a_36_472# _451_/a_36_151# 0.096503f
C6874 _060_ net21 0.074356f
C6875 _320_/a_1568_472# state\[1\] 0.001531f
C6876 _412_/a_36_151# valid 0.009757f
C6877 FILLER_0_7_104/a_124_375# vdd 0.031505f
C6878 _101_ _045_ 0.001111f
C6879 _070_ net47 0.071795f
C6880 ctln[2] vss 0.256543f
C6881 _085_ _071_ 0.127349f
C6882 net68 FILLER_0_6_47/a_1828_472# 0.009096f
C6883 _227_/a_36_160# vss 0.010455f
C6884 net74 _370_/a_848_380# 0.004546f
C6885 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_484_472# 0.013276f
C6886 net38 _034_ 0.025823f
C6887 FILLER_0_18_107/a_1020_375# vdd -0.008765f
C6888 _434_/a_36_151# _023_ 0.035162f
C6889 _413_/a_36_151# vdd 0.130213f
C6890 net1 net2 0.624657f
C6891 trim_mask\[1\] FILLER_0_6_47/a_2724_472# 0.003645f
C6892 _161_ _310_/a_49_472# 0.022411f
C6893 output28/a_224_472# FILLER_0_11_282/a_36_472# 0.008834f
C6894 FILLER_0_19_187/a_36_472# _434_/a_36_151# 0.002398f
C6895 net79 net4 0.386068f
C6896 _049_ FILLER_0_22_128/a_2812_375# 0.001905f
C6897 result[4] net60 0.244453f
C6898 _431_/a_36_151# _131_ 0.03645f
C6899 net54 FILLER_0_22_128/a_572_375# 0.048634f
C6900 net19 _082_ 0.029316f
C6901 FILLER_0_16_89/a_36_472# _451_/a_2225_156# 0.001329f
C6902 result[9] FILLER_0_24_274/a_36_472# 0.009425f
C6903 mask\[3\] FILLER_0_17_161/a_124_375# 0.032905f
C6904 output8/a_224_472# vdd 0.023187f
C6905 net76 FILLER_0_5_198/a_484_472# 0.00169f
C6906 _141_ net23 0.782974f
C6907 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_36_472# 0.016748f
C6908 FILLER_0_21_28/a_2276_472# _423_/a_448_472# 0.008036f
C6909 _144_ _354_/a_665_69# 0.001518f
C6910 _421_/a_796_472# net19 0.009462f
C6911 _030_ _367_/a_36_68# 0.015584f
C6912 net37 _160_ 0.003563f
C6913 FILLER_0_9_28/a_2276_472# _042_ 0.002496f
C6914 FILLER_0_9_28/a_1828_472# net51 0.001502f
C6915 FILLER_0_20_15/a_1020_375# net40 0.005742f
C6916 _446_/a_2665_112# vdd 0.044081f
C6917 _421_/a_2665_112# _419_/a_2248_156# 0.001545f
C6918 output21/a_224_472# output35/a_224_472# 0.001374f
C6919 net65 output48/a_224_472# 0.015306f
C6920 _414_/a_36_151# vss 0.002101f
C6921 _414_/a_448_472# vdd 0.013377f
C6922 FILLER_0_22_86/a_36_472# _437_/a_36_151# 0.059367f
C6923 net69 _384_/a_224_472# 0.002407f
C6924 FILLER_0_5_72/a_484_472# vss 0.003738f
C6925 FILLER_0_5_72/a_932_472# vdd 0.002735f
C6926 FILLER_0_5_164/a_572_375# _386_/a_848_380# 0.001121f
C6927 _319_/a_672_472# _125_ 0.002725f
C6928 _128_ _223_/a_36_160# 0.012824f
C6929 FILLER_0_12_136/a_1468_375# state\[2\] 0.035275f
C6930 net16 _054_ 0.044357f
C6931 output9/a_224_472# net76 0.002042f
C6932 _432_/a_2560_156# net63 0.00227f
C6933 trim_val\[3\] _168_ 0.271475f
C6934 _303_/a_36_472# _098_ 0.021192f
C6935 _091_ mask\[2\] 2.252217f
C6936 _308_/a_124_24# _439_/a_2665_112# 0.002245f
C6937 net16 cal_count\[2\] 0.041089f
C6938 _029_ _154_ 0.116532f
C6939 FILLER_0_9_28/a_1468_375# _444_/a_2248_156# 0.001074f
C6940 _078_ _122_ 0.185069f
C6941 _083_ calibrate 0.001446f
C6942 _095_ _043_ 2.807456f
C6943 _077_ _062_ 0.037598f
C6944 _323_/a_36_113# _015_ 0.003795f
C6945 _449_/a_36_151# FILLER_0_12_50/a_124_375# 0.017882f
C6946 _016_ vss 0.069165f
C6947 result[7] ctlp[1] 0.07619f
C6948 _415_/a_1308_423# vdd 0.004258f
C6949 _124_ FILLER_0_10_107/a_572_375# 0.002135f
C6950 net41 net72 0.319547f
C6951 net53 mask\[2\] 0.005907f
C6952 _067_ cal_count\[0\] 0.201595f
C6953 net38 _445_/a_2248_156# 0.029721f
C6954 net16 FILLER_0_8_37/a_124_375# 0.010358f
C6955 _095_ _185_ 0.034457f
C6956 _079_ net21 0.065561f
C6957 _119_ _120_ 0.036534f
C6958 _420_/a_448_472# _009_ 0.061681f
C6959 net74 _390_/a_244_472# 0.001317f
C6960 _411_/a_36_151# FILLER_0_0_232/a_124_375# 0.059049f
C6961 _176_ _451_/a_2225_156# 0.030788f
C6962 ctln[7] _442_/a_2560_156# 0.001742f
C6963 _072_ _247_/a_36_160# 0.005008f
C6964 _093_ FILLER_0_17_142/a_484_472# 0.011974f
C6965 FILLER_0_15_150/a_36_472# vss 0.00975f
C6966 _286_/a_224_472# vdd 0.00154f
C6967 fanout72/a_36_113# _449_/a_36_151# 0.032681f
C6968 FILLER_0_6_90/a_572_375# _439_/a_2665_112# 0.001646f
C6969 FILLER_0_8_24/a_572_375# vdd 0.011353f
C6970 _016_ net74 0.568682f
C6971 _443_/a_36_151# net23 0.012359f
C6972 FILLER_0_5_54/a_1380_472# _440_/a_36_151# 0.001723f
C6973 FILLER_0_11_142/a_484_472# _120_ 0.007893f
C6974 FILLER_0_17_72/a_1380_472# _027_ 0.00378f
C6975 FILLER_0_17_72/a_2276_472# _150_ 0.003968f
C6976 net50 _441_/a_1308_423# 0.032656f
C6977 net52 _441_/a_1000_472# 0.011506f
C6978 _175_ _095_ 0.041931f
C6979 FILLER_0_12_220/a_124_375# vdd -0.008946f
C6980 FILLER_0_4_49/a_124_375# net66 0.017584f
C6981 FILLER_0_13_212/a_1020_375# net79 0.009597f
C6982 _176_ fanout55/a_36_160# 0.070942f
C6983 ctln[6] vss 0.45431f
C6984 net23 _433_/a_2665_112# 0.015555f
C6985 FILLER_0_4_107/a_572_375# _160_ 0.008945f
C6986 net26 vdd 0.487733f
C6987 _155_ vdd 0.193832f
C6988 state\[0\] _223_/a_36_160# 0.070065f
C6989 _093_ FILLER_0_18_76/a_36_472# 0.129892f
C6990 _345_/a_36_160# FILLER_0_19_111/a_572_375# 0.132282f
C6991 FILLER_0_11_124/a_124_375# vdd 0.016626f
C6992 _176_ _401_/a_36_68# 0.004263f
C6993 net52 _440_/a_2560_156# 0.004924f
C6994 FILLER_0_23_274/a_36_472# vss 0.002346f
C6995 output29/a_224_472# _416_/a_36_151# 0.07368f
C6996 fanout74/a_36_113# _443_/a_36_151# 0.032681f
C6997 net50 _439_/a_448_472# 0.020872f
C6998 net52 _439_/a_796_472# 0.003099f
C6999 _115_ vdd 0.455713f
C7000 output44/a_224_472# FILLER_0_18_2/a_1916_375# 0.032639f
C7001 _053_ FILLER_0_7_72/a_1828_472# 0.013271f
C7002 _425_/a_1308_423# net37 0.002601f
C7003 mask\[4\] FILLER_0_18_177/a_484_472# 0.016924f
C7004 output36/a_224_472# _417_/a_2665_112# 0.008243f
C7005 net29 _006_ 0.135646f
C7006 _063_ _166_ 0.025402f
C7007 _110_ net36 0.002287f
C7008 FILLER_0_6_239/a_124_375# _074_ 0.010359f
C7009 net41 _424_/a_36_151# 0.00413f
C7010 FILLER_0_12_136/a_124_375# vss 0.004063f
C7011 FILLER_0_12_136/a_572_375# vdd 0.016972f
C7012 _417_/a_36_151# vdd 0.140703f
C7013 ctln[1] net19 0.001327f
C7014 _133_ _059_ 0.039848f
C7015 net69 FILLER_0_2_111/a_36_472# 0.010759f
C7016 _031_ FILLER_0_2_111/a_1020_375# 0.016661f
C7017 _065_ trim_val\[2\] 0.002278f
C7018 FILLER_0_12_124/a_36_472# _017_ 0.004641f
C7019 ctln[4] FILLER_0_0_198/a_36_472# 0.02582f
C7020 net27 mask\[0\] 0.067038f
C7021 result[8] output19/a_224_472# 0.001465f
C7022 output35/a_224_472# ctlp[2] 0.001465f
C7023 result[6] net61 0.120359f
C7024 _000_ cal_itt\[1\] 0.012692f
C7025 _178_ _402_/a_2172_497# 0.003871f
C7026 _008_ _006_ 0.02963f
C7027 _065_ _447_/a_796_472# 0.007495f
C7028 output36/a_224_472# _045_ 0.041236f
C7029 mask\[3\] _098_ 0.026156f
C7030 FILLER_0_5_54/a_932_472# vss 0.003426f
C7031 FILLER_0_5_54/a_1380_472# vdd 0.008983f
C7032 cal_count\[2\] _452_/a_1353_112# 0.002558f
C7033 _105_ _422_/a_36_151# 0.030571f
C7034 _072_ net48 0.037795f
C7035 _254_/a_448_472# net22 0.009088f
C7036 _195_/a_67_603# vdd 0.022493f
C7037 net64 _043_ 0.004021f
C7038 ctln[1] input2/a_36_113# 0.05197f
C7039 _424_/a_36_151# FILLER_0_18_37/a_572_375# 0.002807f
C7040 net57 _163_ 0.759175f
C7041 _096_ _320_/a_1568_472# 0.001632f
C7042 net73 FILLER_0_17_104/a_1380_472# 0.003206f
C7043 FILLER_0_14_91/a_484_472# _136_ 0.038919f
C7044 _432_/a_2665_112# _019_ 0.002852f
C7045 mask\[1\] _043_ 0.027561f
C7046 _101_ _285_/a_244_68# 0.001153f
C7047 mask\[5\] result[8] 0.003797f
C7048 result[2] _044_ 0.393081f
C7049 _256_/a_2960_68# _056_ 0.001168f
C7050 FILLER_0_15_212/a_36_472# net22 0.003143f
C7051 valid _425_/a_2248_156# 0.00154f
C7052 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_124_375# 0.004426f
C7053 _440_/a_2665_112# _164_ 0.067034f
C7054 cal_itt\[2\] _000_ 0.042235f
C7055 net44 net6 0.005889f
C7056 output21/a_224_472# mask\[7\] 0.032297f
C7057 _258_/a_36_160# vss 0.005039f
C7058 _151_ vss 0.050544f
C7059 _322_/a_1152_472# _118_ 0.001235f
C7060 _322_/a_124_24# _124_ 0.041337f
C7061 output34/a_224_472# vss 0.011966f
C7062 en net18 0.32189f
C7063 _363_/a_36_68# FILLER_0_7_104/a_572_375# 0.002308f
C7064 _422_/a_36_151# _010_ 0.006787f
C7065 net16 FILLER_0_17_38/a_484_472# 0.032356f
C7066 trimb[1] vss 0.048527f
C7067 _233_/a_36_160# _445_/a_2248_156# 0.00136f
C7068 _253_/a_1732_68# cal_itt\[1\] 0.001829f
C7069 _063_ trim_mask\[1\] 0.127216f
C7070 net54 _433_/a_36_151# 0.00661f
C7071 net81 FILLER_0_15_212/a_36_472# 0.003945f
C7072 FILLER_0_7_72/a_1380_472# net50 0.077411f
C7073 result[7] FILLER_0_23_282/a_124_375# 0.016009f
C7074 FILLER_0_2_177/a_36_472# net59 0.007582f
C7075 _100_ FILLER_0_12_236/a_484_472# 0.00195f
C7076 _119_ _227_/a_36_160# 0.01123f
C7077 FILLER_0_10_28/a_124_375# net40 0.047331f
C7078 _165_ _033_ 0.022734f
C7079 _431_/a_36_151# FILLER_0_15_116/a_572_375# 0.001543f
C7080 net70 FILLER_0_14_107/a_484_472# 0.010987f
C7081 net63 mask\[3\] 0.37365f
C7082 _053_ FILLER_0_7_59/a_36_472# 0.073877f
C7083 FILLER_0_14_91/a_484_472# _070_ 0.001773f
C7084 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1468_375# 0.086635f
C7085 ctln[5] net22 0.072969f
C7086 cal_itt\[3\] net59 0.018616f
C7087 FILLER_0_8_263/a_124_375# calibrate 0.006928f
C7088 _070_ state\[1\] 0.032046f
C7089 FILLER_0_19_47/a_484_472# FILLER_0_18_37/a_1468_375# 0.001684f
C7090 _412_/a_36_151# net59 0.003938f
C7091 FILLER_0_4_177/a_572_375# net76 0.009573f
C7092 output32/a_224_472# vdd 0.082664f
C7093 _103_ _094_ 0.280781f
C7094 FILLER_0_16_57/a_1380_472# _131_ 0.008223f
C7095 fanout73/a_36_113# net53 0.047141f
C7096 ctlp[8] mask\[8\] 0.001554f
C7097 FILLER_0_17_38/a_572_375# vss 0.007503f
C7098 FILLER_0_17_38/a_36_472# vdd 0.01637f
C7099 FILLER_0_5_109/a_484_472# net47 0.002299f
C7100 net46 FILLER_0_20_15/a_1020_375# 0.0302f
C7101 trimb[3] FILLER_0_20_15/a_124_375# 0.001391f
C7102 _321_/a_2034_472# _120_ 0.002489f
C7103 _345_/a_36_160# vss 0.003697f
C7104 trim_val\[4\] _443_/a_36_151# 0.009986f
C7105 cal_itt\[0\] _082_ 0.018597f
C7106 _098_ _433_/a_1000_472# 0.0184f
C7107 FILLER_0_18_2/a_36_472# net44 0.011079f
C7108 output37/a_224_472# fanout59/a_36_160# 0.021845f
C7109 _093_ net54 0.003211f
C7110 mask\[1\] net21 0.023956f
C7111 _104_ _199_/a_36_160# 0.095519f
C7112 _340_/a_36_160# _140_ 0.062613f
C7113 _043_ vss 1.362912f
C7114 FILLER_0_13_65/a_36_472# _043_ 0.013651f
C7115 net34 FILLER_0_22_177/a_932_472# 0.003953f
C7116 _091_ _339_/a_36_160# 0.031941f
C7117 net47 _452_/a_36_151# 0.021978f
C7118 _367_/a_36_68# _156_ 0.096366f
C7119 _307_/a_672_472# _113_ 0.006607f
C7120 mask\[9\] _438_/a_1000_472# 0.056239f
C7121 fanout59/a_36_160# net5 0.05829f
C7122 _121_ _314_/a_224_472# 0.00323f
C7123 FILLER_0_3_172/a_2364_375# net22 0.013028f
C7124 ctlp[8] vss 0.107975f
C7125 FILLER_0_18_171/a_36_472# mask\[3\] 0.00262f
C7126 net54 FILLER_0_19_134/a_124_375# 0.002681f
C7127 FILLER_0_17_72/a_2724_472# _438_/a_36_151# 0.002529f
C7128 comp FILLER_0_15_2/a_124_375# 0.034135f
C7129 _185_ vss 0.021437f
C7130 _285_/a_36_472# mask\[2\] 0.002447f
C7131 _429_/a_448_472# _018_ 0.035489f
C7132 _346_/a_49_472# mask\[5\] 0.037629f
C7133 _085_ net23 0.020463f
C7134 net74 _043_ 0.65119f
C7135 _424_/a_2665_112# _423_/a_2248_156# 0.001314f
C7136 output7/a_224_472# trim[2] 0.008581f
C7137 ctln[0] output40/a_224_472# 0.017541f
C7138 FILLER_0_15_142/a_484_472# _427_/a_36_151# 0.001723f
C7139 FILLER_0_14_81/a_124_375# _175_ 0.005719f
C7140 FILLER_0_21_133/a_36_472# vdd 0.092168f
C7141 FILLER_0_21_133/a_124_375# vss 0.015693f
C7142 _322_/a_1152_472# _068_ 0.001502f
C7143 _175_ vss 0.162988f
C7144 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_36_472# 0.009654f
C7145 cal_count\[3\] _408_/a_728_93# 0.040643f
C7146 _413_/a_36_151# FILLER_0_3_172/a_2724_472# 0.001723f
C7147 FILLER_0_10_78/a_1380_472# _308_/a_124_24# 0.037778f
C7148 _411_/a_2665_112# _073_ 0.009313f
C7149 net50 FILLER_0_7_59/a_572_375# 0.009554f
C7150 cal_count\[1\] _043_ 0.002223f
C7151 net44 FILLER_0_15_10/a_124_375# 0.009108f
C7152 _062_ _060_ 0.032472f
C7153 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_36_472# 0.012267f
C7154 ctln[7] output15/a_224_472# 0.00838f
C7155 _265_/a_244_68# cal_itt\[0\] 0.003127f
C7156 ctlp[2] mask\[7\] 0.036719f
C7157 output44/a_224_472# output46/a_224_472# 0.005749f
C7158 _131_ _182_ 0.113302f
C7159 _053_ _028_ 0.891578f
C7160 _087_ FILLER_0_3_172/a_1916_375# 0.001223f
C7161 net21 vss 1.123312f
C7162 _261_/a_36_160# vss 0.05095f
C7163 _081_ cal_itt\[1\] 0.009747f
C7164 _431_/a_36_151# _137_ 0.011412f
C7165 _233_/a_36_160# FILLER_0_6_37/a_124_375# 0.001713f
C7166 net50 net14 0.192231f
C7167 _064_ net49 0.377675f
C7168 _122_ _160_ 0.004488f
C7169 FILLER_0_19_47/a_36_472# _012_ 0.001667f
C7170 FILLER_0_17_200/a_484_472# _069_ 0.001396f
C7171 _006_ result[3] 0.016909f
C7172 _053_ _359_/a_1492_488# 0.001437f
C7173 _185_ cal_count\[1\] 0.001949f
C7174 _430_/a_1308_423# _429_/a_36_151# 0.001722f
C7175 net69 _441_/a_36_151# 0.035817f
C7176 _120_ _389_/a_36_148# 0.022887f
C7177 net52 FILLER_0_3_142/a_124_375# 0.002239f
C7178 FILLER_0_10_107/a_484_472# vss 0.00298f
C7179 _093_ FILLER_0_18_139/a_484_472# 0.008683f
C7180 _447_/a_2248_156# _030_ 0.001588f
C7181 _064_ net68 0.059889f
C7182 trim_val\[2\] _036_ 0.279133f
C7183 _321_/a_170_472# _121_ 0.007364f
C7184 _176_ _055_ 0.001694f
C7185 net71 _437_/a_448_472# 0.060858f
C7186 FILLER_0_12_136/a_484_472# _127_ 0.005549f
C7187 net41 _407_/a_36_472# 0.003257f
C7188 FILLER_0_15_235/a_36_472# FILLER_0_15_228/a_36_472# 0.002765f
C7189 _447_/a_796_472# _036_ 0.006511f
C7190 _064_ _445_/a_1204_472# 0.007445f
C7191 _306_/a_36_68# _055_ 0.006686f
C7192 FILLER_0_7_72/a_484_472# _077_ 0.001332f
C7193 result[5] net19 0.003542f
C7194 _175_ cal_count\[1\] 0.203153f
C7195 _088_ FILLER_0_3_221/a_484_472# 0.002245f
C7196 FILLER_0_20_177/a_932_472# vdd 0.035019f
C7197 FILLER_0_20_177/a_484_472# vss 0.001256f
C7198 _436_/a_36_151# net54 0.004179f
C7199 _091_ FILLER_0_15_212/a_1380_472# 0.002787f
C7200 _232_/a_67_603# vdd 0.007565f
C7201 FILLER_0_14_263/a_36_472# vdd 0.02759f
C7202 FILLER_0_14_263/a_124_375# vss 0.007923f
C7203 _002_ net22 0.038848f
C7204 cal_itt\[2\] _081_ 0.003204f
C7205 _450_/a_1353_112# output6/a_224_472# 0.008732f
C7206 FILLER_0_16_107/a_36_472# _451_/a_36_151# 0.059367f
C7207 ctln[1] cal_itt\[0\] 0.003349f
C7208 _079_ _001_ 0.082209f
C7209 FILLER_0_12_136/a_572_375# FILLER_0_11_142/a_36_472# 0.001543f
C7210 cal_itt\[3\] FILLER_0_5_198/a_124_375# 0.01268f
C7211 _096_ _136_ 0.022182f
C7212 FILLER_0_4_144/a_484_472# vss 0.033414f
C7213 FILLER_0_18_177/a_124_375# vss 0.00364f
C7214 FILLER_0_18_177/a_572_375# vdd 0.031241f
C7215 _093_ FILLER_0_18_107/a_1020_375# 0.006376f
C7216 _081_ FILLER_0_6_177/a_36_472# 0.00483f
C7217 _418_/a_36_151# vdd 0.155643f
C7218 _411_/a_796_472# net75 0.006358f
C7219 _411_/a_448_472# _000_ 0.073053f
C7220 _074_ _312_/a_234_472# 0.005755f
C7221 _420_/a_36_151# FILLER_0_23_290/a_124_375# 0.026277f
C7222 output12/a_224_472# FILLER_0_1_192/a_124_375# 0.032639f
C7223 net41 _444_/a_1308_423# 0.015841f
C7224 _070_ _385_/a_36_68# 0.049178f
C7225 _014_ FILLER_0_7_233/a_124_375# 0.00143f
C7226 FILLER_0_14_91/a_124_375# vdd -0.010114f
C7227 _413_/a_2248_156# cal_itt\[2\] 0.002527f
C7228 _053_ FILLER_0_6_90/a_36_472# 0.002495f
C7229 net52 FILLER_0_9_72/a_1380_472# 0.003507f
C7230 FILLER_0_20_2/a_572_375# net43 0.051705f
C7231 output48/a_224_472# _079_ 0.003556f
C7232 _138_ vdd 0.090752f
C7233 net47 _039_ 0.042757f
C7234 _106_ FILLER_0_17_218/a_36_472# 0.002777f
C7235 _116_ _061_ 0.04837f
C7236 _149_ _437_/a_36_151# 0.037766f
C7237 trim_mask\[3\] net14 0.142743f
C7238 _095_ _451_/a_448_472# 0.002474f
C7239 net60 _417_/a_36_151# 0.007446f
C7240 _000_ net59 0.004356f
C7241 FILLER_0_15_212/a_1020_375# mask\[1\] 0.017527f
C7242 FILLER_0_19_171/a_1380_472# vss 0.004488f
C7243 _425_/a_796_472# calibrate 0.025807f
C7244 net52 fanout52/a_36_160# 0.036543f
C7245 _253_/a_36_68# net82 0.016638f
C7246 FILLER_0_18_107/a_3172_472# FILLER_0_17_133/a_124_375# 0.001543f
C7247 _000_ net4 0.036895f
C7248 _072_ _311_/a_66_473# 0.031716f
C7249 mask\[5\] _098_ 1.316993f
C7250 FILLER_0_20_169/a_124_375# _098_ 0.019219f
C7251 FILLER_0_18_177/a_1828_472# net21 0.001887f
C7252 _438_/a_2248_156# vdd 0.024595f
C7253 _131_ _040_ 0.211618f
C7254 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_124_375# 0.001597f
C7255 FILLER_0_13_212/a_124_375# net62 0.001597f
C7256 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_572_375# 0.001597f
C7257 _011_ _422_/a_1000_472# 0.005583f
C7258 _308_/a_124_24# net50 0.02221f
C7259 FILLER_0_17_72/a_3260_375# _451_/a_1040_527# 0.001117f
C7260 _431_/a_36_151# net56 0.001371f
C7261 FILLER_0_12_124/a_124_375# _127_ 0.003767f
C7262 FILLER_0_15_282/a_36_472# _006_ 0.003055f
C7263 net15 FILLER_0_15_59/a_484_472# 0.015199f
C7264 _070_ FILLER_0_7_233/a_124_375# 0.004917f
C7265 _072_ _374_/a_244_472# 0.001816f
C7266 net73 FILLER_0_18_107/a_2724_472# 0.02814f
C7267 trim_mask\[4\] _241_/a_224_472# 0.009431f
C7268 net15 _453_/a_448_472# 0.040851f
C7269 output34/a_224_472# _103_ 0.027876f
C7270 FILLER_0_7_72/a_2724_472# trim_mask\[0\] 0.006975f
C7271 _133_ _134_ 0.015205f
C7272 _137_ FILLER_0_19_155/a_572_375# 0.030256f
C7273 fanout53/a_36_160# fanout56/a_36_113# 0.001636f
C7274 net75 FILLER_0_6_231/a_572_375# 0.002577f
C7275 net34 net61 0.037731f
C7276 _432_/a_2665_112# net80 0.041304f
C7277 _242_/a_36_160# _169_ 0.051038f
C7278 _104_ net33 0.037008f
C7279 result[8] FILLER_0_24_274/a_1468_375# 0.00726f
C7280 _092_ mask\[4\] 0.072581f
C7281 FILLER_0_21_125/a_36_472# mask\[7\] 0.00344f
C7282 _178_ net40 0.029542f
C7283 _028_ _164_ 0.019799f
C7284 net50 FILLER_0_6_90/a_572_375# 0.010099f
C7285 result[0] net64 0.09782f
C7286 output8/a_224_472# output11/a_224_472# 0.003437f
C7287 FILLER_0_6_47/a_2364_375# vdd 0.015888f
C7288 FILLER_0_6_47/a_1916_375# vss 0.005279f
C7289 _176_ _315_/a_36_68# 0.003811f
C7290 mask\[5\] net63 0.112147f
C7291 FILLER_0_15_212/a_1020_375# vss 0.035883f
C7292 output47/a_224_472# net40 0.002339f
C7293 FILLER_0_15_212/a_1468_375# vdd 0.010445f
C7294 _449_/a_36_151# FILLER_0_13_72/a_484_472# 0.001723f
C7295 net10 net8 0.003331f
C7296 _402_/a_728_93# vdd 0.050988f
C7297 _322_/a_692_472# net74 0.003192f
C7298 net73 FILLER_0_17_133/a_124_375# 0.022541f
C7299 result[5] fanout78/a_36_113# 0.018989f
C7300 result[5] fanout60/a_36_160# 0.001585f
C7301 output32/a_224_472# net78 0.002901f
C7302 output32/a_224_472# net60 0.191561f
C7303 net31 _094_ 0.203395f
C7304 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_1020_375# 0.026339f
C7305 net23 FILLER_0_16_154/a_484_472# 0.001369f
C7306 net53 _451_/a_3129_107# 0.002806f
C7307 net57 _067_ 0.018966f
C7308 FILLER_0_8_247/a_1020_375# calibrate 0.008393f
C7309 _398_/a_36_113# net3 0.099638f
C7310 net16 FILLER_0_18_53/a_36_472# 0.001532f
C7311 FILLER_0_17_104/a_36_472# net14 0.012286f
C7312 _061_ _117_ 0.046662f
C7313 _419_/a_448_472# net77 0.007659f
C7314 output47/a_224_472# input3/a_36_113# 0.001371f
C7315 _293_/a_36_472# vss 0.014842f
C7316 net52 _443_/a_448_472# 0.050192f
C7317 _057_ _267_/a_1792_472# 0.003005f
C7318 output42/a_224_472# net44 0.079084f
C7319 _384_/a_224_472# vss 0.004801f
C7320 net34 _108_ 0.297364f
C7321 FILLER_0_14_107/a_1020_375# FILLER_0_16_115/a_36_472# 0.001512f
C7322 _077_ FILLER_0_9_72/a_1468_375# 0.008273f
C7323 _023_ mask\[6\] 0.077441f
C7324 _453_/a_1308_423# _042_ 0.001778f
C7325 _453_/a_448_472# net51 0.006397f
C7326 _402_/a_1296_93# cal_count\[1\] 0.004472f
C7327 net73 mask\[9\] 0.383862f
C7328 FILLER_0_18_53/a_572_375# vdd 0.018416f
C7329 cal net18 0.123815f
C7330 _415_/a_36_151# result[1] 0.012965f
C7331 _187_ _181_ 0.001158f
C7332 FILLER_0_16_73/a_484_472# vss 0.007212f
C7333 FILLER_0_16_89/a_124_375# _131_ 0.017319f
C7334 _086_ _375_/a_692_497# 0.002565f
C7335 _433_/a_1308_423# _022_ 0.015376f
C7336 net81 FILLER_0_15_228/a_36_472# 0.003953f
C7337 FILLER_0_4_107/a_124_375# net47 0.004586f
C7338 FILLER_0_1_266/a_36_472# net9 0.041635f
C7339 FILLER_0_3_172/a_1916_375# vdd -0.010166f
C7340 result[0] vss 0.291352f
C7341 _077_ _188_ 0.1656f
C7342 FILLER_0_21_206/a_124_375# net21 0.035287f
C7343 output48/a_224_472# net64 0.002845f
C7344 _422_/a_2665_112# vss 0.006352f
C7345 _065_ net52 0.017184f
C7346 _449_/a_796_472# net72 0.00138f
C7347 _449_/a_36_151# net55 0.003388f
C7348 _033_ vss 0.019158f
C7349 _438_/a_36_151# net14 0.008367f
C7350 FILLER_0_2_111/a_124_375# _157_ 0.028285f
C7351 output14/a_224_472# vdd 0.054725f
C7352 FILLER_0_10_78/a_484_472# _176_ 0.001731f
C7353 _431_/a_36_151# FILLER_0_18_107/a_2276_472# 0.002799f
C7354 _413_/a_448_472# net82 0.004927f
C7355 net55 FILLER_0_17_72/a_1020_375# 0.049648f
C7356 _077_ fanout67/a_36_160# 0.017322f
C7357 _446_/a_1000_472# net66 0.006158f
C7358 _081_ net59 0.185504f
C7359 net73 FILLER_0_19_111/a_36_472# 0.001412f
C7360 FILLER_0_5_72/a_124_375# net49 0.001158f
C7361 _414_/a_2560_156# _074_ 0.001344f
C7362 _005_ _416_/a_36_151# 0.018752f
C7363 fanout50/a_36_160# _164_ 0.08721f
C7364 FILLER_0_3_221/a_932_472# vss 0.002881f
C7365 FILLER_0_3_221/a_1380_472# vdd 0.003819f
C7366 _432_/a_36_151# _141_ 0.008193f
C7367 net4 _081_ 0.02226f
C7368 net54 FILLER_0_18_139/a_1020_375# 0.003589f
C7369 _056_ _310_/a_49_472# 0.003286f
C7370 FILLER_0_16_73/a_484_472# cal_count\[1\] 0.001135f
C7371 FILLER_0_19_47/a_124_375# _052_ 0.019401f
C7372 FILLER_0_16_73/a_572_375# net15 0.002076f
C7373 FILLER_0_20_193/a_36_472# _098_ 0.006652f
C7374 _451_/a_1353_112# vdd 0.009693f
C7375 ctln[1] _411_/a_1308_423# 0.037098f
C7376 FILLER_0_5_72/a_484_472# _029_ 0.004625f
C7377 FILLER_0_5_72/a_1020_375# trim_mask\[1\] 0.010728f
C7378 FILLER_0_3_172/a_3172_472# net21 0.037958f
C7379 _086_ _267_/a_1120_472# 0.004245f
C7380 mask\[9\] FILLER_0_19_111/a_484_472# 0.041744f
C7381 _001_ vss 0.004381f
C7382 _065_ net41 0.001765f
C7383 net19 _009_ 0.055383f
C7384 net26 _423_/a_796_472# 0.001077f
C7385 _413_/a_2248_156# net59 0.05485f
C7386 FILLER_0_4_123/a_36_472# net69 0.001015f
C7387 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1380_472# 0.013276f
C7388 FILLER_0_9_270/a_484_472# FILLER_0_9_282/a_36_472# 0.002296f
C7389 _431_/a_1000_472# _136_ 0.024253f
C7390 net22 _435_/a_36_151# 0.001559f
C7391 net57 _121_ 0.004182f
C7392 FILLER_0_21_133/a_36_472# _433_/a_36_151# 0.001723f
C7393 _059_ net37 0.011845f
C7394 output37/a_224_472# net37 0.011407f
C7395 _350_/a_49_472# vdd 0.026837f
C7396 FILLER_0_17_218/a_124_375# _069_ 0.003162f
C7397 net51 _450_/a_3129_107# 0.030082f
C7398 _004_ net64 0.001495f
C7399 FILLER_0_2_111/a_484_472# vdd 0.005951f
C7400 _142_ FILLER_0_17_133/a_36_472# 0.069383f
C7401 _077_ _256_/a_36_68# 0.027906f
C7402 _188_ _453_/a_36_151# 0.03354f
C7403 FILLER_0_21_286/a_124_375# net18 0.015582f
C7404 _062_ vss 0.58133f
C7405 _431_/a_448_472# fanout70/a_36_113# 0.001157f
C7406 output48/a_224_472# vss 0.006655f
C7407 _396_/a_224_472# net36 0.00114f
C7408 _098_ FILLER_0_16_154/a_1020_375# 0.003386f
C7409 _004_ mask\[1\] 0.052788f
C7410 _414_/a_2665_112# net59 0.010265f
C7411 _449_/a_448_472# FILLER_0_11_64/a_36_472# 0.001462f
C7412 _036_ _167_ 0.003223f
C7413 net78 _418_/a_36_151# 0.003648f
C7414 net60 _418_/a_36_151# 0.016348f
C7415 net28 _195_/a_67_603# 0.012984f
C7416 ctln[6] _442_/a_448_472# 0.003039f
C7417 net20 _419_/a_1308_423# 0.022245f
C7418 net60 _419_/a_1204_472# 0.023544f
C7419 net61 _419_/a_2665_112# 0.022394f
C7420 _136_ FILLER_0_15_180/a_124_375# 0.002442f
C7421 _053_ _251_/a_906_472# 0.001696f
C7422 net3 cal_count\[2\] 0.119728f
C7423 net63 FILLER_0_20_193/a_36_472# 0.048818f
C7424 FILLER_0_7_162/a_36_472# _081_ 0.002493f
C7425 mask\[3\] _137_ 0.231419f
C7426 net76 net22 0.118787f
C7427 net17 vdd 2.139315f
C7428 net74 _062_ 0.062376f
C7429 FILLER_0_17_200/a_124_375# net63 0.008905f
C7430 _142_ net73 0.090025f
C7431 FILLER_0_21_28/a_2276_472# _012_ 0.023696f
C7432 FILLER_0_21_150/a_124_375# vdd 0.020581f
C7433 _031_ _154_ 0.037238f
C7434 net69 _153_ 0.003678f
C7435 net81 net76 0.236554f
C7436 FILLER_0_12_136/a_484_472# net23 0.002172f
C7437 net47 clkc 0.002956f
C7438 _150_ net36 0.108945f
C7439 FILLER_0_4_49/a_124_375# _232_/a_67_603# 0.002082f
C7440 _308_/a_1152_472# trim_mask\[0\] 0.004076f
C7441 FILLER_0_9_28/a_2364_375# trim_val\[0\] 0.006639f
C7442 FILLER_0_15_142/a_572_375# net36 0.006382f
C7443 _104_ _046_ 0.035267f
C7444 FILLER_0_17_200/a_484_472# net22 0.020589f
C7445 _176_ FILLER_0_15_72/a_572_375# 0.005529f
C7446 net38 FILLER_0_20_2/a_484_472# 0.006727f
C7447 net75 _015_ 0.025217f
C7448 net52 _176_ 0.004215f
C7449 net72 FILLER_0_12_50/a_36_472# 0.002007f
C7450 mask\[2\] net23 0.431197f
C7451 _004_ vss 0.115789f
C7452 _052_ net15 0.001074f
C7453 net4 FILLER_0_12_220/a_932_472# 0.050731f
C7454 _086_ _074_ 0.186795f
C7455 _100_ _094_ 0.031066f
C7456 _423_/a_36_151# FILLER_0_23_44/a_1468_375# 0.059049f
C7457 FILLER_0_7_104/a_484_472# _058_ 0.006506f
C7458 _064_ net47 0.110169f
C7459 _099_ net30 0.05959f
C7460 FILLER_0_15_116/a_124_375# net36 0.003055f
C7461 net31 output34/a_224_472# 0.165772f
C7462 _427_/a_448_472# _095_ 0.063616f
C7463 net75 FILLER_0_0_232/a_36_472# 0.001514f
C7464 net68 FILLER_0_5_54/a_572_375# 0.040374f
C7465 FILLER_0_17_200/a_36_472# FILLER_0_18_177/a_2724_472# 0.026657f
C7466 net19 cal_itt\[0\] 0.111163f
C7467 mask\[0\] cal_count\[3\] 0.002612f
C7468 FILLER_0_5_54/a_1468_375# trim_mask\[1\] 0.010901f
C7469 FILLER_0_5_54/a_932_472# _029_ 0.014976f
C7470 FILLER_0_5_212/a_36_472# net37 0.007858f
C7471 _304_/a_224_472# _013_ 0.002769f
C7472 net50 net49 0.238748f
C7473 FILLER_0_21_142/a_124_375# vss 0.009345f
C7474 FILLER_0_21_142/a_572_375# vdd 0.002442f
C7475 _441_/a_36_151# _440_/a_448_472# 0.002538f
C7476 net52 _442_/a_2560_156# 0.008682f
C7477 _058_ FILLER_0_10_94/a_124_375# 0.001597f
C7478 result[7] FILLER_0_23_290/a_124_375# 0.018455f
C7479 FILLER_0_9_28/a_1380_472# _054_ 0.004017f
C7480 _019_ net21 0.065941f
C7481 net17 _452_/a_1040_527# 0.034254f
C7482 fanout50/a_36_160# trim_val\[3\] 0.017252f
C7483 net52 _036_ 0.013473f
C7484 net50 net68 0.224698f
C7485 net35 _023_ 0.008361f
C7486 FILLER_0_17_72/a_1828_472# vss 0.001443f
C7487 FILLER_0_17_72/a_2276_472# vdd 0.001409f
C7488 fanout79/a_36_160# _060_ 0.005814f
C7489 net7 _065_ 0.0295f
C7490 FILLER_0_7_195/a_36_472# vss 0.002568f
C7491 _091_ net4 0.125608f
C7492 FILLER_0_21_206/a_36_472# _204_/a_67_603# 0.003123f
C7493 _068_ FILLER_0_5_148/a_484_472# 0.016952f
C7494 FILLER_0_16_37/a_124_375# vss 0.021237f
C7495 FILLER_0_16_37/a_36_472# vdd 0.142203f
C7496 _429_/a_2248_156# _043_ 0.001001f
C7497 FILLER_0_3_142/a_36_472# _081_ 0.001386f
C7498 FILLER_0_8_127/a_124_375# _133_ 0.001928f
C7499 FILLER_0_8_127/a_36_472# _070_ 0.005078f
C7500 ctlp[4] mask\[5\] 0.001643f
C7501 FILLER_0_19_195/a_124_375# net21 0.039225f
C7502 net33 _434_/a_2665_112# 0.001043f
C7503 mask\[2\] FILLER_0_15_180/a_484_472# 0.00848f
C7504 _440_/a_2665_112# FILLER_0_4_91/a_124_375# 0.006271f
C7505 net76 _076_ 0.003124f
C7506 _144_ net23 0.091811f
C7507 _013_ FILLER_0_18_53/a_484_472# 0.012916f
C7508 FILLER_0_19_187/a_484_472# vss 0.004504f
C7509 _011_ vss 0.003987f
C7510 _136_ _337_/a_49_472# 0.058704f
C7511 mask\[3\] net56 0.002632f
C7512 FILLER_0_1_192/a_124_375# vss 0.049811f
C7513 FILLER_0_1_192/a_36_472# vdd 0.011806f
C7514 _140_ FILLER_0_21_150/a_36_472# 0.015502f
C7515 FILLER_0_4_213/a_36_472# net59 0.044235f
C7516 FILLER_0_13_212/a_572_375# _070_ 0.003986f
C7517 net15 mask\[9\] 0.128816f
C7518 FILLER_0_18_171/a_124_375# mask\[4\] 0.008445f
C7519 FILLER_0_3_2/a_124_375# net66 0.027628f
C7520 FILLER_0_11_124/a_124_375# _135_ 0.004831f
C7521 net25 _012_ 0.001747f
C7522 _171_ _172_ 0.104216f
C7523 _255_/a_224_552# FILLER_0_6_177/a_572_375# 0.001776f
C7524 FILLER_0_4_107/a_484_472# _031_ 0.002521f
C7525 net20 FILLER_0_6_239/a_124_375# 0.004897f
C7526 _131_ FILLER_0_9_105/a_484_472# 0.004364f
C7527 _115_ _135_ 0.004345f
C7528 FILLER_0_17_72/a_932_472# net15 0.001122f
C7529 en fanout59/a_36_160# 0.242369f
C7530 net18 output30/a_224_472# 0.08667f
C7531 net41 _445_/a_2665_112# 0.056125f
C7532 _012_ net36 0.053654f
C7533 _205_/a_36_160# _047_ 0.013528f
C7534 FILLER_0_19_125/a_124_375# _334_/a_36_160# 0.001633f
C7535 _093_ _438_/a_2248_156# 0.004221f
C7536 _083_ FILLER_0_3_221/a_572_375# 0.001072f
C7537 _441_/a_448_472# vdd 0.007984f
C7538 _441_/a_36_151# vss 0.015116f
C7539 _098_ _434_/a_1000_472# 0.00725f
C7540 _340_/a_36_160# _098_ 0.019601f
C7541 _235_/a_67_603# vdd 0.026582f
C7542 net53 _427_/a_2248_156# 0.038716f
C7543 net49 trim_mask\[3\] 0.03723f
C7544 _444_/a_2665_112# net67 0.03521f
C7545 net72 _452_/a_36_151# 0.040035f
C7546 _442_/a_2248_156# trim_mask\[3\] 0.003039f
C7547 _015_ _426_/a_36_151# 0.01243f
C7548 output17/a_224_472# net17 0.09023f
C7549 FILLER_0_15_228/a_124_375# vdd 0.013701f
C7550 _431_/a_36_151# vss 0.00849f
C7551 _431_/a_448_472# vdd 0.001932f
C7552 _104_ net18 0.039321f
C7553 _440_/a_1000_472# vss 0.031704f
C7554 net34 _049_ 0.048403f
C7555 FILLER_0_19_142/a_124_375# vdd 0.022448f
C7556 _430_/a_36_151# _069_ 0.026308f
C7557 _439_/a_36_151# vdd 0.095368f
C7558 _254_/a_244_472# _072_ 0.001552f
C7559 net80 _434_/a_1308_423# 0.006837f
C7560 _044_ vss 0.038421f
C7561 _157_ vdd 0.419501f
C7562 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_36_472# 0.086743f
C7563 _091_ FILLER_0_13_212/a_1020_375# 0.00799f
C7564 net34 _435_/a_2665_112# 0.009214f
C7565 _119_ _062_ 0.080398f
C7566 _432_/a_2248_156# net21 0.002329f
C7567 trim_mask\[2\] FILLER_0_2_93/a_572_375# 0.002818f
C7568 _420_/a_36_151# net18 0.001426f
C7569 _176_ _172_ 0.043154f
C7570 _098_ _437_/a_36_151# 0.092841f
C7571 _086_ _124_ 0.063099f
C7572 FILLER_0_21_142/a_36_472# _140_ 0.009261f
C7573 net36 FILLER_0_15_235/a_484_472# 0.019725f
C7574 _277_/a_36_160# vss 0.030147f
C7575 _250_/a_36_68# _427_/a_2665_112# 0.002152f
C7576 FILLER_0_7_104/a_572_375# _131_ 0.003031f
C7577 FILLER_0_19_47/a_572_375# vss 0.055293f
C7578 FILLER_0_19_47/a_36_472# vdd 0.072773f
C7579 comp _043_ 0.003867f
C7580 net36 _438_/a_448_472# 0.034338f
C7581 _015_ FILLER_0_8_239/a_124_375# 0.007342f
C7582 FILLER_0_14_91/a_36_472# en_co_clk 0.007733f
C7583 net63 _434_/a_1000_472# 0.002404f
C7584 _132_ FILLER_0_18_107/a_2364_375# 0.006403f
C7585 _316_/a_124_24# vss 0.00516f
C7586 _316_/a_848_380# vdd 0.048727f
C7587 net39 vdd 0.2282f
C7588 _053_ FILLER_0_7_104/a_36_472# 0.01752f
C7589 _089_ FILLER_0_5_198/a_36_472# 0.001314f
C7590 _444_/a_2560_156# _054_ 0.003269f
C7591 mask\[5\] FILLER_0_20_177/a_1020_375# 0.013294f
C7592 FILLER_0_16_57/a_124_375# net72 0.052543f
C7593 _385_/a_244_472# net37 0.001593f
C7594 _144_ net33 0.042826f
C7595 FILLER_0_24_96/a_36_472# net25 0.040228f
C7596 input4/a_36_68# vss 0.058179f
C7597 FILLER_0_17_72/a_3260_375# net14 0.040606f
C7598 _423_/a_2560_156# _012_ 0.004165f
C7599 net15 _440_/a_1308_423# 0.015192f
C7600 _430_/a_2665_112# net36 0.003477f
C7601 _412_/a_2248_156# net1 0.044934f
C7602 FILLER_0_9_28/a_1468_375# net16 0.005202f
C7603 net79 _005_ 1.006306f
C7604 net75 fanout75/a_36_113# 0.035159f
C7605 FILLER_0_22_86/a_36_472# net14 0.003007f
C7606 _308_/a_848_380# FILLER_0_10_94/a_484_472# 0.019491f
C7607 net79 FILLER_0_12_220/a_932_472# 0.005532f
C7608 FILLER_0_18_2/a_2812_375# _452_/a_36_151# 0.001597f
C7609 _448_/a_1000_472# net59 0.007647f
C7610 _053_ _414_/a_1204_472# 0.003935f
C7611 _395_/a_36_488# state\[1\] 0.002702f
C7612 _116_ _267_/a_36_472# 0.029316f
C7613 _122_ _059_ 0.190023f
C7614 mask\[5\] _137_ 0.002972f
C7615 _427_/a_448_472# vss 0.040679f
C7616 _427_/a_1308_423# vdd 0.002814f
C7617 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_36_472# 0.086742f
C7618 FILLER_0_16_241/a_124_375# mask\[2\] 0.027201f
C7619 FILLER_0_7_72/a_484_472# vss 0.003793f
C7620 net20 _088_ 0.001704f
C7621 ctln[3] net75 0.066513f
C7622 vss FILLER_0_5_148/a_36_472# 0.029152f
C7623 net35 net15 0.01797f
C7624 _412_/a_448_472# _082_ 0.022743f
C7625 FILLER_0_9_28/a_1020_375# vdd 0.033815f
C7626 _430_/a_36_151# FILLER_0_18_209/a_484_472# 0.001043f
C7627 _405_/a_67_603# cal_count\[2\] 0.021962f
C7628 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1380_472# 0.013277f
C7629 FILLER_0_20_169/a_124_375# FILLER_0_19_171/a_36_472# 0.001543f
C7630 mask\[5\] FILLER_0_19_171/a_36_472# 0.002923f
C7631 ctln[1] FILLER_0_0_232/a_124_375# 0.012033f
C7632 _028_ _133_ 0.007084f
C7633 _002_ FILLER_0_3_172/a_2276_472# 0.030358f
C7634 net48 net37 0.081653f
C7635 ctlp[1] net79 0.002676f
C7636 _131_ cal_count\[2\] 0.044147f
C7637 FILLER_0_24_130/a_124_375# _050_ 0.007643f
C7638 FILLER_0_21_28/a_36_472# net17 0.00347f
C7639 _427_/a_448_472# net74 0.051943f
C7640 _437_/a_2560_156# net14 0.00349f
C7641 output27/a_224_472# FILLER_0_8_263/a_124_375# 0.011584f
C7642 net44 _450_/a_448_472# 0.050752f
C7643 state\[1\] _228_/a_36_68# 0.024977f
C7644 _091_ net79 0.052824f
C7645 net62 output30/a_224_472# 0.074425f
C7646 _076_ _083_ 0.006023f
C7647 _359_/a_1492_488# _133_ 0.003815f
C7648 _068_ _078_ 0.002973f
C7649 net16 _173_ 0.029412f
C7650 _072_ _085_ 0.408915f
C7651 FILLER_0_22_177/a_1020_375# net33 0.013731f
C7652 _028_ _376_/a_36_160# 0.026437f
C7653 FILLER_0_22_177/a_1380_472# _435_/a_36_151# 0.001723f
C7654 output15/a_224_472# net52 0.007862f
C7655 _163_ FILLER_0_6_79/a_36_472# 0.001789f
C7656 FILLER_0_16_73/a_36_472# _394_/a_1336_472# 0.00108f
C7657 FILLER_0_19_155/a_572_375# vss 0.004538f
C7658 _442_/a_1308_423# _031_ 0.003679f
C7659 _131_ FILLER_0_11_124/a_36_472# 0.015445f
C7660 result[0] FILLER_0_9_290/a_36_472# 0.020103f
C7661 FILLER_0_5_72/a_124_375# net47 0.006974f
C7662 _115_ _129_ 0.021405f
C7663 net14 FILLER_0_4_91/a_572_375# 0.047331f
C7664 _053_ FILLER_0_8_37/a_484_472# 0.002095f
C7665 _350_/a_49_472# _147_ 0.016114f
C7666 net34 FILLER_0_22_128/a_2724_472# 0.004465f
C7667 mask\[0\] _429_/a_2665_112# 0.016053f
C7668 cal_itt\[3\] _081_ 0.03503f
C7669 FILLER_0_16_107/a_572_375# _040_ 0.001244f
C7670 net24 FILLER_0_22_86/a_1020_375# 0.022658f
C7671 _140_ _207_/a_67_603# 0.014923f
C7672 FILLER_0_18_177/a_3172_472# vss 0.002639f
C7673 net80 net21 0.016911f
C7674 FILLER_0_7_59/a_124_375# vdd -0.006113f
C7675 _132_ net70 0.534228f
C7676 trimb[4] FILLER_0_15_2/a_36_472# 0.006046f
C7677 net16 _444_/a_36_151# 0.010514f
C7678 FILLER_0_20_177/a_1380_472# _098_ 0.00679f
C7679 net81 FILLER_0_8_263/a_124_375# 0.026195f
C7680 net35 FILLER_0_22_128/a_1916_375# 0.014552f
C7681 net77 vss 0.327705f
C7682 FILLER_0_5_212/a_36_472# _122_ 0.002272f
C7683 FILLER_0_3_204/a_124_375# FILLER_0_3_172/a_3260_375# 0.012001f
C7684 _114_ FILLER_0_12_136/a_1020_375# 0.006974f
C7685 _077_ FILLER_0_9_105/a_484_472# 0.002951f
C7686 net31 _293_/a_36_472# 0.005692f
C7687 _046_ mask\[2\] 0.003147f
C7688 _256_/a_2552_68# _076_ 0.00144f
C7689 FILLER_0_16_241/a_36_472# _282_/a_36_160# 0.006647f
C7690 _376_/a_36_160# FILLER_0_6_90/a_36_472# 0.195478f
C7691 _085_ FILLER_0_13_142/a_1468_375# 0.001153f
C7692 FILLER_0_9_105/a_484_472# FILLER_0_10_107/a_124_375# 0.001543f
C7693 _255_/a_224_552# _374_/a_36_68# 0.00191f
C7694 FILLER_0_16_57/a_1380_472# vss 0.011192f
C7695 trim_mask\[1\] FILLER_0_6_47/a_572_375# 0.007164f
C7696 _303_/a_36_472# vss 0.011549f
C7697 result[6] _419_/a_36_151# 0.001968f
C7698 _102_ vss 0.068703f
C7699 net52 _449_/a_448_472# 0.001042f
C7700 FILLER_0_22_128/a_2812_375# vdd 0.003766f
C7701 FILLER_0_22_128/a_2364_375# vss 0.017496f
C7702 _162_ _058_ 0.015239f
C7703 _415_/a_2248_156# net18 0.057604f
C7704 result[7] _046_ 0.003397f
C7705 FILLER_0_17_72/a_572_375# FILLER_0_15_72/a_484_472# 0.001512f
C7706 _414_/a_2665_112# cal_itt\[3\] 0.02392f
C7707 _126_ _390_/a_36_68# 0.044675f
C7708 net50 FILLER_0_8_37/a_36_472# 0.059367f
C7709 _421_/a_36_151# _419_/a_36_151# 0.561555f
C7710 ctlp[0] vdd 0.08832f
C7711 net55 _451_/a_3129_107# 0.098091f
C7712 _177_ _131_ 0.058938f
C7713 FILLER_0_21_142/a_124_375# _433_/a_448_472# 0.006782f
C7714 fanout79/a_36_160# vss 0.002268f
C7715 net63 FILLER_0_20_177/a_1380_472# 0.011079f
C7716 net82 _159_ 0.001393f
C7717 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3260_375# 0.001597f
C7718 _140_ FILLER_0_19_155/a_484_472# 0.004155f
C7719 _217_/a_36_160# FILLER_0_19_28/a_484_472# 0.006053f
C7720 net65 _413_/a_448_472# 0.044062f
C7721 net38 net40 1.103743f
C7722 vss output41/a_224_472# -0.007739f
C7723 net27 FILLER_0_9_270/a_124_375# 0.079454f
C7724 mask\[3\] net64 0.002654f
C7725 net23 _386_/a_124_24# 0.010805f
C7726 FILLER_0_10_78/a_124_375# vdd -0.011193f
C7727 _408_/a_728_93# _043_ 0.029183f
C7728 output38/a_224_472# _064_ 0.017666f
C7729 _176_ FILLER_0_11_101/a_572_375# 0.00389f
C7730 _428_/a_796_472# _017_ 0.025239f
C7731 _116_ _113_ 0.179616f
C7732 FILLER_0_21_28/a_2364_375# _424_/a_36_151# 0.059049f
C7733 FILLER_0_4_123/a_36_472# vss 0.004542f
C7734 FILLER_0_16_107/a_124_375# net36 0.001706f
C7735 FILLER_0_16_57/a_1380_472# cal_count\[1\] 0.001568f
C7736 FILLER_0_16_57/a_484_472# net15 0.008573f
C7737 _098_ _438_/a_2665_112# 0.004321f
C7738 _104_ _109_ 0.029532f
C7739 net63 FILLER_0_18_177/a_1020_375# 0.007516f
C7740 FILLER_0_5_54/a_572_375# net47 0.009717f
C7741 net42 vdd 0.178782f
C7742 FILLER_0_2_111/a_932_472# _158_ 0.00264f
C7743 _277_/a_36_160# _103_ 0.032112f
C7744 FILLER_0_9_72/a_36_472# vdd 0.109576f
C7745 FILLER_0_9_72/a_1468_375# vss 0.013085f
C7746 output29/a_224_472# _005_ 0.021351f
C7747 net29 _101_ 0.007132f
C7748 net82 FILLER_0_3_172/a_2364_375# 0.010439f
C7749 output14/a_224_472# _442_/a_36_151# 0.172111f
C7750 net58 _082_ 0.004276f
C7751 _171_ FILLER_0_10_94/a_36_472# 0.001514f
C7752 _172_ FILLER_0_10_94/a_124_375# 0.003341f
C7753 FILLER_0_4_123/a_36_472# net74 0.001578f
C7754 FILLER_0_4_144/a_36_472# _370_/a_848_380# 0.15783f
C7755 net75 FILLER_0_8_247/a_1380_472# 0.020589f
C7756 net55 FILLER_0_13_72/a_572_375# 0.005919f
C7757 _093_ FILLER_0_17_72/a_2276_472# 0.017114f
C7758 _165_ trim_mask\[1\] 0.002231f
C7759 _182_ vss 0.068928f
C7760 _359_/a_36_488# vdd 0.083138f
C7761 _078_ vdd 0.181583f
C7762 _130_ FILLER_0_11_124/a_36_472# 0.003572f
C7763 _198_/a_67_603# vss 0.003647f
C7764 net50 net47 0.040157f
C7765 _028_ FILLER_0_7_72/a_1468_375# 0.003785f
C7766 _115_ _219_/a_36_160# 0.001218f
C7767 _394_/a_56_524# _095_ 0.10007f
C7768 _137_ FILLER_0_16_154/a_1020_375# 0.010692f
C7769 _081_ FILLER_0_5_164/a_36_472# 0.001603f
C7770 _188_ vss 0.032923f
C7771 net43 FILLER_0_20_15/a_124_375# 0.005925f
C7772 FILLER_0_6_90/a_36_472# FILLER_0_4_91/a_124_375# 0.001188f
C7773 net76 FILLER_0_5_172/a_124_375# 0.001526f
C7774 net18 _417_/a_1000_472# 0.056791f
C7775 fanout70/a_36_113# net36 0.007807f
C7776 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_124_375# 0.012267f
C7777 _127_ _332_/a_36_472# 0.00288f
C7778 trim[0] trim[1] 0.001567f
C7779 net75 _426_/a_1000_472# 0.002727f
C7780 _273_/a_36_68# net4 0.06843f
C7781 FILLER_0_16_89/a_36_472# _136_ 0.00722f
C7782 result[6] _420_/a_2248_156# 0.003418f
C7783 net26 FILLER_0_18_37/a_932_472# 0.002613f
C7784 FILLER_0_17_200/a_572_375# vdd 0.006861f
C7785 FILLER_0_15_282/a_572_375# output30/a_224_472# 0.029138f
C7786 FILLER_0_2_171/a_36_472# FILLER_0_2_165/a_36_472# 0.003468f
C7787 FILLER_0_9_223/a_124_375# _246_/a_36_68# 0.005308f
C7788 FILLER_0_18_107/a_1020_375# FILLER_0_17_104/a_1380_472# 0.001597f
C7789 fanout67/a_36_160# vss 0.005344f
C7790 FILLER_0_12_136/a_1020_375# _126_ 0.012732f
C7791 _098_ FILLER_0_15_212/a_36_472# 0.011079f
C7792 _176_ _318_/a_224_472# 0.003019f
C7793 _116_ _118_ 0.054068f
C7794 _136_ _171_ 0.008792f
C7795 net52 _032_ 0.009879f
C7796 _153_ vss 0.256017f
C7797 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_36_472# 0.001963f
C7798 _088_ _073_ 0.001254f
C7799 FILLER_0_14_50/a_36_472# _180_ 0.153222f
C7800 _104_ _422_/a_448_472# 0.001955f
C7801 _153_ _365_/a_692_472# 0.002377f
C7802 mask\[8\] _050_ 0.001479f
C7803 mask\[3\] vss 0.664467f
C7804 net10 vdd 0.227004f
C7805 _443_/a_36_151# trim_mask\[4\] 0.002625f
C7806 calibrate _385_/a_36_68# 0.001996f
C7807 _176_ FILLER_0_10_94/a_36_472# 0.009089f
C7808 _140_ FILLER_0_22_128/a_3260_375# 0.003524f
C7809 trimb[3] FILLER_0_20_2/a_484_472# 0.001829f
C7810 _427_/a_2248_156# _071_ 0.001131f
C7811 fanout49/a_36_160# _160_ 0.009662f
C7812 _275_/a_224_472# _092_ 0.002138f
C7813 FILLER_0_17_72/a_36_472# net36 0.001121f
C7814 _132_ FILLER_0_14_107/a_572_375# 0.007439f
C7815 FILLER_0_10_214/a_124_375# _055_ 0.001419f
C7816 _042_ net51 0.026776f
C7817 _441_/a_36_151# FILLER_0_3_78/a_36_472# 0.001723f
C7818 ctlp[1] FILLER_0_21_286/a_36_472# 0.014043f
C7819 _423_/a_36_151# FILLER_0_23_60/a_36_472# 0.001723f
C7820 _182_ cal_count\[1\] 0.166348f
C7821 _442_/a_1308_423# FILLER_0_2_111/a_1468_375# 0.001048f
C7822 FILLER_0_8_138/a_36_472# _059_ 0.02252f
C7823 _257_/a_36_472# _070_ 0.002295f
C7824 trim_val\[0\] _220_/a_67_603# 0.005346f
C7825 _060_ _223_/a_36_160# 0.002922f
C7826 net73 FILLER_0_17_142/a_36_472# 0.002925f
C7827 net15 cal_count\[3\] 0.045013f
C7828 _070_ _171_ 0.084342f
C7829 FILLER_0_21_28/a_2276_472# vdd 0.002733f
C7830 FILLER_0_21_28/a_1828_472# vss -0.001894f
C7831 FILLER_0_6_90/a_124_375# vdd 0.020992f
C7832 fanout51/a_36_113# cal_count\[3\] 0.054567f
C7833 _050_ vss 0.26237f
C7834 result[7] net18 0.098317f
C7835 _163_ _365_/a_36_68# 0.004035f
C7836 _061_ _247_/a_36_160# 0.009993f
C7837 _431_/a_448_472# _093_ 0.002095f
C7838 output9/a_224_472# FILLER_0_1_266/a_36_472# 0.001007f
C7839 _117_ _113_ 0.09166f
C7840 result[6] _421_/a_2560_156# 0.006943f
C7841 _430_/a_36_151# net22 0.005321f
C7842 _004_ _416_/a_2665_112# 0.002631f
C7843 net63 FILLER_0_15_212/a_36_472# 0.059367f
C7844 FILLER_0_11_282/a_124_375# vdd 0.026044f
C7845 _320_/a_36_472# _090_ 0.001941f
C7846 _176_ _136_ 0.114837f
C7847 _093_ FILLER_0_19_142/a_124_375# 0.00346f
C7848 _002_ net82 0.034599f
C7849 _256_/a_36_68# vss 0.055568f
C7850 net58 fanout64/a_36_160# 0.002438f
C7851 net50 FILLER_0_9_60/a_124_375# 0.001715f
C7852 FILLER_0_18_2/a_2276_472# net17 0.037088f
C7853 _233_/a_36_160# net40 0.001875f
C7854 _004_ FILLER_0_10_247/a_36_472# 0.001551f
C7855 _035_ net49 0.018245f
C7856 _115_ FILLER_0_10_107/a_572_375# 0.040198f
C7857 _163_ FILLER_0_5_148/a_124_375# 0.001706f
C7858 FILLER_0_19_55/a_124_375# _052_ 0.053626f
C7859 _136_ _335_/a_49_472# 0.039074f
C7860 _253_/a_36_68# FILLER_0_3_221/a_1468_375# 0.014131f
C7861 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_124_375# 0.012222f
C7862 _430_/a_36_151# net81 0.017255f
C7863 FILLER_0_5_117/a_36_472# vss 0.001215f
C7864 fanout49/a_36_160# _030_ 0.017759f
C7865 trim_mask\[0\] FILLER_0_10_94/a_572_375# 0.003359f
C7866 _068_ _160_ 0.003424f
C7867 fanout64/a_36_160# _425_/a_2665_112# 0.005704f
C7868 calibrate FILLER_0_7_233/a_124_375# 0.011958f
C7869 output17/a_224_472# ctlp[0] 0.018696f
C7870 FILLER_0_19_142/a_124_375# FILLER_0_19_134/a_124_375# 0.003732f
C7871 mask\[9\] FILLER_0_18_76/a_36_472# 0.002584f
C7872 net48 _122_ 0.110769f
C7873 trim_val\[4\] FILLER_0_3_172/a_36_472# 0.006208f
C7874 net76 FILLER_0_3_172/a_2276_472# 0.002531f
C7875 trim_val\[4\] _386_/a_124_24# 0.001172f
C7876 _426_/a_36_151# FILLER_0_8_247/a_1380_472# 0.001723f
C7877 net72 _423_/a_36_151# 0.024965f
C7878 trim_mask\[1\] FILLER_0_6_79/a_124_375# 0.0042f
C7879 FILLER_0_7_72/a_124_375# net52 0.029774f
C7880 FILLER_0_7_162/a_36_472# FILLER_0_8_156/a_572_375# 0.001543f
C7881 _040_ vss 0.216709f
C7882 ctln[1] net58 0.014147f
C7883 vss _433_/a_1000_472# 0.002059f
C7884 _320_/a_36_472# net22 0.005964f
C7885 _116_ _068_ 0.011673f
C7886 _176_ _070_ 0.467961f
C7887 net56 FILLER_0_18_139/a_932_472# 0.011079f
C7888 _070_ FILLER_0_5_164/a_572_375# 0.001083f
C7889 _334_/a_36_160# vdd 0.041716f
C7890 FILLER_0_20_177/a_932_472# _434_/a_36_151# 0.001723f
C7891 FILLER_0_15_290/a_36_472# net18 0.002452f
C7892 net56 FILLER_0_16_154/a_1020_375# 0.002321f
C7893 fanout53/a_36_160# FILLER_0_16_154/a_484_472# 0.014774f
C7894 net52 FILLER_0_2_93/a_124_375# 0.007787f
C7895 ctlp[1] ctlp[2] 0.002331f
C7896 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1468_375# 0.001597f
C7897 _149_ net14 0.102004f
C7898 _118_ _117_ 0.032074f
C7899 _432_/a_36_151# mask\[2\] 0.031341f
C7900 cal_count\[3\] net51 0.042416f
C7901 net67 FILLER_0_6_47/a_124_375# 0.005516f
C7902 output24/a_224_472# net24 0.005559f
C7903 net55 net40 0.043962f
C7904 net55 _424_/a_448_472# 0.005273f
C7905 _020_ fanout70/a_36_113# 0.001266f
C7906 _239_/a_36_160# vdd 0.042369f
C7907 mask\[3\] FILLER_0_18_177/a_1828_472# 0.004274f
C7908 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_484_472# 0.026657f
C7909 output36/a_224_472# net29 0.077505f
C7910 FILLER_0_4_107/a_1380_472# vss 0.004455f
C7911 _103_ net77 0.004691f
C7912 _417_/a_1000_472# net62 0.005762f
C7913 net67 _450_/a_836_156# 0.008805f
C7914 _415_/a_2665_112# net58 0.005219f
C7915 FILLER_0_12_20/a_484_472# vdd 0.003108f
C7916 _058_ FILLER_0_8_156/a_124_375# 0.006325f
C7917 FILLER_0_18_2/a_3260_375# net55 0.004262f
C7918 vss FILLER_0_12_196/a_36_472# 0.003551f
C7919 ctln[6] _031_ 0.004486f
C7920 _413_/a_448_472# output12/a_224_472# 0.001495f
C7921 _232_/a_67_603# FILLER_0_5_54/a_36_472# 0.025312f
C7922 FILLER_0_24_130/a_36_472# net54 0.06125f
C7923 _049_ _146_ 0.042698f
C7924 cal_count\[1\] _040_ 0.019478f
C7925 _079_ _253_/a_36_68# 0.002433f
C7926 _112_ FILLER_0_8_247/a_932_472# 0.001185f
C7927 net4 _246_/a_36_68# 0.003771f
C7928 net18 FILLER_0_17_282/a_36_472# 0.036965f
C7929 mask\[5\] FILLER_0_19_187/a_124_375# 0.007169f
C7930 _321_/a_3662_472# net74 0.00253f
C7931 _072_ FILLER_0_12_220/a_36_472# 0.01861f
C7932 _431_/a_448_472# FILLER_0_17_142/a_124_375# 0.006782f
C7933 _103_ _102_ 0.392644f
C7934 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_124_375# 0.012001f
C7935 _414_/a_36_151# _074_ 0.070632f
C7936 net20 _260_/a_36_68# 0.033776f
C7937 _424_/a_36_151# _423_/a_36_151# 0.006746f
C7938 FILLER_0_20_87/a_124_375# vdd 0.008846f
C7939 FILLER_0_14_81/a_36_472# _394_/a_728_93# 0.005826f
C7940 FILLER_0_11_78/a_572_375# _171_ 0.001028f
C7941 _287_/a_36_472# _099_ 0.030964f
C7942 _363_/a_692_472# _028_ 0.001416f
C7943 net25 vdd 0.195306f
C7944 _322_/a_1152_472# _129_ 0.002978f
C7945 FILLER_0_9_223/a_572_375# _055_ 0.022619f
C7946 _440_/a_36_151# _160_ 0.002966f
C7947 _028_ FILLER_0_6_47/a_2276_472# 0.002066f
C7948 _394_/a_56_524# vss 0.003797f
C7949 fanout55/a_36_160# FILLER_0_13_80/a_36_472# 0.003699f
C7950 net36 vdd 0.939735f
C7951 _142_ FILLER_0_17_142/a_484_472# 0.01467f
C7952 output35/a_224_472# net33 0.170613f
C7953 net5 net8 0.001288f
C7954 net38 _444_/a_796_472# 0.002641f
C7955 FILLER_0_14_99/a_36_472# _095_ 0.011772f
C7956 _044_ _416_/a_2665_112# 0.01372f
C7957 _214_/a_36_160# FILLER_0_23_88/a_124_375# 0.005398f
C7958 FILLER_0_19_28/a_572_375# vss 0.002775f
C7959 FILLER_0_19_28/a_36_472# vdd 0.052986f
C7960 FILLER_0_4_91/a_36_472# _160_ 0.007864f
C7961 _050_ FILLER_0_22_128/a_1020_375# 0.002647f
C7962 output38/a_224_472# _446_/a_448_472# 0.007649f
C7963 _449_/a_2560_156# _067_ 0.007511f
C7964 _098_ FILLER_0_21_150/a_36_472# 0.002964f
C7965 _093_ FILLER_0_19_155/a_36_472# 0.001737f
C7966 FILLER_0_15_2/a_36_472# vss 0.002136f
C7967 FILLER_0_9_223/a_36_472# net4 0.014911f
C7968 _115_ _322_/a_124_24# 0.019655f
C7969 FILLER_0_12_2/a_484_472# vss 0.001748f
C7970 _394_/a_56_524# net74 0.005616f
C7971 _012_ FILLER_0_23_44/a_1020_375# 0.002827f
C7972 _053_ FILLER_0_6_47/a_484_472# 0.006301f
C7973 _080_ net37 0.005467f
C7974 _068_ _117_ 0.011659f
C7975 _436_/a_1000_472# mask\[8\] 0.001091f
C7976 _436_/a_796_472# net35 0.002146f
C7977 _140_ _433_/a_2248_156# 0.003337f
C7978 FILLER_0_20_193/a_572_375# mask\[6\] 0.001262f
C7979 FILLER_0_16_89/a_572_375# vdd 0.005006f
C7980 ctln[4] vdd 0.210384f
C7981 net64 FILLER_0_9_270/a_572_375# 0.017924f
C7982 _417_/a_1204_472# net30 0.001496f
C7983 _417_/a_796_472# result[3] 0.001206f
C7984 net18 rstn 0.015842f
C7985 mask\[2\] FILLER_0_15_235/a_572_375# 0.003879f
C7986 _119_ _153_ 0.001741f
C7987 cal_itt\[3\] _161_ 0.20195f
C7988 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3172_472# 0.013277f
C7989 _430_/a_796_472# _091_ 0.005465f
C7990 _176_ FILLER_0_11_78/a_572_375# 0.013887f
C7991 net54 mask\[9\] 0.094381f
C7992 net31 _277_/a_36_160# 0.053915f
C7993 _030_ _440_/a_36_151# 0.001187f
C7994 _394_/a_56_524# cal_count\[1\] 0.022487f
C7995 mask\[8\] _423_/a_2665_112# 0.004281f
C7996 net35 _423_/a_2248_156# 0.003899f
C7997 net18 _418_/a_1000_472# 0.050485f
C7998 output8/a_224_472# FILLER_0_3_221/a_36_472# 0.001699f
C7999 _394_/a_1336_472# net15 0.01144f
C8000 _103_ _198_/a_67_603# 0.005362f
C8001 _436_/a_1204_472# vdd 0.003143f
C8002 output32/a_224_472# _419_/a_1308_423# 0.005111f
C8003 FILLER_0_14_123/a_124_375# vdd 0.034436f
C8004 output19/a_224_472# vss 0.048948f
C8005 _415_/a_1308_423# net27 0.02437f
C8006 ctlp[1] _420_/a_1308_423# 0.001418f
C8007 mask\[7\] net23 0.225177f
C8008 _440_/a_1000_472# _029_ 0.004334f
C8009 FILLER_0_15_290/a_36_472# net62 0.009046f
C8010 vss _166_ 0.011302f
C8011 vdd _160_ 0.606139f
C8012 net55 FILLER_0_21_60/a_484_472# 0.098472f
C8013 FILLER_0_18_76/a_484_472# vss 0.005065f
C8014 net54 FILLER_0_22_86/a_1380_472# 0.059367f
C8015 _165_ _054_ 0.001337f
C8016 _086_ _163_ 0.413768f
C8017 _069_ state\[1\] 0.003884f
C8018 FILLER_0_21_142/a_36_472# _098_ 0.002964f
C8019 output39/a_224_472# net66 0.009679f
C8020 trim_mask\[1\] FILLER_0_4_91/a_484_472# 0.002806f
C8021 _423_/a_2665_112# vss 0.016881f
C8022 net54 FILLER_0_19_111/a_36_472# 0.003467f
C8023 net72 FILLER_0_17_56/a_124_375# 0.018942f
C8024 FILLER_0_2_101/a_124_375# net14 0.0239f
C8025 trim_val\[4\] FILLER_0_2_165/a_124_375# 0.009193f
C8026 _412_/a_448_472# net19 0.001526f
C8027 net16 net49 0.055931f
C8028 FILLER_0_8_107/a_124_375# FILLER_0_9_105/a_484_472# 0.001684f
C8029 _116_ vdd 0.399137f
C8030 _414_/a_1000_472# net22 0.001649f
C8031 _414_/a_2665_112# _081_ 0.00247f
C8032 mask\[3\] _103_ 0.055796f
C8033 net16 net68 0.275467f
C8034 mask\[5\] vss 0.528441f
C8035 FILLER_0_20_169/a_36_472# vdd 0.010522f
C8036 FILLER_0_20_169/a_124_375# vss 0.017635f
C8037 _136_ FILLER_0_16_154/a_932_472# 0.008185f
C8038 output39/a_224_472# _445_/a_1308_423# 0.010408f
C8039 FILLER_0_1_266/a_484_472# net18 0.010423f
C8040 FILLER_0_1_266/a_572_375# net8 0.016292f
C8041 trimb[4] cal_count\[2\] 0.146942f
C8042 FILLER_0_5_117/a_36_472# _119_ 0.002628f
C8043 FILLER_0_5_117/a_124_375# _086_ 0.003725f
C8044 FILLER_0_12_136/a_1380_472# FILLER_0_13_142/a_572_375# 0.001684f
C8045 net73 FILLER_0_18_139/a_36_472# 0.002491f
C8046 FILLER_0_9_270/a_36_472# vdd 0.008742f
C8047 FILLER_0_9_270/a_572_375# vss 0.017196f
C8048 net64 _223_/a_36_160# 0.007842f
C8049 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1380_472# 0.013276f
C8050 FILLER_0_12_220/a_572_375# _060_ 0.00145f
C8051 net55 FILLER_0_13_80/a_124_375# 0.069951f
C8052 _413_/a_36_151# _088_ 0.001289f
C8053 _163_ _154_ 0.190662f
C8054 FILLER_0_22_128/a_2724_472# _146_ 0.002471f
C8055 _030_ vdd 0.244909f
C8056 fanout82/a_36_113# net37 0.046126f
C8057 ctlp[1] _421_/a_1000_472# 0.007039f
C8058 _427_/a_2248_156# net23 0.033973f
C8059 fanout49/a_36_160# _156_ 0.002871f
C8060 net53 FILLER_0_13_142/a_572_375# 0.001597f
C8061 _442_/a_1204_472# vdd 0.001128f
C8062 _446_/a_1000_472# net17 0.031119f
C8063 _316_/a_124_24# _123_ 0.009391f
C8064 _063_ _444_/a_36_151# 0.030369f
C8065 _020_ vdd 0.194776f
C8066 trim_mask\[1\] vss 0.449335f
C8067 FILLER_0_9_28/a_36_472# net40 0.020589f
C8068 net20 _256_/a_1164_497# 0.001462f
C8069 net47 _382_/a_224_472# 0.001795f
C8070 FILLER_0_5_117/a_124_375# _154_ 0.005866f
C8071 FILLER_0_4_197/a_1380_472# net76 0.003767f
C8072 _424_/a_2248_156# FILLER_0_21_60/a_124_375# 0.001068f
C8073 FILLER_0_15_290/a_124_375# result[3] 0.020277f
C8074 _187_ vdd 0.194575f
C8075 _148_ _025_ 0.007252f
C8076 _055_ _311_/a_1212_473# 0.004259f
C8077 _211_/a_36_160# _050_ 0.010927f
C8078 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_36_472# 0.026657f
C8079 _169_ _163_ 0.013133f
C8080 _086_ _321_/a_3126_472# 0.001522f
C8081 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_124_375# 0.012222f
C8082 FILLER_0_3_54/a_124_375# _164_ 0.008654f
C8083 net73 FILLER_0_18_107/a_572_375# 0.008889f
C8084 FILLER_0_7_72/a_2276_472# _439_/a_2665_112# 0.001167f
C8085 FILLER_0_18_177/a_124_375# FILLER_0_20_177/a_36_472# 0.0027f
C8086 _372_/a_2590_472# _062_ 0.0012f
C8087 mask\[7\] net33 0.02491f
C8088 _425_/a_1308_423# vdd 0.021703f
C8089 _077_ _453_/a_1204_472# 0.011124f
C8090 _104_ result[9] 0.169685f
C8091 _098_ FILLER_0_15_228/a_36_472# 0.022074f
C8092 vdd FILLER_0_3_212/a_124_375# 0.025095f
C8093 net54 _352_/a_49_472# 0.003941f
C8094 FILLER_0_4_177/a_572_375# FILLER_0_5_181/a_124_375# 0.05841f
C8095 mask\[7\] _435_/a_1204_472# 0.007888f
C8096 input1/a_36_113# en 0.036849f
C8097 net70 FILLER_0_11_101/a_484_472# 0.001474f
C8098 net82 net76 0.061682f
C8099 net54 net35 0.114666f
C8100 FILLER_0_18_107/a_1020_375# mask\[9\] 0.005758f
C8101 _091_ FILLER_0_16_154/a_1380_472# 0.00133f
C8102 net72 _174_ 0.199504f
C8103 net65 FILLER_0_1_266/a_124_375# 0.002654f
C8104 _070_ FILLER_0_10_94/a_124_375# 0.008294f
C8105 _223_/a_36_160# vss 0.007187f
C8106 _164_ FILLER_0_6_47/a_484_472# 0.012286f
C8107 _056_ net59 0.001756f
C8108 cal_count\[3\] FILLER_0_12_196/a_124_375# 0.007717f
C8109 mask\[0\] _043_ 0.929722f
C8110 net26 _052_ 0.100927f
C8111 ctln[7] net52 0.06558f
C8112 FILLER_0_5_128/a_36_472# _160_ 0.006214f
C8113 FILLER_0_17_200/a_572_375# _093_ 0.002355f
C8114 _315_/a_716_497# net23 0.004725f
C8115 _117_ vdd 0.050188f
C8116 _056_ net4 0.002408f
C8117 _420_/a_36_151# FILLER_0_23_282/a_36_472# 0.001723f
C8118 FILLER_0_4_107/a_36_472# _153_ 0.042459f
C8119 FILLER_0_4_107/a_932_472# _154_ 0.017867f
C8120 FILLER_0_14_99/a_36_472# vss 0.003598f
C8121 mask\[5\] FILLER_0_18_177/a_1828_472# 0.001038f
C8122 _253_/a_36_68# vss 0.002481f
C8123 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_484_472# 0.001723f
C8124 _415_/a_36_151# _004_ 0.013592f
C8125 _057_ _116_ 0.028033f
C8126 FILLER_0_7_162/a_124_375# calibrate 0.014255f
C8127 _149_ FILLER_0_20_87/a_36_472# 0.001938f
C8128 net32 _421_/a_2665_112# 0.019532f
C8129 _061_ _311_/a_66_473# 0.030169f
C8130 _073_ _260_/a_36_68# 0.079772f
C8131 net63 FILLER_0_15_228/a_36_472# 0.001669f
C8132 trim_val\[4\] net59 0.062701f
C8133 _053_ FILLER_0_6_177/a_36_472# 0.00572f
C8134 _170_ _241_/a_224_472# 0.001199f
C8135 FILLER_0_16_57/a_124_375# _176_ 0.015872f
C8136 _095_ cal_count\[2\] 0.270066f
C8137 _414_/a_36_151# FILLER_0_7_195/a_124_375# 0.059049f
C8138 output45/a_224_472# vdd -0.026726f
C8139 FILLER_0_24_63/a_36_472# ctlp[9] 0.012298f
C8140 FILLER_0_18_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001684f
C8141 result[6] vdd 0.513079f
C8142 _434_/a_796_472# mask\[6\] 0.004416f
C8143 FILLER_0_16_255/a_36_472# _094_ 0.005892f
C8144 net31 _102_ 0.060034f
C8145 FILLER_0_20_193/a_572_375# net35 0.002196f
C8146 result[9] _421_/a_1308_423# 0.011854f
C8147 output25/a_224_472# _051_ 0.019651f
C8148 net79 _416_/a_1308_423# 0.030119f
C8149 net70 FILLER_0_18_107/a_1380_472# 0.00116f
C8150 FILLER_0_3_142/a_36_472# net23 0.043034f
C8151 FILLER_0_8_247/a_124_375# vss 0.002674f
C8152 _058_ _055_ 0.070216f
C8153 FILLER_0_8_247/a_572_375# vdd -0.007963f
C8154 _421_/a_36_151# vdd -0.053849f
C8155 _032_ _152_ 0.001206f
C8156 mask\[0\] net21 0.050431f
C8157 _155_ FILLER_0_8_107/a_36_472# 0.002068f
C8158 net44 _039_ 0.15647f
C8159 _074_ net21 0.186175f
C8160 mask\[3\] _019_ 0.001403f
C8161 _189_/a_67_603# net79 0.008944f
C8162 net15 _120_ 0.028275f
C8163 FILLER_0_12_220/a_484_472# _070_ 0.004091f
C8164 output36/a_224_472# FILLER_0_15_282/a_36_472# 0.008834f
C8165 _225_/a_36_160# vdd 0.058272f
C8166 ctlp[3] _422_/a_2560_156# 0.001006f
C8167 output12/a_224_472# net11 0.009336f
C8168 cal_count\[3\] _389_/a_428_148# 0.001072f
C8169 _444_/a_1204_472# net40 0.017496f
C8170 fanout51/a_36_113# _120_ 0.014349f
C8171 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_572_375# 0.086635f
C8172 cal_itt\[1\] net18 0.026586f
C8173 FILLER_0_20_193/a_484_472# vdd 0.00749f
C8174 FILLER_0_20_193/a_36_472# vss 0.001978f
C8175 net19 net30 0.311153f
C8176 net58 net19 0.044785f
C8177 fanout74/a_36_113# FILLER_0_3_142/a_36_472# 0.016516f
C8178 FILLER_0_16_73/a_36_472# _175_ 0.006803f
C8179 _446_/a_36_151# net40 0.015376f
C8180 output42/a_224_472# net6 0.010571f
C8181 FILLER_0_17_72/a_2724_472# _131_ 0.004095f
C8182 _074_ _375_/a_960_497# 0.004175f
C8183 _035_ net47 0.101683f
C8184 _116_ _279_/a_244_68# 0.001752f
C8185 FILLER_0_9_105/a_484_472# vss 0.004412f
C8186 net32 net22 0.042885f
C8187 _196_/a_36_160# FILLER_0_14_263/a_36_472# 0.004828f
C8188 _410_/a_36_68# net51 0.014342f
C8189 FILLER_0_5_198/a_36_472# net59 0.059378f
C8190 _305_/a_36_159# _316_/a_124_24# 0.003478f
C8191 net10 output11/a_224_472# 0.095679f
C8192 _058_ _313_/a_67_603# 0.010094f
C8193 FILLER_0_18_139/a_932_472# vss 0.041568f
C8194 FILLER_0_18_139/a_1380_472# vdd 0.005855f
C8195 trim[2] trim[3] 0.056575f
C8196 _093_ _334_/a_36_160# 0.014676f
C8197 net65 FILLER_0_3_172/a_2364_375# 0.003745f
C8198 fanout57/a_36_113# FILLER_0_3_172/a_36_472# 0.19419f
C8199 valid net18 0.03851f
C8200 net63 _435_/a_36_151# 0.017194f
C8201 FILLER_0_16_154/a_1020_375# vss 0.001453f
C8202 FILLER_0_16_154/a_1468_375# vdd 0.017574f
C8203 _412_/a_1308_423# cal_itt\[1\] 0.009991f
C8204 FILLER_0_5_72/a_1020_375# _440_/a_2248_156# 0.001068f
C8205 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_124_375# 0.012001f
C8206 _091_ FILLER_0_12_220/a_932_472# 0.001638f
C8207 FILLER_0_7_72/a_3172_472# _058_ 0.001085f
C8208 mask\[7\] FILLER_0_22_128/a_1828_472# 0.004503f
C8209 _057_ _117_ 0.120323f
C8210 FILLER_0_17_64/a_36_472# net36 0.00195f
C8211 FILLER_0_8_127/a_36_472# _125_ 0.003088f
C8212 ctlp[7] net54 0.004355f
C8213 FILLER_0_7_104/a_1020_375# vdd 0.010571f
C8214 mask\[5\] FILLER_0_21_206/a_124_375# 0.011644f
C8215 trim_val\[2\] _167_ 0.011787f
C8216 _076_ net47 0.00115f
C8217 _144_ _348_/a_257_69# 0.001978f
C8218 net20 _429_/a_2665_112# 0.062922f
C8219 FILLER_0_7_146/a_124_375# calibrate 0.014163f
C8220 FILLER_0_12_2/a_124_375# net67 0.003339f
C8221 _436_/a_448_472# _050_ 0.064832f
C8222 FILLER_0_5_164/a_124_375# _066_ 0.006762f
C8223 _120_ net51 1.716752f
C8224 FILLER_0_17_72/a_1916_375# net53 0.001657f
C8225 trim[0] _034_ 0.044322f
C8226 vdd _156_ 0.178622f
C8227 FILLER_0_18_107/a_1916_375# vdd 0.018831f
C8228 trim_val\[1\] FILLER_0_6_47/a_124_375# 0.002577f
C8229 _413_/a_1308_423# vdd 0.002686f
C8230 net65 _264_/a_224_472# 0.001866f
C8231 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_124_375# 0.012552f
C8232 net82 _083_ 0.010347f
C8233 _365_/a_244_472# _156_ 0.003847f
C8234 _177_ _095_ 0.004392f
C8235 _207_/a_67_603# FILLER_0_22_128/a_3172_472# 0.005759f
C8236 mask\[4\] vdd 0.794539f
C8237 _432_/a_2560_156# net80 0.01523f
C8238 net52 FILLER_0_2_165/a_36_472# 0.002601f
C8239 _448_/a_448_472# net22 0.085004f
C8240 net54 FILLER_0_22_128/a_1468_375# 0.004731f
C8241 net9 _082_ 0.001006f
C8242 _432_/a_2248_156# mask\[3\] 0.002775f
C8243 net67 vdd 0.638702f
C8244 result[9] FILLER_0_24_274/a_932_472# 0.001826f
C8245 trim[4] net39 0.004535f
C8246 FILLER_0_16_57/a_124_375# _183_ 0.005825f
C8247 _317_/a_36_113# vdd 0.054289f
C8248 FILLER_0_10_37/a_36_472# net16 0.012905f
C8249 net16 _408_/a_1936_472# 0.022235f
C8250 net69 _159_ 0.010086f
C8251 _187_ cal_count\[0\] 0.645851f
C8252 FILLER_0_24_274/a_36_472# vdd 0.107635f
C8253 FILLER_0_24_274/a_1468_375# vss 0.060201f
C8254 _093_ net36 0.214976f
C8255 FILLER_0_22_86/a_484_472# _437_/a_448_472# 0.008036f
C8256 _430_/a_2248_156# FILLER_0_15_212/a_932_472# 0.035805f
C8257 _414_/a_796_472# vdd 0.001497f
C8258 FILLER_0_5_72/a_1380_472# vss 0.004538f
C8259 _422_/a_36_151# net19 0.033614f
C8260 _098_ net14 0.061285f
C8261 net63 FILLER_0_17_200/a_484_472# 0.003767f
C8262 _057_ _225_/a_36_160# 0.026341f
C8263 FILLER_0_24_274/a_932_472# FILLER_0_23_282/a_36_472# 0.05841f
C8264 net16 _184_ 0.028159f
C8265 _029_ _153_ 0.023421f
C8266 output45/a_224_472# output17/a_224_472# 0.071473f
C8267 _345_/a_36_160# net73 0.032139f
C8268 net65 _002_ 0.042811f
C8269 FILLER_0_5_164/a_124_375# net37 0.008158f
C8270 sample fanout64/a_36_160# 0.007266f
C8271 _390_/a_36_68# vss 0.002334f
C8272 net79 _056_ 0.022406f
C8273 _118_ _059_ 0.022651f
C8274 _025_ FILLER_0_22_107/a_124_375# 0.001891f
C8275 _093_ FILLER_0_16_89/a_572_375# 0.002889f
C8276 FILLER_0_10_37/a_124_375# vdd 0.048346f
C8277 _415_/a_1000_472# vdd 0.002497f
C8278 _092_ FILLER_0_17_218/a_572_375# 0.006125f
C8279 _053_ net59 0.145863f
C8280 _124_ FILLER_0_10_107/a_484_472# 0.00438f
C8281 net10 _411_/a_2665_112# 0.007912f
C8282 state\[1\] _090_ 0.087906f
C8283 _397_/a_36_472# net55 0.039732f
C8284 output10/a_224_472# FILLER_0_0_266/a_36_472# 0.023414f
C8285 fanout82/a_36_113# _122_ 0.007118f
C8286 net16 FILLER_0_8_37/a_36_472# 0.012905f
C8287 cal_count\[3\] _067_ 0.478427f
C8288 _420_/a_796_472# _009_ 0.012395f
C8289 mask\[0\] FILLER_0_15_212/a_1020_375# 0.001158f
C8290 _054_ vss 0.176655f
C8291 _016_ _427_/a_36_151# 0.00483f
C8292 _053_ net4 0.013559f
C8293 net74 _390_/a_36_68# 0.008011f
C8294 cal_count\[2\] vss 0.361185f
C8295 _099_ FILLER_0_14_235/a_572_375# 0.013281f
C8296 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_124_375# 0.026339f
C8297 net18 _416_/a_36_151# 0.027435f
C8298 FILLER_0_8_24/a_36_472# vss 0.001239f
C8299 FILLER_0_8_24/a_484_472# vdd 0.009032f
C8300 _443_/a_36_151# net13 0.001896f
C8301 _443_/a_1308_423# net23 0.034115f
C8302 FILLER_0_3_78/a_572_375# _160_ 0.003506f
C8303 net50 _441_/a_1000_472# 0.02354f
C8304 net52 _441_/a_2248_156# 0.023959f
C8305 FILLER_0_12_220/a_1020_375# vdd -0.014642f
C8306 FILLER_0_12_220/a_572_375# vss 0.007775f
C8307 _104_ net61 1.149805f
C8308 _015_ net4 0.003985f
C8309 FILLER_0_15_150/a_124_375# _427_/a_448_472# 0.008952f
C8310 FILLER_0_4_49/a_36_472# net66 0.012791f
C8311 FILLER_0_13_212/a_36_472# net79 0.006158f
C8312 net55 FILLER_0_18_37/a_124_375# 0.005899f
C8313 FILLER_0_4_107/a_1468_375# _160_ 0.028099f
C8314 net50 _447_/a_448_472# 0.001219f
C8315 state\[1\] net22 0.007096f
C8316 FILLER_0_17_72/a_124_375# vdd 0.0132f
C8317 FILLER_0_8_37/a_124_375# vss 0.00252f
C8318 FILLER_0_8_37/a_572_375# vdd 0.013575f
C8319 _155_ _365_/a_36_68# 0.053708f
C8320 _345_/a_36_160# FILLER_0_19_111/a_484_472# 0.007907f
C8321 net47 FILLER_0_4_91/a_572_375# 0.008167f
C8322 net75 net37 0.07785f
C8323 FILLER_0_11_124/a_36_472# vss 0.002545f
C8324 _274_/a_1612_497# net4 0.00807f
C8325 net50 _439_/a_796_472# 0.002389f
C8326 net52 _439_/a_1204_472# 0.027632f
C8327 output12/a_224_472# ctln[5] 0.069673f
C8328 _070_ FILLER_0_11_109/a_124_375# 0.002358f
C8329 trimb[1] FILLER_0_18_2/a_572_375# 0.010125f
C8330 _053_ FILLER_0_7_72/a_2724_472# 0.016187f
C8331 _141_ _049_ 0.0035f
C8332 _425_/a_1000_472# net37 0.002879f
C8333 mask\[4\] FILLER_0_18_177/a_1380_472# 0.016924f
C8334 net38 _450_/a_36_151# 0.035458f
C8335 output18/a_224_472# vss 0.086897f
C8336 fanout57/a_36_113# FILLER_0_2_165/a_124_375# 0.008057f
C8337 net28 net36 0.002537f
C8338 cal_count\[2\] cal_count\[1\] 0.067712f
C8339 net16 net47 0.089651f
C8340 _434_/a_1204_472# vdd 0.005382f
C8341 _340_/a_36_160# vss 0.029871f
C8342 net74 FILLER_0_11_124/a_36_472# 0.020589f
C8343 output11/a_224_472# ctln[4] 0.072677f
C8344 mask\[8\] _437_/a_36_151# 0.005179f
C8345 FILLER_0_12_136/a_1468_375# vdd 0.026145f
C8346 _422_/a_36_151# _009_ 0.015085f
C8347 ctlp[1] FILLER_0_23_282/a_124_375# 0.00324f
C8348 _417_/a_448_472# vss 0.005289f
C8349 _417_/a_1308_423# vdd 0.002263f
C8350 FILLER_0_12_136/a_1020_375# vss 0.018233f
C8351 net49 FILLER_0_3_78/a_124_375# 0.001597f
C8352 _030_ FILLER_0_3_78/a_572_375# 0.007667f
C8353 _053_ FILLER_0_7_162/a_36_472# 0.004888f
C8354 _068_ _059_ 0.255081f
C8355 _012_ FILLER_0_23_60/a_124_375# 0.002827f
C8356 net69 FILLER_0_2_111/a_932_472# 0.011453f
C8357 _031_ FILLER_0_2_111/a_36_472# 0.034656f
C8358 _065_ _064_ 0.007356f
C8359 _144_ _437_/a_2665_112# 0.001186f
C8360 net58 fanout58/a_36_160# 0.013794f
C8361 result[6] net60 0.094624f
C8362 result[6] net78 0.027123f
C8363 net58 cal_itt\[0\] 0.229955f
C8364 _132_ _145_ 0.010994f
C8365 _065_ _447_/a_1204_472# 0.017675f
C8366 _069_ FILLER_0_13_206/a_36_472# 0.005793f
C8367 _072_ FILLER_0_7_233/a_36_472# 0.00241f
C8368 FILLER_0_7_195/a_124_375# net21 0.007906f
C8369 _104_ _108_ 0.02837f
C8370 FILLER_0_4_123/a_36_472# _370_/a_124_24# 0.003595f
C8371 net78 _421_/a_36_151# 0.001368f
C8372 net60 _421_/a_36_151# 0.224039f
C8373 _020_ _093_ 0.015474f
C8374 _164_ net40 0.048933f
C8375 _086_ _121_ 0.049499f
C8376 _437_/a_448_472# vdd 0.010432f
C8377 _437_/a_36_151# vss 0.006865f
C8378 FILLER_0_10_28/a_36_472# net6 0.038613f
C8379 trim_mask\[2\] _164_ 1.859062f
C8380 cal input1/a_36_113# 0.025739f
C8381 output19/a_224_472# _295_/a_36_472# 0.003896f
C8382 _424_/a_448_472# FILLER_0_18_37/a_1020_375# 0.001674f
C8383 _447_/a_1308_423# _164_ 0.001422f
C8384 result[7] result[9] 1.21288f
C8385 _063_ net49 0.002854f
C8386 _079_ FILLER_0_5_212/a_124_375# 0.005363f
C8387 net18 net59 0.695067f
C8388 _322_/a_848_380# _062_ 0.001872f
C8389 net80 mask\[3\] 0.02972f
C8390 net44 clkc 0.184915f
C8391 cal_count\[3\] _121_ 0.011368f
C8392 FILLER_0_14_91/a_572_375# _095_ 0.011885f
C8393 _322_/a_1084_68# _118_ 0.002515f
C8394 FILLER_0_14_81/a_124_375# _177_ 0.002725f
C8395 net34 vdd 1.161282f
C8396 _424_/a_2665_112# net36 0.028938f
C8397 net4 net18 0.034592f
C8398 _086_ FILLER_0_7_104/a_124_375# 0.001629f
C8399 _326_/a_36_160# vdd 0.066545f
C8400 FILLER_0_7_72/a_2276_472# net50 0.030391f
C8401 FILLER_0_23_44/a_1020_375# vdd -0.014642f
C8402 net54 _433_/a_1308_423# 0.004372f
C8403 mask\[5\] FILLER_0_19_195/a_124_375# 0.007169f
C8404 net81 FILLER_0_15_212/a_932_472# 0.003953f
C8405 result[7] FILLER_0_23_282/a_36_472# 0.014869f
C8406 _177_ vss 0.074896f
C8407 _446_/a_36_151# trim[3] 0.00699f
C8408 mask\[5\] _295_/a_36_472# 0.034027f
C8409 net38 _178_ 0.123812f
C8410 _017_ FILLER_0_14_107/a_484_472# 0.004583f
C8411 _354_/a_49_472# net71 0.010421f
C8412 net70 FILLER_0_14_107/a_1380_472# 0.003355f
C8413 output47/a_224_472# net38 0.082174f
C8414 FILLER_0_16_57/a_36_472# cal_count\[2\] 0.001952f
C8415 FILLER_0_18_2/a_3172_472# FILLER_0_19_28/a_124_375# 0.001684f
C8416 ctln[5] net12 0.41364f
C8417 net15 FILLER_0_5_54/a_932_472# 0.008904f
C8418 _067_ FILLER_0_12_20/a_124_375# 0.017026f
C8419 _105_ net22 0.01308f
C8420 FILLER_0_20_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001543f
C8421 net72 FILLER_0_15_59/a_124_375# 0.022905f
C8422 _412_/a_1308_423# net59 0.00291f
C8423 _131_ net14 0.037705f
C8424 FILLER_0_4_177/a_484_472# net76 0.006746f
C8425 FILLER_0_4_152/a_124_375# net47 0.009228f
C8426 _074_ _062_ 0.005012f
C8427 net20 _094_ 0.677838f
C8428 _416_/a_36_151# net62 0.054002f
C8429 output21/a_224_472# net33 0.001166f
C8430 FILLER_0_17_38/a_484_472# vss 0.001229f
C8431 _084_ _082_ 0.044645f
C8432 _100_ _283_/a_36_472# 0.033597f
C8433 _098_ _433_/a_2248_156# 0.034774f
C8434 FILLER_0_18_2/a_932_472# net44 0.012286f
C8435 FILLER_0_1_98/a_36_472# net52 0.005688f
C8436 net17 _450_/a_3129_107# 0.004255f
C8437 _430_/a_36_151# _139_ 0.012035f
C8438 _028_ FILLER_0_5_72/a_572_375# 0.00123f
C8439 _230_/a_244_68# _070_ 0.001641f
C8440 FILLER_0_16_241/a_36_472# _099_ 0.158391f
C8441 _114_ net14 0.127764f
C8442 _077_ _439_/a_448_472# 0.052962f
C8443 net47 _452_/a_1353_112# 0.003681f
C8444 _442_/a_2248_156# _158_ 0.001288f
C8445 _096_ _090_ 0.026104f
C8446 mask\[9\] _438_/a_2248_156# 0.036436f
C8447 _236_/a_36_160# net39 0.052649f
C8448 FILLER_0_5_181/a_124_375# net22 0.00205f
C8449 _395_/a_36_488# _176_ 0.010116f
C8450 _395_/a_1044_488# _085_ 0.00391f
C8451 net19 _417_/a_2665_112# 0.042961f
C8452 _177_ cal_count\[1\] 0.03631f
C8453 FILLER_0_3_172/a_3260_375# net22 0.015274f
C8454 _136_ FILLER_0_16_115/a_124_375# 0.006372f
C8455 ctln[8] _168_ 0.001145f
C8456 trim[4] net42 0.016428f
C8457 _427_/a_36_151# _043_ 0.002267f
C8458 fanout57/a_36_113# net59 0.00178f
C8459 comp FILLER_0_15_2/a_36_472# 0.001941f
C8460 net31 mask\[5\] 0.017182f
C8461 _429_/a_796_472# _018_ 0.002291f
C8462 cal_itt\[3\] _056_ 0.023192f
C8463 _053_ FILLER_0_7_146/a_36_472# 0.001014f
C8464 fanout75/a_36_113# net59 0.00817f
C8465 _322_/a_1084_68# _068_ 0.001022f
C8466 _052_ FILLER_0_18_53/a_572_375# 0.001631f
C8467 trimb[1] _452_/a_3129_107# 0.007229f
C8468 _095_ _402_/a_56_567# 0.010012f
C8469 ctln[3] _411_/a_448_472# 0.00336f
C8470 output10/a_224_472# _411_/a_2248_156# 0.019736f
C8471 FILLER_0_19_171/a_1380_472# FILLER_0_19_187/a_36_472# 0.013277f
C8472 FILLER_0_10_37/a_124_375# cal_count\[0\] 0.016543f
C8473 FILLER_0_5_128/a_572_375# net47 0.010055f
C8474 net50 FILLER_0_7_59/a_484_472# 0.011974f
C8475 _412_/a_1204_472# net76 0.020975f
C8476 net15 _043_ 0.042278f
C8477 _448_/a_36_151# vdd 0.133302f
C8478 output38/a_224_472# _035_ 0.091395f
C8479 _265_/a_244_68# _084_ 0.016463f
C8480 _359_/a_36_488# _129_ 0.002527f
C8481 _098_ FILLER_0_20_87/a_36_472# 0.016138f
C8482 net57 net36 0.087967f
C8483 net11 vss 0.057193f
C8484 net19 _192_/a_67_603# 0.003106f
C8485 net36 FILLER_0_15_205/a_36_472# 0.005101f
C8486 FILLER_0_14_107/a_124_375# vdd 0.013327f
C8487 _059_ vdd 0.161836f
C8488 _431_/a_1308_423# _137_ 0.008805f
C8489 output37/a_224_472# vdd 0.082206f
C8490 _086_ FILLER_0_11_124/a_124_375# 0.016039f
C8491 FILLER_0_22_177/a_124_375# vdd 0.001293f
C8492 net69 _441_/a_1308_423# 0.016223f
C8493 _086_ _115_ 0.4112f
C8494 _185_ _180_ 0.001053f
C8495 _414_/a_36_151# _163_ 0.001186f
C8496 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_572_375# 0.086635f
C8497 _093_ FILLER_0_18_139/a_1380_472# 0.007013f
C8498 cal_itt\[2\] FILLER_0_3_221/a_124_375# 0.006217f
C8499 _064_ _036_ 0.003286f
C8500 trim_mask\[2\] trim_val\[3\] 0.003342f
C8501 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_124_375# 0.012222f
C8502 _375_/a_36_68# vdd 0.010344f
C8503 net71 _437_/a_796_472# 0.006933f
C8504 net5 vdd 0.516129f
C8505 FILLER_0_12_136/a_1380_472# _127_ 0.001432f
C8506 net63 FILLER_0_17_218/a_124_375# 0.040329f
C8507 _445_/a_448_472# net66 0.010949f
C8508 _064_ _445_/a_2665_112# 0.004701f
C8509 cal_count\[3\] FILLER_0_11_124/a_124_375# 0.002147f
C8510 FILLER_0_7_72/a_1380_472# _077_ 0.001315f
C8511 FILLER_0_18_107/a_1916_375# _433_/a_36_151# 0.002709f
C8512 FILLER_0_20_177/a_1380_472# vss 0.004504f
C8513 _127_ FILLER_0_9_142/a_124_375# 0.005447f
C8514 _115_ cal_count\[3\] 0.004426f
C8515 _175_ net15 0.052586f
C8516 net65 net76 0.14935f
C8517 FILLER_0_7_195/a_36_472# _074_ 0.008706f
C8518 ctlp[2] net33 0.004972f
C8519 _436_/a_1308_423# net54 0.002665f
C8520 FILLER_0_18_100/a_36_472# _136_ 0.003419f
C8521 _127_ net53 0.00917f
C8522 _155_ _154_ 0.18488f
C8523 _029_ trim_mask\[1\] 1.002118f
C8524 _450_/a_448_472# net6 0.041113f
C8525 _308_/a_124_24# _114_ 0.052818f
C8526 FILLER_0_12_136/a_1020_375# FILLER_0_11_142/a_484_472# 0.001543f
C8527 _439_/a_2248_156# trim_mask\[0\] 0.005416f
C8528 cal_itt\[3\] FILLER_0_5_198/a_36_472# 0.07099f
C8529 FILLER_0_10_78/a_484_472# net52 0.004421f
C8530 FILLER_0_12_136/a_572_375# cal_count\[3\] 0.005006f
C8531 _126_ net14 0.238336f
C8532 _068_ _247_/a_36_160# 0.003213f
C8533 FILLER_0_18_177/a_1468_375# vdd 0.024167f
C8534 _132_ _428_/a_448_472# 0.034825f
C8535 _350_/a_49_472# mask\[6\] 0.033488f
C8536 FILLER_0_2_101/a_36_472# _156_ 0.001487f
C8537 net82 FILLER_0_3_212/a_36_472# 0.011542f
C8538 result[7] FILLER_0_24_290/a_124_375# 0.005026f
C8539 _418_/a_448_472# vss 0.005772f
C8540 _418_/a_1308_423# vdd 0.002258f
C8541 _411_/a_796_472# _000_ 0.044697f
C8542 _411_/a_1204_472# net75 0.008304f
C8543 _070_ FILLER_0_8_156/a_124_375# 0.004329f
C8544 _419_/a_2665_112# vdd 0.030085f
C8545 _136_ _451_/a_2225_156# 0.01289f
C8546 _076_ _385_/a_36_68# 0.006512f
C8547 net41 _444_/a_1000_472# 0.002179f
C8548 FILLER_0_14_91/a_36_472# vdd 0.08739f
C8549 FILLER_0_14_91/a_572_375# vss 0.054783f
C8550 mask\[4\] _093_ 0.469687f
C8551 net79 net18 0.222939f
C8552 FILLER_0_20_2/a_484_472# net43 0.005543f
C8553 FILLER_0_12_136/a_1380_472# _071_ 0.004003f
C8554 FILLER_0_18_100/a_36_472# _356_/a_36_472# 0.010679f
C8555 _453_/a_2248_156# vdd 0.010767f
C8556 _026_ _437_/a_36_151# 0.012193f
C8557 _149_ _437_/a_1308_423# 0.015677f
C8558 net57 _116_ 0.069858f
C8559 _095_ _451_/a_1040_527# 0.002316f
C8560 _091_ _273_/a_36_68# 0.00155f
C8561 _144_ net71 0.039862f
C8562 _012_ FILLER_0_21_60/a_572_375# 0.011991f
C8563 output47/a_224_472# net55 0.160037f
C8564 net75 _122_ 0.052177f
C8565 _002_ _079_ 0.051048f
C8566 _077_ _319_/a_672_472# 0.001602f
C8567 FILLER_0_10_214/a_124_375# _070_ 0.017713f
C8568 _072_ net4 0.097916f
C8569 FILLER_0_15_212/a_36_472# mask\[1\] 0.006865f
C8570 FILLER_0_13_142/a_572_375# net23 0.009573f
C8571 _425_/a_1204_472# calibrate 0.009749f
C8572 _089_ net37 0.0326f
C8573 FILLER_0_20_2/a_124_375# vss 0.002737f
C8574 FILLER_0_20_2/a_572_375# vdd 0.010844f
C8575 _290_/a_224_472# net18 0.00868f
C8576 FILLER_0_5_212/a_124_375# vss 0.006344f
C8577 FILLER_0_5_212/a_36_472# vdd 0.107657f
C8578 FILLER_0_18_177/a_2724_472# net21 0.048803f
C8579 _438_/a_2560_156# vdd 0.001166f
C8580 _438_/a_2665_112# vss 0.001389f
C8581 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_36_472# 0.026657f
C8582 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_572_375# 0.001597f
C8583 FILLER_0_13_212/a_1020_375# net62 0.001597f
C8584 trim_val\[1\] vdd 0.173304f
C8585 FILLER_0_1_266/a_572_375# vdd 0.030477f
C8586 _087_ FILLER_0_6_177/a_124_375# 0.001151f
C8587 _408_/a_56_524# FILLER_0_12_20/a_572_375# 0.009967f
C8588 FILLER_0_9_28/a_1380_472# net68 0.008573f
C8589 mask\[5\] net80 0.036014f
C8590 net80 FILLER_0_20_169/a_124_375# 0.054969f
C8591 net20 _258_/a_36_160# 0.041584f
C8592 mask\[7\] _109_ 0.028117f
C8593 _255_/a_224_552# _162_ 0.010564f
C8594 _057_ _375_/a_36_68# 0.003063f
C8595 _077_ net14 0.03359f
C8596 _091_ FILLER_0_10_214/a_36_472# 0.001357f
C8597 net20 output34/a_224_472# 0.023142f
C8598 net75 FILLER_0_6_231/a_484_472# 0.003485f
C8599 result[7] net61 0.021122f
C8600 net48 _068_ 0.054333f
C8601 _074_ _316_/a_124_24# 0.018608f
C8602 _176_ _125_ 0.089769f
C8603 result[8] FILLER_0_24_274/a_484_472# 0.005458f
C8604 net50 FILLER_0_6_90/a_484_472# 0.012286f
C8605 net72 _217_/a_36_160# 0.068583f
C8606 FILLER_0_6_47/a_2812_375# vss 0.035758f
C8607 FILLER_0_6_47/a_3260_375# vdd 0.003435f
C8608 _067_ _120_ 0.031156f
C8609 FILLER_0_7_195/a_124_375# _062_ 0.001983f
C8610 FILLER_0_15_212/a_36_472# vss 0.002853f
C8611 FILLER_0_1_98/a_124_375# trim_val\[3\] 0.001628f
C8612 _151_ _163_ 0.501188f
C8613 trim_mask\[4\] _386_/a_124_24# 0.040347f
C8614 net2 net5 0.47659f
C8615 _053_ cal_itt\[3\] 0.471909f
C8616 _182_ FILLER_0_18_37/a_1380_472# 0.004074f
C8617 FILLER_0_18_2/a_484_472# output47/a_224_472# 0.00175f
C8618 net53 _451_/a_2449_156# 0.015332f
C8619 FILLER_0_6_239/a_36_472# _316_/a_124_24# 0.002228f
C8620 _009_ FILLER_0_23_282/a_572_375# 0.016879f
C8621 FILLER_0_4_197/a_572_375# net22 0.016547f
C8622 _323_/a_36_113# _426_/a_2248_156# 0.001661f
C8623 _127_ FILLER_0_11_135/a_36_472# 0.044488f
C8624 FILLER_0_8_247/a_36_472# calibrate 0.008647f
C8625 net19 net9 0.342451f
C8626 _421_/a_2248_156# mask\[7\] 0.016229f
C8627 net19 _418_/a_2665_112# 0.040822f
C8628 _081_ net23 0.081773f
C8629 _077_ FILLER_0_10_78/a_572_375# 0.001886f
C8630 FILLER_0_17_104/a_932_472# net14 0.002113f
C8631 output25/a_224_472# net24 0.002325f
C8632 _419_/a_796_472# net77 0.001053f
C8633 ctln[5] vss 0.132862f
C8634 net20 _043_ 0.094689f
C8635 _422_/a_448_472# mask\[7\] 0.048658f
C8636 _159_ vss 0.102545f
C8637 net52 _443_/a_796_472# 0.004334f
C8638 net72 _038_ 0.013821f
C8639 _168_ vdd 0.083621f
C8640 _426_/a_448_472# calibrate 0.002745f
C8641 _176_ _174_ 0.00677f
C8642 output26/a_224_472# vdd 0.047141f
C8643 net29 _099_ 0.358926f
C8644 result[7] _108_ 0.063624f
C8645 FILLER_0_13_206/a_36_472# net22 0.053292f
C8646 _077_ FILLER_0_9_72/a_484_472# 0.004472f
C8647 net15 FILLER_0_6_47/a_1916_375# 0.029774f
C8648 _453_/a_1000_472# _042_ 0.004985f
C8649 fanout53/a_36_160# _427_/a_2248_156# 0.027388f
C8650 net74 _159_ 0.129233f
C8651 net79 net62 1.615103f
C8652 FILLER_0_18_53/a_36_472# vss 0.001471f
C8653 FILLER_0_18_53/a_484_472# vdd 0.002358f
C8654 cal net8 0.271166f
C8655 _415_/a_1308_423# result[1] 0.00761f
C8656 FILLER_0_16_89/a_1020_375# _131_ 0.015706f
C8657 output33/a_224_472# result[6] 0.035032f
C8658 _433_/a_1000_472# _022_ 0.05526f
C8659 fanout68/a_36_113# net68 0.027807f
C8660 FILLER_0_4_107/a_1020_375# net47 0.011446f
C8661 _008_ _099_ 0.006163f
C8662 _430_/a_36_151# net63 0.026607f
C8663 FILLER_0_3_221/a_124_375# net59 0.008996f
C8664 _247_/a_36_160# vdd 0.060423f
C8665 FILLER_0_4_197/a_36_472# _270_/a_36_472# 0.004546f
C8666 _217_/a_36_160# _424_/a_36_151# 0.035111f
C8667 _104_ FILLER_0_17_226/a_36_472# 0.013926f
C8668 FILLER_0_21_28/a_124_375# vdd 0.014155f
C8669 _178_ FILLER_0_15_10/a_36_472# 0.001356f
C8670 net69 net14 0.056927f
C8671 output12/a_224_472# net76 0.00803f
C8672 FILLER_0_3_172/a_2812_375# vdd -0.012025f
C8673 valid fanout59/a_36_160# 0.029107f
C8674 net34 _147_ 0.144404f
C8675 _065_ net50 0.123581f
C8676 _449_/a_1308_423# net55 0.001985f
C8677 output47/a_224_472# FILLER_0_15_10/a_36_472# 0.038484f
C8678 _429_/a_36_151# _136_ 0.001188f
C8679 FILLER_0_4_177/a_36_472# FILLER_0_2_177/a_124_375# 0.001512f
C8680 _053_ _257_/a_244_68# 0.001138f
C8681 net4 FILLER_0_3_221/a_124_375# 0.015788f
C8682 _438_/a_1308_423# net14 0.005201f
C8683 FILLER_0_8_239/a_36_472# calibrate 0.008683f
C8684 FILLER_0_10_78/a_1380_472# _176_ 0.009351f
C8685 _431_/a_36_151# FILLER_0_18_107/a_3172_472# 0.00271f
C8686 fanout62/a_36_160# net64 0.052109f
C8687 FILLER_0_17_56/a_124_375# _183_ 0.019253f
C8688 net50 FILLER_0_5_88/a_124_375# 0.03181f
C8689 _077_ _308_/a_124_24# 0.018118f
C8690 _068_ _229_/a_224_472# 0.002601f
C8691 _131_ FILLER_0_14_123/a_36_472# 0.029747f
C8692 net34 _093_ 0.005701f
C8693 FILLER_0_17_72/a_2276_472# mask\[9\] 0.006767f
C8694 _446_/a_2248_156# net66 0.002766f
C8695 net57 _225_/a_36_160# 0.022745f
C8696 _063_ net47 0.142088f
C8697 net52 _387_/a_36_113# 0.02405f
C8698 _112_ calibrate 0.024557f
C8699 FILLER_0_5_72/a_1020_375# net49 0.002208f
C8700 _062_ _226_/a_452_68# 0.001697f
C8701 _129_ _160_ 0.001631f
C8702 _005_ _416_/a_1308_423# 0.020096f
C8703 _443_/a_36_151# _170_ 0.014771f
C8704 fanout64/a_36_160# calibrate 0.001117f
C8705 _132_ FILLER_0_17_104/a_124_375# 0.001918f
C8706 _297_/a_36_472# vss 0.003601f
C8707 net76 FILLER_0_3_172/a_124_375# 0.001186f
C8708 en_co_clk FILLER_0_13_100/a_36_472# 0.001752f
C8709 FILLER_0_19_47/a_36_472# _052_ 0.015772f
C8710 FILLER_0_16_73/a_484_472# net15 0.001946f
C8711 _121_ _120_ 0.069685f
C8712 _451_/a_836_156# vdd 0.003786f
C8713 ctln[1] _411_/a_1000_472# 0.040782f
C8714 fanout49/a_36_160# _440_/a_2665_112# 0.00631f
C8715 _431_/a_36_151# FILLER_0_17_133/a_36_472# 0.001723f
C8716 FILLER_0_5_72/a_36_472# trim_mask\[1\] 0.015775f
C8717 FILLER_0_5_72/a_1380_472# _029_ 0.007385f
C8718 _086_ _267_/a_1792_472# 0.002715f
C8719 _261_/a_36_160# _163_ 0.002002f
C8720 net26 _423_/a_1204_472# 0.001069f
C8721 output29/a_224_472# net18 0.010345f
C8722 _413_/a_2560_156# net59 0.016463f
C8723 _412_/a_36_151# net18 0.011383f
C8724 _431_/a_2248_156# _136_ 0.030673f
C8725 output39/a_224_472# net17 0.041253f
C8726 net57 FILLER_0_16_154/a_1468_375# 0.217874f
C8727 FILLER_0_17_218/a_36_472# _069_ 0.001246f
C8728 _118_ _311_/a_66_473# 0.008528f
C8729 net51 _450_/a_2449_156# 0.008215f
C8730 FILLER_0_2_111/a_932_472# vss -0.001894f
C8731 FILLER_0_2_111/a_1380_472# vdd 0.002688f
C8732 cal_count\[3\] _453_/a_1000_472# 0.001123f
C8733 FILLER_0_21_286/a_36_472# net18 0.18097f
C8734 _053_ _220_/a_255_603# 0.001311f
C8735 _134_ vdd 0.482157f
C8736 _431_/a_36_151# net73 0.015086f
C8737 net48 vdd 0.35704f
C8738 trimb[1] FILLER_0_19_28/a_124_375# 0.00285f
C8739 _043_ FILLER_0_12_196/a_124_375# 0.003935f
C8740 _065_ trim_mask\[3\] 0.020092f
C8741 _187_ _408_/a_1336_472# 0.002191f
C8742 _103_ _418_/a_448_472# 0.002678f
C8743 _091_ _429_/a_448_472# 0.034713f
C8744 net60 _418_/a_1308_423# 0.016365f
C8745 _002_ vss 0.08396f
C8746 fanout62/a_36_160# vss 0.01343f
C8747 net20 _419_/a_1000_472# 0.022734f
C8748 net60 _419_/a_2665_112# 0.059916f
C8749 _136_ FILLER_0_15_180/a_36_472# 0.006924f
C8750 FILLER_0_5_88/a_36_472# _164_ 0.011718f
C8751 net31 output18/a_224_472# 0.04975f
C8752 output44/a_224_472# net44 0.051347f
C8753 FILLER_0_24_63/a_36_472# output25/a_224_472# 0.002338f
C8754 _146_ vdd 0.031209f
C8755 net32 result[8] 0.024881f
C8756 net58 FILLER_0_9_282/a_124_375# 0.021949f
C8757 FILLER_0_21_28/a_3172_472# _012_ 0.018785f
C8758 _390_/a_244_472# _067_ 0.004031f
C8759 trim_mask\[4\] FILLER_0_2_165/a_124_375# 0.011181f
C8760 _320_/a_1792_472# net79 0.002091f
C8761 FILLER_0_21_150/a_36_472# vss 0.012815f
C8762 _174_ _183_ 0.008231f
C8763 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_572_375# 0.086635f
C8764 _031_ _153_ 0.009316f
C8765 FILLER_0_23_60/a_124_375# vdd 0.031398f
C8766 FILLER_0_6_177/a_124_375# vdd 0.017329f
C8767 _053_ trim_mask\[0\] 0.007667f
C8768 FILLER_0_12_136/a_1380_472# net23 0.011488f
C8769 _394_/a_728_93# _043_ 0.00355f
C8770 ctlp[1] FILLER_0_23_290/a_124_375# 0.053745f
C8771 _027_ net36 0.185347f
C8772 _408_/a_56_524# _067_ 0.003678f
C8773 _070_ _055_ 0.516713f
C8774 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1380_472# 0.013276f
C8775 comp cal_count\[2\] 0.015029f
C8776 net55 FILLER_0_11_78/a_124_375# 0.001597f
C8777 _308_/a_1084_68# trim_mask\[0\] 0.001592f
C8778 _258_/a_36_160# _073_ 0.079254f
C8779 net53 net23 0.501857f
C8780 FILLER_0_15_142/a_484_472# net36 0.012033f
C8781 net16 net72 0.367221f
C8782 _176_ FILLER_0_15_72/a_484_472# 0.00753f
C8783 _152_ _058_ 0.00259f
C8784 net21 FILLER_0_12_196/a_124_375# 0.005374f
C8785 _444_/a_2665_112# FILLER_0_6_37/a_124_375# 0.005477f
C8786 FILLER_0_24_96/a_124_375# net24 0.040364f
C8787 _079_ net76 2.404004f
C8788 net66 FILLER_0_5_54/a_932_472# 0.001419f
C8789 _423_/a_36_151# FILLER_0_23_44/a_484_472# 0.001723f
C8790 net50 _220_/a_67_603# 0.005566f
C8791 _068_ _311_/a_66_473# 0.071325f
C8792 _394_/a_728_93# _175_ 0.010801f
C8793 _089_ _122_ 0.006163f
C8794 FILLER_0_15_116/a_36_472# net36 0.013546f
C8795 _427_/a_796_472# _095_ 0.007281f
C8796 _431_/a_2665_112# net53 0.004057f
C8797 _334_/a_36_160# FILLER_0_17_104/a_1380_472# 0.004111f
C8798 net73 _427_/a_448_472# 0.00132f
C8799 _070_ _313_/a_67_603# 0.004265f
C8800 net9 cal_itt\[0\] 0.110446f
C8801 _216_/a_67_603# FILLER_0_18_61/a_124_375# 0.014522f
C8802 FILLER_0_5_54/a_484_472# trim_mask\[1\] 0.013584f
C8803 FILLER_0_4_99/a_124_375# vdd 0.029154f
C8804 FILLER_0_0_266/a_124_375# rstn 0.073089f
C8805 FILLER_0_21_142/a_36_472# vss 0.009084f
C8806 FILLER_0_21_142/a_484_472# vdd 0.004917f
C8807 _260_/a_36_68# FILLER_0_3_221/a_1380_472# 0.001652f
C8808 _080_ FILLER_0_3_221/a_1020_375# 0.001414f
C8809 _091_ FILLER_0_15_180/a_484_472# 0.001757f
C8810 _058_ FILLER_0_10_94/a_36_472# 0.009346f
C8811 net79 FILLER_0_15_282/a_572_375# 0.01043f
C8812 net20 FILLER_0_15_212/a_1020_375# 0.001629f
C8813 net17 _452_/a_1293_527# 0.001011f
C8814 _374_/a_36_68# _076_ 0.026674f
C8815 net50 _036_ 0.002727f
C8816 FILLER_0_17_72/a_3172_472# vdd 0.002712f
C8817 FILLER_0_11_124/a_124_375# _120_ 0.012164f
C8818 net7 net41 0.243942f
C8819 trim_mask\[2\] FILLER_0_4_91/a_124_375# 0.003591f
C8820 _115_ _120_ 0.076035f
C8821 mask\[1\] FILLER_0_15_228/a_36_472# 0.02055f
C8822 FILLER_0_4_49/a_124_375# trim_val\[1\] 0.024557f
C8823 _069_ _176_ 0.766885f
C8824 output29/a_224_472# net62 0.138536f
C8825 net58 fanout76/a_36_160# 0.055026f
C8826 ctlp[1] net33 0.11288f
C8827 mask\[0\] _283_/a_36_472# 0.004645f
C8828 net16 _424_/a_36_151# 0.002969f
C8829 _440_/a_2665_112# FILLER_0_4_91/a_36_472# 0.007491f
C8830 vdd output6/a_224_472# 0.009312f
C8831 FILLER_0_12_136/a_572_375# _120_ 0.001584f
C8832 net43 net40 0.018193f
C8833 _257_/a_36_472# _075_ 0.005709f
C8834 _136_ _337_/a_665_69# 0.001794f
C8835 _006_ vss 0.111492f
C8836 net16 _447_/a_448_472# 0.063057f
C8837 FILLER_0_4_197/a_124_375# vdd 0.011327f
C8838 fanout59/a_36_160# net59 0.021522f
C8839 _015_ FILLER_0_8_247/a_484_472# 0.005458f
C8840 trim_mask\[4\] net59 0.012971f
C8841 FILLER_0_16_107/a_572_375# net14 0.002308f
C8842 net75 net8 0.553872f
C8843 _343_/a_49_472# mask\[4\] 0.036987f
C8844 _186_ _407_/a_244_68# 0.001153f
C8845 output35/a_224_472# _048_ 0.009509f
C8846 vss output40/a_224_472# 0.002459f
C8847 _441_/a_1308_423# vss 0.016854f
C8848 _066_ _386_/a_124_24# 0.059053f
C8849 _098_ _434_/a_2248_156# 0.016991f
C8850 _070_ _058_ 0.07307f
C8851 net53 _427_/a_2560_156# 0.004594f
C8852 _015_ _426_/a_1308_423# 0.029444f
C8853 FILLER_0_13_206/a_124_375# vdd 0.034528f
C8854 _447_/a_36_151# vdd 0.067176f
C8855 FILLER_0_4_123/a_36_472# FILLER_0_2_111/a_1468_375# 0.00189f
C8856 FILLER_0_18_2/a_2364_375# vdd 0.002983f
C8857 FILLER_0_15_228/a_36_472# vss 0.006585f
C8858 _070_ _315_/a_36_68# 0.031892f
C8859 output39/a_224_472# net39 0.129913f
C8860 _115_ FILLER_0_9_105/a_572_375# 0.003191f
C8861 _286_/a_224_472# _094_ 0.008468f
C8862 cal_itt\[3\] _072_ 2.019868f
C8863 output31/a_224_472# FILLER_0_17_282/a_36_472# 0.008834f
C8864 _431_/a_1308_423# vss 0.003472f
C8865 _440_/a_2248_156# vss 0.010006f
C8866 _440_/a_2665_112# vdd -0.002297f
C8867 FILLER_0_19_142/a_36_472# vss 0.011026f
C8868 _430_/a_1308_423# _069_ 0.024499f
C8869 _439_/a_448_472# vss 0.036535f
C8870 _439_/a_1308_423# vdd 0.002368f
C8871 net80 _434_/a_1000_472# 0.01421f
C8872 net80 _340_/a_36_160# 0.004225f
C8873 FILLER_0_20_87/a_36_472# _438_/a_1308_423# 0.010224f
C8874 _091_ FILLER_0_13_212/a_36_472# 0.007355f
C8875 _095_ net14 0.043065f
C8876 _412_/a_448_472# net58 0.044616f
C8877 _323_/a_36_113# vdd 0.009958f
C8878 fanout56/a_36_113# vdd 0.078814f
C8879 _430_/a_2665_112# FILLER_0_17_218/a_572_375# 0.002362f
C8880 trim_mask\[2\] FILLER_0_2_93/a_484_472# 0.001424f
C8881 _098_ _437_/a_1308_423# 0.005568f
C8882 net20 FILLER_0_3_221/a_932_472# 0.054476f
C8883 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_124_375# 0.016748f
C8884 _273_/a_36_68# FILLER_0_10_214/a_36_472# 0.003036f
C8885 _053_ _081_ 0.698311f
C8886 FILLER_0_7_104/a_1468_375# _131_ 0.029718f
C8887 FILLER_0_19_47/a_484_472# vss 0.001338f
C8888 _402_/a_1948_68# _401_/a_36_68# 0.012664f
C8889 FILLER_0_5_181/a_36_472# net37 0.010376f
C8890 net36 _438_/a_796_472# 0.016855f
C8891 output33/a_224_472# net34 0.077682f
C8892 trim[4] net67 0.06366f
C8893 _386_/a_124_24# net37 0.00431f
C8894 net27 FILLER_0_11_282/a_124_375# 0.002857f
C8895 output28/a_224_472# net19 0.101711f
C8896 _067_ _043_ 0.189767f
C8897 net63 _434_/a_2248_156# 0.063346f
C8898 trim[1] vdd 0.089624f
C8899 net15 _441_/a_36_151# 0.01821f
C8900 _053_ FILLER_0_7_104/a_932_472# 0.002529f
C8901 mask\[5\] FILLER_0_20_177/a_36_472# 0.017871f
C8902 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_124_375# 0.009654f
C8903 FILLER_0_16_57/a_1020_375# net72 0.002937f
C8904 _126_ _320_/a_36_472# 0.026216f
C8905 _077_ _251_/a_468_472# 0.002497f
C8906 _144_ _049_ 0.100508f
C8907 _093_ _304_/a_224_472# 0.002907f
C8908 en vdd 0.282941f
C8909 _077_ net68 0.003823f
C8910 net15 _440_/a_1000_472# 0.056791f
C8911 _079_ _083_ 0.872842f
C8912 _088_ _078_ 0.047558f
C8913 _412_/a_2560_156# net1 0.005618f
C8914 _115_ _227_/a_36_160# 0.00124f
C8915 cal_count\[3\] net17 0.068527f
C8916 _063_ FILLER_0_6_47/a_36_472# 0.007244f
C8917 _311_/a_66_473# vdd 0.106886f
C8918 _452_/a_448_472# net40 0.047031f
C8919 _207_/a_67_603# vss 0.00837f
C8920 _444_/a_2665_112# FILLER_0_8_37/a_484_472# 0.001167f
C8921 FILLER_0_7_146/a_124_375# _076_ 0.00688f
C8922 FILLER_0_7_146/a_36_472# _133_ 0.009796f
C8923 FILLER_0_22_86/a_932_472# net14 0.020589f
C8924 net81 _099_ 0.140011f
C8925 net36 FILLER_0_15_212/a_124_375# 0.004391f
C8926 _435_/a_448_472# vdd 0.029967f
C8927 _448_/a_2248_156# net59 0.005684f
C8928 _053_ _414_/a_2665_112# 0.032254f
C8929 _085_ _267_/a_36_472# 0.034055f
C8930 net31 _419_/a_2248_156# 0.001521f
C8931 net36 _196_/a_36_160# 0.024527f
C8932 _176_ FILLER_0_15_59/a_124_375# 0.007169f
C8933 _094_ _195_/a_67_603# 0.043278f
C8934 _408_/a_728_93# cal_count\[2\] 0.001568f
C8935 _427_/a_796_472# vss 0.001131f
C8936 _256_/a_3368_68# net22 0.001285f
C8937 _140_ _024_ 0.00287f
C8938 _221_/a_36_160# _054_ 0.02124f
C8939 FILLER_0_21_133/a_124_375# net54 0.013027f
C8940 FILLER_0_7_72/a_1380_472# vss 0.001117f
C8941 _062_ _163_ 0.001206f
C8942 ctln[3] _000_ 0.008418f
C8943 FILLER_0_9_28/a_1916_375# vdd 0.01295f
C8944 _405_/a_67_603# _184_ 0.010046f
C8945 FILLER_0_8_127/a_124_375# vdd 0.019587f
C8946 vdd FILLER_0_21_60/a_572_375# 0.022291f
C8947 vss FILLER_0_21_60/a_124_375# 0.003723f
C8948 _162_ calibrate 0.228839f
C8949 mask\[5\] FILLER_0_19_171/a_932_472# 0.007596f
C8950 _451_/a_36_151# _040_ 0.018648f
C8951 _002_ FILLER_0_3_172/a_3172_472# 0.002313f
C8952 valid net37 0.051518f
C8953 net22 _202_/a_36_160# 0.052766f
C8954 _427_/a_796_472# net74 0.020124f
C8955 net76 vss 0.436111f
C8956 net44 _450_/a_1040_527# 0.002267f
C8957 _105_ result[8] 0.011678f
C8958 _273_/a_36_68# _246_/a_36_68# 0.001168f
C8959 cal_itt\[0\] _084_ 0.061227f
C8960 FILLER_0_12_28/a_36_472# net40 0.020589f
C8961 FILLER_0_13_290/a_124_375# _416_/a_36_151# 0.026277f
C8962 FILLER_0_22_177/a_36_472# net33 0.013661f
C8963 net68 _453_/a_36_151# 0.039234f
C8964 ctlp[5] net22 0.001542f
C8965 _282_/a_36_160# _098_ 0.00388f
C8966 FILLER_0_13_212/a_124_375# vdd 0.010978f
C8967 net52 FILLER_0_2_127/a_36_472# 0.001964f
C8968 output15/a_224_472# net50 0.00515f
C8969 ctln[8] fanout50/a_36_160# 0.004838f
C8970 net69 net49 0.051235f
C8971 FILLER_0_19_155/a_484_472# vss 0.004002f
C8972 net16 _407_/a_36_472# 0.027354f
C8973 output32/a_224_472# _094_ 0.005545f
C8974 FILLER_0_17_72/a_572_375# _131_ 0.006224f
C8975 _442_/a_1000_472# _031_ 0.004174f
C8976 FILLER_0_16_255/a_36_472# _102_ 0.004641f
C8977 _016_ FILLER_0_12_136/a_572_375# 0.00332f
C8978 net68 net69 0.053856f
C8979 FILLER_0_3_142/a_36_472# trim_mask\[4\] 0.008297f
C8980 FILLER_0_5_72/a_1020_375# net47 0.006974f
C8981 net14 FILLER_0_4_91/a_484_472# 0.020589f
C8982 net19 calibrate 0.043159f
C8983 ctlp[2] _109_ 0.059999f
C8984 net46 net43 0.215092f
C8985 _429_/a_2665_112# FILLER_0_15_212/a_1468_375# 0.010688f
C8986 FILLER_0_17_200/a_484_472# vss 0.003134f
C8987 _173_ vss 0.063821f
C8988 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_124_375# 0.003228f
C8989 fanout61/a_36_113# FILLER_0_21_286/a_572_375# 0.015816f
C8990 _161_ _056_ 0.065732f
C8991 _127_ net23 0.069001f
C8992 FILLER_0_9_223/a_36_472# _273_/a_36_68# 0.015795f
C8993 _039_ net6 0.104745f
C8994 FILLER_0_10_214/a_36_472# _246_/a_36_68# 0.001844f
C8995 _274_/a_36_68# FILLER_0_12_220/a_484_472# 0.001048f
C8996 FILLER_0_16_107/a_484_472# _040_ 0.003828f
C8997 mask\[8\] net14 0.040566f
C8998 net38 net55 0.10956f
C8999 _057_ _311_/a_66_473# 0.042545f
C9000 output46/a_224_472# vss 0.00432f
C9001 FILLER_0_20_193/a_572_375# net21 0.002103f
C9002 _132_ _017_ 0.155924f
C9003 FILLER_0_7_59/a_36_472# vdd 0.016778f
C9004 FILLER_0_7_59/a_572_375# vss 0.017487f
C9005 _147_ _146_ 0.001164f
C9006 net16 _444_/a_1308_423# 0.002172f
C9007 net70 _131_ 0.57653f
C9008 _405_/a_67_603# net47 0.004116f
C9009 net35 FILLER_0_22_128/a_2812_375# 0.010399f
C9010 _137_ _333_/a_36_160# 0.022811f
C9011 _007_ vss 0.017377f
C9012 FILLER_0_1_204/a_36_472# vdd 0.009339f
C9013 FILLER_0_1_204/a_124_375# vss 0.018397f
C9014 net2 en 0.067828f
C9015 _114_ FILLER_0_12_136/a_36_472# 0.003953f
C9016 _009_ FILLER_0_23_290/a_36_472# 0.002345f
C9017 mask\[5\] _204_/a_67_603# 0.023791f
C9018 net68 FILLER_0_6_47/a_572_375# 0.007672f
C9019 _256_/a_3368_68# _076_ 0.001183f
C9020 FILLER_0_12_20/a_124_375# net17 0.002167f
C9021 vss net14 1.003274f
C9022 _013_ _424_/a_448_472# 0.043803f
C9023 net58 _425_/a_2665_112# 0.069807f
C9024 FILLER_0_9_72/a_572_375# _439_/a_36_151# 0.059049f
C9025 _103_ _006_ 0.00205f
C9026 trim_mask\[1\] FILLER_0_6_47/a_1468_375# 0.007169f
C9027 output19/a_224_472# _422_/a_2248_156# 0.011418f
C9028 ctlp[2] _422_/a_448_472# 0.011383f
C9029 output31/a_224_472# _289_/a_36_472# 0.00101f
C9030 output15/a_224_472# trim_mask\[3\] 0.024718f
C9031 net63 FILLER_0_22_177/a_572_375# 0.001597f
C9032 _071_ net23 0.027895f
C9033 _080_ vdd 0.123811f
C9034 net72 FILLER_0_17_64/a_124_375# 0.002236f
C9035 FILLER_0_22_128/a_36_472# vdd 0.004601f
C9036 FILLER_0_22_128/a_3260_375# vss 0.006346f
C9037 _297_/a_36_472# _295_/a_36_472# 0.004259f
C9038 FILLER_0_7_72/a_2812_375# net14 0.025092f
C9039 _444_/a_36_151# vss 0.003795f
C9040 _444_/a_448_472# vdd 0.03285f
C9041 FILLER_0_21_28/a_1468_375# _423_/a_36_151# 0.001543f
C9042 _415_/a_2560_156# net18 0.010318f
C9043 net74 net14 0.034568f
C9044 trim_mask\[2\] _367_/a_36_68# 0.001302f
C9045 fanout75/a_36_113# _081_ 0.015843f
C9046 _187_ _450_/a_3129_107# 0.00126f
C9047 fanout62/a_36_160# FILLER_0_9_290/a_36_472# 0.001961f
C9048 _155_ _151_ 0.10611f
C9049 FILLER_0_19_47/a_124_375# _182_ 0.001771f
C9050 _052_ net36 0.005689f
C9051 _005_ net18 0.073455f
C9052 net16 _404_/a_36_472# 0.001126f
C9053 net65 _413_/a_796_472# 0.006888f
C9054 trim[0] net40 0.005988f
C9055 net27 FILLER_0_9_270/a_36_472# 0.041681f
C9056 FILLER_0_10_78/a_572_375# vss 0.004588f
C9057 FILLER_0_10_78/a_1020_375# vdd 0.002901f
C9058 _176_ FILLER_0_11_101/a_484_472# 0.001777f
C9059 _154_ _157_ 0.447829f
C9060 _236_/a_36_160# net67 0.009332f
C9061 _428_/a_1204_472# _017_ 0.005148f
C9062 _085_ _113_ 0.084246f
C9063 _104_ _420_/a_2248_156# 0.027923f
C9064 FILLER_0_21_28/a_3260_375# _424_/a_36_151# 0.035849f
C9065 _413_/a_36_151# net21 0.012223f
C9066 FILLER_0_16_107/a_36_472# net36 0.001245f
C9067 FILLER_0_16_57/a_1380_472# net15 0.017841f
C9068 FILLER_0_18_2/a_484_472# net38 0.003391f
C9069 FILLER_0_8_2/a_124_375# net40 0.002839f
C9070 net63 FILLER_0_18_177/a_1916_375# 0.040551f
C9071 FILLER_0_5_54/a_1468_375# net47 0.005049f
C9072 _255_/a_224_552# _058_ 0.06267f
C9073 _132_ FILLER_0_12_124/a_36_472# 0.00101f
C9074 FILLER_0_9_72/a_484_472# vss 0.008087f
C9075 FILLER_0_9_72/a_932_472# vdd 0.00604f
C9076 _277_/a_36_160# net20 0.015569f
C9077 _028_ vdd 0.626868f
C9078 net82 FILLER_0_3_172/a_3260_375# 0.007693f
C9079 net68 _165_ 0.002748f
C9080 _066_ net59 0.002935f
C9081 _414_/a_448_472# net21 0.040301f
C9082 _328_/a_36_113# vdd 0.136098f
C9083 net55 FILLER_0_13_72/a_484_472# 0.004375f
C9084 FILLER_0_16_107/a_124_375# FILLER_0_16_89/a_1468_375# 0.005439f
C9085 net61 mask\[7\] 0.071542f
C9086 _093_ FILLER_0_17_72/a_3172_472# 0.012002f
C9087 _083_ vss 0.0284f
C9088 _094_ _418_/a_36_151# 0.041823f
C9089 ctlp[1] net18 0.088706f
C9090 _028_ FILLER_0_7_72/a_2364_375# 0.003884f
C9091 _137_ FILLER_0_16_154/a_36_472# 0.005011f
C9092 FILLER_0_5_164/a_572_375# net22 0.002238f
C9093 net64 FILLER_0_11_282/a_36_472# 0.003938f
C9094 _376_/a_36_160# FILLER_0_5_88/a_36_472# 0.001448f
C9095 _414_/a_2248_156# _075_ 0.044302f
C9096 _253_/a_36_68# _074_ 0.026327f
C9097 FILLER_0_6_90/a_484_472# FILLER_0_4_91/a_572_375# 0.00108f
C9098 net18 _417_/a_2248_156# 0.001601f
C9099 _126_ FILLER_0_13_100/a_124_375# 0.00134f
C9100 mask\[9\] FILLER_0_20_87/a_124_375# 0.004793f
C9101 fanout82/a_36_113# vdd 0.083174f
C9102 FILLER_0_16_89/a_932_472# _136_ 0.045229f
C9103 FILLER_0_15_282/a_484_472# output30/a_224_472# 0.001711f
C9104 FILLER_0_15_282/a_124_375# net30 0.00123f
C9105 _122_ FILLER_0_5_181/a_36_472# 0.003016f
C9106 _132_ FILLER_0_11_109/a_124_375# 0.008627f
C9107 _359_/a_1044_488# net74 0.005311f
C9108 _308_/a_848_380# vdd 0.013895f
C9109 FILLER_0_9_223/a_36_472# _246_/a_36_68# 0.006596f
C9110 output9/a_224_472# net19 0.070689f
C9111 FILLER_0_12_136/a_932_472# _069_ 0.002161f
C9112 FILLER_0_12_136/a_36_472# _126_ 0.014981f
C9113 _098_ FILLER_0_15_212/a_932_472# 0.011837f
C9114 _136_ _172_ 0.024344f
C9115 _053_ FILLER_0_7_72/a_572_375# 0.014569f
C9116 _130_ FILLER_0_12_136/a_36_472# 0.082451f
C9117 mask\[9\] net36 1.116767f
C9118 FILLER_0_20_15/a_124_375# vdd 0.006513f
C9119 FILLER_0_10_256/a_124_375# _015_ 0.001151f
C9120 _141_ vdd 0.439746f
C9121 net38 FILLER_0_15_10/a_36_472# 0.020589f
C9122 _316_/a_1084_68# net37 0.001574f
C9123 net37 net59 0.03883f
C9124 FILLER_0_17_72/a_932_472# net36 0.00356f
C9125 _132_ FILLER_0_14_107/a_1468_375# 0.019517f
C9126 _182_ _180_ 0.090106f
C9127 _129_ _059_ 0.005414f
C9128 net4 net37 0.021795f
C9129 FILLER_0_5_136/a_36_472# vdd 0.092379f
C9130 FILLER_0_5_136/a_124_375# vss 0.053395f
C9131 _105_ _098_ 0.055065f
C9132 _095_ FILLER_0_14_123/a_36_472# 0.014431f
C9133 mask\[7\] _108_ 0.785154f
C9134 _070_ _172_ 0.237178f
C9135 _190_/a_36_160# net47 0.001489f
C9136 FILLER_0_21_28/a_2724_472# vss -0.001553f
C9137 FILLER_0_6_90/a_36_472# vdd 0.00366f
C9138 FILLER_0_6_90/a_572_375# vss 0.006421f
C9139 output32/a_224_472# output34/a_224_472# 0.001691f
C9140 _428_/a_36_151# vdd 0.131612f
C9141 _119_ _319_/a_672_472# 0.00488f
C9142 mask\[4\] FILLER_0_19_171/a_484_472# 0.004669f
C9143 _142_ _334_/a_36_160# 0.009001f
C9144 FILLER_0_18_107/a_124_375# _438_/a_2665_112# 0.029834f
C9145 _430_/a_1308_423# net22 0.035518f
C9146 net63 FILLER_0_15_212/a_932_472# 0.002269f
C9147 FILLER_0_11_282/a_36_472# vss 0.007114f
C9148 _320_/a_224_472# _113_ 0.00871f
C9149 _176_ _038_ 0.039948f
C9150 _053_ _161_ 0.001047f
C9151 _051_ _098_ 0.006332f
C9152 net50 FILLER_0_9_60/a_36_472# 0.001914f
C9153 FILLER_0_18_2/a_3172_472# net17 0.002402f
C9154 FILLER_0_13_142/a_1380_472# _225_/a_36_160# 0.004111f
C9155 FILLER_0_4_107/a_484_472# _157_ 0.027364f
C9156 _115_ FILLER_0_10_107/a_484_472# 0.017642f
C9157 mask\[5\] _201_/a_67_603# 0.001222f
C9158 _163_ FILLER_0_5_148/a_36_472# 0.002454f
C9159 FILLER_0_8_263/a_124_375# net64 0.004793f
C9160 _445_/a_448_472# net17 0.038794f
C9161 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_36_472# 0.086742f
C9162 cal vdd 0.318671f
C9163 FILLER_0_15_116/a_572_375# net70 0.050592f
C9164 fanout50/a_36_160# vdd 0.009536f
C9165 trim_mask\[0\] FILLER_0_10_94/a_484_472# 0.015575f
C9166 _181_ _402_/a_2172_497# 0.001555f
C9167 net57 _385_/a_244_472# 0.001506f
C9168 _005_ net62 0.097739f
C9169 output48/a_224_472# _425_/a_36_151# 0.004037f
C9170 _443_/a_36_151# vdd 0.175472f
C9171 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_36_472# 0.002296f
C9172 net1 _001_ 0.300335f
C9173 ctlp[4] net32 0.001413f
C9174 _432_/a_36_151# _091_ 0.054497f
C9175 trim_val\[4\] FILLER_0_3_172/a_932_472# 0.001407f
C9176 FILLER_0_10_37/a_36_472# _453_/a_36_151# 0.003462f
C9177 _065_ net16 0.068602f
C9178 FILLER_0_7_72/a_124_375# net50 0.009304f
C9179 FILLER_0_7_72/a_1020_375# net52 0.00799f
C9180 vss _433_/a_2248_156# 0.034403f
C9181 vdd _433_/a_2665_112# 0.002569f
C9182 _414_/a_2665_112# _072_ 0.025361f
C9183 _176_ _076_ 0.046873f
C9184 _070_ FILLER_0_5_164/a_484_472# 0.003424f
C9185 FILLER_0_7_162/a_36_472# net37 0.090785f
C9186 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_124_375# 0.012552f
C9187 net52 FILLER_0_2_93/a_36_472# 0.009026f
C9188 net50 FILLER_0_2_93/a_124_375# 0.007132f
C9189 _096_ _098_ 0.00638f
C9190 _088_ FILLER_0_3_212/a_124_375# 0.0042f
C9191 _159_ _370_/a_124_24# 0.021983f
C9192 net79 FILLER_0_13_290/a_124_375# 0.043673f
C9193 output48/a_224_472# net1 0.006536f
C9194 _026_ net14 0.010792f
C9195 _147_ _435_/a_448_472# 0.001008f
C9196 ctlp[2] _300_/a_224_472# 0.002954f
C9197 _188_ net51 0.044278f
C9198 result[5] _008_ 0.165753f
C9199 _083_ _260_/a_244_472# 0.00134f
C9200 _251_/a_906_472# _068_ 0.001762f
C9201 output36/a_224_472# result[2] 0.002356f
C9202 _091_ net62 0.019946f
C9203 FILLER_0_2_177/a_124_375# vdd 0.019296f
C9204 net6 clkc 0.036083f
C9205 _114_ state\[1\] 0.087216f
C9206 _103_ _007_ 0.002514f
C9207 _417_/a_2248_156# net62 0.005537f
C9208 _058_ FILLER_0_8_156/a_36_472# 0.011885f
C9209 _310_/a_49_472# _113_ 0.020387f
C9210 _292_/a_36_160# _048_ 0.008475f
C9211 FILLER_0_17_218/a_572_375# vdd 0.019414f
C9212 FILLER_0_17_218/a_124_375# vss 0.012673f
C9213 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001597f
C9214 net71 FILLER_0_22_107/a_124_375# 0.018295f
C9215 net35 net25 0.129685f
C9216 trimb[3] net38 0.002836f
C9217 FILLER_0_8_263/a_36_472# vdd 0.092694f
C9218 FILLER_0_8_263/a_124_375# vss 0.007944f
C9219 fanout82/a_36_113# net2 0.008681f
C9220 net81 _082_ 0.001633f
C9221 _426_/a_2248_156# FILLER_0_8_239/a_124_375# 0.001068f
C9222 FILLER_0_24_63/a_124_375# vdd 0.029514f
C9223 mask\[5\] FILLER_0_19_187/a_36_472# 0.007596f
C9224 FILLER_0_20_31/a_36_472# vdd 0.097195f
C9225 FILLER_0_20_31/a_124_375# vss 0.049142f
C9226 net31 _006_ 0.307613f
C9227 _383_/a_36_472# vdd -0.002154f
C9228 FILLER_0_17_142/a_36_472# FILLER_0_19_142/a_124_375# 0.001512f
C9229 _414_/a_1308_423# _074_ 0.005458f
C9230 net20 _102_ 0.081029f
C9231 FILLER_0_21_286/a_124_375# vdd 0.026138f
C9232 _093_ FILLER_0_21_60/a_572_375# 0.011177f
C9233 _424_/a_36_151# _423_/a_1308_423# 0.001722f
C9234 FILLER_0_4_144/a_124_375# net47 0.012023f
C9235 _135_ _134_ 0.038135f
C9236 FILLER_0_20_87/a_36_472# vss 0.006244f
C9237 FILLER_0_5_198/a_124_375# net37 0.009149f
C9238 output27/a_224_472# fanout64/a_36_160# 0.027335f
C9239 FILLER_0_10_78/a_124_375# cal_count\[3\] 0.012197f
C9240 _408_/a_728_93# _402_/a_56_567# 0.001359f
C9241 _322_/a_1084_68# _129_ 0.00419f
C9242 _091_ FILLER_0_19_171/a_572_375# 0.013568f
C9243 FILLER_0_9_223/a_484_472# _055_ 0.026026f
C9244 _440_/a_1308_423# _160_ 0.002554f
C9245 _028_ FILLER_0_6_47/a_3172_472# 0.015585f
C9246 net81 _426_/a_448_472# 0.003907f
C9247 output42/a_224_472# _039_ 0.001254f
C9248 _394_/a_718_524# vss 0.002666f
C9249 _211_/a_36_160# net14 0.005761f
C9250 _429_/a_2665_112# FILLER_0_15_228/a_124_375# 0.001077f
C9251 FILLER_0_9_223/a_572_375# calibrate 0.002082f
C9252 _132_ FILLER_0_16_115/a_124_375# 0.033245f
C9253 _413_/a_36_151# FILLER_0_3_172/a_1468_375# 0.001252f
C9254 FILLER_0_2_93/a_124_375# trim_mask\[3\] 0.003033f
C9255 net38 _444_/a_1204_472# 0.018432f
C9256 net61 net79 0.159f
C9257 _056_ _246_/a_36_68# 0.017953f
C9258 FILLER_0_19_28/a_484_472# vss 0.001207f
C9259 FILLER_0_3_204/a_36_472# net59 0.001606f
C9260 FILLER_0_6_239/a_124_375# _317_/a_36_113# 0.002437f
C9261 _448_/a_36_151# _037_ 0.012725f
C9262 output35/a_224_472# _435_/a_2665_112# 0.008469f
C9263 _091_ _072_ 0.162027f
C9264 _269_/a_36_472# _083_ 0.015096f
C9265 _115_ _322_/a_692_472# 0.00171f
C9266 _077_ FILLER_0_9_60/a_124_375# 0.051389f
C9267 _412_/a_2248_156# output37/a_224_472# 0.001141f
C9268 _323_/a_36_113# FILLER_0_10_247/a_124_375# 0.001846f
C9269 _053_ FILLER_0_6_47/a_1380_472# 0.004472f
C9270 _259_/a_455_68# net37 0.0023f
C9271 _436_/a_1204_472# net35 0.005186f
C9272 _441_/a_36_151# net66 0.057618f
C9273 fanout74/a_36_113# net23 0.005294f
C9274 result[7] _419_/a_36_151# 0.001036f
C9275 FILLER_0_16_89/a_1468_375# vdd 0.038266f
C9276 net64 FILLER_0_9_270/a_484_472# 0.017924f
C9277 _417_/a_2665_112# net30 0.015638f
C9278 net41 _452_/a_36_151# 0.036301f
C9279 _002_ FILLER_0_4_185/a_36_472# 0.004231f
C9280 ctlp[5] _140_ 0.002123f
C9281 mask\[2\] FILLER_0_15_235/a_484_472# 0.004683f
C9282 trim[0] trim[3] 0.012429f
C9283 _121_ _062_ 0.001616f
C9284 _430_/a_1204_472# _091_ 0.007301f
C9285 _412_/a_2248_156# net5 0.048919f
C9286 _395_/a_36_488# _055_ 0.002775f
C9287 net76 FILLER_0_5_206/a_36_472# 0.00169f
C9288 _176_ FILLER_0_11_78/a_484_472# 0.008724f
C9289 FILLER_0_21_142/a_124_375# net54 0.027551f
C9290 cal net2 0.081236f
C9291 output9/a_224_472# cal_itt\[0\] 0.008307f
C9292 net49 _440_/a_448_472# 0.049861f
C9293 result[9] ctlp[2] 0.105977f
C9294 FILLER_0_15_116/a_124_375# FILLER_0_14_107/a_1020_375# 0.026339f
C9295 FILLER_0_7_146/a_36_472# net37 0.00208f
C9296 ctln[1] FILLER_0_3_221/a_572_375# 0.001554f
C9297 output8/a_224_472# FILLER_0_3_221/a_932_472# 0.001699f
C9298 _394_/a_718_524# cal_count\[1\] 0.009499f
C9299 _394_/a_56_524# net15 0.006099f
C9300 output10/a_224_472# vss 0.014205f
C9301 net65 _448_/a_448_472# 0.001006f
C9302 net68 _440_/a_448_472# 0.02254f
C9303 net32 _419_/a_448_472# 0.011757f
C9304 _436_/a_2248_156# vss 0.002799f
C9305 _436_/a_2665_112# vdd 0.007946f
C9306 net20 _198_/a_67_603# 0.013603f
C9307 _415_/a_1000_472# net27 0.017938f
C9308 FILLER_0_4_197/a_932_472# net59 0.003599f
C9309 FILLER_0_22_128/a_36_472# _433_/a_36_151# 0.001653f
C9310 ctlp[1] _420_/a_1000_472# 0.001106f
C9311 vdd _034_ 0.424437f
C9312 FILLER_0_17_200/a_36_472# mask\[4\] 0.001242f
C9313 _430_/a_2665_112# mask\[2\] 0.028551f
C9314 _126_ state\[1\] 1.191746f
C9315 _178_ _186_ 0.020123f
C9316 _174_ _401_/a_36_68# 0.033989f
C9317 net29 net19 0.305661f
C9318 output7/a_224_472# vdd 0.086699f
C9319 net72 FILLER_0_17_56/a_36_472# 0.008058f
C9320 _138_ _043_ 0.005826f
C9321 _020_ _142_ 0.010094f
C9322 _139_ _337_/a_49_472# 0.024331f
C9323 net41 FILLER_0_12_28/a_124_375# 0.003909f
C9324 _085_ vdd 0.227153f
C9325 _414_/a_2248_156# net22 0.062122f
C9326 FILLER_0_5_164/a_124_375# vdd 0.00419f
C9327 FILLER_0_19_55/a_124_375# FILLER_0_19_47/a_572_375# 0.012001f
C9328 net16 _036_ 0.637538f
C9329 net20 mask\[3\] 0.047107f
C9330 net39 _445_/a_448_472# 0.014537f
C9331 _372_/a_170_472# _385_/a_36_68# 0.009691f
C9332 FILLER_0_1_266/a_484_472# net8 0.016327f
C9333 _008_ net19 0.027093f
C9334 _008_ _418_/a_1204_472# 0.002933f
C9335 net16 _445_/a_2665_112# 0.061595f
C9336 _326_/a_36_160# _322_/a_124_24# 0.004397f
C9337 FILLER_0_11_101/a_572_375# _070_ 0.011557f
C9338 ctln[6] output14/a_224_472# 0.007421f
C9339 ctlp[7] net25 0.003141f
C9340 net38 FILLER_0_20_15/a_36_472# 0.070475f
C9341 _018_ vdd 0.048119f
C9342 FILLER_0_12_220/a_1468_375# _060_ 0.001429f
C9343 FILLER_0_12_220/a_484_472# _090_ 0.006993f
C9344 input5/a_36_113# net5 0.061819f
C9345 _163_ _153_ 0.243815f
C9346 ctlp[1] _421_/a_2248_156# 0.012937f
C9347 net49 vss 0.689397f
C9348 _427_/a_2560_156# net23 0.042069f
C9349 _251_/a_468_472# vss 0.001679f
C9350 calibrate _055_ 0.006584f
C9351 state\[2\] FILLER_0_13_142/a_572_375# 0.007511f
C9352 fanout53/a_36_160# net53 0.014917f
C9353 net53 FILLER_0_13_142/a_1468_375# 0.002334f
C9354 _442_/a_2665_112# vdd 0.056153f
C9355 _425_/a_36_151# _316_/a_124_24# 0.036238f
C9356 result[7] _420_/a_2248_156# 0.034866f
C9357 _446_/a_2248_156# net17 0.008375f
C9358 net68 vss 0.635359f
C9359 _122_ net59 0.041453f
C9360 _076_ FILLER_0_8_239/a_36_472# 0.029514f
C9361 net15 _423_/a_2665_112# 0.061217f
C9362 _144_ FILLER_0_19_125/a_124_375# 0.012834f
C9363 FILLER_0_16_57/a_1380_472# _394_/a_728_93# 0.001627f
C9364 _445_/a_2248_156# vdd 0.018573f
C9365 net20 _256_/a_36_68# 0.02797f
C9366 _114_ _096_ 0.066848f
C9367 FILLER_0_5_117/a_124_375# _153_ 0.079379f
C9368 _424_/a_2665_112# FILLER_0_21_60/a_572_375# 0.001077f
C9369 _070_ _152_ 0.114651f
C9370 _133_ _081_ 0.002847f
C9371 net4 _122_ 0.03487f
C9372 trim_val\[4\] net23 0.014503f
C9373 _048_ FILLER_0_18_209/a_124_375# 0.001615f
C9374 vdd output30/a_224_472# 0.068123f
C9375 _138_ net21 0.003242f
C9376 net75 vdd 1.265616f
C9377 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_36_472# 0.086742f
C9378 net32 _420_/a_2665_112# 0.002753f
C9379 net73 FILLER_0_18_107/a_1468_375# 0.024898f
C9380 FILLER_0_7_104/a_932_472# _133_ 0.019721f
C9381 _346_/a_49_472# _145_ 0.001141f
C9382 _372_/a_3662_472# _062_ 0.0012f
C9383 _408_/a_56_524# net17 0.048018f
C9384 FILLER_0_18_177/a_572_375# FILLER_0_20_177/a_484_472# 0.0027f
C9385 mask\[7\] _049_ 0.234746f
C9386 _430_/a_448_472# vdd 0.002959f
C9387 _430_/a_36_151# vss 0.011779f
C9388 _077_ _453_/a_2665_112# 0.002824f
C9389 _425_/a_1000_472# vdd 0.019072f
C9390 vss FILLER_0_3_212/a_36_472# 0.00838f
C9391 net57 fanout56/a_36_113# 0.079542f
C9392 calibrate _313_/a_67_603# 0.021436f
C9393 net41 _039_ 0.030362f
C9394 mask\[7\] _435_/a_2665_112# 0.030393f
C9395 net1 input4/a_36_68# 0.056389f
C9396 _285_/a_36_472# net62 0.001288f
C9397 _104_ vdd 0.662413f
C9398 net65 FILLER_0_1_266/a_36_472# 0.003529f
C9399 FILLER_0_5_117/a_36_472# _163_ 0.007418f
C9400 _070_ FILLER_0_10_94/a_36_472# 0.001866f
C9401 FILLER_0_8_24/a_124_375# net17 0.039695f
C9402 ctlp[4] _105_ 0.002221f
C9403 net15 trim_mask\[1\] 0.042093f
C9404 _443_/a_2248_156# _386_/a_124_24# 0.001257f
C9405 net34 _422_/a_1204_472# 0.001029f
C9406 _420_/a_36_151# vdd 0.137919f
C9407 _185_ _402_/a_728_93# 0.007151f
C9408 fanout65/a_36_113# vdd 0.10473f
C9409 net63 _024_ 0.001348f
C9410 net16 _183_ 0.001103f
C9411 _041_ net40 0.082688f
C9412 _333_/a_36_160# vss 0.030799f
C9413 _320_/a_224_472# vdd 0.001757f
C9414 fanout66/a_36_113# net69 0.001345f
C9415 _436_/a_2665_112# FILLER_0_22_128/a_572_375# 0.001092f
C9416 _436_/a_2560_156# FILLER_0_22_128/a_124_375# 0.001178f
C9417 _208_/a_36_160# vss 0.012188f
C9418 _098_ FILLER_0_15_180/a_124_375# 0.019007f
C9419 net58 sample 0.006906f
C9420 _415_/a_1308_423# _004_ 0.002098f
C9421 _057_ _085_ 0.543871f
C9422 _026_ FILLER_0_20_87/a_36_472# 0.004568f
C9423 _199_/a_36_160# _046_ 0.017122f
C9424 _141_ _093_ 0.396041f
C9425 _072_ _161_ 0.048567f
C9426 result[4] net77 0.003336f
C9427 FILLER_0_18_2/a_3260_375# _041_ 0.001024f
C9428 net76 _123_ 0.003431f
C9429 net57 _311_/a_66_473# 0.013777f
C9430 net16 FILLER_0_6_37/a_36_472# 0.013074f
C9431 FILLER_0_21_125/a_124_375# vdd -0.010326f
C9432 _089_ _087_ 0.002217f
C9433 _136_ _070_ 0.010577f
C9434 _449_/a_448_472# _038_ 0.064169f
C9435 _058_ _439_/a_2665_112# 0.001029f
C9436 FILLER_0_16_57/a_1020_375# _176_ 0.006334f
C9437 _095_ _184_ 0.265966f
C9438 _136_ _356_/a_36_472# 0.004667f
C9439 _267_/a_224_472# state\[1\] 0.001937f
C9440 FILLER_0_18_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001684f
C9441 _434_/a_36_151# _146_ 0.003818f
C9442 _434_/a_1204_472# mask\[6\] 0.006692f
C9443 mask\[4\] FILLER_0_19_187/a_572_375# 0.00553f
C9444 result[9] _421_/a_1000_472# 0.012144f
C9445 FILLER_0_17_72/a_2364_375# _136_ 0.047331f
C9446 net79 _416_/a_1000_472# 0.024811f
C9447 FILLER_0_8_247/a_1468_375# vdd 0.011086f
C9448 result[5] fanout61/a_36_113# 0.001866f
C9449 _421_/a_448_472# vss -0.001027f
C9450 _421_/a_1308_423# vdd 0.021664f
C9451 trim_mask\[4\] _081_ 0.111668f
C9452 vdd FILLER_0_6_37/a_124_375# 0.041381f
C9453 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1380_472# 0.013276f
C9454 _058_ calibrate 0.075294f
C9455 net23 FILLER_0_22_128/a_1828_472# 0.003857f
C9456 output43/a_224_472# vss -0.005182f
C9457 _170_ _386_/a_124_24# 0.008511f
C9458 FILLER_0_21_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001723f
C9459 net72 _131_ 0.186396f
C9460 FILLER_0_10_214/a_124_375# _069_ 0.014379f
C9461 _096_ _126_ 0.258912f
C9462 cal_itt\[3\] net37 0.03677f
C9463 FILLER_0_5_117/a_124_375# FILLER_0_4_107/a_1380_472# 0.001684f
C9464 _426_/a_36_151# vdd 0.086652f
C9465 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_484_472# 0.013277f
C9466 FILLER_0_16_107/a_572_375# net70 0.002193f
C9467 cal_itt\[1\] net8 0.040042f
C9468 net58 net9 0.018829f
C9469 _029_ net14 0.042032f
C9470 output21/a_224_472# _108_ 0.005356f
C9471 ctln[7] trim_mask\[3\] 0.059414f
C9472 _095_ FILLER_0_13_100/a_124_375# 0.001989f
C9473 net82 FILLER_0_3_142/a_124_375# 0.018696f
C9474 _446_/a_1308_423# net40 0.038281f
C9475 output42/a_224_472# clkc 0.004924f
C9476 trim[4] output6/a_224_472# 0.004337f
C9477 _086_ _160_ 0.007038f
C9478 FILLER_0_5_172/a_124_375# FILLER_0_5_164/a_572_375# 0.012001f
C9479 _074_ _375_/a_1612_497# 0.004567f
C9480 net80 _435_/a_36_151# 0.035259f
C9481 _310_/a_49_472# vdd 0.043164f
C9482 _281_/a_672_472# _098_ 0.002084f
C9483 _122_ FILLER_0_5_198/a_124_375# 0.001352f
C9484 _187_ _042_ 0.009526f
C9485 _128_ _176_ 0.180252f
C9486 _210_/a_67_603# vss 0.038142f
C9487 _287_/a_36_472# net30 0.005402f
C9488 _086_ _116_ 1.316798f
C9489 net34 mask\[6\] 0.231853f
C9490 net65 FILLER_0_3_172/a_3260_375# 0.002696f
C9491 trimb[1] net17 0.084269f
C9492 net66 output41/a_224_472# 0.015427f
C9493 net63 _435_/a_1308_423# 0.003621f
C9494 FILLER_0_16_154/a_484_472# vdd 0.001006f
C9495 FILLER_0_16_154/a_36_472# vss 0.005098f
C9496 net70 _095_ 0.222423f
C9497 _412_/a_1000_472# cal_itt\[1\] 0.012926f
C9498 FILLER_0_5_72/a_1468_375# _440_/a_2665_112# 0.001077f
C9499 FILLER_0_8_239/a_124_375# vdd 0.035205f
C9500 _098_ _145_ 0.007514f
C9501 cal_itt\[2\] net8 0.057335f
C9502 net19 _420_/a_1204_472# 0.001828f
C9503 _095_ net47 0.508892f
C9504 _116_ cal_count\[3\] 0.384121f
C9505 mask\[7\] FILLER_0_22_128/a_2724_472# 0.001055f
C9506 net61 ctlp[2] 0.022612f
C9507 _154_ _160_ 0.395185f
C9508 net44 FILLER_0_8_2/a_36_472# 0.005851f
C9509 _144_ FILLER_0_18_107/a_1828_472# 0.001169f
C9510 output39/a_224_472# net67 0.008957f
C9511 FILLER_0_4_185/a_36_472# net76 0.023698f
C9512 _093_ FILLER_0_17_218/a_572_375# 0.0029f
C9513 fanout81/a_36_160# vdd 0.095319f
C9514 FILLER_0_21_125/a_572_375# _140_ 0.01659f
C9515 FILLER_0_7_104/a_36_472# vdd 0.096343f
C9516 FILLER_0_7_104/a_1468_375# vss 0.003442f
C9517 _053_ net23 0.031487f
C9518 _436_/a_796_472# _050_ 0.007055f
C9519 net74 _370_/a_1084_68# 0.001301f
C9520 FILLER_0_5_164/a_36_472# _066_ 0.00611f
C9521 net17 _043_ 0.571818f
C9522 FILLER_0_18_107/a_2812_375# vdd 0.004212f
C9523 _413_/a_1000_472# vdd 0.002781f
C9524 _365_/a_36_68# _156_ 0.027744f
C9525 result[1] FILLER_0_11_282/a_124_375# 0.018322f
C9526 _346_/a_257_69# _141_ 0.002092f
C9527 net56 state\[1\] 0.007364f
C9528 net64 FILLER_0_12_220/a_1468_375# 0.01836f
C9529 _005_ _192_/a_255_603# 0.001058f
C9530 FILLER_0_18_139/a_572_375# _145_ 0.00346f
C9531 _101_ mask\[1\] 0.033941f
C9532 _141_ FILLER_0_17_161/a_36_472# 0.011708f
C9533 _111_ _438_/a_36_151# 0.003619f
C9534 net82 fanout52/a_36_160# 0.026154f
C9535 trim[4] trim[1] 0.001879f
C9536 _185_ net17 0.270086f
C9537 _421_/a_2665_112# net19 0.01849f
C9538 _030_ _154_ 0.004803f
C9539 _305_/a_36_159# net76 0.010842f
C9540 net16 _408_/a_2215_68# 0.002096f
C9541 FILLER_0_20_15/a_932_472# net40 0.002705f
C9542 _010_ _419_/a_448_472# 0.003295f
C9543 _069_ _047_ 0.001975f
C9544 _053_ _439_/a_2248_156# 0.002486f
C9545 _187_ cal_count\[3\] 0.031898f
C9546 _430_/a_2665_112# FILLER_0_15_212/a_1380_472# 0.021761f
C9547 _058_ _125_ 0.016525f
C9548 FILLER_0_12_136/a_1380_472# state\[2\] 0.005779f
C9549 FILLER_0_24_274/a_1380_472# FILLER_0_23_282/a_484_472# 0.058411f
C9550 FILLER_0_17_200/a_124_375# FILLER_0_18_177/a_2724_472# 0.001597f
C9551 ctlp[2] _108_ 0.034027f
C9552 FILLER_0_18_2/a_2812_375# FILLER_0_20_15/a_1380_472# 0.001338f
C9553 net63 _337_/a_49_472# 0.001801f
C9554 FILLER_0_4_49/a_36_472# _160_ 0.00202f
C9555 FILLER_0_5_164/a_36_472# net37 0.008378f
C9556 FILLER_0_10_78/a_124_375# _120_ 0.006134f
C9557 _072_ _071_ 0.296543f
C9558 _354_/a_49_472# vdd -0.001073f
C9559 net53 state\[2\] 0.001982f
C9560 _254_/a_448_472# _074_ 0.002163f
C9561 _134_ FILLER_0_10_107/a_572_375# 0.047331f
C9562 _057_ _310_/a_49_472# 0.015839f
C9563 net55 _216_/a_255_603# 0.001011f
C9564 _093_ FILLER_0_16_89/a_1468_375# 0.003988f
C9565 FILLER_0_10_37/a_36_472# vss 0.003659f
C9566 _086_ _117_ 0.010287f
C9567 _415_/a_2248_156# vdd 0.009114f
C9568 _092_ FILLER_0_17_218/a_484_472# 0.007838f
C9569 state\[1\] _060_ 0.003973f
C9570 fanout60/a_36_160# result[3] 0.00188f
C9571 _188_ _067_ 0.001554f
C9572 _420_/a_1204_472# _009_ 0.009314f
C9573 FILLER_0_22_177/a_124_375# mask\[6\] 0.002672f
C9574 _450_/a_448_472# _039_ 0.047559f
C9575 _184_ vss 0.068129f
C9576 net22 _205_/a_36_160# 0.109939f
C9577 _176_ _451_/a_3081_151# 0.001255f
C9578 _379_/a_36_472# _160_ 0.023459f
C9579 _099_ FILLER_0_14_235/a_484_472# 0.00281f
C9580 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_36_472# 0.001723f
C9581 _101_ vss 0.05721f
C9582 trim_mask\[1\] _163_ 0.166315f
C9583 cal_count\[3\] _117_ 0.00114f
C9584 net18 _416_/a_1308_423# 0.021956f
C9585 FILLER_0_18_177/a_2812_375# net22 0.010501f
C9586 FILLER_0_8_138/a_124_375# _313_/a_67_603# 0.00744f
C9587 _443_/a_1308_423# net13 0.004098f
C9588 _443_/a_1000_472# net23 0.034596f
C9589 _449_/a_36_151# vdd 0.09324f
C9590 FILLER_0_3_78/a_484_472# _160_ 0.004988f
C9591 FILLER_0_13_65/a_124_375# _449_/a_36_151# 0.059049f
C9592 _106_ FILLER_0_17_226/a_124_375# 0.061857f
C9593 net52 _441_/a_2560_156# 0.004721f
C9594 net50 _441_/a_2248_156# 0.027849f
C9595 _440_/a_448_472# net47 0.016997f
C9596 FILLER_0_12_220/a_36_472# vdd 0.027911f
C9597 FILLER_0_12_220/a_1468_375# vss 0.057853f
C9598 _104_ net78 0.049954f
C9599 _104_ net60 0.063407f
C9600 FILLER_0_13_212/a_932_472# net79 0.006824f
C9601 _105_ _420_/a_2665_112# 0.001159f
C9602 FILLER_0_4_49/a_572_375# net49 0.004345f
C9603 net20 _223_/a_36_160# 0.066119f
C9604 net55 FILLER_0_18_37/a_1020_375# 0.005661f
C9605 _333_/a_36_160# _097_ 0.001332f
C9606 FILLER_0_4_107/a_484_472# _160_ 0.008194f
C9607 net41 _423_/a_36_151# 0.001134f
C9608 FILLER_0_17_72/a_572_375# vss 0.008057f
C9609 FILLER_0_17_72/a_1020_375# vdd 0.002541f
C9610 FILLER_0_8_37/a_484_472# vdd 0.009603f
C9611 _069_ _429_/a_36_151# 0.010076f
C9612 _443_/a_36_151# _442_/a_36_151# 0.06169f
C9613 FILLER_0_4_49/a_572_375# net68 0.023227f
C9614 net81 net19 0.786284f
C9615 net47 FILLER_0_4_91/a_484_472# 0.007531f
C9616 _274_/a_2124_68# net4 0.00137f
C9617 ctln[7] FILLER_0_0_130/a_36_472# 0.012298f
C9618 net74 _372_/a_1194_69# 0.002006f
C9619 _072_ FILLER_0_10_214/a_36_472# 0.015199f
C9620 net82 _443_/a_448_472# 0.007335f
C9621 _089_ vdd 0.087336f
C9622 net52 _439_/a_2665_112# 0.00117f
C9623 trimb[1] FILLER_0_18_2/a_1468_375# 0.002041f
C9624 _095_ FILLER_0_14_107/a_572_375# 0.01418f
C9625 result[9] ctlp[1] 0.074012f
C9626 FILLER_0_8_127/a_124_375# _129_ 0.056784f
C9627 result[8] _107_ 0.041984f
C9628 FILLER_0_17_56/a_36_472# _404_/a_36_472# 0.004546f
C9629 _425_/a_2248_156# net37 0.01491f
C9630 _371_/a_36_113# _159_ 0.021612f
C9631 mask\[4\] FILLER_0_18_177/a_2276_472# 0.016876f
C9632 _328_/a_36_113# _135_ 0.005635f
C9633 FILLER_0_13_100/a_124_375# vss 0.00513f
C9634 FILLER_0_13_100/a_36_472# vdd 0.021826f
C9635 net38 _450_/a_1353_112# 0.02208f
C9636 FILLER_0_18_209/a_484_472# _047_ 0.002188f
C9637 result[9] _417_/a_2248_156# 0.046399f
C9638 _131_ _331_/a_448_472# 0.007271f
C9639 _010_ _420_/a_2665_112# 0.029378f
C9640 _165_ FILLER_0_6_47/a_36_472# 0.077573f
C9641 cal_count\[2\] _180_ 0.153207f
C9642 _434_/a_2665_112# vdd 0.030225f
C9643 _071_ FILLER_0_13_142/a_1468_375# 0.007453f
C9644 net79 _284_/a_224_472# 0.009327f
C9645 FILLER_0_18_107/a_124_375# net14 0.005202f
C9646 ctlp[1] FILLER_0_23_282/a_36_472# 0.003169f
C9647 mask\[8\] _437_/a_1308_423# 0.001928f
C9648 fanout70/a_36_113# fanout73/a_36_113# 0.001578f
C9649 fanout81/a_36_160# net2 0.044793f
C9650 FILLER_0_12_136/a_36_472# vss 0.003185f
C9651 FILLER_0_12_136/a_484_472# vdd 0.005304f
C9652 _422_/a_1308_423# _009_ 0.008875f
C9653 _417_/a_796_472# vss 0.001608f
C9654 net49 FILLER_0_3_78/a_36_472# 0.059367f
C9655 _030_ FILLER_0_3_78/a_484_472# 0.007736f
C9656 _031_ FILLER_0_2_111/a_932_472# 0.017509f
C9657 net41 _064_ 0.301777f
C9658 _173_ _408_/a_728_93# 0.022838f
C9659 net58 _084_ 0.141836f
C9660 _036_ FILLER_0_3_78/a_124_375# 0.00215f
C9661 _065_ _447_/a_2665_112# 0.034757f
C9662 net74 FILLER_0_13_100/a_124_375# 0.005049f
C9663 _126_ FILLER_0_13_206/a_36_472# 0.026561f
C9664 net54 _050_ 0.040506f
C9665 net36 FILLER_0_18_76/a_572_375# 0.005153f
C9666 _443_/a_2248_156# net59 0.002471f
C9667 net70 vss 0.175272f
C9668 _272_/a_36_472# net76 0.04597f
C9669 _162_ _076_ 0.008623f
C9670 _411_/a_448_472# net8 0.04545f
C9671 net82 FILLER_0_2_177/a_572_375# 0.003837f
C9672 net34 net35 2.497277f
C9673 ctlp[6] mask\[7\] 0.011418f
C9674 cal_count\[2\] _452_/a_3129_107# 0.008853f
C9675 net78 _421_/a_1308_423# 0.015694f
C9676 net60 _421_/a_1308_423# 0.020693f
C9677 mask\[2\] vdd 0.433058f
C9678 net47 vss 0.919407f
C9679 _213_/a_67_603# _051_ 0.015959f
C9680 _099_ _098_ 0.018316f
C9681 _441_/a_2665_112# _164_ 0.021931f
C9682 FILLER_0_8_138/a_124_375# _058_ 0.009863f
C9683 _193_/a_36_160# result[3] 0.002218f
C9684 net47 _365_/a_692_472# 0.002051f
C9685 net57 _428_/a_36_151# 0.023215f
C9686 FILLER_0_4_213/a_124_375# vdd 0.009037f
C9687 net70 net74 0.017928f
C9688 net8 net59 0.062623f
C9689 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_36_472# 0.012267f
C9690 _069_ _055_ 0.741952f
C9691 net55 FILLER_0_18_61/a_36_472# 0.022296f
C9692 _440_/a_3041_156# _164_ 0.001221f
C9693 FILLER_0_14_91/a_484_472# _095_ 0.011772f
C9694 FILLER_0_1_192/a_36_472# net21 0.016033f
C9695 net74 net47 0.030815f
C9696 _095_ state\[1\] 0.069906f
C9697 result[7] vdd 0.500292f
C9698 net4 net8 0.00647f
C9699 _126_ FILLER_0_15_180/a_124_375# 0.001238f
C9700 _086_ FILLER_0_7_104/a_1020_375# 0.00757f
C9701 _119_ FILLER_0_7_104/a_1468_375# 0.022368f
C9702 FILLER_0_10_37/a_124_375# _042_ 0.002437f
C9703 _428_/a_36_151# _135_ 0.030608f
C9704 _063_ _445_/a_2665_112# 0.009759f
C9705 FILLER_0_7_72/a_3172_472# net50 0.001428f
C9706 FILLER_0_23_44/a_36_472# vdd 0.01833f
C9707 FILLER_0_23_44/a_1468_375# vss 0.055902f
C9708 net54 _433_/a_1000_472# 0.0025f
C9709 net64 _282_/a_36_160# 0.014431f
C9710 _255_/a_224_552# _070_ 0.001333f
C9711 _104_ _093_ 0.109158f
C9712 FILLER_0_21_125/a_124_375# _433_/a_36_151# 0.059049f
C9713 FILLER_0_17_64/a_124_375# _183_ 0.001236f
C9714 net57 _443_/a_36_151# 0.003322f
C9715 _072_ _246_/a_36_68# 0.064797f
C9716 cal_itt\[3\] _122_ 0.03282f
C9717 net18 net33 0.001671f
C9718 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1380_472# 0.013277f
C9719 _067_ FILLER_0_12_20/a_36_472# 0.015608f
C9720 _412_/a_1000_472# net59 0.00147f
C9721 mask\[3\] FILLER_0_16_154/a_572_375# 0.027873f
C9722 net72 FILLER_0_15_59/a_36_472# 0.049812f
C9723 _170_ net59 0.002301f
C9724 net72 _453_/a_36_151# 0.001607f
C9725 net32 vss 0.824307f
C9726 _098_ _202_/a_36_160# 0.006831f
C9727 _081_ _066_ 0.061358f
C9728 _416_/a_1308_423# net62 0.002665f
C9729 net73 _438_/a_2665_112# 0.001708f
C9730 _412_/a_2248_156# en 0.022108f
C9731 _429_/a_448_472# net62 0.002713f
C9732 _144_ vdd 0.40911f
C9733 _098_ _433_/a_2560_156# 0.004273f
C9734 FILLER_0_7_104/a_124_375# _153_ 0.001205f
C9735 FILLER_0_7_104/a_1020_375# _154_ 0.005051f
C9736 net65 _411_/a_36_151# 0.001415f
C9737 net17 _450_/a_2449_156# 0.05017f
C9738 _430_/a_36_151# _019_ 0.019296f
C9739 _028_ FILLER_0_5_72/a_1468_375# 0.00123f
C9740 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3260_375# 0.086635f
C9741 _091_ FILLER_0_18_177/a_484_472# 0.004272f
C9742 _189_/a_67_603# net62 0.001695f
C9743 FILLER_0_12_124/a_124_375# vdd -0.00168f
C9744 FILLER_0_18_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001684f
C9745 output36/a_224_472# vss -0.002521f
C9746 FILLER_0_9_60/a_124_375# vss 0.003217f
C9747 FILLER_0_9_60/a_572_375# vdd 0.031403f
C9748 _077_ _439_/a_796_472# 0.007471f
C9749 net47 _452_/a_836_156# 0.002075f
C9750 _154_ _156_ 0.019471f
C9751 FILLER_0_10_214/a_124_375# _090_ 0.072741f
C9752 net44 net3 0.195171f
C9753 mask\[9\] _438_/a_2560_156# 0.008709f
C9754 _236_/a_36_160# trim[1] 0.003604f
C9755 FILLER_0_15_290/a_36_472# vdd 0.092839f
C9756 FILLER_0_15_290/a_124_375# vss 0.032056f
C9757 FILLER_0_7_146/a_124_375# _372_/a_170_472# 0.001188f
C9758 output11/a_224_472# net75 0.015211f
C9759 FILLER_0_3_172/a_484_472# net22 0.012284f
C9760 _418_/a_2665_112# _417_/a_2665_112# 0.00131f
C9761 _386_/a_848_380# net22 0.00429f
C9762 FILLER_0_9_28/a_484_472# net41 0.042989f
C9763 _226_/a_1044_68# net21 0.001903f
C9764 net66 _166_ 0.011066f
C9765 _081_ FILLER_0_8_156/a_484_472# 0.001772f
C9766 cal_itt\[3\] _061_ 0.001311f
C9767 _343_/a_49_472# _141_ 0.04106f
C9768 _424_/a_448_472# _012_ 0.007299f
C9769 _081_ net37 1.274337f
C9770 net63 _202_/a_36_160# 0.004414f
C9771 net7 _064_ 0.001538f
C9772 _095_ _402_/a_718_527# 0.002109f
C9773 trimb[1] _452_/a_2449_156# 0.001681f
C9774 _282_/a_36_160# vss 0.005221f
C9775 FILLER_0_8_24/a_124_375# net42 0.032303f
C9776 net35 FILLER_0_22_177/a_124_375# 0.0073f
C9777 _044_ FILLER_0_14_263/a_36_472# 0.002013f
C9778 FILLER_0_22_86/a_572_375# net71 0.002239f
C9779 FILLER_0_5_128/a_484_472# net47 0.009309f
C9780 net44 _245_/a_672_472# 0.001285f
C9781 _178_ _179_ 0.063494f
C9782 FILLER_0_10_78/a_1468_375# _114_ 0.01836f
C9783 _131_ _404_/a_36_472# 0.031567f
C9784 FILLER_0_17_282/a_124_375# vss 0.024404f
C9785 FILLER_0_17_282/a_36_472# vdd 0.107351f
C9786 _448_/a_1308_423# vdd 0.006042f
C9787 output9/a_224_472# fanout76/a_36_160# 0.016067f
C9788 _087_ FILLER_0_5_181/a_36_472# 0.154469f
C9789 _033_ net17 0.028529f
C9790 FILLER_0_14_235/a_124_375# net62 0.015659f
C9791 _088_ FILLER_0_3_172/a_2812_375# 0.002239f
C9792 FILLER_0_14_107/a_1020_375# vdd 0.008956f
C9793 ctlp[1] FILLER_0_24_290/a_124_375# 0.050488f
C9794 _431_/a_1000_472# _137_ 0.010168f
C9795 _063_ FILLER_0_6_37/a_36_472# 0.014315f
C9796 FILLER_0_22_177/a_1020_375# vdd 0.001695f
C9797 _115_ FILLER_0_9_72/a_1468_375# 0.025664f
C9798 _114_ FILLER_0_9_72/a_1380_472# 0.001043f
C9799 FILLER_0_1_98/a_36_472# trim_mask\[3\] 0.106084f
C9800 net69 _441_/a_1000_472# 0.018209f
C9801 _304_/a_224_472# mask\[9\] 0.003125f
C9802 net81 fanout58/a_36_160# 0.005575f
C9803 _072_ net23 0.006278f
C9804 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_484_472# 0.013277f
C9805 cal_itt\[2\] FILLER_0_3_221/a_1020_375# 0.010951f
C9806 FILLER_0_5_109/a_124_375# vdd 0.060786f
C9807 net81 cal_itt\[0\] 0.001048f
C9808 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_36_472# 0.086742f
C9809 fanout73/a_36_113# vdd 0.048166f
C9810 FILLER_0_16_37/a_36_472# _402_/a_1296_93# 0.001477f
C9811 _447_/a_448_472# net69 0.001694f
C9812 _069_ _315_/a_36_68# 0.002242f
C9813 _077_ _374_/a_36_68# 0.012411f
C9814 net63 FILLER_0_17_218/a_36_472# 0.003889f
C9815 net49 _029_ 0.004408f
C9816 FILLER_0_7_72/a_2276_472# _077_ 0.00475f
C9817 _059_ FILLER_0_5_148/a_124_375# 0.007657f
C9818 fanout66/a_36_113# vss 0.014789f
C9819 _122_ FILLER_0_5_164/a_36_472# 0.002232f
C9820 fanout57/a_36_113# trim_val\[4\] 0.078297f
C9821 net34 FILLER_0_22_128/a_1468_375# 0.003214f
C9822 _436_/a_1000_472# net54 0.002051f
C9823 net68 _029_ 0.094915f
C9824 FILLER_0_9_28/a_2364_375# _077_ 0.00397f
C9825 _137_ FILLER_0_15_180/a_124_375# 0.003108f
C9826 FILLER_0_8_127/a_36_472# _077_ 0.003023f
C9827 net20 FILLER_0_12_220/a_572_375# 0.007386f
C9828 _253_/a_36_68# _073_ 0.027664f
C9829 net52 FILLER_0_5_72/a_124_375# 0.029702f
C9830 _155_ _153_ 0.033366f
C9831 _450_/a_448_472# clkc 0.003011f
C9832 _450_/a_1040_527# net6 0.019715f
C9833 fanout68/a_36_113# _065_ 0.005586f
C9834 _415_/a_448_472# FILLER_0_11_282/a_124_375# 0.008952f
C9835 vdd rstn 0.160093f
C9836 FILLER_0_20_107/a_124_375# FILLER_0_20_98/a_124_375# 0.003228f
C9837 FILLER_0_12_136/a_1468_375# cal_count\[3\] 0.004337f
C9838 result[9] _418_/a_2248_156# 0.043716f
C9839 FILLER_0_18_177/a_2364_375# vdd 0.020562f
C9840 _410_/a_36_68# _187_ 0.038745f
C9841 _132_ _428_/a_796_472# 0.001472f
C9842 _350_/a_665_69# mask\[6\] 0.001069f
C9843 _339_/a_36_160# vdd 0.01226f
C9844 _372_/a_358_69# _163_ 0.001427f
C9845 _116_ _120_ 0.005759f
C9846 _428_/a_448_472# _131_ 0.041178f
C9847 _093_ FILLER_0_18_107/a_2812_375# 0.00626f
C9848 ctln[1] FILLER_0_0_266/a_36_472# 0.011046f
C9849 _291_/a_36_160# output18/a_224_472# 0.001175f
C9850 _418_/a_796_472# vss 0.00145f
C9851 _096_ _095_ 0.086147f
C9852 _411_/a_1204_472# _000_ 0.002575f
C9853 _411_/a_2665_112# net75 0.005223f
C9854 _076_ FILLER_0_8_156/a_124_375# 0.0062f
C9855 _070_ FILLER_0_8_156/a_36_472# 0.001338f
C9856 _106_ _069_ 0.006716f
C9857 _354_/a_49_472# _433_/a_36_151# 0.001715f
C9858 output9/a_224_472# _412_/a_448_472# 0.001025f
C9859 net26 FILLER_0_21_28/a_1828_472# 0.010367f
C9860 net41 _444_/a_2248_156# 0.028267f
C9861 FILLER_0_2_171/a_36_472# net22 0.081357f
C9862 FILLER_0_14_91/a_484_472# vss 0.003257f
C9863 net61 ctlp[1] 2.770871f
C9864 state\[1\] vss 0.294171f
C9865 net36 _094_ 0.086414f
C9866 _453_/a_2665_112# vss 0.037567f
C9867 _026_ _437_/a_1308_423# 0.018479f
C9868 _149_ _437_/a_1000_472# 0.019115f
C9869 net41 _446_/a_448_472# 0.040165f
C9870 _053_ FILLER_0_5_54/a_124_375# 0.001571f
C9871 net67 FILLER_0_12_20/a_124_375# 0.007044f
C9872 net57 _085_ 0.211414f
C9873 net57 FILLER_0_5_164/a_124_375# 0.040872f
C9874 net28 _426_/a_36_151# 0.004878f
C9875 _012_ FILLER_0_21_60/a_484_472# 0.01517f
C9876 net22 _047_ 0.132529f
C9877 net58 calibrate 0.205792f
C9878 _086_ _326_/a_36_160# 0.063565f
C9879 FILLER_0_15_212/a_932_472# mask\[1\] 0.014799f
C9880 state\[2\] _071_ 0.04575f
C9881 mask\[6\] _146_ 0.181681f
C9882 fanout53/a_36_160# net23 0.007461f
C9883 FILLER_0_13_142/a_1468_375# net23 0.011746f
C9884 _258_/a_36_160# _078_ 0.006096f
C9885 output13/a_224_472# net52 0.018089f
C9886 _425_/a_2665_112# calibrate 0.029064f
C9887 _008_ _106_ 0.034748f
C9888 FILLER_0_20_2/a_484_472# vdd 0.001049f
C9889 FILLER_0_9_28/a_2364_375# _453_/a_36_151# 0.001597f
C9890 _018_ FILLER_0_15_205/a_36_472# 0.00273f
C9891 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_484_472# 0.026657f
C9892 FILLER_0_13_212/a_36_472# net62 0.015187f
C9893 _335_/a_49_472# _098_ 0.001047f
C9894 fanout52/a_36_160# _443_/a_2665_112# 0.007884f
C9895 FILLER_0_1_266/a_484_472# vdd 0.003622f
C9896 _077_ FILLER_0_7_59/a_484_472# 0.001371f
C9897 FILLER_0_8_107/a_36_472# _134_ 0.005632f
C9898 _187_ _120_ 0.144679f
C9899 FILLER_0_2_165/a_36_472# net22 0.028367f
C9900 mask\[5\] FILLER_0_20_193/a_572_375# 0.036451f
C9901 FILLER_0_3_54/a_124_375# vdd 0.029897f
C9902 FILLER_0_9_28/a_2276_472# net68 0.023299f
C9903 _072_ _056_ 0.061377f
C9904 net82 _082_ 0.286003f
C9905 _415_/a_36_151# FILLER_0_8_263/a_124_375# 0.001619f
C9906 result[7] net78 0.019651f
C9907 result[7] net60 0.778099f
C9908 result[8] FILLER_0_24_274/a_1380_472# 0.005458f
C9909 FILLER_0_12_2/a_572_375# net67 0.007509f
C9910 mask\[4\] FILLER_0_19_195/a_36_472# 0.004669f
C9911 FILLER_0_6_47/a_36_472# vss 0.002433f
C9912 FILLER_0_6_47/a_484_472# vdd 0.005065f
C9913 FILLER_0_15_212/a_1380_472# vdd 0.003213f
C9914 FILLER_0_15_212/a_932_472# vss 0.019114f
C9915 _429_/a_36_151# net22 0.020582f
C9916 _093_ FILLER_0_17_72/a_1020_375# 0.001994f
C9917 net32 _103_ 0.038496f
C9918 _337_/a_49_472# _137_ 0.046633f
C9919 _308_/a_848_380# _219_/a_36_160# 0.001045f
C9920 _323_/a_36_113# net27 0.010949f
C9921 _104_ output33/a_224_472# 0.032929f
C9922 FILLER_0_14_181/a_124_375# _098_ 0.005696f
C9923 FILLER_0_4_49/a_572_375# net47 0.00654f
C9924 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_932_472# 0.001723f
C9925 output13/a_224_472# _387_/a_36_113# 0.020974f
C9926 _425_/a_36_151# FILLER_0_8_247/a_124_375# 0.001597f
C9927 FILLER_0_7_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001723f
C9928 net81 _429_/a_36_151# 0.018551f
C9929 _009_ FILLER_0_23_282/a_484_472# 0.009744f
C9930 FILLER_0_4_197/a_1468_375# net22 0.009108f
C9931 FILLER_0_8_247/a_932_472# calibrate 0.008694f
C9932 _053_ _164_ 0.058788f
C9933 _418_/a_36_151# net77 0.019316f
C9934 net52 net50 0.702793f
C9935 mask\[8\] _051_ 0.003475f
C9936 FILLER_0_15_150/a_36_472# net36 0.012318f
C9937 _105_ vss 0.485198f
C9938 _422_/a_796_472# mask\[7\] 0.001755f
C9939 net38 net43 0.016358f
C9940 net52 _443_/a_1204_472# 0.005165f
C9941 _096_ mask\[1\] 0.010488f
C9942 net39 _033_ 0.607942f
C9943 cal_count\[2\] FILLER_0_15_2/a_572_375# 0.015401f
C9944 FILLER_0_19_125/a_36_472# _145_ 0.004858f
C9945 _430_/a_36_151# net80 0.082603f
C9946 net2 rstn 0.002598f
C9947 _289_/a_36_472# vdd 0.006886f
C9948 _446_/a_2248_156# _160_ 0.002464f
C9949 _055_ _090_ 0.040233f
C9950 _077_ FILLER_0_9_72/a_1380_472# 0.006408f
C9951 net15 FILLER_0_6_47/a_2812_375# 0.002944f
C9952 net72 _095_ 0.136566f
C9953 _051_ vss 0.050185f
C9954 _415_/a_1000_472# result[1] 0.005365f
C9955 FILLER_0_16_89/a_36_472# _131_ 0.013616f
C9956 _074_ net76 0.026801f
C9957 _086_ _375_/a_36_68# 0.038443f
C9958 fanout68/a_36_113# _036_ 0.007847f
C9959 FILLER_0_4_107/a_36_472# net47 0.002982f
C9960 _010_ vss 0.064717f
C9961 _430_/a_1308_423# net63 0.01125f
C9962 FILLER_0_21_125/a_572_375# _098_ 0.006462f
C9963 _093_ mask\[2\] 0.009354f
C9964 FILLER_0_2_93/a_572_375# _367_/a_36_68# 0.001069f
C9965 FILLER_0_5_181/a_124_375# vss 0.011456f
C9966 FILLER_0_5_181/a_36_472# vdd 0.081434f
C9967 FILLER_0_4_197/a_124_375# _088_ 0.024641f
C9968 FILLER_0_21_28/a_1020_375# vdd 0.04353f
C9969 _031_ net14 0.00913f
C9970 FILLER_0_3_172/a_36_472# vdd 0.006145f
C9971 FILLER_0_3_172/a_3260_375# vss 0.054783f
C9972 _386_/a_124_24# vdd 0.014293f
C9973 FILLER_0_16_241/a_36_472# net30 0.001025f
C9974 FILLER_0_9_223/a_572_375# _076_ 0.034523f
C9975 FILLER_0_9_223/a_124_375# _068_ 0.010485f
C9976 net80 _333_/a_36_160# 0.001594f
C9977 net41 net50 0.002438f
C9978 _449_/a_1000_472# net55 0.001617f
C9979 FILLER_0_4_177/a_484_472# FILLER_0_2_177/a_572_375# 0.001512f
C9980 FILLER_0_17_200/a_572_375# net21 0.011557f
C9981 net4 FILLER_0_3_221/a_1020_375# 0.006974f
C9982 _438_/a_1000_472# net14 0.003275f
C9983 FILLER_0_2_111/a_36_472# _157_ 0.104961f
C9984 FILLER_0_5_54/a_124_375# _164_ 0.004076f
C9985 _055_ net22 0.084669f
C9986 output25/a_224_472# _214_/a_36_160# 0.027335f
C9987 _385_/a_36_68# vss 0.002408f
C9988 net60 FILLER_0_17_282/a_36_472# 0.009978f
C9989 FILLER_0_18_100/a_124_375# vdd 0.044014f
C9990 _413_/a_1204_472# net82 0.00291f
C9991 FILLER_0_17_56/a_36_472# _183_ 0.056523f
C9992 _077_ _308_/a_692_472# 0.002268f
C9993 _081_ _122_ 2.557248f
C9994 _152_ calibrate 0.020369f
C9995 result[7] _093_ 0.001096f
C9996 _446_/a_2560_156# net66 0.002649f
C9997 output9/a_224_472# net58 0.050634f
C9998 _144_ _433_/a_36_151# 0.086558f
C9999 _114_ _171_ 0.203692f
C10000 FILLER_0_6_239/a_36_472# net76 0.011803f
C10001 ctlp[4] ctlp[5] 0.001257f
C10002 ctln[1] net82 0.001141f
C10003 _062_ _226_/a_1044_68# 0.001944f
C10004 _096_ vss 0.126096f
C10005 trim_mask\[2\] fanout49/a_36_160# 0.12844f
C10006 net52 trim_mask\[3\] 0.666362f
C10007 _005_ _416_/a_1000_472# 0.027013f
C10008 net56 _145_ 0.009307f
C10009 net54 FILLER_0_18_139/a_932_472# 0.003365f
C10010 _443_/a_1308_423# _170_ 0.043472f
C10011 _092_ _091_ 0.028594f
C10012 _132_ FILLER_0_17_104/a_1020_375# 0.009251f
C10013 net76 FILLER_0_3_172/a_1020_375# 0.007439f
C10014 _415_/a_448_472# FILLER_0_9_270/a_36_472# 0.012285f
C10015 _131_ FILLER_0_17_104/a_124_375# 0.006681f
C10016 _144_ _147_ 0.057955f
C10017 FILLER_0_11_64/a_36_472# _038_ 0.001822f
C10018 _451_/a_3129_107# vdd 0.008569f
C10019 ctln[1] _411_/a_2248_156# 0.013381f
C10020 FILLER_0_5_72/a_932_472# trim_mask\[1\] 0.014619f
C10021 _395_/a_36_488# _070_ 0.005165f
C10022 _176_ _131_ 1.798819f
C10023 cal_itt\[1\] vdd 0.410279f
C10024 FILLER_0_13_212/a_572_375# _248_/a_36_68# 0.030745f
C10025 FILLER_0_4_152/a_36_472# _386_/a_124_24# 0.004755f
C10026 _431_/a_2560_156# _136_ 0.013111f
C10027 _325_/a_224_472# _130_ 0.001685f
C10028 net57 FILLER_0_16_154/a_484_472# 0.001532f
C10029 ctln[3] FILLER_0_0_232/a_36_472# 0.015594f
C10030 FILLER_0_7_233/a_36_472# vdd 0.016804f
C10031 FILLER_0_7_233/a_124_375# vss 0.003952f
C10032 en_co_clk net53 0.001712f
C10033 net35 _146_ 0.096468f
C10034 net38 _452_/a_448_472# 0.016895f
C10035 _014_ calibrate 0.403103f
C10036 _114_ _176_ 0.147182f
C10037 _431_/a_1308_423# net73 0.039024f
C10038 _414_/a_2665_112# _122_ 0.007441f
C10039 valid vdd 0.148392f
C10040 FILLER_0_12_28/a_124_375# _039_ 0.004669f
C10041 trimb[1] FILLER_0_19_28/a_36_472# 0.01233f
C10042 mask\[3\] FILLER_0_18_177/a_572_375# 0.002924f
C10043 _098_ FILLER_0_16_154/a_932_472# 0.001701f
C10044 _114_ _306_/a_36_68# 0.032258f
C10045 state\[1\] _097_ 0.004171f
C10046 net60 _418_/a_1000_472# 0.007557f
C10047 cal_itt\[2\] vdd 0.267121f
C10048 _207_/a_255_603# mask\[6\] 0.003114f
C10049 vdd FILLER_0_13_72/a_572_375# -0.001166f
C10050 vss FILLER_0_13_72/a_124_375# 0.043492f
C10051 net58 FILLER_0_9_282/a_36_472# 0.062389f
C10052 trimb[0] trimb[3] 0.549457f
C10053 result[4] _417_/a_448_472# 0.003485f
C10054 output31/a_224_472# _417_/a_2248_156# 0.024448f
C10055 _390_/a_36_68# _067_ 0.029588f
C10056 net47 _380_/a_224_472# 0.001405f
C10057 _432_/a_796_472# _091_ 0.018082f
C10058 _155_ trim_mask\[1\] 0.006536f
C10059 FILLER_0_23_60/a_36_472# vss 0.006794f
C10060 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_484_472# 0.013276f
C10061 _053_ _072_ 0.001774f
C10062 _178_ _181_ 0.188669f
C10063 FILLER_0_6_177/a_572_375# vss 0.008666f
C10064 FILLER_0_6_177/a_36_472# vdd 0.109918f
C10065 trim_mask\[4\] _369_/a_36_68# 0.00407f
C10066 _408_/a_718_524# _067_ 0.006516f
C10067 _076_ _055_ 0.056585f
C10068 net74 FILLER_0_13_72/a_124_375# 0.014594f
C10069 ctlp[8] net25 0.055914f
C10070 net65 FILLER_0_2_177/a_572_375# 0.017058f
C10071 FILLER_0_2_171/a_124_375# vdd 0.042659f
C10072 net55 FILLER_0_11_78/a_36_472# 0.059367f
C10073 _127_ FILLER_0_11_142/a_124_375# 0.00205f
C10074 net32 _295_/a_36_472# 0.002637f
C10075 _070_ calibrate 0.675125f
C10076 _068_ net59 0.001388f
C10077 state\[2\] net23 0.331644f
C10078 output35/a_224_472# vdd 0.064053f
C10079 ctlp[4] _107_ 0.080312f
C10080 net4 _068_ 0.040977f
C10081 _126_ _171_ 0.01633f
C10082 FILLER_0_16_255/a_36_472# _006_ 0.006621f
C10083 FILLER_0_4_123/a_124_375# _159_ 0.023643f
C10084 _399_/a_224_472# _179_ 0.002288f
C10085 _402_/a_728_93# _182_ 0.00263f
C10086 net44 _190_/a_36_160# 0.015628f
C10087 FILLER_0_15_72/a_124_375# FILLER_0_15_59/a_572_375# 0.003228f
C10088 _423_/a_36_151# FILLER_0_23_44/a_1380_472# 0.001723f
C10089 FILLER_0_7_104/a_1380_472# _125_ 0.001279f
C10090 _068_ _311_/a_692_473# 0.002377f
C10091 _427_/a_1204_472# _095_ 0.006692f
C10092 net68 FILLER_0_5_54/a_484_472# 0.047601f
C10093 _144_ _436_/a_36_151# 0.029716f
C10094 _074_ _083_ 0.035769f
C10095 FILLER_0_5_198/a_572_375# net22 0.029657f
C10096 _076_ _313_/a_67_603# 0.024219f
C10097 net18 net62 0.089041f
C10098 FILLER_0_18_2/a_2724_472# net47 0.001551f
C10099 FILLER_0_4_99/a_36_472# vss 0.002273f
C10100 trim_mask\[4\] net23 0.180803f
C10101 FILLER_0_5_54/a_1380_472# trim_mask\[1\] 0.01205f
C10102 net72 vss 0.472104f
C10103 FILLER_0_2_165/a_124_375# vdd 0.020315f
C10104 _118_ _315_/a_716_497# 0.001968f
C10105 FILLER_0_9_223/a_124_375# vdd 0.006153f
C10106 FILLER_0_13_65/a_36_472# net72 0.00272f
C10107 _445_/a_36_151# net47 0.002364f
C10108 FILLER_0_4_99/a_124_375# _365_/a_36_68# 0.001918f
C10109 _029_ net47 2.210804f
C10110 _451_/a_36_151# net14 0.037503f
C10111 _095_ _281_/a_672_472# 0.00134f
C10112 _076_ FILLER_0_6_231/a_124_375# 0.001382f
C10113 _070_ FILLER_0_6_231/a_36_472# 0.001096f
C10114 net79 FILLER_0_15_282/a_484_472# 0.006575f
C10115 net36 net21 0.034415f
C10116 _369_/a_244_472# vdd 0.001255f
C10117 _021_ _143_ 0.007778f
C10118 net17 _452_/a_2225_156# 0.001943f
C10119 net82 FILLER_0_4_213/a_572_375# 0.00123f
C10120 _443_/a_448_472# net69 0.068491f
C10121 net79 _113_ 0.002432f
C10122 net32 net31 0.023293f
C10123 FILLER_0_9_142/a_124_375# _122_ 0.004711f
C10124 _093_ FILLER_0_18_177/a_2364_375# 0.001989f
C10125 _131_ _183_ 0.227229f
C10126 trim_mask\[2\] FILLER_0_4_91/a_36_472# 0.003327f
C10127 _126_ _176_ 0.057877f
C10128 net82 _032_ 0.014269f
C10129 fanout74/a_36_113# trim_mask\[4\] 0.026261f
C10130 net72 net74 0.035298f
C10131 net2 cal_itt\[1\] 0.284695f
C10132 _033_ net42 0.002707f
C10133 _144_ _346_/a_257_69# 0.001089f
C10134 _306_/a_36_68# _126_ 0.01893f
C10135 vdd _416_/a_36_151# 0.142481f
C10136 _116_ _043_ 0.002037f
C10137 output27/a_224_472# FILLER_0_9_282/a_124_375# 0.029138f
C10138 ctln[4] net21 0.009947f
C10139 _114_ FILLER_0_13_142/a_124_375# 0.00191f
C10140 net52 FILLER_0_0_130/a_36_472# 0.002743f
C10141 _430_/a_2665_112# fanout63/a_36_160# 0.010365f
C10142 net16 trim_val\[2\] 0.124462f
C10143 _257_/a_36_472# _077_ 0.019883f
C10144 _025_ _437_/a_2665_112# 0.001245f
C10145 output16/a_224_472# _447_/a_2248_156# 0.001937f
C10146 ctln[9] _447_/a_448_472# 0.003564f
C10147 net16 _447_/a_796_472# 0.003278f
C10148 net57 FILLER_0_13_100/a_36_472# 0.077963f
C10149 _013_ FILLER_0_21_28/a_1916_375# 0.006025f
C10150 net72 cal_count\[1\] 0.13509f
C10151 valid net2 0.062523f
C10152 _065_ net69 0.051511f
C10153 _379_/a_36_472# trim_val\[1\] 0.00909f
C10154 FILLER_0_4_197/a_1020_375# vdd 0.002455f
C10155 mask\[1\] FILLER_0_15_180/a_124_375# 0.004011f
C10156 FILLER_0_22_86/a_124_375# _098_ 0.011864f
C10157 FILLER_0_16_107/a_484_472# net14 0.001528f
C10158 _000_ net8 0.021422f
C10159 _449_/a_2248_156# FILLER_0_13_80/a_124_375# 0.001068f
C10160 _024_ vss 0.132549f
C10161 _424_/a_36_151# vss 0.030774f
C10162 _424_/a_448_472# vdd 0.014219f
C10163 vdd net40 1.984115f
C10164 _083_ FILLER_0_3_221/a_484_472# 0.02695f
C10165 _441_/a_1000_472# vss 0.01858f
C10166 _066_ _386_/a_692_472# 0.001958f
C10167 net54 _437_/a_36_151# 0.019307f
C10168 _098_ _434_/a_2560_156# 0.003888f
C10169 trim_mask\[2\] vdd 0.376424f
C10170 FILLER_0_11_64/a_124_375# vdd 0.045435f
C10171 _088_ _080_ 0.003418f
C10172 _070_ _125_ 0.125523f
C10173 _076_ _058_ 0.912225f
C10174 _428_/a_2665_112# FILLER_0_13_142/a_124_375# 0.003325f
C10175 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_572_375# 0.086635f
C10176 net55 _452_/a_448_472# 0.05323f
C10177 _015_ _426_/a_1000_472# 0.033582f
C10178 FILLER_0_13_206/a_36_472# vss 0.003985f
C10179 _193_/a_36_160# FILLER_0_13_290/a_36_472# 0.004828f
C10180 _447_/a_1308_423# vdd 0.004739f
C10181 FILLER_0_18_2/a_3260_375# vdd 0.046682f
C10182 trim_val\[3\] _164_ 0.018411f
C10183 _068_ _315_/a_716_497# 0.00217f
C10184 _076_ _315_/a_36_68# 0.001568f
C10185 _070_ _315_/a_1657_68# 0.001601f
C10186 output39/a_224_472# trim[1] 0.061797f
C10187 _115_ FILLER_0_9_105/a_484_472# 0.004075f
C10188 _187_ _043_ 0.011995f
C10189 _101_ _100_ 0.012073f
C10190 _431_/a_1000_472# vss 0.002491f
C10191 _096_ _097_ 0.038778f
C10192 net57 mask\[2\] 0.022012f
C10193 _440_/a_2560_156# vss 0.002793f
C10194 _126_ FILLER_0_14_181/a_124_375# 0.004632f
C10195 _116_ net21 0.036746f
C10196 mask\[2\] FILLER_0_15_205/a_36_472# 0.001204f
C10197 net29 net30 0.053996f
C10198 _430_/a_1000_472# _069_ 0.00929f
C10199 _439_/a_796_472# vss 0.003859f
C10200 input3/a_36_113# vdd 0.117445f
C10201 _091_ FILLER_0_13_212/a_932_472# 0.008749f
C10202 FILLER_0_10_78/a_1380_472# FILLER_0_10_94/a_36_472# 0.013277f
C10203 _077_ _176_ 0.00497f
C10204 net17 output41/a_224_472# 0.030456f
C10205 _412_/a_796_472# net58 0.001182f
C10206 _431_/a_1308_423# _427_/a_36_151# 0.001256f
C10207 _086_ _134_ 0.020487f
C10208 _411_/a_36_151# vss 0.035447f
C10209 _176_ FILLER_0_10_107/a_124_375# 0.013408f
C10210 _098_ _437_/a_1000_472# 0.007963f
C10211 FILLER_0_7_72/a_36_472# _439_/a_448_472# 0.008036f
C10212 FILLER_0_7_104/a_484_472# _131_ 0.00432f
C10213 _008_ net30 1.112351f
C10214 _359_/a_36_488# _062_ 0.005596f
C10215 net36 _438_/a_1204_472# 0.012234f
C10216 _132_ _318_/a_224_472# 0.001097f
C10217 mask\[7\] vdd 1.098711f
C10218 _316_/a_1084_68# vdd 0.001166f
C10219 cal_count\[3\] _134_ 0.011364f
C10220 net63 _434_/a_2560_156# 0.014333f
C10221 FILLER_0_15_180/a_572_375# vdd 0.068901f
C10222 net15 _441_/a_1308_423# 0.009697f
C10223 _155_ FILLER_0_7_104/a_572_375# 0.002336f
C10224 net59 vdd 2.180407f
C10225 mask\[5\] FILLER_0_20_177/a_932_472# 0.016114f
C10226 FILLER_0_16_57/a_572_375# net55 0.004559f
C10227 FILLER_0_16_57/a_36_472# net72 0.040135f
C10228 _126_ _320_/a_672_472# 0.003662f
C10229 _148_ vdd 0.01565f
C10230 ctlp[3] _104_ 0.025066f
C10231 net35 _435_/a_448_472# 0.007865f
C10232 net4 vdd 1.218939f
C10233 trim_val\[4\] trim_mask\[4\] 0.152123f
C10234 _028_ FILLER_0_6_79/a_36_472# 0.016281f
C10235 _086_ FILLER_0_6_177/a_124_375# 0.043788f
C10236 _035_ _167_ 0.01574f
C10237 net7 ctln[0] 0.001209f
C10238 net15 _439_/a_448_472# 0.038829f
C10239 _452_/a_1040_527# net40 0.007832f
C10240 mask\[5\] FILLER_0_18_177/a_572_375# 0.002653f
C10241 FILLER_0_7_146/a_36_472# _068_ 0.012745f
C10242 _114_ FILLER_0_10_94/a_124_375# 0.040691f
C10243 _432_/a_1308_423# FILLER_0_18_177/a_36_472# 0.009119f
C10244 result[4] _418_/a_448_472# 0.004918f
C10245 output31/a_224_472# _418_/a_2248_156# 0.023576f
C10246 net36 FILLER_0_15_212/a_1020_375# 0.004863f
C10247 _435_/a_796_472# vdd 0.003478f
C10248 _448_/a_2560_156# net59 0.007516f
C10249 fanout66/a_36_113# _029_ 0.001684f
C10250 _085_ _267_/a_672_472# 0.006682f
C10251 _116_ _267_/a_1568_472# 0.001147f
C10252 _326_/a_36_160# FILLER_0_9_105/a_572_375# 0.005489f
C10253 _132_ _136_ 0.034253f
C10254 _176_ FILLER_0_15_59/a_36_472# 0.00622f
C10255 FILLER_0_18_171/a_124_375# _091_ 0.034351f
C10256 _370_/a_124_24# net47 0.017609f
C10257 _408_/a_728_93# _184_ 0.001389f
C10258 _028_ FILLER_0_8_107/a_36_472# 0.002173f
C10259 _374_/a_36_68# vss 0.047832f
C10260 FILLER_0_24_274/a_36_472# FILLER_0_23_274/a_36_472# 0.05841f
C10261 _427_/a_2248_156# vdd -0.002315f
C10262 _427_/a_1204_472# vss 0.0041f
C10263 sample calibrate 0.001861f
C10264 _141_ mask\[6\] 0.009844f
C10265 _232_/a_67_603# trim_mask\[1\] 0.022808f
C10266 FILLER_0_7_72/a_2724_472# vdd 0.007669f
C10267 _335_/a_49_472# _137_ 0.03139f
C10268 FILLER_0_15_235/a_572_375# net62 0.001315f
C10269 FILLER_0_15_282/a_572_375# net18 0.00298f
C10270 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_124_375# 0.026339f
C10271 FILLER_0_9_28/a_2812_375# vdd 0.016637f
C10272 FILLER_0_9_223/a_572_375# _128_ 0.006559f
C10273 net52 net22 0.017993f
C10274 FILLER_0_8_24/a_572_375# _054_ 0.004858f
C10275 FILLER_0_8_127/a_36_472# vss 0.004344f
C10276 vss FILLER_0_21_60/a_36_472# 0.001384f
C10277 vdd FILLER_0_21_60/a_484_472# 0.005181f
C10278 _276_/a_36_160# FILLER_0_17_218/a_36_472# 0.035111f
C10279 _451_/a_1353_112# _040_ 0.005265f
C10280 net81 fanout76/a_36_160# 0.041089f
C10281 _117_ net21 0.016722f
C10282 _043_ _225_/a_36_160# 0.007958f
C10283 FILLER_0_7_162/a_124_375# vss 0.018732f
C10284 FILLER_0_7_162/a_36_472# vdd 0.026981f
C10285 net82 net19 1.14585f
C10286 _093_ FILLER_0_18_100/a_124_375# 0.011632f
C10287 _427_/a_1204_472# net74 0.003057f
C10288 _332_/a_36_472# vdd 0.017097f
C10289 net27 FILLER_0_8_263/a_36_472# 0.003956f
C10290 FILLER_0_8_138/a_124_375# _070_ 0.002997f
C10291 _059_ _120_ 0.0127f
C10292 FILLER_0_22_177/a_932_472# net33 0.014021f
C10293 net68 _453_/a_1308_423# 0.002195f
C10294 FILLER_0_7_104/a_1020_375# _151_ 0.002336f
C10295 FILLER_0_1_98/a_124_375# vdd 0.036865f
C10296 FILLER_0_8_127/a_36_472# net74 0.063481f
C10297 _411_/a_2248_156# net19 0.001197f
C10298 FILLER_0_13_212/a_1020_375# vdd -0.014642f
C10299 FILLER_0_13_212/a_572_375# vss 0.007991f
C10300 _053_ _133_ 0.288819f
C10301 _013_ net55 0.239055f
C10302 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_124_375# 0.003228f
C10303 FILLER_0_17_72/a_1468_375# _131_ 0.006871f
C10304 ctln[1] clk 0.551557f
C10305 vss _145_ 0.399701f
C10306 _105_ _295_/a_36_472# 0.031356f
C10307 ctlp[2] _420_/a_2248_156# 0.001156f
C10308 _036_ net69 0.353233f
C10309 FILLER_0_13_80/a_124_375# vdd 0.018971f
C10310 FILLER_0_5_72/a_36_472# net47 0.003953f
C10311 net50 trim_val\[0\] 0.390586f
C10312 _053_ _376_/a_36_160# 0.005109f
C10313 mask\[4\] output34/a_224_472# 0.001777f
C10314 FILLER_0_18_107/a_2364_375# _022_ 0.001902f
C10315 trimb[3] net43 0.221036f
C10316 FILLER_0_14_181/a_124_375# _137_ 0.006021f
C10317 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_36_472# 0.007947f
C10318 _448_/a_2248_156# trim_val\[4\] 0.001534f
C10319 FILLER_0_2_177/a_484_472# net22 0.001324f
C10320 _161_ _061_ 0.026347f
C10321 _337_/a_257_69# vdd 0.002972f
C10322 _369_/a_36_68# _367_/a_36_68# 0.038188f
C10323 FILLER_0_24_130/a_124_375# output23/a_224_472# 0.006051f
C10324 FILLER_0_9_223/a_572_375# state\[0\] 0.079258f
C10325 _428_/a_448_472# _095_ 0.008804f
C10326 _315_/a_244_497# vss 0.008724f
C10327 _274_/a_36_68# _070_ 0.032424f
C10328 _039_ clkc 0.003104f
C10329 net33 _048_ 0.017633f
C10330 _352_/a_49_472# FILLER_0_22_128/a_36_472# 0.063744f
C10331 mask\[7\] FILLER_0_22_128/a_572_375# 0.01909f
C10332 _057_ _311_/a_692_473# 0.002083f
C10333 net52 _038_ 0.001152f
C10334 net46 vdd 0.255965f
C10335 FILLER_0_20_193/a_484_472# net21 0.00371f
C10336 FILLER_0_5_198/a_124_375# vdd 0.010749f
C10337 net47 _221_/a_36_160# 0.012197f
C10338 FILLER_0_7_59/a_484_472# vss 0.005804f
C10339 _384_/a_224_472# _160_ 0.00324f
C10340 net2 net59 0.334636f
C10341 net55 FILLER_0_21_28/a_2812_375# 0.004005f
C10342 net41 _217_/a_36_160# 0.004517f
C10343 _412_/a_448_472# net81 0.047334f
C10344 _017_ _131_ 0.005879f
C10345 net80 FILLER_0_22_177/a_572_375# 0.005202f
C10346 FILLER_0_11_142/a_124_375# net23 0.002992f
C10347 net35 FILLER_0_22_128/a_36_472# 0.00784f
C10348 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_124_375# 0.012001f
C10349 net30 result[3] 0.002746f
C10350 net36 _451_/a_448_472# 0.042223f
C10351 _114_ FILLER_0_12_136/a_932_472# 0.003953f
C10352 net2 net4 0.854661f
C10353 _238_/a_67_603# net14 0.004718f
C10354 _395_/a_1044_488# _071_ 0.001198f
C10355 net31 _105_ 0.054065f
C10356 trimb[4] net44 0.127019f
C10357 net68 FILLER_0_6_47/a_1468_375# 0.022624f
C10358 _025_ net71 0.030824f
C10359 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_572_375# 0.007947f
C10360 _013_ _424_/a_796_472# 0.032857f
C10361 net41 _035_ 0.048883f
C10362 FILLER_0_9_72/a_1468_375# _439_/a_36_151# 0.005577f
C10363 net20 _006_ 0.014721f
C10364 _294_/a_224_472# mask\[3\] 0.00233f
C10365 trim_mask\[1\] FILLER_0_6_47/a_2364_375# 0.007169f
C10366 net67 _043_ 0.003726f
C10367 _098_ _205_/a_36_160# 0.033853f
C10368 FILLER_0_3_142/a_36_472# vdd 0.10948f
C10369 FILLER_0_3_142/a_124_375# vss 0.008128f
C10370 _114_ _017_ 0.071595f
C10371 net63 FILLER_0_22_177/a_1468_375# 0.005028f
C10372 _074_ _251_/a_468_472# 0.001217f
C10373 FILLER_0_0_96/a_36_472# net14 0.009584f
C10374 net23 _066_ 0.031928f
C10375 _128_ _055_ 1.887595f
C10376 cal_itt\[3\] _087_ 0.002881f
C10377 FILLER_0_22_128/a_932_472# vdd 0.004405f
C10378 FILLER_0_22_128/a_484_472# vss 0.002338f
C10379 FILLER_0_16_89/a_572_375# _451_/a_448_472# 0.001597f
C10380 _033_ _160_ 0.020281f
C10381 FILLER_0_16_73/a_124_375# _176_ 0.006386f
C10382 _077_ FILLER_0_8_239/a_36_472# 0.001289f
C10383 FILLER_0_9_28/a_1916_375# _042_ 0.002352f
C10384 FILLER_0_9_28/a_1468_375# net51 0.00111f
C10385 net54 _438_/a_2665_112# 0.032855f
C10386 _030_ _384_/a_224_472# 0.003019f
C10387 net65 fanout64/a_36_160# 0.214347f
C10388 FILLER_0_7_59/a_572_375# net15 0.033245f
C10389 FILLER_0_15_282/a_572_375# net62 0.007699f
C10390 net79 vdd 1.283563f
C10391 FILLER_0_7_146/a_36_472# vdd 0.072981f
C10392 FILLER_0_7_146/a_124_375# vss 0.050543f
C10393 net26 FILLER_0_23_44/a_572_375# 0.003172f
C10394 net20 FILLER_0_15_228/a_36_472# 0.020589f
C10395 FILLER_0_16_57/a_124_375# FILLER_0_17_56/a_124_375# 0.026339f
C10396 trim[0] trim[2] 0.002289f
C10397 net16 _167_ 0.001124f
C10398 fanout67/a_36_160# _439_/a_36_151# 0.00246f
C10399 _114_ _250_/a_36_68# 0.017773f
C10400 net22 FILLER_0_18_209/a_572_375# 0.005202f
C10401 vdd trim[3] 0.147228f
C10402 net65 _413_/a_1204_472# 0.017514f
C10403 _165_ _220_/a_67_603# 0.004199f
C10404 _059_ _227_/a_36_160# 0.099735f
C10405 FILLER_0_10_78/a_36_472# vdd 0.001865f
C10406 FILLER_0_10_78/a_1468_375# vss 0.054053f
C10407 _153_ _157_ 0.050552f
C10408 _428_/a_2248_156# net53 0.001188f
C10409 FILLER_0_15_142/a_124_375# _136_ 0.001706f
C10410 _104_ _420_/a_2560_156# 0.002734f
C10411 _413_/a_1308_423# net21 0.065716f
C10412 FILLER_0_21_28/a_36_472# net40 0.032105f
C10413 _274_/a_244_497# net64 0.004085f
C10414 net64 _099_ 0.007017f
C10415 ctln[1] net65 0.073241f
C10416 net23 net37 0.01763f
C10417 _086_ _311_/a_66_473# 0.007295f
C10418 FILLER_0_18_2/a_1380_472# net38 0.029747f
C10419 _069_ _070_ 0.257147f
C10420 mask\[4\] net21 0.049513f
C10421 FILLER_0_5_54/a_484_472# net47 0.006652f
C10422 ctln[2] net5 0.001249f
C10423 FILLER_0_4_99/a_36_472# FILLER_0_4_107/a_36_472# 0.002296f
C10424 output38/a_224_472# _445_/a_36_151# 0.199812f
C10425 _099_ mask\[1\] 0.19135f
C10426 _097_ FILLER_0_15_180/a_124_375# 0.007065f
C10427 _242_/a_36_160# net47 0.028264f
C10428 FILLER_0_9_72/a_1380_472# vss 0.007254f
C10429 FILLER_0_12_124/a_36_472# _131_ 0.028609f
C10430 net82 FILLER_0_3_172/a_484_472# 0.008052f
C10431 _360_/a_36_160# _133_ 0.001878f
C10432 _142_ _141_ 0.200324f
C10433 net75 FILLER_0_6_239/a_124_375# 0.013962f
C10434 state\[0\] _055_ 0.042917f
C10435 net78 mask\[7\] 0.001437f
C10436 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1468_375# 0.016748f
C10437 _173_ net51 0.016607f
C10438 net60 mask\[7\] 0.001053f
C10439 vdd FILLER_0_22_107/a_124_375# 0.029828f
C10440 _094_ _418_/a_1308_423# 0.029276f
C10441 _119_ _374_/a_36_68# 0.001756f
C10442 _086_ _374_/a_244_472# 0.001496f
C10443 _137_ FILLER_0_16_154/a_932_472# 0.004753f
C10444 _320_/a_36_472# mask\[0\] 0.001026f
C10445 _028_ FILLER_0_7_72/a_3260_375# 0.003505f
C10446 _062_ _160_ 0.001024f
C10447 net75 net27 0.037524f
C10448 net58 output27/a_224_472# 0.121438f
C10449 _141_ net35 0.003655f
C10450 mask\[4\] FILLER_0_20_177/a_484_472# 0.001215f
C10451 _253_/a_672_68# _074_ 0.001857f
C10452 net43 FILLER_0_20_15/a_36_472# 0.002803f
C10453 fanout52/a_36_160# vss 0.010082f
C10454 _114_ FILLER_0_12_124/a_36_472# 0.003953f
C10455 _119_ FILLER_0_8_127/a_36_472# 0.053962f
C10456 _144_ _434_/a_36_151# 0.004055f
C10457 _376_/a_36_160# _164_ 0.004503f
C10458 output27/a_224_472# _425_/a_2665_112# 0.021504f
C10459 FILLER_0_15_282/a_36_472# net30 0.001692f
C10460 FILLER_0_15_282/a_124_375# result[3] 0.004601f
C10461 net24 vss 0.172755f
C10462 FILLER_0_18_107/a_36_472# FILLER_0_17_104/a_484_472# 0.026657f
C10463 _432_/a_448_472# _136_ 0.001892f
C10464 _119_ FILLER_0_7_162/a_124_375# 0.059009f
C10465 _131_ FILLER_0_11_109/a_124_375# 0.001048f
C10466 FILLER_0_12_136/a_932_472# _126_ 0.014483f
C10467 _086_ _331_/a_244_472# 0.001991f
C10468 _038_ _172_ 0.050158f
C10469 _053_ FILLER_0_7_72/a_1468_375# 0.014569f
C10470 calibrate FILLER_0_8_156/a_36_472# 0.001283f
C10471 _122_ FILLER_0_8_156/a_572_375# 0.002572f
C10472 net61 net33 0.043271f
C10473 FILLER_0_20_15/a_1020_375# vdd 0.005198f
C10474 mask\[4\] FILLER_0_18_177/a_124_375# 0.016093f
C10475 _069_ FILLER_0_9_142/a_36_472# 0.035528f
C10476 output34/a_224_472# net34 0.031833f
C10477 _000_ FILLER_0_3_221/a_1020_375# 0.016709f
C10478 net82 cal_itt\[0\] 0.063072f
C10479 net29 _417_/a_2665_112# 0.002977f
C10480 FILLER_0_14_181/a_36_472# _113_ 0.004214f
C10481 _111_ _098_ 0.014998f
C10482 _126_ _017_ 0.071134f
C10483 FILLER_0_17_72/a_1828_472# net36 0.028046f
C10484 _099_ vss 0.255039f
C10485 _431_/a_36_151# _334_/a_36_160# 0.032942f
C10486 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_572_375# 0.026339f
C10487 _132_ FILLER_0_14_107/a_484_472# 0.005391f
C10488 _421_/a_2248_156# _109_ 0.001349f
C10489 trim_mask\[2\] FILLER_0_3_78/a_572_375# 0.011713f
C10490 _131_ FILLER_0_14_107/a_1468_375# 0.051201f
C10491 _114_ FILLER_0_11_109/a_124_375# 0.009676f
C10492 _292_/a_36_160# vdd 0.01694f
C10493 fanout59/a_36_160# net18 0.003981f
C10494 net81 FILLER_0_15_235/a_124_375# 0.008139f
C10495 _281_/a_672_472# _097_ 0.002131f
C10496 _411_/a_2248_156# cal_itt\[0\] 0.006897f
C10497 _075_ _070_ 0.009314f
C10498 _422_/a_448_472# _109_ 0.006344f
C10499 FILLER_0_6_90/a_484_472# vss 0.00243f
C10500 _128_ _315_/a_36_68# 0.04902f
C10501 _428_/a_1308_423# vdd 0.004352f
C10502 net29 _045_ 0.344478f
C10503 FILLER_0_15_142/a_572_375# net53 0.021481f
C10504 mask\[7\] _433_/a_36_151# 0.001832f
C10505 _260_/a_36_68# _080_ 0.001888f
C10506 mask\[4\] FILLER_0_19_171/a_1380_472# 0.002581f
C10507 trim_val\[4\] _066_ 0.015621f
C10508 ctln[2] FILLER_0_1_266/a_572_375# 0.012126f
C10509 _430_/a_1000_472# net22 0.032221f
C10510 net20 net76 0.021613f
C10511 net58 net81 0.375649f
C10512 _126_ _250_/a_36_68# 0.022134f
C10513 net57 FILLER_0_3_172/a_36_472# 0.001007f
C10514 net57 _386_/a_124_24# 0.037058f
C10515 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_124_375# 0.026339f
C10516 _061_ FILLER_0_8_156/a_572_375# 0.023346f
C10517 FILLER_0_15_72/a_124_375# vdd 0.020511f
C10518 net37 FILLER_0_6_231/a_572_375# 0.001989f
C10519 fanout63/a_36_160# vdd 0.020165f
C10520 _428_/a_448_472# net74 0.019814f
C10521 mask\[7\] _147_ 0.295801f
C10522 FILLER_0_15_116/a_484_472# net70 0.049569f
C10523 _176_ _095_ 0.064978f
C10524 FILLER_0_15_116/a_124_375# net53 0.009286f
C10525 net81 _425_/a_2665_112# 0.010188f
C10526 net29 _192_/a_67_603# 0.017997f
C10527 _377_/a_36_472# trim_mask\[1\] 0.001763f
C10528 _123_ FILLER_0_7_233/a_124_375# 0.007717f
C10529 FILLER_0_22_177/a_124_375# _434_/a_1308_423# 0.001064f
C10530 net33 _108_ 0.001901f
C10531 _306_/a_36_68# _095_ 0.001366f
C10532 vss _202_/a_36_160# 0.010418f
C10533 _443_/a_1308_423# vdd 0.00203f
C10534 _443_/a_448_472# vss 0.030448f
C10535 FILLER_0_14_99/a_124_375# _451_/a_1040_527# 0.010005f
C10536 _422_/a_36_151# _421_/a_2665_112# 0.001725f
C10537 _065_ ctln[9] 0.123393f
C10538 net55 _423_/a_448_472# 0.00206f
C10539 net41 net16 2.918931f
C10540 net82 FILLER_0_2_171/a_36_472# 0.001777f
C10541 FILLER_0_7_72/a_1916_375# net52 0.001608f
C10542 FILLER_0_7_72/a_1020_375# net50 0.014749f
C10543 vss _433_/a_2560_156# 0.003477f
C10544 output23/a_224_472# vss 0.075684f
C10545 _449_/a_2665_112# _176_ 0.048319f
C10546 result[9] net18 0.019413f
C10547 ctlp[5] vss 0.032166f
C10548 net27 _426_/a_36_151# 0.008613f
C10549 trim_val\[4\] net37 0.003661f
C10550 output22/a_224_472# _435_/a_36_151# 0.12978f
C10551 _136_ _438_/a_36_151# 0.030558f
C10552 _431_/a_36_151# net36 0.006618f
C10553 net50 FILLER_0_2_93/a_36_472# 0.008147f
C10554 net56 FILLER_0_16_154/a_932_472# 0.001401f
C10555 _062_ _117_ 0.042699f
C10556 FILLER_0_17_200/a_572_375# FILLER_0_18_177/a_3172_472# 0.001597f
C10557 FILLER_0_12_124/a_36_472# _126_ 0.056268f
C10558 net52 _448_/a_2665_112# 0.039348f
C10559 FILLER_0_1_212/a_124_375# vdd 0.020159f
C10560 FILLER_0_7_59/a_124_375# fanout67/a_36_160# 0.001597f
C10561 _134_ _120_ 0.047627f
C10562 fanout57/a_36_113# trim_mask\[4\] 0.002404f
C10563 output21/a_224_472# vdd 0.028725f
C10564 net16 FILLER_0_18_37/a_572_375# 0.03477f
C10565 _065_ vss 0.230397f
C10566 _397_/a_36_472# vdd 0.094023f
C10567 FILLER_0_2_177/a_572_375# vss 0.008507f
C10568 FILLER_0_2_177/a_36_472# vdd 0.110255f
C10569 net34 net21 0.036237f
C10570 _417_/a_2560_156# net62 0.003361f
C10571 FILLER_0_17_218/a_36_472# vss 0.006061f
C10572 FILLER_0_17_218/a_484_472# vdd 0.004777f
C10573 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001597f
C10574 FILLER_0_18_2/a_1380_472# net55 0.007469f
C10575 FILLER_0_5_88/a_124_375# vss 0.015423f
C10576 FILLER_0_5_88/a_36_472# vdd 0.090268f
C10577 net71 FILLER_0_22_107/a_36_472# 0.034505f
C10578 output29/a_224_472# vdd 0.103437f
C10579 FILLER_0_5_206/a_124_375# net59 0.008027f
C10580 ctlp[1] _419_/a_36_151# 0.015335f
C10581 _356_/a_36_472# _438_/a_36_151# 0.004432f
C10582 cal_itt\[3\] vdd 0.571239f
C10583 _412_/a_36_151# vdd 0.080326f
C10584 FILLER_0_14_181/a_124_375# _095_ 0.005538f
C10585 FILLER_0_24_63/a_36_472# vss 0.008178f
C10586 _293_/a_36_472# mask\[4\] 0.023203f
C10587 net46 FILLER_0_21_28/a_36_472# 0.051176f
C10588 result[4] _006_ 0.271278f
C10589 _441_/a_36_151# _160_ 0.030777f
C10590 _414_/a_1000_472# _074_ 0.00222f
C10591 net54 FILLER_0_21_150/a_36_472# 0.005439f
C10592 _433_/a_448_472# _145_ 0.045046f
C10593 FILLER_0_18_37/a_124_375# vdd 0.024546f
C10594 _431_/a_36_151# FILLER_0_14_123/a_124_375# 0.002807f
C10595 net79 FILLER_0_12_236/a_572_375# 0.010684f
C10596 FILLER_0_21_286/a_36_472# vdd 0.008714f
C10597 FILLER_0_21_286/a_572_375# vss 0.031895f
C10598 _093_ FILLER_0_21_60/a_484_472# 0.001396f
C10599 FILLER_0_4_144/a_36_472# net47 0.008498f
C10600 _126_ FILLER_0_11_135/a_124_375# 0.008245f
C10601 FILLER_0_5_198/a_36_472# net37 0.0114f
C10602 _130_ FILLER_0_11_135/a_124_375# 0.001198f
C10603 output11/a_224_472# net59 0.002364f
C10604 FILLER_0_7_72/a_1468_375# _164_ 0.003223f
C10605 _028_ _086_ 0.011526f
C10606 _091_ FILLER_0_19_171/a_1468_375# 0.002731f
C10607 _394_/a_1936_472# vss 0.006085f
C10608 _163_ net14 0.040169f
C10609 net23 net13 0.018808f
C10610 _413_/a_36_151# FILLER_0_3_172/a_2364_375# 0.059049f
C10611 _079_ _082_ 0.709481f
C10612 FILLER_0_2_93/a_36_472# trim_mask\[3\] 0.003417f
C10613 net78 net79 0.009641f
C10614 net60 net79 0.113281f
C10615 _131_ FILLER_0_16_115/a_124_375# 0.016715f
C10616 cal_count\[2\] _402_/a_728_93# 0.036871f
C10617 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_124_375# 0.012001f
C10618 _134_ FILLER_0_9_105/a_572_375# 0.02163f
C10619 _448_/a_2665_112# _387_/a_36_113# 0.010064f
C10620 _448_/a_1308_423# _037_ 0.034533f
C10621 FILLER_0_10_28/a_124_375# vdd 0.039012f
C10622 _436_/a_36_151# mask\[7\] 0.030028f
C10623 trim[0] _446_/a_36_151# 0.044586f
C10624 net38 _446_/a_1308_423# 0.010331f
C10625 _077_ FILLER_0_9_60/a_36_472# 0.038809f
C10626 _033_ net67 0.148585f
C10627 _328_/a_36_113# cal_count\[3\] 0.006392f
C10628 _012_ FILLER_0_23_44/a_932_472# 0.001572f
C10629 _053_ FILLER_0_6_47/a_2276_472# 0.004472f
C10630 _436_/a_36_151# _148_ 0.032004f
C10631 _436_/a_2665_112# net35 0.012468f
C10632 _441_/a_36_151# _030_ 0.005324f
C10633 result[7] _419_/a_1308_423# 0.015718f
C10634 output34/a_224_472# _419_/a_2665_112# 0.010731f
C10635 FILLER_0_16_89/a_36_472# vss 0.001289f
C10636 net44 vss 0.477283f
C10637 output39/a_224_472# _034_ 0.002236f
C10638 _257_/a_36_472# vss 0.023401f
C10639 _398_/a_36_113# net17 0.002702f
C10640 input2/a_36_113# clk 0.021981f
C10641 _335_/a_49_472# mask\[1\] 0.032497f
C10642 _028_ _154_ 0.174927f
C10643 vss _107_ 0.186994f
C10644 _189_/a_67_603# FILLER_0_14_235/a_36_472# 0.002778f
C10645 mask\[0\] FILLER_0_12_220/a_1468_375# 0.001484f
C10646 _171_ vss 0.004501f
C10647 _072_ state\[2\] 0.002629f
C10648 _412_/a_2560_156# net5 0.007446f
C10649 _430_/a_2665_112# _091_ 0.016404f
C10650 _098_ _047_ 0.062495f
C10651 FILLER_0_19_134/a_36_472# _145_ 0.080913f
C10652 FILLER_0_14_91/a_124_375# _177_ 0.00134f
C10653 FILLER_0_21_142/a_36_472# net54 0.02217f
C10654 net49 _440_/a_796_472# 0.003597f
C10655 FILLER_0_18_209/a_124_375# vdd 0.023676f
C10656 net7 net16 0.033509f
C10657 FILLER_0_15_116/a_572_375# FILLER_0_14_107/a_1468_375# 0.026339f
C10658 FILLER_0_15_116/a_36_472# FILLER_0_14_107/a_1020_375# 0.001723f
C10659 ctln[1] FILLER_0_3_221/a_1468_375# 0.001235f
C10660 _394_/a_1936_472# cal_count\[1\] 0.008364f
C10661 _394_/a_718_524# net15 0.027444f
C10662 output32/a_224_472# _418_/a_448_472# 0.008149f
C10663 net68 _440_/a_796_472# 0.021463f
C10664 net20 _083_ 0.230786f
C10665 result[5] _419_/a_448_472# 0.00232f
C10666 _032_ net69 0.347645f
C10667 _431_/a_36_151# _020_ 0.023081f
C10668 net57 FILLER_0_2_165/a_124_375# 0.007153f
C10669 ctlp[2] vdd 0.617599f
C10670 _415_/a_2248_156# net27 0.022666f
C10671 FILLER_0_22_128/a_932_472# _433_/a_36_151# 0.002841f
C10672 FILLER_0_7_104/a_1020_375# _062_ 0.003073f
C10673 trimb[1] FILLER_0_20_2/a_572_375# 0.003431f
C10674 result[9] net62 0.339372f
C10675 _122_ net23 0.276617f
C10676 _079_ _265_/a_244_68# 0.021777f
C10677 _427_/a_36_151# FILLER_0_14_123/a_36_472# 0.004032f
C10678 _261_/a_36_160# _059_ 0.004993f
C10679 FILLER_0_17_200/a_572_375# mask\[3\] 0.013879f
C10680 FILLER_0_14_81/a_124_375# _176_ 0.001549f
C10681 _087_ _081_ 0.002169f
C10682 FILLER_0_17_104/a_572_375# vdd 0.03661f
C10683 result[2] net19 0.065763f
C10684 net55 FILLER_0_17_56/a_572_375# 0.020564f
C10685 FILLER_0_5_128/a_124_375# _360_/a_36_160# 0.005705f
C10686 _057_ cal_itt\[3\] 0.014849f
C10687 FILLER_0_14_91/a_36_472# _043_ 0.001779f
C10688 _176_ vss 0.761803f
C10689 FILLER_0_5_164/a_572_375# vss 0.055055f
C10690 FILLER_0_5_164/a_36_472# vdd 0.004144f
C10691 _079_ _112_ 0.004464f
C10692 FILLER_0_5_148/a_36_472# _160_ 0.001025f
C10693 _306_/a_36_68# vss 0.008326f
C10694 FILLER_0_14_181/a_124_375# mask\[1\] 0.044784f
C10695 _413_/a_36_151# _002_ 0.0076f
C10696 net39 _445_/a_796_472# 0.002296f
C10697 net23 _049_ 0.215528f
C10698 _429_/a_36_151# FILLER_0_15_205/a_124_375# 0.059049f
C10699 _220_/a_67_603# vss 0.001485f
C10700 _077_ _162_ 0.013298f
C10701 net47 _450_/a_2225_156# 0.057106f
C10702 _008_ _418_/a_2665_112# 0.010862f
C10703 _103_ _099_ 0.025799f
C10704 net29 _287_/a_36_472# 0.002936f
C10705 fanout54/a_36_160# net23 0.05522f
C10706 FILLER_0_11_101/a_484_472# _070_ 0.017841f
C10707 net52 FILLER_0_6_47/a_2724_472# 0.011079f
C10708 _274_/a_1164_497# state\[0\] 0.002914f
C10709 _070_ _090_ 0.369847f
C10710 net24 _211_/a_36_160# 0.021941f
C10711 _073_ net76 0.040554f
C10712 _074_ net47 0.012724f
C10713 _053_ net37 0.080949f
C10714 FILLER_0_12_220/a_484_472# _060_ 0.003379f
C10715 _176_ net74 0.067915f
C10716 FILLER_0_16_107/a_124_375# FILLER_0_18_107/a_36_472# 0.001512f
C10717 net18 FILLER_0_13_290/a_124_375# 0.007717f
C10718 _412_/a_36_151# net2 0.003823f
C10719 FILLER_0_13_228/a_36_472# net79 0.006824f
C10720 ctlp[1] _421_/a_2560_156# 0.001062f
C10721 _251_/a_1130_472# vss 0.001211f
C10722 state\[2\] FILLER_0_13_142/a_1468_375# 0.018691f
C10723 net81 _136_ 0.021146f
C10724 net53 FILLER_0_13_142/a_484_472# 0.059444f
C10725 net3 FILLER_0_15_10/a_124_375# 0.035504f
C10726 result[7] _420_/a_2560_156# 0.001179f
C10727 net55 _041_ 0.972122f
C10728 _446_/a_2560_156# net17 0.00101f
C10729 net65 net19 0.044106f
C10730 _270_/a_36_472# _087_ 0.02676f
C10731 _036_ vss 0.161195f
C10732 _131_ _451_/a_2225_156# 0.008232f
C10733 _445_/a_2560_156# vdd 0.002586f
C10734 _445_/a_2665_112# vss 0.004455f
C10735 net54 FILLER_0_19_142/a_36_472# 0.07544f
C10736 FILLER_0_8_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001597f
C10737 _303_/a_36_472# net36 0.006675f
C10738 _176_ cal_count\[1\] 0.297763f
C10739 _163_ FILLER_0_5_136/a_124_375# 0.009765f
C10740 _070_ net22 0.032551f
C10741 trim_mask\[0\] vdd 0.154098f
C10742 _102_ net36 0.003446f
C10743 _076_ _152_ 0.063574f
C10744 _068_ _081_ 0.006663f
C10745 input5/a_36_113# rstn 0.019149f
C10746 _000_ vdd 0.215988f
C10747 mask\[4\] _201_/a_255_603# 0.002111f
C10748 FILLER_0_6_90/a_572_375# _163_ 0.007844f
C10749 net73 FILLER_0_18_107/a_2364_375# 0.015484f
C10750 _091_ _113_ 0.006236f
C10751 FILLER_0_2_93/a_124_375# net69 0.015032f
C10752 _408_/a_718_524# net17 0.012884f
C10753 FILLER_0_18_177/a_1020_375# FILLER_0_20_177/a_932_472# 0.0027f
C10754 FILLER_0_14_181/a_36_472# vdd 0.027265f
C10755 FILLER_0_14_181/a_124_375# vss 0.009291f
C10756 _430_/a_1308_423# vss 0.003054f
C10757 _425_/a_2248_156# vdd 0.010067f
C10758 net63 _429_/a_36_151# 0.0144f
C10759 ctlp[4] _009_ 0.004522f
C10760 _161_ _267_/a_36_472# 0.043279f
C10761 net17 _054_ 0.034759f
C10762 net15 net49 0.057277f
C10763 FILLER_0_12_2/a_124_375# _450_/a_36_151# 0.001543f
C10764 net80 _024_ 0.064854f
C10765 net32 _204_/a_67_603# 0.037639f
C10766 cal_count\[2\] net17 0.074204f
C10767 _122_ FILLER_0_6_231/a_572_375# 0.016091f
C10768 net68 net15 0.205016f
C10769 result[7] _421_/a_1456_156# 0.001009f
C10770 FILLER_0_8_24/a_36_472# net17 0.045619f
C10771 _136_ _038_ 0.061274f
C10772 FILLER_0_4_177/a_124_375# net37 0.00459f
C10773 _426_/a_448_472# net64 0.054931f
C10774 net61 net18 0.71051f
C10775 net34 _422_/a_2665_112# 0.006103f
C10776 _420_/a_1308_423# vdd 0.00284f
C10777 _420_/a_448_472# vss 0.007371f
C10778 vdd _450_/a_36_151# 0.08588f
C10779 _063_ _167_ 0.002201f
C10780 net70 _451_/a_36_151# 0.04524f
C10781 _320_/a_1120_472# vdd 0.001676f
C10782 _414_/a_2665_112# _068_ 0.002324f
C10783 FILLER_0_16_57/a_572_375# FILLER_0_18_61/a_36_472# 0.001512f
C10784 _098_ FILLER_0_15_180/a_36_472# 0.101593f
C10785 _415_/a_1000_472# _004_ 0.005004f
C10786 net33 _435_/a_2665_112# 0.005831f
C10787 _013_ FILLER_0_18_37/a_1020_375# 0.023067f
C10788 net19 _419_/a_448_472# 0.037199f
C10789 output20/a_224_472# _422_/a_36_151# 0.053592f
C10790 FILLER_0_10_78/a_1468_375# _389_/a_36_148# 0.001699f
C10791 FILLER_0_21_125/a_36_472# vdd 0.007233f
C10792 FILLER_0_21_125/a_572_375# vss 0.054783f
C10793 net28 net79 0.116857f
C10794 _003_ _079_ 0.035497f
C10795 _089_ _088_ 0.009863f
C10796 _038_ _070_ 0.075667f
C10797 _449_/a_796_472# _038_ 0.018626f
C10798 mask\[9\] _354_/a_49_472# 0.032687f
C10799 FILLER_0_13_142/a_572_375# vdd 0.017472f
C10800 FILLER_0_16_57/a_36_472# _176_ 0.075537f
C10801 FILLER_0_13_142/a_124_375# vss 0.009543f
C10802 output38/a_224_472# FILLER_0_3_2/a_36_472# 0.035046f
C10803 net45 vss 0.028798f
C10804 trimb[0] net43 0.109028f
C10805 _324_/a_224_472# _129_ 0.009728f
C10806 FILLER_0_9_142/a_124_375# _118_ 0.06224f
C10807 net64 FILLER_0_8_239/a_36_472# 0.002666f
C10808 _413_/a_448_472# FILLER_0_1_192/a_36_472# 0.001462f
C10809 _434_/a_2665_112# mask\[6\] 0.026286f
C10810 mask\[4\] FILLER_0_19_187/a_484_472# 0.004669f
C10811 _183_ vss 0.009822f
C10812 _082_ vss 0.053349f
C10813 _056_ _061_ 0.445098f
C10814 net76 net1 0.059026f
C10815 net57 _427_/a_2248_156# 0.002706f
C10816 net79 _416_/a_2248_156# 0.026136f
C10817 FILLER_0_8_247/a_36_472# vss 0.003706f
C10818 FILLER_0_8_247/a_484_472# vdd 0.005485f
C10819 _421_/a_1000_472# vdd 0.006281f
C10820 FILLER_0_7_59/a_124_375# trim_mask\[1\] 0.001548f
C10821 fanout77/a_36_113# vss 0.004099f
C10822 net74 FILLER_0_13_142/a_124_375# 0.002722f
C10823 vss FILLER_0_6_37/a_36_472# 0.006755f
C10824 FILLER_0_10_247/a_124_375# net79 0.00498f
C10825 net23 FILLER_0_22_128/a_2724_472# 0.054521f
C10826 net52 FILLER_0_3_78/a_124_375# 0.017889f
C10827 FILLER_0_4_123/a_36_472# _160_ 0.050308f
C10828 fanout64/a_36_160# net64 0.043709f
C10829 _070_ _076_ 0.198272f
C10830 mask\[3\] net36 0.002974f
C10831 FILLER_0_13_290/a_124_375# net62 0.032026f
C10832 net68 net51 0.008885f
C10833 _426_/a_1308_423# vdd 0.008509f
C10834 FILLER_0_16_107/a_484_472# net70 0.002732f
C10835 net52 FILLER_0_2_101/a_124_375# 0.007787f
C10836 FILLER_0_7_162/a_36_472# net57 0.015199f
C10837 _173_ _067_ 0.011854f
C10838 _430_/a_36_151# FILLER_0_18_177/a_2724_472# 0.001512f
C10839 FILLER_0_16_37/a_36_472# cal_count\[2\] 0.008691f
C10840 _326_/a_36_160# _062_ 0.007797f
C10841 _446_/a_1000_472# net40 0.0368f
C10842 _436_/a_36_151# FILLER_0_22_107/a_124_375# 0.026916f
C10843 _178_ vdd 0.440802f
C10844 FILLER_0_11_101/a_124_375# vdd 0.024363f
C10845 FILLER_0_24_96/a_124_375# output24/a_224_472# 0.00363f
C10846 _064_ _446_/a_448_472# 0.01156f
C10847 _122_ FILLER_0_5_198/a_36_472# 0.00305f
C10848 output47/a_224_472# vdd 0.028666f
C10849 _088_ FILLER_0_4_213/a_124_375# 0.016013f
C10850 _073_ _083_ 0.097365f
C10851 _086_ _085_ 0.374127f
C10852 net65 FILLER_0_3_172/a_484_472# 0.003678f
C10853 net65 _386_/a_848_380# 0.00123f
C10854 net17 FILLER_0_23_44/a_572_375# 0.001332f
C10855 _013_ FILLER_0_18_61/a_36_472# 0.01628f
C10856 net63 _435_/a_1000_472# 0.002536f
C10857 _247_/a_36_160# net21 0.002254f
C10858 _017_ _095_ 0.002789f
C10859 FILLER_0_16_154/a_1380_472# vdd 0.001901f
C10860 FILLER_0_16_154/a_932_472# vss 0.001652f
C10861 _412_/a_2248_156# cal_itt\[1\] 0.005868f
C10862 FILLER_0_3_172/a_2812_375# net21 0.015743f
C10863 FILLER_0_8_239/a_36_472# vss 0.003115f
C10864 _265_/a_244_68# vss 0.009604f
C10865 trim[4] net40 0.017911f
C10866 net73 net70 0.040702f
C10867 fanout70/a_36_113# net53 0.031633f
C10868 _408_/a_1336_472# net40 0.020063f
C10869 net19 _420_/a_2665_112# 0.012322f
C10870 ctln[8] output16/a_224_472# 0.006971f
C10871 sample output27/a_224_472# 0.006116f
C10872 ctln[2] en 0.001355f
C10873 _081_ vdd 0.729534f
C10874 _085_ cal_count\[3\] 0.653405f
C10875 _076_ FILLER_0_9_142/a_36_472# 0.038562f
C10876 _068_ FILLER_0_9_142/a_124_375# 0.008226f
C10877 ctlp[2] net78 0.369805f
C10878 _153_ _160_ 0.304792f
C10879 _093_ _397_/a_36_472# 0.001509f
C10880 fanout75/a_36_113# net37 0.010418f
C10881 _077_ FILLER_0_8_156/a_124_375# 0.00407f
C10882 result[2] _193_/a_36_160# 0.040932f
C10883 _112_ vss 0.145781f
C10884 net16 trim_val\[0\] 0.00463f
C10885 _415_/a_2665_112# net64 0.074373f
C10886 _093_ FILLER_0_17_218/a_484_472# 0.004665f
C10887 result[0] net5 0.001104f
C10888 FILLER_0_21_125/a_484_472# _140_ 0.013936f
C10889 mask\[0\] state\[1\] 0.064758f
C10890 FILLER_0_7_104/a_932_472# vdd 0.020291f
C10891 fanout64/a_36_160# vss 0.007097f
C10892 net61 net62 0.874859f
C10893 net36 _040_ 0.429029f
C10894 _144_ mask\[6\] 0.230129f
C10895 net81 FILLER_0_10_256/a_36_472# 0.089055f
C10896 FILLER_0_14_99/a_124_375# net14 0.04852f
C10897 _436_/a_1204_472# _050_ 0.006724f
C10898 net54 net14 0.121719f
C10899 net68 _381_/a_36_472# 0.003421f
C10900 FILLER_0_2_127/a_124_375# vdd 0.013496f
C10901 FILLER_0_18_107/a_3260_375# vss 0.056926f
C10902 FILLER_0_18_107/a_36_472# vdd 0.116746f
C10903 output15/a_224_472# vss 0.067969f
C10904 _413_/a_2248_156# vdd -0.006767f
C10905 net65 cal_itt\[0\] 0.07564f
C10906 net41 _063_ 0.105528f
C10907 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_36_472# 0.086905f
C10908 _267_/a_36_472# _071_ 0.001682f
C10909 result[6] net77 0.111093f
C10910 FILLER_0_19_195/a_124_375# _202_/a_36_160# 0.005489f
C10911 _161_ _113_ 0.201931f
C10912 FILLER_0_14_107/a_572_375# _451_/a_36_151# 0.02627f
C10913 vdd FILLER_0_10_94/a_572_375# 0.02784f
C10914 _448_/a_1204_472# net22 0.002283f
C10915 FILLER_0_18_139/a_1468_375# _145_ 0.002318f
C10916 mask\[8\] _354_/a_257_69# 0.003809f
C10917 net80 _337_/a_49_472# 0.015686f
C10918 FILLER_0_16_89/a_572_375# _040_ 0.004252f
C10919 net31 _099_ 0.01086f
C10920 _417_/a_36_151# _006_ 0.015561f
C10921 ctln[1] vss 0.27233f
C10922 FILLER_0_21_28/a_1916_375# _012_ 0.023886f
C10923 _270_/a_36_472# vdd 0.09815f
C10924 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_124_375# 0.001597f
C10925 _443_/a_2665_112# FILLER_0_2_165/a_36_472# 0.007491f
C10926 net52 _158_ 0.001338f
C10927 _030_ _153_ 0.026157f
C10928 _421_/a_36_151# net77 0.028951f
C10929 net57 FILLER_0_3_142/a_36_472# 0.002298f
C10930 FILLER_0_16_57/a_36_472# _183_ 0.004107f
C10931 _010_ _419_/a_796_472# 0.001613f
C10932 _187_ _188_ 0.001453f
C10933 FILLER_0_24_274/a_1380_472# vss 0.005744f
C10934 net39 _054_ 0.049797f
C10935 _414_/a_2248_156# vss 0.00384f
C10936 _414_/a_2665_112# vdd 0.006496f
C10937 FILLER_0_11_135/a_36_472# _118_ 0.002496f
C10938 FILLER_0_5_117/a_36_472# _160_ 0.005314f
C10939 _059_ _062_ 0.161331f
C10940 FILLER_0_8_138/a_124_375# calibrate 0.013177f
C10941 FILLER_0_10_78/a_1020_375# _120_ 0.003403f
C10942 _413_/a_36_151# net76 0.084453f
C10943 output37/a_224_472# output48/a_224_472# 0.005147f
C10944 _255_/a_224_552# _090_ 0.001598f
C10945 _149_ FILLER_0_20_98/a_124_375# 0.020028f
C10946 _134_ FILLER_0_10_107/a_484_472# 0.020725f
C10947 _093_ FILLER_0_16_89/a_484_472# 0.001526f
C10948 net72 FILLER_0_17_38/a_124_375# 0.041464f
C10949 FILLER_0_14_181/a_124_375# _097_ 0.001668f
C10950 _053_ _122_ 0.368823f
C10951 _375_/a_36_68# _062_ 0.012855f
C10952 _415_/a_2665_112# vss 0.015461f
C10953 _114_ _055_ 0.071738f
C10954 _144_ mask\[9\] 0.001909f
C10955 ctln[3] FILLER_0_0_266/a_124_375# 0.002726f
C10956 _120_ FILLER_0_9_72/a_932_472# 0.001709f
C10957 _161_ _118_ 0.023939f
C10958 _420_/a_2665_112# _009_ 0.001752f
C10959 FILLER_0_22_177/a_1020_375# mask\[6\] 0.002657f
C10960 _093_ FILLER_0_18_209/a_124_375# 0.00333f
C10961 _414_/a_448_472# net76 0.002346f
C10962 net1 _083_ 0.30074f
C10963 mask\[4\] FILLER_0_19_155/a_572_375# 0.020261f
C10964 _450_/a_1040_527# _039_ 0.015478f
C10965 FILLER_0_16_107/a_484_472# FILLER_0_14_107/a_572_375# 0.001404f
C10966 net65 FILLER_0_2_171/a_36_472# 0.023858f
C10967 _005_ vdd 0.506158f
C10968 net18 _416_/a_1000_472# 0.046085f
C10969 _449_/a_1308_423# vdd 0.002584f
C10970 _449_/a_448_472# vss 0.032274f
C10971 net28 output29/a_224_472# 0.028512f
C10972 net50 _441_/a_2560_156# 0.008865f
C10973 _440_/a_796_472# net47 0.002508f
C10974 _230_/a_244_68# _060_ 0.002039f
C10975 FILLER_0_12_220/a_484_472# vss 0.006724f
C10976 FILLER_0_12_220/a_932_472# vdd 0.003359f
C10977 mask\[8\] FILLER_0_22_86/a_124_375# 0.014263f
C10978 FILLER_0_4_49/a_484_472# net49 0.006499f
C10979 net82 fanout76/a_36_160# 0.001033f
C10980 FILLER_0_5_128/a_572_375# _152_ 0.00813f
C10981 FILLER_0_9_28/a_1020_375# _054_ 0.002273f
C10982 ctlp[6] net23 0.006951f
C10983 net55 FILLER_0_18_37/a_36_472# 0.006084f
C10984 _106_ net63 0.034574f
C10985 FILLER_0_4_107/a_1380_472# _160_ 0.020979f
C10986 net35 _434_/a_2665_112# 0.024254f
C10987 output31/a_224_472# net18 0.009938f
C10988 output32/a_224_472# _006_ 0.001009f
C10989 FILLER_0_17_72/a_1916_375# vdd 0.002595f
C10990 FILLER_0_17_72/a_1468_375# vss 0.003461f
C10991 net52 net82 0.108202f
C10992 _069_ _429_/a_1308_423# 0.027468f
C10993 FILLER_0_4_49/a_484_472# net68 0.027016f
C10994 FILLER_0_16_89/a_124_375# net36 0.011956f
C10995 _093_ FILLER_0_17_104/a_572_375# 0.01418f
C10996 FILLER_0_21_142/a_36_472# FILLER_0_21_133/a_36_472# 0.001963f
C10997 _321_/a_2034_472# _176_ 0.002722f
C10998 _069_ _395_/a_36_488# 0.042974f
C10999 output29/a_224_472# _416_/a_2248_156# 0.024448f
C11000 result[2] _416_/a_448_472# 0.003015f
C11001 net82 _443_/a_796_472# 0.00219f
C11002 _003_ vss 0.095366f
C11003 net50 _439_/a_2665_112# 0.007973f
C11004 trimb[1] FILLER_0_18_2/a_2364_375# 0.001523f
C11005 _095_ FILLER_0_14_107/a_1468_375# 0.010523f
C11006 _105_ _204_/a_67_603# 0.061486f
C11007 _142_ mask\[2\] 0.093231f
C11008 _401_/a_36_68# FILLER_0_15_59/a_36_472# 0.019798f
C11009 FILLER_0_7_72/a_1468_375# _376_/a_36_160# 0.02985f
C11010 _425_/a_2560_156# net37 0.002508f
C11011 FILLER_0_22_86/a_124_375# vss 0.00285f
C11012 FILLER_0_22_86/a_572_375# vdd 0.017472f
C11013 mask\[4\] FILLER_0_18_177/a_3172_472# 0.014657f
C11014 _116_ FILLER_0_12_196/a_36_472# 0.010951f
C11015 result[9] _417_/a_2560_156# 0.00263f
C11016 net38 _450_/a_836_156# 0.0039f
C11017 _143_ _140_ 0.00806f
C11018 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_124_375# 0.026339f
C11019 ctlp[1] vdd 0.942436f
C11020 _140_ _348_/a_49_472# 0.023816f
C11021 _091_ vdd 1.011371f
C11022 _384_/a_224_472# _168_ 0.003461f
C11023 FILLER_0_12_136/a_932_472# vss 0.008682f
C11024 FILLER_0_12_136/a_1380_472# vdd 0.006419f
C11025 mask\[8\] _437_/a_1000_472# 0.00112f
C11026 _422_/a_1000_472# _009_ 0.007191f
C11027 _417_/a_2248_156# vdd 0.004032f
C11028 _086_ _310_/a_49_472# 0.013039f
C11029 FILLER_0_9_142/a_124_375# vdd 0.015952f
C11030 net25 _423_/a_2665_112# 0.007096f
C11031 _389_/a_36_148# _171_ 0.023988f
C11032 net36 FILLER_0_18_76/a_484_472# 0.005765f
C11033 _069_ _228_/a_36_68# 0.001676f
C11034 net23 _170_ 0.107532f
C11035 _178_ cal_count\[0\] 0.011488f
C11036 FILLER_0_17_72/a_572_375# net15 0.003021f
C11037 FILLER_0_15_142/a_572_375# net23 0.006327f
C11038 net53 vdd 0.78288f
C11039 _017_ vss 0.022624f
C11040 _161_ _068_ 0.026092f
C11041 FILLER_0_13_206/a_124_375# _043_ 0.014212f
C11042 net82 FILLER_0_2_177/a_484_472# 0.001777f
C11043 net20 _421_/a_448_472# 0.015767f
C11044 fanout77/a_36_113# _103_ 0.006045f
C11045 cal_count\[3\] _310_/a_49_472# 0.00277f
C11046 net78 _421_/a_1000_472# 0.022212f
C11047 net60 _421_/a_1000_472# 0.035511f
C11048 net70 _427_/a_36_151# 0.029237f
C11049 _131_ _058_ 0.031061f
C11050 FILLER_0_8_138/a_124_375# _125_ 0.001589f
C11051 net57 _428_/a_1308_423# 0.018725f
C11052 _096_ mask\[0\] 0.052773f
C11053 _029_ FILLER_0_5_88/a_124_375# 0.006771f
C11054 net61 _422_/a_448_472# 0.006042f
C11055 _412_/a_448_472# net82 0.030379f
C11056 FILLER_0_4_213/a_36_472# vdd 0.087733f
C11057 FILLER_0_4_213/a_572_375# vss 0.017689f
C11058 _017_ net74 0.041246f
C11059 _109_ _108_ 0.001806f
C11060 _126_ _055_ 0.01647f
C11061 net47 FILLER_0_5_148/a_572_375# 0.062581f
C11062 FILLER_0_9_28/a_124_375# net47 0.006757f
C11063 _144_ _352_/a_49_472# 0.00176f
C11064 _127_ _118_ 0.141388f
C11065 _250_/a_36_68# vss 0.005108f
C11066 _032_ vss 0.02257f
C11067 _236_/a_36_160# net40 0.035082f
C11068 _114_ _058_ 0.013316f
C11069 FILLER_0_10_37/a_36_472# net51 0.002346f
C11070 FILLER_0_4_197/a_124_375# net21 0.018398f
C11071 net55 _012_ 0.060122f
C11072 _214_/a_36_160# _098_ 0.001496f
C11073 net54 _433_/a_2248_156# 0.04755f
C11074 _176_ _389_/a_36_148# 0.060256f
C11075 _144_ net35 0.036236f
C11076 _255_/a_224_552# _076_ 0.081663f
C11077 _446_/a_1000_472# trim[3] 0.001257f
C11078 input1/a_36_113# net18 0.004922f
C11079 FILLER_0_21_125/a_36_472# _433_/a_36_151# 0.001723f
C11080 FILLER_0_11_78/a_124_375# vdd -0.011022f
C11081 _166_ _160_ 0.492224f
C11082 _412_/a_2248_156# net59 0.008792f
C11083 net15 net47 0.035839f
C11084 fanout69/a_36_113# trim_mask\[4\] 0.027938f
C11085 net74 _032_ 0.208799f
C11086 _074_ FILLER_0_7_233/a_124_375# 0.003081f
C11087 ctlp[3] mask\[7\] 0.103955f
C11088 _037_ net59 0.799647f
C11089 FILLER_0_4_177/a_36_472# trim_val\[4\] 0.001889f
C11090 FILLER_0_19_55/a_36_472# net36 0.001068f
C11091 result[5] vss 0.307366f
C11092 output16/a_224_472# vdd 0.006151f
C11093 _077_ FILLER_0_11_64/a_36_472# 0.076102f
C11094 _416_/a_1000_472# net62 0.002399f
C11095 _301_/a_36_472# vdd 0.013061f
C11096 _412_/a_2560_156# en 0.049213f
C11097 FILLER_0_12_50/a_124_375# vdd 0.039185f
C11098 _155_ net14 0.10433f
C11099 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_124_375# 0.012001f
C11100 trim_val\[4\] _443_/a_2248_156# 0.050943f
C11101 _100_ _099_ 0.03589f
C11102 FILLER_0_7_104/a_1020_375# _153_ 0.026997f
C11103 net65 _411_/a_1308_423# 0.004122f
C11104 _028_ FILLER_0_5_72/a_484_472# 0.003042f
C11105 _422_/a_448_472# _108_ 0.03293f
C11106 _115_ net14 0.037635f
C11107 FILLER_0_12_124/a_36_472# vss 0.001443f
C11108 FILLER_0_18_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001684f
C11109 output31/a_224_472# net62 0.030092f
C11110 _370_/a_848_380# FILLER_0_5_136/a_36_472# 0.001177f
C11111 FILLER_0_9_60/a_36_472# vss 0.001327f
C11112 FILLER_0_9_60/a_484_472# vdd 0.005181f
C11113 _077_ _439_/a_1204_472# 0.016471f
C11114 _153_ _156_ 0.539362f
C11115 _053_ _444_/a_2665_112# 0.001698f
C11116 FILLER_0_7_72/a_2724_472# _219_/a_36_160# 0.001448f
C11117 fanout72/a_36_113# vdd -0.002193f
C11118 FILLER_0_13_65/a_124_375# fanout72/a_36_113# 0.005467f
C11119 net15 FILLER_0_23_44/a_1468_375# 0.001307f
C11120 result[9] FILLER_0_23_282/a_36_472# 0.001324f
C11121 output11/a_224_472# _000_ 0.006606f
C11122 FILLER_0_3_172/a_1380_472# net22 0.012284f
C11123 FILLER_0_10_256/a_124_375# vdd 0.041848f
C11124 _074_ FILLER_0_6_177/a_572_375# 0.012642f
C11125 fanout67/a_36_160# net67 0.017633f
C11126 _022_ _145_ 0.199016f
C11127 FILLER_0_23_282/a_124_375# vdd -0.003896f
C11128 mask\[5\] FILLER_0_20_169/a_36_472# 0.016469f
C11129 cal_itt\[3\] net57 0.001586f
C11130 net42 _054_ 0.006314f
C11131 _077_ _055_ 0.083808f
C11132 FILLER_0_12_124/a_36_472# net74 0.021369f
C11133 mask\[4\] mask\[3\] 1.118454f
C11134 _343_/a_665_69# _141_ 0.002451f
C11135 fanout75/a_36_113# _122_ 0.001035f
C11136 _247_/a_36_160# _062_ 0.011327f
C11137 FILLER_0_7_72/a_124_375# vss 0.044754f
C11138 FILLER_0_7_72/a_572_375# vdd 0.004039f
C11139 _075_ calibrate 0.022901f
C11140 _127_ _068_ 0.052712f
C11141 _128_ _070_ 1.279188f
C11142 comp net44 0.079931f
C11143 ctln[3] _411_/a_1204_472# 0.00185f
C11144 FILLER_0_8_24/a_36_472# net42 0.010665f
C11145 _267_/a_36_472# net23 0.001178f
C11146 _445_/a_448_472# _034_ 0.03826f
C11147 net35 FILLER_0_22_177/a_1020_375# 0.008333f
C11148 trim_mask\[1\] _160_ 0.051511f
C11149 FILLER_0_22_86/a_1468_375# net71 0.010224f
C11150 FILLER_0_11_109/a_124_375# vss 0.006764f
C11151 FILLER_0_11_109/a_36_472# vdd 0.109453f
C11152 FILLER_0_2_93/a_572_375# vdd 0.022073f
C11153 _002_ FILLER_0_3_172/a_1916_375# 0.047331f
C11154 FILLER_0_10_78/a_572_375# _115_ 0.004573f
C11155 input5/a_36_113# net59 0.257143f
C11156 _311_/a_66_473# net21 0.02018f
C11157 FILLER_0_11_135/a_36_472# vdd 0.091206f
C11158 FILLER_0_11_135/a_124_375# vss 0.02843f
C11159 _443_/a_36_151# _370_/a_848_380# 0.001568f
C11160 _105_ _201_/a_67_603# 0.003335f
C11161 net47 net51 0.007412f
C11162 net64 net19 0.029763f
C11163 _448_/a_1000_472# vdd 0.004267f
C11164 trim_val\[4\] _170_ 0.281942f
C11165 FILLER_0_11_64/a_36_472# _453_/a_36_151# 0.001723f
C11166 net15 FILLER_0_9_60/a_124_375# 0.003602f
C11167 _327_/a_36_472# _114_ 0.019746f
C11168 FILLER_0_13_212/a_124_375# _043_ 0.011912f
C11169 _095_ _280_/a_224_472# 0.001416f
C11170 input4/a_36_68# net5 0.004765f
C11171 FILLER_0_14_235/a_36_472# net62 0.00534f
C11172 _087_ FILLER_0_3_172/a_932_472# 0.001947f
C11173 ctln[2] cal 0.009784f
C11174 _431_/a_2248_156# _137_ 0.01617f
C11175 FILLER_0_14_107/a_1468_375# vss 0.055167f
C11176 FILLER_0_14_107/a_36_472# vdd 0.114495f
C11177 FILLER_0_22_177/a_1468_375# vss 0.028064f
C11178 FILLER_0_22_177/a_36_472# vdd 0.111906f
C11179 net66 net49 0.657679f
C11180 _077_ _313_/a_67_603# 0.007446f
C11181 _449_/a_36_151# cal_count\[3\] 0.018365f
C11182 net69 _441_/a_2248_156# 0.036635f
C11183 FILLER_0_5_109/a_572_375# vss 0.055343f
C11184 FILLER_0_5_109/a_36_472# vdd 0.042799f
C11185 net68 net66 0.81104f
C11186 cal_itt\[2\] FILLER_0_3_221/a_36_472# 0.003825f
C11187 FILLER_0_5_109/a_124_375# _365_/a_36_68# 0.004633f
C11188 _162_ vss 0.08357f
C11189 _077_ FILLER_0_6_231/a_124_375# 0.009235f
C11190 _161_ vdd 0.262564f
C11191 net71 _437_/a_2665_112# 0.039687f
C11192 net48 _001_ 0.006122f
C11193 _399_/a_224_472# vdd 0.001593f
C11194 net50 _444_/a_2248_156# 0.005539f
C11195 FILLER_0_7_72/a_3172_472# _077_ 0.001923f
C11196 _059_ FILLER_0_5_148/a_36_472# 0.010977f
C11197 _258_/a_36_160# _080_ 0.261387f
C11198 FILLER_0_0_130/a_124_375# net13 0.009149f
C11199 _128_ FILLER_0_9_142/a_36_472# 0.005101f
C11200 net34 FILLER_0_22_128/a_2364_375# 0.009656f
C11201 _436_/a_2248_156# net54 0.043158f
C11202 FILLER_0_9_28/a_3260_375# _077_ 0.01495f
C11203 _016_ _428_/a_36_151# 0.001824f
C11204 result[8] _422_/a_36_151# 0.001488f
C11205 FILLER_0_22_86/a_124_375# _026_ 0.001024f
C11206 _008_ FILLER_0_17_226/a_124_375# 0.006576f
C11207 _137_ FILLER_0_15_180/a_36_472# 0.004437f
C11208 state\[0\] _070_ 0.009608f
C11209 net20 FILLER_0_12_220/a_1468_375# 0.016974f
C11210 net52 FILLER_0_5_72/a_1020_375# 0.00799f
C11211 _436_/a_36_151# FILLER_0_21_125/a_36_472# 0.001695f
C11212 _450_/a_1040_527# clkc 0.001412f
C11213 state\[0\] FILLER_0_12_220/a_1380_472# 0.003733f
C11214 FILLER_0_4_123/a_124_375# net47 0.011322f
C11215 _062_ _134_ 0.024038f
C11216 _285_/a_36_472# vdd 0.073338f
C11217 output48/a_224_472# net48 0.001786f
C11218 _308_/a_124_24# _115_ 0.039354f
C11219 _079_ cal_itt\[0\] 0.018495f
C11220 net58 net82 0.022761f
C11221 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_36_472# 0.001963f
C11222 _205_/a_36_160# vss 0.003612f
C11223 FILLER_0_12_136/a_484_472# cal_count\[3\] 0.007275f
C11224 net16 FILLER_0_12_28/a_124_375# 0.002225f
C11225 result[6] output19/a_224_472# 0.001526f
C11226 output33/a_224_472# ctlp[2] 0.00175f
C11227 _098_ FILLER_0_18_209/a_572_375# 0.001352f
C11228 FILLER_0_21_206/a_36_472# _434_/a_2665_112# 0.00243f
C11229 fanout71/a_36_113# net71 0.087994f
C11230 FILLER_0_18_177/a_3260_375# vdd 0.003399f
C11231 _132_ _428_/a_1204_472# 0.025555f
C11232 _372_/a_1194_69# _163_ 0.001328f
C11233 _085_ _120_ 0.032964f
C11234 _093_ FILLER_0_18_107/a_36_472# 0.008683f
C11235 net19 vss 1.140787f
C11236 _418_/a_2248_156# vdd 0.00423f
C11237 _411_/a_2248_156# net58 0.014884f
C11238 _068_ FILLER_0_8_156/a_572_375# 0.00185f
C11239 _076_ FILLER_0_8_156/a_36_472# 0.006989f
C11240 FILLER_0_9_60/a_124_375# net51 0.002346f
C11241 FILLER_0_9_223/a_572_375# _426_/a_2665_112# 0.005202f
C11242 _155_ FILLER_0_6_90/a_572_375# 0.001562f
C11243 _450_/a_3129_107# net40 0.034729f
C11244 net60 ctlp[1] 0.073021f
C11245 ctlp[1] net78 0.025929f
C11246 FILLER_0_23_88/a_124_375# vss 0.014165f
C11247 FILLER_0_23_88/a_36_472# vdd 0.002576f
C11248 FILLER_0_18_100/a_124_375# mask\[9\] 0.005751f
C11249 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_36_472# 0.086635f
C11250 FILLER_0_5_206/a_124_375# _081_ 0.031751f
C11251 _149_ _437_/a_2248_156# 0.031905f
C11252 _026_ _437_/a_1000_472# 0.042316f
C11253 fanout66/a_36_113# net15 0.024302f
C11254 net67 FILLER_0_12_20/a_36_472# 0.054453f
C11255 _095_ _451_/a_2225_156# 0.001102f
C11256 _440_/a_36_151# FILLER_0_6_47/a_1380_472# 0.001512f
C11257 net57 FILLER_0_5_164/a_36_472# 0.032208f
C11258 _028_ _151_ 0.020076f
C11259 FILLER_0_17_56/a_572_375# FILLER_0_18_61/a_36_472# 0.001597f
C11260 _439_/a_36_151# FILLER_0_6_47/a_2812_375# 0.001512f
C11261 cal_itt\[2\] _088_ 0.010847f
C11262 _077_ _058_ 3.018054f
C11263 _432_/a_448_472# _021_ 0.032563f
C11264 mask\[0\] FILLER_0_13_206/a_36_472# 0.012766f
C11265 FILLER_0_13_142/a_484_472# net23 0.006746f
C11266 input2/a_36_113# vss 0.055539f
C11267 fanout55/a_36_160# _095_ 0.00409f
C11268 _444_/a_2665_112# _164_ 0.015644f
C11269 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_36_472# 0.086635f
C11270 _441_/a_36_151# _168_ 0.033578f
C11271 FILLER_0_13_212/a_932_472# net62 0.059367f
C11272 _063_ trim_val\[0\] 0.001978f
C11273 _095_ _401_/a_36_68# 0.001398f
C11274 _327_/a_36_472# _126_ 0.011444f
C11275 FILLER_0_5_72/a_572_375# _164_ 0.005919f
C11276 _327_/a_36_472# _130_ 0.001474f
C11277 FILLER_0_1_204/a_36_472# net21 0.076466f
C11278 _431_/a_2248_156# net56 0.013627f
C11279 FILLER_0_3_204/a_124_375# net22 0.031438f
C11280 mask\[5\] FILLER_0_20_193/a_484_472# 0.02147f
C11281 _098_ FILLER_0_19_171/a_124_375# 0.040575f
C11282 FILLER_0_3_54/a_36_472# vss 0.002818f
C11283 FILLER_0_9_28/a_3172_472# net68 0.007929f
C11284 _072_ _061_ 0.448032f
C11285 trim_mask\[4\] _066_ 0.396509f
C11286 net15 _453_/a_2665_112# 0.011775f
C11287 output35/a_224_472# mask\[6\] 0.069819f
C11288 _057_ _161_ 1.09228f
C11289 net16 _039_ 0.031852f
C11290 _095_ FILLER_0_13_72/a_36_472# 0.00819f
C11291 _098_ FILLER_0_15_235/a_124_375# 0.012702f
C11292 output44/a_224_472# FILLER_0_20_15/a_484_472# 0.0323f
C11293 net47 _163_ 0.64626f
C11294 _127_ vdd 0.155954f
C11295 _432_/a_36_151# FILLER_0_18_171/a_124_375# 0.001597f
C11296 FILLER_0_12_50/a_124_375# cal_count\[0\] 0.002359f
C11297 _413_/a_448_472# ctln[4] 0.001072f
C11298 FILLER_0_2_111/a_124_375# _369_/a_36_68# 0.001176f
C11299 net81 output28/a_224_472# 0.01335f
C11300 FILLER_0_12_2/a_484_472# net67 0.006435f
C11301 vss FILLER_0_16_115/a_124_375# 0.006358f
C11302 vdd FILLER_0_16_115/a_36_472# 0.093403f
C11303 _389_/a_36_148# FILLER_0_10_94/a_124_375# 0.004673f
C11304 _136_ _139_ 0.394888f
C11305 FILLER_0_6_47/a_1380_472# vdd 0.002735f
C11306 _429_/a_1308_423# net22 0.001856f
C11307 _093_ FILLER_0_17_72/a_1916_375# 0.017467f
C11308 net52 FILLER_0_5_54/a_1468_375# 0.003649f
C11309 _415_/a_2665_112# FILLER_0_9_290/a_36_472# 0.007376f
C11310 result[5] _103_ 0.425479f
C11311 net34 _050_ 0.004662f
C11312 FILLER_0_5_117/a_124_375# net47 0.011773f
C11313 net32 net20 0.006161f
C11314 _009_ vss 0.105833f
C11315 _228_/a_36_68# _090_ 0.018462f
C11316 FILLER_0_4_49/a_484_472# net47 0.002964f
C11317 FILLER_0_18_2/a_36_472# trimb[4] 0.001673f
C11318 net81 _429_/a_1308_423# 0.008913f
C11319 FILLER_0_7_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001723f
C11320 _111_ vss 0.233815f
C11321 FILLER_0_4_197/a_484_472# net22 0.007955f
C11322 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_36_472# 0.086635f
C11323 _098_ FILLER_0_20_98/a_124_375# 0.012779f
C11324 _418_/a_36_151# _007_ 0.007397f
C11325 _077_ FILLER_0_10_78/a_484_472# 0.002486f
C11326 _068_ _246_/a_36_68# 0.059106f
C11327 _274_/a_36_68# _069_ 0.02257f
C11328 _091_ FILLER_0_13_228/a_36_472# 0.001826f
C11329 output27/a_224_472# calibrate 0.010614f
C11330 _422_/a_1204_472# mask\[7\] 0.025592f
C11331 result[9] net61 0.014374f
C11332 _426_/a_2665_112# _055_ 0.00142f
C11333 _449_/a_36_151# _394_/a_1336_472# 0.001582f
C11334 _091_ _093_ 0.035503f
C11335 net52 _443_/a_2665_112# 0.05031f
C11336 _367_/a_244_472# vdd 0.001113f
C11337 FILLER_0_4_144/a_36_472# FILLER_0_3_142/a_124_375# 0.001543f
C11338 _074_ _374_/a_36_68# 0.001447f
C11339 _071_ vdd 0.074299f
C11340 trim[1] _033_ 0.015549f
C11341 cal_count\[2\] FILLER_0_15_2/a_484_472# 0.015036f
C11342 _426_/a_1204_472# calibrate 0.00182f
C11343 fanout78/a_36_113# vss 0.031944f
C11344 fanout60/a_36_160# vss 0.035381f
C11345 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_36_472# 0.002765f
C11346 _228_/a_36_68# net22 0.052558f
C11347 _055_ _060_ 0.181186f
C11348 _273_/a_36_68# vdd 0.041825f
C11349 net27 net4 0.025834f
C11350 net44 _221_/a_36_160# 0.013363f
C11351 _118_ net23 0.108864f
C11352 net82 _152_ 0.001896f
C11353 _453_/a_2665_112# net51 0.046426f
C11354 _174_ FILLER_0_15_59/a_124_375# 0.00622f
C11355 net56 _427_/a_2665_112# 0.012193f
C11356 _363_/a_36_68# FILLER_0_5_109/a_484_472# 0.001709f
C11357 mask\[5\] mask\[4\] 0.176881f
C11358 net57 FILLER_0_13_142/a_572_375# 0.011369f
C11359 FILLER_0_7_162/a_124_375# _074_ 0.007213f
C11360 _415_/a_2248_156# result[1] 0.010922f
C11361 net38 vdd 0.906502f
C11362 _428_/a_36_151# _043_ 0.027757f
C11363 FILLER_0_16_89/a_932_472# _131_ 0.008223f
C11364 _119_ _162_ 0.036701f
C11365 net20 _282_/a_36_160# 0.016884f
C11366 FILLER_0_4_107/a_932_472# net47 0.008252f
C11367 _430_/a_1000_472# net63 0.016386f
C11368 FILLER_0_21_125/a_484_472# _098_ 0.002964f
C11369 FILLER_0_3_221/a_36_472# net59 0.075858f
C11370 FILLER_0_12_20/a_572_375# net47 0.00139f
C11371 FILLER_0_4_197/a_1020_375# _088_ 0.013641f
C11372 FILLER_0_21_28/a_1916_375# vdd -0.009753f
C11373 _052_ _424_/a_448_472# 0.017551f
C11374 FILLER_0_3_172/a_932_472# vdd 0.009887f
C11375 _386_/a_848_380# vss 0.012638f
C11376 _442_/a_36_151# FILLER_0_2_127/a_124_375# 0.001597f
C11377 FILLER_0_9_223/a_36_472# _068_ 0.076678f
C11378 FILLER_0_9_223/a_484_472# _076_ 0.001736f
C11379 net17 output40/a_224_472# 0.00187f
C11380 _449_/a_2248_156# net55 0.052445f
C11381 net4 FILLER_0_3_221/a_36_472# 0.010517f
C11382 vss FILLER_0_8_156/a_124_375# 0.001766f
C11383 vdd FILLER_0_8_156/a_572_375# 0.014611f
C11384 _438_/a_2248_156# net14 0.045909f
C11385 net28 _005_ 0.080653f
C11386 FILLER_0_8_239/a_36_472# _123_ 0.011767f
C11387 ctln[7] vss 0.132613f
C11388 FILLER_0_18_100/a_36_472# vss 0.002412f
C11389 _413_/a_2665_112# net82 0.004306f
C11390 trim_mask\[1\] _156_ 0.007519f
C11391 calibrate net22 0.036525f
C11392 net55 FILLER_0_17_72/a_36_472# 0.020422f
C11393 FILLER_0_18_2/a_1916_375# net17 0.013121f
C11394 net81 FILLER_0_14_235/a_572_375# 0.029643f
C11395 net10 net11 0.007522f
C11396 _064_ _035_ 0.02225f
C11397 _446_/a_2665_112# net49 0.006979f
C11398 _144_ _433_/a_1308_423# 0.027969f
C11399 net18 net8 0.072251f
C11400 _114_ _172_ 0.045798f
C11401 net54 _210_/a_67_603# 0.001108f
C11402 result[9] _108_ 0.015443f
C11403 FILLER_0_5_109/a_124_375# _154_ 0.058658f
C11404 FILLER_0_10_214/a_124_375# vss 0.013034f
C11405 FILLER_0_10_214/a_36_472# vdd 0.026621f
C11406 FILLER_0_20_87/a_124_375# _437_/a_36_151# 0.059049f
C11407 net50 trim_mask\[3\] 0.001654f
C11408 net67 trim_mask\[1\] 0.01761f
C11409 _372_/a_358_69# _160_ 0.001562f
C11410 _005_ _416_/a_2248_156# 0.036714f
C11411 net81 calibrate 0.047274f
C11412 FILLER_0_14_81/a_36_472# _451_/a_3129_107# 0.001557f
C11413 _443_/a_1000_472# _170_ 0.012879f
C11414 _056_ _113_ 0.052362f
C11415 net1 _265_/a_468_472# 0.002612f
C11416 net48 _316_/a_124_24# 0.068708f
C11417 _261_/a_36_160# FILLER_0_5_136/a_36_472# 0.00304f
C11418 net76 FILLER_0_3_172/a_1916_375# 0.019901f
C11419 _131_ FILLER_0_17_104/a_1020_375# 0.006574f
C11420 net36 _437_/a_36_151# 0.002694f
C11421 _451_/a_2225_156# vss 0.003848f
C11422 ctln[1] _411_/a_2560_156# 0.001413f
C11423 fanout58/a_36_160# vss 0.039959f
C11424 cal_itt\[0\] vss 0.11965f
C11425 output48/a_224_472# en 0.003074f
C11426 FILLER_0_21_206/a_124_375# _205_/a_36_160# 0.03126f
C11427 mask\[7\] mask\[6\] 0.227476f
C11428 net65 fanout76/a_36_160# 0.018025f
C11429 fanout55/a_36_160# vss 0.005203f
C11430 net22 _435_/a_2248_156# 0.003453f
C11431 _062_ _311_/a_66_473# 0.027039f
C11432 net57 FILLER_0_16_154/a_1380_472# 0.041458f
C11433 _068_ net23 0.432092f
C11434 _088_ net59 0.270902f
C11435 net38 _452_/a_1040_527# 0.002024f
C11436 _193_/a_36_160# vss 0.035228f
C11437 net57 _081_ 0.023513f
C11438 _431_/a_1000_472# net73 0.035816f
C11439 _177_ net36 0.371814f
C11440 mask\[3\] FILLER_0_18_177/a_1468_375# 0.002924f
C11441 output21/a_224_472# ctlp[3] 0.021951f
C11442 _088_ net4 0.096522f
C11443 _057_ _071_ 0.139904f
C11444 _103_ net19 0.047895f
C11445 _077_ net52 0.047585f
C11446 _103_ _418_/a_1204_472# 0.00582f
C11447 _091_ _429_/a_1204_472# 0.024554f
C11448 fanout55/a_36_160# net74 0.016856f
C11449 FILLER_0_5_212/a_124_375# _078_ 0.002018f
C11450 net60 _418_/a_2248_156# 0.045472f
C11451 net60 _419_/a_3041_156# 0.001022f
C11452 FILLER_0_14_107/a_124_375# _040_ 0.001861f
C11453 _056_ _118_ 0.028015f
C11454 vss FILLER_0_13_72/a_36_472# 0.034188f
C11455 cal_count\[1\] _451_/a_2225_156# 0.006336f
C11456 FILLER_0_13_65/a_36_472# FILLER_0_13_72/a_36_472# 0.002765f
C11457 _095_ _055_ 0.002933f
C11458 _340_/a_36_160# FILLER_0_20_169/a_36_472# 0.195478f
C11459 FILLER_0_24_63/a_124_375# ctlp[8] 0.005758f
C11460 FILLER_0_8_127/a_124_375# _062_ 0.046401f
C11461 _432_/a_1204_472# _091_ 0.00563f
C11462 net65 FILLER_0_1_212/a_36_472# 0.004414f
C11463 output35/a_224_472# net35 0.007217f
C11464 fanout55/a_36_160# cal_count\[1\] 0.007256f
C11465 _233_/a_36_160# vdd 0.064615f
C11466 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_36_472# 0.086635f
C11467 _024_ _023_ 0.005966f
C11468 _408_/a_1936_472# _067_ 0.003007f
C11469 _199_/a_36_160# vdd 0.036579f
C11470 net74 FILLER_0_13_72/a_36_472# 0.007448f
C11471 net65 FILLER_0_2_177/a_484_472# 0.01675f
C11472 FILLER_0_2_171/a_36_472# vss 0.002909f
C11473 net34 output19/a_224_472# 0.122464f
C11474 _246_/a_36_68# vdd 0.047419f
C11475 _127_ FILLER_0_11_142/a_36_472# 0.004538f
C11476 _401_/a_36_68# cal_count\[1\] 0.006747f
C11477 _095_ FILLER_0_15_10/a_124_375# 0.023187f
C11478 _076_ calibrate 1.005804f
C11479 _098_ _348_/a_49_472# 0.011096f
C11480 vss _047_ 0.070755f
C11481 net65 _412_/a_448_472# 0.043862f
C11482 _276_/a_36_160# _106_ 0.009097f
C11483 output14/a_224_472# net14 0.018674f
C11484 mask\[9\] _148_ 0.01635f
C11485 _429_/a_36_151# mask\[1\] 0.001021f
C11486 FILLER_0_4_144/a_484_472# _443_/a_36_151# 0.002841f
C11487 ctln[3] net8 0.003753f
C11488 _126_ _172_ 0.017618f
C11489 FILLER_0_5_109/a_124_375# FILLER_0_4_107/a_484_472# 0.001684f
C11490 net15 FILLER_0_13_72/a_124_375# 0.006403f
C11491 FILLER_0_18_107/a_3172_472# _145_ 0.002415f
C11492 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_572_375# 0.007947f
C11493 _033_ _444_/a_448_472# 0.047424f
C11494 _069_ FILLER_0_18_209/a_484_472# 0.013944f
C11495 _053_ FILLER_0_6_47/a_124_375# 0.002541f
C11496 net66 net47 0.238874f
C11497 _068_ _311_/a_1660_473# 0.003542f
C11498 _104_ FILLER_0_23_274/a_36_472# 0.001642f
C11499 mask\[5\] net34 0.041303f
C11500 _427_/a_2665_112# _095_ 0.039612f
C11501 FILLER_0_5_198/a_484_472# net22 0.012457f
C11502 net27 net79 0.059863f
C11503 _068_ _313_/a_255_603# 0.001149f
C11504 net15 FILLER_0_23_60/a_36_472# 0.004561f
C11505 _136_ _098_ 0.049635f
C11506 FILLER_0_9_223/a_572_375# vss 0.00704f
C11507 FILLER_0_9_223/a_36_472# vdd 0.030289f
C11508 net55 vdd 1.248648f
C11509 FILLER_0_2_165/a_36_472# vss 0.001099f
C11510 _420_/a_36_151# FILLER_0_23_274/a_36_472# 0.001723f
C11511 _080_ FILLER_0_3_221/a_932_472# 0.003217f
C11512 _451_/a_1353_112# net14 0.041814f
C11513 net52 net69 0.372114f
C11514 _305_/a_36_159# _112_ 0.001664f
C11515 _076_ FILLER_0_6_231/a_36_472# 0.005517f
C11516 _369_/a_36_68# vdd 0.042534f
C11517 net82 FILLER_0_4_213/a_484_472# 0.002255f
C11518 _056_ _068_ 0.127175f
C11519 _302_/a_224_472# vss 0.005149f
C11520 net18 _419_/a_36_151# 0.021491f
C11521 _443_/a_448_472# _031_ 0.001143f
C11522 _032_ _442_/a_448_472# 0.001977f
C11523 _443_/a_796_472# net69 0.020234f
C11524 FILLER_0_10_256/a_124_375# net28 0.034928f
C11525 fanout71/a_36_113# FILLER_0_20_107/a_36_472# 0.001645f
C11526 _093_ FILLER_0_18_177/a_3260_375# 0.002695f
C11527 ctlp[3] ctlp[2] 0.006764f
C11528 _280_/a_224_472# _097_ 0.007508f
C11529 ctln[2] fanout81/a_36_160# 0.003798f
C11530 output9/a_224_472# net81 0.02825f
C11531 _086_ FILLER_0_5_181/a_36_472# 0.013437f
C11532 _105_ _291_/a_36_160# 0.002075f
C11533 output39/a_224_472# net40 0.087367f
C11534 vdd _416_/a_1308_423# 0.002623f
C11535 vss _416_/a_448_472# 0.004806f
C11536 output46/a_224_472# net17 0.082914f
C11537 _436_/a_2248_156# FILLER_0_21_133/a_36_472# 0.001148f
C11538 output27/a_224_472# FILLER_0_9_282/a_36_472# 0.001711f
C11539 mask\[0\] _099_ 0.00418f
C11540 ctln[4] net11 0.194506f
C11541 _114_ FILLER_0_13_142/a_1020_375# 0.001964f
C11542 _429_/a_36_151# vss 0.026298f
C11543 _429_/a_448_472# vdd 0.008822f
C11544 _119_ FILLER_0_8_156/a_124_375# 0.025304f
C11545 FILLER_0_4_49/a_572_375# FILLER_0_3_54/a_36_472# 0.001597f
C11546 vss net6 0.096009f
C11547 output31/a_224_472# result[9] 0.082001f
C11548 net16 _064_ 0.121797f
C11549 _079_ FILLER_0_5_198/a_572_375# 0.011369f
C11550 _088_ FILLER_0_5_198/a_124_375# 0.001374f
C11551 net73 _145_ 0.009144f
C11552 net64 _055_ 0.00384f
C11553 _095_ FILLER_0_13_80/a_36_472# 0.004187f
C11554 state\[1\] FILLER_0_12_196/a_124_375# 0.063785f
C11555 _289_/a_244_68# _103_ 0.001153f
C11556 FILLER_0_10_256/a_124_375# FILLER_0_10_247/a_124_375# 0.002036f
C11557 _067_ net47 0.0609f
C11558 _189_/a_67_603# vdd 0.01494f
C11559 net72 _180_ 0.040135f
C11560 net16 _447_/a_1204_472# 0.00194f
C11561 net72 net15 0.157843f
C11562 _018_ _043_ 0.0022f
C11563 FILLER_0_4_197/a_36_472# vdd 0.042721f
C11564 FILLER_0_4_197/a_1468_375# vss 0.057762f
C11565 result[6] output18/a_224_472# 0.003068f
C11566 output33/a_224_472# ctlp[1] 0.018552f
C11567 FILLER_0_18_171/a_36_472# _143_ 0.005167f
C11568 net70 FILLER_0_14_99/a_124_375# 0.002922f
C11569 FILLER_0_8_107/a_124_375# _058_ 0.01823f
C11570 mask\[1\] FILLER_0_15_180/a_36_472# 0.001145f
C11571 _091_ net57 0.006076f
C11572 cal_itt\[2\] _260_/a_36_68# 0.004081f
C11573 net23 vdd 1.576398f
C11574 _104_ output34/a_224_472# 0.112239f
C11575 _424_/a_796_472# vdd 0.001951f
C11576 _186_ _181_ 0.018817f
C11577 vdd trim[2] 0.166648f
C11578 net20 _010_ 0.016197f
C11579 FILLER_0_23_290/a_124_375# vdd 0.030435f
C11580 _083_ FILLER_0_3_221/a_1380_472# 0.00181f
C11581 _441_/a_2248_156# vss 0.005663f
C11582 _441_/a_2665_112# vdd 0.012404f
C11583 _444_/a_36_151# net17 0.001435f
C11584 _219_/a_36_160# trim_mask\[0\] 0.395762f
C11585 trim_val\[2\] vss 0.027243f
C11586 FILLER_0_11_64/a_36_472# vss 0.006069f
C11587 _076_ _125_ 0.009254f
C11588 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_484_472# 0.013276f
C11589 _071_ _314_/a_224_472# 0.001359f
C11590 _352_/a_49_472# mask\[7\] 0.001066f
C11591 net55 _452_/a_1040_527# 0.021721f
C11592 _015_ _426_/a_2248_156# 0.021465f
C11593 net57 net53 0.053565f
C11594 _447_/a_1000_472# vdd 0.003392f
C11595 FILLER_0_18_2/a_484_472# vdd 0.003495f
C11596 FILLER_0_18_2/a_36_472# vss 0.001872f
C11597 _114_ FILLER_0_11_101/a_572_375# 0.051108f
C11598 fanout74/a_36_113# vdd 0.099021f
C11599 _066_ net37 0.006164f
C11600 net34 _299_/a_36_472# 0.003396f
C11601 result[4] FILLER_0_17_282/a_124_375# 0.018106f
C11602 _431_/a_2248_156# vss 0.041929f
C11603 _431_/a_2665_112# vdd 0.015335f
C11604 net76 FILLER_0_1_192/a_36_472# 0.003817f
C11605 _148_ _352_/a_49_472# 0.003082f
C11606 net35 mask\[7\] 0.954332f
C11607 _446_/a_448_472# _035_ 0.018273f
C11608 FILLER_0_14_50/a_124_375# _401_/a_36_68# 0.001129f
C11609 _430_/a_2248_156# _069_ 0.042876f
C11610 result[2] net30 0.019568f
C11611 _439_/a_1204_472# vss 0.006567f
C11612 _127_ _321_/a_170_472# 0.023836f
C11613 _372_/a_170_472# _152_ 0.037088f
C11614 _131_ _152_ 0.002949f
C11615 _412_/a_1204_472# net58 0.018724f
C11616 net35 _148_ 0.114816f
C11617 _214_/a_36_160# _213_/a_67_603# 0.002505f
C11618 _411_/a_1308_423# vss 0.0013f
C11619 output13/a_224_472# net22 0.022308f
C11620 _176_ FILLER_0_10_107/a_36_472# 0.009019f
C11621 _386_/a_124_24# _169_ 0.02709f
C11622 _098_ _437_/a_2248_156# 0.008669f
C11623 vdd FILLER_0_14_235/a_124_375# -0.011193f
C11624 FILLER_0_7_104/a_1380_472# _131_ 0.043557f
C11625 FILLER_0_24_96/a_124_375# output25/a_224_472# 0.002633f
C11626 _093_ FILLER_0_16_115/a_36_472# 0.001526f
C11627 input4/a_36_68# en 0.064323f
C11628 FILLER_0_21_125/a_572_375# _022_ 0.006025f
C11629 _018_ net21 0.077174f
C11630 _055_ vss 0.365503f
C11631 net61 _108_ 0.030767f
C11632 FILLER_0_4_152/a_36_472# net23 0.047194f
C11633 _163_ _385_/a_36_68# 0.012699f
C11634 FILLER_0_15_180/a_36_472# vss 0.00138f
C11635 FILLER_0_15_180/a_484_472# vdd 0.037927f
C11636 _132_ FILLER_0_18_107/a_1380_472# 0.034976f
C11637 net15 _441_/a_1000_472# 0.025912f
C11638 net67 _054_ 0.391592f
C11639 FILLER_0_16_57/a_1468_375# net55 0.006307f
C11640 FILLER_0_16_57/a_932_472# net72 0.004262f
C11641 _025_ vdd 0.259346f
C11642 _447_/a_448_472# net15 0.001766f
C11643 fanout82/a_36_113# output48/a_224_472# 0.009784f
C11644 _164_ FILLER_0_6_47/a_124_375# 0.069738f
C11645 net67 FILLER_0_8_24/a_36_472# 0.001252f
C11646 _086_ FILLER_0_6_177/a_36_472# 0.064045f
C11647 net65 net58 1.468105f
C11648 FILLER_0_15_10/a_36_472# vdd 0.086171f
C11649 FILLER_0_15_10/a_124_375# vss 0.002173f
C11650 net19 _416_/a_2665_112# 0.059453f
C11651 net20 FILLER_0_7_233/a_124_375# 0.017217f
C11652 net15 _439_/a_796_472# 0.001822f
C11653 fanout66/a_36_113# net66 0.032757f
C11654 _311_/a_1660_473# vdd 0.001435f
C11655 FILLER_0_9_28/a_484_472# net16 0.021584f
C11656 net65 _425_/a_2665_112# 0.00628f
C11657 mask\[5\] FILLER_0_18_177/a_1468_375# 0.002726f
C11658 net33 vdd 0.42212f
C11659 _274_/a_36_68# net81 0.014689f
C11660 _313_/a_67_603# vss 0.016047f
C11661 _114_ FILLER_0_10_94/a_36_472# 0.08191f
C11662 _137_ FILLER_0_17_104/a_1020_375# 0.001676f
C11663 mask\[2\] FILLER_0_16_154/a_124_375# 0.087247f
C11664 net31 net19 0.023019f
C11665 FILLER_0_18_2/a_1380_472# _452_/a_448_472# 0.059367f
C11666 _430_/a_448_472# net21 0.03842f
C11667 _110_ net71 0.004816f
C11668 net36 FILLER_0_15_212/a_36_472# 0.005396f
C11669 _435_/a_1204_472# vdd 0.013805f
C11670 _326_/a_36_160# FILLER_0_9_105/a_484_472# 0.002647f
C11671 _062_ FILLER_0_5_136/a_36_472# 0.001404f
C11672 _094_ mask\[2\] 0.089828f
C11673 net68 _232_/a_67_603# 0.00184f
C11674 _131_ _136_ 1.42765f
C11675 _370_/a_692_472# net47 0.001021f
C11676 vss FILLER_0_6_231/a_124_375# 0.00353f
C11677 vdd FILLER_0_6_231/a_572_375# 0.018694f
C11678 _056_ vdd 0.423512f
C11679 _427_/a_2665_112# vss 0.01229f
C11680 mask\[4\] output18/a_224_472# 0.017718f
C11681 FILLER_0_7_72/a_3172_472# vss 0.002425f
C11682 _414_/a_36_151# _089_ 0.039611f
C11683 FILLER_0_15_282/a_484_472# net18 0.018113f
C11684 _337_/a_665_69# mask\[1\] 0.002125f
C11685 FILLER_0_4_177/a_572_375# net22 0.006125f
C11686 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_572_375# 0.026339f
C11687 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_36_472# 0.001723f
C11688 trim_val\[1\] _166_ 0.06773f
C11689 FILLER_0_9_28/a_36_472# vdd 0.086674f
C11690 FILLER_0_9_28/a_3260_375# vss 0.05542f
C11691 FILLER_0_9_223/a_484_472# _128_ 0.005152f
C11692 FILLER_0_10_28/a_124_375# _450_/a_3129_107# 0.010735f
C11693 FILLER_0_8_24/a_484_472# _054_ 0.009315f
C11694 FILLER_0_14_263/a_124_375# output30/a_224_472# 0.011584f
C11695 _451_/a_836_156# _040_ 0.016371f
C11696 output35/a_224_472# FILLER_0_21_206/a_36_472# 0.0323f
C11697 _114_ _136_ 0.003405f
C11698 _032_ _370_/a_124_24# 0.007035f
C11699 net82 net9 0.004599f
C11700 trim_val\[4\] vdd 0.245329f
C11701 net52 FILLER_0_2_111/a_572_375# 0.00245f
C11702 _372_/a_170_472# _070_ 0.024545f
C11703 _131_ _070_ 0.161861f
C11704 _069_ _090_ 1.067281f
C11705 FILLER_0_8_138/a_124_375# _076_ 0.031436f
C11706 fanout62/a_36_160# FILLER_0_11_282/a_124_375# 0.058702f
C11707 _392_/a_36_68# vdd 0.036386f
C11708 FILLER_0_8_37/a_572_375# _054_ 0.137749f
C11709 net68 _453_/a_1000_472# 0.001816f
C11710 result[2] FILLER_0_15_282/a_124_375# 0.001114f
C11711 _257_/a_36_472# _074_ 0.011352f
C11712 FILLER_0_1_98/a_36_472# vss 0.002275f
C11713 _072_ _267_/a_36_472# 0.024239f
C11714 FILLER_0_13_212/a_1468_375# vss 0.062822f
C11715 FILLER_0_13_212/a_36_472# vdd 0.105926f
C11716 FILLER_0_6_177/a_572_375# _163_ 0.001839f
C11717 _053_ _068_ 0.066662f
C11718 fanout80/a_36_113# vdd 0.033884f
C11719 ctln[4] ctln[5] 0.031901f
C11720 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_36_472# 0.007947f
C11721 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_124_375# 0.001597f
C11722 FILLER_0_20_107/a_36_472# net71 0.004375f
C11723 FILLER_0_17_72/a_2364_375# _131_ 0.006037f
C11724 _096_ FILLER_0_12_196/a_124_375# 0.002309f
C11725 _157_ net14 0.026868f
C11726 _106_ net64 0.001587f
C11727 _016_ FILLER_0_12_136/a_484_472# 0.001516f
C11728 FILLER_0_11_109/a_36_472# _135_ 0.001891f
C11729 FILLER_0_13_80/a_36_472# vss 0.009445f
C11730 FILLER_0_5_72/a_932_472# net47 0.003953f
C11731 FILLER_0_4_177/a_124_375# _087_ 0.002288f
C11732 _114_ _070_ 0.507391f
C11733 _275_/a_224_472# mask\[3\] 0.002528f
C11734 FILLER_0_4_99/a_124_375# _153_ 0.030839f
C11735 _106_ mask\[1\] 0.005728f
C11736 _069_ net22 0.327999f
C11737 _430_/a_36_151# _138_ 0.001123f
C11738 _058_ vss 0.19427f
C11739 FILLER_0_24_290/a_36_472# FILLER_0_23_290/a_36_472# 0.05841f
C11740 net52 FILLER_0_6_79/a_124_375# 0.010099f
C11741 FILLER_0_9_223/a_484_472# state\[0\] 0.007034f
C11742 _111_ FILLER_0_18_76/a_124_375# 0.002494f
C11743 _428_/a_796_472# _095_ 0.00117f
C11744 trim_val\[1\] trim_mask\[1\] 0.519723f
C11745 _315_/a_36_68# vss 0.02467f
C11746 _274_/a_2552_68# _070_ 0.001238f
C11747 result[7] FILLER_0_24_274/a_572_375# 0.006125f
C11748 net74 FILLER_0_13_80/a_36_472# 0.00679f
C11749 net81 _069_ 0.034401f
C11750 _272_/a_36_472# _003_ 0.001634f
C11751 _408_/a_244_524# net47 0.001066f
C11752 net16 _174_ 0.022224f
C11753 mask\[7\] FILLER_0_22_128/a_1468_375# 0.0178f
C11754 _159_ _160_ 0.021804f
C11755 _057_ _311_/a_1660_473# 0.004637f
C11756 trimb[3] vdd 0.283005f
C11757 FILLER_0_5_198/a_572_375# vss 0.055087f
C11758 FILLER_0_5_198/a_36_472# vdd 0.088893f
C11759 _260_/a_36_68# net59 0.004346f
C11760 net74 _058_ 0.026905f
C11761 FILLER_0_16_241/a_124_375# vdd 0.035603f
C11762 net39 _444_/a_36_151# 0.14155f
C11763 _074_ FILLER_0_5_164/a_572_375# 0.001307f
C11764 net72 FILLER_0_21_28/a_1380_472# 0.048287f
C11765 _095_ FILLER_0_15_72/a_572_375# 0.00352f
C11766 _412_/a_796_472# net81 0.038712f
C11767 net16 _444_/a_2248_156# 0.065914f
C11768 FILLER_0_11_142/a_36_472# net23 0.002015f
C11769 net35 FILLER_0_22_128/a_932_472# 0.007806f
C11770 _276_/a_36_160# FILLER_0_18_209/a_572_375# 0.004736f
C11771 net36 _451_/a_1040_527# 0.00974f
C11772 FILLER_0_8_24/a_572_375# net47 0.0353f
C11773 output21/a_224_472# mask\[6\] 0.013037f
C11774 _149_ FILLER_0_20_107/a_124_375# 0.001244f
C11775 cal_count\[1\] FILLER_0_13_80/a_36_472# 0.001559f
C11776 FILLER_0_19_155/a_124_375# _145_ 0.006057f
C11777 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_484_472# 0.001963f
C11778 cal_count\[3\] net40 0.080767f
C11779 _057_ _056_ 0.167928f
C11780 FILLER_0_9_72/a_484_472# _439_/a_36_151# 0.001723f
C11781 net64 FILLER_0_9_282/a_124_375# 0.046477f
C11782 FILLER_0_11_64/a_124_375# cal_count\[3\] 0.002495f
C11783 trim_mask\[1\] FILLER_0_6_47/a_3260_375# 0.003764f
C11784 _155_ net47 0.009532f
C11785 _274_/a_2960_68# _091_ 0.001338f
C11786 net63 FILLER_0_22_177/a_484_472# 0.059367f
C11787 result[6] _419_/a_2248_156# 0.002634f
C11788 _106_ vss 0.180823f
C11789 _074_ _251_/a_1130_472# 0.00237f
C11790 FILLER_0_22_128/a_1828_472# vdd 0.005724f
C11791 FILLER_0_22_128/a_1380_472# vss 0.007305f
C11792 net55 FILLER_0_17_64/a_36_472# 0.034504f
C11793 _052_ FILLER_0_18_37/a_124_375# 0.03242f
C11794 _093_ _199_/a_36_160# 0.05226f
C11795 _444_/a_1204_472# vdd 0.001086f
C11796 FILLER_0_16_73/a_36_472# _176_ 0.013449f
C11797 _128_ calibrate 0.039365f
C11798 _446_/a_36_151# vdd 0.06703f
C11799 _126_ _136_ 0.086459f
C11800 _421_/a_36_151# _419_/a_2248_156# 0.001203f
C11801 _075_ net22 0.180274f
C11802 FILLER_0_7_59/a_484_472# net15 0.015199f
C11803 FILLER_0_21_142/a_572_375# _433_/a_2248_156# 0.006739f
C11804 FILLER_0_21_142/a_124_375# _433_/a_2665_112# 0.004834f
C11805 FILLER_0_15_282/a_484_472# net62 0.009524f
C11806 _452_/a_448_472# _041_ 0.007f
C11807 net41 _095_ 0.641184f
C11808 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2724_472# 0.026657f
C11809 result[7] FILLER_0_23_274/a_36_472# 0.014434f
C11810 _016_ FILLER_0_12_124/a_124_375# 0.007335f
C11811 FILLER_0_16_57/a_572_375# FILLER_0_17_56/a_572_375# 0.026339f
C11812 net65 _413_/a_2665_112# 0.033675f
C11813 net22 FILLER_0_18_209/a_484_472# 0.005297f
C11814 FILLER_0_10_78/a_484_472# vss 0.005854f
C11815 FILLER_0_10_78/a_932_472# vdd 0.005517f
C11816 output38/a_224_472# net66 0.148811f
C11817 FILLER_0_7_72/a_124_375# FILLER_0_5_72/a_36_472# 0.001512f
C11818 FILLER_0_15_142/a_36_472# _136_ 0.003745f
C11819 _428_/a_2560_156# net53 0.002265f
C11820 FILLER_0_21_28/a_1380_472# _424_/a_36_151# 0.001723f
C11821 _413_/a_1000_472# net21 0.041643f
C11822 mask\[8\] FILLER_0_22_107/a_572_375# 0.030641f
C11823 net35 FILLER_0_22_107/a_124_375# 0.010439f
C11824 _314_/a_224_472# net23 0.001238f
C11825 _274_/a_1164_497# net64 0.002049f
C11826 output42/a_224_472# vss 0.00418f
C11827 _307_/a_234_472# _085_ 0.001966f
C11828 net34 output18/a_224_472# 0.17524f
C11829 FILLER_0_18_2/a_2276_472# net38 0.002313f
C11830 _069_ _076_ 0.033276f
C11831 _126_ _070_ 0.089475f
C11832 net63 FILLER_0_18_177/a_36_472# 0.015187f
C11833 net20 _411_/a_36_151# 0.011179f
C11834 _245_/a_672_472# _039_ 0.001025f
C11835 FILLER_0_5_54/a_1380_472# net47 0.003924f
C11836 _097_ FILLER_0_15_180/a_36_472# 0.005242f
C11837 _095_ _406_/a_36_159# 0.131137f
C11838 _093_ net55 0.182194f
C11839 _077_ FILLER_0_10_94/a_36_472# 0.001114f
C11840 _119_ _313_/a_67_603# 0.015457f
C11841 net82 FILLER_0_3_172/a_1380_472# 0.007879f
C11842 _449_/a_36_151# _043_ 0.001572f
C11843 FILLER_0_15_116/a_572_375# _136_ 0.001706f
C11844 net4 FILLER_0_12_236/a_484_472# 0.014212f
C11845 _176_ _451_/a_36_151# 0.003176f
C11846 output14/a_224_472# _442_/a_2248_156# 0.001723f
C11847 FILLER_0_9_282/a_124_375# vss 0.00451f
C11848 FILLER_0_9_282/a_572_375# vdd 0.002928f
C11849 _122_ _066_ 0.001217f
C11850 FILLER_0_4_144/a_572_375# _081_ 0.002236f
C11851 vss _167_ 0.043544f
C11852 FILLER_0_4_144/a_124_375# _152_ 0.007333f
C11853 _414_/a_1204_472# net21 0.007637f
C11854 _327_/a_36_472# net74 0.009344f
C11855 vdd FILLER_0_22_107/a_36_472# 0.114332f
C11856 vss FILLER_0_22_107/a_572_375# 0.001944f
C11857 _094_ _418_/a_1000_472# 0.053462f
C11858 state\[0\] calibrate 0.001061f
C11859 state\[1\] _121_ 0.006184f
C11860 _046_ vdd 0.041841f
C11861 _394_/a_2215_68# _095_ 0.001134f
C11862 mask\[4\] FILLER_0_20_177/a_1380_472# 0.001215f
C11863 ctln[2] rstn 0.017812f
C11864 _053_ vdd 1.467835f
C11865 _127_ _135_ 0.00622f
C11866 net27 _425_/a_2248_156# 0.027078f
C11867 net52 _440_/a_448_472# 0.067294f
C11868 output22/a_224_472# _024_ 0.029795f
C11869 FILLER_0_18_171/a_36_472# FILLER_0_18_177/a_36_472# 0.003468f
C11870 FILLER_0_13_100/a_36_472# _043_ 0.012726f
C11871 FILLER_0_18_107/a_484_472# FILLER_0_17_104/a_932_472# 0.026657f
C11872 _176_ _124_ 0.036117f
C11873 _189_/a_67_603# FILLER_0_13_228/a_36_472# 0.005759f
C11874 _053_ FILLER_0_7_72/a_2364_375# 0.015932f
C11875 _147_ net23 0.011375f
C11876 _015_ vdd 0.27747f
C11877 _122_ FILLER_0_8_156/a_484_472# 0.007378f
C11878 net60 net33 0.008865f
C11879 _104_ _422_/a_2665_112# 0.040586f
C11880 FILLER_0_20_15/a_1468_375# vss 0.055156f
C11881 FILLER_0_20_15/a_36_472# vdd 0.086947f
C11882 mask\[4\] FILLER_0_18_177/a_1020_375# 0.015941f
C11883 _129_ FILLER_0_11_135/a_36_472# 0.078373f
C11884 net69 _152_ 0.002532f
C11885 _443_/a_2248_156# trim_mask\[4\] 0.002315f
C11886 net50 FILLER_0_4_91/a_572_375# 0.007234f
C11887 output34/a_224_472# result[7] 0.057094f
C11888 net82 _084_ 0.020793f
C11889 _122_ net37 3.870625f
C11890 _016_ fanout73/a_36_113# 0.001731f
C11891 net76 _078_ 0.029213f
C11892 FILLER_0_17_72/a_1020_375# _175_ 0.028592f
C11893 _321_/a_170_472# net23 0.025371f
C11894 _140_ FILLER_0_22_128/a_2276_472# 0.002954f
C11895 _074_ _082_ 0.069835f
C11896 _093_ net23 0.042838f
C11897 mask\[8\] _214_/a_36_160# 0.001264f
C11898 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_1020_375# 0.026339f
C11899 _132_ FILLER_0_14_107/a_1380_472# 0.049391f
C11900 net57 _071_ 0.12089f
C11901 trimb[3] output17/a_224_472# 0.047604f
C11902 FILLER_0_0_232/a_36_472# vdd 0.050082f
C11903 FILLER_0_0_232/a_124_375# vss 0.019863f
C11904 _441_/a_2665_112# FILLER_0_3_78/a_572_375# 0.010688f
C11905 output13/a_224_472# _448_/a_2665_112# 0.027303f
C11906 trim_mask\[2\] FILLER_0_3_78/a_484_472# 0.008122f
C11907 _392_/a_36_68# cal_count\[0\] 0.038691f
C11908 _013_ FILLER_0_17_56/a_572_375# 0.001047f
C11909 result[0] fanout65/a_36_113# 0.001816f
C11910 mask\[5\] _146_ 0.051687f
C11911 _143_ _137_ 0.009932f
C11912 net81 FILLER_0_15_235/a_36_472# 0.001855f
C11913 net75 _001_ 0.056236f
C11914 _077_ _070_ 0.29321f
C11915 _256_/a_1164_497# net4 0.004729f
C11916 _128_ _125_ 0.017316f
C11917 _411_/a_2248_156# _084_ 0.002258f
C11918 _422_/a_796_472# _109_ 0.002086f
C11919 net50 net16 0.015448f
C11920 _070_ FILLER_0_10_107/a_124_375# 0.009848f
C11921 trim_val\[0\] _453_/a_36_151# 0.001629f
C11922 _449_/a_2665_112# _172_ 0.003296f
C11923 _128_ _315_/a_1657_68# 0.0013f
C11924 _428_/a_1000_472# vdd 0.005345f
C11925 cal input4/a_36_68# 0.054357f
C11926 net69 FILLER_0_2_127/a_36_472# 0.019383f
C11927 _119_ _058_ 0.692466f
C11928 FILLER_0_15_142/a_484_472# net53 0.044267f
C11929 FILLER_0_5_54/a_124_375# vdd 0.007387f
C11930 ctln[8] trim_val\[3\] 0.007f
C11931 ctln[2] FILLER_0_1_266/a_484_472# 0.019076f
C11932 net49 net17 0.029142f
C11933 _089_ net21 0.006605f
C11934 _214_/a_36_160# vss 0.007045f
C11935 _072_ _118_ 0.120452f
C11936 net36 _006_ 0.001331f
C11937 net57 _386_/a_692_472# 0.00409f
C11938 net68 net17 0.601273f
C11939 net75 output48/a_224_472# 0.070114f
C11940 fanout76/a_36_160# vss 0.028897f
C11941 net68 _377_/a_36_472# 0.001305f
C11942 _061_ FILLER_0_8_156/a_484_472# 0.00255f
C11943 net31 _047_ 0.029502f
C11944 FILLER_0_4_177/a_124_375# vdd 0.021637f
C11945 FILLER_0_17_282/a_124_375# _417_/a_36_151# 0.059049f
C11946 FILLER_0_15_72/a_572_375# vss 0.007579f
C11947 FILLER_0_15_72/a_36_472# vdd 0.108844f
C11948 net37 FILLER_0_6_231/a_484_472# 0.004323f
C11949 net57 FILLER_0_8_156/a_572_375# 0.014948f
C11950 _415_/a_36_151# net19 0.05689f
C11951 _136_ _137_ 0.417639f
C11952 FILLER_0_15_116/a_36_472# net53 0.005099f
C11953 net52 vss 1.608047f
C11954 net21 _434_/a_2665_112# 0.004945f
C11955 _013_ _041_ 0.00271f
C11956 output32/a_224_472# net32 0.014826f
C11957 net20 FILLER_0_13_212/a_572_375# 0.002085f
C11958 net48 _425_/a_448_472# 0.013011f
C11959 _141_ FILLER_0_19_155/a_572_375# 0.033271f
C11960 _440_/a_36_151# _164_ 0.003699f
C11961 _443_/a_796_472# vss 0.001654f
C11962 trim_mask\[4\] _170_ 0.09738f
C11963 _132_ _140_ 0.019255f
C11964 _033_ FILLER_0_6_37/a_124_375# 0.018812f
C11965 result[8] FILLER_0_23_290/a_36_472# 0.001414f
C11966 FILLER_0_7_72/a_1916_375# net50 0.059471f
C11967 result[1] _416_/a_36_151# 0.007739f
C11968 _345_/a_36_160# _144_ 0.00465f
C11969 net36 FILLER_0_15_228/a_36_472# 0.008225f
C11970 net27 _426_/a_1308_423# 0.00384f
C11971 output22/a_224_472# _435_/a_1308_423# 0.005111f
C11972 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_36_472# 0.086904f
C11973 _431_/a_1308_423# net36 0.002865f
C11974 mask\[2\] net21 0.033368f
C11975 _444_/a_36_151# net42 0.006866f
C11976 _350_/a_49_472# _208_/a_36_160# 0.078981f
C11977 _147_ net33 0.001686f
C11978 net18 vdd 1.496006f
C11979 _289_/a_36_472# _094_ 0.00922f
C11980 FILLER_0_16_57/a_124_375# _131_ 0.012982f
C11981 FILLER_0_3_204/a_36_472# FILLER_0_4_197/a_932_472# 0.026657f
C11982 _065_ _238_/a_67_603# 0.005075f
C11983 FILLER_0_1_212/a_36_472# vss 0.00858f
C11984 FILLER_0_7_59/a_36_472# fanout67/a_36_160# 0.013068f
C11985 _067_ FILLER_0_13_72/a_124_375# 0.001782f
C11986 _216_/a_67_603# vss 0.012211f
C11987 net19 FILLER_0_23_274/a_124_375# 0.01233f
C11988 trim_val\[0\] FILLER_0_6_47/a_572_375# 0.03235f
C11989 net55 _424_/a_2665_112# 0.056555f
C11990 FILLER_0_15_72/a_572_375# cal_count\[1\] 0.135344f
C11991 _114_ _255_/a_224_552# 0.005131f
C11992 net16 FILLER_0_18_37/a_1468_375# 0.002269f
C11993 net41 vss 0.810444f
C11994 _448_/a_2248_156# _443_/a_2248_156# 0.006556f
C11995 FILLER_0_18_2/a_572_375# net44 0.072627f
C11996 _004_ net75 0.003999f
C11997 FILLER_0_18_2/a_2276_472# net55 0.006033f
C11998 _360_/a_36_160# vdd 0.006439f
C11999 _144_ FILLER_0_21_133/a_124_375# 0.001885f
C12000 ctlp[1] _419_/a_1308_423# 0.00678f
C12001 FILLER_0_10_78/a_36_472# FILLER_0_9_72/a_572_375# 0.001543f
C12002 _412_/a_1308_423# vdd 0.003842f
C12003 _232_/a_67_603# net47 0.014888f
C12004 _072_ _068_ 0.185471f
C12005 _387_/a_36_113# vss 0.047621f
C12006 FILLER_0_3_204/a_124_375# net82 0.014222f
C12007 FILLER_0_5_109/a_124_375# _151_ 0.003377f
C12008 _164_ vdd 0.711488f
C12009 _431_/a_2248_156# FILLER_0_17_142/a_572_375# 0.006739f
C12010 _431_/a_2665_112# FILLER_0_17_142/a_124_375# 0.004834f
C12011 _406_/a_36_159# vss 0.002509f
C12012 _414_/a_2248_156# _074_ 0.013023f
C12013 FILLER_0_21_286/a_484_472# vss 0.008522f
C12014 FILLER_0_18_37/a_1020_375# vdd 0.020683f
C12015 net79 FILLER_0_12_236/a_484_472# 0.009305f
C12016 net81 output27/a_224_472# 0.011872f
C12017 FILLER_0_10_78/a_36_472# cal_count\[3\] 0.266339f
C12018 output44/a_224_472# _452_/a_1353_112# 0.001321f
C12019 _090_ net22 0.032492f
C12020 _127_ _129_ 0.716384f
C12021 _091_ FILLER_0_19_171/a_484_472# 0.013944f
C12022 FILLER_0_6_90/a_124_375# net14 0.005361f
C12023 _065_ net15 0.065255f
C12024 _095_ _450_/a_448_472# 0.001393f
C12025 _077_ FILLER_0_12_50/a_36_472# 0.177624f
C12026 _413_/a_36_151# FILLER_0_3_172/a_3260_375# 0.059049f
C12027 net38 _444_/a_1288_156# 0.001147f
C12028 cal_count\[2\] _402_/a_244_567# 0.004411f
C12029 _411_/a_36_151# _073_ 0.00135f
C12030 fanout57/a_36_113# vdd 0.005473f
C12031 _134_ FILLER_0_9_105/a_484_472# 0.011499f
C12032 output43/a_224_472# net17 0.083607f
C12033 _448_/a_2248_156# _170_ 0.00254f
C12034 _448_/a_1000_472# _037_ 0.03564f
C12035 FILLER_0_10_28/a_36_472# vss 0.001102f
C12036 _062_ _310_/a_49_472# 0.020509f
C12037 _050_ FILLER_0_22_128/a_36_472# 0.001098f
C12038 _265_/a_916_472# _001_ 0.001719f
C12039 net72 _067_ 0.055817f
C12040 net56 _136_ 0.462275f
C12041 _442_/a_36_151# net23 0.00157f
C12042 _078_ _083_ 0.01015f
C12043 _132_ _149_ 0.087289f
C12044 _165_ trim_val\[0\] 0.164683f
C12045 _053_ FILLER_0_6_47/a_3172_472# 0.001777f
C12046 _436_/a_36_151# _025_ 0.026707f
C12047 fanout75/a_36_113# vdd 0.028614f
C12048 _441_/a_448_472# net49 0.001245f
C12049 result[7] _419_/a_1000_472# 0.015362f
C12050 FILLER_0_16_89/a_1380_472# vdd 0.010554f
C12051 _432_/a_36_151# vdd 0.173104f
C12052 FILLER_0_18_2/a_3172_472# net40 0.046864f
C12053 _028_ _153_ 0.008011f
C12054 _172_ vss 0.054608f
C12055 _235_/a_67_603# net68 0.027525f
C12056 _445_/a_448_472# net40 0.044285f
C12057 _181_ _179_ 0.011848f
C12058 _009_ FILLER_0_23_274/a_124_375# 0.010723f
C12059 FILLER_0_18_209/a_572_375# vss 0.007545f
C12060 FILLER_0_18_209/a_36_472# vdd 0.089327f
C12061 net49 _440_/a_1204_472# 0.006692f
C12062 net81 net22 0.064261f
C12063 net7 ctln[9] 0.005103f
C12064 _414_/a_2560_156# cal_itt\[3\] 0.007141f
C12065 trim[4] net38 0.095379f
C12066 FILLER_0_15_116/a_484_472# FILLER_0_14_107/a_1468_375# 0.001723f
C12067 net64 FILLER_0_15_235/a_124_375# 0.025203f
C12068 output36/a_224_472# FILLER_0_14_263/a_36_472# 0.001711f
C12069 _394_/a_1936_472# net15 0.001592f
C12070 ctln[3] vdd 0.167569f
C12071 _104_ _011_ 0.021454f
C12072 _442_/a_2248_156# _157_ 0.002731f
C12073 _032_ _031_ 0.013851f
C12074 net57 net55 0.001926f
C12075 _091_ FILLER_0_15_212/a_124_375# 0.025529f
C12076 _431_/a_1308_423# _020_ 0.001997f
C12077 _003_ _074_ 0.00476f
C12078 FILLER_0_15_235/a_124_375# mask\[1\] 0.013103f
C12079 _415_/a_2560_156# net27 0.008433f
C12080 net74 _172_ 0.006643f
C12081 _440_/a_2665_112# trim_mask\[1\] 0.007959f
C12082 trimb[1] FILLER_0_20_2/a_484_472# 0.003628f
C12083 net65 sample 0.148853f
C12084 FILLER_0_18_61/a_36_472# vdd 0.08828f
C12085 FILLER_0_18_61/a_124_375# vss 0.021307f
C12086 FILLER_0_12_50/a_36_472# _453_/a_36_151# 0.001748f
C12087 net58 net64 0.590523f
C12088 vdd net62 1.53102f
C12089 _070_ _248_/a_36_68# 0.007095f
C12090 net39 net49 0.158007f
C12091 FILLER_0_17_104/a_1468_375# vdd 0.022331f
C12092 net2 net18 0.030437f
C12093 net55 FILLER_0_17_56/a_484_472# 0.023554f
C12094 net7 vss 0.117948f
C12095 _044_ output30/a_224_472# 0.00717f
C12096 FILLER_0_5_128/a_36_472# _360_/a_36_160# 0.195479f
C12097 FILLER_0_5_164/a_484_472# vss 0.003257f
C12098 net82 calibrate 0.002345f
C12099 mask\[3\] _141_ 0.361692f
C12100 _413_/a_1308_423# _002_ 0.002178f
C12101 net39 _445_/a_1204_472# 0.002681f
C12102 net52 FILLER_0_9_72/a_124_375# 0.029702f
C12103 FILLER_0_21_286/a_124_375# net77 0.00301f
C12104 net20 _099_ 0.011124f
C12105 _070_ _060_ 0.822179f
C12106 _274_/a_36_68# state\[0\] 0.001852f
C12107 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_572_375# 0.086635f
C12108 net75 _316_/a_124_24# 0.003078f
C12109 FILLER_0_12_220/a_1380_472# _060_ 0.01563f
C12110 net44 _452_/a_3129_107# 0.067848f
C12111 FILLER_0_16_107/a_572_375# FILLER_0_18_107/a_484_472# 0.001512f
C12112 FILLER_0_11_64/a_124_375# _120_ 0.004514f
C12113 FILLER_0_19_171/a_572_375# vdd 0.022516f
C12114 _323_/a_36_113# _223_/a_36_160# 0.238626f
C12115 state\[2\] FILLER_0_13_142/a_484_472# 0.004186f
C12116 net57 net23 0.324262f
C12117 net53 FILLER_0_13_142/a_1380_472# 0.041222f
C12118 _442_/a_3041_156# vdd 0.001178f
C12119 FILLER_0_15_235/a_124_375# vss 0.001993f
C12120 FILLER_0_15_235/a_572_375# vdd -0.005887f
C12121 trim_val\[3\] vdd 0.211478f
C12122 net65 net9 0.061456f
C12123 FILLER_0_18_177/a_2364_375# net21 0.018463f
C12124 net36 net14 0.037175f
C12125 _091_ net27 0.023019f
C12126 _072_ vdd 0.715894f
C12127 _128_ _069_ 0.018491f
C12128 _176_ _180_ 0.030701f
C12129 _076_ net22 0.03249f
C12130 _176_ net15 0.038396f
C12131 FILLER_0_20_107/a_124_375# _098_ 0.01186f
C12132 ctln[4] FILLER_0_1_204/a_124_375# 0.008283f
C12133 _077_ _255_/a_224_552# 0.025141f
C12134 vss net30 0.17209f
C12135 _032_ _371_/a_36_113# 0.030245f
C12136 net58 vss 0.589419f
C12137 FILLER_0_6_90/a_484_472# _163_ 0.011711f
C12138 FILLER_0_9_28/a_1020_375# net68 0.004803f
C12139 net73 FILLER_0_18_107/a_3260_375# 0.001629f
C12140 FILLER_0_0_130/a_124_375# vdd 0.012493f
C12141 FILLER_0_2_93/a_36_472# net69 0.010977f
C12142 FILLER_0_16_107/a_572_375# _136_ 0.006445f
C12143 FILLER_0_16_89/a_572_375# net14 0.00106f
C12144 _070_ _330_/a_224_472# 0.001096f
C12145 FILLER_0_18_177/a_1468_375# FILLER_0_20_177/a_1380_472# 0.0027f
C12146 _430_/a_1000_472# vss 0.001626f
C12147 _425_/a_2560_156# vdd 0.001827f
C12148 _425_/a_2665_112# vss 0.002983f
C12149 _069_ FILLER_0_11_142/a_572_375# 0.020472f
C12150 _086_ cal_itt\[3\] 0.046874f
C12151 _093_ _046_ 0.061989f
C12152 FILLER_0_20_98/a_36_472# vdd 0.095266f
C12153 FILLER_0_20_98/a_124_375# vss 0.013019f
C12154 _184_ net17 0.007958f
C12155 FILLER_0_18_107/a_36_472# mask\[9\] 0.005458f
C12156 result[9] _420_/a_2248_156# 0.046636f
C12157 _190_/a_36_160# _039_ 0.003926f
C12158 _036_ net15 0.036489f
C12159 _122_ FILLER_0_6_231/a_484_472# 0.017477f
C12160 _123_ FILLER_0_6_231/a_124_375# 0.001259f
C12161 _164_ FILLER_0_6_47/a_3172_472# 0.001058f
C12162 FILLER_0_4_177/a_36_472# net37 0.004017f
C12163 net60 net18 0.949607f
C12164 net78 net18 1.351707f
C12165 _426_/a_796_472# net64 0.006933f
C12166 _420_/a_796_472# vss 0.001659f
C12167 vss _450_/a_448_472# -0.001661f
C12168 _136_ _095_ 0.043768f
C12169 net70 _451_/a_1353_112# 0.00194f
C12170 net14 _160_ 0.034023f
C12171 _320_/a_1792_472# vdd 0.001113f
C12172 _109_ vdd 0.059259f
C12173 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_36_472# 0.026657f
C12174 FILLER_0_9_290/a_124_375# FILLER_0_9_282/a_572_375# 0.012001f
C12175 output32/a_224_472# _010_ 0.001508f
C12176 output20/a_224_472# _422_/a_1308_423# 0.005632f
C12177 mask\[3\] FILLER_0_17_218/a_572_375# 0.015907f
C12178 FILLER_0_21_125/a_484_472# vss 0.002399f
C12179 result[1] net79 0.25261f
C12180 _170_ _066_ 0.189122f
C12181 _449_/a_1204_472# _038_ 0.005899f
C12182 output33/a_224_472# net33 0.151281f
C12183 FILLER_0_13_142/a_1468_375# vdd 0.028002f
C12184 fanout53/a_36_160# vdd 0.016868f
C12185 FILLER_0_16_57/a_932_472# _176_ 0.010635f
C12186 FILLER_0_13_142/a_1020_375# vss 0.005307f
C12187 trimb[2] vss 0.102375f
C12188 net41 FILLER_0_21_28/a_484_472# 0.060027f
C12189 net34 _297_/a_36_472# 0.005603f
C12190 _187_ _173_ 0.03421f
C12191 FILLER_0_16_57/a_124_375# FILLER_0_15_59/a_36_472# 0.001543f
C12192 FILLER_0_8_107/a_124_375# _070_ 0.003069f
C12193 net31 _106_ 0.035117f
C12194 FILLER_0_7_59/a_124_375# net68 0.019553f
C12195 _012_ net71 0.004946f
C12196 net79 _416_/a_2560_156# 0.013576f
C12197 FILLER_0_8_247/a_1380_472# vdd 0.036604f
C12198 _421_/a_2248_156# vdd 0.035239f
C12199 _030_ net14 0.079892f
C12200 _077_ _039_ 0.104126f
C12201 trimb[0] vdd 0.10929f
C12202 ctln[5] _448_/a_36_151# 0.009209f
C12203 _133_ _068_ 0.002552f
C12204 net52 FILLER_0_3_78/a_36_472# 0.034084f
C12205 _422_/a_36_151# vss 0.014056f
C12206 output22/a_224_472# ctlp[5] 0.024131f
C12207 _422_/a_448_472# vdd 0.032865f
C12208 output9/a_224_472# net82 0.003636f
C12209 _378_/a_224_472# vdd 0.002263f
C12210 _057_ _072_ 0.048392f
C12211 FILLER_0_10_256/a_124_375# net27 0.006216f
C12212 net17 net47 2.009509f
C12213 _426_/a_1000_472# vdd 0.007031f
C12214 net26 net72 0.868238f
C12215 net57 trim_val\[4\] 0.295336f
C12216 _232_/a_67_603# FILLER_0_6_47/a_36_472# 0.010206f
C12217 FILLER_0_15_282/a_124_375# vss 0.004893f
C12218 FILLER_0_16_37/a_36_472# _184_ 0.001522f
C12219 FILLER_0_15_282/a_572_375# vdd 0.002928f
C12220 net54 _145_ 0.087336f
C12221 _446_/a_2248_156# net40 0.037373f
C12222 _074_ _162_ 0.112872f
C12223 FILLER_0_11_101/a_36_472# vdd 0.093852f
C12224 FILLER_0_11_101/a_572_375# vss 0.055325f
C12225 net80 _435_/a_1000_472# 0.001079f
C12226 net76 _263_/a_224_472# 0.00132f
C12227 _088_ FILLER_0_4_213/a_36_472# 0.01735f
C12228 net15 _183_ 0.007353f
C12229 _183_ _180_ 0.002621f
C12230 _285_/a_36_472# _196_/a_36_160# 0.004619f
C12231 net8 FILLER_0_0_266/a_124_375# 0.001181f
C12232 FILLER_0_3_221/a_124_375# vdd 0.008869f
C12233 _438_/a_448_472# net71 0.044454f
C12234 fanout80/a_36_113# FILLER_0_15_205/a_36_472# 0.010419f
C12235 FILLER_0_4_49/a_124_375# _164_ 0.017213f
C12236 _000_ _260_/a_36_68# 0.004354f
C12237 output11/a_224_472# FILLER_0_0_232/a_36_472# 0.023414f
C12238 _315_/a_716_497# _120_ 0.001321f
C12239 net63 _435_/a_2248_156# 0.045342f
C12240 ctln[2] net59 0.009218f
C12241 _412_/a_2665_112# fanout58/a_36_160# 0.001221f
C12242 output8/a_224_472# _411_/a_36_151# 0.12978f
C12243 _412_/a_2560_156# cal_itt\[1\] 0.00454f
C12244 _408_/a_56_524# net40 0.001367f
C12245 _394_/a_1336_472# FILLER_0_15_72/a_124_375# 0.016876f
C12246 output10/a_224_472# net10 0.012455f
C12247 _420_/a_36_151# net77 0.023469f
C12248 _013_ _012_ 0.003113f
C12249 ctln[2] net4 0.039098f
C12250 _152_ vss 0.140215f
C12251 net16 _217_/a_36_160# 0.00629f
C12252 _074_ net19 0.035973f
C12253 _077_ FILLER_0_8_156/a_36_472# 0.00563f
C12254 _136_ mask\[1\] 0.407932f
C12255 _021_ _098_ 0.014179f
C12256 _175_ _451_/a_3129_107# 0.021546f
C12257 FILLER_0_7_104/a_1380_472# vss 0.003236f
C12258 FILLER_0_8_24/a_124_375# net40 0.002431f
C12259 _114_ _395_/a_36_488# 0.005314f
C12260 net78 net62 0.001947f
C12261 net60 net62 0.002144f
C12262 _015_ FILLER_0_10_247/a_124_375# 0.001261f
C12263 FILLER_0_13_290/a_36_472# result[3] 0.001069f
C12264 net16 _035_ 0.034977f
C12265 FILLER_0_3_78/a_572_375# _164_ 0.055492f
C12266 _238_/a_67_603# output15/a_224_472# 0.019027f
C12267 _081_ FILLER_0_5_148/a_124_375# 0.021583f
C12268 _436_/a_2665_112# _050_ 0.030939f
C12269 _028_ trim_mask\[1\] 0.148182f
C12270 _036_ _381_/a_36_472# 0.023012f
C12271 net74 _152_ 1.007413f
C12272 _043_ FILLER_0_13_72/a_572_375# 0.013294f
C12273 net26 _424_/a_36_151# 0.062638f
C12274 _038_ FILLER_0_11_78/a_484_472# 0.001782f
C12275 FILLER_0_2_101/a_124_375# trim_mask\[3\] 0.033692f
C12276 FILLER_0_2_127/a_36_472# vss 0.002567f
C12277 FILLER_0_18_107/a_932_472# vdd 0.009633f
C12278 _413_/a_2665_112# vss 0.012213f
C12279 net65 _084_ 0.031674f
C12280 _267_/a_672_472# _071_ 0.00255f
C12281 FILLER_0_19_187/a_484_472# _434_/a_2665_112# 0.001868f
C12282 mask\[5\] _141_ 0.241158f
C12283 _208_/a_36_160# FILLER_0_22_128/a_2812_375# 0.026361f
C12284 net61 _419_/a_36_151# 0.019141f
C12285 vdd FILLER_0_10_94/a_484_472# 0.008627f
C12286 net54 FILLER_0_22_128/a_484_472# 0.055436f
C12287 _143_ vss 0.02001f
C12288 _448_/a_2665_112# net22 0.010428f
C12289 net64 FILLER_0_12_220/a_1380_472# 0.011079f
C12290 FILLER_0_18_139/a_484_472# _145_ 0.002415f
C12291 FILLER_0_16_89/a_1468_375# _040_ 0.004985f
C12292 FILLER_0_16_37/a_36_472# net47 0.008304f
C12293 output15/a_224_472# FILLER_0_0_96/a_36_472# 0.023414f
C12294 _058_ FILLER_0_9_105/a_124_375# 0.014234f
C12295 _348_/a_49_472# vss 0.002301f
C12296 _417_/a_1308_423# _006_ 0.022704f
C12297 trim_val\[0\] vss 0.11063f
C12298 FILLER_0_21_28/a_2812_375# _012_ 0.016736f
C12299 net74 _318_/a_224_472# 0.001513f
C12300 _014_ vss 0.034646f
C12301 net74 FILLER_0_2_127/a_36_472# 0.001261f
C12302 net63 FILLER_0_17_226/a_124_375# 0.00507f
C12303 FILLER_0_5_164/a_36_472# _169_ 0.00284f
C12304 FILLER_0_5_164/a_572_375# _163_ 0.046852f
C12305 _422_/a_2248_156# net19 0.003451f
C12306 _114_ _439_/a_2665_112# 0.011015f
C12307 FILLER_0_10_78/a_36_472# _120_ 0.004669f
C12308 FILLER_0_7_72/a_1020_375# FILLER_0_6_79/a_124_375# 0.026339f
C12309 _136_ vss 0.947188f
C12310 _104_ _198_/a_67_603# 0.007168f
C12311 _414_/a_2560_156# _081_ 0.008322f
C12312 output15/a_224_472# net15 0.028578f
C12313 net72 FILLER_0_17_38/a_36_472# 0.123542f
C12314 ctln[6] net59 0.001267f
C12315 _103_ net30 0.013544f
C12316 _432_/a_36_151# _093_ 0.018324f
C12317 _430_/a_36_151# FILLER_0_17_200/a_572_375# 0.059049f
C12318 _186_ vdd 0.074983f
C12319 net36 FILLER_0_20_87/a_36_472# 0.074773f
C12320 FILLER_0_22_177/a_36_472# mask\[6\] 0.006882f
C12321 _093_ FILLER_0_18_209/a_36_472# 0.007068f
C12322 net55 _027_ 0.002104f
C12323 mask\[4\] FILLER_0_19_155/a_484_472# 0.024522f
C12324 net74 _136_ 0.042043f
C12325 _431_/a_448_472# net70 0.002293f
C12326 trim_mask\[1\] FILLER_0_6_90/a_36_472# 0.001162f
C12327 net18 _416_/a_2248_156# 0.002106f
C12328 _133_ vdd 0.27652f
C12329 _070_ vss 1.363355f
C12330 _021_ FILLER_0_18_171/a_36_472# 0.103755f
C12331 FILLER_0_9_28/a_1020_375# FILLER_0_10_37/a_36_472# 0.001597f
C12332 _449_/a_796_472# vss 0.00143f
C12333 _104_ mask\[3\] 0.078406f
C12334 _440_/a_1204_472# net47 0.006257f
C12335 FILLER_0_12_220/a_1380_472# vss 0.006172f
C12336 net35 FILLER_0_22_86/a_572_375# 0.010986f
C12337 mask\[8\] FILLER_0_22_86/a_1020_375# 0.009431f
C12338 mask\[4\] FILLER_0_17_200/a_484_472# 0.001701f
C12339 net52 _442_/a_448_472# 0.044149f
C12340 FILLER_0_5_128/a_484_472# _152_ 0.002283f
C12341 FILLER_0_9_28/a_1916_375# _054_ 0.005889f
C12342 _093_ FILLER_0_18_61/a_36_472# 0.004039f
C12343 net55 FILLER_0_18_37/a_932_472# 0.00769f
C12344 _114_ _311_/a_1920_473# 0.005579f
C12345 trimb[1] net40 0.00126f
C12346 _045_ mask\[1\] 0.024178f
C12347 net50 _447_/a_2665_112# 0.015374f
C12348 FILLER_0_17_72/a_2812_375# vdd 0.005986f
C12349 _069_ _429_/a_1000_472# 0.029501f
C12350 _376_/a_36_160# vdd -0.006711f
C12351 output35/a_224_472# net21 0.069263f
C12352 _142_ net53 0.001961f
C12353 _093_ FILLER_0_17_104/a_1468_375# 0.010965f
C12354 _432_/a_448_472# _139_ 0.001772f
C12355 net52 _029_ 0.03261f
C12356 net74 _070_ 0.394108f
C12357 _321_/a_3126_472# _176_ 0.001932f
C12358 _069_ _395_/a_1492_488# 0.002565f
C12359 FILLER_0_3_142/a_36_472# _370_/a_848_380# 0.001207f
C12360 net82 _443_/a_1204_472# 0.004056f
C12361 _095_ FILLER_0_14_107/a_484_472# 0.014431f
C12362 _083_ _263_/a_224_472# 0.003191f
C12363 net78 _109_ 0.001432f
C12364 net60 _109_ 0.021502f
C12365 _132_ _098_ 0.038463f
C12366 _053_ net57 0.037224f
C12367 net44 FILLER_0_15_2/a_572_375# 0.041552f
C12368 FILLER_0_22_86/a_1468_375# vdd 0.035441f
C12369 _192_/a_67_603# mask\[1\] 0.020097f
C12370 net39 net47 0.13057f
C12371 net33 _434_/a_36_151# 0.002776f
C12372 _131_ FILLER_0_17_56/a_124_375# 0.001609f
C12373 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_36_472# 0.001723f
C12374 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_572_375# 0.026339f
C12375 FILLER_0_12_2/a_36_472# net44 0.011079f
C12376 _128_ _090_ 0.018296f
C12377 _178_ FILLER_0_14_50/a_36_472# 0.001492f
C12378 FILLER_0_7_59/a_572_375# net67 0.007538f
C12379 _071_ FILLER_0_13_142/a_1380_472# 0.001617f
C12380 FILLER_0_24_130/a_124_375# output24/a_224_472# 0.00515f
C12381 net14 _156_ 0.184287f
C12382 FILLER_0_3_204/a_124_375# net65 0.003831f
C12383 net79 _094_ 0.301878f
C12384 _300_/a_224_472# vdd 0.001344f
C12385 mask\[8\] _437_/a_2248_156# 0.004415f
C12386 _422_/a_2248_156# _009_ 0.061786f
C12387 _417_/a_2665_112# vss 0.002571f
C12388 _417_/a_2560_156# vdd 0.001658f
C12389 _065_ net66 0.003956f
C12390 _449_/a_448_472# net15 0.040076f
C12391 FILLER_0_10_37/a_124_375# _173_ 0.00262f
C12392 _095_ _452_/a_36_151# 0.002974f
C12393 _074_ FILLER_0_3_172/a_484_472# 0.001763f
C12394 FILLER_0_9_142/a_36_472# vss 0.004305f
C12395 _043_ net40 0.031043f
C12396 _389_/a_36_148# _172_ 0.039684f
C12397 _239_/a_36_160# net68 0.043367f
C12398 net13 _170_ 0.001668f
C12399 _258_/a_36_160# net59 0.003167f
C12400 state\[2\] vdd 0.392508f
C12401 FILLER_0_15_142/a_484_472# net23 0.002884f
C12402 _411_/a_1204_472# net8 0.001768f
C12403 FILLER_0_5_172/a_124_375# net22 0.002388f
C12404 _178_ cal_count\[3\] 0.002061f
C12405 ctln[3] output11/a_224_472# 0.068614f
C12406 FILLER_0_11_101/a_124_375# cal_count\[3\] 0.00419f
C12407 _176_ _394_/a_728_93# 0.002001f
C12408 net60 _421_/a_2248_156# 0.036944f
C12409 _128_ net22 0.03249f
C12410 _290_/a_224_472# _094_ 0.003006f
C12411 _045_ vss 0.032891f
C12412 _437_/a_2665_112# vdd 0.050182f
C12413 _185_ net40 0.048742f
C12414 _444_/a_36_151# net67 0.055072f
C12415 _373_/a_1254_68# _090_ 0.001326f
C12416 _131_ _125_ 0.013932f
C12417 net57 _428_/a_1000_472# 0.024803f
C12418 _420_/a_2248_156# _108_ 0.021735f
C12419 FILLER_0_4_213/a_484_472# vss 0.007857f
C12420 _086_ _081_ 0.033115f
C12421 fanout59/a_36_160# vdd 0.02169f
C12422 _083_ _265_/a_224_472# 0.003404f
C12423 net34 _207_/a_67_603# 0.008585f
C12424 net47 FILLER_0_5_148/a_484_472# 0.009741f
C12425 _192_/a_67_603# vss 0.007021f
C12426 trim_mask\[4\] vdd 0.20602f
C12427 _028_ FILLER_0_7_104/a_572_375# 0.003664f
C12428 _086_ FILLER_0_7_104/a_932_472# 0.001786f
C12429 _119_ FILLER_0_7_104/a_1380_472# 0.002603f
C12430 net34 _435_/a_36_151# 0.011954f
C12431 state\[0\] _090_ 0.003121f
C12432 _301_/a_36_472# net35 0.051887f
C12433 _074_ cal_itt\[0\] 0.076802f
C12434 FILLER_0_23_44/a_1380_472# vss 0.003905f
C12435 net54 _433_/a_2560_156# 0.014333f
C12436 vdd FILLER_0_4_91/a_124_375# 0.019812f
C12437 net28 net62 0.05491f
C12438 _115_ _315_/a_244_497# 0.00153f
C12439 fanout71/a_36_113# vdd 0.028178f
C12440 FILLER_0_5_128/a_36_472# _133_ 0.001217f
C12441 _110_ _012_ 0.046196f
C12442 FILLER_0_11_78/a_36_472# vdd -0.001328f
C12443 FILLER_0_11_78/a_572_375# vss 0.004808f
C12444 _432_/a_36_151# FILLER_0_17_161/a_36_472# 0.004847f
C12445 net31 FILLER_0_18_209/a_572_375# 0.001813f
C12446 _166_ _034_ 0.001936f
C12447 _141_ FILLER_0_16_154/a_1020_375# 0.003441f
C12448 mask\[3\] FILLER_0_16_154/a_484_472# 0.002067f
C12449 net20 FILLER_0_8_239/a_36_472# 0.004483f
C12450 net58 FILLER_0_9_290/a_36_472# 0.005553f
C12451 _444_/a_448_472# _054_ 0.017318f
C12452 _174_ _131_ 0.002314f
C12453 _416_/a_2248_156# net62 0.043158f
C12454 FILLER_0_12_50/a_36_472# vss 0.0027f
C12455 _415_/a_448_472# net79 0.001602f
C12456 net43 vdd 0.210686f
C12457 FILLER_0_21_133/a_124_375# mask\[7\] 0.00145f
C12458 trim_val\[4\] _443_/a_2560_156# 0.049334f
C12459 _448_/a_2560_156# trim_mask\[4\] 0.001306f
C12460 FILLER_0_7_104/a_932_472# _154_ 0.002023f
C12461 sample net64 0.209777f
C12462 output33/a_224_472# net18 0.110644f
C12463 _423_/a_448_472# _012_ 0.038928f
C12464 net65 _411_/a_1000_472# 0.001916f
C12465 _028_ FILLER_0_5_72/a_1380_472# 0.002164f
C12466 _422_/a_796_472# _108_ 0.007356f
C12467 _430_/a_36_151# net36 0.003701f
C12468 result[9] vdd 0.597071f
C12469 _077_ _439_/a_2665_112# 0.035688f
C12470 _031_ _369_/a_692_472# 0.00359f
C12471 FILLER_0_4_152/a_36_472# trim_mask\[4\] 0.011746f
C12472 _069_ FILLER_0_15_205/a_124_375# 0.002728f
C12473 FILLER_0_3_172/a_2276_472# net22 0.012151f
C12474 net65 calibrate 0.012434f
C12475 _307_/a_672_472# _096_ 0.001367f
C12476 _427_/a_2248_156# _043_ 0.001148f
C12477 _081_ _169_ 0.260462f
C12478 FILLER_0_4_144/a_572_375# net23 0.019114f
C12479 output42/a_224_472# _221_/a_36_160# 0.017421f
C12480 FILLER_0_10_256/a_36_472# vss 0.001792f
C12481 net49 _160_ 1.243817f
C12482 _074_ FILLER_0_6_177/a_484_472# 0.002068f
C12483 mask\[7\] net21 0.050718f
C12484 FILLER_0_23_282/a_36_472# vdd 0.106034f
C12485 FILLER_0_23_282/a_572_375# vss 0.058599f
C12486 _430_/a_2665_112# _092_ 0.004778f
C12487 _069_ _098_ 0.029447f
C12488 _424_/a_1204_472# _012_ 0.003572f
C12489 net59 net21 0.157689f
C12490 net68 _160_ 0.072339f
C12491 _057_ state\[2\] 0.054838f
C12492 FILLER_0_7_72/a_1020_375# vss 0.004851f
C12493 FILLER_0_7_72/a_1468_375# vdd 0.001135f
C12494 ctln[1] net20 0.135151f
C12495 _077_ calibrate 0.055446f
C12496 _432_/a_1308_423# _137_ 0.002078f
C12497 _128_ _076_ 0.04562f
C12498 ctln[3] _411_/a_2665_112# 0.003037f
C12499 fanout69/a_36_113# vdd 0.00378f
C12500 _445_/a_796_472# _034_ 0.009261f
C12501 net35 FILLER_0_22_177/a_36_472# 0.005721f
C12502 FILLER_0_22_86/a_484_472# net71 0.00583f
C12503 output38/a_224_472# net17 0.04454f
C12504 FILLER_0_2_93/a_484_472# vdd 0.005163f
C12505 net44 _067_ 0.001203f
C12506 _136_ _097_ 0.002577f
C12507 _002_ FILLER_0_3_172/a_2812_375# 0.006403f
C12508 _119_ _070_ 1.949038f
C12509 _052_ FILLER_0_21_28/a_1916_375# 0.002388f
C12510 FILLER_0_12_2/a_572_375# _450_/a_36_151# 0.001597f
C12511 FILLER_0_10_78/a_1468_375# _115_ 0.032403f
C12512 FILLER_0_10_78/a_1380_472# _114_ 0.011079f
C12513 _144_ FILLER_0_19_155/a_572_375# 0.003611f
C12514 _067_ _171_ 0.007069f
C12515 FILLER_0_21_28/a_572_375# net17 0.001455f
C12516 _437_/a_448_472# net14 0.090442f
C12517 FILLER_0_16_255/a_36_472# net19 0.001273f
C12518 _448_/a_2248_156# vdd 0.008296f
C12519 trim_val\[4\] _037_ 0.258184f
C12520 _001_ cal_itt\[1\] 0.057933f
C12521 _132_ _131_ 0.444097f
C12522 fanout68/a_36_113# net50 0.020067f
C12523 FILLER_0_13_212/a_1020_375# _043_ 0.01418f
C12524 _072_ _395_/a_244_68# 0.001406f
C12525 _178_ _278_/a_36_160# 0.269109f
C12526 _087_ FILLER_0_3_172/a_1828_472# 0.027954f
C12527 FILLER_0_11_142/a_572_375# _076_ 0.031784f
C12528 _102_ mask\[2\] 0.036292f
C12529 result[7] net77 0.005269f
C12530 _431_/a_2560_156# _137_ 0.002967f
C12531 FILLER_0_14_107/a_484_472# vss -0.001894f
C12532 FILLER_0_14_107/a_932_472# vdd 0.006908f
C12533 _104_ output19/a_224_472# 0.064818f
C12534 sample vss 0.276162f
C12535 FILLER_0_22_177/a_484_472# vss -0.001894f
C12536 FILLER_0_22_177/a_932_472# vdd 0.029547f
C12537 _030_ net49 0.046089f
C12538 fanout57/a_36_113# net57 0.004316f
C12539 _115_ FILLER_0_9_72/a_1380_472# 0.007262f
C12540 _043_ FILLER_0_13_80/a_124_375# 0.013485f
C12541 _053_ _372_/a_2034_472# 0.00181f
C12542 FILLER_0_22_177/a_124_375# _435_/a_36_151# 0.059049f
C12543 net69 _441_/a_2560_156# 0.002904f
C12544 _053_ _129_ 0.003479f
C12545 _126_ _125_ 0.032402f
C12546 _087_ net37 0.23484f
C12547 net31 net30 0.130396f
C12548 _439_/a_36_151# _453_/a_2665_112# 0.001738f
C12549 _130_ _125_ 0.002745f
C12550 net63 _069_ 0.04528f
C12551 FILLER_0_5_109/a_484_472# vss 0.00212f
C12552 _036_ net66 0.04474f
C12553 net68 _030_ 0.007737f
C12554 cal_itt\[2\] FILLER_0_3_221/a_932_472# 0.016327f
C12555 FILLER_0_12_220/a_1380_472# FILLER_0_12_236/a_36_472# 0.013277f
C12556 FILLER_0_5_72/a_124_375# FILLER_0_5_54/a_1468_375# 0.005439f
C12557 _132_ _114_ 0.08562f
C12558 output12/a_224_472# FILLER_0_0_198/a_124_375# 0.00515f
C12559 FILLER_0_5_109/a_36_472# _365_/a_36_68# 0.07596f
C12560 _077_ FILLER_0_6_231/a_36_472# 0.075292f
C12561 net50 _444_/a_2560_156# 0.001479f
C12562 result[7] _102_ 0.010818f
C12563 _432_/a_36_151# net57 0.00484f
C12564 _429_/a_36_151# FILLER_0_15_212/a_572_375# 0.059049f
C12565 net34 FILLER_0_22_128/a_3260_375# 0.006974f
C12566 _436_/a_2560_156# net54 0.010748f
C12567 _452_/a_36_151# vss 0.02741f
C12568 _452_/a_448_472# vdd 0.019824f
C12569 _448_/a_36_151# net76 0.03831f
C12570 _016_ _428_/a_1308_423# 0.00107f
C12571 result[8] _422_/a_1308_423# 0.001356f
C12572 FILLER_0_22_86/a_1020_375# _026_ 0.001032f
C12573 mask\[4\] _433_/a_2248_156# 0.001082f
C12574 net20 FILLER_0_12_220/a_484_472# 0.001758f
C12575 output29/a_224_472# _094_ 0.006731f
C12576 net52 FILLER_0_5_72/a_36_472# 0.014911f
C12577 _176_ _067_ 0.046599f
C12578 _450_/a_2225_156# net6 0.001143f
C12579 _432_/a_448_472# _098_ 0.032293f
C12580 output37/a_224_472# net76 0.004028f
C12581 _308_/a_692_472# _115_ 0.001485f
C12582 mask\[0\] _429_/a_36_151# 0.026729f
C12583 FILLER_0_0_130/a_124_375# _442_/a_36_151# 0.059049f
C12584 output48/a_224_472# valid 0.046397f
C12585 _079_ _084_ 0.046584f
C12586 net35 FILLER_0_23_88/a_36_472# 0.00675f
C12587 FILLER_0_16_73/a_572_375# net55 0.015207f
C12588 net42 net47 0.237866f
C12589 _048_ vdd 0.270091f
C12590 FILLER_0_12_136/a_1380_472# cal_count\[3\] 0.00383f
C12591 FILLER_0_18_177/a_484_472# vdd 0.006177f
C12592 FILLER_0_18_177/a_36_472# vss 0.002187f
C12593 FILLER_0_20_177/a_124_375# _098_ 0.018701f
C12594 _428_/a_1204_472# _131_ 0.012968f
C12595 _093_ FILLER_0_18_107/a_932_472# 0.008683f
C12596 net9 vss 0.086497f
C12597 output24/a_224_472# vss 0.004078f
C12598 _418_/a_2560_156# vdd 0.001506f
C12599 _418_/a_2665_112# vss 0.003519f
C12600 _413_/a_36_151# FILLER_0_2_177/a_572_375# 0.073306f
C12601 _255_/a_224_552# vss 0.001019f
C12602 FILLER_0_5_128/a_124_375# vdd 0.008803f
C12603 FILLER_0_9_60/a_36_472# net51 0.059421f
C12604 _073_ _082_ 0.009987f
C12605 _068_ net37 0.006392f
C12606 FILLER_0_9_223/a_484_472# _426_/a_2665_112# 0.004209f
C12607 _450_/a_2449_156# net40 0.010265f
C12608 _155_ FILLER_0_6_90/a_484_472# 0.005297f
C12609 _198_/a_67_603# mask\[2\] 0.005143f
C12610 _141_ _340_/a_36_160# 0.00584f
C12611 _149_ _437_/a_2560_156# 0.008064f
C12612 _053_ FILLER_0_5_54/a_36_472# 0.003309f
C12613 net75 _425_/a_448_472# 0.038993f
C12614 output17/a_224_472# net43 0.006661f
C12615 FILLER_0_16_57/a_124_375# vss 0.001678f
C12616 FILLER_0_16_57/a_572_375# vdd 0.004039f
C12617 _440_/a_36_151# FILLER_0_6_47/a_2276_472# 0.001512f
C12618 FILLER_0_3_2/a_124_375# _446_/a_36_151# 0.023595f
C12619 FILLER_0_9_223/a_484_472# _060_ 0.001529f
C12620 FILLER_0_17_56/a_484_472# FILLER_0_18_61/a_36_472# 0.026657f
C12621 _077_ _125_ 0.017422f
C12622 FILLER_0_12_28/a_36_472# vdd 0.095598f
C12623 FILLER_0_12_28/a_124_375# vss 0.013117f
C12624 result[8] net22 0.278936f
C12625 _432_/a_448_472# net63 0.002757f
C12626 net81 _139_ 0.001762f
C12627 FILLER_0_13_142/a_1380_472# net23 0.026285f
C12628 net79 _043_ 0.393702f
C12629 _072_ _311_/a_3220_473# 0.001995f
C12630 _414_/a_36_151# cal_itt\[3\] 0.049033f
C12631 FILLER_0_5_198/a_124_375# net21 0.029659f
C12632 FILLER_0_21_150/a_36_472# _146_ 0.00236f
C12633 net71 vdd 0.775031f
C12634 _441_/a_1308_423# _168_ 0.044302f
C12635 mask\[3\] mask\[2\] 0.077703f
C12636 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_484_472# 0.026657f
C12637 _189_/a_67_603# net27 0.008028f
C12638 net65 output9/a_224_472# 0.095296f
C12639 net41 _408_/a_728_93# 0.058816f
C12640 FILLER_0_5_72/a_1468_375# _164_ 0.040819f
C12641 FILLER_0_14_50/a_36_472# FILLER_0_12_50/a_124_375# 0.0027f
C12642 FILLER_0_1_204/a_36_472# net11 0.014707f
C12643 net75 _253_/a_36_68# 0.047906f
C12644 _099_ _195_/a_67_603# 0.065049f
C12645 _339_/a_36_160# FILLER_0_19_155/a_572_375# 0.003589f
C12646 _431_/a_2560_156# net56 0.001258f
C12647 cal_count\[3\] FILLER_0_11_78/a_124_375# 0.019818f
C12648 FILLER_0_24_290/a_124_375# vdd 0.026739f
C12649 vdd FILLER_0_13_290/a_124_375# 0.031436f
C12650 net57 _072_ 0.108982f
C12651 _098_ FILLER_0_15_235/a_36_472# 0.093007f
C12652 _132_ _126_ 0.247838f
C12653 FILLER_0_3_142/a_36_472# _261_/a_36_160# 0.001542f
C12654 _033_ net40 0.298492f
C12655 _098_ _438_/a_36_151# 0.009083f
C12656 cal_count\[3\] FILLER_0_12_50/a_124_375# 0.060164f
C12657 net76 FILLER_0_5_212/a_36_472# 0.00377f
C12658 net80 FILLER_0_19_171/a_124_375# 0.024758f
C12659 _053_ _219_/a_36_160# 0.005244f
C12660 _389_/a_36_148# FILLER_0_10_94/a_36_472# 0.001723f
C12661 _176_ _121_ 0.035608f
C12662 net55 _052_ 0.095046f
C12663 _136_ _019_ 0.049263f
C12664 FILLER_0_6_47/a_2276_472# vdd 0.002735f
C12665 FILLER_0_6_47/a_1828_472# vss 0.003457f
C12666 _429_/a_1000_472# net22 0.007429f
C12667 net75 FILLER_0_8_247/a_124_375# 0.002085f
C12668 _021_ _137_ 0.002807f
C12669 _093_ FILLER_0_17_72/a_2812_375# 0.019521f
C12670 net72 net17 0.004503f
C12671 net79 net21 0.645949f
C12672 result[5] net20 0.045364f
C12673 _201_/a_67_603# _047_ 0.013357f
C12674 FILLER_0_11_142/a_124_375# vdd 0.010672f
C12675 _114_ _069_ 0.029875f
C12676 _228_/a_36_68# _060_ 0.016962f
C12677 vss _039_ 0.180364f
C12678 _425_/a_36_151# FILLER_0_8_247/a_36_472# 0.02628f
C12679 _425_/a_1308_423# FILLER_0_8_247/a_1020_375# 0.001064f
C12680 net81 _429_/a_1000_472# 0.011018f
C12681 _131_ FILLER_0_18_37/a_1468_375# 0.001151f
C12682 _013_ vdd 0.372605f
C12683 net27 FILLER_0_14_235/a_124_375# 0.002299f
C12684 FILLER_0_4_197/a_1380_472# net22 0.012286f
C12685 FILLER_0_21_142/a_484_472# FILLER_0_21_150/a_36_472# 0.013277f
C12686 net63 FILLER_0_19_171/a_1020_375# 0.004794f
C12687 net38 output39/a_224_472# 0.036027f
C12688 net82 FILLER_0_3_221/a_572_375# 0.005424f
C12689 _077_ FILLER_0_10_78/a_1380_472# 0.001548f
C12690 _132_ FILLER_0_15_116/a_572_375# 0.003964f
C12691 FILLER_0_21_125/a_572_375# net54 0.024701f
C12692 _086_ FILLER_0_11_135/a_36_472# 0.004074f
C12693 _074_ FILLER_0_6_231/a_124_375# 0.006087f
C12694 _422_/a_2665_112# mask\[7\] 0.028271f
C12695 result[9] net60 0.251903f
C12696 result[9] net78 0.015761f
C12697 _367_/a_36_68# vdd 0.010246f
C12698 ctln[1] _073_ 0.001457f
C12699 _066_ vdd 0.14893f
C12700 _426_/a_2665_112# calibrate 0.004837f
C12701 cal_count\[3\] FILLER_0_11_109/a_36_472# 0.00702f
C12702 ctlp[9] vss 0.013018f
C12703 net1 _082_ 0.033169f
C12704 net61 vdd 0.46584f
C12705 _140_ FILLER_0_22_128/a_124_375# 0.011452f
C12706 output46/a_224_472# FILLER_0_20_2/a_572_375# 0.03228f
C12707 _136_ FILLER_0_17_142/a_572_375# 0.001371f
C12708 cal_count\[3\] FILLER_0_11_135/a_36_472# 0.005101f
C12709 net82 net22 1.960347f
C12710 _002_ FILLER_0_4_197/a_124_375# 0.001406f
C12711 _402_/a_1948_68# cal_count\[1\] 0.037053f
C12712 net57 FILLER_0_13_142/a_1468_375# 0.011369f
C12713 net57 fanout53/a_36_160# 0.009946f
C12714 _428_/a_1308_423# _043_ 0.024052f
C12715 trim[0] vdd 0.125774f
C12716 _415_/a_2560_156# result[1] 0.002282f
C12717 _086_ _161_ 0.077837f
C12718 FILLER_0_8_138/a_124_375# _077_ 0.007238f
C12719 _430_/a_2248_156# net63 0.051057f
C12720 FILLER_0_4_197/a_36_472# _088_ 0.067725f
C12721 net81 net82 0.063498f
C12722 FILLER_0_6_239/a_124_375# FILLER_0_6_231/a_572_375# 0.012001f
C12723 FILLER_0_12_20/a_484_472# net47 0.020293f
C12724 fanout71/a_36_113# _433_/a_36_151# 0.138322f
C12725 _070_ _389_/a_36_148# 0.010534f
C12726 FILLER_0_21_28/a_2812_375# vdd -0.014642f
C12727 _111_ net15 0.049514f
C12728 _052_ _424_/a_796_472# 0.002115f
C12729 FILLER_0_3_172/a_1828_472# vdd 0.0083f
C12730 net23 mask\[6\] 0.025699f
C12731 _442_/a_448_472# FILLER_0_2_127/a_36_472# 0.008634f
C12732 FILLER_0_8_2/a_124_375# vdd 0.016103f
C12733 _449_/a_2560_156# net55 0.004835f
C12734 net4 FILLER_0_3_221/a_932_472# 0.002116f
C12735 vss FILLER_0_8_156/a_36_472# 0.00168f
C12736 vdd FILLER_0_8_156/a_484_472# 0.007249f
C12737 result[1] _005_ 0.001478f
C12738 _438_/a_2560_156# net14 0.049389f
C12739 FILLER_0_5_54/a_36_472# _164_ 0.003923f
C12740 result[6] _421_/a_448_472# 0.038671f
C12741 _161_ cal_count\[3\] 0.047389f
C12742 output43/a_224_472# output45/a_224_472# 0.246888f
C12743 net37 vdd 0.544653f
C12744 _020_ FILLER_0_18_107/a_2364_375# 0.003755f
C12745 _001_ net59 0.001439f
C12746 FILLER_0_11_101/a_124_375# _120_ 0.008016f
C12747 net55 FILLER_0_17_72/a_932_472# 0.024922f
C12748 net81 FILLER_0_14_235/a_484_472# 0.015266f
C12749 FILLER_0_18_2/a_2812_375# net17 0.012909f
C12750 FILLER_0_4_107/a_1468_375# trim_mask\[4\] 0.00157f
C12751 _112_ _425_/a_36_151# 0.032941f
C12752 net68 net67 0.147318f
C12753 _144_ _433_/a_1000_472# 0.029564f
C12754 _115_ _171_ 0.033359f
C12755 ctln[7] FILLER_0_0_96/a_36_472# 0.01317f
C12756 FILLER_0_16_37/a_36_472# net72 0.005134f
C12757 FILLER_0_5_109/a_124_375# _153_ 0.040726f
C12758 FILLER_0_5_109/a_36_472# _154_ 0.070958f
C12759 FILLER_0_10_78/a_124_375# _453_/a_2665_112# 0.006271f
C12760 _005_ _416_/a_2560_156# 0.004273f
C12761 net70 net36 0.066607f
C12762 _443_/a_2248_156# _170_ 0.068179f
C12763 _061_ _113_ 0.012561f
C12764 _132_ FILLER_0_17_104/a_932_472# 0.006091f
C12765 net1 _265_/a_244_68# 0.023821f
C12766 _108_ vdd 0.298249f
C12767 trim_val\[4\] FILLER_0_3_172/a_572_375# 0.001076f
C12768 output48/a_224_472# net59 0.039277f
C12769 _131_ FILLER_0_17_104/a_36_472# 0.004125f
C12770 _426_/a_36_151# FILLER_0_8_247/a_124_375# 0.059049f
C12771 _118_ _122_ 0.046796f
C12772 net41 FILLER_0_17_38/a_124_375# 0.001109f
C12773 FILLER_0_9_72/a_36_472# _453_/a_2665_112# 0.001167f
C12774 _084_ vss 0.082779f
C12775 _140_ _149_ 0.0088f
C12776 _175_ FILLER_0_15_72/a_124_375# 0.009573f
C12777 _112_ net1 0.001653f
C12778 _132_ _137_ 0.023462f
C12779 _412_/a_2248_156# net18 0.05155f
C12780 net22 _435_/a_2560_156# 0.002281f
C12781 _062_ _311_/a_692_473# 0.008632f
C12782 FILLER_0_5_109/a_572_375# _163_ 0.003096f
C12783 FILLER_0_10_37/a_124_375# net68 0.012617f
C12784 _087_ _122_ 0.007241f
C12785 FILLER_0_0_266/a_124_375# vdd 0.006328f
C12786 _162_ _163_ 0.011497f
C12787 _014_ _123_ 0.050082f
C12788 _115_ _176_ 1.300336f
C12789 _179_ vdd 0.049022f
C12790 _431_/a_2248_156# net73 0.003228f
C12791 FILLER_0_15_205/a_124_375# net22 0.049201f
C12792 FILLER_0_12_28/a_36_472# cal_count\[0\] 0.001662f
C12793 mask\[3\] FILLER_0_18_177/a_2364_375# 0.002935f
C12794 net16 _063_ 0.038576f
C12795 FILLER_0_8_247/a_124_375# FILLER_0_8_239/a_124_375# 0.003732f
C12796 _187_ _408_/a_1936_472# 0.017573f
C12797 net29 result[2] 0.001786f
C12798 FILLER_0_4_107/a_124_375# vss 0.00322f
C12799 FILLER_0_4_107/a_572_375# vdd 0.034678f
C12800 _077_ net50 0.312283f
C12801 net54 FILLER_0_18_107/a_3260_375# 0.001619f
C12802 _103_ _418_/a_2665_112# 0.0066f
C12803 _091_ _429_/a_2665_112# 0.002597f
C12804 net70 FILLER_0_14_123/a_124_375# 0.032077f
C12805 net20 net19 0.384932f
C12806 net60 _418_/a_2560_156# 0.020147f
C12807 _098_ net22 0.157058f
C12808 FILLER_0_5_117/a_124_375# FILLER_0_5_109/a_572_375# 0.012001f
C12809 ctln[1] net1 0.003756f
C12810 output20/a_224_472# result[8] 0.038114f
C12811 net81 FILLER_0_15_205/a_124_375# 0.015134f
C12812 _207_/a_67_603# _146_ 0.026192f
C12813 net33 mask\[6\] 0.881813f
C12814 _061_ _118_ 0.268815f
C12815 _436_/a_36_151# _437_/a_2665_112# 0.001466f
C12816 mask\[5\] _434_/a_2665_112# 0.003849f
C12817 output46/a_224_472# FILLER_0_21_28/a_124_375# 0.003337f
C12818 net68 FILLER_0_8_37/a_572_375# 0.011704f
C12819 net81 _098_ 0.029506f
C12820 FILLER_0_3_54/a_36_472# _381_/a_36_472# 0.010679f
C12821 net47 _160_ 0.2966f
C12822 _397_/a_36_472# _175_ 0.004667f
C12823 _289_/a_36_472# _102_ 0.046918f
C12824 _432_/a_2665_112# _091_ 0.002978f
C12825 _086_ _127_ 0.042698f
C12826 FILLER_0_7_162/a_36_472# _062_ 0.016683f
C12827 _132_ FILLER_0_19_125/a_36_472# 0.008568f
C12828 net28 _192_/a_255_603# 0.003166f
C12829 FILLER_0_2_93/a_484_472# FILLER_0_2_101/a_36_472# 0.013277f
C12830 net48 net76 0.069349f
C12831 FILLER_0_11_78/a_572_375# _389_/a_36_148# 0.021545f
C12832 output36/a_224_472# net36 0.009109f
C12833 output21/a_224_472# net21 0.011791f
C12834 _401_/a_36_68# _180_ 0.051459f
C12835 _028_ FILLER_0_6_47/a_2812_375# 0.023189f
C12836 net54 _354_/a_257_69# 0.001135f
C12837 _068_ _122_ 0.096251f
C12838 _127_ cal_count\[3\] 0.306114f
C12839 _192_/a_67_603# _416_/a_2665_112# 0.012638f
C12840 _044_ _416_/a_36_151# 0.032206f
C12841 FILLER_0_7_195/a_124_375# _055_ 0.001597f
C12842 net63 net22 0.223664f
C12843 _449_/a_448_472# _067_ 0.0432f
C12844 cal_itt\[3\] net21 0.175781f
C12845 _189_/a_255_603# net64 0.002455f
C12846 result[8] FILLER_0_23_282/a_484_472# 0.001908f
C12847 FILLER_0_5_109/a_572_375# FILLER_0_4_107/a_932_472# 0.001684f
C12848 net15 FILLER_0_13_72/a_36_472# 0.006713f
C12849 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_484_472# 0.001963f
C12850 _033_ _444_/a_796_472# 0.0099f
C12851 _165_ _444_/a_2248_156# 0.006027f
C12852 _053_ FILLER_0_6_47/a_1020_375# 0.015621f
C12853 net36 _282_/a_36_160# 0.002754f
C12854 _068_ _311_/a_2180_473# 0.001454f
C12855 net76 FILLER_0_6_177/a_124_375# 0.00227f
C12856 _092_ vdd 0.140213f
C12857 _143_ net80 0.023487f
C12858 net2 net37 0.05083f
C12859 FILLER_0_14_81/a_36_472# net55 0.015878f
C12860 _370_/a_124_24# _152_ 0.069015f
C12861 _370_/a_848_380# _081_ 0.035068f
C12862 _020_ net70 0.014391f
C12863 FILLER_0_16_57/a_1020_375# FILLER_0_17_64/a_124_375# 0.026339f
C12864 state\[0\] _128_ 0.228492f
C12865 _086_ _071_ 0.041029f
C12866 FILLER_0_0_198/a_36_472# vdd 0.052226f
C12867 FILLER_0_0_198/a_124_375# vss 0.017602f
C12868 en_co_clk vdd 0.245319f
C12869 FILLER_0_9_223/a_484_472# vss 0.006102f
C12870 cal_count\[3\] _373_/a_438_68# 0.003743f
C12871 _451_/a_836_156# net14 0.00174f
C12872 _104_ output18/a_224_472# 0.08426f
C12873 net50 net69 0.634381f
C12874 net52 _031_ 0.633473f
C12875 FILLER_0_3_204/a_36_472# vdd 0.092654f
C12876 FILLER_0_3_204/a_124_375# vss 0.017795f
C12877 _011_ mask\[7\] 0.043474f
C12878 _143_ FILLER_0_18_139/a_1468_375# 0.001097f
C12879 output28/a_224_472# vss -0.0033f
C12880 _061_ _068_ 1.857322f
C12881 _110_ vdd 0.041979f
C12882 net18 _419_/a_1308_423# 0.013637f
C12883 _289_/a_36_472# _198_/a_67_603# 0.027695f
C12884 FILLER_0_1_192/a_124_375# net59 0.014491f
C12885 _443_/a_1204_472# net69 0.002642f
C12886 cal_count\[3\] _071_ 0.214649f
C12887 result[5] result[4] 0.090472f
C12888 _142_ net23 0.037306f
C12889 net20 _009_ 0.026064f
C12890 net80 _136_ 0.034194f
C12891 FILLER_0_5_172/a_36_472# net37 0.013857f
C12892 net45 net26 0.002978f
C12893 FILLER_0_14_99/a_36_472# FILLER_0_13_100/a_36_472# 0.026657f
C12894 _144_ mask\[5\] 0.38642f
C12895 vss _416_/a_796_472# 0.001468f
C12896 net35 net23 0.04007f
C12897 net71 _433_/a_36_151# 0.014126f
C12898 _134_ net14 0.001303f
C12899 net27 FILLER_0_9_282/a_572_375# 0.002809f
C12900 _178_ _408_/a_56_524# 0.014421f
C12901 _367_/a_244_472# _154_ 0.001775f
C12902 net64 FILLER_0_14_235/a_572_375# 0.008689f
C12903 _429_/a_1308_423# vss 0.008906f
C12904 _119_ FILLER_0_8_156/a_36_472# 0.010504f
C12905 vss clkc 0.0311f
C12906 _423_/a_36_151# vss 0.012999f
C12907 _423_/a_448_472# vdd 0.01351f
C12908 FILLER_0_4_49/a_484_472# FILLER_0_3_54/a_36_472# 0.026657f
C12909 net38 cal_count\[3\] 0.002225f
C12910 _079_ FILLER_0_5_198/a_484_472# 0.008167f
C12911 _335_/a_257_69# _043_ 0.001043f
C12912 _075_ _077_ 0.004518f
C12913 _414_/a_36_151# _081_ 0.016708f
C12914 FILLER_0_10_256/a_36_472# FILLER_0_10_247/a_36_472# 0.001963f
C12915 mask\[3\] _289_/a_36_472# 0.02347f
C12916 output31/a_224_472# vdd 0.083516f
C12917 net64 calibrate 0.096329f
C12918 FILLER_0_9_142/a_124_375# _120_ 0.04442f
C12919 net61 net78 1.588656f
C12920 net61 net60 0.059237f
C12921 FILLER_0_4_197/a_932_472# vdd 0.003395f
C12922 _008_ _419_/a_448_472# 0.01758f
C12923 FILLER_0_15_116/a_36_472# FILLER_0_17_104/a_1468_375# 0.001512f
C12924 net13 vdd 0.264116f
C12925 _070_ FILLER_0_9_105/a_124_375# 0.017687f
C12926 FILLER_0_22_86/a_36_472# _098_ 0.182093f
C12927 FILLER_0_20_107/a_124_375# vss 0.002749f
C12928 FILLER_0_20_107/a_36_472# vdd 0.117841f
C12929 FILLER_0_7_146/a_36_472# _062_ 0.011622f
C12930 _093_ net71 0.133323f
C12931 _424_/a_1204_472# vdd 0.001573f
C12932 FILLER_0_23_290/a_36_472# vss 0.0074f
C12933 _015_ net27 0.103416f
C12934 _444_/a_1308_423# net17 0.028709f
C12935 FILLER_0_22_128/a_3260_375# _146_ 0.004692f
C12936 _441_/a_2560_156# vss 0.001374f
C12937 _064_ vss 0.228443f
C12938 _428_/a_2665_112# FILLER_0_13_142/a_36_472# 0.003706f
C12939 output8/a_224_472# ctln[1] 0.020259f
C12940 net69 trim_mask\[3\] 0.017779f
C12941 _015_ _426_/a_2560_156# 0.024461f
C12942 _228_/a_36_68# vss 0.031389f
C12943 net57 state\[2\] 1.25275f
C12944 _013_ FILLER_0_17_64/a_36_472# 0.001991f
C12945 _447_/a_2248_156# vdd 0.009094f
C12946 net23 FILLER_0_5_148/a_124_375# 0.01836f
C12947 net36 state\[1\] 0.004105f
C12948 _114_ FILLER_0_11_101/a_484_472# 0.025975f
C12949 _114_ _090_ 0.001909f
C12950 _005_ _094_ 0.162984f
C12951 _431_/a_2560_156# vss 0.004767f
C12952 _025_ _352_/a_49_472# 0.003933f
C12953 net34 _208_/a_36_160# 0.002666f
C12954 FILLER_0_9_28/a_572_375# net40 0.001406f
C12955 _446_/a_796_472# _035_ 0.013039f
C12956 result[2] result[3] 0.09741f
C12957 FILLER_0_4_197/a_124_375# net76 0.00811f
C12958 _439_/a_2665_112# vss 0.003954f
C12959 _070_ _370_/a_124_24# 0.00219f
C12960 _412_/a_2665_112# net58 0.006815f
C12961 net35 _025_ 0.02169f
C12962 _431_/a_2248_156# _427_/a_36_151# 0.001081f
C12963 FILLER_0_14_181/a_36_472# _043_ 0.008613f
C12964 fanout66/a_36_113# _160_ 0.015681f
C12965 input4/a_36_68# net59 0.003625f
C12966 _106_ _201_/a_67_603# 0.00327f
C12967 _411_/a_1000_472# vss 0.002964f
C12968 _174_ _095_ 0.977766f
C12969 output13/a_224_472# net12 0.002723f
C12970 _386_/a_692_472# _169_ 0.004014f
C12971 _386_/a_848_380# _163_ 0.026484f
C12972 _098_ _437_/a_2560_156# 0.001174f
C12973 _274_/a_36_68# _060_ 0.02117f
C12974 vss FILLER_0_14_235/a_572_375# 0.017196f
C12975 FILLER_0_21_125/a_484_472# _022_ 0.004649f
C12976 input4/a_36_68# net4 0.004679f
C12977 FILLER_0_11_78/a_124_375# _120_ 0.014367f
C12978 _432_/a_448_472# _137_ 0.008956f
C12979 net57 trim_mask\[4\] 0.259381f
C12980 _359_/a_636_68# _062_ 0.001578f
C12981 net78 _108_ 0.056528f
C12982 net41 _450_/a_2225_156# 0.024042f
C12983 FILLER_0_4_99/a_124_375# net14 0.003714f
C12984 calibrate vss 1.140031f
C12985 _122_ vdd 0.379907f
C12986 _132_ FILLER_0_18_107/a_2276_472# 0.006713f
C12987 _155_ FILLER_0_7_104/a_484_472# 0.003068f
C12988 FILLER_0_11_64/a_36_472# net15 0.020589f
C12989 net35 net33 1.594925f
C12990 _436_/a_448_472# output24/a_224_472# 0.009204f
C12991 FILLER_0_16_57/a_484_472# net55 0.001797f
C12992 fanout51/a_36_113# FILLER_0_11_64/a_36_472# 0.001396f
C12993 FILLER_0_12_50/a_124_375# _120_ 0.002753f
C12994 _004_ net79 0.27387f
C12995 _093_ _013_ 0.064462f
C12996 _164_ FILLER_0_6_47/a_1020_375# 0.004285f
C12997 net50 _165_ 0.056964f
C12998 FILLER_0_17_72/a_3172_472# net14 0.046864f
C12999 _320_/a_1120_472# _043_ 0.002242f
C13000 net32 result[6] 0.048987f
C13001 result[8] FILLER_0_24_290/a_36_472# 0.004676f
C13002 _132_ FILLER_0_16_107/a_572_375# 0.007439f
C13003 fanout66/a_36_113# _030_ 0.038252f
C13004 _311_/a_2180_473# vdd 0.001974f
C13005 input1/a_36_113# vdd 0.099655f
C13006 net53 FILLER_0_16_154/a_124_375# 0.003458f
C13007 FILLER_0_9_28/a_1380_472# net16 0.005297f
C13008 FILLER_0_19_142/a_124_375# _145_ 0.009109f
C13009 ctlp[3] _109_ 0.001371f
C13010 mask\[5\] FILLER_0_18_177/a_2364_375# 0.002726f
C13011 _049_ vdd 0.199608f
C13012 net67 FILLER_0_8_37/a_36_472# 0.001479f
C13013 _346_/a_49_472# _140_ 0.003436f
C13014 mask\[5\] _339_/a_36_160# 0.007734f
C13015 _115_ FILLER_0_10_94/a_124_375# 0.010311f
C13016 _408_/a_1336_472# _186_ 0.010089f
C13017 fanout54/a_36_160# vdd 0.008482f
C13018 FILLER_0_13_142/a_572_375# _043_ 0.009328f
C13019 net32 _421_/a_36_151# 0.008275f
C13020 mask\[2\] FILLER_0_16_154/a_1020_375# 0.020485f
C13021 result[4] net19 0.015095f
C13022 FILLER_0_18_2/a_2724_472# _452_/a_36_151# 0.011733f
C13023 FILLER_0_18_2/a_1828_472# _452_/a_1353_112# 0.001313f
C13024 FILLER_0_18_2/a_36_472# _452_/a_3129_107# 0.035307f
C13025 _430_/a_796_472# net21 0.015066f
C13026 FILLER_0_14_91/a_124_375# _176_ 0.019567f
C13027 net36 FILLER_0_15_212/a_932_472# 0.008239f
C13028 net51 net6 0.142515f
C13029 _435_/a_2665_112# vdd 0.01769f
C13030 _053_ FILLER_0_6_79/a_36_472# 0.001777f
C13031 net27 net18 0.092379f
C13032 _116_ state\[1\] 0.693219f
C13033 _436_/a_36_151# net71 0.03535f
C13034 net34 _210_/a_67_603# 0.01049f
C13035 vss FILLER_0_6_231/a_36_472# 0.0048f
C13036 vdd FILLER_0_6_231/a_484_472# 0.004642f
C13037 net17 FILLER_0_20_15/a_572_375# 0.018398f
C13038 _061_ vdd 0.295557f
C13039 FILLER_0_9_28/a_3172_472# FILLER_0_9_60/a_36_472# 0.013276f
C13040 _069_ _248_/a_36_68# 0.058746f
C13041 _132_ _095_ 0.042874f
C13042 net38 _278_/a_36_160# 0.010587f
C13043 _335_/a_49_472# _138_ 0.005957f
C13044 _414_/a_448_472# _003_ 0.023209f
C13045 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_572_375# 0.086635f
C13046 FILLER_0_4_177/a_484_472# net22 0.006506f
C13047 FILLER_0_11_109/a_36_472# _120_ 0.014554f
C13048 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_484_472# 0.001723f
C13049 FILLER_0_9_28/a_932_472# vdd 0.04397f
C13050 _141_ FILLER_0_21_150/a_36_472# 0.002773f
C13051 output25/a_224_472# _213_/a_67_603# 0.032497f
C13052 ctlp[1] FILLER_0_24_274/a_572_375# 0.002408f
C13053 _451_/a_3129_107# _040_ 0.004116f
C13054 _178_ FILLER_0_17_38/a_572_375# 0.031538f
C13055 FILLER_0_11_135/a_36_472# _120_ 0.012562f
C13056 _258_/a_36_160# _081_ 0.00776f
C13057 _443_/a_2665_112# net22 0.00621f
C13058 net47 _156_ 0.040298f
C13059 FILLER_0_17_56/a_124_375# vss 0.00143f
C13060 FILLER_0_17_56/a_572_375# vdd 0.003489f
C13061 _053_ FILLER_0_8_107/a_36_472# 0.013669f
C13062 FILLER_0_7_59/a_484_472# _439_/a_36_151# 0.001061f
C13063 FILLER_0_11_64/a_36_472# net51 0.009015f
C13064 _126_ FILLER_0_11_101/a_484_472# 0.001488f
C13065 net23 FILLER_0_22_128/a_1468_375# 0.001866f
C13066 _129_ _133_ 0.080636f
C13067 _372_/a_2034_472# _133_ 0.001257f
C13068 _372_/a_170_472# _076_ 0.049892f
C13069 _069_ _060_ 0.538161f
C13070 _126_ _090_ 0.003538f
C13071 FILLER_0_1_98/a_36_472# _238_/a_67_603# 0.02529f
C13072 FILLER_0_8_37/a_484_472# _054_ 0.022621f
C13073 _178_ _043_ 0.130207f
C13074 net25 _051_ 0.090798f
C13075 ctlp[3] _422_/a_448_472# 0.001441f
C13076 FILLER_0_7_104/a_932_472# _151_ 0.002092f
C13077 net55 cal_count\[3\] 0.005157f
C13078 net67 net47 0.126281f
C13079 FILLER_0_13_212/a_484_472# vss 0.002397f
C13080 FILLER_0_6_177/a_484_472# _163_ 0.002256f
C13081 FILLER_0_8_24/a_484_472# FILLER_0_8_37/a_36_472# 0.001963f
C13082 FILLER_0_17_72/a_3260_375# _131_ 0.004986f
C13083 _288_/a_224_472# vdd 0.002071f
C13084 _425_/a_36_151# net19 0.009499f
C13085 _178_ _185_ 0.979797f
C13086 _114_ _076_ 0.088609f
C13087 output47/a_224_472# _185_ 0.001177f
C13088 FILLER_0_17_226/a_124_375# vss 0.025007f
C13089 FILLER_0_17_226/a_36_472# vdd 0.087587f
C13090 ctlp[4] net22 0.257841f
C13091 _196_/a_36_160# net62 0.029171f
C13092 FILLER_0_14_181/a_124_375# _138_ 0.001663f
C13093 FILLER_0_18_139/a_124_375# vdd 0.023256f
C13094 net40 output41/a_224_472# 0.081551f
C13095 _125_ vss 0.149512f
C13096 FILLER_0_22_86/a_1380_472# FILLER_0_22_107/a_36_472# 0.001963f
C13097 _041_ vdd 0.19154f
C13098 net68 trim_val\[1\] 0.006974f
C13099 _021_ vss 0.142648f
C13100 FILLER_0_5_206/a_124_375# net37 0.005485f
C13101 net65 output27/a_224_472# 0.019729f
C13102 FILLER_0_12_2/a_572_375# net38 0.00609f
C13103 ctlp[7] _025_ 0.007483f
C13104 net20 FILLER_0_9_223/a_572_375# 0.03118f
C13105 _132_ FILLER_0_19_111/a_572_375# 0.01675f
C13106 _016_ net53 0.180698f
C13107 _369_/a_36_68# _154_ 0.042308f
C13108 net50 FILLER_0_6_79/a_124_375# 0.004402f
C13109 net66 FILLER_0_3_54/a_36_472# 0.008174f
C13110 _412_/a_36_151# _001_ 0.006762f
C13111 _111_ FILLER_0_18_76/a_36_472# 0.006706f
C13112 FILLER_0_5_72/a_572_375# _440_/a_36_151# 0.035849f
C13113 result[7] FILLER_0_24_274/a_1468_375# 0.006125f
C13114 _181_ vdd 0.209604f
C13115 net79 _044_ 0.013636f
C13116 _086_ net23 0.037804f
C13117 mask\[7\] FILLER_0_22_128/a_2364_375# 0.003632f
C13118 net1 net19 0.024768f
C13119 FILLER_0_5_198/a_484_472# vss 0.001338f
C13120 net74 _125_ 0.071757f
C13121 FILLER_0_16_241/a_36_472# vss 0.004432f
C13122 FILLER_0_15_150/a_36_472# net53 0.016925f
C13123 trim[1] _444_/a_36_151# 0.001391f
C13124 _074_ FILLER_0_5_164/a_484_472# 0.003556f
C13125 _095_ FILLER_0_15_72/a_484_472# 0.002306f
C13126 _412_/a_1204_472# net81 0.003435f
C13127 net16 _444_/a_2560_156# 0.010829f
C13128 net80 FILLER_0_22_177/a_484_472# 0.005297f
C13129 cal_itt\[3\] _062_ 0.009718f
C13130 net35 FILLER_0_22_128/a_1828_472# 0.016187f
C13131 _276_/a_36_160# FILLER_0_18_209/a_484_472# 0.003913f
C13132 mask\[0\] _335_/a_665_69# 0.001711f
C13133 _412_/a_36_151# output48/a_224_472# 0.229574f
C13134 cal_count\[3\] net23 0.045417f
C13135 _065_ net17 0.035195f
C13136 trim_val\[2\] _381_/a_36_472# 0.005253f
C13137 FILLER_0_8_24/a_484_472# net47 0.042018f
C13138 net15 FILLER_0_13_80/a_36_472# 0.001122f
C13139 net20 _429_/a_36_151# 0.002103f
C13140 FILLER_0_19_155/a_36_472# _145_ 0.005521f
C13141 output9/a_224_472# vss 0.007544f
C13142 FILLER_0_11_101/a_572_375# FILLER_0_10_107/a_36_472# 0.001684f
C13143 _013_ _424_/a_2665_112# 0.001222f
C13144 FILLER_0_9_72/a_1380_472# _439_/a_36_151# 0.001723f
C13145 _057_ _061_ 0.030546f
C13146 FILLER_0_18_171/a_124_375# vdd 0.021417f
C13147 net64 FILLER_0_9_282/a_36_472# 0.031302f
C13148 _028_ _439_/a_448_472# 0.017606f
C13149 input1/a_36_113# net2 0.018839f
C13150 trim_mask\[1\] FILLER_0_6_47/a_484_472# 0.022211f
C13151 _174_ vss 0.188373f
C13152 FILLER_0_13_65/a_36_472# _174_ 0.011724f
C13153 result[4] fanout78/a_36_113# 0.001531f
C13154 net67 FILLER_0_9_60/a_124_375# 0.003083f
C13155 net63 FILLER_0_22_177/a_1380_472# 0.062289f
C13156 result[4] fanout60/a_36_160# 0.027276f
C13157 output31/a_224_472# net60 0.216716f
C13158 net65 net22 0.374917f
C13159 _122_ FILLER_0_5_172/a_36_472# 0.003007f
C13160 FILLER_0_22_128/a_2276_472# vss 0.02979f
C13161 FILLER_0_22_128/a_2724_472# vdd 0.005923f
C13162 _140_ _098_ 0.647503f
C13163 FILLER_0_16_89/a_484_472# _451_/a_448_472# 0.059367f
C13164 _052_ FILLER_0_18_37/a_1020_375# 0.001287f
C13165 _444_/a_2248_156# vss 0.001329f
C13166 _444_/a_2665_112# vdd 0.029351f
C13167 net27 net62 0.008623f
C13168 _081_ net21 0.030964f
C13169 trim_mask\[2\] _153_ 0.007934f
C13170 fanout77/a_36_113# _418_/a_36_151# 0.001082f
C13171 _446_/a_1308_423# vdd 0.002346f
C13172 net65 net81 0.083316f
C13173 _081_ _261_/a_36_160# 0.049069f
C13174 FILLER_0_9_28/a_3260_375# net51 0.001597f
C13175 _126_ _038_ 0.031198f
C13176 _421_/a_448_472# _419_/a_2665_112# 0.002393f
C13177 net49 _168_ 0.031157f
C13178 FILLER_0_20_193/a_572_375# _205_/a_36_160# 0.002828f
C13179 _077_ net22 0.049592f
C13180 _174_ net74 0.00916f
C13181 FILLER_0_5_72/a_572_375# vdd -0.00211f
C13182 FILLER_0_5_72/a_124_375# vss 0.041166f
C13183 _119_ calibrate 0.062309f
C13184 FILLER_0_6_79/a_36_472# _164_ 0.008685f
C13185 _452_/a_1040_527# _041_ 0.002066f
C13186 net26 FILLER_0_23_44/a_484_472# 0.003796f
C13187 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3172_472# 0.026657f
C13188 net58 _074_ 0.004651f
C13189 FILLER_0_16_57/a_36_472# FILLER_0_17_56/a_124_375# 0.001723f
C13190 state\[1\] _225_/a_36_160# 0.0535f
C13191 FILLER_0_10_78/a_1380_472# vss 0.002096f
C13192 net23 _169_ 0.00151f
C13193 net25 FILLER_0_23_60/a_36_472# 0.005618f
C13194 FILLER_0_7_72/a_572_375# FILLER_0_5_72/a_484_472# 0.001512f
C13195 _132_ mask\[8\] 0.029292f
C13196 net16 _131_ 0.001308f
C13197 FILLER_0_21_28/a_2276_472# _424_/a_36_151# 0.001723f
C13198 _413_/a_2248_156# net21 0.009186f
C13199 mask\[8\] FILLER_0_22_107/a_484_472# 0.024416f
C13200 net35 FILLER_0_22_107/a_36_472# 0.007196f
C13201 net76 _080_ 0.03728f
C13202 _274_/a_36_68# net64 0.036017f
C13203 _092_ _093_ 0.287983f
C13204 _127_ _120_ 0.198577f
C13205 _174_ cal_count\[1\] 0.081252f
C13206 _096_ _116_ 0.020685f
C13207 output34/a_224_472# ctlp[1] 0.00277f
C13208 _073_ cal_itt\[0\] 0.211566f
C13209 _126_ _076_ 0.005517f
C13210 net63 FILLER_0_18_177/a_932_472# 0.063742f
C13211 net10 _411_/a_36_151# 0.127193f
C13212 _267_/a_36_472# _113_ 0.014178f
C13213 FILLER_0_15_142/a_124_375# _095_ 0.003935f
C13214 _285_/a_36_472# _094_ 0.045394f
C13215 _415_/a_36_151# FILLER_0_10_256/a_36_472# 0.004847f
C13216 net38 _445_/a_448_472# 0.023336f
C13217 net27 FILLER_0_15_235/a_572_375# 0.001554f
C13218 _270_/a_36_472# net21 0.001606f
C13219 net44 net17 0.046636f
C13220 net82 FILLER_0_3_172/a_2276_472# 0.007729f
C13221 net82 _386_/a_1084_68# 0.001068f
C13222 net20 _055_ 0.203142f
C13223 FILLER_0_15_116/a_484_472# _136_ 0.002712f
C13224 FILLER_0_9_282/a_36_472# vss 0.002224f
C13225 FILLER_0_4_107/a_1020_375# _158_ 0.003535f
C13226 FILLER_0_4_107/a_484_472# _369_/a_36_68# 0.001049f
C13227 FILLER_0_4_144/a_36_472# _152_ 0.008211f
C13228 FILLER_0_4_144/a_484_472# _081_ 0.001145f
C13229 _093_ _110_ 0.08348f
C13230 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1380_472# 0.003468f
C13231 _132_ vss 0.492496f
C13232 FILLER_0_5_54/a_1020_375# _440_/a_36_151# 0.059049f
C13233 FILLER_0_9_28/a_124_375# output42/a_224_472# 0.003337f
C13234 vss FILLER_0_22_107/a_484_472# 0.003617f
C13235 _094_ _418_/a_2248_156# 0.028557f
C13236 FILLER_0_8_138/a_124_375# vss 0.00629f
C13237 FILLER_0_8_138/a_36_472# vdd 0.008749f
C13238 _086_ _056_ 0.043494f
C13239 _028_ FILLER_0_7_72/a_1380_472# 0.001777f
C13240 output13/a_224_472# vss 0.108144f
C13241 FILLER_0_21_206/a_36_472# net33 0.001447f
C13242 FILLER_0_7_195/a_36_472# cal_itt\[3\] 0.070665f
C13243 _414_/a_36_151# _161_ 0.033054f
C13244 _053_ _365_/a_36_68# 0.001572f
C13245 _052_ FILLER_0_18_61/a_36_472# 0.001508f
C13246 _144_ _340_/a_36_160# 0.008886f
C13247 _132_ net74 0.031741f
C13248 _056_ cal_count\[3\] 0.186969f
C13249 _050_ mask\[7\] 0.128172f
C13250 FILLER_0_18_107/a_932_472# FILLER_0_17_104/a_1380_472# 0.026657f
C13251 net72 _394_/a_244_524# 0.001083f
C13252 _053_ FILLER_0_7_72/a_3260_375# 0.071059f
C13253 _050_ _148_ 0.002456f
C13254 _091_ _043_ 0.041409f
C13255 _256_/a_1612_497# _055_ 0.001438f
C13256 mask\[4\] FILLER_0_18_177/a_1916_375# 0.013466f
C13257 FILLER_0_20_15/a_932_472# vdd 0.002617f
C13258 net50 FILLER_0_4_91/a_484_472# 0.008749f
C13259 _149_ _098_ 0.398643f
C13260 _000_ FILLER_0_3_221/a_932_472# 0.008308f
C13261 FILLER_0_18_209/a_572_375# _201_/a_67_603# 0.008812f
C13262 _256_/a_716_497# calibrate 0.001066f
C13263 _140_ FILLER_0_22_128/a_3172_472# 0.005458f
C13264 _105_ result[6] 0.001477f
C13265 _432_/a_796_472# _093_ 0.002586f
C13266 _274_/a_36_68# vss 0.052669f
C13267 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001723f
C13268 net20 FILLER_0_6_231/a_124_375# 0.060499f
C13269 net57 _066_ 0.069098f
C13270 _013_ FILLER_0_17_56/a_484_472# 0.002659f
C13271 _131_ FILLER_0_14_107/a_1380_472# 0.01797f
C13272 _065_ _441_/a_448_472# 0.001973f
C13273 _065_ _235_/a_67_603# 0.004135f
C13274 _392_/a_36_68# cal_count\[3\] 0.003072f
C13275 net53 _043_ 0.053033f
C13276 net48 _251_/a_468_472# 0.002731f
C13277 _256_/a_36_68# net4 0.017783f
C13278 _077_ _076_ 1.895143f
C13279 output35/a_224_472# output19/a_224_472# 0.015892f
C13280 output33/a_224_472# net61 0.04987f
C13281 _422_/a_1204_472# _109_ 0.001807f
C13282 _178_ _402_/a_1296_93# 0.062418f
C13283 _070_ FILLER_0_10_107/a_36_472# 0.013252f
C13284 _428_/a_2248_156# vdd 0.006977f
C13285 net32 net34 0.330134f
C13286 net79 net77 0.431572f
C13287 _031_ FILLER_0_2_127/a_36_472# 0.016207f
C13288 _120_ FILLER_0_8_156/a_572_375# 0.030218f
C13289 _119_ _125_ 0.11554f
C13290 FILLER_0_5_54/a_572_375# vss 0.002617f
C13291 FILLER_0_5_54/a_1020_375# vdd -0.014642f
C13292 result[6] _010_ 0.056004f
C13293 _069_ mask\[1\] 0.029447f
C13294 FILLER_0_7_72/a_2276_472# FILLER_0_6_90/a_124_375# 0.001684f
C13295 _036_ net17 0.153479f
C13296 _238_/a_67_603# net52 0.006325f
C13297 FILLER_0_4_177/a_572_375# vss 0.054783f
C13298 FILLER_0_4_177/a_36_472# vdd 0.114788f
C13299 _412_/a_2248_156# fanout59/a_36_160# 0.007753f
C13300 net57 FILLER_0_8_156/a_484_472# 0.008895f
C13301 FILLER_0_15_72/a_484_472# vss 0.010761f
C13302 _415_/a_1308_423# net19 0.001498f
C13303 _445_/a_2665_112# net17 0.006445f
C13304 _428_/a_1204_472# net74 0.009712f
C13305 mask\[5\] output35/a_224_472# 0.003461f
C13306 _414_/a_2560_156# _053_ 0.008732f
C13307 net50 vss 1.178736f
C13308 output29/a_224_472# _044_ 0.087528f
C13309 net29 mask\[1\] 0.023266f
C13310 _421_/a_36_151# _010_ 0.015107f
C13311 output32/a_224_472# result[5] 0.047325f
C13312 _091_ net21 0.030022f
C13313 net20 FILLER_0_13_212/a_1468_375# 0.009573f
C13314 FILLER_0_4_99/a_36_472# _160_ 0.006222f
C13315 _028_ FILLER_0_7_59/a_572_375# 0.00133f
C13316 net57 net37 0.091923f
C13317 _141_ FILLER_0_19_155/a_484_472# 0.015625f
C13318 fanout55/a_36_160# _067_ 0.126784f
C13319 net55 FILLER_0_18_76/a_572_375# 0.002278f
C13320 _181_ cal_count\[0\] 0.001114f
C13321 _443_/a_1204_472# vss 0.005425f
C13322 _443_/a_2248_156# vdd 0.010579f
C13323 net1 fanout58/a_36_160# 0.060243f
C13324 _008_ net64 0.001427f
C13325 _021_ _097_ 0.002219f
C13326 output44/a_224_472# vss 0.014054f
C13327 _253_/a_36_68# cal_itt\[1\] 0.039692f
C13328 FILLER_0_7_72/a_36_472# net52 0.014911f
C13329 FILLER_0_7_72/a_2812_375# net50 0.006598f
C13330 FILLER_0_19_28/a_572_375# net40 0.00139f
C13331 output28/a_224_472# _416_/a_2665_112# 0.008243f
C13332 fanout79/a_36_160# net79 0.011193f
C13333 result[1] _416_/a_1308_423# 0.002597f
C13334 FILLER_0_14_50/a_124_375# _174_ 0.033245f
C13335 ctlp[6] vdd 0.207209f
C13336 _028_ net14 0.066292f
C13337 net70 FILLER_0_14_107/a_124_375# 0.029975f
C13338 net27 _426_/a_1000_472# 0.002971f
C13339 _431_/a_1000_472# net36 0.001771f
C13340 FILLER_0_18_2/a_2812_375# FILLER_0_19_28/a_36_472# 0.001684f
C13341 output12/a_224_472# net22 0.002662f
C13342 _328_/a_36_113# net14 0.002272f
C13343 _248_/a_36_68# _090_ 0.041161f
C13344 _147_ _049_ 0.001131f
C13345 net8 vdd 0.593788f
C13346 _059_ net47 0.00606f
C13347 _371_/a_36_113# _152_ 0.001083f
C13348 FILLER_0_16_57/a_1020_375# _131_ 0.012481f
C13349 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1380_472# 0.026657f
C13350 ctlp[2] _011_ 0.101324f
C13351 output41/a_224_472# trim[3] 0.042209f
C13352 output25/a_224_472# mask\[8\] 0.015742f
C13353 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_572_375# 0.086635f
C13354 net67 FILLER_0_6_47/a_36_472# 0.004607f
C13355 output46/a_224_472# FILLER_0_20_15/a_124_375# 0.029497f
C13356 FILLER_0_15_72/a_484_472# cal_count\[1\] 0.013337f
C13357 _083_ _080_ 0.043927f
C13358 net16 FILLER_0_18_37/a_484_472# 0.054878f
C13359 net15 FILLER_0_15_72/a_572_375# 0.002741f
C13360 _096_ _225_/a_36_160# 0.004807f
C13361 _053_ _042_ 0.00242f
C13362 FILLER_0_4_99/a_36_472# _030_ 0.002699f
C13363 _069_ vss 0.323941f
C13364 net52 net15 0.166073f
C13365 fanout72/a_36_113# _043_ 0.017862f
C13366 _093_ fanout54/a_36_160# 0.003506f
C13367 net52 fanout51/a_36_113# 0.036773f
C13368 cal_itt\[2\] _253_/a_36_68# 0.010756f
C13369 _091_ FILLER_0_18_177/a_124_375# 0.010316f
C13370 _308_/a_848_380# net14 0.021982f
C13371 _150_ vdd 0.05295f
C13372 _090_ _060_ 0.396493f
C13373 net34 FILLER_0_22_177/a_572_375# 0.006974f
C13374 FILLER_0_18_2/a_3172_472# net55 0.00602f
C13375 _189_/a_67_603# _429_/a_2665_112# 0.015187f
C13376 net29 vss 0.259409f
C13377 net36 FILLER_0_15_180/a_124_375# 0.004275f
C13378 ctlp[1] _419_/a_1000_472# 0.005263f
C13379 FILLER_0_10_78/a_484_472# FILLER_0_9_72/a_1020_375# 0.001543f
C13380 _016_ _127_ 0.01898f
C13381 _248_/a_36_68# net22 0.002193f
C13382 _412_/a_1000_472# vdd 0.002008f
C13383 _121_ FILLER_0_8_156/a_124_375# 0.033427f
C13384 ctln[4] _411_/a_36_151# 0.0022f
C13385 _170_ vdd 0.18848f
C13386 FILLER_0_3_172/a_124_375# net22 0.01308f
C13387 output25/a_224_472# vss 0.080847f
C13388 _105_ mask\[4\] 0.025209f
C13389 _106_ _291_/a_36_160# 0.054237f
C13390 FILLER_0_15_142/a_124_375# vss 0.009207f
C13391 FILLER_0_15_142/a_572_375# vdd -0.013698f
C13392 trim_mask\[3\] vss 0.156544f
C13393 _074_ _014_ 0.001557f
C13394 net20 _106_ 0.050151f
C13395 FILLER_0_18_37/a_1468_375# vss 0.054381f
C13396 FILLER_0_18_37/a_36_472# vdd 0.136723f
C13397 net45 net17 0.192181f
C13398 _008_ vss 0.355468f
C13399 _141_ FILLER_0_22_128/a_3260_375# 0.003544f
C13400 output7/a_224_472# output40/a_224_472# 0.038066f
C13401 net39 net44 0.0112f
C13402 _322_/a_848_380# _070_ 0.006182f
C13403 _216_/a_67_603# net15 0.060076f
C13404 mask\[0\] _136_ 0.025838f
C13405 _060_ net22 0.533421f
C13406 _091_ FILLER_0_19_171/a_1380_472# 0.001044f
C13407 net76 FILLER_0_2_177/a_124_375# 0.00439f
C13408 FILLER_0_15_10/a_124_375# FILLER_0_15_2/a_572_375# 0.012001f
C13409 FILLER_0_15_116/a_124_375# vdd 0.012886f
C13410 FILLER_0_6_90/a_36_472# net14 0.002705f
C13411 FILLER_0_15_142/a_124_375# net74 0.005931f
C13412 _428_/a_36_151# net14 0.004485f
C13413 _119_ FILLER_0_8_138/a_124_375# 0.006523f
C13414 mask\[9\] FILLER_0_20_98/a_36_472# 0.005917f
C13415 net81 _060_ 0.019654f
C13416 FILLER_0_14_107/a_36_472# _043_ 0.001661f
C13417 _448_/a_2248_156# _037_ 0.027079f
C13418 _050_ FILLER_0_22_128/a_932_472# 0.001098f
C13419 FILLER_0_4_144/a_572_375# trim_mask\[4\] 0.014071f
C13420 net79 _283_/a_36_472# 0.010249f
C13421 output19/a_224_472# mask\[7\] 0.001181f
C13422 _442_/a_36_151# net13 0.009343f
C13423 _053_ _086_ 0.091538f
C13424 _114_ _128_ 0.047516f
C13425 _118_ _113_ 0.005092f
C13426 FILLER_0_4_197/a_1380_472# net82 0.003084f
C13427 _081_ _001_ 0.012101f
C13428 _429_/a_2665_112# FILLER_0_14_235/a_124_375# 0.006271f
C13429 _436_/a_1308_423# _025_ 0.006243f
C13430 FILLER_0_17_38/a_124_375# _452_/a_36_151# 0.006111f
C13431 FILLER_0_4_152/a_36_472# _170_ 0.005476f
C13432 result[7] _419_/a_2248_156# 0.001916f
C13433 _095_ FILLER_0_13_142/a_36_472# 0.001782f
C13434 net22 net12 0.032084f
C13435 _075_ vss 0.046342f
C13436 net52 net51 0.091698f
C13437 FILLER_0_17_226/a_36_472# _093_ 0.004282f
C13438 _074_ _070_ 0.102481f
C13439 _139_ _098_ 0.026578f
C13440 _093_ FILLER_0_18_139/a_124_375# 0.008393f
C13441 _235_/a_67_603# _036_ 0.043345f
C13442 net55 _120_ 0.001054f
C13443 trim_val\[1\] net47 0.34878f
C13444 FILLER_0_12_136/a_124_375# _127_ 0.004013f
C13445 FILLER_0_18_209/a_484_472# vss 0.005794f
C13446 net49 _440_/a_2665_112# 0.025303f
C13447 _064_ _445_/a_36_151# 0.03209f
C13448 _447_/a_36_151# net68 0.040925f
C13449 trim_mask\[2\] trim_mask\[1\] 0.002186f
C13450 _414_/a_1456_156# cal_itt\[3\] 0.001134f
C13451 net64 FILLER_0_15_235/a_36_472# 0.046292f
C13452 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_124_375# 0.026339f
C13453 output48/a_224_472# _081_ 0.007705f
C13454 output32/a_224_472# net19 0.08441f
C13455 FILLER_0_20_177/a_124_375# vss 0.002674f
C13456 FILLER_0_20_177/a_572_375# vdd -0.001627f
C13457 _088_ FILLER_0_3_221/a_124_375# 0.002378f
C13458 _322_/a_848_380# FILLER_0_9_142/a_36_472# 0.011591f
C13459 mask\[5\] mask\[7\] 0.014384f
C13460 result[5] _418_/a_36_151# 0.009705f
C13461 _067_ net6 0.015232f
C13462 net32 _419_/a_2665_112# 0.027035f
C13463 net57 en_co_clk 0.195533f
C13464 _091_ FILLER_0_15_212/a_1020_375# 0.00799f
C13465 _431_/a_1000_472# _020_ 0.009685f
C13466 FILLER_0_15_235/a_36_472# mask\[1\] 0.009316f
C13467 _053_ _154_ 0.41707f
C13468 FILLER_0_7_104/a_932_472# _062_ 0.001184f
C13469 trim[4] FILLER_0_8_2/a_124_375# 0.028454f
C13470 net16 _453_/a_36_151# 0.001634f
C13471 _028_ FILLER_0_6_90/a_572_375# 0.015802f
C13472 net38 FILLER_0_8_24/a_124_375# 0.001013f
C13473 FILLER_0_16_255/a_36_472# net30 0.00209f
C13474 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_36_472# 0.086635f
C13475 _079_ net22 0.039221f
C13476 net41 net51 0.031531f
C13477 FILLER_0_17_104/a_36_472# vss 0.002744f
C13478 FILLER_0_17_104/a_484_472# vdd 0.020339f
C13479 _318_/a_224_472# _124_ 0.001288f
C13480 _012_ vdd 0.261844f
C13481 result[9] _419_/a_1308_423# 0.012036f
C13482 ctln[0] vss 0.125714f
C13483 _050_ FILLER_0_22_107/a_124_375# 0.002634f
C13484 net63 _139_ 0.003073f
C13485 mask\[2\] FILLER_0_15_212/a_36_472# 0.001181f
C13486 _161_ net21 0.011799f
C13487 net26 FILLER_0_21_28/a_1468_375# 0.041169f
C13488 _419_/a_36_151# vdd -0.110366f
C13489 _136_ _451_/a_36_151# 0.043941f
C13490 net63 result[8] 0.013631f
C13491 _430_/a_2248_156# mask\[1\] 0.001498f
C13492 _413_/a_1000_472# _002_ 0.006249f
C13493 net39 _445_/a_2665_112# 0.002831f
C13494 _086_ FILLER_0_4_177/a_124_375# 0.024433f
C13495 _317_/a_36_113# FILLER_0_7_233/a_124_375# 0.03227f
C13496 net52 FILLER_0_9_72/a_1020_375# 0.00799f
C13497 _267_/a_36_472# vdd 0.005477f
C13498 _053_ _169_ 0.014161f
C13499 FILLER_0_15_59/a_572_375# vdd 0.03104f
C13500 FILLER_0_21_286/a_36_472# net77 0.001557f
C13501 FILLER_0_15_59/a_124_375# vss 0.003806f
C13502 _120_ net23 0.147166f
C13503 net20 _274_/a_1164_497# 0.002879f
C13504 net57 _395_/a_1044_488# 0.002526f
C13505 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_484_472# 0.013276f
C13506 fanout60/a_36_160# _417_/a_36_151# 0.062739f
C13507 net75 _316_/a_692_472# 0.00138f
C13508 net44 _452_/a_2449_156# 0.0059f
C13509 FILLER_0_19_171/a_1468_375# vdd 0.064097f
C13510 _027_ net71 0.057875f
C13511 _131_ FILLER_0_17_64/a_124_375# 0.005913f
C13512 _348_/a_257_69# mask\[6\] 0.00159f
C13513 state\[2\] FILLER_0_13_142/a_1380_472# 0.019965f
C13514 net15 FILLER_0_18_61/a_124_375# 0.001179f
C13515 FILLER_0_15_235/a_484_472# vdd 0.006f
C13516 FILLER_0_15_235/a_36_472# vss 0.003138f
C13517 _178_ FILLER_0_16_37/a_124_375# 0.036901f
C13518 _346_/a_49_472# _098_ 0.028579f
C13519 FILLER_0_17_282/a_36_472# _418_/a_448_472# 0.011962f
C13520 FILLER_0_18_177/a_3260_375# net21 0.005704f
C13521 calibrate _123_ 0.016296f
C13522 _438_/a_448_472# vdd 0.009409f
C13523 _438_/a_36_151# vss 0.014203f
C13524 FILLER_0_17_161/a_124_375# _098_ 0.002013f
C13525 _128_ _126_ 0.008298f
C13526 FILLER_0_10_28/a_36_472# net51 0.00703f
C13527 result[2] FILLER_0_13_290/a_36_472# 0.016496f
C13528 _105_ net34 0.784678f
C13529 mask\[3\] fanout63/a_36_160# 0.002585f
C13530 vss result[3] 0.28152f
C13531 _415_/a_2248_156# fanout62/a_36_160# 0.007753f
C13532 cal_count\[1\] FILLER_0_15_59/a_124_375# 0.010034f
C13533 FILLER_0_9_28/a_1916_375# net68 0.050307f
C13534 _119_ _069_ 0.00226f
C13535 net73 FILLER_0_18_107/a_484_472# 0.0052f
C13536 FILLER_0_0_130/a_36_472# vss 0.00351f
C13537 net4 _223_/a_36_160# 0.020711f
C13538 mask\[7\] _299_/a_36_472# 0.033949f
C13539 FILLER_0_19_125/a_124_375# vdd 0.032954f
C13540 FILLER_0_16_89/a_1468_375# net14 0.022582f
C13541 FILLER_0_24_96/a_124_375# vss 0.017357f
C13542 FILLER_0_24_96/a_36_472# vdd 0.094828f
C13543 FILLER_0_16_107/a_484_472# _136_ 0.013449f
C13544 _430_/a_2248_156# vss 0.030251f
C13545 _432_/a_1308_423# net80 0.030835f
C13546 _430_/a_2665_112# vdd 0.021353f
C13547 _068_ _118_ 1.374452f
C13548 _070_ _124_ 0.114614f
C13549 _069_ FILLER_0_11_142/a_484_472# 0.005789f
C13550 FILLER_0_4_99/a_36_472# _156_ 0.0255f
C13551 FILLER_0_18_107/a_932_472# mask\[9\] 0.005296f
C13552 output27/a_224_472# net64 0.04953f
C13553 result[9] _420_/a_2560_156# 0.002295f
C13554 net19 FILLER_0_14_263/a_36_472# 0.135429f
C13555 FILLER_0_6_47/a_124_375# vdd 0.008011f
C13556 net52 _163_ 0.00157f
C13557 trimb[1] net38 0.161478f
C13558 net57 _122_ 0.034045f
C13559 _420_/a_2248_156# vdd 0.00331f
C13560 _079_ _076_ 0.001575f
C13561 net75 net76 0.106326f
C13562 net20 FILLER_0_1_212/a_36_472# 0.013846f
C13563 net23 FILLER_0_16_154/a_124_375# 0.002689f
C13564 net53 _451_/a_448_472# 0.026909f
C13565 net70 _451_/a_836_156# 0.006451f
C13566 net73 _136_ 0.050578f
C13567 _002_ _089_ 0.002349f
C13568 _370_/a_848_380# net23 0.001196f
C13569 _013_ FILLER_0_18_37/a_932_472# 0.010651f
C13570 mask\[3\] FILLER_0_17_218/a_484_472# 0.017442f
C13571 _057_ _267_/a_36_472# 0.038568f
C13572 _376_/a_36_160# FILLER_0_6_79/a_36_472# 0.003913f
C13573 _077_ _128_ 0.005311f
C13574 _449_/a_2665_112# _038_ 0.024406f
C13575 FILLER_0_13_142/a_36_472# vss 0.005768f
C13576 trim[0] FILLER_0_3_2/a_124_375# 0.020708f
C13577 net16 _165_ 0.021744f
C13578 _431_/a_2665_112# FILLER_0_16_154/a_124_375# 0.006271f
C13579 _004_ _005_ 0.004158f
C13580 _392_/a_244_472# _067_ 0.001893f
C13581 net38 _043_ 0.117134f
C13582 ctlp[3] net61 0.007397f
C13583 _227_/a_36_160# net23 0.055152f
C13584 net25 net24 0.031854f
C13585 _008_ _103_ 0.092504f
C13586 FILLER_0_16_57/a_572_375# FILLER_0_15_59/a_484_472# 0.001543f
C13587 FILLER_0_8_107/a_36_472# _133_ 0.00589f
C13588 FILLER_0_7_59/a_36_472# net68 0.050931f
C13589 net57 _061_ 0.127011f
C13590 _415_/a_36_151# output28/a_224_472# 0.229574f
C13591 _177_ _451_/a_3129_107# 0.043731f
C13592 mask\[1\] net22 0.029526f
C13593 _421_/a_2665_112# vss 0.002792f
C13594 _421_/a_2560_156# vdd 0.001862f
C13595 net74 FILLER_0_13_142/a_36_472# 0.003568f
C13596 _392_/a_36_68# _120_ 0.001738f
C13597 net81 net64 0.455159f
C13598 ctln[5] _448_/a_1308_423# 0.004061f
C13599 _442_/a_2665_112# net14 0.011563f
C13600 output27/a_224_472# vss 0.027374f
C13601 _422_/a_796_472# vdd 0.003546f
C13602 net81 mask\[1\] 2.509493f
C13603 trim_mask\[4\] FILLER_0_2_111/a_1020_375# 0.02806f
C13604 _098_ FILLER_0_15_205/a_124_375# 0.009558f
C13605 _426_/a_2248_156# vdd 0.003943f
C13606 net36 _099_ 0.325141f
C13607 FILLER_0_10_78/a_124_375# _176_ 0.002785f
C13608 FILLER_0_15_282/a_36_472# vss 0.004616f
C13609 _446_/a_2560_156# net40 0.012204f
C13610 _081_ _316_/a_124_24# 0.011421f
C13611 FILLER_0_11_101/a_484_472# vss 0.003923f
C13612 trim_val\[2\] _446_/a_2665_112# 0.012621f
C13613 _090_ vss 0.267577f
C13614 _113_ vdd 0.774039f
C13615 FILLER_0_6_177/a_124_375# net47 0.002925f
C13616 _112_ _316_/a_848_380# 0.022235f
C13617 _305_/a_36_159# calibrate 0.003505f
C13618 fanout61/a_36_113# vss 0.05514f
C13619 _445_/a_2248_156# _444_/a_36_151# 0.001081f
C13620 FILLER_0_3_221/a_572_375# vss 0.003292f
C13621 fanout54/a_36_160# FILLER_0_18_139/a_1020_375# 0.031033f
C13622 FILLER_0_4_49/a_36_472# _164_ 0.033727f
C13623 _438_/a_796_472# net71 0.00514f
C13624 net65 FILLER_0_3_172/a_2276_472# 0.001777f
C13625 ctlp[3] _108_ 0.009437f
C13626 net63 _435_/a_2560_156# 0.023868f
C13627 output8/a_224_472# _411_/a_1308_423# 0.005111f
C13628 FILLER_0_5_72/a_124_375# _029_ 0.010208f
C13629 _408_/a_718_524# net40 0.011463f
C13630 _394_/a_728_93# FILLER_0_15_72/a_572_375# 0.02852f
C13631 _239_/a_36_160# _065_ 0.032139f
C13632 _413_/a_448_472# net59 0.059041f
C13633 output34/a_224_472# _199_/a_36_160# 0.003531f
C13634 FILLER_0_23_60/a_124_375# FILLER_0_23_44/a_1468_375# 0.012001f
C13635 net22 vss 1.28233f
C13636 FILLER_0_15_150/a_36_472# net23 0.010444f
C13637 _054_ net40 0.072879f
C13638 net63 FILLER_0_15_205/a_124_375# 0.001597f
C13639 fanout49/a_36_160# FILLER_0_4_91/a_36_472# 0.001461f
C13640 _074_ net9 0.002862f
C13641 _255_/a_224_552# _074_ 0.005907f
C13642 cal_count\[2\] net40 0.313209f
C13643 _379_/a_36_472# _164_ 0.026812f
C13644 _093_ _150_ 0.406318f
C13645 FILLER_0_2_111/a_124_375# vdd 0.024756f
C13646 net63 _098_ 0.055686f
C13647 net81 vss 0.766885f
C13648 net66 _167_ 0.016569f
C13649 ctln[6] net23 0.003826f
C13650 FILLER_0_3_78/a_484_472# _164_ 0.05311f
C13651 FILLER_0_4_99/a_124_375# net47 0.001409f
C13652 FILLER_0_12_28/a_36_472# _450_/a_3129_107# 0.009814f
C13653 _081_ FILLER_0_5_148/a_36_472# 0.020403f
C13654 _118_ vdd 0.292155f
C13655 _043_ FILLER_0_13_72/a_484_472# 0.016114f
C13656 mask\[9\] _437_/a_2665_112# 0.014146f
C13657 net26 _424_/a_1308_423# 0.001179f
C13658 _431_/a_2665_112# FILLER_0_15_150/a_36_472# 0.035266f
C13659 ctln[8] vdd 0.125219f
C13660 FILLER_0_4_107/a_36_472# trim_mask\[3\] 0.00152f
C13661 _086_ _072_ 0.220767f
C13662 fanout78/a_36_113# _418_/a_36_151# 0.030244f
C13663 FILLER_0_18_107/a_1828_472# vdd 0.004446f
C13664 trim_val\[1\] FILLER_0_6_47/a_36_472# 0.00351f
C13665 fanout60/a_36_160# _418_/a_36_151# 0.029017f
C13666 net78 _419_/a_36_151# 0.007437f
C13667 net60 _419_/a_36_151# 0.016173f
C13668 net61 _419_/a_1308_423# 0.00793f
C13669 input3/a_36_113# cal_count\[2\] 0.00555f
C13670 FILLER_0_14_107/a_484_472# _451_/a_36_151# 0.001723f
C13671 _005_ _044_ 0.50767f
C13672 net54 FILLER_0_22_128/a_1380_472# 0.008765f
C13673 _021_ net80 0.254353f
C13674 _341_/a_49_472# _137_ 0.059288f
C13675 FILLER_0_18_139/a_1380_472# _145_ 0.002077f
C13676 _417_/a_1000_472# _006_ 0.026299f
C13677 FILLER_0_16_89/a_484_472# _040_ 0.009871f
C13678 _058_ FILLER_0_9_105/a_36_472# 0.011426f
C13679 output47/a_224_472# _452_/a_2225_156# 0.012077f
C13680 _087_ vdd 0.281159f
C13681 _072_ cal_count\[3\] 0.028346f
C13682 _292_/a_36_160# mask\[5\] 0.007486f
C13683 FILLER_0_16_107/a_124_375# vdd 0.026251f
C13684 net75 _083_ 0.055491f
C13685 trimb[1] net55 0.017528f
C13686 _035_ vss 0.105648f
C13687 net16 _095_ 0.042842f
C13688 ctlp[4] result[8] 0.151286f
C13689 fanout81/a_36_160# net76 0.001905f
C13690 fanout49/a_36_160# vdd 0.099887f
C13691 FILLER_0_5_164/a_484_472# _163_ 0.029894f
C13692 net47 output6/a_224_472# 0.070584f
C13693 FILLER_0_18_171/a_36_472# _098_ 0.020038f
C13694 fanout71/a_36_113# mask\[9\] 0.044939f
C13695 net20 FILLER_0_15_235/a_124_375# 0.001278f
C13696 net45 ctlp[0] 0.001134f
C13697 _414_/a_36_151# _056_ 0.00356f
C13698 FILLER_0_10_78/a_932_472# _120_ 0.003672f
C13699 _038_ vss 0.373776f
C13700 _315_/a_36_68# _121_ 0.031617f
C13701 _057_ _113_ 0.339862f
C13702 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_36_472# 0.026657f
C13703 net55 FILLER_0_17_38/a_572_375# 0.007646f
C13704 result[1] net18 0.056799f
C13705 _161_ _062_ 0.046903f
C13706 FILLER_0_16_255/a_36_472# _417_/a_2665_112# 0.003221f
C13707 net20 net30 0.033149f
C13708 net4 FILLER_0_12_220/a_572_375# 0.019052f
C13709 _004_ FILLER_0_10_256/a_124_375# 0.006989f
C13710 fanout70/a_36_113# vdd 0.015969f
C13711 FILLER_0_17_104/a_572_375# _040_ 0.001228f
C13712 FILLER_0_7_104/a_124_375# _058_ 0.006125f
C13713 FILLER_0_22_177/a_932_472# mask\[6\] 0.006573f
C13714 _450_/a_2225_156# _039_ 0.034731f
C13715 net55 _043_ 0.053191f
C13716 net74 _038_ 0.055774f
C13717 mask\[4\] _145_ 0.340415f
C13718 _431_/a_36_151# net53 0.001579f
C13719 _431_/a_796_472# net70 0.001754f
C13720 output21/a_224_472# output19/a_224_472# 0.007877f
C13721 net54 FILLER_0_22_107/a_572_375# 0.002239f
C13722 _068_ vdd 0.793549f
C13723 _076_ vss 1.132839f
C13724 _443_/a_1456_156# net23 0.001009f
C13725 FILLER_0_5_54/a_572_375# _029_ 0.00494f
C13726 FILLER_0_18_100/a_124_375# _438_/a_2665_112# 0.010688f
C13727 _449_/a_2248_156# vdd -0.001225f
C13728 _449_/a_1204_472# vss 0.006048f
C13729 FILLER_0_16_255/a_36_472# _045_ 0.001653f
C13730 fanout50/a_36_160# net49 0.030626f
C13731 _440_/a_2665_112# net47 0.014066f
C13732 net34 _024_ 0.009705f
C13733 net35 FILLER_0_22_86/a_1468_375# 0.010438f
C13734 mask\[8\] FILLER_0_22_86/a_36_472# 0.012471f
C13735 net52 _442_/a_796_472# 0.004871f
C13736 _114_ _311_/a_2700_473# 0.005178f
C13737 FILLER_0_17_72/a_3260_375# vss 0.052993f
C13738 FILLER_0_17_72/a_36_472# vdd 0.111688f
C13739 _075_ FILLER_0_5_206/a_36_472# 0.001503f
C13740 FILLER_0_16_89/a_36_472# net36 0.010907f
C13741 net60 _420_/a_2248_156# 0.035104f
C13742 net78 _420_/a_2248_156# 0.001534f
C13743 _093_ FILLER_0_17_104/a_484_472# 0.014431f
C13744 net50 _029_ 0.025102f
C13745 _093_ _012_ 0.141641f
C13746 _429_/a_448_472# _043_ 0.003615f
C13747 trimb[1] FILLER_0_18_2/a_484_472# 0.009245f
C13748 _095_ FILLER_0_14_107/a_1380_472# 0.011439f
C13749 output21/a_224_472# mask\[5\] 0.009585f
C13750 net55 _175_ 0.142124f
C13751 _057_ _118_ 0.055726f
C13752 _128_ _426_/a_2665_112# 0.025626f
C13753 net44 FILLER_0_15_2/a_484_472# 0.047161f
C13754 FILLER_0_22_86/a_36_472# vss 0.002319f
C13755 _189_/a_67_603# _043_ 0.005635f
C13756 _131_ FILLER_0_17_56/a_36_472# 0.001491f
C13757 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_484_472# 0.001723f
C13758 _128_ _060_ 0.022833f
C13759 FILLER_0_7_59/a_484_472# net67 0.03109f
C13760 FILLER_0_19_111/a_124_375# vdd 0.005128f
C13761 net31 net29 0.009564f
C13762 mask\[8\] _437_/a_2560_156# 0.001171f
C13763 _422_/a_2560_156# _009_ 0.002551f
C13764 _341_/a_49_472# net56 0.018486f
C13765 net23 _043_ 0.042095f
C13766 _065_ _030_ 0.001499f
C13767 net41 net66 0.08664f
C13768 _449_/a_796_472# net15 0.006722f
C13769 net69 FILLER_0_3_78/a_124_375# 0.004201f
C13770 _230_/a_652_68# _062_ 0.001144f
C13771 FILLER_0_19_125/a_124_375# _433_/a_36_151# 0.001597f
C13772 _178_ _182_ 0.067534f
C13773 net69 FILLER_0_2_101/a_124_375# 0.015032f
C13774 net31 _008_ 0.292444f
C13775 _089_ net76 0.017609f
C13776 FILLER_0_19_55/a_124_375# _216_/a_67_603# 0.003017f
C13777 _411_/a_2665_112# net8 0.036782f
C13778 _093_ _438_/a_448_472# 0.0106f
C13779 FILLER_0_4_123/a_124_375# _152_ 0.039668f
C13780 FILLER_0_11_101/a_36_472# cal_count\[3\] 0.005101f
C13781 net20 _421_/a_1204_472# 0.019627f
C13782 net60 _421_/a_2560_156# 0.001951f
C13783 _176_ net36 0.336675f
C13784 net53 _427_/a_448_472# 0.047356f
C13785 _444_/a_1308_423# net67 0.021684f
C13786 _373_/a_1458_68# _113_ 0.001257f
C13787 net57 _428_/a_2248_156# 0.022587f
C13788 net20 _422_/a_36_151# 0.083307f
C13789 trim_mask\[1\] FILLER_0_5_88/a_36_472# 0.038642f
C13790 _139_ _137_ 0.093639f
C13791 _429_/a_448_472# net21 0.014792f
C13792 FILLER_0_7_195/a_36_472# _161_ 0.015074f
C13793 net3 _190_/a_36_160# 0.013324f
C13794 FILLER_0_17_282/a_36_472# _006_ 0.002964f
C13795 _440_/a_36_151# vdd 0.117768f
C13796 _127_ _062_ 0.020537f
C13797 state\[0\] _426_/a_2665_112# 0.017088f
C13798 net16 ctln[9] 0.07797f
C13799 net38 _033_ 0.03598f
C13800 FILLER_0_4_197/a_36_472# net21 0.011079f
C13801 FILLER_0_6_239/a_124_375# net37 0.001989f
C13802 net75 FILLER_0_8_263/a_124_375# 0.001386f
C13803 _115_ _058_ 0.038308f
C13804 output19/a_224_472# ctlp[2] 0.04607f
C13805 net34 _435_/a_1308_423# 0.008652f
C13806 state\[0\] _060_ 0.047136f
C13807 _074_ _084_ 0.110937f
C13808 vss FILLER_0_4_91/a_572_375# 0.055113f
C13809 result[1] net62 0.061866f
C13810 net41 _067_ 0.033696f
C13811 _261_/a_36_160# net23 0.005015f
C13812 _115_ _315_/a_36_68# 0.001683f
C13813 _057_ _068_ 0.393271f
C13814 _402_/a_728_93# _401_/a_36_68# 0.002178f
C13815 _087_ FILLER_0_5_172/a_36_472# 0.00443f
C13816 FILLER_0_21_206/a_124_375# net22 0.05301f
C13817 net57 _443_/a_2248_156# 0.001117f
C13818 FILLER_0_11_78/a_484_472# vss 0.004063f
C13819 output20/a_224_472# vss -0.004787f
C13820 net27 net37 0.003648f
C13821 _024_ FILLER_0_22_177/a_124_375# 0.005166f
C13822 _141_ FILLER_0_16_154/a_36_472# 0.00126f
C13823 _432_/a_2560_156# _091_ 0.001542f
C13824 net65 net82 0.630327f
C13825 _444_/a_796_472# _054_ 0.001838f
C13826 output14/a_224_472# ctln[7] 0.076006f
C13827 net16 vss 0.679042f
C13828 _416_/a_2560_156# net62 0.010748f
C13829 _144_ _207_/a_67_603# 0.064623f
C13830 mask\[5\] ctlp[2] 0.104304f
C13831 _429_/a_2665_112# net62 0.02887f
C13832 FILLER_0_12_2/a_124_375# vdd 0.0247f
C13833 _423_/a_796_472# _012_ 0.015809f
C13834 _013_ _052_ 0.284735f
C13835 _422_/a_1204_472# _108_ 0.015401f
C13836 _430_/a_1308_423# net36 0.003317f
C13837 _412_/a_448_472# net1 0.035155f
C13838 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_572_375# 0.086635f
C13839 ctlp[1] net77 0.716304f
C13840 net69 _158_ 0.033459f
C13841 mask\[9\] net71 0.344312f
C13842 _116_ _176_ 0.067051f
C13843 _429_/a_36_151# _138_ 0.002064f
C13844 FILLER_0_13_100/a_36_472# net14 0.046864f
C13845 FILLER_0_3_172/a_3172_472# net22 0.010714f
C13846 FILLER_0_13_65/a_124_375# vdd 0.011301f
C13847 _306_/a_36_68# _116_ 0.00183f
C13848 net79 FILLER_0_12_220/a_572_375# 0.010889f
C13849 _152_ _163_ 0.05157f
C13850 FILLER_0_4_144/a_484_472# net23 0.01239f
C13851 net20 _413_/a_2665_112# 0.015855f
C13852 FILLER_0_17_72/a_932_472# net71 0.001418f
C13853 net49 _034_ 0.031359f
C13854 _053_ _414_/a_36_151# 0.035994f
C13855 FILLER_0_23_282/a_484_472# vss 0.005378f
C13856 _424_/a_2665_112# _012_ 0.01024f
C13857 net59 net11 0.016998f
C13858 FILLER_0_4_123/a_124_375# _070_ 0.001677f
C13859 _036_ _160_ 0.034434f
C13860 net57 _170_ 0.057355f
C13861 FILLER_0_7_72/a_1916_375# vss 0.001259f
C13862 FILLER_0_7_72/a_2364_375# vdd 0.018287f
C13863 net16 cal_count\[1\] 0.007291f
C13864 ctln[1] net10 0.029592f
C13865 _432_/a_1000_472# _137_ 0.008914f
C13866 FILLER_0_17_161/a_124_375# _137_ 0.016092f
C13867 FILLER_0_18_76/a_124_375# _438_/a_36_151# 0.001252f
C13868 _445_/a_1204_472# _034_ 0.003057f
C13869 _062_ FILLER_0_8_156/a_572_375# 0.002944f
C13870 net35 FILLER_0_22_177/a_932_472# 0.00643f
C13871 FILLER_0_22_86/a_1380_472# net71 0.011277f
C13872 _238_/a_67_603# FILLER_0_2_93/a_36_472# 0.002778f
C13873 net20 _014_ 0.008597f
C13874 output26/a_224_472# FILLER_0_23_60/a_36_472# 0.003292f
C13875 result[6] FILLER_0_21_286/a_572_375# 0.015047f
C13876 FILLER_0_8_263/a_124_375# FILLER_0_8_247/a_1468_375# 0.012001f
C13877 cal_count\[3\] _186_ 0.012453f
C13878 _086_ _133_ 0.035637f
C13879 _119_ _076_ 0.083673f
C13880 _052_ FILLER_0_21_28/a_2812_375# 0.002388f
C13881 FILLER_0_12_2/a_484_472# _450_/a_36_151# 0.059367f
C13882 FILLER_0_10_78/a_484_472# _115_ 0.005678f
C13883 _144_ FILLER_0_19_155/a_484_472# 0.006137f
C13884 net58 _073_ 0.057725f
C13885 _067_ _172_ 0.010195f
C13886 _448_/a_2665_112# vss 0.009029f
C13887 net33 net21 0.052426f
C13888 FILLER_0_13_212/a_36_472# _043_ 0.011752f
C13889 FILLER_0_2_93/a_484_472# FILLER_0_0_96/a_124_375# 0.001338f
C13890 _076_ _269_/a_36_472# 0.001618f
C13891 _131_ _372_/a_170_472# 0.002967f
C13892 net79 _417_/a_448_472# 0.028398f
C13893 FILLER_0_8_138/a_36_472# _129_ 0.055537f
C13894 _079_ FILLER_0_3_172/a_2276_472# 0.00261f
C13895 FILLER_0_8_263/a_124_375# _426_/a_36_151# 0.001252f
C13896 FILLER_0_14_107/a_1380_472# vss 0.001338f
C13897 FILLER_0_22_177/a_1380_472# vss 0.001502f
C13898 _444_/a_448_472# net47 0.030563f
C13899 FILLER_0_4_152/a_124_375# vss 0.019426f
C13900 FILLER_0_4_152/a_36_472# vdd 0.087397f
C13901 _053_ _372_/a_3126_472# 0.001056f
C13902 FILLER_0_22_177/a_1020_375# _435_/a_36_151# 0.059049f
C13903 _094_ net18 0.468109f
C13904 _013_ mask\[9\] 0.011224f
C13905 result[4] net30 0.298966f
C13906 _233_/a_36_160# _033_ 0.017573f
C13907 _063_ _165_ 0.021839f
C13908 _056_ net21 0.484506f
C13909 FILLER_0_16_255/a_36_472# _287_/a_36_472# 0.004546f
C13910 _036_ _030_ 0.430683f
C13911 output27/a_224_472# FILLER_0_9_290/a_36_472# 0.001711f
C13912 _447_/a_2665_112# net69 0.002067f
C13913 _114_ _131_ 0.036548f
C13914 net82 net69 0.005307f
C13915 _445_/a_2248_156# net49 0.029744f
C13916 _133_ _154_ 0.0133f
C13917 mask\[4\] _202_/a_36_160# 0.007912f
C13918 net19 _316_/a_848_380# 0.00558f
C13919 ctlp[2] _299_/a_36_472# 0.012937f
C13920 _267_/a_1792_472# _055_ 0.003058f
C13921 mask\[8\] _140_ 0.003375f
C13922 net20 _070_ 0.075448f
C13923 _108_ mask\[6\] 0.032481f
C13924 _452_/a_1040_527# vdd 0.004153f
C13925 result[8] _422_/a_1000_472# 0.001104f
C13926 ctln[2] net18 0.106494f
C13927 FILLER_0_22_86/a_932_472# _149_ 0.001205f
C13928 FILLER_0_22_86/a_36_472# _026_ 0.001503f
C13929 net20 FILLER_0_12_220/a_1380_472# 0.029747f
C13930 net52 FILLER_0_5_72/a_932_472# 0.008749f
C13931 net48 FILLER_0_7_233/a_124_375# 0.013455f
C13932 mask\[0\] _429_/a_1308_423# 0.019225f
C13933 net55 FILLER_0_18_53/a_124_375# 0.011674f
C13934 net72 FILLER_0_18_53/a_484_472# 0.001067f
C13935 FILLER_0_16_73/a_484_472# net55 0.004188f
C13936 _321_/a_170_472# _118_ 0.034852f
C13937 FILLER_0_18_177/a_1380_472# vdd 0.005692f
C13938 FILLER_0_18_177/a_932_472# vss -0.001894f
C13939 _328_/a_36_113# net70 0.00292f
C13940 fanout80/a_36_113# net21 0.021603f
C13941 output47/a_224_472# FILLER_0_15_2/a_36_472# 0.035046f
C13942 _070_ _163_ 1.884485f
C13943 _140_ vss 0.53195f
C13944 FILLER_0_20_177/a_1020_375# _098_ 0.013949f
C13945 _428_/a_2665_112# _131_ 0.006081f
C13946 _128_ net64 0.291788f
C13947 _093_ FILLER_0_18_107/a_1828_472# 0.001872f
C13948 _413_/a_36_151# FILLER_0_2_177/a_484_472# 0.006095f
C13949 _057_ vdd 0.801978f
C13950 _432_/a_448_472# net80 0.045963f
C13951 _402_/a_56_567# net40 0.033835f
C13952 FILLER_0_5_212/a_124_375# net59 0.045135f
C13953 _144_ FILLER_0_22_128/a_3260_375# 0.006444f
C13954 FILLER_0_5_128/a_572_375# vss 0.057605f
C13955 state\[2\] cal_count\[3\] 0.005312f
C13956 net35 net71 0.042275f
C13957 FILLER_0_15_212/a_1380_472# FILLER_0_15_228/a_36_472# 0.013277f
C13958 _431_/a_36_151# FILLER_0_16_115/a_36_472# 0.004847f
C13959 FILLER_0_5_206/a_36_472# net22 0.049294f
C13960 _091_ mask\[3\] 0.044304f
C13961 net41 _446_/a_2665_112# 0.004501f
C13962 _053_ FILLER_0_5_54/a_932_472# 0.001578f
C13963 net75 _425_/a_796_472# 0.001146f
C13964 FILLER_0_16_57/a_1468_375# vdd 0.020146f
C13965 FILLER_0_16_57/a_1020_375# vss 0.004487f
C13966 _440_/a_36_151# FILLER_0_6_47/a_3172_472# 0.001653f
C13967 fanout49/a_36_160# FILLER_0_3_78/a_572_375# 0.00805f
C13968 FILLER_0_6_37/a_36_472# _160_ 0.008686f
C13969 _078_ FILLER_0_4_213/a_572_375# 0.02957f
C13970 FILLER_0_16_107/a_124_375# _093_ 0.003941f
C13971 _114_ _428_/a_2665_112# 0.002329f
C13972 net80 FILLER_0_20_177/a_124_375# 0.001198f
C13973 _292_/a_36_160# output18/a_224_472# 0.009736f
C13974 _315_/a_244_497# _059_ 0.00101f
C13975 net57 _267_/a_36_472# 0.032037f
C13976 FILLER_0_22_128/a_572_375# vdd 0.001473f
C13977 net56 FILLER_0_17_161/a_124_375# 0.001108f
C13978 net81 _019_ 0.004079f
C13979 FILLER_0_5_128/a_572_375# net74 0.050735f
C13980 net2 vdd 0.434557f
C13981 _428_/a_36_151# FILLER_0_13_100/a_124_375# 0.023595f
C13982 _415_/a_448_472# net18 0.057688f
C13983 output34/a_224_472# _046_ 0.006059f
C13984 FILLER_0_5_72/a_1380_472# FILLER_0_5_88/a_36_472# 0.013277f
C13985 net64 FILLER_0_12_236/a_124_375# 0.043517f
C13986 FILLER_0_5_198/a_36_472# net21 0.014911f
C13987 _414_/a_1308_423# cal_itt\[3\] 0.044184f
C13988 _436_/a_2665_112# _210_/a_67_603# 0.007103f
C13989 _132_ _022_ 0.001404f
C13990 _441_/a_1000_472# _168_ 0.036305f
C13991 net31 _421_/a_2665_112# 0.005428f
C13992 output17/a_224_472# vdd 0.026649f
C13993 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_36_472# 0.002296f
C13994 _137_ _098_ 0.07262f
C13995 _053_ _151_ 0.538643f
C13996 net63 FILLER_0_20_177/a_1020_375# 0.005919f
C13997 net58 net1 0.626432f
C13998 _115_ net52 0.022268f
C13999 FILLER_0_5_72/a_484_472# _164_ 0.003769f
C14000 net75 _253_/a_672_68# 0.003771f
C14001 _000_ _253_/a_36_68# 0.005121f
C14002 mask\[0\] FILLER_0_14_235/a_572_375# 0.002003f
C14003 _339_/a_36_160# FILLER_0_19_155/a_484_472# 0.00304f
C14004 cal_count\[3\] FILLER_0_11_78/a_36_472# 0.031399f
C14005 _098_ FILLER_0_19_171/a_36_472# 0.021559f
C14006 net47 FILLER_0_5_136/a_36_472# 0.006139f
C14007 trim_mask\[4\] _154_ 0.014658f
C14008 FILLER_0_24_290/a_36_472# vss 0.007621f
C14009 state\[0\] net64 0.01679f
C14010 _428_/a_36_151# net70 0.040167f
C14011 vss FILLER_0_13_290/a_36_472# 0.009561f
C14012 FILLER_0_5_172/a_124_375# vss 0.028247f
C14013 FILLER_0_5_172/a_36_472# vdd 0.092294f
C14014 net41 FILLER_0_8_24/a_572_375# 0.003909f
C14015 FILLER_0_16_57/a_124_375# net15 0.001594f
C14016 mask\[8\] _149_ 0.0498f
C14017 trimb[1] FILLER_0_20_15/a_36_472# 0.001292f
C14018 FILLER_0_18_2/a_1020_375# net38 0.047331f
C14019 _074_ calibrate 0.046632f
C14020 _128_ vss 0.859962f
C14021 _098_ _438_/a_1308_423# 0.004124f
C14022 _126_ _131_ 0.626666f
C14023 _067_ _450_/a_448_472# 0.003113f
C14024 _188_ FILLER_0_12_50/a_124_375# 0.00157f
C14025 _130_ _131_ 0.005955f
C14026 FILLER_0_2_111/a_572_375# _158_ 0.031641f
C14027 net54 FILLER_0_20_98/a_124_375# 0.001639f
C14028 _363_/a_36_68# vss 0.043707f
C14029 net41 net26 0.057852f
C14030 _094_ net62 0.04063f
C14031 ctln[5] net59 0.030363f
C14032 net82 FILLER_0_3_172/a_124_375# 0.011418f
C14033 ctln[1] ctln[4] 0.002283f
C14034 ctln[3] ctln[2] 0.012289f
C14035 net44 net67 0.08001f
C14036 FILLER_0_6_47/a_2724_472# vss 0.020876f
C14037 FILLER_0_6_47/a_3172_472# vdd 0.002089f
C14038 net75 FILLER_0_8_247/a_1020_375# 0.009573f
C14039 _093_ FILLER_0_17_72/a_36_472# 0.001971f
C14040 net63 _137_ 0.006317f
C14041 net52 FILLER_0_5_54/a_1380_472# 0.00179f
C14042 _128_ net74 0.121254f
C14043 trim_mask\[4\] _169_ 0.042442f
C14044 FILLER_0_11_142/a_36_472# vdd 0.110248f
C14045 FILLER_0_11_142/a_572_375# vss 0.052505f
C14046 _114_ _126_ 3.341247f
C14047 FILLER_0_7_146/a_124_375# _059_ 0.029514f
C14048 _149_ vss 0.005314f
C14049 _130_ _114_ 0.002404f
C14050 vdd cal_count\[0\] 0.491891f
C14051 net31 net22 0.002533f
C14052 net81 _429_/a_2248_156# 0.017036f
C14053 FILLER_0_6_239/a_124_375# _122_ 0.01772f
C14054 net53 _040_ 0.035628f
C14055 FILLER_0_3_204/a_36_472# _088_ 0.004381f
C14056 net27 FILLER_0_14_235/a_36_472# 0.003401f
C14057 net81 FILLER_0_10_247/a_36_472# 0.015109f
C14058 FILLER_0_12_236/a_572_375# vdd 0.024713f
C14059 FILLER_0_12_236/a_124_375# vss 0.001024f
C14060 output38/a_224_472# trim[1] 0.003114f
C14061 _418_/a_1000_472# _007_ 0.001051f
C14062 net82 FILLER_0_3_221/a_1468_375# 0.009095f
C14063 net26 FILLER_0_18_37/a_572_375# 0.00109f
C14064 result[6] _420_/a_448_472# 0.017262f
C14065 _132_ FILLER_0_15_116/a_484_472# 0.010148f
C14066 fanout62/a_36_160# _416_/a_36_151# 0.016215f
C14067 _274_/a_3368_68# _069_ 0.001414f
C14068 _104_ _421_/a_448_472# 0.001106f
C14069 FILLER_0_21_125/a_484_472# net54 0.022347f
C14070 _093_ FILLER_0_19_111/a_124_375# 0.00186f
C14071 FILLER_0_15_116/a_572_375# _131_ 0.051323f
C14072 _074_ FILLER_0_6_231/a_36_472# 0.004325f
C14073 _038_ _389_/a_36_148# 0.003749f
C14074 _341_/a_49_472# vss 0.003485f
C14075 _062_ net23 0.061239f
C14076 net17 net6 0.063494f
C14077 net78 vdd 0.265913f
C14078 net60 vdd 0.575502f
C14079 _035_ _380_/a_224_472# 0.001921f
C14080 state\[0\] vss 0.126943f
C14081 output46/a_224_472# FILLER_0_20_2/a_484_472# 0.001699f
C14082 net15 FILLER_0_6_47/a_1828_472# 0.014911f
C14083 FILLER_0_17_72/a_1468_375# net36 0.047507f
C14084 _130_ _428_/a_2665_112# 0.001241f
C14085 output45/a_224_472# net45 0.019483f
C14086 output23/a_224_472# net34 0.021474f
C14087 _359_/a_244_68# _059_ 0.002986f
C14088 net57 FILLER_0_13_142/a_484_472# 0.011685f
C14089 fanout68/a_36_113# net69 0.046009f
C14090 _428_/a_1000_472# _043_ 0.020031f
C14091 _322_/a_848_380# _125_ 0.013667f
C14092 net25 FILLER_0_22_86/a_124_375# 0.004298f
C14093 _077_ _131_ 0.03465f
C14094 _430_/a_2560_156# net63 0.009628f
C14095 _053_ net21 0.036284f
C14096 FILLER_0_4_197/a_932_472# _088_ 0.014643f
C14097 mask\[7\] _297_/a_36_472# 0.003196f
C14098 FILLER_0_21_28/a_3260_375# vss 0.054959f
C14099 FILLER_0_21_28/a_36_472# vdd 0.090954f
C14100 output34/a_224_472# net18 0.126175f
C14101 _052_ _424_/a_1204_472# 0.002681f
C14102 FILLER_0_3_172/a_2724_472# vdd 0.006405f
C14103 net79 _418_/a_448_472# 0.034736f
C14104 FILLER_0_13_212/a_484_472# mask\[0\] 0.001794f
C14105 FILLER_0_8_2/a_36_472# vss 0.004429f
C14106 FILLER_0_16_89/a_124_375# FILLER_0_17_72/a_1916_375# 0.026339f
C14107 _399_/a_224_472# _182_ 0.002729f
C14108 trim_val\[2\] net17 0.019133f
C14109 result[6] _421_/a_796_472# 0.004697f
C14110 result[6] fanout77/a_36_113# 0.001469f
C14111 _232_/a_67_603# _167_ 0.014152f
C14112 _077_ _114_ 0.047702f
C14113 FILLER_0_11_101/a_36_472# _120_ 0.007656f
C14114 _213_/a_67_603# _098_ 0.018092f
C14115 net55 FILLER_0_17_72/a_1828_472# 0.001217f
C14116 _110_ mask\[9\] 0.00319f
C14117 net41 FILLER_0_23_44/a_124_375# 0.001526f
C14118 _391_/a_245_68# cal_count\[0\] 0.001201f
C14119 _144_ _433_/a_2248_156# 0.021805f
C14120 _114_ FILLER_0_10_107/a_124_375# 0.004825f
C14121 net4 _264_/a_224_472# 0.001408f
C14122 mask\[7\] _350_/a_257_69# 0.001135f
C14123 FILLER_0_5_109/a_36_472# _153_ 0.034328f
C14124 _073_ _070_ 0.001892f
C14125 FILLER_0_17_64/a_124_375# vss 0.022351f
C14126 FILLER_0_17_64/a_36_472# vdd 0.094397f
C14127 FILLER_0_4_49/a_124_375# vdd 0.008637f
C14128 _443_/a_2560_156# _170_ 0.00758f
C14129 _443_/a_2248_156# _037_ 0.005717f
C14130 net76 FILLER_0_5_181/a_36_472# 0.014784f
C14131 _035_ _445_/a_36_151# 0.002276f
C14132 net57 _113_ 0.012056f
C14133 _131_ FILLER_0_17_104/a_932_472# 0.002988f
C14134 _426_/a_36_151# FILLER_0_8_247/a_1020_375# 0.059049f
C14135 output8/a_224_472# net58 0.018549f
C14136 vdd _433_/a_36_151# 0.086874f
C14137 _414_/a_36_151# _072_ 0.033026f
C14138 net41 FILLER_0_17_38/a_36_472# 0.001308f
C14139 net56 FILLER_0_18_139/a_572_375# 0.005919f
C14140 _175_ FILLER_0_15_72/a_36_472# 0.006746f
C14141 _428_/a_36_151# FILLER_0_14_107/a_572_375# 0.001597f
C14142 _002_ net59 0.016205f
C14143 FILLER_0_16_89/a_124_375# net53 0.001032f
C14144 FILLER_0_20_177/a_572_375# _434_/a_36_151# 0.059049f
C14145 _412_/a_2560_156# net18 0.015371f
C14146 _130_ _126_ 0.061836f
C14147 FILLER_0_5_109/a_484_472# _163_ 0.005054f
C14148 _139_ mask\[1\] 0.017315f
C14149 _425_/a_36_151# _014_ 0.12681f
C14150 _147_ vdd 0.09215f
C14151 FILLER_0_0_266/a_36_472# vss 0.003738f
C14152 _118_ _311_/a_3220_473# 0.001133f
C14153 net51 _039_ 0.398642f
C14154 net38 _452_/a_2225_156# 0.034415f
C14155 FILLER_0_3_78/a_572_375# vdd 0.014442f
C14156 FILLER_0_3_78/a_124_375# vss 0.004739f
C14157 mask\[9\] FILLER_0_20_107/a_36_472# 0.006047f
C14158 _150_ _027_ 0.006689f
C14159 _431_/a_2560_156# net73 0.001018f
C14160 FILLER_0_8_37/a_572_375# _220_/a_67_603# 0.00744f
C14161 _321_/a_170_472# vdd 0.060585f
C14162 _398_/a_36_113# _178_ 0.004282f
C14163 net3 _095_ 0.002383f
C14164 FILLER_0_13_228/a_36_472# vdd 0.085375f
C14165 FILLER_0_13_228/a_124_375# vss 0.007465f
C14166 _111_ _303_/a_244_68# 0.001153f
C14167 FILLER_0_2_101/a_124_375# vss 0.04897f
C14168 FILLER_0_2_101/a_36_472# vdd 0.099518f
C14169 FILLER_0_4_107/a_1468_375# vdd 0.023541f
C14170 _114_ _267_/a_224_472# 0.001264f
C14171 _093_ vdd 1.439861f
C14172 output47/a_224_472# _398_/a_36_113# 0.001605f
C14173 FILLER_0_11_101/a_572_375# FILLER_0_9_105/a_36_472# 0.0027f
C14174 net20 _418_/a_2665_112# 0.013517f
C14175 _056_ _062_ 0.320621f
C14176 FILLER_0_18_2/a_1020_375# net55 0.003942f
C14177 net76 cal_itt\[1\] 0.027781f
C14178 FILLER_0_24_274/a_484_472# _420_/a_36_151# 0.002841f
C14179 _170_ _037_ 0.05171f
C14180 net57 _118_ 0.036179f
C14181 net34 _107_ 0.017589f
C14182 mask\[5\] _091_ 0.048311f
C14183 _091_ FILLER_0_20_169/a_124_375# 0.003958f
C14184 net68 FILLER_0_8_37/a_484_472# 0.002696f
C14185 net47 _034_ 0.052602f
C14186 _136_ _067_ 0.051914f
C14187 vdd FILLER_0_19_134/a_124_375# 0.027957f
C14188 _063_ vss 0.157186f
C14189 _369_/a_692_472# _157_ 0.0025f
C14190 _331_/a_448_472# _134_ 0.001126f
C14191 _255_/a_224_552# _163_ 0.002169f
C14192 FILLER_0_1_212/a_124_375# net11 0.029766f
C14193 valid net76 0.285892f
C14194 FILLER_0_11_78/a_484_472# _389_/a_36_148# 0.001043f
C14195 FILLER_0_19_47/a_572_375# net55 0.003447f
C14196 _363_/a_692_472# _086_ 0.001353f
C14197 fanout72/a_36_113# _394_/a_56_524# 0.002775f
C14198 ctln[6] FILLER_0_0_130/a_124_375# 0.026786f
C14199 _448_/a_36_151# FILLER_0_2_177/a_572_375# 0.001597f
C14200 FILLER_0_9_290/a_124_375# vdd 0.028723f
C14201 FILLER_0_4_185/a_36_472# net22 0.006506f
C14202 _136_ FILLER_0_14_99/a_124_375# 0.007209f
C14203 net47 FILLER_0_5_164/a_124_375# 0.011983f
C14204 FILLER_0_5_206/a_124_375# vdd 0.038311f
C14205 _139_ vss 0.052996f
C14206 net80 net81 0.006516f
C14207 net65 _412_/a_1204_472# 0.001629f
C14208 _086_ FILLER_0_11_142/a_124_375# 0.009046f
C14209 _128_ FILLER_0_12_236/a_36_472# 0.001043f
C14210 result[8] vss 0.235206f
C14211 FILLER_0_18_100/a_124_375# net14 0.04037f
C14212 _070_ _067_ 0.001869f
C14213 output35/a_224_472# _435_/a_36_151# 0.001362f
C14214 _449_/a_796_472# _067_ 0.004874f
C14215 FILLER_0_12_220/a_932_472# _223_/a_36_160# 0.001323f
C14216 output40/a_224_472# net40 0.0374f
C14217 output31/a_224_472# FILLER_0_16_255/a_124_375# 0.001274f
C14218 FILLER_0_7_195/a_124_375# calibrate 0.00576f
C14219 _033_ _444_/a_1204_472# 0.002294f
C14220 _053_ FILLER_0_6_47/a_1916_375# 0.008103f
C14221 _110_ net35 0.053239f
C14222 _068_ _311_/a_3220_473# 0.004371f
C14223 _149_ _026_ 0.243704f
C14224 output11/a_224_472# vdd 0.01016f
C14225 _235_/a_255_603# trim_mask\[2\] 0.001488f
C14226 _235_/a_67_603# trim_val\[2\] 0.00747f
C14227 FILLER_0_11_142/a_124_375# cal_count\[3\] 0.010782f
C14228 _417_/a_36_151# net30 0.010021f
C14229 _370_/a_692_472# _152_ 0.005908f
C14230 _370_/a_1152_472# _081_ 0.001901f
C14231 _125_ _124_ 0.085897f
C14232 net16 _380_/a_224_472# 0.008718f
C14233 cal_itt\[3\] _375_/a_1612_497# 0.003901f
C14234 _409_/a_245_68# cal_count\[3\] 0.001164f
C14235 _133_ _120_ 0.003762f
C14236 cal_count\[3\] _373_/a_1060_68# 0.00165f
C14237 net81 _100_ 0.24831f
C14238 _445_/a_2248_156# net47 0.028909f
C14239 FILLER_0_4_185/a_124_375# _087_ 0.120668f
C14240 FILLER_0_15_150/a_36_472# fanout53/a_36_160# 0.002059f
C14241 _095_ _098_ 0.057687f
C14242 _158_ vss 0.007784f
C14243 FILLER_0_17_142/a_124_375# vdd 0.020936f
C14244 net28 vdd 0.489756f
C14245 net18 _419_/a_1000_472# 0.008295f
C14246 net57 _068_ 0.029812f
C14247 _436_/a_36_151# vdd 0.078019f
C14248 _091_ _223_/a_36_160# 0.001976f
C14249 FILLER_0_19_47/a_36_472# _424_/a_1308_423# 0.010224f
C14250 _043_ net62 0.00426f
C14251 _430_/a_36_151# mask\[2\] 0.016265f
C14252 net54 FILLER_0_22_86/a_1020_375# 0.001597f
C14253 FILLER_0_16_73/a_124_375# _131_ 0.015859f
C14254 FILLER_0_8_239/a_36_472# _317_/a_36_113# 0.00191f
C14255 vdd _416_/a_2248_156# 0.004325f
C14256 _256_/a_716_497# _128_ 0.001035f
C14257 net27 FILLER_0_9_282/a_484_472# 0.006955f
C14258 result[0] FILLER_0_9_282/a_572_375# 0.042859f
C14259 _367_/a_36_68# _154_ 0.028801f
C14260 net64 FILLER_0_14_235/a_484_472# 0.012355f
C14261 _429_/a_1000_472# vss 0.006901f
C14262 _423_/a_1308_423# vss 0.001726f
C14263 _423_/a_796_472# vdd 0.001494f
C14264 FILLER_0_10_247/a_124_375# vdd 0.040502f
C14265 _086_ net37 0.039329f
C14266 _414_/a_1308_423# _081_ 0.003429f
C14267 FILLER_0_19_28/a_124_375# _452_/a_36_151# 0.002709f
C14268 _178_ cal_count\[2\] 0.119443f
C14269 _346_/a_49_472# vss 0.0031f
C14270 _136_ FILLER_0_16_154/a_572_375# 0.003842f
C14271 net60 net78 0.030634f
C14272 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_124_375# 0.012001f
C14273 output47/a_224_472# cal_count\[2\] 0.080405f
C14274 FILLER_0_4_197/a_1380_472# vss 0.007979f
C14275 net53 FILLER_0_14_99/a_36_472# 0.004153f
C14276 _432_/a_1204_472# vdd 0.004019f
C14277 FILLER_0_17_161/a_124_375# vss 0.00824f
C14278 FILLER_0_17_161/a_36_472# vdd 0.006972f
C14279 _008_ _419_/a_796_472# 0.013039f
C14280 net52 FILLER_0_6_47/a_2364_375# 0.002577f
C14281 _070_ FILLER_0_9_105/a_36_472# 0.023853f
C14282 _333_/a_36_160# mask\[2\] 0.022517f
C14283 FILLER_0_22_86/a_932_472# _098_ 0.001442f
C14284 FILLER_0_14_123/a_124_375# FILLER_0_14_107/a_1468_375# 0.012001f
C14285 output8/a_224_472# _413_/a_2665_112# 0.010726f
C14286 output32/a_224_472# net30 0.001139f
C14287 _424_/a_2665_112# vdd 0.013636f
C14288 _424_/a_2248_156# vss 0.004855f
C14289 _024_ _435_/a_448_472# 0.039244f
C14290 _444_/a_1000_472# net17 0.02064f
C14291 net54 _437_/a_2248_156# 0.046559f
C14292 _027_ _438_/a_448_472# 0.053901f
C14293 _066_ _169_ 0.222791f
C14294 net36 net19 0.031858f
C14295 _040_ FILLER_0_16_115/a_36_472# 0.001876f
C14296 _427_/a_448_472# net23 0.014853f
C14297 net25 FILLER_0_23_88/a_124_375# 0.010782f
C14298 _442_/a_36_151# vdd 0.102701f
C14299 net55 _452_/a_2225_156# 0.022788f
C14300 _031_ trim_mask\[3\] 0.016747f
C14301 fanout62/a_36_160# net79 0.011515f
C14302 _132_ _451_/a_36_151# 0.007777f
C14303 _447_/a_2665_112# vss 0.012813f
C14304 net23 FILLER_0_5_148/a_36_472# 0.011079f
C14305 FILLER_0_18_2/a_2276_472# vdd 0.004679f
C14306 _070_ _121_ 0.285424f
C14307 net82 vss 0.550252f
C14308 _114_ _060_ 0.003352f
C14309 _415_/a_36_151# net81 0.046145f
C14310 net15 _423_/a_36_151# 0.003422f
C14311 FILLER_0_5_109/a_572_375# _160_ 0.004207f
C14312 _083_ cal_itt\[1\] 0.046464f
C14313 output36/a_224_472# output30/a_224_472# 0.003578f
C14314 net32 _104_ 0.342568f
C14315 FILLER_0_4_197/a_1020_375# net76 0.006026f
C14316 FILLER_0_15_290/a_124_375# output30/a_224_472# 0.02894f
C14317 net3 vss 0.02666f
C14318 _411_/a_2665_112# vdd 0.026095f
C14319 FILLER_0_2_93/a_124_375# _030_ 0.001641f
C14320 _386_/a_1152_472# _163_ 0.004076f
C14321 FILLER_0_12_50/a_36_472# _067_ 0.011087f
C14322 vss FILLER_0_14_235/a_484_472# 0.003246f
C14323 output10/a_224_472# rstn 0.001656f
C14324 net82 net74 0.007059f
C14325 output42/a_224_472# net17 0.047757f
C14326 _116_ _162_ 0.00156f
C14327 FILLER_0_11_78/a_36_472# _120_ 0.014169f
C14328 _131_ _330_/a_224_472# 0.001186f
C14329 net41 _402_/a_728_93# 0.032823f
C14330 _077_ _453_/a_36_151# 0.042928f
C14331 _132_ _124_ 0.005668f
C14332 mask\[1\] FILLER_0_15_205/a_124_375# 0.007883f
C14333 _169_ net37 0.03934f
C14334 FILLER_0_14_263/a_124_375# net62 0.037111f
C14335 net64 _098_ 0.281888f
C14336 _129_ _118_ 0.213736f
C14337 mask\[7\] _435_/a_36_151# 0.037736f
C14338 net63 FILLER_0_19_187/a_124_375# 0.012282f
C14339 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_572_375# 0.001597f
C14340 _053_ _062_ 0.185944f
C14341 net35 _049_ 0.022439f
C14342 FILLER_0_16_57/a_1380_472# net55 0.002219f
C14343 cal_itt\[2\] _083_ 0.10423f
C14344 _098_ mask\[1\] 1.476748f
C14345 _069_ mask\[0\] 0.040599f
C14346 FILLER_0_12_20/a_572_375# _039_ 0.005679f
C14347 _144_ _208_/a_36_160# 0.00717f
C14348 output34/a_224_472# _421_/a_2248_156# 0.001144f
C14349 result[7] _421_/a_448_472# 0.018021f
C14350 _390_/a_692_472# _136_ 0.004782f
C14351 net35 _435_/a_2665_112# 0.007912f
C14352 net44 FILLER_0_20_2/a_572_375# 0.002597f
C14353 _073_ net9 0.005417f
C14354 _320_/a_1792_472# _043_ 0.002235f
C14355 _072_ net21 0.062333f
C14356 FILLER_0_21_142/a_124_375# FILLER_0_22_128/a_1828_472# 0.001543f
C14357 result[5] result[6] 0.065361f
C14358 output14/a_224_472# net52 0.02346f
C14359 _132_ FILLER_0_16_107/a_484_472# 0.005391f
C14360 FILLER_0_16_107/a_572_375# _131_ 0.015859f
C14361 FILLER_0_20_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001543f
C14362 _065_ _168_ 0.020406f
C14363 FILLER_0_4_107/a_572_375# _154_ 0.052251f
C14364 _436_/a_448_472# FILLER_0_22_128/a_124_375# 0.006782f
C14365 net36 FILLER_0_16_115/a_124_375# 0.001706f
C14366 _115_ FILLER_0_10_94/a_36_472# 0.014605f
C14367 _072_ _375_/a_960_497# 0.001322f
C14368 FILLER_0_13_142/a_1468_375# _043_ 0.009636f
C14369 net32 _421_/a_1308_423# 0.005394f
C14370 mask\[2\] FILLER_0_16_154/a_36_472# 0.312123f
C14371 FILLER_0_18_2/a_2276_472# _452_/a_1040_527# 0.008652f
C14372 FILLER_0_18_2/a_484_472# _452_/a_2225_156# 0.019521f
C14373 _430_/a_1204_472# net21 0.006991f
C14374 FILLER_0_14_91/a_36_472# _176_ 0.076419f
C14375 mask\[8\] _098_ 0.096999f
C14376 _435_/a_1288_156# vdd 0.001119f
C14377 net76 net59 3.439686f
C14378 result[0] net18 0.085445f
C14379 _085_ state\[1\] 0.182697f
C14380 output46/a_224_472# net40 0.002542f
C14381 net63 net64 0.002181f
C14382 net17 FILLER_0_20_15/a_1468_375# 0.010099f
C14383 _095_ _405_/a_67_603# 0.012596f
C14384 FILLER_0_24_63/a_36_472# output26/a_224_472# 0.023414f
C14385 net76 net4 0.024291f
C14386 net57 vdd 1.260693f
C14387 output33/a_224_472# vdd -0.031734f
C14388 net63 mask\[1\] 0.120872f
C14389 _414_/a_796_472# _003_ 0.006511f
C14390 _414_/a_1000_472# _089_ 0.001754f
C14391 _111_ net36 0.102444f
C14392 FILLER_0_15_205/a_124_375# vss 0.026372f
C14393 FILLER_0_15_205/a_36_472# vdd 0.010089f
C14394 FILLER_0_23_290/a_124_375# net77 0.001783f
C14395 FILLER_0_18_76/a_572_375# net71 0.006025f
C14396 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_484_472# 0.013276f
C14397 _294_/a_224_472# _106_ 0.001038f
C14398 _131_ _095_ 0.043211f
C14399 _132_ net73 0.460325f
C14400 FILLER_0_9_28/a_1828_472# vdd 0.006263f
C14401 FILLER_0_8_107/a_124_375# _131_ 0.001624f
C14402 ctlp[1] FILLER_0_24_274/a_1468_375# 0.01305f
C14403 net36 _280_/a_224_472# 0.001012f
C14404 FILLER_0_14_263/a_36_472# net30 0.003972f
C14405 _098_ vss 0.958032f
C14406 _451_/a_2449_156# _040_ 0.004434f
C14407 trim_mask\[4\] _370_/a_848_380# 0.027744f
C14408 trim_mask\[2\] net14 0.060278f
C14409 FILLER_0_17_56/a_36_472# vss 0.00167f
C14410 FILLER_0_17_56/a_484_472# vdd 0.002789f
C14411 FILLER_0_3_54/a_36_472# _160_ 0.00702f
C14412 _135_ vdd 0.018662f
C14413 net52 FILLER_0_2_111/a_484_472# 0.061249f
C14414 net23 FILLER_0_22_128/a_2364_375# 0.018463f
C14415 FILLER_0_14_99/a_36_472# FILLER_0_14_107/a_36_472# 0.002296f
C14416 _372_/a_2590_472# _076_ 0.002268f
C14417 _129_ _068_ 0.104827f
C14418 net55 _182_ 0.012838f
C14419 net79 _006_ 0.050445f
C14420 _114_ _095_ 0.001338f
C14421 FILLER_0_12_220/a_124_375# _070_ 0.007554f
C14422 _033_ _164_ 0.007117f
C14423 _075_ _074_ 0.058521f
C14424 _444_/a_36_151# net40 0.032012f
C14425 en_co_clk cal_count\[3\] 0.001359f
C14426 FILLER_0_13_212/a_1380_472# vss 0.010223f
C14427 FILLER_0_17_72/a_484_472# _131_ 0.002672f
C14428 net42 net6 0.166896f
C14429 FILLER_0_4_185/a_124_375# vdd 0.02924f
C14430 _425_/a_1308_423# net19 0.058462f
C14431 _115_ _070_ 0.890903f
C14432 FILLER_0_4_152/a_36_472# net57 0.015332f
C14433 FILLER_0_18_139/a_1020_375# vdd 0.001285f
C14434 FILLER_0_18_139/a_572_375# vss 0.009977f
C14435 trim[2] output41/a_224_472# 0.005452f
C14436 output40/a_224_472# trim[3] 0.122003f
C14437 FILLER_0_1_204/a_124_375# net59 0.00999f
C14438 _086_ _395_/a_1044_488# 0.001091f
C14439 net65 FILLER_0_3_172/a_124_375# 0.021073f
C14440 FILLER_0_12_2/a_484_472# net38 0.002706f
C14441 net63 vss 0.566021f
C14442 net20 FILLER_0_9_223/a_484_472# 0.002601f
C14443 _016_ state\[2\] 0.002937f
C14444 _132_ FILLER_0_19_111/a_484_472# 0.004619f
C14445 result[9] _094_ 0.03984f
C14446 _369_/a_36_68# _153_ 0.008048f
C14447 FILLER_0_24_130/a_36_472# ctlp[6] 0.005932f
C14448 _445_/a_2665_112# trim_val\[1\] 0.015206f
C14449 _428_/a_2665_112# _095_ 0.001471f
C14450 net15 FILLER_0_17_56/a_124_375# 0.001854f
C14451 result[7] FILLER_0_24_274/a_484_472# 0.006641f
C14452 _091_ FILLER_0_12_220/a_572_375# 0.003075f
C14453 net68 FILLER_0_3_54/a_124_375# 0.022559f
C14454 mask\[7\] FILLER_0_22_128/a_3260_375# 0.00186f
C14455 _116_ _373_/a_244_68# 0.001213f
C14456 _144_ FILLER_0_18_107/a_2364_375# 0.002388f
C14457 net39 _444_/a_1000_472# 0.001323f
C14458 FILLER_0_10_78/a_484_472# _439_/a_36_151# 0.00271f
C14459 _077_ _426_/a_2665_112# 0.001392f
C14460 _067_ FILLER_0_12_28/a_124_375# 0.012779f
C14461 output24/a_224_472# net54 0.177947f
C14462 net65 FILLER_0_3_221/a_1468_375# 0.001695f
C14463 net35 FILLER_0_22_128/a_2724_472# 0.012359f
C14464 fanout68/a_36_113# vss 0.006152f
C14465 net41 net17 0.911377f
C14466 net36 _451_/a_2225_156# 0.044144f
C14467 net20 _429_/a_1308_423# 0.001186f
C14468 net68 FILLER_0_6_47/a_484_472# 0.005391f
C14469 output18/a_224_472# ctlp[1] 0.039734f
C14470 FILLER_0_18_61/a_124_375# FILLER_0_18_53/a_572_375# 0.012001f
C14471 FILLER_0_18_171/a_36_472# vss 0.0032f
C14472 output38/a_224_472# _034_ 0.039873f
C14473 FILLER_0_9_72/a_1468_375# _439_/a_2248_156# 0.001901f
C14474 _115_ FILLER_0_9_142/a_36_472# 0.00336f
C14475 _028_ _439_/a_796_472# 0.013039f
C14476 result[6] net19 0.834308f
C14477 _057_ net57 0.873864f
C14478 trim_mask\[1\] FILLER_0_6_47/a_1380_472# 0.006166f
C14479 _093_ FILLER_0_19_134/a_124_375# 0.003473f
C14480 net56 _137_ 0.0313f
C14481 _343_/a_49_472# vdd 0.089707f
C14482 FILLER_0_22_128/a_3172_472# vss 0.006339f
C14483 FILLER_0_7_72/a_2724_472# net14 0.012436f
C14484 result[9] FILLER_0_24_274/a_572_375# 0.003576f
C14485 net76 FILLER_0_5_198/a_124_375# 0.006974f
C14486 output42/a_224_472# net39 0.027208f
C14487 net70 FILLER_0_13_100/a_36_472# 0.00585f
C14488 _406_/a_36_159# net17 0.053547f
C14489 _421_/a_36_151# net19 0.016842f
C14490 _446_/a_1000_472# vdd 0.001598f
C14491 FILLER_0_9_28/a_484_472# net51 0.001023f
C14492 net16 _408_/a_728_93# 0.107634f
C14493 net55 _040_ 0.107198f
C14494 FILLER_0_20_193/a_484_472# _205_/a_36_160# 0.001684f
C14495 FILLER_0_5_72/a_1020_375# vss 0.004157f
C14496 FILLER_0_5_72/a_1468_375# vdd 0.001826f
C14497 _086_ _122_ 0.033097f
C14498 FILLER_0_12_136/a_124_375# state\[2\] 0.001029f
C14499 FILLER_0_12_136/a_1020_375# net53 0.002709f
C14500 _036_ _168_ 0.01699f
C14501 net80 _140_ 0.188514f
C14502 FILLER_0_16_57/a_484_472# FILLER_0_17_56/a_572_375# 0.001723f
C14503 output37/a_224_472# fanout64/a_36_160# 0.017421f
C14504 _050_ net23 0.003752f
C14505 _186_ _043_ 0.045082f
C14506 _083_ net59 0.408831f
C14507 _077_ _330_/a_224_472# 0.001921f
C14508 FILLER_0_7_72/a_1020_375# FILLER_0_5_72/a_932_472# 0.001512f
C14509 FILLER_0_1_98/a_124_375# net14 0.049552f
C14510 FILLER_0_21_28/a_3172_472# _424_/a_36_151# 0.001723f
C14511 _413_/a_2560_156# net21 0.002416f
C14512 FILLER_0_10_28/a_36_472# net17 0.012954f
C14513 _174_ net15 0.090215f
C14514 _174_ _180_ 0.102241f
C14515 trim[4] vdd 0.198218f
C14516 _096_ _085_ 0.0099f
C14517 net4 _083_ 0.135165f
C14518 _086_ _311_/a_2180_473# 0.001744f
C14519 _408_/a_1336_472# vdd 0.040992f
C14520 _073_ _084_ 0.048469f
C14521 net63 FILLER_0_18_177/a_1828_472# 0.047684f
C14522 _115_ FILLER_0_11_78/a_572_375# 0.034089f
C14523 _067_ _039_ 0.221585f
C14524 FILLER_0_15_142/a_36_472# _095_ 0.001526f
C14525 _186_ _185_ 0.007962f
C14526 _195_/a_67_603# _045_ 0.004028f
C14527 net82 FILLER_0_3_172/a_3172_472# 0.007677f
C14528 trim_val\[1\] FILLER_0_6_37/a_36_472# 0.011347f
C14529 _139_ _019_ 0.094494f
C14530 _405_/a_67_603# vss 0.008564f
C14531 _405_/a_255_603# vdd 0.001044f
C14532 _150_ mask\[9\] 0.162185f
C14533 _105_ _104_ 0.931514f
C14534 _093_ FILLER_0_17_142/a_124_375# 0.009328f
C14535 output46/a_224_472# net46 0.008691f
C14536 net20 calibrate 0.044792f
C14537 net41 FILLER_0_16_37/a_36_472# 0.009425f
C14538 _372_/a_170_472# vss 0.027819f
C14539 FILLER_0_11_142/a_124_375# _120_ 0.036088f
C14540 _129_ vdd 0.314544f
C14541 _094_ _418_/a_2560_156# 0.011088f
C14542 _131_ vss 0.549133f
C14543 FILLER_0_15_116/a_572_375# _095_ 0.00152f
C14544 FILLER_0_5_72/a_124_375# net15 0.006403f
C14545 _086_ _061_ 0.152228f
C14546 net52 _441_/a_448_472# 0.04874f
C14547 _028_ FILLER_0_7_72/a_2276_472# 0.001777f
C14548 net72 FILLER_0_20_31/a_36_472# 0.002751f
C14549 ctln[1] net5 0.050549f
C14550 FILLER_0_20_177/a_572_375# mask\[6\] 0.001158f
C14551 result[9] FILLER_0_23_274/a_36_472# 0.0064f
C14552 fanout63/a_36_160# FILLER_0_15_228/a_36_472# 0.014197f
C14553 _273_/a_36_68# _223_/a_36_160# 0.002786f
C14554 result[6] _009_ 0.095754f
C14555 net52 _440_/a_1204_472# 0.003916f
C14556 _176_ _134_ 0.035146f
C14557 _061_ cal_count\[3\] 0.003415f
C14558 _104_ _010_ 0.252687f
C14559 net74 _372_/a_170_472# 0.079123f
C14560 _114_ vss 0.365613f
C14561 _131_ net74 0.227843f
C14562 net52 _439_/a_36_151# 0.01388f
C14563 output44/a_224_472# FILLER_0_18_2/a_572_375# 0.001296f
C14564 _122_ _169_ 0.014463f
C14565 calibrate _163_ 0.026892f
C14566 net52 _157_ 0.005889f
C14567 _053_ FILLER_0_7_72/a_484_472# 0.00887f
C14568 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_36_472# 0.002296f
C14569 _050_ _025_ 0.033887f
C14570 mask\[4\] FILLER_0_18_177/a_2812_375# 0.013557f
C14571 FILLER_0_20_15/a_1380_472# vss 0.003678f
C14572 _026_ _098_ 0.197713f
C14573 net55 FILLER_0_19_28/a_572_375# 0.002115f
C14574 net7 net17 0.050676f
C14575 _077_ FILLER_0_8_107/a_124_375# 0.010439f
C14576 FILLER_0_18_209/a_484_472# _201_/a_67_603# 0.001605f
C14577 _010_ _420_/a_36_151# 0.001838f
C14578 _421_/a_36_151# _009_ 0.00246f
C14579 _434_/a_36_151# vdd 0.104871f
C14580 FILLER_0_5_212/a_124_375# _081_ 0.01149f
C14581 FILLER_0_18_107/a_2276_472# _137_ 0.001752f
C14582 _274_/a_2552_68# vss 0.003123f
C14583 _093_ FILLER_0_17_161/a_36_472# 0.006224f
C14584 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001723f
C14585 net20 FILLER_0_6_231/a_36_472# 0.045553f
C14586 _114_ net74 0.559239f
C14587 _098_ FILLER_0_21_206/a_124_375# 0.001882f
C14588 _131_ cal_count\[1\] 0.001497f
C14589 net69 FILLER_0_2_111/a_572_375# 0.015789f
C14590 state\[2\] _043_ 0.028842f
C14591 _093_ _424_/a_2665_112# 0.001854f
C14592 _098_ _097_ 0.034041f
C14593 output33/a_224_472# net60 0.002526f
C14594 _065_ _447_/a_36_151# 0.043351f
C14595 _133_ FILLER_0_10_107/a_484_472# 0.001798f
C14596 net18 _044_ 0.174456f
C14597 net32 result[7] 0.103491f
C14598 net79 _007_ 0.096772f
C14599 _428_/a_2665_112# vss 0.005991f
C14600 FILLER_0_5_54/a_36_472# vdd 0.006056f
C14601 FILLER_0_5_54/a_1468_375# vss 0.053407f
C14602 _072_ _062_ 0.025795f
C14603 FILLER_0_14_50/a_36_472# _181_ 0.001514f
C14604 FILLER_0_20_31/a_124_375# net40 0.011967f
C14605 _075_ FILLER_0_7_195/a_124_375# 0.008178f
C14606 _004_ net62 0.001201f
C14607 clk vss 0.210484f
C14608 _441_/a_36_151# _164_ 0.008955f
C14609 trimb[1] net43 0.004299f
C14610 FILLER_0_7_72/a_2724_472# FILLER_0_6_90/a_572_375# 0.001684f
C14611 net29 FILLER_0_16_255/a_36_472# 0.086886f
C14612 _096_ _320_/a_224_472# 0.001285f
C14613 _440_/a_2665_112# FILLER_0_5_88/a_124_375# 0.02132f
C14614 FILLER_0_14_91/a_124_375# _136_ 0.013064f
C14615 _238_/a_67_603# net50 0.002229f
C14616 FILLER_0_4_177/a_484_472# vss 0.002399f
C14617 _432_/a_2248_156# _139_ 0.002904f
C14618 FILLER_0_12_2/a_36_472# clkc 0.004826f
C14619 _415_/a_1000_472# net19 0.001125f
C14620 _136_ _138_ 0.186242f
C14621 FILLER_0_21_28/a_3172_472# FILLER_0_21_60/a_36_472# 0.013276f
C14622 _428_/a_2665_112# net74 0.048822f
C14623 _256_/a_36_68# _056_ 0.008305f
C14624 net20 FILLER_0_13_212/a_484_472# 0.001273f
C14625 net44 output6/a_224_472# 0.078248f
C14626 _282_/a_36_160# mask\[2\] 0.023533f
C14627 ctln[1] FILLER_0_1_266/a_572_375# 0.004319f
C14628 _141_ _145_ 0.094128f
C14629 net55 FILLER_0_18_76/a_484_472# 0.003745f
C14630 _322_/a_124_24# _118_ 0.04952f
C14631 _443_/a_2665_112# vss 0.007913f
C14632 _414_/a_2248_156# FILLER_0_5_212/a_36_472# 0.035805f
C14633 net1 _084_ 0.008356f
C14634 net41 net39 0.003649f
C14635 net16 FILLER_0_17_38/a_124_375# 0.046435f
C14636 FILLER_0_16_241/a_124_375# _198_/a_67_603# 0.002082f
C14637 net55 _423_/a_2665_112# 0.002379f
C14638 FILLER_0_7_72/a_36_472# net50 0.011974f
C14639 FILLER_0_7_72/a_932_472# net52 0.008749f
C14640 mask\[9\] _012_ 0.008145f
C14641 FILLER_0_19_28/a_484_472# net40 0.020293f
C14642 net81 FILLER_0_15_212/a_572_375# 0.006974f
C14643 result[1] _416_/a_1000_472# 0.001529f
C14644 net28 _416_/a_2248_156# 0.001082f
C14645 net20 FILLER_0_17_226/a_124_375# 0.001895f
C14646 mask\[0\] net22 0.054097f
C14647 net38 _398_/a_36_113# 0.061273f
C14648 _446_/a_36_151# output41/a_224_472# 0.135198f
C14649 _074_ net22 0.079421f
C14650 net70 FILLER_0_14_107/a_1020_375# 0.011157f
C14651 net27 _426_/a_2248_156# 0.002303f
C14652 _431_/a_2248_156# net36 0.001441f
C14653 net15 FILLER_0_5_54/a_572_375# 0.002259f
C14654 FILLER_0_18_2/a_3260_375# FILLER_0_19_28/a_484_472# 0.001684f
C14655 output12/a_224_472# net12 0.007193f
C14656 _248_/a_36_68# _060_ 0.004581f
C14657 net22 _204_/a_67_603# 0.006495f
C14658 net81 mask\[0\] 0.320022f
C14659 _159_ _081_ 0.003646f
C14660 net65 net64 0.119915f
C14661 FILLER_0_16_57/a_36_472# _131_ 0.00864f
C14662 fanout73/a_36_113# net70 0.00238f
C14663 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_484_472# 0.013277f
C14664 FILLER_0_5_109/a_124_375# net47 0.010784f
C14665 output46/a_224_472# FILLER_0_20_15/a_1020_375# 0.001274f
C14666 ctlp[4] vss 0.102044f
C14667 net16 FILLER_0_18_37/a_1380_472# 0.002932f
C14668 net15 FILLER_0_15_72/a_484_472# 0.002925f
C14669 _219_/a_36_160# vdd 0.013125f
C14670 mask\[3\] FILLER_0_16_241/a_124_375# 0.006824f
C14671 net20 FILLER_0_16_241/a_36_472# 0.001528f
C14672 _098_ _433_/a_448_472# 0.027678f
C14673 _126_ vss 0.399848f
C14674 net50 net15 0.177988f
C14675 FILLER_0_3_2/a_124_375# vdd 0.021963f
C14676 net17 _450_/a_448_472# 0.017832f
C14677 _130_ vss 0.090346f
C14678 cal_itt\[2\] _253_/a_672_68# 0.0016f
C14679 _091_ FILLER_0_18_177/a_1020_375# 0.002226f
C14680 _027_ vdd 0.146607f
C14681 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2724_472# 0.026657f
C14682 _140_ _434_/a_448_472# 0.00128f
C14683 net34 FILLER_0_22_177/a_1468_375# 0.006974f
C14684 net36 FILLER_0_15_180/a_36_472# 0.007275f
C14685 result[2] vss 0.327009f
C14686 _159_ FILLER_0_2_127/a_124_375# 0.020951f
C14687 ctlp[1] _419_/a_2248_156# 0.028734f
C14688 mask\[9\] _438_/a_448_472# 0.046823f
C14689 FILLER_0_10_78/a_932_472# FILLER_0_9_72/a_1468_375# 0.001543f
C14690 _412_/a_2248_156# vdd 0.005671f
C14691 _238_/a_67_603# trim_mask\[3\] 0.028437f
C14692 _037_ vdd 0.158731f
C14693 FILLER_0_3_172/a_1020_375# net22 0.013048f
C14694 output42/a_224_472# net42 0.117956f
C14695 FILLER_0_19_55/a_36_472# net55 0.062683f
C14696 FILLER_0_15_142/a_484_472# vdd 0.001097f
C14697 FILLER_0_15_142/a_36_472# vss 0.006166f
C14698 _126_ net74 1.001749f
C14699 ctlp[3] vdd 0.251098f
C14700 net48 _082_ 0.003853f
C14701 _056_ FILLER_0_12_196/a_36_472# 0.039555f
C14702 FILLER_0_17_72/a_1380_472# _438_/a_36_151# 0.001221f
C14703 _130_ net74 0.001655f
C14704 trim_val\[2\] _160_ 0.051804f
C14705 _433_/a_2665_112# _145_ 0.018359f
C14706 FILLER_0_18_37/a_932_472# vdd 0.01019f
C14707 trimb[2] net17 0.007637f
C14708 FILLER_0_15_142/a_124_375# _427_/a_36_151# 0.059049f
C14709 FILLER_0_0_96/a_36_472# trim_mask\[3\] 0.005343f
C14710 FILLER_0_7_195/a_36_472# _072_ 0.008357f
C14711 mask\[5\] net23 0.002188f
C14712 _322_/a_848_380# _076_ 0.006699f
C14713 net76 FILLER_0_2_177/a_36_472# 0.003526f
C14714 FILLER_0_14_91/a_572_375# net53 0.063988f
C14715 FILLER_0_15_116/a_36_472# vdd 0.013454f
C14716 FILLER_0_15_142/a_36_472# net74 0.003166f
C14717 _236_/a_36_160# vdd 0.023428f
C14718 _119_ _372_/a_170_472# 0.003159f
C14719 _119_ _131_ 0.073868f
C14720 cal_itt\[3\] net76 0.017174f
C14721 _044_ net62 0.101165f
C14722 _412_/a_36_151# net76 0.001169f
C14723 FILLER_0_14_107/a_932_472# _043_ 0.0017f
C14724 net65 vss 0.471168f
C14725 _448_/a_2560_156# _037_ 0.011661f
C14726 _127_ FILLER_0_11_124/a_36_472# 0.001641f
C14727 FILLER_0_4_144/a_484_472# trim_mask\[4\] 0.015778f
C14728 _436_/a_2248_156# mask\[7\] 0.003615f
C14729 _427_/a_2665_112# net36 0.009904f
C14730 _198_/a_67_603# _046_ 0.007349f
C14731 net49 net40 0.093233f
C14732 net34 net19 0.039959f
C14733 _429_/a_2665_112# FILLER_0_14_235/a_36_472# 0.007491f
C14734 _436_/a_1000_472# _025_ 0.061189f
C14735 FILLER_0_17_38/a_36_472# _452_/a_36_151# 0.096503f
C14736 _441_/a_2248_156# _030_ 0.003495f
C14737 trim_mask\[2\] net49 0.041781f
C14738 _064_ net66 0.304028f
C14739 _140_ _022_ 0.001997f
C14740 net56 _095_ 0.004847f
C14741 _095_ FILLER_0_13_142/a_932_472# 0.001782f
C14742 _077_ vss 1.071923f
C14743 _119_ _114_ 0.001581f
C14744 _074_ _076_ 0.03553f
C14745 net68 net40 0.036106f
C14746 _019_ _098_ 0.010193f
C14747 _137_ mask\[1\] 0.782055f
C14748 ctlp[6] ctlp[7] 0.002504f
C14749 _093_ FILLER_0_18_139/a_1020_375# 0.003529f
C14750 FILLER_0_10_107/a_124_375# vss 0.003015f
C14751 FILLER_0_10_107/a_572_375# vdd 0.043678f
C14752 trim_mask\[2\] net68 0.099597f
C14753 en_co_clk _120_ 0.008507f
C14754 _445_/a_1204_472# net40 0.003916f
C14755 _116_ _055_ 0.72331f
C14756 net48 _265_/a_244_68# 0.00365f
C14757 input5/a_36_113# vdd 0.026855f
C14758 FILLER_0_3_142/a_124_375# _443_/a_36_151# 0.059049f
C14759 FILLER_0_15_235/a_124_375# FILLER_0_15_228/a_124_375# 0.002868f
C14760 _064_ _445_/a_1308_423# 0.01485f
C14761 _447_/a_1308_423# net68 0.006686f
C14762 _447_/a_36_151# _036_ 0.007244f
C14763 FILLER_0_7_72/a_2812_375# _077_ 0.002969f
C14764 net79 FILLER_0_11_282/a_36_472# 0.004358f
C14765 net18 net77 0.378783f
C14766 net35 _012_ 0.007543f
C14767 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_36_472# 0.001723f
C14768 FILLER_0_20_177/a_1468_375# vdd 0.016422f
C14769 result[9] FILLER_0_14_263/a_124_375# 0.003706f
C14770 output32/a_224_472# _418_/a_2665_112# 0.011048f
C14771 output19/a_224_472# net33 0.126671f
C14772 _077_ net74 0.025882f
C14773 mask\[3\] _046_ 0.018595f
C14774 net38 _054_ 0.640545f
C14775 _091_ FILLER_0_15_212/a_36_472# 0.007355f
C14776 FILLER_0_1_212/a_124_375# FILLER_0_1_204/a_124_375# 0.003732f
C14777 net48 _112_ 0.284235f
C14778 _053_ fanout67/a_36_160# 0.05724f
C14779 net80 _139_ 0.178583f
C14780 _053_ _153_ 0.015583f
C14781 ctln[2] FILLER_0_0_266/a_124_375# 0.041898f
C14782 calibrate FILLER_0_9_270/a_124_375# 0.002292f
C14783 net38 cal_count\[2\] 0.047195f
C14784 _114_ _097_ 0.004412f
C14785 ctlp[9] net26 0.02213f
C14786 _028_ FILLER_0_6_90/a_484_472# 0.01566f
C14787 net38 FILLER_0_8_24/a_36_472# 0.015829f
C14788 FILLER_0_10_78/a_124_375# net52 0.008557f
C14789 FILLER_0_4_144/a_124_375# vss 0.017638f
C14790 FILLER_0_4_144/a_572_375# vdd -0.013698f
C14791 _073_ FILLER_0_6_231/a_36_472# 0.001898f
C14792 _011_ _109_ 0.055905f
C14793 FILLER_0_17_104/a_1380_472# vdd 0.010877f
C14794 result[9] _419_/a_1000_472# 0.012469f
C14795 _050_ FILLER_0_22_107/a_36_472# 0.001098f
C14796 net63 _019_ 0.004471f
C14797 mask\[5\] net33 0.251971f
C14798 _411_/a_36_151# net75 0.033786f
C14799 net26 FILLER_0_21_28/a_2364_375# 0.003691f
C14800 _419_/a_1308_423# vdd 0.007543f
C14801 _136_ _451_/a_1353_112# 0.058703f
C14802 _086_ FILLER_0_4_177/a_36_472# 0.001464f
C14803 _343_/a_49_472# _093_ 0.001926f
C14804 net52 FILLER_0_9_72/a_36_472# 0.014911f
C14805 _137_ vss 0.343959f
C14806 FILLER_0_15_59/a_484_472# vdd 0.010447f
C14807 FILLER_0_15_59/a_36_472# vss 0.00459f
C14808 net20 _274_/a_36_68# 0.021022f
C14809 _453_/a_36_151# vss 0.007105f
C14810 _453_/a_448_472# vdd 0.010005f
C14811 _098_ FILLER_0_18_76/a_124_375# 0.001831f
C14812 net10 FILLER_0_0_232/a_124_375# 0.022977f
C14813 comp net3 0.05248f
C14814 _345_/a_36_160# net71 0.002396f
C14815 net54 FILLER_0_20_107/a_124_375# 0.072539f
C14816 net22 _201_/a_67_603# 0.004491f
C14817 _375_/a_36_68# _162_ 0.011065f
C14818 _375_/a_1612_497# _161_ 0.003325f
C14819 net63 FILLER_0_19_195/a_124_375# 0.017284f
C14820 _076_ FILLER_0_3_221/a_484_472# 0.001225f
C14821 FILLER_0_19_171/a_484_472# vdd 0.009225f
C14822 FILLER_0_19_171/a_36_472# vss 0.001338f
C14823 _377_/a_36_472# trim_val\[0\] 0.135527f
C14824 net69 vss 0.34555f
C14825 _425_/a_36_151# calibrate 0.071513f
C14826 FILLER_0_9_28/a_1916_375# _220_/a_67_603# 0.014522f
C14827 net34 _009_ 0.325819f
C14828 _087_ _088_ 0.001219f
C14829 net59 FILLER_0_3_212/a_36_472# 0.058623f
C14830 FILLER_0_24_96/a_36_472# net35 0.002526f
C14831 _394_/a_728_93# _174_ 0.012471f
C14832 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_572_375# 0.086635f
C14833 _011_ _422_/a_448_472# 0.044695f
C14834 net74 net69 0.143604f
C14835 _360_/a_36_160# FILLER_0_4_123/a_36_472# 0.001165f
C14836 _055_ _117_ 0.242156f
C14837 mask\[4\] _047_ 0.080091f
C14838 cal_count\[1\] FILLER_0_15_59/a_36_472# 0.00544f
C14839 FILLER_0_18_177/a_3172_472# FILLER_0_18_209/a_36_472# 0.013276f
C14840 net15 FILLER_0_15_59/a_124_375# 0.007439f
C14841 _180_ FILLER_0_15_59/a_124_375# 0.009926f
C14842 FILLER_0_9_28/a_2812_375# net68 0.012462f
C14843 net73 FILLER_0_18_107/a_1380_472# 0.039646f
C14844 output43/a_224_472# net40 0.014984f
C14845 FILLER_0_19_125/a_36_472# vss 0.001056f
C14846 net16 _450_/a_2225_156# 0.001015f
C14847 _133_ _062_ 1.210949f
C14848 mask\[7\] _208_/a_36_160# 0.105845f
C14849 output34/a_224_472# net61 0.008309f
C14850 _432_/a_1000_472# net80 0.033803f
C14851 _430_/a_2560_156# vss 0.002924f
C14852 net47 _386_/a_124_24# 0.024696f
C14853 _322_/a_124_24# vdd 0.01572f
C14854 net80 FILLER_0_17_161/a_124_375# 0.021914f
C14855 _321_/a_170_472# _129_ 0.024601f
C14856 _122_ _120_ 0.143427f
C14857 output26/a_224_472# FILLER_0_23_44/a_484_472# 0.0323f
C14858 result[8] FILLER_0_24_274/a_124_375# 0.00726f
C14859 _395_/a_36_488# _121_ 0.009689f
C14860 FILLER_0_6_47/a_1020_375# vdd 0.016637f
C14861 net50 _163_ 0.068547f
C14862 result[7] _010_ 0.054533f
C14863 FILLER_0_15_212/a_124_375# vdd -0.004549f
C14864 _311_/a_1212_473# _117_ 0.001673f
C14865 _449_/a_36_151# FILLER_0_13_72/a_124_375# 0.059049f
C14866 FILLER_0_3_204/a_124_375# _413_/a_36_151# 0.035849f
C14867 _155_ FILLER_0_4_107/a_124_375# 0.00162f
C14868 _432_/a_2248_156# net63 0.047337f
C14869 _196_/a_36_160# vdd 0.106963f
C14870 _426_/a_2665_112# net64 0.01548f
C14871 _420_/a_2560_156# vdd 0.001652f
C14872 _420_/a_2665_112# vss 0.001749f
C14873 net2 input5/a_36_113# 0.007518f
C14874 input2/a_36_113# net5 0.001761f
C14875 net77 net62 0.122747f
C14876 output31/a_224_472# _094_ 0.004668f
C14877 vdd _450_/a_3129_107# 0.039939f
C14878 net53 _451_/a_1040_527# 0.023651f
C14879 _147_ _434_/a_36_151# 0.001817f
C14880 _258_/a_36_160# net37 0.006865f
C14881 net64 _060_ 0.05104f
C14882 _360_/a_36_160# _153_ 0.006561f
C14883 mask\[8\] _213_/a_67_603# 0.039626f
C14884 net19 _419_/a_2665_112# 0.00276f
C14885 FILLER_0_17_104/a_572_375# net14 0.004285f
C14886 output12/a_224_472# vss 0.013728f
C14887 FILLER_0_18_2/a_3172_472# _041_ 0.001503f
C14888 en_co_clk _390_/a_244_472# 0.001238f
C14889 net56 vss 0.367812f
C14890 FILLER_0_13_142/a_1380_472# vdd 0.001977f
C14891 FILLER_0_13_142/a_932_472# vss 0.005192f
C14892 _017_ _134_ 0.017998f
C14893 net67 net6 0.345681f
C14894 fanout66/a_36_113# FILLER_0_3_54/a_124_375# 0.002853f
C14895 _077_ FILLER_0_9_72/a_124_375# 0.008103f
C14896 _119_ _077_ 2.584241f
C14897 FILLER_0_17_72/a_2276_472# _136_ 0.055635f
C14898 net82 _370_/a_124_24# 0.001011f
C14899 _413_/a_36_151# FILLER_0_4_197/a_484_472# 0.001512f
C14900 net20 _008_ 0.153014f
C14901 FILLER_0_6_239/a_124_375# vdd 0.031271f
C14902 _213_/a_67_603# vss 0.019344f
C14903 _210_/a_67_603# mask\[7\] 0.039004f
C14904 FILLER_0_5_88/a_124_375# FILLER_0_6_90/a_36_472# 0.001543f
C14905 FILLER_0_16_73/a_124_375# vss 0.026383f
C14906 FILLER_0_16_73/a_572_375# vdd 0.005054f
C14907 _177_ _451_/a_2449_156# 0.002085f
C14908 net55 cal_count\[2\] 0.022989f
C14909 _248_/a_36_68# vss 0.027935f
C14910 _276_/a_36_160# vss 0.02914f
C14911 ctln[5] _448_/a_1000_472# 0.007584f
C14912 FILLER_0_3_172/a_572_375# vdd 0.007121f
C14913 net27 vdd 0.88294f
C14914 _065_ fanout50/a_36_160# 0.022932f
C14915 _422_/a_1204_472# vdd 0.001062f
C14916 _165_ vss 0.048027f
C14917 _449_/a_36_151# net72 0.039436f
C14918 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001597f
C14919 _426_/a_2665_112# vss 0.006288f
C14920 FILLER_0_10_78/a_1020_375# _176_ 0.020379f
C14921 FILLER_0_5_117/a_36_472# _360_/a_36_160# 0.003913f
C14922 trim_mask\[0\] net14 0.499565f
C14923 _427_/a_2665_112# _225_/a_36_160# 0.001394f
C14924 FILLER_0_4_107/a_572_375# _151_ 0.00162f
C14925 _064_ _446_/a_2665_112# 0.039211f
C14926 _446_/a_448_472# net66 0.017696f
C14927 _060_ vss 0.318005f
C14928 FILLER_0_24_96/a_36_472# ctlp[7] 0.001551f
C14929 trimb[4] vss 0.039934f
C14930 FILLER_0_6_177/a_36_472# net47 0.011891f
C14931 _058_ _117_ 0.003932f
C14932 _114_ _389_/a_36_148# 0.009465f
C14933 _167_ _160_ 0.157458f
C14934 _112_ _316_/a_1152_472# 0.001449f
C14935 _445_/a_2665_112# _444_/a_448_472# 0.001178f
C14936 _432_/a_36_151# mask\[3\] 0.002148f
C14937 FILLER_0_3_221/a_36_472# vdd 0.018263f
C14938 FILLER_0_3_221/a_1468_375# vss 0.004085f
C14939 net25 _214_/a_36_160# 0.019894f
C14940 net65 FILLER_0_3_172/a_3172_472# 0.001777f
C14941 ctln[4] FILLER_0_0_232/a_124_375# 0.002726f
C14942 _122_ _227_/a_36_160# 0.005128f
C14943 FILLER_0_17_38/a_572_375# _179_ 0.002825f
C14944 FILLER_0_5_72/a_1020_375# _029_ 0.010208f
C14945 _086_ _267_/a_36_472# 0.070088f
C14946 net80 _098_ 1.289178f
C14947 mask\[9\] FILLER_0_19_111/a_124_375# 0.031474f
C14948 _239_/a_36_160# net41 0.006002f
C14949 net26 _423_/a_36_151# 0.067024f
C14950 _413_/a_796_472# net59 0.006163f
C14951 FILLER_0_17_200/a_36_472# vdd 0.001039f
C14952 net12 vss 0.043754f
C14953 _059_ FILLER_0_8_156/a_124_375# 0.00593f
C14954 _431_/a_448_472# _136_ 0.064724f
C14955 net37 net21 0.03272f
C14956 _174_ _067_ 0.002678f
C14957 _184_ net40 0.122833f
C14958 _093_ _027_ 0.047164f
C14959 FILLER_0_2_111/a_1020_375# vdd 0.007918f
C14960 ctln[6] net13 0.065837f
C14961 output44/a_224_472# FILLER_0_19_28/a_124_375# 0.005166f
C14962 _065_ _383_/a_36_472# 0.02518f
C14963 _095_ mask\[1\] 0.001297f
C14964 _137_ _097_ 0.001654f
C14965 _283_/a_36_472# net62 0.002309f
C14966 net26 _424_/a_1000_472# 0.003207f
C14967 FILLER_0_18_107/a_2724_472# vdd 0.004677f
C14968 _103_ _419_/a_448_472# 0.001207f
C14969 net78 _419_/a_1308_423# 0.018598f
C14970 _052_ vdd 0.264744f
C14971 net61 _419_/a_1000_472# 0.017712f
C14972 net60 _419_/a_1308_423# 0.029697f
C14973 FILLER_0_24_130/a_36_472# vdd 0.050082f
C14974 FILLER_0_24_130/a_124_375# vss 0.018125f
C14975 net76 _081_ 0.706096f
C14976 _322_/a_848_380# _128_ 0.012288f
C14977 net63 net80 0.337396f
C14978 _300_/a_224_472# _011_ 0.007508f
C14979 mask\[6\] vdd 0.573103f
C14980 _216_/a_67_603# net36 0.028132f
C14981 _417_/a_2248_156# _006_ 0.039121f
C14982 FILLER_0_16_89/a_1380_472# _040_ 0.008446f
C14983 ctln[8] FILLER_0_0_96/a_124_375# 0.002726f
C14984 net32 output35/a_224_472# 0.072991f
C14985 output43/a_224_472# net46 0.0215f
C14986 FILLER_0_11_109/a_124_375# _134_ 0.027704f
C14987 _088_ vdd 0.140259f
C14988 _079_ vss 0.124667f
C14989 _320_/a_36_472# net79 0.029189f
C14990 FILLER_0_16_107/a_572_375# vss 0.055104f
C14991 FILLER_0_16_107/a_36_472# vdd 0.110244f
C14992 _000_ _083_ 0.017601f
C14993 _053_ trim_mask\[1\] 0.110786f
C14994 FILLER_0_6_79/a_124_375# vss 0.007008f
C14995 FILLER_0_6_79/a_36_472# vdd 0.087807f
C14996 FILLER_0_12_136/a_1020_375# net23 0.005919f
C14997 net55 _177_ 0.327874f
C14998 fanout58/a_36_160# net5 0.003758f
C14999 FILLER_0_17_133/a_124_375# vdd 0.010519f
C15000 net20 FILLER_0_15_235/a_36_472# 0.002227f
C15001 net52 _160_ 0.133292f
C15002 ctln[4] FILLER_0_1_212/a_36_472# 0.006408f
C15003 _308_/a_124_24# trim_mask\[0\] 0.018998f
C15004 _115_ _439_/a_2665_112# 0.003617f
C15005 _074_ FILLER_0_5_172/a_124_375# 0.068565f
C15006 FILLER_0_14_81/a_124_375# _095_ 0.009791f
C15007 cal_count\[2\] FILLER_0_15_10/a_36_472# 0.015502f
C15008 net55 FILLER_0_17_38/a_484_472# 0.013624f
C15009 _126_ _389_/a_36_148# 0.007813f
C15010 FILLER_0_18_171/a_36_472# net80 0.041571f
C15011 _095_ vss 1.465527f
C15012 _270_/a_36_472# net76 0.009569f
C15013 FILLER_0_13_65/a_36_472# _095_ 0.003171f
C15014 FILLER_0_11_101/a_124_375# net14 0.011983f
C15015 FILLER_0_8_107/a_124_375# vss 0.031335f
C15016 FILLER_0_8_107/a_36_472# vdd 0.117254f
C15017 _284_/a_224_472# _094_ 0.001731f
C15018 FILLER_0_18_107/a_2812_375# _145_ 0.030158f
C15019 net66 FILLER_0_5_54/a_572_375# 0.002203f
C15020 net47 net40 0.635497f
C15021 _423_/a_36_151# FILLER_0_23_44/a_124_375# 0.059049f
C15022 en_co_clk _043_ 0.041355f
C15023 _450_/a_1284_156# _039_ 0.001226f
C15024 _450_/a_3129_107# cal_count\[0\] 0.020971f
C15025 _430_/a_2248_156# net20 0.001893f
C15026 _132_ net54 0.016007f
C15027 FILLER_0_18_177/a_2724_472# net22 0.004297f
C15028 FILLER_0_8_138/a_36_472# _120_ 0.006759f
C15029 net54 FILLER_0_22_107/a_484_472# 0.005897f
C15030 FILLER_0_5_54/a_124_375# trim_mask\[1\] 0.024065f
C15031 FILLER_0_5_54/a_1468_375# _029_ 0.008339f
C15032 _304_/a_224_472# _111_ 0.003461f
C15033 _449_/a_2665_112# vss 0.007395f
C15034 net74 _095_ 0.04188f
C15035 mask\[9\] vdd 0.940144f
C15036 net50 net66 0.016385f
C15037 net52 _030_ 0.035783f
C15038 net41 _160_ 0.006523f
C15039 net35 FILLER_0_22_86/a_484_472# 0.008347f
C15040 mask\[8\] FILLER_0_22_86/a_932_472# 0.012284f
C15041 net52 _442_/a_1204_472# 0.005558f
C15042 _256_/a_36_68# _072_ 0.027152f
C15043 net17 _452_/a_36_151# 0.041497f
C15044 _162_ FILLER_0_6_177/a_124_375# 0.031168f
C15045 FILLER_0_17_72/a_484_472# vss 0.005334f
C15046 net7 _239_/a_36_160# 0.068281f
C15047 net15 _038_ 0.078028f
C15048 _150_ FILLER_0_18_76/a_572_375# 0.008337f
C15049 FILLER_0_16_89/a_932_472# net36 0.001709f
C15050 net60 _420_/a_2560_156# 0.001358f
C15051 _093_ FILLER_0_17_104/a_1380_472# 0.014431f
C15052 _068_ FILLER_0_5_148/a_124_375# 0.003986f
C15053 net18 FILLER_0_9_270/a_572_375# 0.005977f
C15054 _449_/a_2665_112# net74 0.001185f
C15055 _095_ cal_count\[1\] 0.853949f
C15056 net64 mask\[1\] 0.038611f
C15057 _164_ _166_ 0.002368f
C15058 output18/a_224_472# net33 0.135766f
C15059 FILLER_0_22_86/a_1380_472# vdd 0.008224f
C15060 FILLER_0_22_86/a_932_472# vss -0.001553f
C15061 FILLER_0_19_111/a_572_375# vss 0.003337f
C15062 FILLER_0_19_111/a_36_472# vdd 0.034386f
C15063 _013_ FILLER_0_18_53/a_124_375# 0.015996f
C15064 FILLER_0_7_59/a_124_375# trim_val\[0\] 0.002169f
C15065 FILLER_0_19_187/a_572_375# vdd 0.023383f
C15066 FILLER_0_18_107/a_36_472# net14 0.005297f
C15067 mask\[3\] fanout53/a_36_160# 0.001205f
C15068 _449_/a_1204_472# net15 0.01349f
C15069 net69 FILLER_0_3_78/a_36_472# 0.002068f
C15070 _086_ _113_ 0.072034f
C15071 FILLER_0_3_204/a_36_472# net21 0.01535f
C15072 net14 FILLER_0_10_94/a_572_375# 0.047331f
C15073 net27 FILLER_0_12_236/a_572_375# 0.083731f
C15074 _258_/a_36_160# _122_ 0.00102f
C15075 _015_ FILLER_0_8_247/a_124_375# 0.00706f
C15076 result[4] _008_ 0.134001f
C15077 _031_ FILLER_0_2_101/a_124_375# 0.00179f
C15078 _106_ mask\[4\] 0.091207f
C15079 net17 FILLER_0_12_28/a_124_375# 0.009108f
C15080 _093_ _438_/a_796_472# 0.001924f
C15081 cal_count\[3\] _113_ 0.093684f
C15082 _098_ _434_/a_448_472# 0.015893f
C15083 _079_ _260_/a_244_472# 0.00325f
C15084 _070_ _319_/a_234_472# 0.004015f
C15085 net41 _187_ 0.002046f
C15086 state\[2\] _427_/a_448_472# 0.00237f
C15087 net53 _427_/a_796_472# 0.001983f
C15088 _444_/a_1000_472# net67 0.025169f
C15089 FILLER_0_12_236/a_36_472# _060_ 0.014046f
C15090 net57 _428_/a_2560_156# 0.010877f
C15091 net61 _422_/a_2665_112# 0.023601f
C15092 FILLER_0_18_2/a_124_375# vdd 0.008721f
C15093 net32 mask\[7\] 0.01969f
C15094 FILLER_0_16_255/a_124_375# vdd 0.029925f
C15095 net64 vss 0.636644f
C15096 _440_/a_1308_423# vdd 0.00218f
C15097 _440_/a_448_472# vss 0.032037f
C15098 FILLER_0_18_2/a_3172_472# FILLER_0_18_37/a_36_472# 0.002765f
C15099 trim_mask\[1\] _164_ 0.195956f
C15100 _083_ _081_ 0.03934f
C15101 _359_/a_36_488# _152_ 0.032195f
C15102 _128_ _124_ 0.111918f
C15103 mask\[1\] vss 0.46268f
C15104 _028_ FILLER_0_7_104/a_484_472# 0.00499f
C15105 FILLER_0_4_197/a_932_472# net21 0.00663f
C15106 _115_ _125_ 0.049021f
C15107 net34 _435_/a_1000_472# 0.007444f
C15108 vss FILLER_0_4_91/a_484_472# 0.003328f
C15109 net20 FILLER_0_3_221/a_572_375# 0.004331f
C15110 net36 FILLER_0_15_235/a_124_375# 0.007232f
C15111 _086_ _118_ 0.166544f
C15112 _402_/a_1296_93# _179_ 0.001692f
C15113 comp _190_/a_36_160# 0.001891f
C15114 _142_ vdd 0.090938f
C15115 output42/a_224_472# net67 0.05585f
C15116 _352_/a_49_472# vdd 0.077542f
C15117 net63 _434_/a_448_472# 0.008139f
C15118 output39/a_224_472# vdd 0.022593f
C15119 _053_ FILLER_0_7_104/a_572_375# 0.005239f
C15120 ctln[9] vss 0.167242f
C15121 FILLER_0_10_214/a_124_375# _247_/a_36_160# 0.005732f
C15122 cal_count\[3\] _118_ 0.009058f
C15123 FILLER_0_12_20/a_484_472# _450_/a_448_472# 0.04564f
C15124 FILLER_0_17_142/a_572_375# _137_ 0.006974f
C15125 mask\[8\] vss 0.378558f
C15126 net35 vdd 1.0365f
C15127 _086_ _087_ 0.015938f
C15128 _098_ _022_ 0.013131f
C15129 FILLER_0_2_111/a_124_375# _154_ 0.004032f
C15130 _423_/a_1204_472# _012_ 0.003181f
C15131 net17 _039_ 0.079171f
C15132 _422_/a_2665_112# _108_ 0.023365f
C15133 _430_/a_1000_472# net36 0.001836f
C15134 _412_/a_796_472# net1 0.002922f
C15135 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3172_472# 0.013276f
C15136 net20 net81 0.036173f
C15137 _140_ _023_ 0.079452f
C15138 trim_mask\[2\] fanout66/a_36_113# 0.015961f
C15139 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_484_472# 0.013276f
C15140 _081_ FILLER_0_5_136/a_124_375# 0.025819f
C15141 net79 _101_ 0.014383f
C15142 FILLER_0_14_81/a_124_375# vss 0.03341f
C15143 FILLER_0_14_81/a_36_472# vdd 0.00958f
C15144 _031_ _158_ 0.015116f
C15145 _085_ _176_ 0.024708f
C15146 _337_/a_49_472# mask\[2\] 0.00188f
C15147 FILLER_0_22_86/a_572_375# net14 0.009573f
C15148 _163_ net22 0.005017f
C15149 _306_/a_36_68# _085_ 0.00755f
C15150 net79 FILLER_0_12_220/a_1468_375# 0.012754f
C15151 FILLER_0_13_65/a_36_472# vss 0.007545f
C15152 FILLER_0_14_50/a_124_375# _095_ 0.052375f
C15153 _448_/a_448_472# net59 0.050956f
C15154 _365_/a_36_68# vdd 0.004308f
C15155 _053_ _414_/a_1308_423# 0.029387f
C15156 _122_ net21 0.026632f
C15157 mask\[7\] FILLER_0_22_177/a_572_375# 0.001315f
C15158 FILLER_0_0_96/a_124_375# vdd 0.034959f
C15159 FILLER_0_7_72/a_3260_375# vdd 0.008342f
C15160 net16 _180_ 0.00101f
C15161 _432_/a_2248_156# _137_ 0.001775f
C15162 _326_/a_36_160# _058_ 0.003897f
C15163 vdd FILLER_0_5_148/a_124_375# -0.011369f
C15164 _062_ FILLER_0_8_156/a_484_472# 0.006123f
C15165 net74 vss 0.589483f
C15166 FILLER_0_13_65/a_36_472# net74 0.014937f
C15167 _104_ _107_ 0.021508f
C15168 result[6] FILLER_0_21_286/a_484_472# 0.011149f
C15169 net53 net14 0.04525f
C15170 _062_ net37 0.082701f
C15171 mask\[5\] FILLER_0_19_171/a_572_375# 0.007169f
C15172 output48/a_224_472# net37 0.095886f
C15173 _086_ _068_ 0.080666f
C15174 FILLER_0_10_78/a_1380_472# _115_ 0.051132f
C15175 _144_ _145_ 0.671767f
C15176 _105_ output35/a_224_472# 0.013092f
C15177 _437_/a_1204_472# net14 0.004949f
C15178 FILLER_0_14_81/a_124_375# cal_count\[1\] 0.070473f
C15179 _053_ _054_ 0.015389f
C15180 _359_/a_36_488# _070_ 0.028563f
C15181 FILLER_0_13_212/a_932_472# _043_ 0.014431f
C15182 _095_ _097_ 0.030222f
C15183 net79 _417_/a_796_472# 0.001042f
C15184 _088_ FILLER_0_3_172/a_2724_472# 0.005827f
C15185 net68 _220_/a_255_603# 0.001908f
C15186 _059_ _313_/a_67_603# 0.061666f
C15187 cal_count\[1\] vss 0.307993f
C15188 FILLER_0_13_65/a_36_472# cal_count\[1\] 0.016393f
C15189 _435_/a_2665_112# net21 0.067461f
C15190 output22/a_224_472# net22 0.032714f
C15191 FILLER_0_17_38/a_572_375# _041_ 0.021754f
C15192 _449_/a_2248_156# cal_count\[3\] 0.002041f
C15193 net28 _196_/a_36_160# 0.060575f
C15194 output15/a_224_472# fanout50/a_36_160# 0.003531f
C15195 _293_/a_36_472# _092_ 0.004828f
C15196 result[4] result[3] 0.089939f
C15197 _061_ net21 0.049282f
C15198 _442_/a_448_472# net69 0.004308f
C15199 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1468_375# 0.016748f
C15200 net27 FILLER_0_9_290/a_124_375# 0.002657f
C15201 _069_ _121_ 0.137961f
C15202 net48 cal_itt\[0\] 0.006171f
C15203 _445_/a_2560_156# net49 0.001208f
C15204 ctln[1] cal 0.123834f
C15205 _106_ net34 0.013009f
C15206 _429_/a_36_151# FILLER_0_15_212/a_484_472# 0.001723f
C15207 net34 FILLER_0_22_128/a_1380_472# 0.001011f
C15208 FILLER_0_4_152/a_124_375# FILLER_0_5_148/a_572_375# 0.05841f
C15209 net20 _076_ 0.228128f
C15210 FILLER_0_9_28/a_2276_472# _077_ 0.003256f
C15211 FILLER_0_17_200/a_36_472# _093_ 0.005101f
C15212 _016_ _428_/a_2248_156# 0.048889f
C15213 ctln[2] net8 0.057281f
C15214 FILLER_0_22_86/a_932_472# _026_ 0.001587f
C15215 net56 FILLER_0_17_142/a_572_375# 0.014948f
C15216 net16 net51 0.035455f
C15217 mask\[0\] _429_/a_1000_472# 0.020553f
C15218 FILLER_0_4_107/a_484_472# FILLER_0_2_111/a_124_375# 0.001404f
C15219 net4 state\[1\] 0.010195f
C15220 net55 FILLER_0_18_53/a_36_472# 0.00953f
C15221 _181_ _185_ 0.061846f
C15222 _321_/a_2590_472# _118_ 0.002396f
C15223 FILLER_0_18_177/a_1828_472# vss -0.001107f
C15224 FILLER_0_18_177/a_2276_472# vdd 0.005211f
C15225 _328_/a_36_113# _017_ 0.006485f
C15226 _147_ mask\[6\] 0.103475f
C15227 net72 FILLER_0_21_28/a_1020_375# 0.040811f
C15228 _076_ _163_ 0.030003f
C15229 FILLER_0_20_177/a_36_472# _098_ 0.015061f
C15230 net35 FILLER_0_22_128/a_572_375# 0.010439f
C15231 _093_ FILLER_0_18_107/a_2724_472# 0.00308f
C15232 _044_ FILLER_0_13_290/a_124_375# 0.001855f
C15233 ctlp[7] vdd 0.481613f
C15234 FILLER_0_4_123/a_36_472# trim_mask\[4\] 0.003692f
C15235 input2/a_36_113# en 0.002108f
C15236 FILLER_0_5_128/a_484_472# vss 0.004051f
C15237 net41 net67 0.03408f
C15238 FILLER_0_4_144/a_572_375# net57 0.001254f
C15239 _077_ FILLER_0_9_105/a_124_375# 0.007189f
C15240 _256_/a_2124_68# _070_ 0.002444f
C15241 _256_/a_1612_497# _076_ 0.001111f
C15242 net75 _425_/a_1204_472# 0.015778f
C15243 _042_ vdd 0.261947f
C15244 _136_ _334_/a_36_160# 0.005574f
C15245 FILLER_0_16_57/a_484_472# vdd 0.005894f
C15246 FILLER_0_16_57/a_36_472# vss 0.003789f
C15247 _058_ _059_ 0.990213f
C15248 output15/a_224_472# _383_/a_36_472# 0.001154f
C15249 fanout49/a_36_160# FILLER_0_3_78/a_484_472# 0.003699f
C15250 _078_ FILLER_0_4_213/a_484_472# 0.003702f
C15251 FILLER_0_16_107/a_36_472# _093_ 0.001526f
C15252 net50 FILLER_0_8_24/a_572_375# 0.001597f
C15253 FILLER_0_18_100/a_36_472# FILLER_0_17_72/a_3172_472# 0.05841f
C15254 _427_/a_2248_156# state\[1\] 0.001849f
C15255 _260_/a_36_68# vdd 0.011119f
C15256 net57 _267_/a_672_472# 0.004637f
C15257 FILLER_0_22_128/a_1020_375# vss 0.003747f
C15258 FILLER_0_22_128/a_1468_375# vdd 0.016807f
C15259 FILLER_0_5_128/a_484_472# net74 0.025425f
C15260 _093_ FILLER_0_17_133/a_124_375# 0.009649f
C15261 _074_ net82 0.123449f
C15262 _155_ net50 0.012085f
C15263 net64 FILLER_0_12_236/a_36_472# 0.052381f
C15264 _414_/a_1000_472# cal_itt\[3\] 0.08528f
C15265 FILLER_0_9_28/a_2276_472# _453_/a_36_151# 0.059367f
C15266 net27 FILLER_0_10_247/a_124_375# 0.015466f
C15267 FILLER_0_15_290/a_124_375# net79 0.051113f
C15268 FILLER_0_2_93/a_572_375# net14 0.044606f
C15269 _115_ net50 0.008628f
C15270 net66 _382_/a_224_472# 0.001902f
C15271 FILLER_0_5_72/a_1380_472# _164_ 0.049427f
C15272 _099_ mask\[2\] 0.776725f
C15273 _097_ mask\[1\] 0.001232f
C15274 mask\[0\] FILLER_0_14_235/a_484_472# 0.004688f
C15275 output38/a_224_472# net40 0.072234f
C15276 FILLER_0_19_47/a_572_375# _013_ 0.012993f
C15277 output27/a_224_472# FILLER_0_9_270/a_124_375# 0.001274f
C15278 _098_ FILLER_0_19_171/a_932_472# 0.003573f
C15279 _088_ FILLER_0_5_206/a_124_375# 0.001374f
C15280 _079_ FILLER_0_5_206/a_36_472# 0.008243f
C15281 _428_/a_36_151# _017_ 0.021229f
C15282 FILLER_0_21_28/a_1020_375# _424_/a_36_151# 0.001252f
C15283 FILLER_0_21_28/a_572_375# net40 0.001406f
C15284 FILLER_0_16_57/a_36_472# cal_count\[1\] 0.002116f
C15285 net80 _137_ 0.260786f
C15286 FILLER_0_16_57/a_1020_375# net15 0.048731f
C15287 mask\[8\] _026_ 0.001638f
C15288 trimb[1] FILLER_0_20_15/a_932_472# 0.001069f
C15289 FILLER_0_18_2/a_1916_375# net38 0.006403f
C15290 _098_ _438_/a_1000_472# 0.001492f
C15291 _413_/a_2665_112# ctln[4] 0.001394f
C15292 _067_ _450_/a_1040_527# 0.007414f
C15293 FILLER_0_14_50/a_36_472# vdd 0.081414f
C15294 FILLER_0_14_50/a_124_375# vss 0.002412f
C15295 _105_ mask\[7\] 0.486236f
C15296 FILLER_0_9_72/a_124_375# vss 0.047932f
C15297 FILLER_0_9_72/a_572_375# vdd -0.014642f
C15298 _011_ _108_ 0.036521f
C15299 _152_ _160_ 0.286108f
C15300 _093_ mask\[9\] 0.460108f
C15301 net82 FILLER_0_3_172/a_1020_375# 0.010679f
C15302 _119_ vss 0.22921f
C15303 _086_ vdd 1.212255f
C15304 net80 FILLER_0_19_171/a_36_472# 0.040915f
C15305 net75 _082_ 0.417366f
C15306 net20 output20/a_224_472# 0.024692f
C15307 FILLER_0_18_139/a_1468_375# _137_ 0.004111f
C15308 _136_ net36 1.151311f
C15309 FILLER_0_4_123/a_36_472# fanout69/a_36_113# 0.007864f
C15310 FILLER_0_15_150/a_36_472# FILLER_0_15_142/a_572_375# 0.086635f
C15311 FILLER_0_16_37/a_124_375# _179_ 0.005434f
C15312 net75 FILLER_0_8_247/a_36_472# 0.002992f
C15313 _093_ FILLER_0_17_72/a_932_472# 0.004367f
C15314 _269_/a_36_472# vss 0.014227f
C15315 mask\[4\] FILLER_0_18_209/a_572_375# 0.032112f
C15316 _299_/a_36_472# _109_ 0.030751f
C15317 output18/a_224_472# net18 0.01698f
C15318 _028_ FILLER_0_7_72/a_124_375# 0.017052f
C15319 _115_ _069_ 0.022355f
C15320 FILLER_0_11_142/a_484_472# vss 0.033416f
C15321 _414_/a_448_472# _075_ 0.020304f
C15322 _026_ vss 0.005992f
C15323 ctln[6] _170_ 0.005146f
C15324 trim[4] _236_/a_36_160# 0.004514f
C15325 cal_count\[3\] vdd 1.020669f
C15326 _131_ FILLER_0_18_37/a_1380_472# 0.035078f
C15327 net81 _429_/a_2560_156# 0.003888f
C15328 net18 _417_/a_448_472# 0.03772f
C15329 _119_ net74 0.02813f
C15330 FILLER_0_12_236/a_36_472# vss 0.001526f
C15331 FILLER_0_12_236/a_484_472# vdd 0.00923f
C15332 net63 FILLER_0_19_171/a_932_472# 0.00128f
C15333 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_124_375# 0.007947f
C15334 net32 _292_/a_36_160# 0.011466f
C15335 net75 _426_/a_448_472# 0.041705f
C15336 FILLER_0_21_206/a_36_472# vdd 0.00971f
C15337 FILLER_0_21_206/a_124_375# vss 0.05074f
C15338 FILLER_0_16_89/a_572_375# _136_ 0.069752f
C15339 net82 FILLER_0_3_221/a_484_472# 0.013492f
C15340 result[6] _420_/a_796_472# 0.002296f
C15341 _097_ vss 0.00839f
C15342 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_124_375# 0.005439f
C15343 FILLER_0_15_116/a_484_472# _131_ 0.042796f
C15344 _098_ FILLER_0_15_212/a_572_375# 0.009099f
C15345 FILLER_0_17_142/a_124_375# FILLER_0_17_133/a_124_375# 0.003228f
C15346 _154_ vdd 0.639978f
C15347 _350_/a_257_69# net23 0.003052f
C15348 FILLER_0_14_50/a_124_375# cal_count\[1\] 0.023752f
C15349 _091_ FILLER_0_17_218/a_124_375# 0.013726f
C15350 net81 FILLER_0_9_270/a_124_375# 0.014206f
C15351 _356_/a_36_472# net36 0.004539f
C15352 _103_ vss 0.098913f
C15353 _423_/a_36_151# net17 0.002865f
C15354 _443_/a_36_151# _032_ 0.0737f
C15355 net69 _370_/a_124_24# 0.001491f
C15356 _316_/a_124_24# net37 0.011141f
C15357 FILLER_0_23_88/a_36_472# net14 0.003077f
C15358 net15 FILLER_0_6_47/a_2724_472# 0.006158f
C15359 FILLER_0_17_72/a_2364_375# net36 0.005483f
C15360 _002_ FILLER_0_4_197/a_36_472# 0.006574f
C15361 output45/a_224_472# trimb[2] 0.045907f
C15362 net57 FILLER_0_13_142/a_1380_472# 0.011768f
C15363 FILLER_0_12_124/a_36_472# _428_/a_36_151# 0.001723f
C15364 _428_/a_2248_156# _043_ 0.011841f
C15365 _096_ FILLER_0_15_180/a_572_375# 0.001972f
C15366 _343_/a_257_69# _137_ 0.003494f
C15367 net75 _265_/a_244_68# 0.046186f
C15368 _098_ _204_/a_67_603# 0.00539f
C15369 _008_ _417_/a_36_151# 0.001136f
C15370 _052_ _424_/a_2665_112# 0.003027f
C15371 FILLER_0_21_28/a_932_472# vdd 0.04815f
C15372 FILLER_0_3_172/a_3172_472# vss 0.003689f
C15373 _211_/a_36_160# vss 0.002041f
C15374 FILLER_0_5_88/a_36_472# net47 0.003953f
C15375 _169_ vdd 0.055642f
C15376 net29 _195_/a_67_603# 0.048817f
C15377 FILLER_0_13_212/a_1380_472# mask\[0\] 0.002361f
C15378 cal_itt\[3\] net47 0.00247f
C15379 FILLER_0_16_89/a_572_375# FILLER_0_17_72/a_2364_375# 0.026339f
C15380 mask\[4\] FILLER_0_19_171/a_124_375# 0.001988f
C15381 net75 _112_ 0.041092f
C15382 net23 FILLER_0_21_150/a_36_472# 0.016375f
C15383 _064_ net17 0.108825f
C15384 net79 state\[1\] 0.005861f
C15385 result[6] _421_/a_1204_472# 0.005361f
C15386 net63 FILLER_0_15_212/a_572_375# 0.001597f
C15387 FILLER_0_4_107/a_124_375# _157_ 0.001427f
C15388 FILLER_0_4_107/a_1380_472# trim_mask\[4\] 0.011766f
C15389 _035_ net66 1.624557f
C15390 _112_ _425_/a_1000_472# 0.001973f
C15391 _144_ _433_/a_2560_156# 0.01064f
C15392 fanout58/a_36_160# en 0.00568f
C15393 _114_ FILLER_0_10_107/a_36_472# 0.00263f
C15394 net81 _425_/a_36_151# 0.014663f
C15395 _073_ _076_ 0.011358f
C15396 FILLER_0_10_78/a_36_472# _453_/a_2665_112# 0.007491f
C15397 _181_ _402_/a_1296_93# 0.040412f
C15398 _070_ _160_ 0.065914f
C15399 FILLER_0_4_49/a_36_472# vdd 0.090733f
C15400 FILLER_0_4_49/a_572_375# vss 0.008729f
C15401 net33 _297_/a_36_472# 0.00521f
C15402 _122_ _062_ 0.190871f
C15403 _142_ _093_ 0.492191f
C15404 _086_ _057_ 0.82902f
C15405 output21/a_224_472# net32 0.017976f
C15406 net76 FILLER_0_3_172/a_932_472# 0.005391f
C15407 net36 _045_ 0.091033f
C15408 _426_/a_36_151# FILLER_0_8_247/a_36_472# 0.001723f
C15409 ctln[1] net75 0.159105f
C15410 fanout63/a_36_160# _282_/a_36_160# 0.23939f
C15411 _413_/a_2665_112# FILLER_0_3_212/a_124_375# 0.001077f
C15412 vss _433_/a_448_472# 0.005349f
C15413 _116_ _070_ 0.166494f
C15414 net56 FILLER_0_18_139/a_1468_375# 0.065206f
C15415 _093_ net35 0.00127f
C15416 FILLER_0_20_177/a_1468_375# _434_/a_36_151# 0.001822f
C15417 _020_ _136_ 0.022753f
C15418 _057_ cal_count\[3\] 0.416063f
C15419 net81 net1 0.03613f
C15420 fanout64/a_36_160# fanout65/a_36_113# 0.001627f
C15421 _379_/a_36_472# vdd 0.004183f
C15422 net25 FILLER_0_23_44/a_1380_472# 0.0014f
C15423 _019_ mask\[1\] 0.007797f
C15424 fanout82/a_36_113# net19 0.021188f
C15425 _042_ cal_count\[0\] 0.006265f
C15426 FILLER_0_21_142/a_36_472# net23 0.001629f
C15427 FILLER_0_3_78/a_36_472# vss 0.004461f
C15428 net72 _424_/a_448_472# 0.011745f
C15429 net72 net40 0.001815f
C15430 output32/a_224_472# _008_ 0.074809f
C15431 _431_/a_1456_156# net73 0.001304f
C15432 FILLER_0_8_37/a_484_472# _220_/a_67_603# 0.005759f
C15433 mask\[9\] _424_/a_2665_112# 0.015491f
C15434 mask\[3\] FILLER_0_18_177/a_484_472# 0.005654f
C15435 _118_ _120_ 0.339442f
C15436 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_124_375# 0.009654f
C15437 output36/a_224_472# output29/a_224_472# 0.007726f
C15438 output6/a_224_472# net6 0.076605f
C15439 net15 FILLER_0_17_64/a_124_375# 0.047331f
C15440 FILLER_0_4_107/a_36_472# vss 0.002634f
C15441 FILLER_0_4_107/a_484_472# vdd 0.03151f
C15442 vdd _278_/a_36_160# 0.016488f
C15443 _417_/a_448_472# net62 0.011318f
C15444 net53 FILLER_0_14_123/a_36_472# 0.062713f
C15445 net67 _450_/a_448_472# 0.068692f
C15446 FILLER_0_12_20/a_124_375# vdd 0.017452f
C15447 net61 net77 0.986569f
C15448 _061_ _062_ 0.344031f
C15449 FILLER_0_18_2/a_1916_375# net55 0.008235f
C15450 output46/a_224_472# net38 0.003296f
C15451 _053_ FILLER_0_5_212/a_124_375# 0.048501f
C15452 _038_ _067_ 0.503045f
C15453 vss FILLER_0_19_134/a_36_472# 0.005204f
C15454 _376_/a_36_160# trim_mask\[1\] 0.003111f
C15455 FILLER_0_19_47/a_484_472# net55 0.061087f
C15456 FILLER_0_19_171/a_484_472# _434_/a_36_151# 0.002841f
C15457 FILLER_0_5_128/a_572_375# _163_ 0.007391f
C15458 _322_/a_124_24# _129_ 0.017754f
C15459 _429_/a_36_151# FILLER_0_13_206/a_124_375# 0.001597f
C15460 _448_/a_448_472# FILLER_0_2_177/a_36_472# 0.001927f
C15461 _448_/a_36_151# FILLER_0_2_177/a_484_472# 0.059367f
C15462 FILLER_0_9_290/a_36_472# vss 0.011755f
C15463 net47 FILLER_0_5_164/a_36_472# 0.046908f
C15464 _394_/a_1336_472# vdd 0.003226f
C15465 FILLER_0_5_206/a_36_472# vss 0.003493f
C15466 _019_ vss 0.10954f
C15467 _142_ FILLER_0_17_142/a_124_375# 0.011387f
C15468 net42 _039_ 0.001096f
C15469 net38 _444_/a_36_151# 0.009033f
C15470 FILLER_0_10_247/a_36_472# net64 0.059367f
C15471 _086_ FILLER_0_11_142/a_36_472# 0.006774f
C15472 _449_/a_1204_472# _067_ 0.014354f
C15473 _436_/a_36_151# _352_/a_49_472# 0.005127f
C15474 FILLER_0_15_2/a_124_375# vdd 0.010829f
C15475 output40/a_224_472# trim[2] 0.025041f
C15476 _081_ _265_/a_468_472# 0.005156f
C15477 _412_/a_448_472# output37/a_224_472# 0.001155f
C15478 _033_ _444_/a_2665_112# 0.004024f
C15479 FILLER_0_12_2/a_572_375# vdd 0.022401f
C15480 net32 ctlp[2] 0.097138f
C15481 _053_ FILLER_0_6_47/a_2812_375# 0.003818f
C15482 _058_ _134_ 0.034211f
C15483 _070_ _117_ 0.080445f
C15484 _050_ net71 0.033192f
C15485 _436_/a_36_151# net35 0.014669f
C15486 FILLER_0_19_195/a_124_375# vss 0.020433f
C15487 FILLER_0_19_195/a_36_472# vdd 0.094409f
C15488 _013_ _182_ 0.001681f
C15489 _235_/a_67_603# _064_ 0.003796f
C15490 net52 _453_/a_2248_156# 0.011419f
C15491 FILLER_0_11_142/a_36_472# cal_count\[3\] 0.008454f
C15492 _417_/a_36_151# result[3] 0.006379f
C15493 _417_/a_1308_423# net30 0.007538f
C15494 net20 _128_ 0.041f
C15495 cal_count\[3\] cal_count\[0\] 0.098735f
C15496 FILLER_0_18_2/a_2812_375# net40 0.018463f
C15497 FILLER_0_16_57/a_932_472# FILLER_0_17_64/a_124_375# 0.001723f
C15498 trim[0] output41/a_224_472# 0.018464f
C15499 vss _295_/a_36_472# 0.009751f
C15500 _432_/a_2248_156# mask\[1\] 0.002293f
C15501 _447_/a_2248_156# _441_/a_36_151# 0.035837f
C15502 _068_ _120_ 0.447243f
C15503 _389_/a_36_148# vss 0.001935f
C15504 trim_mask\[2\] _447_/a_448_472# 0.002533f
C15505 trim_val\[2\] _447_/a_36_151# 0.022122f
C15506 _430_/a_36_151# _091_ 0.02228f
C15507 _098_ _201_/a_67_603# 0.005932f
C15508 _445_/a_2560_156# net47 0.014069f
C15509 FILLER_0_15_150/a_124_375# net56 0.011873f
C15510 net18 _418_/a_448_472# 0.026048f
C15511 _143_ FILLER_0_18_139/a_1380_472# 0.002226f
C15512 output8/a_224_472# FILLER_0_3_221/a_572_375# 0.03228f
C15513 FILLER_0_17_142/a_572_375# vss 0.049716f
C15514 FILLER_0_17_142/a_36_472# vdd 0.108843f
C15515 result[1] vdd 0.221634f
C15516 FILLER_0_5_172/a_124_375# _163_ 0.006403f
C15517 net18 _419_/a_2248_156# 0.014287f
C15518 net73 _098_ 0.004745f
C15519 _142_ FILLER_0_17_161/a_36_472# 0.00657f
C15520 _436_/a_1308_423# vdd 0.005258f
C15521 _143_ FILLER_0_16_154/a_1468_375# 0.002033f
C15522 FILLER_0_4_197/a_572_375# net59 0.001512f
C15523 _096_ net79 0.015605f
C15524 _440_/a_448_472# _029_ 0.043511f
C15525 _232_/a_255_603# _164_ 0.001274f
C15526 mask\[7\] _024_ 0.122185f
C15527 net55 FILLER_0_21_60/a_124_375# 0.015315f
C15528 _430_/a_1308_423# mask\[2\] 0.020226f
C15529 _363_/a_36_68# _163_ 0.005627f
C15530 FILLER_0_18_76/a_572_375# vdd -0.009037f
C15531 FILLER_0_18_76/a_124_375# vss 0.006877f
C15532 FILLER_0_16_73/a_36_472# _131_ 0.008223f
C15533 vdd _416_/a_2560_156# 0.00165f
C15534 vss _416_/a_2665_112# 0.002676f
C15535 _091_ _333_/a_36_160# 0.031262f
C15536 result[0] FILLER_0_9_282/a_484_472# 0.018647f
C15537 _367_/a_36_68# _153_ 0.019803f
C15538 _118_ _227_/a_36_160# 0.017547f
C15539 _429_/a_2248_156# vss 0.040729f
C15540 _429_/a_2665_112# vdd 0.010552f
C15541 trim_mask\[1\] FILLER_0_4_91/a_124_375# 0.006803f
C15542 _064_ net39 0.558387f
C15543 _086_ _314_/a_224_472# 0.003715f
C15544 net16 net66 0.030521f
C15545 FILLER_0_20_98/a_36_472# _437_/a_36_151# 0.001723f
C15546 FILLER_0_10_247/a_36_472# vss 0.002828f
C15547 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_36_472# 0.026657f
C15548 FILLER_0_8_263/a_36_472# net19 0.047387f
C15549 _414_/a_448_472# net22 0.047364f
C15550 _414_/a_1000_472# _081_ 0.006091f
C15551 _178_ _184_ 0.436202f
C15552 net31 vss 0.562041f
C15553 _013_ FILLER_0_21_28/a_1828_472# 0.003978f
C15554 _136_ FILLER_0_16_154/a_1468_375# 0.0028f
C15555 fanout52/a_36_160# _386_/a_124_24# 0.004695f
C15556 net20 state\[0\] 0.396139f
C15557 _292_/a_36_160# _105_ 0.027405f
C15558 net23 _207_/a_67_603# 0.002734f
C15559 net47 _450_/a_36_151# 0.029201f
C15560 _008_ _418_/a_36_151# 0.016984f
C15561 cal_count\[3\] _314_/a_224_472# 0.002143f
C15562 FILLER_0_19_125/a_36_472# _022_ 0.013011f
C15563 _432_/a_2665_112# vdd 0.009104f
C15564 _289_/a_36_472# _099_ 0.035055f
C15565 FILLER_0_12_136/a_572_375# FILLER_0_13_142/a_36_472# 0.001684f
C15566 net52 FILLER_0_6_47/a_3260_375# 0.040612f
C15567 mask\[4\] _143_ 0.352305f
C15568 net41 trim_val\[1\] 0.001912f
C15569 FILLER_0_12_220/a_124_375# _090_ 0.001521f
C15570 _424_/a_2560_156# vss 0.001554f
C15571 _024_ _435_/a_796_472# 0.006511f
C15572 mask\[4\] _348_/a_49_472# 0.001241f
C15573 ctlp[1] _421_/a_448_472# 0.011026f
C15574 net54 _437_/a_2560_156# 0.009745f
C15575 _098_ _023_ 0.004191f
C15576 _027_ _438_/a_796_472# 0.031292f
C15577 _150_ _438_/a_1204_472# 0.003696f
C15578 FILLER_0_21_28/a_124_375# FILLER_0_20_15/a_1468_375# 0.026339f
C15579 net67 trim_val\[0\] 0.382079f
C15580 _442_/a_1308_423# vdd 0.00782f
C15581 _442_/a_448_472# vss 0.001428f
C15582 result[7] _420_/a_448_472# 0.003274f
C15583 _446_/a_448_472# net17 0.026011f
C15584 FILLER_0_18_2/a_3172_472# vdd 0.011201f
C15585 _316_/a_124_24# _122_ 0.040082f
C15586 _316_/a_848_380# calibrate 0.012121f
C15587 _076_ _121_ 0.013717f
C15588 net15 _423_/a_1308_423# 0.001999f
C15589 _345_/a_36_160# FILLER_0_19_125/a_124_375# 0.005398f
C15590 FILLER_0_5_109/a_484_472# _160_ 0.001598f
C15591 _233_/a_36_160# _444_/a_36_151# 0.032942f
C15592 _445_/a_36_151# vss 0.009726f
C15593 _445_/a_448_472# vdd 0.007946f
C15594 _029_ vss 0.11129f
C15595 _414_/a_36_151# _087_ 0.010359f
C15596 _317_/a_36_113# _014_ 0.037134f
C15597 _016_ _118_ 0.001549f
C15598 _322_/a_848_380# _126_ 0.002519f
C15599 _029_ _365_/a_692_472# 0.001426f
C15600 FILLER_0_4_197/a_36_472# net76 0.003914f
C15601 _410_/a_36_68# vdd 0.039824f
C15602 net16 _067_ 0.039705f
C15603 net52 _168_ 0.726039f
C15604 _055_ _311_/a_66_473# 0.040326f
C15605 _086_ _321_/a_170_472# 0.046783f
C15606 _182_ _179_ 0.109377f
C15607 FILLER_0_16_37/a_124_375# _181_ 0.001198f
C15608 FILLER_0_8_138/a_36_472# _062_ 0.001109f
C15609 _077_ _453_/a_1308_423# 0.071515f
C15610 _068_ _227_/a_36_160# 0.053563f
C15611 net15 _424_/a_2248_156# 0.00415f
C15612 _131_ _124_ 0.002448f
C15613 _123_ vss 0.016878f
C15614 mask\[7\] _435_/a_1308_423# 0.028235f
C15615 input1/a_36_113# input4/a_36_68# 0.015796f
C15616 comp vss 0.148428f
C15617 _436_/a_36_151# ctlp[7] 0.002655f
C15618 net63 FILLER_0_19_187/a_36_472# 0.006753f
C15619 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_1020_375# 0.001597f
C15620 _126_ mask\[0\] 0.067513f
C15621 FILLER_0_12_20/a_484_472# _039_ 0.006288f
C15622 _178_ net47 0.09023f
C15623 _447_/a_2665_112# net15 0.063341f
C15624 net44 FILLER_0_20_2/a_484_472# 0.039736f
C15625 output47/a_224_472# net47 0.023797f
C15626 output21/a_224_472# _105_ 0.034631f
C15627 FILLER_0_21_142/a_572_375# FILLER_0_22_128/a_2276_472# 0.001543f
C15628 _144_ FILLER_0_21_125/a_572_375# 0.003787f
C15629 net26 _217_/a_36_160# 0.021067f
C15630 net34 _422_/a_36_151# 0.032272f
C15631 _303_/a_36_472# _110_ 0.001606f
C15632 FILLER_0_16_107/a_484_472# _131_ 0.008223f
C15633 _207_/a_67_603# net33 0.005153f
C15634 FILLER_0_20_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001543f
C15635 mask\[5\] _048_ 0.062788f
C15636 net53 FILLER_0_16_154/a_36_472# 0.006261f
C15637 FILLER_0_4_107/a_1468_375# _154_ 0.005202f
C15638 FILLER_0_4_107/a_572_375# _153_ 0.010165f
C15639 FILLER_0_21_286/a_124_375# _009_ 0.001024f
C15640 mask\[5\] FILLER_0_18_177/a_484_472# 0.001063f
C15641 net80 mask\[1\] 0.015535f
C15642 net20 FILLER_0_13_228/a_124_375# 0.047331f
C15643 net58 output37/a_224_472# 0.099539f
C15644 _255_/a_224_552# _116_ 0.027303f
C15645 _120_ vdd 0.750809f
C15646 _408_/a_728_93# _095_ 0.040366f
C15647 mask\[2\] FILLER_0_16_154/a_932_472# 0.021665f
C15648 _072_ _375_/a_1612_497# 0.002646f
C15649 FILLER_0_13_142/a_484_472# _043_ 0.011974f
C15650 net32 _421_/a_1000_472# 0.002275f
C15651 _432_/a_2248_156# FILLER_0_18_177/a_1828_472# 0.035805f
C15652 FILLER_0_18_107/a_572_375# FILLER_0_19_111/a_124_375# 0.058411f
C15653 _272_/a_36_472# _079_ 0.0237f
C15654 output37/a_224_472# _425_/a_2665_112# 0.022027f
C15655 _376_/a_36_160# FILLER_0_5_72/a_1380_472# 0.035111f
C15656 _081_ net47 1.302193f
C15657 net17 FILLER_0_20_15/a_484_472# 0.011079f
C15658 net58 net5 0.387314f
C15659 _186_ cal_count\[2\] 0.001605f
C15660 FILLER_0_15_150/a_124_375# _095_ 0.003939f
C15661 net41 FILLER_0_21_28/a_124_375# 0.003254f
C15662 cal fanout58/a_36_160# 0.047586f
C15663 _434_/a_36_151# mask\[6\] 0.048644f
C15664 FILLER_0_18_76/a_484_472# net71 0.004649f
C15665 net64 _100_ 0.001674f
C15666 FILLER_0_9_28/a_2276_472# vss -0.001894f
C15667 net81 _195_/a_67_603# 0.002322f
C15668 FILLER_0_17_104/a_36_472# _438_/a_2248_156# 0.001731f
C15669 net73 _131_ 0.022043f
C15670 ctlp[1] FILLER_0_24_274/a_484_472# 0.001875f
C15671 net65 _074_ 0.002666f
C15672 _100_ mask\[1\] 0.002229f
C15673 _101_ _005_ 0.003946f
C15674 trim_mask\[4\] _370_/a_1152_472# 0.001449f
C15675 _441_/a_2665_112# net14 0.00104f
C15676 net23 FILLER_0_22_128/a_3260_375# 0.012171f
C15677 net52 FILLER_0_2_111/a_1380_472# 0.050754f
C15678 _372_/a_3126_472# _068_ 0.005304f
C15679 _444_/a_1308_423# net40 0.043396f
C15680 _077_ _074_ 0.148596f
C15681 _043_ _113_ 0.048005f
C15682 net20 result[8] 0.014571f
C15683 FILLER_0_20_193/a_124_375# vdd 0.009092f
C15684 net75 net19 1.345314f
C15685 _326_/a_36_160# FILLER_0_7_104/a_1380_472# 0.002051f
C15686 output14/a_224_472# trim_mask\[3\] 0.001155f
C15687 net80 vss 0.347557f
C15688 output42/a_224_472# output6/a_224_472# 0.292612f
C15689 FILLER_0_17_72/a_1380_472# _131_ 0.006873f
C15690 _439_/a_2248_156# net14 0.001279f
C15691 net69 _031_ 0.450281f
C15692 FILLER_0_9_105/a_572_375# vdd 0.074717f
C15693 FILLER_0_4_185/a_36_472# vss 0.002627f
C15694 net50 net17 0.010654f
C15695 _425_/a_1000_472# net19 0.020388f
C15696 _115_ _076_ 0.051404f
C15697 _092_ mask\[3\] 0.040554f
C15698 FILLER_0_13_206/a_36_472# net79 0.00402f
C15699 FILLER_0_18_139/a_1468_375# vss 0.009191f
C15700 FILLER_0_18_139/a_36_472# vdd 0.089771f
C15701 _104_ net19 0.159483f
C15702 net65 FILLER_0_3_172/a_1020_375# 0.006035f
C15703 output44/a_224_472# net17 0.07836f
C15704 net15 _098_ 0.003965f
C15705 _105_ ctlp[2] 0.223601f
C15706 FILLER_0_16_154/a_124_375# vdd 0.00439f
C15707 FILLER_0_5_72/a_484_472# _440_/a_36_151# 0.001723f
C15708 result[7] FILLER_0_24_274/a_1380_472# 0.006454f
C15709 fanout62/a_36_160# net18 0.008106f
C15710 net19 _420_/a_36_151# 0.016882f
C15711 _094_ vdd 0.717159f
C15712 _100_ vss 0.020176f
C15713 _036_ FILLER_0_3_54/a_124_375# 0.010221f
C15714 _089_ _003_ 0.014763f
C15715 _370_/a_124_24# vss 0.005764f
C15716 _370_/a_848_380# vdd -0.001256f
C15717 mask\[7\] FILLER_0_22_128/a_484_472# 0.010605f
C15718 _126_ _124_ 0.012466f
C15719 net61 output19/a_224_472# 0.077658f
C15720 FILLER_0_8_127/a_124_375# _058_ 0.007791f
C15721 net54 _140_ 1.37516f
C15722 _305_/a_36_159# vss 0.003366f
C15723 net55 FILLER_0_21_28/a_2724_472# 0.049771f
C15724 _415_/a_36_151# net64 0.001735f
C15725 _320_/a_1120_472# state\[1\] 0.001998f
C15726 mask\[0\] _137_ 0.009052f
C15727 _259_/a_271_68# net4 0.003663f
C15728 _254_/a_448_472# _072_ 0.002611f
C15729 net16 _446_/a_2665_112# 0.045966f
C15730 ctln[2] vdd 0.245598f
C15731 net68 FILLER_0_6_47/a_1380_472# 0.049638f
C15732 _227_/a_36_160# vdd 0.007828f
C15733 net74 _370_/a_124_24# 0.083426f
C15734 FILLER_0_18_107/a_572_375# vdd 0.00419f
C15735 FILLER_0_18_107/a_124_375# vss 0.003425f
C15736 trim_mask\[1\] FILLER_0_6_47/a_2276_472# 0.006166f
C15737 net31 _103_ 0.227588f
C15738 _132_ _431_/a_448_472# 0.003024f
C15739 output28/a_224_472# FILLER_0_11_282/a_124_375# 0.002977f
C15740 net33 FILLER_0_22_128/a_3260_375# 0.001178f
C15741 net54 FILLER_0_22_128/a_124_375# 0.032013f
C15742 _052_ FILLER_0_18_37/a_932_472# 0.002749f
C15743 net76 FILLER_0_5_198/a_36_472# 0.003987f
C15744 FILLER_0_21_28/a_2276_472# _423_/a_36_151# 0.013806f
C15745 FILLER_0_5_117/a_124_375# _158_ 0.001068f
C15746 _421_/a_1308_423# net19 0.055838f
C15747 _030_ _367_/a_692_472# 0.002082f
C15748 _326_/a_36_160# _070_ 0.018037f
C15749 _152_ _059_ 0.038141f
C15750 cal_itt\[3\] FILLER_0_6_177/a_572_375# 0.00225f
C15751 net69 _371_/a_36_113# 0.016091f
C15752 _446_/a_2248_156# vdd 0.059236f
C15753 FILLER_0_9_28/a_1828_472# _042_ 0.001809f
C15754 FILLER_0_9_28/a_1380_472# net51 0.002012f
C15755 _187_ _039_ 0.228074f
C15756 _410_/a_36_68# cal_count\[0\] 0.007618f
C15757 _421_/a_2248_156# _419_/a_2248_156# 0.001364f
C15758 FILLER_0_19_55/a_36_472# _013_ 0.005889f
C15759 FILLER_0_11_282/a_36_472# _416_/a_1308_423# 0.001295f
C15760 FILLER_0_24_274/a_124_375# vss 0.002674f
C15761 _414_/a_36_151# vdd 0.166006f
C15762 FILLER_0_5_164/a_124_375# _386_/a_848_380# 0.014613f
C15763 FILLER_0_5_72/a_36_472# vss 0.031034f
C15764 FILLER_0_5_72/a_484_472# vdd 0.002735f
C15765 FILLER_0_12_136/a_1020_375# state\[2\] 0.001952f
C15766 net80 FILLER_0_18_177/a_1828_472# 0.00195f
C15767 _426_/a_36_151# net19 0.04851f
C15768 output19/a_224_472# _108_ 0.005075f
C15769 _155_ FILLER_0_4_91/a_572_375# 0.004038f
C15770 _308_/a_124_24# _439_/a_2248_156# 0.01963f
C15771 FILLER_0_8_107/a_36_472# _219_/a_36_160# 0.002767f
C15772 net20 net82 0.026007f
C15773 FILLER_0_5_164/a_36_472# _385_/a_36_68# 0.001674f
C15774 _118_ net21 0.007371f
C15775 net16 FILLER_0_8_24/a_572_375# 0.002225f
C15776 net38 net49 0.117427f
C15777 FILLER_0_7_72/a_1468_375# FILLER_0_5_72/a_1380_472# 0.00108f
C15778 net70 net53 1.170795f
C15779 _104_ _009_ 0.284256f
C15780 _016_ vdd 0.114288f
C15781 fanout61/a_36_113# _418_/a_36_151# 0.001442f
C15782 _415_/a_448_472# vdd 0.005273f
C15783 _415_/a_36_151# vss 0.003124f
C15784 _408_/a_56_524# vdd 0.003158f
C15785 _408_/a_728_93# vss 0.001345f
C15786 net16 net26 0.273031f
C15787 net63 FILLER_0_18_177/a_2724_472# 0.001857f
C15788 _115_ FILLER_0_11_78/a_484_472# 0.003641f
C15789 trimb[0] FILLER_0_20_2/a_124_375# 0.006864f
C15790 _096_ _335_/a_257_69# 0.001084f
C15791 _420_/a_36_151# _009_ 0.018171f
C15792 FILLER_0_15_142/a_36_472# net73 0.001893f
C15793 _221_/a_36_160# vss 0.037067f
C15794 net82 _163_ 0.00269f
C15795 mask\[5\] _108_ 0.036539f
C15796 _027_ mask\[9\] 0.050723f
C15797 _288_/a_224_472# _102_ 0.002528f
C15798 _176_ _451_/a_3129_107# 0.021559f
C15799 ctln[7] _442_/a_2665_112# 0.01075f
C15800 _093_ FILLER_0_17_142/a_36_472# 0.011974f
C15801 FILLER_0_15_150/a_36_472# vdd 0.088307f
C15802 FILLER_0_15_150/a_124_375# vss 0.01957f
C15803 FILLER_0_4_107/a_932_472# _158_ 0.029116f
C15804 output46/a_224_472# trimb[3] 0.050924f
C15805 FILLER_0_8_24/a_124_375# vdd 0.01166f
C15806 FILLER_0_5_54/a_932_472# _440_/a_36_151# 0.001723f
C15807 _372_/a_2590_472# vss 0.00106f
C15808 FILLER_0_11_142/a_36_472# _120_ 0.040786f
C15809 FILLER_0_15_116/a_484_472# _095_ 0.001069f
C15810 _120_ cal_count\[0\] 0.014209f
C15811 net54 _149_ 0.212511f
C15812 net32 ctlp[1] 0.032275f
C15813 net50 _441_/a_448_472# 0.074088f
C15814 _028_ FILLER_0_7_72/a_3172_472# 0.001873f
C15815 _086_ net57 0.126563f
C15816 FILLER_0_13_212/a_572_375# net79 0.009626f
C15817 ctln[6] vdd 0.116327f
C15818 FILLER_0_5_128/a_484_472# _370_/a_124_24# 0.00171f
C15819 net23 _433_/a_2248_156# 0.005588f
C15820 _078_ FILLER_0_6_231/a_36_472# 0.013046f
C15821 FILLER_0_20_177/a_1468_375# mask\[6\] 0.001162f
C15822 net72 FILLER_0_18_37/a_124_375# 0.05632f
C15823 net18 _006_ 0.082256f
C15824 FILLER_0_4_107/a_124_375# _160_ 0.005906f
C15825 _093_ FILLER_0_18_76/a_572_375# 0.025143f
C15826 _131_ _427_/a_36_151# 0.0012f
C15827 net52 _440_/a_2665_112# 0.005084f
C15828 FILLER_0_23_274/a_124_375# vss 0.017196f
C15829 FILLER_0_23_274/a_36_472# vdd 0.010289f
C15830 fanout62/a_36_160# net62 0.02201f
C15831 output14/a_224_472# FILLER_0_0_130/a_36_472# 0.023414f
C15832 net57 cal_count\[3\] 0.02848f
C15833 net50 _439_/a_36_151# 0.009774f
C15834 net52 _439_/a_1308_423# 0.033366f
C15835 output44/a_224_472# FILLER_0_18_2/a_1468_375# 0.032639f
C15836 _086_ _135_ 0.005637f
C15837 net81 _138_ 0.006815f
C15838 _053_ FILLER_0_7_72/a_1380_472# 0.01339f
C15839 _425_/a_448_472# net37 0.002755f
C15840 FILLER_0_16_37/a_124_375# FILLER_0_18_37/a_36_472# 0.001512f
C15841 mask\[4\] FILLER_0_18_177/a_36_472# 0.018019f
C15842 ctln[1] rstn 0.62944f
C15843 net55 FILLER_0_19_28/a_484_472# 0.001426f
C15844 output36/a_224_472# _417_/a_2248_156# 0.023576f
C15845 _033_ FILLER_0_6_47/a_124_375# 0.002521f
C15846 _321_/a_786_69# net23 0.001073f
C15847 _434_/a_1308_423# vdd 0.033494f
C15848 _432_/a_2665_112# _093_ 0.02266f
C15849 FILLER_0_8_107/a_124_375# FILLER_0_10_107/a_36_472# 0.0027f
C15850 _274_/a_3368_68# vss 0.001714f
C15851 _096_ FILLER_0_14_181/a_36_472# 0.028078f
C15852 _068_ net21 0.030836f
C15853 cal_count\[3\] _135_ 0.039115f
C15854 FILLER_0_12_136/a_124_375# vdd 0.004378f
C15855 _068_ _261_/a_36_160# 0.008557f
C15856 _070_ _059_ 0.041498f
C15857 _131_ _180_ 0.016104f
C15858 _131_ net15 0.037758f
C15859 _031_ FILLER_0_2_111/a_572_375# 0.023633f
C15860 net69 FILLER_0_2_111/a_1468_375# 0.021524f
C15861 _239_/a_36_160# _064_ 0.001292f
C15862 _065_ trim_mask\[2\] 0.002792f
C15863 _053_ net76 0.022571f
C15864 ctln[4] FILLER_0_0_198/a_124_375# 0.015879f
C15865 ctln[2] net2 0.004284f
C15866 net75 cal_itt\[0\] 0.032053f
C15867 _065_ _447_/a_1308_423# 0.024822f
C15868 _414_/a_36_151# _057_ 0.003902f
C15869 _028_ _058_ 0.041158f
C15870 _128_ _121_ 0.051501f
C15871 result[5] result[7] 0.016166f
C15872 net20 _098_ 0.087341f
C15873 output23/a_224_472# mask\[7\] 0.046766f
C15874 FILLER_0_5_54/a_484_472# vss 0.001929f
C15875 FILLER_0_5_54/a_932_472# vdd 0.003166f
C15876 cal_count\[2\] _452_/a_448_472# 0.003314f
C15877 FILLER_0_18_107/a_1468_375# net71 0.001292f
C15878 _242_/a_36_160# vss 0.032884f
C15879 ctlp[5] mask\[7\] 0.131468f
C15880 FILLER_0_17_133/a_36_472# _137_ 0.001963f
C15881 mask\[0\] _060_ 0.002039f
C15882 _428_/a_2665_112# _427_/a_36_151# 0.028591f
C15883 _441_/a_1308_423# _164_ 0.001807f
C15884 FILLER_0_10_28/a_36_472# output6/a_224_472# 0.010475f
C15885 _182_ _041_ 0.08834f
C15886 _193_/a_36_160# output30/a_224_472# 0.018f
C15887 net57 _169_ 0.033365f
C15888 _096_ _320_/a_1120_472# 0.004315f
C15889 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_36_472# 0.026657f
C15890 FILLER_0_14_91/a_36_472# _136_ 0.008573f
C15891 _233_/a_36_160# net49 0.035342f
C15892 FILLER_0_11_142/a_572_375# _121_ 0.003107f
C15893 _421_/a_1000_472# _010_ 0.01379f
C15894 _181_ _182_ 0.02735f
C15895 net20 FILLER_0_13_212/a_1380_472# 0.006746f
C15896 ctln[1] FILLER_0_1_266/a_484_472# 0.002068f
C15897 _440_/a_2248_156# _164_ 0.054298f
C15898 _258_/a_36_160# vdd 0.00617f
C15899 _151_ vdd 0.157764f
C15900 _322_/a_692_472# _118_ 0.002849f
C15901 output34/a_224_472# vdd 0.094191f
C15902 net16 FILLER_0_17_38/a_36_472# 0.014381f
C15903 _308_/a_848_380# _058_ 0.031449f
C15904 trimb[1] vdd 0.225206f
C15905 trim_mask\[3\] _157_ 0.052956f
C15906 net73 _137_ 0.047989f
C15907 _253_/a_1528_68# cal_itt\[1\] 0.002251f
C15908 FILLER_0_7_72/a_1828_472# net52 0.00159f
C15909 FILLER_0_7_72/a_932_472# net50 0.074005f
C15910 net81 FILLER_0_15_212/a_1468_375# 0.006906f
C15911 vss _022_ 0.067509f
C15912 FILLER_0_2_177/a_572_375# net59 0.005397f
C15913 result[1] _416_/a_2248_156# 0.001888f
C15914 FILLER_0_17_226/a_36_472# mask\[3\] 0.011509f
C15915 _017_ FILLER_0_14_107/a_1020_375# 0.001363f
C15916 net70 FILLER_0_14_107/a_36_472# 0.054561f
C15917 FILLER_0_9_28/a_1020_375# net50 0.001512f
C15918 net27 _426_/a_2560_156# 0.004199f
C15919 _110_ _423_/a_2665_112# 0.001668f
C15920 net20 net63 0.045207f
C15921 _053_ FILLER_0_7_59/a_572_375# 0.014569f
C15922 _431_/a_2560_156# net36 0.001858f
C15923 net15 FILLER_0_5_54/a_1468_375# 0.039975f
C15924 FILLER_0_24_290/a_124_375# FILLER_0_24_274/a_1468_375# 0.012001f
C15925 FILLER_0_20_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001543f
C15926 _341_/a_49_472# FILLER_0_16_154/a_572_375# 0.001643f
C15927 FILLER_0_4_177/a_124_375# net76 0.003962f
C15928 net44 net40 0.003336f
C15929 _449_/a_1308_423# _453_/a_2665_112# 0.001066f
C15930 FILLER_0_16_57/a_932_472# _131_ 0.007885f
C15931 net78 _094_ 0.050187f
C15932 net60 _094_ 0.579872f
C15933 _412_/a_448_472# en 0.011052f
C15934 FILLER_0_17_38/a_572_375# vdd 0.01525f
C15935 FILLER_0_5_109/a_36_472# net47 0.005565f
C15936 net67 FILLER_0_6_47/a_1828_472# 0.001175f
C15937 net46 FILLER_0_20_15/a_572_375# 0.029486f
C15938 _321_/a_170_472# _120_ 0.040613f
C15939 _053_ net14 0.713784f
C15940 _345_/a_36_160# vdd 0.100094f
C15941 cal_itt\[1\] _082_ 0.921465f
C15942 net3 FILLER_0_15_2/a_572_375# 0.004377f
C15943 _098_ _433_/a_796_472# 0.002825f
C15944 FILLER_0_3_2/a_36_472# vss 0.004076f
C15945 net67 _039_ 0.302826f
C15946 _006_ net62 0.136418f
C15947 _308_/a_1084_68# net14 0.002892f
C15948 _043_ vdd 0.827689f
C15949 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3172_472# 0.026657f
C15950 FILLER_0_13_65/a_124_375# _043_ 0.013045f
C15951 net34 FILLER_0_22_177/a_484_472# 0.003953f
C15952 net44 input3/a_36_113# 0.016865f
C15953 _307_/a_234_472# _113_ 0.007518f
C15954 ctlp[1] _419_/a_2560_156# 0.002551f
C15955 mask\[9\] _438_/a_796_472# 0.004751f
C15956 _130_ _427_/a_36_151# 0.001056f
C15957 _236_/a_36_160# output39/a_224_472# 0.042231f
C15958 _395_/a_36_488# _116_ 0.033784f
C15959 _412_/a_2665_112# vss 0.011887f
C15960 _079_ _074_ 0.025058f
C15961 FILLER_0_19_125/a_36_472# net73 0.004017f
C15962 FILLER_0_3_172/a_1916_375# net22 0.00941f
C15963 ctlp[8] vdd 0.115254f
C15964 FILLER_0_18_171/a_124_375# mask\[3\] 0.001156f
C15965 net76 net18 0.002264f
C15966 _064_ _160_ 0.006705f
C15967 _185_ vdd 0.325358f
C15968 _429_/a_36_151# _018_ 0.118135f
C15969 cal_itt\[3\] _374_/a_36_68# 0.001569f
C15970 FILLER_0_18_37/a_1380_472# vss 0.002042f
C15971 _081_ _385_/a_36_68# 0.006303f
C15972 FILLER_0_15_142/a_36_472# _427_/a_36_151# 0.001723f
C15973 cal_itt\[2\] _082_ 0.032565f
C15974 FILLER_0_21_133/a_124_375# vdd 0.010519f
C15975 _073_ net82 0.028504f
C15976 mask\[7\] _107_ 0.13732f
C15977 FILLER_0_14_91/a_484_472# net53 0.00544f
C15978 FILLER_0_15_228/a_36_472# net62 0.002128f
C15979 FILLER_0_15_116/a_484_472# vss 0.003923f
C15980 net53 state\[1\] 0.00554f
C15981 _175_ vdd 0.147794f
C15982 net7 _447_/a_36_151# 0.002494f
C15983 FILLER_0_1_98/a_124_375# _065_ 0.001136f
C15984 cal_count\[3\] _408_/a_1336_472# 0.010351f
C15985 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_124_375# 0.003732f
C15986 _413_/a_36_151# FILLER_0_3_172/a_2276_472# 0.001723f
C15987 _116_ _228_/a_36_68# 0.013091f
C15988 _086_ _129_ 0.051553f
C15989 net63 output22/a_224_472# 0.017997f
C15990 mask\[0\] _095_ 0.006711f
C15991 net50 FILLER_0_7_59/a_124_375# 0.002292f
C15992 _411_/a_2248_156# _073_ 0.003809f
C15993 _412_/a_1308_423# net76 0.023786f
C15994 FILLER_0_11_101/a_572_375# _134_ 0.0024f
C15995 _062_ _113_ 0.020368f
C15996 _265_/a_244_68# cal_itt\[1\] 0.024108f
C15997 net79 _099_ 0.010543f
C15998 _155_ _363_/a_36_68# 0.013915f
C15999 _115_ _128_ 0.263909f
C16000 net21 vdd 1.653552f
C16001 result[7] net19 0.087363f
C16002 _261_/a_36_160# vdd 0.0109f
C16003 _436_/a_2248_156# _025_ 0.001054f
C16004 _441_/a_2665_112# net49 0.062459f
C16005 _129_ cal_count\[3\] 0.005967f
C16006 _053_ _359_/a_1044_488# 0.001474f
C16007 _036_ net40 0.599505f
C16008 _093_ FILLER_0_18_139/a_36_472# 0.008761f
C16009 FILLER_0_10_107/a_36_472# vss 0.003894f
C16010 FILLER_0_10_107/a_484_472# vdd 0.034172f
C16011 trim_val\[3\] _441_/a_1308_423# 0.001312f
C16012 trim_mask\[2\] _036_ 0.466145f
C16013 _085_ _055_ 0.240451f
C16014 _375_/a_960_497# vdd 0.004471f
C16015 net24 FILLER_0_22_107/a_124_375# 0.001023f
C16016 net71 _437_/a_36_151# 0.055761f
C16017 FILLER_0_12_136/a_36_472# _127_ 0.023927f
C16018 _064_ _445_/a_1000_472# 0.015908f
C16019 _447_/a_1000_472# net68 0.006223f
C16020 _447_/a_1308_423# _036_ 0.003079f
C16021 _116_ calibrate 0.018482f
C16022 net18 _007_ 0.060872f
C16023 FILLER_0_20_177/a_36_472# vss 0.003944f
C16024 FILLER_0_20_177/a_484_472# vdd 0.010805f
C16025 _093_ _094_ 0.003586f
C16026 _091_ FILLER_0_15_212/a_932_472# 0.008749f
C16027 _335_/a_49_472# FILLER_0_15_180/a_572_375# 0.001126f
C16028 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_36_472# 0.002296f
C16029 net80 _019_ 0.265857f
C16030 FILLER_0_14_263/a_124_375# vdd 0.026205f
C16031 calibrate FILLER_0_9_270/a_36_472# 0.00119f
C16032 fanout75/a_36_113# net76 0.040306f
C16033 valid fanout64/a_36_160# 0.001811f
C16034 _118_ _062_ 0.029651f
C16035 FILLER_0_8_2/a_124_375# _054_ 0.001055f
C16036 net70 FILLER_0_16_115/a_36_472# 0.003407f
C16037 FILLER_0_2_111/a_1380_472# FILLER_0_2_127/a_36_472# 0.013276f
C16038 FILLER_0_10_78/a_1020_375# net52 0.001158f
C16039 _057_ _043_ 0.02152f
C16040 FILLER_0_4_144/a_36_472# vss 0.008308f
C16041 FILLER_0_4_144/a_484_472# vdd 0.004027f
C16042 _070_ _247_/a_36_160# 0.0169f
C16043 FILLER_0_18_177/a_124_375# vdd 0.033102f
C16044 output37/a_224_472# sample 0.015298f
C16045 _077_ net15 0.238832f
C16046 _105_ ctlp[1] 0.158795f
C16047 FILLER_0_4_107/a_124_375# _156_ 0.00268f
C16048 net82 _425_/a_36_151# 0.002959f
C16049 _093_ FILLER_0_18_107/a_572_375# 0.008393f
C16050 mask\[5\] _049_ 0.008296f
C16051 _081_ FILLER_0_6_177/a_572_375# 0.007285f
C16052 _411_/a_36_151# _000_ 0.023297f
C16053 _411_/a_1308_423# net75 0.028281f
C16054 _419_/a_1000_472# vdd 0.004107f
C16055 net41 _444_/a_448_472# 0.031876f
C16056 _053_ FILLER_0_6_90/a_572_375# 0.073688f
C16057 sample net5 0.359975f
C16058 net52 FILLER_0_9_72/a_932_472# 0.008749f
C16059 net23 _208_/a_36_160# 0.112626f
C16060 net61 output18/a_224_472# 0.059062f
C16061 FILLER_0_20_2/a_124_375# net43 0.001563f
C16062 _028_ net52 0.150861f
C16063 _106_ FILLER_0_17_218/a_572_375# 0.022684f
C16064 FILLER_0_4_144/a_572_375# FILLER_0_5_148/a_124_375# 0.05841f
C16065 FILLER_0_21_133/a_36_472# _140_ 0.008378f
C16066 _453_/a_1308_423# vss 0.003012f
C16067 _178_ net72 0.007093f
C16068 net48 _014_ 0.276733f
C16069 _095_ _451_/a_36_151# 0.008311f
C16070 _003_ FILLER_0_5_181/a_36_472# 0.003545f
C16071 FILLER_0_16_241/a_36_472# net36 0.001988f
C16072 ctln[1] cal_itt\[2\] 0.053339f
C16073 FILLER_0_15_212/a_572_375# mask\[1\] 0.012463f
C16074 FILLER_0_19_171/a_932_472# vss 0.001256f
C16075 FILLER_0_19_171/a_1380_472# vdd 0.03086f
C16076 _348_/a_49_472# _146_ 0.001552f
C16077 ctlp[1] _010_ 0.002794f
C16078 net82 net1 0.029512f
C16079 FILLER_0_14_181/a_36_472# FILLER_0_15_180/a_124_375# 0.001723f
C16080 _031_ vss 0.18315f
C16081 _425_/a_448_472# _122_ 0.002863f
C16082 _425_/a_1308_423# calibrate 0.022697f
C16083 mask\[0\] net64 0.45093f
C16084 net58 en 0.029072f
C16085 result[7] _009_ 0.697145f
C16086 _035_ net17 0.021052f
C16087 net45 net40 0.029947f
C16088 _438_/a_1000_472# vss 0.001536f
C16089 FILLER_0_16_57/a_1468_375# _175_ 0.001654f
C16090 mask\[0\] mask\[1\] 0.01742f
C16091 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_484_472# 0.013276f
C16092 _011_ _422_/a_796_472# 0.009261f
C16093 _132_ _334_/a_36_160# 0.026495f
C16094 _057_ net21 0.143214f
C16095 net79 FILLER_0_21_286/a_572_375# 0.001476f
C16096 cal_count\[2\] _179_ 0.404284f
C16097 trim_mask\[4\] _159_ 0.049552f
C16098 FILLER_0_15_282/a_572_375# _006_ 0.001054f
C16099 net38 net47 0.352245f
C16100 net28 _094_ 0.007842f
C16101 net15 FILLER_0_15_59/a_36_472# 0.00464f
C16102 _180_ FILLER_0_15_59/a_36_472# 0.087308f
C16103 net16 _402_/a_728_93# 0.040925f
C16104 net73 FILLER_0_18_107/a_2276_472# 0.016723f
C16105 net15 _453_/a_36_151# 0.009841f
C16106 FILLER_0_16_89/a_1380_472# net14 0.049391f
C16107 _255_/a_224_552# _375_/a_36_68# 0.00229f
C16108 _068_ _062_ 0.089152f
C16109 _070_ _134_ 0.087767f
C16110 _137_ FILLER_0_19_155/a_124_375# 0.00129f
C16111 net48 _070_ 0.264809f
C16112 _077_ net51 0.76967f
C16113 _432_/a_2248_156# net80 0.059406f
C16114 net47 _386_/a_692_472# 0.003299f
C16115 _322_/a_848_380# vss 0.026127f
C16116 _321_/a_2590_472# _129_ 0.005391f
C16117 _161_ state\[1\] 0.002512f
C16118 output26/a_224_472# FILLER_0_23_44/a_1380_472# 0.0323f
C16119 result[8] FILLER_0_24_274/a_1020_375# 0.00726f
C16120 net15 net69 0.034091f
C16121 FILLER_0_1_98/a_36_472# _442_/a_2665_112# 0.002597f
C16122 _210_/a_67_603# net23 0.005398f
C16123 net50 FILLER_0_6_90/a_124_375# 0.041764f
C16124 _395_/a_1492_488# _121_ 0.002537f
C16125 FILLER_0_6_47/a_1916_375# vdd -0.014642f
C16126 FILLER_0_6_47/a_1468_375# vss 0.003462f
C16127 _043_ cal_count\[0\] 0.019077f
C16128 FILLER_0_19_55/a_124_375# FILLER_0_17_56/a_36_472# 0.001338f
C16129 FILLER_0_15_212/a_572_375# vss 0.005835f
C16130 FILLER_0_15_212/a_1020_375# vdd -0.00211f
C16131 _052_ mask\[9\] 0.007224f
C16132 _449_/a_36_151# FILLER_0_13_72/a_36_472# 0.001723f
C16133 _402_/a_1296_93# vdd 0.017239f
C16134 FILLER_0_17_200/a_572_375# _069_ 0.011239f
C16135 _322_/a_848_380# net74 0.00168f
C16136 vdd _450_/a_2449_156# 0.003646f
C16137 net23 FILLER_0_16_154/a_36_472# 0.035678f
C16138 ctlp[6] _050_ 0.100418f
C16139 mask\[0\] vss 0.694674f
C16140 _185_ cal_count\[0\] 0.008096f
C16141 _082_ net59 0.004251f
C16142 _074_ vss 0.404343f
C16143 FILLER_0_8_247/a_572_375# calibrate 0.008498f
C16144 fanout50/a_36_160# net52 0.037383f
C16145 _301_/a_36_472# _051_ 0.001277f
C16146 net35 _213_/a_255_603# 0.001597f
C16147 _419_/a_36_151# net77 0.163616f
C16148 _204_/a_67_603# vss 0.010366f
C16149 net4 _082_ 0.004529f
C16150 _293_/a_36_472# vdd 0.087136f
C16151 net73 _095_ 0.003688f
C16152 _132_ net36 0.029615f
C16153 _057_ _267_/a_1568_472# 0.002083f
C16154 net52 _443_/a_36_151# 0.020518f
C16155 _303_/a_36_472# _012_ 0.001735f
C16156 en_co_clk _390_/a_36_68# 0.086301f
C16157 input2/a_36_113# rstn 0.002202f
C16158 _430_/a_36_151# fanout80/a_36_113# 0.018169f
C16159 net57 _120_ 0.012391f
C16160 _431_/a_2665_112# FILLER_0_16_154/a_36_472# 0.007491f
C16161 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1468_375# 0.086635f
C16162 _055_ _310_/a_49_472# 0.00384f
C16163 net18 FILLER_0_11_282/a_36_472# 0.048657f
C16164 net67 clkc 0.102244f
C16165 _077_ FILLER_0_9_72/a_1020_375# 0.008103f
C16166 FILLER_0_9_28/a_1828_472# _120_ 0.00108f
C16167 FILLER_0_17_72/a_3172_472# _136_ 0.002925f
C16168 _453_/a_448_472# _042_ 0.053209f
C16169 _453_/a_36_151# net51 0.012537f
C16170 fanout68/a_36_113# net66 0.042828f
C16171 FILLER_0_6_239/a_36_472# vss 0.003177f
C16172 fanout75/a_36_113# _083_ 0.002133f
C16173 _086_ FILLER_0_10_107/a_572_375# 0.001179f
C16174 net54 _098_ 0.116416f
C16175 fanout69/a_36_113# _159_ 0.005623f
C16176 net74 _371_/a_36_113# 0.027966f
C16177 FILLER_0_18_53/a_124_375# vdd 0.022f
C16178 FILLER_0_16_73/a_36_472# vss 0.035175f
C16179 FILLER_0_16_73/a_484_472# vdd 0.003462f
C16180 _075_ _078_ 0.001896f
C16181 _433_/a_448_472# _022_ 0.074451f
C16182 _135_ _120_ 0.017522f
C16183 net81 FILLER_0_15_228/a_124_375# 0.006974f
C16184 FILLER_0_3_172/a_1468_375# vdd 0.045181f
C16185 ctln[5] _448_/a_2248_156# 0.004396f
C16186 result[0] vdd 0.193436f
C16187 _422_/a_2248_156# vss 0.001755f
C16188 _422_/a_2665_112# vdd 0.008306f
C16189 trim_val\[3\] net14 0.01035f
C16190 _033_ vdd 0.509957f
C16191 net20 net65 0.335083f
C16192 _415_/a_2665_112# _416_/a_36_151# 0.001602f
C16193 fanout60/a_36_160# FILLER_0_17_282/a_36_472# 0.002647f
C16194 _431_/a_36_151# FILLER_0_18_107/a_1828_472# 0.001221f
C16195 _413_/a_36_151# net82 0.00601f
C16196 _265_/a_244_68# net59 0.001147f
C16197 _064_ net67 0.006691f
C16198 net55 FILLER_0_17_72/a_572_375# 0.023585f
C16199 output34/a_224_472# _093_ 0.012298f
C16200 _446_/a_796_472# net66 0.002296f
C16201 _345_/a_36_160# _433_/a_36_151# 0.015565f
C16202 _233_/a_36_160# net47 0.054273f
C16203 net4 FILLER_0_8_239/a_36_472# 0.008503f
C16204 _187_ _174_ 0.001321f
C16205 ctlp[4] output22/a_224_472# 0.008275f
C16206 net73 FILLER_0_19_111/a_572_375# 0.04458f
C16207 output8/a_224_472# net82 0.002936f
C16208 _112_ _316_/a_1084_68# 0.005773f
C16209 _307_/a_234_472# vdd 0.001209f
C16210 net20 _077_ 0.094476f
C16211 net56 FILLER_0_19_155/a_124_375# 0.006762f
C16212 _112_ net59 0.002846f
C16213 _092_ output18/a_224_472# 0.002205f
C16214 FILLER_0_3_221/a_484_472# vss 0.005602f
C16215 FILLER_0_3_221/a_932_472# vdd 0.005654f
C16216 net54 FILLER_0_18_139/a_572_375# 0.00217f
C16217 net65 _163_ 0.013462f
C16218 _142_ FILLER_0_18_107/a_2724_472# 0.001549f
C16219 FILLER_0_16_73/a_124_375# net15 0.005202f
C16220 FILLER_0_20_193/a_572_375# _098_ 0.078973f
C16221 _451_/a_36_151# vss 0.028073f
C16222 _451_/a_448_472# vdd 0.04463f
C16223 ctln[1] _411_/a_448_472# 0.039538f
C16224 FILLER_0_5_72/a_36_472# _029_ 0.007282f
C16225 FILLER_0_5_72/a_572_375# trim_mask\[1\] 0.010714f
C16226 FILLER_0_3_172/a_2724_472# net21 0.009426f
C16227 _086_ _267_/a_672_472# 0.004515f
C16228 mask\[9\] FILLER_0_19_111/a_36_472# 0.285112f
C16229 _001_ vdd 0.122898f
C16230 FILLER_0_20_98/a_36_472# net14 0.024154f
C16231 _189_/a_67_603# FILLER_0_12_220/a_1468_375# 0.029786f
C16232 _321_/a_3126_472# _126_ 0.002939f
C16233 _321_/a_358_69# _069_ 0.001124f
C16234 _059_ FILLER_0_8_156/a_36_472# 0.18373f
C16235 _431_/a_796_472# _136_ 0.009889f
C16236 _104_ _106_ 0.17237f
C16237 net16 net17 0.034209f
C16238 FILLER_0_21_133/a_124_375# _433_/a_36_151# 0.059049f
C16239 FILLER_0_13_228/a_36_472# _043_ 0.02119f
C16240 ctln[1] net59 0.053978f
C16241 _126_ FILLER_0_12_196/a_124_375# 0.001392f
C16242 FILLER_0_2_111/a_36_472# vdd 0.033758f
C16243 FILLER_0_2_111/a_1468_375# vss 0.055168f
C16244 net35 mask\[6\] 0.041818f
C16245 fanout56/a_36_113# _136_ 0.002316f
C16246 _317_/a_36_113# calibrate 0.011799f
C16247 _077_ _256_/a_1612_497# 0.002724f
C16248 cal_count\[3\] _453_/a_448_472# 0.001494f
C16249 _142_ FILLER_0_17_133/a_124_375# 0.022066f
C16250 net45 net46 0.038161f
C16251 _062_ vdd 0.393862f
C16252 _431_/a_36_151# fanout70/a_36_113# 0.016241f
C16253 output48/a_224_472# vdd 0.038342f
C16254 output44/a_224_472# FILLER_0_19_28/a_36_472# 0.023414f
C16255 _098_ FILLER_0_16_154/a_572_375# 0.001791f
C16256 ctln[1] net4 0.009703f
C16257 _414_/a_2248_156# net59 0.004437f
C16258 net41 FILLER_0_20_31/a_36_472# 0.030033f
C16259 net55 net47 0.049398f
C16260 _449_/a_36_151# FILLER_0_11_64/a_36_472# 0.046516f
C16261 FILLER_0_5_128/a_124_375# _159_ 0.003644f
C16262 _124_ vss 0.110847f
C16263 net61 _418_/a_448_472# 0.001253f
C16264 FILLER_0_18_107/a_3172_472# vss 0.006614f
C16265 FILLER_0_7_72/a_3172_472# FILLER_0_7_104/a_36_472# 0.013276f
C16266 state\[1\] _071_ 0.196063f
C16267 net20 _419_/a_448_472# 0.025583f
C16268 _132_ _020_ 0.037636f
C16269 ctln[6] _442_/a_36_151# 0.007031f
C16270 net78 _419_/a_1000_472# 0.040603f
C16271 net60 _419_/a_1000_472# 0.028992f
C16272 net61 _419_/a_2248_156# 0.022159f
C16273 _110_ _437_/a_36_151# 0.00125f
C16274 net63 FILLER_0_20_193/a_572_375# 0.015818f
C16275 net74 FILLER_0_2_111/a_1468_375# 0.003854f
C16276 _096_ _161_ 0.00104f
C16277 _417_/a_2560_156# _006_ 0.007804f
C16278 _053_ net68 0.239882f
C16279 output43/a_224_472# trimb[3] 0.070044f
C16280 trimb[0] output46/a_224_472# 0.048191f
C16281 trimb[4] _452_/a_3129_107# 0.004943f
C16282 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_36_472# 0.026657f
C16283 FILLER_0_21_28/a_1828_472# _012_ 0.021162f
C16284 output31/a_224_472# _417_/a_448_472# 0.008149f
C16285 net74 _124_ 0.180235f
C16286 _069_ net36 0.032818f
C16287 FILLER_0_16_107/a_484_472# vss 0.004223f
C16288 _178_ _407_/a_36_472# 0.001699f
C16289 FILLER_0_11_282/a_36_472# net62 0.00149f
C16290 FILLER_0_16_57/a_124_375# FILLER_0_18_53/a_484_472# 0.001512f
C16291 _076_ _226_/a_1044_68# 0.0023f
C16292 FILLER_0_17_133/a_36_472# vss 0.006791f
C16293 output25/a_224_472# net25 0.179738f
C16294 net29 net36 0.370099f
C16295 net50 _160_ 0.048787f
C16296 _308_/a_692_472# trim_mask\[0\] 0.004377f
C16297 _093_ net21 0.032584f
C16298 FILLER_0_15_142/a_124_375# net36 0.006533f
C16299 vss _201_/a_67_603# 0.012925f
C16300 FILLER_0_16_89/a_36_472# _397_/a_36_472# 0.004546f
C16301 output21/a_224_472# _107_ 0.086601f
C16302 net38 FILLER_0_20_2/a_36_472# 0.002204f
C16303 net72 FILLER_0_12_50/a_124_375# 0.011077f
C16304 net23 net47 0.090948f
C16305 _004_ vdd 0.448886f
C16306 FILLER_0_11_101/a_36_472# net14 0.04522f
C16307 net4 FILLER_0_12_220/a_484_472# 0.022264f
C16308 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_124_375# 0.012222f
C16309 _119_ _074_ 0.153267f
C16310 net73 vss 0.342554f
C16311 _423_/a_36_151# FILLER_0_23_44/a_1020_375# 0.059049f
C16312 FILLER_0_7_104/a_36_472# _058_ 0.006613f
C16313 _257_/a_36_472# cal_itt\[3\] 0.136487f
C16314 net16 FILLER_0_16_37/a_36_472# 0.015199f
C16315 _016_ net57 0.028276f
C16316 _427_/a_36_151# _095_ 0.029048f
C16317 net75 FILLER_0_0_232/a_124_375# 0.00217f
C16318 _430_/a_2665_112# mask\[3\] 0.002697f
C16319 net68 FILLER_0_5_54/a_124_375# 0.018458f
C16320 fanout72/a_36_113# net72 0.02315f
C16321 net19 cal_itt\[1\] 0.044717f
C16322 _129_ _120_ 0.017802f
C16323 FILLER_0_5_212/a_124_375# net37 0.005414f
C16324 FILLER_0_5_54/a_1020_375# trim_mask\[1\] 0.010745f
C16325 net50 _030_ 0.073046f
C16326 net41 _034_ 0.026084f
C16327 FILLER_0_21_142/a_124_375# vdd 0.020936f
C16328 _441_/a_36_151# _440_/a_36_151# 0.003983f
C16329 mask\[0\] FILLER_0_12_236/a_36_472# 0.002801f
C16330 net35 FILLER_0_22_86/a_1380_472# 0.00813f
C16331 _091_ FILLER_0_15_180/a_124_375# 0.001415f
C16332 net73 net74 0.016949f
C16333 net52 _442_/a_2665_112# 0.031179f
C16334 _140_ _350_/a_49_472# 0.028997f
C16335 _021_ mask\[4\] 0.018108f
C16336 _256_/a_2552_68# _072_ 0.001213f
C16337 net17 _452_/a_1353_112# 0.038603f
C16338 _162_ FILLER_0_6_177/a_36_472# 0.001723f
C16339 _161_ FILLER_0_6_177/a_572_375# 0.004064f
C16340 FILLER_0_17_72/a_1828_472# vdd 0.001969f
C16341 FILLER_0_17_72/a_1380_472# vss 0.003698f
C16342 output7/a_224_472# net41 0.003942f
C16343 net20 _420_/a_2665_112# 0.030202f
C16344 _027_ FILLER_0_18_76/a_572_375# 0.08501f
C16345 _150_ FILLER_0_18_76/a_484_472# 0.003548f
C16346 FILLER_0_7_195/a_36_472# vdd 0.04565f
C16347 FILLER_0_7_195/a_124_375# vss 0.006314f
C16348 FILLER_0_21_206/a_124_375# _204_/a_67_603# 0.003591f
C16349 _068_ FILLER_0_5_148/a_36_472# 0.003015f
C16350 _057_ _062_ 0.062063f
C16351 FILLER_0_16_37/a_124_375# vdd 0.038329f
C16352 valid net19 0.00646f
C16353 output35/a_224_472# FILLER_0_22_177/a_1468_375# 0.018187f
C16354 net18 FILLER_0_9_270/a_484_472# 0.004375f
C16355 _069_ _116_ 0.390834f
C16356 net2 _001_ 0.081616f
C16357 _095_ _180_ 0.013383f
C16358 FILLER_0_8_127/a_124_375# _070_ 0.003265f
C16359 net15 _095_ 0.056214f
C16360 net58 cal 0.001209f
C16361 _063_ _232_/a_67_603# 0.005404f
C16362 result[9] _006_ 0.05748f
C16363 FILLER_0_19_111/a_484_472# vss 0.003811f
C16364 _013_ FILLER_0_18_53/a_36_472# 0.013138f
C16365 net16 _235_/a_67_603# 0.038585f
C16366 FILLER_0_7_59/a_36_472# trim_val\[0\] 0.003014f
C16367 _023_ vss 0.114191f
C16368 FILLER_0_24_130/a_36_472# ctlp[7] 0.012298f
C16369 FILLER_0_19_187/a_36_472# vss 0.001951f
C16370 FILLER_0_19_187/a_484_472# vdd 0.011023f
C16371 FILLER_0_0_198/a_36_472# net11 0.056269f
C16372 _011_ vdd 0.182751f
C16373 output16/a_224_472# _447_/a_448_472# 0.003175f
C16374 FILLER_0_1_192/a_124_375# vdd 0.017212f
C16375 output26/a_224_472# ctlp[9] 0.034572f
C16376 FILLER_0_4_213/a_572_375# net59 0.061684f
C16377 _140_ FILLER_0_21_150/a_124_375# 0.019084f
C16378 output48/a_224_472# net2 0.06309f
C16379 net14 FILLER_0_10_94/a_484_472# 0.020589f
C16380 _173_ _186_ 0.002111f
C16381 net27 FILLER_0_12_236/a_484_472# 0.042937f
C16382 FILLER_0_1_266/a_124_375# FILLER_0_0_266/a_124_375# 0.05841f
C16383 _015_ FILLER_0_8_247/a_1020_375# 0.006994f
C16384 net4 FILLER_0_4_213/a_572_375# 0.001015f
C16385 FILLER_0_12_136/a_124_375# net57 0.001727f
C16386 net65 _073_ 0.775972f
C16387 FILLER_0_17_72/a_484_472# net15 0.002925f
C16388 net41 _445_/a_2248_156# 0.065247f
C16389 output35/a_224_472# _205_/a_36_160# 0.002043f
C16390 _276_/a_36_160# _291_/a_36_160# 0.239422f
C16391 cal_count\[2\] _041_ 0.02197f
C16392 cal_itt\[3\] _251_/a_1130_472# 0.001099f
C16393 _399_/a_224_472# net72 0.002538f
C16394 _098_ _434_/a_796_472# 0.001383f
C16395 _441_/a_36_151# vdd 0.098562f
C16396 _088_ _260_/a_36_68# 0.003476f
C16397 net49 _164_ 0.428468f
C16398 net53 _427_/a_1204_472# 0.004293f
C16399 _444_/a_2248_156# net67 0.028782f
C16400 net16 FILLER_0_19_47/a_36_472# 0.009509f
C16401 _077_ _073_ 0.009611f
C16402 _394_/a_56_524# FILLER_0_15_59/a_572_375# 0.003413f
C16403 _181_ cal_count\[2\] 0.375819f
C16404 _139_ _138_ 0.00256f
C16405 output38/a_224_472# net38 0.018882f
C16406 net68 _164_ 0.189377f
C16407 net20 _426_/a_2665_112# 0.018602f
C16408 FILLER_0_16_255/a_36_472# vss 0.00184f
C16409 _431_/a_36_151# vdd 0.145005f
C16410 output10/a_224_472# ctln[3] 0.064347f
C16411 _440_/a_796_472# vss 0.001285f
C16412 net35 _352_/a_49_472# 0.02594f
C16413 mask\[8\] _352_/a_257_69# 0.003259f
C16414 FILLER_0_9_28/a_36_472# net47 0.006712f
C16415 fanout62/a_36_160# FILLER_0_13_290/a_124_375# 0.001138f
C16416 _044_ vdd 0.406979f
C16417 net80 _434_/a_448_472# 0.113898f
C16418 FILLER_0_16_89/a_484_472# _176_ 0.004026f
C16419 _091_ FILLER_0_13_212/a_572_375# 0.022882f
C16420 net20 _060_ 0.0426f
C16421 net58 FILLER_0_8_263/a_36_472# 0.059769f
C16422 _017_ _332_/a_36_472# 0.033837f
C16423 net34 _435_/a_2248_156# 0.01519f
C16424 trim_mask\[2\] FILLER_0_2_93/a_124_375# 0.046032f
C16425 net20 FILLER_0_3_221/a_1468_375# 0.007234f
C16426 net36 FILLER_0_15_235/a_36_472# 0.00664f
C16427 _114_ _121_ 0.002513f
C16428 FILLER_0_21_142/a_572_375# _140_ 0.018708f
C16429 _277_/a_36_160# vdd 0.115507f
C16430 FILLER_0_7_104/a_124_375# _131_ 0.001291f
C16431 FILLER_0_19_47/a_572_375# vdd 0.019566f
C16432 FILLER_0_19_47/a_124_375# vss 0.002211f
C16433 trim_val\[4\] net47 0.003977f
C16434 net36 _438_/a_36_151# 0.076525f
C16435 FILLER_0_17_200/a_572_375# net22 0.047331f
C16436 _024_ FILLER_0_22_177/a_36_472# 0.003242f
C16437 net32 net33 0.467071f
C16438 ctlp[3] _296_/a_224_472# 0.005335f
C16439 _316_/a_124_24# vdd 0.033047f
C16440 _132_ FILLER_0_18_107/a_1916_375# 0.019011f
C16441 _053_ FILLER_0_7_104/a_1468_375# 0.001492f
C16442 _091_ _337_/a_49_472# 0.014992f
C16443 _444_/a_2665_112# _054_ 0.003576f
C16444 _069_ _117_ 0.041311f
C16445 mask\[5\] FILLER_0_20_177/a_572_375# 0.013294f
C16446 FILLER_0_17_142/a_484_472# _137_ 0.003953f
C16447 FILLER_0_24_96/a_124_375# net25 0.008342f
C16448 input4/a_36_68# vdd 0.09828f
C16449 FILLER_0_17_72/a_2812_375# net14 0.018463f
C16450 _009_ _298_/a_224_472# 0.002441f
C16451 net15 _440_/a_448_472# 0.036624f
C16452 _423_/a_2665_112# _012_ 0.014394f
C16453 _430_/a_2248_156# net36 0.001198f
C16454 output7/a_224_472# net7 0.01565f
C16455 _412_/a_1204_472# net1 0.019647f
C16456 _293_/a_36_472# _093_ 0.004121f
C16457 _152_ FILLER_0_5_136/a_36_472# 0.049485f
C16458 FILLER_0_9_28/a_1020_375# net16 0.012909f
C16459 FILLER_0_21_286/a_484_472# _420_/a_36_151# 0.027236f
C16460 _238_/a_67_603# vss 0.008203f
C16461 FILLER_0_21_206/a_36_472# mask\[6\] 0.015735f
C16462 FILLER_0_22_86/a_1468_375# net14 0.024975f
C16463 net79 FILLER_0_12_220/a_484_472# 0.005464f
C16464 net57 _043_ 1.955053f
C16465 _448_/a_796_472# net59 0.004855f
C16466 _053_ _414_/a_1000_472# 0.029433f
C16467 _143_ _141_ 0.192528f
C16468 mask\[7\] FILLER_0_22_177/a_1468_375# 0.001315f
C16469 FILLER_0_0_96/a_36_472# vss 0.00344f
C16470 calibrate _059_ 0.506928f
C16471 _427_/a_36_151# vss 0.019281f
C16472 output37/a_224_472# calibrate 0.013149f
C16473 _141_ _348_/a_49_472# 0.037821f
C16474 FILLER_0_7_72/a_36_472# vss 0.033878f
C16475 ctln[9] net15 0.01475f
C16476 _016_ _129_ 0.002216f
C16477 _297_/a_36_472# _108_ 0.011437f
C16478 net20 _079_ 0.177911f
C16479 _326_/a_36_160# _125_ 0.050008f
C16480 mask\[8\] net15 0.02403f
C16481 state\[1\] net23 0.075055f
C16482 vdd FILLER_0_5_148/a_36_472# 0.001227f
C16483 vss FILLER_0_5_148/a_572_375# 0.042687f
C16484 _412_/a_36_151# _082_ 0.016538f
C16485 FILLER_0_9_28/a_572_375# vdd 0.023246f
C16486 _430_/a_36_151# FILLER_0_18_209/a_36_472# 0.002841f
C16487 FILLER_0_12_124/a_36_472# _332_/a_36_472# 0.004546f
C16488 net65 net1 0.035488f
C16489 sample en 0.001572f
C16490 _375_/a_36_68# calibrate 0.048799f
C16491 mask\[5\] FILLER_0_19_171/a_1468_375# 0.007169f
C16492 _077_ _067_ 0.090648f
C16493 _002_ FILLER_0_3_172/a_1828_472# 0.016749f
C16494 fanout81/a_36_160# fanout76/a_36_160# 0.01081f
C16495 _443_/a_36_151# _152_ 0.002345f
C16496 _427_/a_36_151# net74 0.04306f
C16497 FILLER_0_19_55/a_36_472# _012_ 0.001667f
C16498 _437_/a_2665_112# net14 0.002936f
C16499 fanout58/a_36_160# cal_itt\[1\] 0.010654f
C16500 net44 _450_/a_36_151# 0.026203f
C16501 _328_/a_36_113# _070_ 0.016264f
C16502 cal_itt\[1\] cal_itt\[0\] 0.055355f
C16503 _076_ _078_ 0.012626f
C16504 _359_/a_1044_488# _133_ 0.001894f
C16505 _359_/a_1492_488# _070_ 0.0043f
C16506 _359_/a_36_488# _076_ 0.005184f
C16507 _432_/a_36_151# _333_/a_36_160# 0.032942f
C16508 FILLER_0_22_177/a_572_375# net33 0.013337f
C16509 FILLER_0_21_133/a_36_472# _098_ 0.002964f
C16510 _106_ mask\[2\] 0.039965f
C16511 _180_ vss 0.106022f
C16512 FILLER_0_6_177/a_484_472# FILLER_0_5_181/a_36_472# 0.05841f
C16513 net15 vss 1.330044f
C16514 FILLER_0_17_38/a_484_472# _041_ 0.009607f
C16515 FILLER_0_13_65/a_36_472# net15 0.036527f
C16516 net50 _156_ 0.020099f
C16517 _444_/a_1204_472# net47 0.007847f
C16518 fanout51/a_36_113# vss 0.0844f
C16519 _113_ FILLER_0_12_196/a_36_472# 0.002495f
C16520 FILLER_0_22_177/a_932_472# _435_/a_36_151# 0.001723f
C16521 net69 net66 0.09789f
C16522 _120_ FILLER_0_10_107/a_572_375# 0.002214f
C16523 FILLER_0_19_155/a_572_375# vdd 0.01384f
C16524 FILLER_0_19_155/a_124_375# vss 0.00336f
C16525 FILLER_0_20_107/a_36_472# _438_/a_2665_112# 0.035266f
C16526 _442_/a_448_472# _031_ 0.019293f
C16527 trim_val\[3\] net49 0.009336f
C16528 _131_ FILLER_0_11_124/a_124_375# 0.008946f
C16529 result[0] FILLER_0_9_290/a_124_375# 0.030628f
C16530 _443_/a_36_151# FILLER_0_2_127/a_36_472# 0.006095f
C16531 FILLER_0_15_205/a_36_472# net21 0.007503f
C16532 ctln[5] FILLER_0_0_198/a_36_472# 0.012298f
C16533 _308_/a_848_380# _070_ 0.033275f
C16534 _115_ _131_ 0.410424f
C16535 net14 FILLER_0_4_91/a_124_375# 0.009573f
C16536 net50 net67 0.518421f
C16537 mask\[7\] net19 0.003605f
C16538 _053_ FILLER_0_8_37/a_36_472# 0.001011f
C16539 net15 net74 0.05717f
C16540 output46/a_224_472# net43 0.10562f
C16541 net19 net59 0.0206f
C16542 net34 FILLER_0_22_128/a_2276_472# 0.005532f
C16543 _452_/a_3129_107# vss 0.00145f
C16544 _452_/a_2225_156# vdd 0.005612f
C16545 FILLER_0_9_28/a_3172_472# _077_ 0.011059f
C16546 _432_/a_2560_156# vdd 0.003219f
C16547 FILLER_0_3_54/a_36_472# net40 0.069702f
C16548 cal_itt\[2\] cal_itt\[0\] 0.011453f
C16549 _016_ _428_/a_2560_156# 0.003934f
C16550 _005_ _099_ 0.001603f
C16551 trim_mask\[2\] FILLER_0_3_54/a_36_472# 0.004063f
C16552 net4 net19 0.050898f
C16553 _412_/a_36_151# _265_/a_244_68# 0.072351f
C16554 _119_ _312_/a_672_472# 0.00145f
C16555 _039_ output6/a_224_472# 0.012051f
C16556 net56 FILLER_0_17_142/a_484_472# 0.008895f
C16557 _114_ _115_ 0.148291f
C16558 FILLER_0_16_107/a_124_375# _040_ 0.008721f
C16559 mask\[0\] _429_/a_2248_156# 0.016246f
C16560 FILLER_0_4_107/a_932_472# FILLER_0_2_111/a_572_375# 0.001512f
C16561 _070_ FILLER_0_5_136/a_36_472# 0.029293f
C16562 _255_/a_224_552# _311_/a_66_473# 0.002588f
C16563 cal_count\[1\] _180_ 0.300952f
C16564 net15 cal_count\[1\] 0.089855f
C16565 FILLER_0_18_177/a_3172_472# vdd 0.002358f
C16566 FILLER_0_20_177/a_932_472# _098_ 0.008366f
C16567 _412_/a_448_472# fanout81/a_36_160# 0.00998f
C16568 net35 FILLER_0_22_128/a_1468_375# 0.015932f
C16569 output30/a_224_472# net30 0.043557f
C16570 FILLER_0_5_212/a_124_375# _122_ 0.001352f
C16571 net77 vdd 0.526632f
C16572 net75 net58 0.061787f
C16573 mask\[4\] _069_ 0.001182f
C16574 _114_ FILLER_0_12_136/a_572_375# 0.006974f
C16575 net2 input4/a_36_68# 0.031809f
C16576 FILLER_0_4_144/a_484_472# net57 0.003724f
C16577 _077_ FILLER_0_9_105/a_36_472# 0.003177f
C16578 net27 result[1] 0.187252f
C16579 output26/a_224_472# _423_/a_36_151# 0.011936f
C16580 output47/a_224_472# net44 0.077292f
C16581 _256_/a_36_68# _068_ 0.029112f
C16582 result[5] net79 0.036275f
C16583 FILLER_0_16_241/a_124_375# _282_/a_36_160# 0.005398f
C16584 FILLER_0_9_105/a_124_375# FILLER_0_10_107/a_36_472# 0.001543f
C16585 FILLER_0_11_101/a_124_375# _171_ 0.00105f
C16586 net51 vss 0.21065f
C16587 net36 net22 0.034258f
C16588 trim_mask\[3\] _156_ 0.002638f
C16589 FILLER_0_16_57/a_932_472# vss 0.003388f
C16590 FILLER_0_16_57/a_1380_472# vdd 0.005673f
C16591 trim_mask\[1\] FILLER_0_6_47/a_124_375# 0.005902f
C16592 net60 _011_ 0.003094f
C16593 _011_ net78 0.002956f
C16594 FILLER_0_20_193/a_124_375# FILLER_0_20_177/a_1468_375# 0.012222f
C16595 _053_ net47 0.011652f
C16596 _303_/a_36_472# vdd 0.015964f
C16597 net50 FILLER_0_8_24/a_484_472# 0.059367f
C16598 _102_ vdd 0.211559f
C16599 _056_ state\[1\] 0.219625f
C16600 _104_ net30 0.001375f
C16601 FILLER_0_22_128/a_1916_375# vss 0.018094f
C16602 FILLER_0_22_128/a_2364_375# vdd 0.015888f
C16603 net81 net36 0.030215f
C16604 _415_/a_1204_472# net18 0.001828f
C16605 _414_/a_2248_156# cal_itt\[3\] 0.032294f
C16606 FILLER_0_9_28/a_2724_472# _453_/a_448_472# 0.008036f
C16607 result[5] _290_/a_224_472# 0.001638f
C16608 FILLER_0_2_93/a_484_472# net14 0.019214f
C16609 fanout79/a_36_160# vdd 0.099877f
C16610 net63 FILLER_0_20_177/a_932_472# 0.004375f
C16611 _073_ FILLER_0_3_221/a_1468_375# 0.006377f
C16612 net65 _413_/a_36_151# 0.033028f
C16613 trim[0] output40/a_224_472# 0.005306f
C16614 FILLER_0_19_47/a_484_472# _013_ 0.009677f
C16615 vdd output41/a_224_472# 0.003282f
C16616 mask\[7\] _009_ 0.078131f
C16617 _408_/a_1336_472# _043_ 0.023648f
C16618 net20 net64 0.374636f
C16619 _428_/a_1308_423# _017_ 0.005962f
C16620 _428_/a_448_472# net53 0.001959f
C16621 _116_ _090_ 0.122467f
C16622 FILLER_0_21_28/a_1916_375# _424_/a_36_151# 0.059049f
C16623 FILLER_0_4_123/a_36_472# vdd 0.091386f
C16624 FILLER_0_4_123/a_124_375# vss 0.009712f
C16625 FILLER_0_16_57/a_932_472# cal_count\[1\] 0.002217f
C16626 net20 mask\[1\] 0.09671f
C16627 output8/a_224_472# net65 0.084944f
C16628 _074_ _123_ 0.157299f
C16629 _098_ _438_/a_2248_156# 0.002798f
C16630 net63 FILLER_0_18_177/a_572_375# 0.004407f
C16631 _247_/a_36_160# _228_/a_36_68# 0.001919f
C16632 FILLER_0_2_111/a_484_472# _158_ 0.003604f
C16633 FILLER_0_5_54/a_124_375# net47 0.012889f
C16634 output9/a_224_472# net5 0.005189f
C16635 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_124_375# 0.003732f
C16636 FILLER_0_9_72/a_1020_375# vss 0.005622f
C16637 FILLER_0_9_72/a_1468_375# vdd 0.026475f
C16638 net82 FILLER_0_3_172/a_1916_375# 0.010202f
C16639 _397_/a_36_472# FILLER_0_17_72/a_1468_375# 0.001295f
C16640 FILLER_0_4_123/a_124_375# net74 0.002449f
C16641 FILLER_0_15_150/a_36_472# FILLER_0_15_142/a_484_472# 0.013277f
C16642 net58 FILLER_0_8_247/a_1468_375# 0.001669f
C16643 net75 FILLER_0_8_247/a_932_472# 0.006746f
C16644 net55 FILLER_0_13_72/a_124_375# 0.00281f
C16645 _093_ FILLER_0_17_72/a_1828_472# 0.053526f
C16646 _126_ FILLER_0_11_124/a_124_375# 0.038971f
C16647 _185_ _405_/a_255_603# 0.002565f
C16648 _182_ vdd 0.161134f
C16649 _130_ FILLER_0_11_124/a_124_375# 0.001943f
C16650 mask\[4\] FILLER_0_18_209/a_484_472# 0.021522f
C16651 _120_ _450_/a_3129_107# 0.001598f
C16652 _267_/a_224_472# _121_ 0.0029f
C16653 _394_/a_728_93# _095_ 0.035417f
C16654 _198_/a_67_603# vdd 0.015843f
C16655 _137_ FILLER_0_16_154/a_572_375# 0.010132f
C16656 _028_ FILLER_0_7_72/a_1020_375# 0.003837f
C16657 _116_ net22 0.122052f
C16658 _173_ FILLER_0_12_28/a_36_472# 0.001633f
C16659 ctln[6] _037_ 0.031407f
C16660 _193_/a_36_160# _416_/a_36_151# 0.065269f
C16661 _188_ vdd 0.022839f
C16662 FILLER_0_6_239/a_36_472# _123_ 0.004433f
C16663 net18 _417_/a_796_472# 0.006722f
C16664 net58 _426_/a_36_151# 0.002612f
C16665 net75 _426_/a_796_472# 0.003146f
C16666 FILLER_0_17_200/a_36_472# _432_/a_2665_112# 0.007491f
C16667 _105_ net33 0.202272f
C16668 FILLER_0_16_89/a_1468_375# _136_ 0.005791f
C16669 net82 FILLER_0_3_221/a_1380_472# 0.008049f
C16670 _003_ cal_itt\[3\] 0.054183f
C16671 result[6] _420_/a_1204_472# 0.002681f
C16672 _046_ _282_/a_36_160# 0.005584f
C16673 FILLER_0_15_282/a_124_375# output30/a_224_472# 0.029138f
C16674 _098_ FILLER_0_15_212/a_1468_375# 0.008327f
C16675 fanout67/a_36_160# vdd 0.018829f
C16676 FILLER_0_12_136/a_572_375# _126_ 0.01289f
C16677 _291_/a_36_160# vss 0.012222f
C16678 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_124_375# 0.007947f
C16679 _153_ vdd 0.672318f
C16680 _079_ _073_ 0.234533f
C16681 net39 FILLER_0_8_2/a_36_472# 0.010296f
C16682 FILLER_0_14_50/a_124_375# _180_ 0.022435f
C16683 net56 net54 0.018493f
C16684 _091_ FILLER_0_17_218/a_36_472# 0.066133f
C16685 _154_ _365_/a_36_68# 0.02267f
C16686 net81 FILLER_0_9_270/a_36_472# 0.084422f
C16687 _104_ _422_/a_36_151# 0.032235f
C16688 net15 FILLER_0_9_72/a_124_375# 0.006492f
C16689 net20 vss 1.402494f
C16690 mask\[3\] vdd 0.340612f
C16691 _035_ _160_ 0.120469f
C16692 _176_ FILLER_0_10_94/a_572_375# 0.011743f
C16693 _140_ FILLER_0_22_128/a_2812_375# 0.003154f
C16694 _283_/a_36_472# vdd 0.092097f
C16695 _132_ FILLER_0_14_107/a_124_375# 0.003315f
C16696 ctlp[1] FILLER_0_21_286/a_572_375# 0.026009f
C16697 _423_/a_36_151# FILLER_0_23_60/a_124_375# 0.005577f
C16698 FILLER_0_8_138/a_124_375# _059_ 0.007966f
C16699 _428_/a_2560_156# _043_ 0.009909f
C16700 _004_ net28 0.082388f
C16701 net25 FILLER_0_22_86/a_36_472# 0.001265f
C16702 _396_/a_224_472# _177_ 0.001254f
C16703 _050_ vdd 0.484554f
C16704 FILLER_0_21_28/a_1380_472# vss 0.001688f
C16705 FILLER_0_21_28/a_1828_472# vdd 0.004227f
C16706 net79 net19 0.03862f
C16707 _360_/a_36_160# net47 0.011731f
C16708 _163_ vss 0.638066f
C16709 net72 net55 0.233515f
C16710 FILLER_0_16_89/a_1020_375# FILLER_0_17_72/a_2812_375# 0.026339f
C16711 FILLER_0_16_89/a_36_472# FILLER_0_17_72/a_1916_375# 0.001723f
C16712 net71 net14 0.147175f
C16713 mask\[4\] FILLER_0_19_171/a_1020_375# 0.006236f
C16714 _117_ _090_ 0.041465f
C16715 _431_/a_36_151# _093_ 0.004862f
C16716 result[6] _421_/a_2665_112# 0.034452f
C16717 fanout58/a_36_160# net59 0.048057f
C16718 _004_ _416_/a_2248_156# 0.001078f
C16719 net47 _164_ 0.118311f
C16720 net58 fanout81/a_36_160# 0.013959f
C16721 _256_/a_1612_497# vss 0.004265f
C16722 _077_ _115_ 0.131611f
C16723 FILLER_0_18_2/a_1828_472# net17 0.008573f
C16724 FILLER_0_2_101/a_124_375# _157_ 0.002818f
C16725 net41 FILLER_0_23_44/a_36_472# 0.001116f
C16726 _004_ FILLER_0_10_247/a_124_375# 0.004573f
C16727 net31 _201_/a_67_603# 0.015773f
C16728 _115_ FILLER_0_10_107/a_124_375# 0.011098f
C16729 net74 _163_ 0.042013f
C16730 net4 cal_itt\[0\] 0.054266f
C16731 FILLER_0_5_117/a_124_375# vss 0.001764f
C16732 FILLER_0_5_117/a_36_472# vdd 0.092171f
C16733 net81 _425_/a_1308_423# 0.004202f
C16734 net32 net18 0.028135f
C16735 FILLER_0_17_56/a_124_375# FILLER_0_18_53/a_484_472# 0.001597f
C16736 _076_ _160_ 0.006506f
C16737 _101_ net62 0.023932f
C16738 _094_ _196_/a_36_160# 0.001668f
C16739 FILLER_0_4_49/a_484_472# vss 0.002751f
C16740 _277_/a_36_160# _093_ 0.018101f
C16741 net3 net17 0.045911f
C16742 _177_ _150_ 0.002507f
C16743 _136_ _018_ 0.002892f
C16744 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_572_375# 0.086635f
C16745 mask\[9\] FILLER_0_18_76/a_572_375# 0.006158f
C16746 net48 calibrate 0.482314f
C16747 output43/a_224_472# trimb[0] 0.043402f
C16748 net76 FILLER_0_3_172/a_1828_472# 0.051851f
C16749 _096_ _056_ 0.001946f
C16750 _065_ output16/a_224_472# 0.049052f
C16751 _239_/a_36_160# net16 0.003137f
C16752 _426_/a_36_151# FILLER_0_8_247/a_932_472# 0.001723f
C16753 mask\[0\] _100_ 0.005921f
C16754 _040_ vdd 0.065702f
C16755 ctln[1] _000_ 0.223573f
C16756 fanout49/a_36_160# trim_mask\[1\] 0.00358f
C16757 result[6] fanout61/a_36_113# 0.003917f
C16758 _116_ _076_ 0.008283f
C16759 _085_ _070_ 0.058787f
C16760 FILLER_0_17_72/a_484_472# FILLER_0_18_76/a_36_472# 0.05841f
C16761 net56 FILLER_0_18_139/a_484_472# 0.004375f
C16762 output36/a_224_472# net18 0.010751f
C16763 net75 _014_ 0.204357f
C16764 _428_/a_36_151# FILLER_0_14_107/a_484_472# 0.059367f
C16765 net76 net37 0.549565f
C16766 FILLER_0_20_177/a_484_472# _434_/a_36_151# 0.001723f
C16767 FILLER_0_16_89/a_36_472# net53 0.004701f
C16768 net56 FILLER_0_16_154/a_572_375# 0.002321f
C16769 _074_ _305_/a_36_159# 0.012602f
C16770 FILLER_0_1_98/a_124_375# ctln[7] 0.004533f
C16771 _371_/a_36_113# _370_/a_124_24# 0.008354f
C16772 _245_/a_672_472# net17 0.00121f
C16773 cal_count\[3\] _042_ 0.001716f
C16774 net55 _424_/a_36_151# 0.007344f
C16775 net39 _063_ 0.004732f
C16776 mask\[3\] FILLER_0_18_177/a_1380_472# 0.005654f
C16777 _285_/a_36_472# _099_ 0.040922f
C16778 _321_/a_3662_472# vdd 0.001229f
C16779 _251_/a_906_472# _070_ 0.002124f
C16780 FILLER_0_7_233/a_36_472# FILLER_0_6_231/a_124_375# 0.001684f
C16781 output6/a_224_472# clkc 0.017846f
C16782 FILLER_0_4_107/a_1380_472# vdd 0.007022f
C16783 _415_/a_2248_156# net58 0.001869f
C16784 FILLER_0_12_20/a_572_375# vss 0.054934f
C16785 FILLER_0_12_20/a_36_472# vdd 0.068477f
C16786 net24 FILLER_0_23_88/a_36_472# 0.006289f
C16787 FILLER_0_2_171/a_36_472# net59 0.066486f
C16788 _081_ _082_ 0.008298f
C16789 net67 _450_/a_1040_527# 0.032098f
C16790 net60 net77 0.046792f
C16791 net78 net77 0.252376f
C16792 _292_/a_36_160# _205_/a_36_160# 0.105676f
C16793 FILLER_0_18_2/a_2812_375# net55 0.007169f
C16794 vdd FILLER_0_12_196/a_36_472# 0.019648f
C16795 vss FILLER_0_12_196/a_124_375# 0.042104f
C16796 _413_/a_36_151# output12/a_224_472# 0.006251f
C16797 _367_/a_36_68# net14 0.055776f
C16798 net57 _062_ 0.067654f
C16799 _079_ net1 0.099822f
C16800 FILLER_0_24_130/a_124_375# net54 0.001269f
C16801 net18 FILLER_0_17_282/a_124_375# 0.048177f
C16802 output31/a_224_472# _006_ 0.090006f
C16803 net60 _102_ 0.008212f
C16804 net20 _260_/a_244_472# 0.001593f
C16805 FILLER_0_13_80/a_36_472# _451_/a_3129_107# 0.001115f
C16806 net40 net6 0.00772f
C16807 net28 _044_ 0.481924f
C16808 _158_ _157_ 0.001663f
C16809 _176_ net53 0.083005f
C16810 FILLER_0_14_81/a_124_375# _394_/a_728_93# 0.004587f
C16811 _095_ _067_ 0.00784f
C16812 _363_/a_244_472# _028_ 0.002693f
C16813 FILLER_0_5_128/a_484_472# _163_ 0.009861f
C16814 FILLER_0_19_171/a_1380_472# _434_/a_36_151# 0.00271f
C16815 _322_/a_692_472# _129_ 0.004891f
C16816 FILLER_0_9_223/a_124_375# _055_ 0.014525f
C16817 _394_/a_56_524# vdd 0.010692f
C16818 _394_/a_728_93# vss 0.024106f
C16819 _408_/a_728_93# _450_/a_2225_156# 0.00128f
C16820 fanout55/a_36_160# FILLER_0_13_80/a_124_375# 0.00805f
C16821 _069_ _059_ 0.002034f
C16822 _142_ FILLER_0_17_142/a_36_472# 0.011216f
C16823 FILLER_0_2_165/a_36_472# net59 0.067972f
C16824 net38 _444_/a_1308_423# 0.007915f
C16825 FILLER_0_14_50/a_36_472# cal_count\[3\] 0.005814f
C16826 _024_ net23 0.001994f
C16827 fanout78/a_36_113# net79 0.029496f
C16828 fanout60/a_36_160# net79 0.069956f
C16829 _044_ _416_/a_2248_156# 0.005198f
C16830 FILLER_0_14_99/a_124_375# _095_ 0.012128f
C16831 FILLER_0_19_28/a_572_375# vdd 0.034691f
C16832 FILLER_0_18_177/a_3260_375# _202_/a_36_160# 0.001948f
C16833 FILLER_0_4_91/a_572_375# _160_ 0.007391f
C16834 _050_ FILLER_0_22_128/a_572_375# 0.002607f
C16835 _086_ cal_count\[3\] 0.259095f
C16836 _449_/a_2665_112# _067_ 0.03661f
C16837 output38/a_224_472# _446_/a_36_151# 0.117966f
C16838 _098_ FILLER_0_21_150/a_124_375# 0.006526f
C16839 FILLER_0_15_2/a_36_472# vdd 0.104741f
C16840 FILLER_0_15_2/a_572_375# vss 0.055203f
C16841 FILLER_0_9_223/a_572_375# net4 0.02077f
C16842 net31 FILLER_0_16_255/a_36_472# 0.003056f
C16843 _081_ _265_/a_244_68# 0.03338f
C16844 FILLER_0_12_2/a_36_472# vss 0.003757f
C16845 _012_ FILLER_0_23_44/a_572_375# 0.002827f
C16846 trim_val\[2\] net40 0.06019f
C16847 _436_/a_1308_423# net35 0.008773f
C16848 _125_ _134_ 0.00437f
C16849 FILLER_0_16_89/a_124_375# vdd 0.01011f
C16850 net64 FILLER_0_9_270/a_124_375# 0.013532f
C16851 trim_mask\[2\] trim_val\[2\] 0.21814f
C16852 _417_/a_1000_472# net30 0.004556f
C16853 net16 _160_ 0.354736f
C16854 cal_itt\[3\] _162_ 0.141474f
C16855 _086_ _154_ 0.102849f
C16856 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_572_375# 0.086635f
C16857 _432_/a_2560_156# _093_ 0.007613f
C16858 _064_ _447_/a_36_151# 0.004185f
C16859 _430_/a_1308_423# _091_ 0.023198f
C16860 _112_ _081_ 0.037903f
C16861 _176_ FILLER_0_11_78/a_124_375# 0.004803f
C16862 _438_/a_448_472# _437_/a_36_151# 0.00198f
C16863 _451_/a_1697_156# net14 0.001298f
C16864 net66 _440_/a_448_472# 0.023934f
C16865 mask\[8\] _423_/a_2248_156# 0.001648f
C16866 net18 _418_/a_796_472# 0.003044f
C16867 output8/a_224_472# FILLER_0_3_221/a_1468_375# 0.032044f
C16868 _394_/a_728_93# cal_count\[1\] 0.057049f
C16869 FILLER_0_17_142/a_484_472# vss 0.030872f
C16870 fanout66/a_36_113# _164_ 0.010496f
C16871 net18 _419_/a_2560_156# 0.008155f
C16872 result[2] FILLER_0_14_263/a_36_472# 0.001134f
C16873 _436_/a_1000_472# vdd 0.006522f
C16874 output32/a_224_472# _419_/a_448_472# 0.010723f
C16875 mask\[2\] net30 0.089173f
C16876 _415_/a_448_472# net27 0.05785f
C16877 output19/a_224_472# vdd 0.063651f
C16878 net50 trim_val\[1\] 0.002079f
C16879 FILLER_0_4_197/a_1468_375# net59 0.050218f
C16880 ctlp[1] _420_/a_448_472# 0.038053f
C16881 _093_ FILLER_0_18_177/a_3172_472# 0.003708f
C16882 _440_/a_796_472# _029_ 0.009261f
C16883 output36/a_224_472# net62 0.317201f
C16884 _073_ vss 0.216342f
C16885 vdd _166_ 0.108744f
C16886 net55 FILLER_0_21_60/a_36_472# 0.06794f
C16887 FILLER_0_15_290/a_124_375# net62 0.034614f
C16888 net20 FILLER_0_12_236/a_36_472# 0.003143f
C16889 mask\[4\] net22 0.075713f
C16890 _430_/a_1000_472# mask\[2\] 0.00785f
C16891 FILLER_0_18_76/a_36_472# vss 0.007456f
C16892 _119_ _163_ 0.009297f
C16893 net54 FILLER_0_22_86/a_932_472# 0.047897f
C16894 _126_ _138_ 0.003253f
C16895 FILLER_0_21_142/a_572_375# _098_ 0.006558f
C16896 _429_/a_2560_156# vss 0.005255f
C16897 output29/a_224_472# net19 0.09445f
C16898 trim_mask\[1\] FILLER_0_4_91/a_36_472# 0.26171f
C16899 _064_ trim[1] 0.166575f
C16900 _423_/a_2665_112# vdd 0.022696f
C16901 _423_/a_2248_156# vss 0.010039f
C16902 _412_/a_36_151# net19 0.03393f
C16903 FILLER_0_12_220/a_124_375# _248_/a_36_68# 0.005308f
C16904 fanout68/a_36_113# net17 0.001252f
C16905 _414_/a_2248_156# _081_ 0.002027f
C16906 _093_ _303_/a_36_472# 0.096502f
C16907 net20 _103_ 0.261438f
C16908 net82 _316_/a_848_380# 0.087022f
C16909 result[4] vss 0.306116f
C16910 _093_ _102_ 0.008937f
C16911 _136_ FILLER_0_16_154/a_484_472# 0.007583f
C16912 mask\[5\] vdd 0.79138f
C16913 FILLER_0_20_169/a_124_375# vdd 0.03036f
C16914 output39/a_224_472# _445_/a_448_472# 0.009352f
C16915 FILLER_0_1_266/a_124_375# net8 0.012703f
C16916 FILLER_0_5_117/a_124_375# _119_ 0.002747f
C16917 _008_ _418_/a_1308_423# 0.027229f
C16918 net47 _450_/a_1353_112# 0.018879f
C16919 FILLER_0_12_136/a_1020_375# FILLER_0_13_142/a_484_472# 0.001684f
C16920 _024_ net33 0.001047f
C16921 FILLER_0_9_270/a_572_375# vdd 0.02345f
C16922 _070_ _310_/a_49_472# 0.00564f
C16923 _053_ _385_/a_36_68# 0.018437f
C16924 net79 _193_/a_36_160# 0.010228f
C16925 _413_/a_36_151# _079_ 0.0017f
C16926 _187_ net16 0.161791f
C16927 _176_ FILLER_0_11_109/a_36_472# 0.002951f
C16928 ctlp[1] _421_/a_796_472# 0.001754f
C16929 net66 vss 0.265973f
C16930 ctlp[1] fanout77/a_36_113# 0.012793f
C16931 net53 FILLER_0_13_142/a_124_375# 0.001599f
C16932 _442_/a_1000_472# vdd 0.003088f
C16933 _316_/a_692_472# _122_ 0.002929f
C16934 _316_/a_1152_472# calibrate 0.001604f
C16935 net15 _423_/a_1000_472# 0.001786f
C16936 fanout54/a_36_160# FILLER_0_19_142/a_36_472# 0.002647f
C16937 trim_mask\[1\] vdd 0.241393f
C16938 net20 _256_/a_716_497# 0.007413f
C16939 net4 _055_ 0.216844f
C16940 _114_ _307_/a_672_472# 0.0018f
C16941 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1468_375# 0.086635f
C16942 FILLER_0_4_197/a_932_472# net76 0.003693f
C16943 FILLER_0_19_55/a_124_375# vss 0.001882f
C16944 FILLER_0_19_55/a_36_472# vdd 0.085984f
C16945 FILLER_0_11_101/a_36_472# FILLER_0_13_100/a_124_375# 0.001436f
C16946 _372_/a_1602_69# _152_ 0.00262f
C16947 net80 _023_ 0.261119f
C16948 FILLER_0_20_87/a_36_472# net71 0.003995f
C16949 net50 _168_ 0.306226f
C16950 _055_ _311_/a_692_473# 0.003127f
C16951 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001597f
C16952 FILLER_0_15_282/a_36_472# _417_/a_1308_423# 0.001295f
C16953 _086_ _321_/a_2590_472# 0.001522f
C16954 net73 FILLER_0_18_107/a_124_375# 0.003742f
C16955 net75 FILLER_0_10_256/a_36_472# 0.010024f
C16956 _288_/a_224_472# _006_ 0.001278f
C16957 FILLER_0_7_104/a_1468_375# _133_ 0.003206f
C16958 _132_ _134_ 0.029512f
C16959 FILLER_0_7_72/a_2276_472# _439_/a_2248_156# 0.013656f
C16960 _129_ _062_ 0.20212f
C16961 _098_ FILLER_0_15_228/a_124_375# 0.080662f
C16962 _425_/a_36_151# vss 0.00158f
C16963 _425_/a_448_472# vdd 0.029071f
C16964 _077_ _453_/a_1000_472# 0.033726f
C16965 net32 _109_ 0.038411f
C16966 output21/a_224_472# _009_ 0.004164f
C16967 net23 _145_ 0.035734f
C16968 _003_ _081_ 0.041822f
C16969 mask\[7\] _435_/a_1000_472# 0.024725f
C16970 _093_ _198_/a_67_603# 0.004447f
C16971 _405_/a_67_603# net17 0.014714f
C16972 ctlp[2] net19 0.017506f
C16973 net54 mask\[8\] 0.162104f
C16974 FILLER_0_18_107/a_572_375# mask\[9\] 0.005368f
C16975 net52 _386_/a_124_24# 0.001051f
C16976 cal_count\[3\] _278_/a_36_160# 0.008398f
C16977 _223_/a_36_160# vdd 0.018653f
C16978 cal_count\[3\] FILLER_0_12_20/a_124_375# 0.008038f
C16979 net34 _421_/a_2665_112# 0.001056f
C16980 result[7] _421_/a_1204_472# 0.014927f
C16981 _164_ FILLER_0_6_47/a_36_472# 0.047981f
C16982 _067_ vss 0.20904f
C16983 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_36_472# 0.003468f
C16984 FILLER_0_11_124/a_36_472# _118_ 0.002798f
C16985 FILLER_0_17_282/a_36_472# net30 0.001189f
C16986 net15 _029_ 0.111797f
C16987 _144_ FILLER_0_21_125/a_484_472# 0.001616f
C16988 net4 FILLER_0_6_231/a_124_375# 0.002212f
C16989 net1 vss 0.161208f
C16990 _207_/a_67_603# _049_ 0.003205f
C16991 _299_/a_36_472# vdd 0.098451f
C16992 FILLER_0_4_107/a_484_472# _154_ 0.040595f
C16993 _420_/a_36_151# FILLER_0_23_282/a_572_375# 0.059049f
C16994 FILLER_0_21_286/a_36_472# _009_ 0.003266f
C16995 FILLER_0_14_99/a_124_375# vss 0.017196f
C16996 FILLER_0_14_99/a_36_472# vdd 0.095251f
C16997 _253_/a_36_68# vdd 0.016219f
C16998 mask\[5\] FILLER_0_18_177/a_1380_472# 0.001063f
C16999 net54 vss 0.715177f
C17000 FILLER_0_20_169/a_36_472# _140_ 0.023696f
C17001 _149_ FILLER_0_20_87/a_124_375# 0.004191f
C17002 mask\[3\] _093_ 2.443356f
C17003 net74 _067_ 0.674895f
C17004 FILLER_0_13_142/a_1380_472# _043_ 0.011974f
C17005 net32 _421_/a_2248_156# 0.038586f
C17006 _432_/a_2665_112# FILLER_0_18_177/a_2276_472# 0.021761f
C17007 net76 _122_ 0.028025f
C17008 _056_ _311_/a_254_473# 0.005937f
C17009 _053_ FILLER_0_6_177/a_572_375# 0.01663f
C17010 net28 fanout79/a_36_160# 0.036675f
C17011 FILLER_0_18_107/a_1020_375# FILLER_0_19_111/a_572_375# 0.05841f
C17012 FILLER_0_18_139/a_572_375# FILLER_0_19_142/a_124_375# 0.026339f
C17013 FILLER_0_15_72/a_572_375# _451_/a_3129_107# 0.007026f
C17014 net17 FILLER_0_20_15/a_1380_472# 0.012286f
C17015 _186_ _184_ 0.047995f
C17016 FILLER_0_24_63/a_124_375# ctlp[9] 0.002726f
C17017 output43/a_224_472# net43 0.11662f
C17018 _168_ trim_mask\[3\] 0.007154f
C17019 _069_ _247_/a_36_160# 0.046764f
C17020 net41 FILLER_0_21_28/a_1020_375# 0.010649f
C17021 _137_ _138_ 0.045916f
C17022 _339_/a_36_160# FILLER_0_19_171/a_124_375# 0.006021f
C17023 _434_/a_1308_423# mask\[6\] 0.022677f
C17024 FILLER_0_16_255/a_124_375# _094_ 0.004398f
C17025 FILLER_0_9_28/a_3172_472# vss 0.001977f
C17026 result[9] _421_/a_448_472# 0.015264f
C17027 _374_/a_36_68# _056_ 0.011052f
C17028 net79 _416_/a_448_472# 0.078357f
C17029 ctlp[1] FILLER_0_24_274/a_1380_472# 0.008573f
C17030 FILLER_0_20_107/a_36_472# net14 0.002543f
C17031 FILLER_0_3_142/a_124_375# net23 0.25251f
C17032 _429_/a_36_151# net79 0.02414f
C17033 net34 net22 0.031404f
C17034 trim_mask\[4\] _370_/a_1084_68# 0.005157f
C17035 net55 _404_/a_36_472# 0.001746f
C17036 FILLER_0_10_247/a_124_375# fanout79/a_36_160# 0.010334f
C17037 sample fanout65/a_36_113# 0.050978f
C17038 _142_ FILLER_0_16_154/a_124_375# 0.004001f
C17039 _136_ FILLER_0_13_100/a_36_472# 0.005029f
C17040 _307_/a_672_472# _126_ 0.00121f
C17041 FILLER_0_12_220/a_36_472# _070_ 0.087648f
C17042 ctlp[3] _422_/a_2665_112# 0.001024f
C17043 _444_/a_1000_472# net40 0.038229f
C17044 FILLER_0_15_290/a_124_375# FILLER_0_15_282/a_572_375# 0.012001f
C17045 FILLER_0_20_193/a_572_375# vss 0.005887f
C17046 FILLER_0_20_193/a_36_472# vdd 0.091886f
C17047 net75 net9 0.006945f
C17048 _072_ state\[1\] 0.267762f
C17049 fanout74/a_36_113# FILLER_0_3_142/a_124_375# 0.002073f
C17050 FILLER_0_10_256/a_36_472# _426_/a_36_151# 0.059238f
C17051 FILLER_0_16_73/a_572_375# _175_ 0.138524f
C17052 FILLER_0_17_200/a_124_375# vdd -0.010938f
C17053 FILLER_0_17_72/a_2276_472# _131_ 0.004125f
C17054 FILLER_0_7_146/a_124_375# net23 0.00129f
C17055 _074_ _375_/a_692_497# 0.004556f
C17056 _398_/a_36_113# vdd 0.030449f
C17057 FILLER_0_15_72/a_124_375# FILLER_0_13_72/a_36_472# 0.001418f
C17058 FILLER_0_9_105/a_36_472# vss 0.002744f
C17059 FILLER_0_9_105/a_484_472# vdd 0.03152f
C17060 _292_/a_36_160# _047_ 0.001291f
C17061 _196_/a_36_160# FILLER_0_14_263/a_124_375# 0.005732f
C17062 _032_ FILLER_0_2_127/a_124_375# 0.002221f
C17063 _410_/a_36_68# _042_ 0.041079f
C17064 _425_/a_2248_156# net19 0.010557f
C17065 _128_ _116_ 0.069335f
C17066 _127_ _176_ 0.319517f
C17067 ctlp[2] _009_ 0.220631f
C17068 FILLER_0_5_198/a_572_375# net59 0.00183f
C17069 _115_ _449_/a_2665_112# 0.00947f
C17070 FILLER_0_4_91/a_572_375# _156_ 0.004958f
C17071 FILLER_0_18_139/a_484_472# vss 0.006719f
C17072 FILLER_0_18_139/a_932_472# vdd 0.002904f
C17073 net65 FILLER_0_3_172/a_1916_375# 0.003745f
C17074 _136_ mask\[2\] 1.822289f
C17075 _121_ vss 0.082882f
C17076 FILLER_0_16_154/a_1020_375# vdd 0.004279f
C17077 FILLER_0_16_154/a_572_375# vss 0.003976f
C17078 _412_/a_448_472# cal_itt\[1\] 0.043203f
C17079 _086_ _268_/a_245_68# 0.001044f
C17080 net38 net44 0.523774f
C17081 output42/a_224_472# net40 0.003278f
C17082 _091_ FILLER_0_12_220/a_484_472# 0.001453f
C17083 net19 _420_/a_1308_423# 0.010051f
C17084 output37/a_224_472# output27/a_224_472# 0.012653f
C17085 output9/a_224_472# en 0.011047f
C17086 mask\[7\] FILLER_0_22_128/a_1380_472# 0.015814f
C17087 FILLER_0_8_127/a_124_375# _125_ 0.003105f
C17088 output29/a_224_472# _193_/a_36_160# 0.006363f
C17089 net16 net67 0.038448f
C17090 net40 _167_ 0.020177f
C17091 output27/a_224_472# net5 0.008663f
C17092 _320_/a_1792_472# state\[1\] 0.001901f
C17093 FILLER_0_7_104/a_572_375# vdd 0.038253f
C17094 _144_ _143_ 0.001774f
C17095 trim_mask\[2\] _167_ 0.027204f
C17096 _144_ _348_/a_49_472# 0.037768f
C17097 net20 _429_/a_2248_156# 0.027661f
C17098 fanout52/a_36_160# net23 0.009496f
C17099 _176_ _071_ 0.002542f
C17100 _436_/a_36_151# _050_ 0.037103f
C17101 net74 _370_/a_692_472# 0.005066f
C17102 _120_ _042_ 0.031451f
C17103 net31 _291_/a_36_160# 0.005683f
C17104 _306_/a_36_68# _071_ 0.054312f
C17105 net17 _190_/a_36_160# 0.04702f
C17106 FILLER_0_18_107/a_1468_375# vdd 0.004726f
C17107 _434_/a_448_472# _023_ 0.03093f
C17108 _413_/a_448_472# vdd 0.016117f
C17109 _413_/a_36_151# vss 0.003285f
C17110 trim_mask\[1\] FILLER_0_6_47/a_3172_472# 0.004605f
C17111 net82 _078_ 0.00197f
C17112 net31 net20 0.238809f
C17113 _049_ FILLER_0_22_128/a_3260_375# 0.16381f
C17114 _431_/a_448_472# _131_ 0.006194f
C17115 state\[1\] FILLER_0_13_142/a_1468_375# 0.010245f
C17116 net73 _022_ 0.003246f
C17117 net52 FILLER_0_2_165/a_124_375# 0.002214f
C17118 net54 FILLER_0_22_128/a_1020_375# 0.010068f
C17119 _448_/a_36_151# net22 0.027581f
C17120 FILLER_0_16_89/a_36_472# _451_/a_2449_156# 0.001571f
C17121 mask\[3\] FILLER_0_17_161/a_36_472# 0.13873f
C17122 result[9] FILLER_0_24_274/a_484_472# 0.003507f
C17123 FILLER_0_2_171/a_36_472# FILLER_0_2_177/a_36_472# 0.003468f
C17124 output8/a_224_472# vss 0.076244f
C17125 FILLER_0_17_200/a_36_472# net21 0.036768f
C17126 _421_/a_1000_472# net19 0.03394f
C17127 FILLER_0_20_15/a_1468_375# net40 0.030032f
C17128 _446_/a_2560_156# vdd 0.003959f
C17129 _446_/a_2665_112# vss 0.001781f
C17130 FILLER_0_10_37/a_124_375# net16 0.010358f
C17131 _421_/a_2665_112# _419_/a_2665_112# 0.002588f
C17132 _410_/a_36_68# cal_count\[3\] 0.001096f
C17133 FILLER_0_24_274/a_1020_375# vss 0.003553f
C17134 _414_/a_1308_423# vdd 0.004897f
C17135 FILLER_0_22_86/a_484_472# _437_/a_36_151# 0.013806f
C17136 FILLER_0_5_164/a_36_472# _386_/a_848_380# 0.001177f
C17137 FILLER_0_7_146/a_36_472# _313_/a_67_603# 0.002287f
C17138 FILLER_0_5_72/a_932_472# vss 0.003084f
C17139 FILLER_0_5_72/a_1380_472# vdd 0.001438f
C17140 net81 output37/a_224_472# 0.00641f
C17141 _128_ _117_ 0.045015f
C17142 _390_/a_36_68# vdd 0.012472f
C17143 _275_/a_224_472# _069_ 0.004466f
C17144 _148_ FILLER_0_22_107/a_572_375# 0.00652f
C17145 _093_ FILLER_0_16_89/a_124_375# 0.004086f
C17146 _449_/a_36_151# FILLER_0_12_50/a_36_472# 0.003462f
C17147 net81 net5 0.006276f
C17148 _289_/a_36_472# net30 0.009623f
C17149 _415_/a_796_472# vdd 0.001842f
C17150 _408_/a_718_524# vdd 0.002635f
C17151 _092_ FILLER_0_17_218/a_124_375# 0.020704f
C17152 net10 _411_/a_2248_156# 0.002419f
C17153 output10/a_224_472# FILLER_0_0_266/a_124_375# 0.00515f
C17154 fanout82/a_36_113# calibrate 0.004982f
C17155 net21 mask\[6\] 0.634881f
C17156 trimb[0] FILLER_0_20_2/a_36_472# 0.005458f
C17157 net16 FILLER_0_8_37/a_572_375# 0.004285f
C17158 _054_ vdd 0.360345f
C17159 _086_ _120_ 0.408014f
C17160 _420_/a_1308_423# _009_ 0.014359f
C17161 mask\[0\] FILLER_0_15_212/a_572_375# 0.001158f
C17162 _088_ net21 0.053843f
C17163 cal_count\[2\] vdd 0.932907f
C17164 _139_ net36 0.024268f
C17165 _176_ _451_/a_2449_156# 0.038547f
C17166 _411_/a_36_151# FILLER_0_0_232/a_36_472# 0.001723f
C17167 _029_ _163_ 0.007545f
C17168 FILLER_0_8_24/a_572_375# vss 0.012859f
C17169 FILLER_0_8_24/a_36_472# vdd 0.007423f
C17170 net20 _123_ 0.034801f
C17171 _443_/a_448_472# net23 0.038188f
C17172 FILLER_0_5_72/a_36_472# net15 0.006713f
C17173 FILLER_0_3_78/a_124_375# _160_ 0.003276f
C17174 net54 _026_ 0.006401f
C17175 net50 _441_/a_796_472# 0.010626f
C17176 net52 trim_mask\[2\] 0.036196f
C17177 FILLER_0_12_220/a_572_375# vdd -0.014642f
C17178 FILLER_0_12_220/a_124_375# vss 0.040895f
C17179 cal_count\[3\] _120_ 4.687877f
C17180 FILLER_0_15_150/a_124_375# _427_/a_36_151# 0.001822f
C17181 FILLER_0_13_212/a_1468_375# net79 0.009597f
C17182 FILLER_0_4_49/a_572_375# net66 0.074393f
C17183 FILLER_0_2_101/a_124_375# _160_ 0.001047f
C17184 net26 vss 0.263774f
C17185 output23/a_224_472# net23 0.122379f
C17186 FILLER_0_4_107/a_1020_375# _160_ 0.015684f
C17187 trim_mask\[4\] net47 0.264421f
C17188 _195_/a_67_603# mask\[1\] 0.016836f
C17189 _155_ vss 0.13648f
C17190 _093_ FILLER_0_18_76/a_484_472# 0.024853f
C17191 _105_ _109_ 0.107328f
C17192 ctlp[5] net23 0.025206f
C17193 FILLER_0_8_37/a_124_375# vdd 0.029725f
C17194 fanout81/a_36_160# net9 0.002274f
C17195 FILLER_0_11_124/a_36_472# vdd 0.005222f
C17196 FILLER_0_11_124/a_124_375# vss 0.017354f
C17197 net47 FILLER_0_4_91/a_124_375# 0.009482f
C17198 net50 _440_/a_2665_112# 0.009767f
C17199 _115_ vss 0.372063f
C17200 output29/a_224_472# _416_/a_448_472# 0.008149f
C17201 FILLER_0_4_49/a_124_375# trim_mask\[1\] 0.006676f
C17202 net52 _439_/a_1000_472# 0.03537f
C17203 net50 _439_/a_1308_423# 0.008832f
C17204 output44/a_224_472# FILLER_0_18_2/a_2364_375# 0.032639f
C17205 trimb[1] FILLER_0_18_2/a_124_375# 0.01352f
C17206 _053_ FILLER_0_7_72/a_2276_472# 0.016004f
C17207 fanout73/a_36_113# _136_ 0.002661f
C17208 mask\[4\] FILLER_0_18_177/a_932_472# 0.016924f
C17209 FILLER_0_9_28/a_2364_375# _053_ 0.029866f
C17210 mask\[4\] _140_ 0.001697f
C17211 FILLER_0_18_209/a_124_375# _047_ 0.006317f
C17212 _143_ _339_/a_36_160# 0.00507f
C17213 output18/a_224_472# vdd -0.01545f
C17214 FILLER_0_17_72/a_932_472# _175_ 0.003281f
C17215 _063_ _160_ 0.091185f
C17216 FILLER_0_5_212/a_36_472# net22 0.0015f
C17217 FILLER_0_6_239/a_36_472# _074_ 0.004715f
C17218 _434_/a_1000_472# vdd 0.032431f
C17219 net74 FILLER_0_11_124/a_124_375# 0.047331f
C17220 _340_/a_36_160# vdd 0.006001f
C17221 FILLER_0_12_136/a_1020_375# vdd 0.017472f
C17222 FILLER_0_12_136/a_572_375# vss 0.006091f
C17223 net41 net40 2.687418f
C17224 _417_/a_36_151# vss 0.040392f
C17225 _030_ FILLER_0_3_78/a_124_375# 0.010439f
C17226 _053_ FILLER_0_7_162/a_124_375# 0.007494f
C17227 _115_ net74 0.033145f
C17228 net69 FILLER_0_2_111/a_484_472# 0.010567f
C17229 _031_ FILLER_0_2_111/a_1468_375# 0.013595f
C17230 _076_ _059_ 1.03702f
C17231 _065_ _441_/a_2665_112# 0.003318f
C17232 fanout52/a_36_160# trim_val\[4\] 0.019286f
C17233 net75 _084_ 0.045583f
C17234 net58 cal_itt\[1\] 0.79493f
C17235 net55 net44 0.018961f
C17236 fanout76/a_36_160# net4 0.002206f
C17237 net54 _211_/a_36_160# 0.001244f
C17238 _069_ FILLER_0_13_206/a_124_375# 0.009695f
C17239 _065_ _447_/a_1000_472# 0.03162f
C17240 net41 FILLER_0_18_2/a_3260_375# 0.042057f
C17241 _072_ FILLER_0_7_233/a_124_375# 0.002279f
C17242 FILLER_0_5_54/a_1380_472# vss 0.007301f
C17243 FILLER_0_4_123/a_124_375# _370_/a_124_24# 0.007188f
C17244 cal_count\[2\] _452_/a_1040_527# 0.002003f
C17245 _195_/a_67_603# vss 0.002638f
C17246 _119_ _121_ 0.007336f
C17247 _437_/a_36_151# vdd 0.115376f
C17248 FILLER_0_10_28/a_124_375# net6 0.007948f
C17249 _096_ _320_/a_1792_472# 0.001419f
C17250 net58 valid 0.149817f
C17251 _003_ _161_ 0.004981f
C17252 cal_itt\[2\] net58 0.003431f
C17253 valid _425_/a_2665_112# 0.001839f
C17254 _440_/a_2560_156# _164_ 0.003934f
C17255 _242_/a_36_160# FILLER_0_5_148/a_572_375# 0.00805f
C17256 FILLER_0_14_91/a_124_375# _095_ 0.01418f
C17257 FILLER_0_1_212/a_36_472# net59 0.002567f
C17258 _424_/a_2248_156# net36 0.017101f
C17259 FILLER_0_17_200/a_572_375# net63 0.007512f
C17260 _158_ _160_ 0.018681f
C17261 _151_ _365_/a_36_68# 0.001944f
C17262 _005_ net19 0.033451f
C17263 _253_/a_1100_68# _084_ 0.001651f
C17264 FILLER_0_7_72/a_1828_472# net50 0.094122f
C17265 net27 result[0] 0.106157f
C17266 net54 _433_/a_448_472# 0.008777f
C17267 FILLER_0_23_44/a_572_375# vdd -0.011314f
C17268 result[7] FILLER_0_23_282/a_572_375# 0.015853f
C17269 fanout54/a_36_160# _433_/a_2248_156# 0.012122f
C17270 net81 FILLER_0_15_212/a_484_472# 0.00169f
C17271 FILLER_0_2_177/a_484_472# net59 0.007829f
C17272 FILLER_0_10_28/a_36_472# net40 0.020589f
C17273 _177_ vdd 0.111636f
C17274 cal_itt\[3\] _055_ 0.007428f
C17275 net55 _176_ 0.300149f
C17276 net70 FILLER_0_14_107/a_932_472# 0.008396f
C17277 net53 FILLER_0_14_107/a_1468_375# 0.001642f
C17278 net32 result[9] 0.001371f
C17279 _021_ _141_ 0.047816f
C17280 FILLER_0_17_72/a_3172_472# FILLER_0_17_104/a_36_472# 0.013277f
C17281 _053_ FILLER_0_7_59/a_484_472# 0.013665f
C17282 net15 FILLER_0_5_54/a_484_472# 0.002186f
C17283 FILLER_0_8_263/a_36_472# calibrate 0.006968f
C17284 FILLER_0_20_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001543f
C17285 FILLER_0_19_47/a_124_375# FILLER_0_18_37/a_1380_472# 0.001684f
C17286 _412_/a_448_472# net59 0.001462f
C17287 _247_/a_36_160# _090_ 0.010285f
C17288 FILLER_0_4_177/a_36_472# net76 0.003007f
C17289 output32/a_224_472# vss -0.003023f
C17290 ctlp[8] net35 0.001859f
C17291 FILLER_0_17_38/a_484_472# vdd 0.009211f
C17292 trim_val\[0\] FILLER_0_6_47/a_484_472# 0.001215f
C17293 trim_val\[4\] _443_/a_448_472# 0.038063f
C17294 FILLER_0_14_81/a_36_472# _043_ 0.001714f
C17295 output36/a_224_472# result[9] 0.059164f
C17296 net3 FILLER_0_15_2/a_484_472# 0.002224f
C17297 _098_ _433_/a_1204_472# 0.014374f
C17298 FILLER_0_18_2/a_484_472# net44 0.047503f
C17299 FILLER_0_1_98/a_124_375# net52 0.001167f
C17300 _414_/a_36_151# _086_ 0.002687f
C17301 FILLER_0_16_241/a_124_375# _099_ 0.040547f
C17302 ctlp[1] net19 0.029153f
C17303 net34 FILLER_0_22_177/a_1380_472# 0.003953f
C17304 _077_ _439_/a_36_151# 0.035432f
C17305 net47 _452_/a_448_472# 0.005335f
C17306 mask\[9\] _438_/a_1204_472# 0.03521f
C17307 _395_/a_36_488# _085_ 0.020572f
C17308 _247_/a_36_160# net22 0.048614f
C17309 FILLER_0_22_86/a_124_375# FILLER_0_23_88/a_36_472# 0.001684f
C17310 FILLER_0_3_172/a_2812_375# net22 0.013048f
C17311 net54 FILLER_0_19_134/a_36_472# 0.061344f
C17312 _064_ _034_ 1.397143f
C17313 _346_/a_257_69# mask\[5\] 0.001764f
C17314 output22/a_224_472# net80 0.00955f
C17315 _430_/a_36_151# _092_ 0.002363f
C17316 _053_ FILLER_0_7_146/a_124_375# 0.005844f
C17317 _176_ net23 0.036283f
C17318 net7 net40 0.025164f
C17319 comp FILLER_0_12_2/a_36_472# 0.003875f
C17320 FILLER_0_14_81/a_36_472# _175_ 0.076977f
C17321 FILLER_0_21_133/a_36_472# vss 0.004298f
C17322 net35 net21 0.001845f
C17323 net75 output28/a_224_472# 0.00151f
C17324 _052_ FILLER_0_18_53/a_124_375# 0.001585f
C17325 ctln[3] _411_/a_36_151# 0.004014f
C17326 _016_ cal_count\[3\] 0.004588f
C17327 state\[2\] state\[1\] 0.229832f
C17328 net20 FILLER_0_24_274/a_124_375# 0.002751f
C17329 FILLER_0_3_204/a_36_472# FILLER_0_3_212/a_36_472# 0.002296f
C17330 FILLER_0_5_128/a_124_375# net47 0.011156f
C17331 cal_count\[3\] _408_/a_56_524# 0.001685f
C17332 _413_/a_36_151# FILLER_0_3_172/a_3172_472# 0.001723f
C17333 _438_/a_2665_112# FILLER_0_19_111/a_124_375# 0.006271f
C17334 _069_ FILLER_0_13_212/a_124_375# 0.070185f
C17335 net50 FILLER_0_7_59/a_36_472# 0.01018f
C17336 _411_/a_2560_156# _073_ 0.002649f
C17337 _412_/a_1000_472# net76 0.024114f
C17338 _204_/a_67_603# _201_/a_67_603# 0.001129f
C17339 _067_ _389_/a_36_148# 0.002789f
C17340 _328_/a_36_113# _132_ 0.006002f
C17341 net44 FILLER_0_15_10/a_36_472# 0.012286f
C17342 FILLER_0_17_200/a_124_375# _093_ 0.00419f
C17343 FILLER_0_18_100/a_36_472# FILLER_0_18_107/a_36_472# 0.002764f
C17344 net58 _416_/a_36_151# 0.001558f
C17345 _359_/a_36_488# _131_ 0.006398f
C17346 net34 _140_ 0.033459f
C17347 _098_ FILLER_0_20_87/a_124_375# 0.019333f
C17348 net11 vdd 0.330644f
C17349 _165_ _377_/a_36_472# 0.025689f
C17350 _287_/a_36_472# mask\[2\] 0.00492f
C17351 output9/a_224_472# cal 0.011495f
C17352 net36 FILLER_0_15_205/a_124_375# 0.004337f
C17353 _081_ cal_itt\[0\] 0.036569f
C17354 _431_/a_448_472# _137_ 0.008493f
C17355 _233_/a_36_160# FILLER_0_6_37/a_36_472# 0.012692f
C17356 net25 _098_ 0.001267f
C17357 net33 _107_ 0.001322f
C17358 FILLER_0_19_47/a_484_472# _012_ 0.001667f
C17359 net69 _441_/a_448_472# 0.028545f
C17360 _119_ _115_ 0.06747f
C17361 _138_ mask\[1\] 0.085445f
C17362 net36 _098_ 3.387566f
C17363 FILLER_0_17_226/a_124_375# FILLER_0_17_218/a_572_375# 0.012001f
C17364 _106_ fanout63/a_36_160# 0.00715f
C17365 net52 FILLER_0_3_142/a_36_472# 0.001122f
C17366 trimb[4] net17 0.004628f
C17367 _447_/a_2665_112# _030_ 0.001226f
C17368 net32 _048_ 0.008647f
C17369 net71 _437_/a_1308_423# 0.023981f
C17370 FILLER_0_12_136/a_932_472# _127_ 0.002804f
C17371 _445_/a_36_151# net66 0.058093f
C17372 net66 _029_ 0.056971f
C17373 _064_ _445_/a_2248_156# 0.013127f
C17374 _447_/a_1000_472# _036_ 0.002902f
C17375 _261_/a_36_160# FILLER_0_5_148/a_124_375# 0.005705f
C17376 cal_itt\[3\] _058_ 0.002207f
C17377 FILLER_0_7_72/a_932_472# _077_ 0.001315f
C17378 result[5] _418_/a_2248_156# 0.001309f
C17379 FILLER_0_20_177/a_1380_472# vdd 0.009871f
C17380 FILLER_0_20_177/a_932_472# vss 0.001272f
C17381 net41 net46 0.061224f
C17382 FILLER_0_7_195/a_124_375# _074_ 0.019559f
C17383 _436_/a_448_472# net54 0.006129f
C17384 net69 _157_ 0.112249f
C17385 _232_/a_67_603# vss 0.00988f
C17386 _004_ net27 0.080285f
C17387 FILLER_0_18_100/a_124_375# _136_ 0.002528f
C17388 _127_ _017_ 0.005836f
C17389 ctlp[1] _009_ 0.085933f
C17390 net55 _183_ 0.024948f
C17391 FILLER_0_14_263/a_36_472# vss 0.003195f
C17392 _450_/a_1040_527# output6/a_224_472# 0.005581f
C17393 _450_/a_36_151# net6 0.035997f
C17394 _046_ _099_ 0.005245f
C17395 FILLER_0_16_107/a_484_472# _451_/a_36_151# 0.027244f
C17396 _116_ _311_/a_2700_473# 0.001555f
C17397 FILLER_0_10_78/a_36_472# net52 0.014225f
C17398 FILLER_0_12_136/a_124_375# cal_count\[3\] 0.005006f
C17399 output33/a_224_472# output19/a_224_472# 0.115114f
C17400 FILLER_0_18_177/a_1020_375# vdd 0.040478f
C17401 _132_ _428_/a_36_151# 0.013691f
C17402 FILLER_0_20_193/a_124_375# FILLER_0_19_195/a_36_472# 0.001543f
C17403 FILLER_0_2_101/a_124_375# _156_ 0.022015f
C17404 net82 FILLER_0_3_212/a_124_375# 0.015932f
C17405 net63 net36 0.010544f
C17406 _081_ FILLER_0_6_177/a_484_472# 0.010037f
C17407 _418_/a_36_151# vss 0.041728f
C17408 _150_ net14 0.001303f
C17409 _411_/a_1308_423# _000_ 0.004012f
C17410 _411_/a_1000_472# net75 0.03227f
C17411 _074_ _312_/a_672_472# 0.005399f
C17412 _419_/a_2248_156# vdd 0.040646f
C17413 FILLER_0_10_256/a_124_375# net19 0.002884f
C17414 _420_/a_36_151# FILLER_0_23_290/a_36_472# 0.001723f
C17415 FILLER_0_14_91/a_572_375# vdd -0.011429f
C17416 _413_/a_2665_112# cal_itt\[2\] 0.003007f
C17417 _053_ FILLER_0_6_90/a_484_472# 0.011443f
C17418 _014_ FILLER_0_7_233/a_36_472# 0.002089f
C17419 _450_/a_448_472# net40 0.00222f
C17420 net19 FILLER_0_23_282/a_124_375# 0.001668f
C17421 net60 output18/a_224_472# 0.001518f
C17422 _028_ net50 0.087995f
C17423 _106_ FILLER_0_17_218/a_484_472# 0.012952f
C17424 _138_ vss 0.006962f
C17425 net16 trim_val\[1\] 0.164715f
C17426 _326_/a_36_160# _128_ 0.02761f
C17427 _149_ _437_/a_448_472# 0.009274f
C17428 _453_/a_1000_472# vss 0.001738f
C17429 _095_ _451_/a_1353_112# 0.00475f
C17430 _012_ FILLER_0_21_60/a_124_375# 0.016032f
C17431 _086_ _151_ 0.002442f
C17432 net75 calibrate 0.101912f
C17433 _002_ _087_ 0.00636f
C17434 mask\[5\] output33/a_224_472# 0.0238f
C17435 net58 net59 0.066534f
C17436 FILLER_0_15_212/a_1468_375# mask\[1\] 0.045287f
C17437 _348_/a_665_69# _146_ 0.001153f
C17438 _432_/a_36_151# _337_/a_49_472# 0.002462f
C17439 FILLER_0_13_142/a_124_375# net23 0.003962f
C17440 _425_/a_796_472# _122_ 0.001701f
C17441 _425_/a_36_151# _123_ 0.006319f
C17442 _425_/a_1000_472# calibrate 0.027245f
C17443 net41 trim[3] 0.005906f
C17444 FILLER_0_20_2/a_124_375# vdd 0.010886f
C17445 net58 net4 0.858616f
C17446 net47 _066_ 0.096823f
C17447 FILLER_0_20_169/a_36_472# _098_ 0.007354f
C17448 FILLER_0_3_2/a_124_375# output41/a_224_472# 0.030009f
C17449 FILLER_0_5_212/a_124_375# vdd 0.024541f
C17450 FILLER_0_18_177/a_2276_472# net21 0.01016f
C17451 _438_/a_2665_112# vdd 0.00587f
C17452 _438_/a_2248_156# vss 0.002607f
C17453 FILLER_0_17_72/a_124_375# FILLER_0_17_64/a_124_375# 0.003732f
C17454 FILLER_0_13_212/a_572_375# net62 0.001597f
C17455 _063_ net67 0.039144f
C17456 _011_ _422_/a_1204_472# 0.002176f
C17457 FILLER_0_1_266/a_124_375# vdd -0.002281f
C17458 FILLER_0_8_107/a_36_472# _062_ 0.001832f
C17459 _410_/a_36_68# _120_ 0.073688f
C17460 _431_/a_448_472# net56 0.001464f
C17461 FILLER_0_12_124/a_36_472# _127_ 0.01468f
C17462 net56 FILLER_0_19_142/a_124_375# 0.003154f
C17463 FILLER_0_15_282/a_484_472# _006_ 0.00444f
C17464 _151_ _154_ 0.108571f
C17465 _250_/a_36_68# _071_ 0.199512f
C17466 _070_ FILLER_0_7_233/a_36_472# 0.07194f
C17467 FILLER_0_9_28/a_932_472# net68 0.003603f
C17468 _072_ _374_/a_36_68# 0.061028f
C17469 _005_ _193_/a_36_160# 0.009892f
C17470 net73 FILLER_0_18_107/a_3172_472# 0.00533f
C17471 net15 _453_/a_1308_423# 0.00293f
C17472 FILLER_0_7_72/a_3172_472# trim_mask\[0\] 0.001438f
C17473 _229_/a_224_472# net22 0.007346f
C17474 _091_ FILLER_0_10_214/a_124_375# 0.006331f
C17475 _095_ net17 0.172789f
C17476 net48 _076_ 0.077031f
C17477 result[8] FILLER_0_24_274/a_36_472# 0.005458f
C17478 FILLER_0_13_228/a_124_375# FILLER_0_12_220/a_1020_375# 0.05841f
C17479 FILLER_0_21_125/a_484_472# mask\[7\] 0.003404f
C17480 net47 net37 0.057409f
C17481 net50 FILLER_0_6_90/a_36_472# 0.049285f
C17482 FILLER_0_6_47/a_2364_375# vss 0.008275f
C17483 FILLER_0_6_47/a_2812_375# vdd 0.002455f
C17484 FILLER_0_15_212/a_1468_375# vss 0.060206f
C17485 FILLER_0_15_212/a_36_472# vdd 0.105575f
C17486 cal_count\[3\] _043_ 0.721078f
C17487 FILLER_0_18_177/a_3260_375# _205_/a_36_160# 0.001313f
C17488 output32/a_224_472# _103_ 0.090957f
C17489 _402_/a_56_567# vdd 0.014708f
C17490 _426_/a_3041_156# net64 0.001046f
C17491 net73 FILLER_0_17_133/a_36_472# 0.049294f
C17492 net32 net61 0.056005f
C17493 _208_/a_36_160# _049_ 0.04568f
C17494 FILLER_0_6_239/a_124_375# _316_/a_124_24# 0.003524f
C17495 net53 _451_/a_2225_156# 0.011677f
C17496 _009_ FILLER_0_23_282/a_124_375# 0.012402f
C17497 _127_ FILLER_0_11_135/a_124_375# 0.040456f
C17498 FILLER_0_4_197/a_124_375# net22 0.00145f
C17499 FILLER_0_8_247/a_1468_375# calibrate 0.006404f
C17500 fanout50/a_36_160# net50 0.052685f
C17501 _077_ FILLER_0_10_78/a_124_375# 0.001886f
C17502 FILLER_0_17_104/a_484_472# net14 0.004272f
C17503 ctln[5] vdd 0.256793f
C17504 _422_/a_36_151# mask\[7\] 0.043316f
C17505 _159_ vdd 0.025131f
C17506 net52 _443_/a_1308_423# 0.02003f
C17507 _131_ net36 0.068899f
C17508 output39/a_224_472# _033_ 0.045759f
C17509 _058_ trim_mask\[0\] 0.076069f
C17510 _426_/a_36_151# calibrate 0.004525f
C17511 _324_/a_224_472# _070_ 0.00142f
C17512 FILLER_0_13_206/a_124_375# net22 0.024537f
C17513 _077_ FILLER_0_9_72/a_36_472# 0.006408f
C17514 net15 FILLER_0_6_47/a_1468_375# 0.007439f
C17515 result[9] _010_ 0.121471f
C17516 _453_/a_796_472# _042_ 0.005463f
C17517 _453_/a_1308_423# net51 0.001804f
C17518 mask\[5\] _343_/a_49_472# 0.002228f
C17519 _346_/a_49_472# mask\[4\] 0.079347f
C17520 _402_/a_728_93# cal_count\[1\] 0.057043f
C17521 FILLER_0_18_53/a_572_375# vss 0.057185f
C17522 FILLER_0_18_53/a_36_472# vdd 0.089087f
C17523 _415_/a_448_472# result[1] 0.005209f
C17524 FILLER_0_16_89/a_572_375# _131_ 0.012481f
C17525 _086_ _375_/a_960_497# 0.001454f
C17526 _077_ _078_ 0.069858f
C17527 _433_/a_796_472# _022_ 0.025882f
C17528 FILLER_0_4_107/a_572_375# net47 0.006041f
C17529 _093_ _437_/a_36_151# 0.056554f
C17530 _104_ FILLER_0_17_226/a_124_375# 0.024833f
C17531 FILLER_0_3_172/a_2364_375# vdd -0.010717f
C17532 _178_ FILLER_0_15_10/a_124_375# 0.002355f
C17533 FILLER_0_21_206/a_36_472# net21 0.132984f
C17534 net32 _108_ 0.035815f
C17535 FILLER_0_9_223/a_124_375# _070_ 0.002989f
C17536 _449_/a_1000_472# net72 0.001247f
C17537 _449_/a_448_472# net55 0.004439f
C17538 net7 trim[3] 0.044017f
C17539 _053_ _257_/a_36_472# 0.00507f
C17540 _438_/a_448_472# net14 0.020612f
C17541 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1380_472# 0.026657f
C17542 FILLER_0_8_239/a_124_375# calibrate 0.008393f
C17543 output14/a_224_472# vss 0.012129f
C17544 FILLER_0_10_78/a_932_472# _176_ 0.0109f
C17545 _431_/a_36_151# FILLER_0_18_107/a_2724_472# 0.00271f
C17546 _413_/a_1308_423# net82 0.003079f
C17547 net55 FILLER_0_17_72/a_1468_375# 0.014449f
C17548 _131_ FILLER_0_14_123/a_124_375# 0.016964f
C17549 _446_/a_1204_472# net66 0.001885f
C17550 _305_/a_36_159# _425_/a_36_151# 0.001404f
C17551 _115_ _389_/a_36_148# 0.029505f
C17552 net73 FILLER_0_19_111/a_484_472# 0.007404f
C17553 FILLER_0_5_72/a_572_375# net49 0.001158f
C17554 _062_ _226_/a_276_68# 0.001286f
C17555 _005_ _416_/a_448_472# 0.04044f
C17556 net56 FILLER_0_19_155/a_36_472# 0.00611f
C17557 _093_ _177_ 0.001194f
C17558 FILLER_0_3_221/a_1380_472# vss 0.002804f
C17559 _131_ _160_ 0.003984f
C17560 FILLER_0_24_96/a_36_472# net14 0.002882f
C17561 _297_/a_36_472# vdd 0.042391f
C17562 en_co_clk FILLER_0_13_100/a_124_375# 0.002325f
C17563 FILLER_0_16_73/a_36_472# net15 0.005297f
C17564 FILLER_0_19_47/a_572_375# _052_ 0.020156f
C17565 FILLER_0_20_193/a_484_472# _098_ 0.012457f
C17566 _431_/a_36_151# FILLER_0_17_133/a_124_375# 0.059049f
C17567 _451_/a_1040_527# vdd 0.004038f
C17568 FILLER_0_5_72/a_932_472# _029_ 0.007801f
C17569 FILLER_0_5_72/a_1468_375# trim_mask\[1\] 0.017105f
C17570 net81 en 0.071123f
C17571 _086_ _267_/a_1568_472# 0.002143f
C17572 net26 _423_/a_1000_472# 0.001338f
C17573 _413_/a_2665_112# net59 0.066623f
C17574 _305_/a_36_159# net1 0.013619f
C17575 _431_/a_1204_472# _136_ 0.007382f
C17576 net22 _435_/a_448_472# 0.001929f
C17577 _105_ _048_ 0.02699f
C17578 net57 FILLER_0_16_154/a_1020_375# 0.001902f
C17579 FILLER_0_17_218/a_572_375# _069_ 0.001464f
C17580 _350_/a_49_472# vss 0.001319f
C17581 net51 _450_/a_2225_156# 0.009822f
C17582 FILLER_0_15_116/a_36_472# _040_ 0.002896f
C17583 FILLER_0_2_111/a_932_472# vdd 0.003808f
C17584 FILLER_0_2_111/a_484_472# vss -0.001894f
C17585 _043_ _278_/a_36_160# 0.004357f
C17586 _053_ _220_/a_67_603# 0.065611f
C17587 _114_ _116_ 0.038641f
C17588 net45 trimb[3] 0.001109f
C17589 net34 result[8] 0.076645f
C17590 _098_ FILLER_0_16_154/a_1468_375# 0.009042f
C17591 _065_ _164_ 0.006953f
C17592 _099_ net62 0.062012f
C17593 _103_ _418_/a_36_151# 0.032388f
C17594 net54 FILLER_0_18_107/a_124_375# 0.001636f
C17595 net41 FILLER_0_18_37/a_124_375# 0.004639f
C17596 _091_ _429_/a_36_151# 0.006557f
C17597 net60 _418_/a_448_472# 0.055895f
C17598 fanout62/a_36_160# vdd 0.059299f
C17599 _002_ vdd 0.152662f
C17600 _185_ _278_/a_36_160# 0.001237f
C17601 net60 _419_/a_2248_156# 0.047724f
C17602 net78 _419_/a_2248_156# 0.001614f
C17603 net61 _419_/a_2560_156# 0.008214f
C17604 _136_ FILLER_0_15_180/a_572_375# 0.001571f
C17605 FILLER_0_5_88/a_124_375# _164_ 0.006288f
C17606 _020_ _131_ 0.011012f
C17607 net63 FILLER_0_20_193/a_484_472# 0.015851f
C17608 net17 vss 0.940703f
C17609 _322_/a_1084_68# _128_ 0.002629f
C17610 FILLER_0_20_169/a_124_375# _434_/a_36_151# 0.026916f
C17611 mask\[5\] _434_/a_36_151# 0.00104f
C17612 FILLER_0_11_101/a_124_375# _058_ 0.002209f
C17613 FILLER_0_24_63/a_124_375# output25/a_224_472# 0.007304f
C17614 FILLER_0_21_28/a_2724_472# _012_ 0.020109f
C17615 _383_/a_36_472# trim_mask\[3\] 0.003193f
C17616 _320_/a_1568_472# net79 0.001157f
C17617 _155_ _029_ 0.174512f
C17618 FILLER_0_21_150/a_124_375# vss 0.013882f
C17619 FILLER_0_21_150/a_36_472# vdd 0.092128f
C17620 FILLER_0_4_99/a_124_375# FILLER_0_4_91/a_572_375# 0.012001f
C17621 FILLER_0_12_136/a_932_472# net23 0.004375f
C17622 net41 FILLER_0_10_28/a_124_375# 0.003909f
C17623 _408_/a_728_93# _067_ 0.006262f
C17624 _414_/a_2248_156# _056_ 0.001452f
C17625 mask\[4\] _098_ 0.041526f
C17626 sample valid 0.103192f
C17627 FILLER_0_7_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001723f
C17628 FILLER_0_15_142/a_36_472# net36 0.015456f
C17629 _099_ FILLER_0_15_235/a_572_375# 0.001327f
C17630 _176_ FILLER_0_15_72/a_36_472# 0.002101f
C17631 _051_ net71 0.001617f
C17632 _444_/a_2248_156# FILLER_0_6_37/a_124_375# 0.001101f
C17633 net4 _070_ 0.169392f
C17634 FILLER_0_21_142/a_124_375# net35 0.00123f
C17635 output10/a_224_472# net8 0.010088f
C17636 _087_ net76 0.529571f
C17637 net4 FILLER_0_12_220/a_1380_472# 0.016375f
C17638 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_36_472# 0.086743f
C17639 net57 _390_/a_36_68# 0.001112f
C17640 net66 FILLER_0_5_54/a_484_472# 0.001863f
C17641 _423_/a_36_151# FILLER_0_23_44/a_36_472# 0.001723f
C17642 FILLER_0_7_104/a_932_472# _058_ 0.002096f
C17643 _394_/a_1336_472# _175_ 0.002792f
C17644 _076_ _311_/a_66_473# 0.003077f
C17645 FILLER_0_15_116/a_572_375# net36 0.007321f
C17646 _427_/a_1308_423# _095_ 0.022677f
C17647 _000_ FILLER_0_0_232/a_124_375# 0.001391f
C17648 net68 FILLER_0_5_54/a_1020_375# 0.00648f
C17649 _431_/a_2248_156# net53 0.003335f
C17650 net73 _427_/a_36_151# 0.006328f
C17651 net9 cal_itt\[1\] 0.028339f
C17652 _081_ FILLER_0_5_198/a_572_375# 0.001285f
C17653 _091_ _055_ 0.003332f
C17654 _250_/a_36_68# net23 0.002628f
C17655 _032_ net23 0.019676f
C17656 FILLER_0_5_54/a_36_472# trim_mask\[1\] 0.101342f
C17657 FILLER_0_5_54/a_1380_472# _029_ 0.01027f
C17658 FILLER_0_9_28/a_932_472# FILLER_0_10_37/a_36_472# 0.026657f
C17659 FILLER_0_21_142/a_572_375# vss 0.097474f
C17660 FILLER_0_21_142/a_36_472# vdd 0.111749f
C17661 _441_/a_36_151# _440_/a_1308_423# 0.001736f
C17662 _091_ FILLER_0_15_180/a_36_472# 0.00375f
C17663 result[7] FILLER_0_23_290/a_36_472# 0.013403f
C17664 FILLER_0_9_28/a_1828_472# _054_ 0.003145f
C17665 net79 FILLER_0_15_282/a_124_375# 0.001058f
C17666 net63 mask\[4\] 0.043339f
C17667 _137_ _334_/a_36_160# 0.015722f
C17668 net17 _452_/a_836_156# 0.002817f
C17669 _374_/a_244_472# _076_ 0.001567f
C17670 _114_ _117_ 0.008886f
C17671 _161_ FILLER_0_6_177/a_484_472# 0.001723f
C17672 _128_ _247_/a_36_160# 0.00163f
C17673 FILLER_0_17_72/a_2724_472# vdd 0.007064f
C17674 FILLER_0_17_72/a_2276_472# vss -0.001288f
C17675 _027_ FILLER_0_18_76/a_484_472# 0.00705f
C17676 mask\[1\] FILLER_0_15_228/a_124_375# 0.013558f
C17677 FILLER_0_16_37/a_36_472# vss 0.005874f
C17678 fanout74/a_36_113# _032_ 0.012909f
C17679 _069_ _085_ 0.032519f
C17680 _429_/a_2665_112# _043_ 0.007641f
C17681 output9/a_224_472# fanout81/a_36_160# 0.012218f
C17682 net20 mask\[0\] 0.103301f
C17683 net65 ctln[4] 0.020799f
C17684 FILLER_0_8_127/a_36_472# _133_ 0.004423f
C17685 net20 _074_ 0.038279f
C17686 _122_ net47 0.030693f
C17687 FILLER_0_19_195/a_36_472# net21 0.009159f
C17688 output11/a_224_472# net11 0.003448f
C17689 output31/a_224_472# output36/a_224_472# 0.00289f
C17690 _140_ _146_ 0.135012f
C17691 _105_ net61 0.020753f
C17692 cal_itt\[3\] FILLER_0_5_164/a_484_472# 0.001518f
C17693 FILLER_0_21_286/a_572_375# net62 0.003744f
C17694 _431_/a_36_151# _142_ 0.030496f
C17695 _069_ _018_ 0.002777f
C17696 ctln[8] net14 0.001447f
C17697 _245_/a_234_472# net47 0.00188f
C17698 _006_ vdd 0.632993f
C17699 _294_/a_224_472# vss 0.001022f
C17700 _136_ _337_/a_257_69# 0.002933f
C17701 net16 _447_/a_36_151# 0.133348f
C17702 FILLER_0_1_192/a_36_472# vss 0.004422f
C17703 FILLER_0_4_213/a_484_472# net59 0.048997f
C17704 FILLER_0_9_142/a_124_375# _313_/a_67_603# 0.029786f
C17705 output33/a_224_472# output18/a_224_472# 0.111946f
C17706 FILLER_0_18_171/a_36_472# mask\[4\] 0.01222f
C17707 FILLER_0_3_2/a_36_472# net66 0.011419f
C17708 _328_/a_36_113# FILLER_0_11_101/a_484_472# 0.001826f
C17709 _074_ _163_ 0.446493f
C17710 FILLER_0_11_124/a_36_472# _135_ 0.110114f
C17711 _065_ trim_val\[3\] 1.235816f
C17712 _015_ FILLER_0_8_247/a_36_472# 0.005458f
C17713 net20 FILLER_0_6_239/a_36_472# 0.005138f
C17714 FILLER_0_18_177/a_1468_375# _139_ 0.001359f
C17715 FILLER_0_16_107/a_124_375# net14 0.004684f
C17716 net41 _445_/a_2560_156# 0.002221f
C17717 mask\[4\] FILLER_0_22_128/a_3172_472# 0.001484f
C17718 _093_ _438_/a_2665_112# 0.003293f
C17719 vdd output40/a_224_472# 0.079607f
C17720 FILLER_0_18_177/a_3260_375# _047_ 0.030543f
C17721 _114_ _225_/a_36_160# 0.003628f
C17722 _098_ _434_/a_1204_472# 0.006257f
C17723 _441_/a_1308_423# vdd 0.002837f
C17724 _441_/a_448_472# vss 0.025073f
C17725 _235_/a_67_603# vss 0.002019f
C17726 _444_/a_2560_156# net67 0.012781f
C17727 net53 _427_/a_2665_112# 0.042564f
C17728 net72 _452_/a_448_472# 0.001296f
C17729 _442_/a_2665_112# trim_mask\[3\] 0.019514f
C17730 _015_ _426_/a_448_472# 0.035938f
C17731 _394_/a_56_524# FILLER_0_15_59/a_484_472# 0.001033f
C17732 _394_/a_718_524# FILLER_0_15_59/a_572_375# 0.001447f
C17733 _181_ _184_ 0.022711f
C17734 output38/a_224_472# trim[0] 0.026911f
C17735 FILLER_0_15_228/a_124_375# vss 0.006435f
C17736 _019_ _138_ 0.003734f
C17737 FILLER_0_15_228/a_36_472# vdd 0.084606f
C17738 _066_ _385_/a_36_68# 0.001405f
C17739 net36 _137_ 0.048198f
C17740 _036_ _164_ 0.011115f
C17741 _115_ FILLER_0_9_105/a_124_375# 0.002316f
C17742 net27 _283_/a_36_472# 0.023243f
C17743 output31/a_224_472# FILLER_0_17_282/a_124_375# 0.002977f
C17744 _431_/a_1308_423# vdd 0.002397f
C17745 _431_/a_448_472# vss 0.005583f
C17746 _440_/a_1204_472# vss 0.007007f
C17747 _440_/a_2248_156# vdd -0.003421f
C17748 FILLER_0_19_142/a_36_472# vdd 0.107105f
C17749 FILLER_0_19_142/a_124_375# vss 0.032026f
C17750 _430_/a_448_472# _069_ 0.047845f
C17751 output29/a_224_472# net30 0.044542f
C17752 _439_/a_36_151# vss 0.032466f
C17753 _439_/a_448_472# vdd 0.006996f
C17754 net80 _434_/a_796_472# 0.039593f
C17755 _091_ FILLER_0_13_212/a_1468_375# 0.003576f
C17756 _157_ vss 0.039512f
C17757 FILLER_0_20_87/a_36_472# _438_/a_448_472# 0.004782f
C17758 _412_/a_36_151# net58 0.010226f
C17759 net34 _435_/a_2560_156# 0.002967f
C17760 _105_ _108_ 0.548284f
C17761 _063_ trim_val\[1\] 0.038045f
C17762 _086_ _062_ 0.066419f
C17763 FILLER_0_2_93/a_124_375# _441_/a_2665_112# 0.006271f
C17764 trim_mask\[2\] FILLER_0_2_93/a_36_472# 0.281054f
C17765 net54 _022_ 0.004106f
C17766 _432_/a_2665_112# net21 0.005773f
C17767 _098_ _437_/a_448_472# 0.050691f
C17768 _273_/a_36_68# FILLER_0_10_214/a_124_375# 0.003707f
C17769 FILLER_0_5_212/a_124_375# FILLER_0_5_206/a_124_375# 0.005439f
C17770 FILLER_0_21_142/a_484_472# _140_ 0.011035f
C17771 FILLER_0_7_104/a_1020_375# _131_ 0.016404f
C17772 FILLER_0_19_47/a_484_472# vdd 0.001133f
C17773 FILLER_0_19_47/a_36_472# vss 0.001559f
C17774 FILLER_0_5_181/a_124_375# net37 0.005396f
C17775 net36 _438_/a_1308_423# 0.012976f
C17776 _015_ FILLER_0_8_239/a_36_472# 0.002627f
C17777 _316_/a_692_472# vdd 0.001634f
C17778 cal_count\[3\] _062_ 0.004405f
C17779 _132_ FILLER_0_18_107/a_2812_375# 0.002706f
C17780 net79 _136_ 0.00111f
C17781 net39 vss 0.170972f
C17782 _053_ FILLER_0_7_104/a_484_472# 0.005353f
C17783 net50 FILLER_0_6_37/a_124_375# 0.003821f
C17784 mask\[5\] FILLER_0_20_177/a_1468_375# 0.013222f
C17785 FILLER_0_16_57/a_572_375# net72 0.012909f
C17786 _385_/a_36_68# net37 0.047762f
C17787 _449_/a_36_151# _174_ 0.002252f
C17788 net81 fanout82/a_36_113# 0.061162f
C17789 _077_ _251_/a_244_472# 0.002492f
C17790 FILLER_0_17_200/a_36_472# mask\[3\] 0.27914f
C17791 _303_/a_36_472# mask\[9\] 0.013976f
C17792 _010_ _108_ 0.002048f
C17793 _076_ _080_ 0.005433f
C17794 _104_ _008_ 0.135471f
C17795 FILLER_0_16_73/a_572_375# _040_ 0.014453f
C17796 net15 _440_/a_796_472# 0.005848f
C17797 mask\[0\] FILLER_0_12_196/a_124_375# 0.034009f
C17798 FILLER_0_9_142/a_124_375# _315_/a_36_68# 0.028077f
C17799 _079_ _078_ 0.03338f
C17800 _430_/a_2560_156# net36 0.00164f
C17801 output7/a_224_472# ctln[0] 0.081823f
C17802 _412_/a_2665_112# net1 0.063655f
C17803 FILLER_0_3_78/a_124_375# _168_ 0.009374f
C17804 _452_/a_36_151# net40 0.012138f
C17805 FILLER_0_9_28/a_1916_375# net16 0.001431f
C17806 net65 FILLER_0_3_212/a_124_375# 0.003807f
C17807 _207_/a_67_603# vdd 0.034688f
C17808 _444_/a_2248_156# FILLER_0_8_37/a_484_472# 0.013656f
C17809 _077_ _187_ 0.058967f
C17810 net79 _070_ 0.009715f
C17811 FILLER_0_7_146/a_124_375# _133_ 0.001577f
C17812 FILLER_0_22_86/a_484_472# net14 0.006746f
C17813 net79 FILLER_0_12_220/a_1380_472# 0.010583f
C17814 fanout77/a_36_113# net18 0.060158f
C17815 FILLER_0_18_2/a_2364_375# _452_/a_1353_112# 0.001068f
C17816 FILLER_0_18_2/a_3260_375# _452_/a_36_151# 0.001597f
C17817 FILLER_0_18_2/a_572_375# _452_/a_3129_107# 0.001073f
C17818 _435_/a_36_151# vdd 0.059103f
C17819 _132_ _354_/a_49_472# 0.034372f
C17820 FILLER_0_19_111/a_124_375# net14 0.001837f
C17821 trim[4] _054_ 0.005511f
C17822 _053_ _414_/a_2248_156# 0.013478f
C17823 net69 _160_ 0.077526f
C17824 _106_ ctlp[1] 0.002631f
C17825 _427_/a_1308_423# vss 0.030292f
C17826 FILLER_0_16_241/a_36_472# mask\[2\] 0.025337f
C17827 FILLER_0_7_72/a_932_472# vss 0.002763f
C17828 sample net59 0.001181f
C17829 _106_ _091_ 0.001188f
C17830 net63 net34 0.050865f
C17831 _161_ _055_ 0.078364f
C17832 vss FILLER_0_5_148/a_484_472# 0.009015f
C17833 FILLER_0_9_28/a_1468_375# vdd 0.009854f
C17834 _405_/a_255_603# cal_count\[2\] 0.001576f
C17835 vdd FILLER_0_21_60/a_124_375# 0.014029f
C17836 mask\[5\] FILLER_0_19_171/a_484_472# 0.007647f
C17837 ctln[1] FILLER_0_0_232/a_36_472# 0.005158f
C17838 _002_ FILLER_0_3_172/a_2724_472# 0.006713f
C17839 output34/a_224_472# _094_ 0.002719f
C17840 net41 _178_ 0.019945f
C17841 FILLER_0_24_130/a_36_472# _050_ 0.008605f
C17842 _427_/a_1308_423# net74 0.005627f
C17843 net76 vdd 1.272072f
C17844 output27/a_224_472# FILLER_0_8_263/a_36_472# 0.002002f
C17845 _164_ FILLER_0_6_37/a_36_472# 0.001049f
C17846 net56 net36 0.772486f
C17847 cal_itt\[1\] _084_ 0.495918f
C17848 _069_ _310_/a_49_472# 0.023925f
C17849 FILLER_0_12_28/a_124_375# net40 0.047331f
C17850 _072_ _176_ 0.298077f
C17851 FILLER_0_22_177/a_1468_375# net33 0.017455f
C17852 net25 _213_/a_67_603# 0.027452f
C17853 _072_ _306_/a_36_68# 0.042843f
C17854 _020_ _137_ 0.228674f
C17855 _161_ _311_/a_1212_473# 0.004138f
C17856 _111_ net55 0.002855f
C17857 _013_ net72 0.006579f
C17858 ctln[4] output12/a_224_472# 0.041517f
C17859 net69 _030_ 0.49547f
C17860 _105_ _092_ 0.006701f
C17861 FILLER_0_19_155/a_36_472# vss 0.004125f
C17862 FILLER_0_19_155/a_484_472# vdd 0.003341f
C17863 FILLER_0_17_72/a_124_375# _131_ 0.006224f
C17864 _442_/a_796_472# _031_ 0.013039f
C17865 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1380_472# 0.003468f
C17866 _187_ _453_/a_36_151# 0.001829f
C17867 _016_ FILLER_0_12_136/a_124_375# 0.008914f
C17868 _178_ _406_/a_36_159# 0.007052f
C17869 FILLER_0_5_72/a_572_375# net47 0.006974f
C17870 net14 FILLER_0_4_91/a_36_472# 0.005793f
C17871 FILLER_0_3_142/a_124_375# trim_mask\[4\] 0.002514f
C17872 _072_ _251_/a_1130_472# 0.004007f
C17873 _429_/a_2248_156# FILLER_0_15_212/a_1468_375# 0.001068f
C17874 net34 FILLER_0_22_128/a_3172_472# 0.003953f
C17875 FILLER_0_17_200/a_484_472# vdd 0.008335f
C17876 fanout75/a_36_113# _082_ 0.016843f
C17877 _173_ vdd 0.080629f
C17878 _162_ _056_ 0.018616f
C17879 FILLER_0_2_177/a_124_375# net22 0.001318f
C17880 cal_itt\[2\] _084_ 0.061303f
C17881 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_572_375# 0.001597f
C17882 _053_ _003_ 0.021223f
C17883 _074_ _073_ 0.040339f
C17884 net4 net9 0.008183f
C17885 FILLER_0_16_107/a_36_472# _040_ 0.015026f
C17886 mask\[0\] _429_/a_2560_156# 0.010913f
C17887 net79 _192_/a_67_603# 0.017688f
C17888 FILLER_0_4_107/a_1380_472# FILLER_0_2_111/a_1020_375# 0.001512f
C17889 trimb[0] net44 0.00246f
C17890 _413_/a_2248_156# FILLER_0_1_212/a_36_472# 0.035805f
C17891 _321_/a_3126_472# _124_ 0.001072f
C17892 net24 FILLER_0_22_86/a_1468_375# 0.008075f
C17893 output46/a_224_472# vdd 0.043652f
C17894 FILLER_0_7_59/a_572_375# vdd 0.005991f
C17895 FILLER_0_7_59/a_124_375# vss 0.002006f
C17896 fanout51/a_36_113# net15 0.001562f
C17897 net19 net33 0.254336f
C17898 ctln[1] net18 0.004646f
C17899 net16 _444_/a_448_472# 0.038803f
C17900 net81 FILLER_0_8_263/a_36_472# 0.007373f
C17901 net35 FILLER_0_22_128/a_2364_375# 0.012732f
C17902 output30/a_224_472# result[3] 0.019025f
C17903 _007_ vdd 0.129966f
C17904 FILLER_0_1_204/a_124_375# vdd 0.047704f
C17905 _000_ net58 0.00389f
C17906 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3260_375# 0.086635f
C17907 _114_ FILLER_0_12_136/a_1468_375# 0.006974f
C17908 _009_ FILLER_0_23_290/a_124_375# 0.002666f
C17909 result[0] result[1] 0.06045f
C17910 _039_ net40 0.036781f
C17911 net68 FILLER_0_6_47/a_124_375# 0.002491f
C17912 _256_/a_2960_68# _076_ 0.001292f
C17913 _323_/a_36_113# _128_ 0.014377f
C17914 FILLER_0_9_105/a_572_375# FILLER_0_10_107/a_484_472# 0.001543f
C17915 vdd net14 2.23064f
C17916 _013_ _424_/a_36_151# 0.012928f
C17917 net58 _425_/a_2248_156# 0.051603f
C17918 FILLER_0_9_72/a_124_375# _439_/a_36_151# 0.059049f
C17919 FILLER_0_7_195/a_124_375# _163_ 0.001308f
C17920 ctlp[2] _422_/a_36_151# 0.068086f
C17921 trim_mask\[1\] FILLER_0_6_47/a_1020_375# 0.007169f
C17922 _365_/a_244_472# net14 0.001257f
C17923 net67 _190_/a_36_160# 0.023989f
C17924 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1468_375# 0.086742f
C17925 net60 _006_ 0.006254f
C17926 output15/a_224_472# _164_ 0.031363f
C17927 _061_ state\[1\] 0.02716f
C17928 net38 net6 0.071232f
C17929 FILLER_0_22_128/a_2812_375# vss 0.004347f
C17930 FILLER_0_22_128/a_3260_375# vdd 0.005207f
C17931 _165_ _160_ 0.008705f
C17932 FILLER_0_7_72/a_2364_375# net14 0.005919f
C17933 _444_/a_36_151# vdd 0.071209f
C17934 _053_ FILLER_0_4_213/a_572_375# 0.003451f
C17935 _161_ _058_ 0.101968f
C17936 _415_/a_2665_112# net18 0.004988f
C17937 _326_/a_36_160# _131_ 0.023688f
C17938 _116_ _248_/a_36_68# 0.007314f
C17939 net50 FILLER_0_8_37/a_484_472# 0.003311f
C17940 _421_/a_36_151# _419_/a_448_472# 0.002098f
C17941 ctlp[0] vss 0.005302f
C17942 net55 _451_/a_2225_156# 0.031243f
C17943 fanout52/a_36_160# trim_mask\[4\] 0.014356f
C17944 _230_/a_244_68# _056_ 0.001844f
C17945 _447_/a_2665_112# _168_ 0.001107f
C17946 _016_ _043_ 0.030341f
C17947 net65 _413_/a_1308_423# 0.022097f
C17948 net55 fanout55/a_36_160# 0.028425f
C17949 _052_ FILLER_0_19_28/a_572_375# 0.011078f
C17950 net27 FILLER_0_9_270/a_572_375# 0.043797f
C17951 FILLER_0_10_78/a_124_375# vss 0.006775f
C17952 FILLER_0_10_78/a_572_375# vdd -0.014642f
C17953 _408_/a_56_524# _043_ 0.10151f
C17954 _428_/a_1000_472# _017_ 0.012268f
C17955 _085_ _090_ 0.001012f
C17956 _116_ _060_ 0.020653f
C17957 FILLER_0_21_28/a_2812_375# _424_/a_36_151# 0.059049f
C17958 net15 net51 0.191328f
C17959 FILLER_0_16_107/a_572_375# net36 0.001706f
C17960 _132_ _144_ 0.185339f
C17961 net80 _138_ 0.002053f
C17962 FILLER_0_16_57/a_932_472# net15 0.037807f
C17963 fanout51/a_36_113# net51 0.013081f
C17964 net72 _179_ 0.083699f
C17965 net76 net2 0.039533f
C17966 net63 FILLER_0_18_177/a_1468_375# 0.020059f
C17967 _067_ _450_/a_2225_156# 0.002584f
C17968 net42 vss 0.017902f
C17969 state\[0\] _323_/a_36_113# 0.016796f
C17970 FILLER_0_5_54/a_1020_375# net47 0.005159f
C17971 _408_/a_56_524# _185_ 0.002484f
C17972 _071_ _055_ 0.002641f
C17973 FILLER_0_9_72/a_36_472# vss 0.0392f
C17974 FILLER_0_9_72/a_484_472# vdd 0.005654f
C17975 net82 FILLER_0_3_172/a_2812_375# 0.010439f
C17976 _171_ FILLER_0_10_94/a_484_472# 0.001446f
C17977 output14/a_224_472# _442_/a_448_472# 0.008149f
C17978 _077_ net67 0.073924f
C17979 _273_/a_36_68# _055_ 0.081216f
C17980 _414_/a_36_151# net21 0.007791f
C17981 net55 FILLER_0_13_72/a_36_472# 0.002172f
C17982 _093_ FILLER_0_17_72/a_2724_472# 0.02416f
C17983 FILLER_0_2_111/a_572_375# _160_ 0.001049f
C17984 _083_ vdd 0.157549f
C17985 _359_/a_36_488# vss 0.002427f
C17986 _078_ vss 0.367953f
C17987 _137_ FILLER_0_16_154/a_1468_375# 0.014214f
C17988 _074_ net1 0.128466f
C17989 _028_ FILLER_0_7_72/a_1916_375# 0.003862f
C17990 net64 FILLER_0_11_282/a_124_375# 0.023042f
C17991 _081_ FILLER_0_5_164/a_484_472# 0.001105f
C17992 _095_ net36 0.127549f
C17993 net43 FILLER_0_20_15/a_572_375# 0.003924f
C17994 net18 _417_/a_1204_472# 0.01349f
C17995 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_36_472# 0.002765f
C17996 ctln[3] ctln[1] 0.926618f
C17997 net75 _426_/a_1204_472# 0.001592f
C17998 FILLER_0_16_89/a_484_472# _136_ 0.032722f
C17999 _122_ FILLER_0_5_181/a_124_375# 0.001352f
C18000 _050_ _352_/a_49_472# 0.005393f
C18001 FILLER_0_17_200/a_572_375# vss 0.017327f
C18002 FILLER_0_15_282/a_36_472# output30/a_224_472# 0.001711f
C18003 _359_/a_36_488# net74 0.037211f
C18004 _308_/a_124_24# vdd 0.011014f
C18005 _018_ net22 0.141743f
C18006 _098_ FILLER_0_15_212/a_484_472# 0.00912f
C18007 FILLER_0_12_136/a_1468_375# _126_ 0.012732f
C18008 _056_ _373_/a_244_68# 0.00229f
C18009 _053_ FILLER_0_7_72/a_124_375# 0.014569f
C18010 _153_ _365_/a_36_68# 0.056496f
C18011 net35 _050_ 0.28822f
C18012 net38 FILLER_0_15_10/a_124_375# 0.047331f
C18013 net10 vss 0.324553f
C18014 _122_ _385_/a_36_68# 0.003549f
C18015 _035_ _034_ 1.26804f
C18016 net81 _018_ 0.081888f
C18017 _176_ FILLER_0_10_94/a_484_472# 0.009483f
C18018 _140_ FILLER_0_22_128/a_36_472# 0.050084f
C18019 FILLER_0_17_72/a_484_472# net36 0.001629f
C18020 FILLER_0_10_214/a_36_472# _055_ 0.027657f
C18021 net52 FILLER_0_11_78/a_124_375# 0.006273f
C18022 _132_ FILLER_0_14_107/a_1020_375# 0.029702f
C18023 _372_/a_170_472# _059_ 0.033956f
C18024 ctlp[1] FILLER_0_21_286/a_484_472# 0.045536f
C18025 output27/a_224_472# fanout65/a_36_113# 0.011564f
C18026 FILLER_0_5_136/a_124_375# vdd 0.035814f
C18027 _004_ result[1] 0.005653f
C18028 FILLER_0_20_169/a_124_375# mask\[6\] 0.001178f
C18029 mask\[5\] mask\[6\] 0.140269f
C18030 mask\[4\] _137_ 0.086066f
C18031 _069_ mask\[2\] 0.032781f
C18032 net73 FILLER_0_17_142/a_484_472# 0.001122f
C18033 _095_ FILLER_0_14_123/a_124_375# 0.014486f
C18034 FILLER_0_21_28/a_2724_472# vdd 0.001342f
C18035 net69 _156_ 0.008057f
C18036 FILLER_0_6_90/a_572_375# vdd 0.028324f
C18037 net29 mask\[2\] 0.122202f
C18038 output29/a_224_472# _045_ 0.002303f
C18039 _119_ _319_/a_234_472# 0.004559f
C18040 FILLER_0_16_89/a_1468_375# FILLER_0_17_72/a_3260_375# 0.026339f
C18041 FILLER_0_16_89/a_484_472# FILLER_0_17_72/a_2364_375# 0.001723f
C18042 mask\[4\] FILLER_0_19_171/a_36_472# 0.001776f
C18043 output15/a_224_472# trim_val\[3\] 0.042209f
C18044 output9/a_224_472# FILLER_0_1_266/a_484_472# 0.0323f
C18045 net47 _170_ 0.010131f
C18046 _117_ _060_ 0.149558f
C18047 _430_/a_448_472# net22 0.036303f
C18048 _415_/a_2665_112# net62 0.003644f
C18049 _320_/a_36_472# _113_ 0.030365f
C18050 _093_ FILLER_0_19_142/a_36_472# 0.002415f
C18051 net63 FILLER_0_15_212/a_484_472# 0.059367f
C18052 net75 net81 0.420021f
C18053 FILLER_0_11_282/a_36_472# vdd 0.106843f
C18054 FILLER_0_11_282/a_124_375# vss 0.005415f
C18055 _020_ FILLER_0_18_107/a_2276_472# 0.004069f
C18056 FILLER_0_7_72/a_1916_375# FILLER_0_6_90/a_36_472# 0.001684f
C18057 _053_ _162_ 0.00209f
C18058 FILLER_0_18_2/a_2724_472# net17 0.017841f
C18059 FILLER_0_4_107/a_36_472# _157_ 0.005289f
C18060 _374_/a_36_68# FILLER_0_8_156/a_484_472# 0.002559f
C18061 _173_ cal_count\[0\] 0.517178f
C18062 _008_ mask\[2\] 0.003475f
C18063 _115_ FILLER_0_10_107/a_36_472# 0.016715f
C18064 _163_ FILLER_0_5_148/a_572_375# 0.001706f
C18065 FILLER_0_19_55/a_36_472# _052_ 0.019665f
C18066 _430_/a_448_472# net81 0.003775f
C18067 net4 _084_ 0.029194f
C18068 _445_/a_36_151# net17 0.009838f
C18069 result[5] net18 0.173673f
C18070 FILLER_0_15_116/a_124_375# net70 0.02416f
C18071 fanout49/a_36_160# net49 0.032999f
C18072 FILLER_0_17_56/a_36_472# FILLER_0_18_53/a_484_472# 0.026657f
C18073 _181_ _402_/a_718_527# 0.00461f
C18074 calibrate FILLER_0_7_233/a_36_472# 0.013262f
C18075 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_124_375# 0.009654f
C18076 FILLER_0_19_125/a_36_472# FILLER_0_18_107/a_1916_375# 0.001684f
C18077 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_484_472# 0.013276f
C18078 mask\[9\] FILLER_0_18_76/a_484_472# 0.002672f
C18079 FILLER_0_14_99/a_124_375# _451_/a_36_151# 0.001441f
C18080 valid calibrate 0.002363f
C18081 FILLER_0_10_37/a_124_375# _453_/a_36_151# 0.017882f
C18082 trim_val\[4\] FILLER_0_3_172/a_484_472# 0.002633f
C18083 trim_val\[4\] _386_/a_848_380# 0.007605f
C18084 trim_mask\[1\] FILLER_0_6_79/a_36_472# 0.006265f
C18085 FILLER_0_7_72/a_572_375# net52 0.022624f
C18086 mask\[9\] _423_/a_2665_112# 0.001735f
C18087 vdd _433_/a_2248_156# 0.008127f
C18088 FILLER_0_17_72/a_932_472# FILLER_0_18_76/a_484_472# 0.05841f
C18089 FILLER_0_7_162/a_124_375# net37 0.011644f
C18090 net56 FILLER_0_18_139/a_1380_472# 0.048069f
C18091 _428_/a_448_472# FILLER_0_14_107/a_932_472# 0.007f
C18092 _091_ FILLER_0_18_209/a_572_375# 0.001343f
C18093 _334_/a_36_160# vss 0.002713f
C18094 net64 net36 0.037523f
C18095 FILLER_0_16_89/a_932_472# net53 0.012534f
C18096 fanout53/a_36_160# FILLER_0_16_154/a_932_472# 0.001426f
C18097 net52 FILLER_0_2_93/a_572_375# 0.007787f
C18098 _147_ _207_/a_67_603# 0.001123f
C18099 comp net17 0.02802f
C18100 net36 mask\[1\] 0.28584f
C18101 _147_ _435_/a_36_151# 0.003096f
C18102 _188_ _042_ 0.015684f
C18103 net55 _424_/a_1308_423# 0.00168f
C18104 _239_/a_36_160# vss 0.001596f
C18105 _246_/a_36_68# _055_ 0.028938f
C18106 mask\[3\] FILLER_0_18_177/a_2276_472# 0.01204f
C18107 FILLER_0_7_233/a_124_375# FILLER_0_6_231/a_484_472# 0.001684f
C18108 _187_ _095_ 0.00765f
C18109 _141_ _140_ 0.131685f
C18110 _415_/a_2560_156# net58 0.002325f
C18111 FILLER_0_12_20/a_484_472# vss 0.001783f
C18112 _417_/a_1204_472# net62 0.001941f
C18113 net5 clk 0.042578f
C18114 _058_ FILLER_0_8_156/a_572_375# 0.007692f
C18115 _310_/a_49_472# _090_ 0.059827f
C18116 net78 _007_ 0.054904f
C18117 net60 _007_ 0.025806f
C18118 FILLER_0_17_218/a_124_375# vdd 0.00593f
C18119 mask\[8\] net25 0.035648f
C18120 _327_/a_36_472# _127_ 0.002934f
C18121 FILLER_0_8_263/a_124_375# vdd 0.032664f
C18122 _070_ trim_mask\[0\] 0.006144f
C18123 _326_/a_36_160# _077_ 0.00419f
C18124 output46/a_224_472# FILLER_0_21_28/a_36_472# 0.010684f
C18125 mask\[5\] FILLER_0_19_187/a_572_375# 0.005529f
C18126 _072_ FILLER_0_12_220/a_484_472# 0.028355f
C18127 FILLER_0_20_31/a_124_375# vdd 0.04619f
C18128 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_36_472# 0.086635f
C18129 _414_/a_448_472# _074_ 0.008725f
C18130 mask\[4\] net56 0.006006f
C18131 _423_/a_36_151# net40 0.004045f
C18132 ctlp[7] _050_ 0.153673f
C18133 _175_ _043_ 0.001037f
C18134 net24 net71 0.015101f
C18135 FILLER_0_20_87/a_36_472# vdd 0.006784f
C18136 FILLER_0_20_87/a_124_375# vss 0.00279f
C18137 _363_/a_36_68# _028_ 0.015609f
C18138 net25 vss 0.528437f
C18139 FILLER_0_9_223/a_36_472# _055_ 0.014713f
C18140 _091_ FILLER_0_19_171/a_124_375# 0.028992f
C18141 net81 _426_/a_36_151# 0.060652f
C18142 _440_/a_448_472# _160_ 0.004748f
C18143 _028_ FILLER_0_6_47/a_2724_472# 0.023218f
C18144 _429_/a_2248_156# FILLER_0_15_228/a_124_375# 0.030666f
C18145 net36 vss 1.788802f
C18146 FILLER_0_0_198/a_124_375# net59 0.004565f
C18147 _079_ _263_/a_224_472# 0.002505f
C18148 _098_ _146_ 0.004276f
C18149 _119_ _359_/a_36_488# 0.003263f
C18150 net38 _444_/a_1000_472# 0.027886f
C18151 _043_ net21 0.033824f
C18152 FILLER_0_19_28/a_484_472# vdd 0.010504f
C18153 _214_/a_36_160# FILLER_0_23_88/a_36_472# 0.006647f
C18154 FILLER_0_3_204/a_124_375# net59 0.007104f
C18155 _276_/a_36_160# mask\[4\] 0.025336f
C18156 FILLER_0_4_91/a_484_472# _160_ 0.009925f
C18157 _050_ FILLER_0_22_128/a_1468_375# 0.001661f
C18158 output35/a_224_472# _435_/a_2248_156# 0.019736f
C18159 _093_ FILLER_0_19_155/a_484_472# 0.001236f
C18160 FILLER_0_15_2/a_484_472# vss 0.003267f
C18161 FILLER_0_4_123/a_36_472# _154_ 0.001043f
C18162 _269_/a_36_472# _078_ 0.033601f
C18163 FILLER_0_9_223/a_484_472# net4 0.047334f
C18164 _115_ _322_/a_848_380# 0.011372f
C18165 _165_ net67 0.045827f
C18166 _012_ FILLER_0_23_44/a_1468_375# 0.002827f
C18167 _064_ net40 0.141744f
C18168 _053_ FILLER_0_6_47/a_932_472# 0.011457f
C18169 _436_/a_1000_472# net35 0.009213f
C18170 net74 net36 0.012494f
C18171 FILLER_0_16_89/a_1020_375# vdd 0.007416f
C18172 net64 FILLER_0_9_270/a_36_472# 0.014971f
C18173 _140_ _433_/a_2665_112# 0.001108f
C18174 ctln[4] vss 0.244634f
C18175 _002_ FILLER_0_4_185/a_124_375# 0.013895f
C18176 _417_/a_2248_156# net30 0.048831f
C18177 _081_ _152_ 0.172002f
C18178 _093_ FILLER_0_17_200/a_484_472# 0.007492f
C18179 net16 _034_ 0.096088f
C18180 cal_count\[3\] _188_ 0.048745f
C18181 _086_ _153_ 0.017325f
C18182 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_484_472# 0.013277f
C18183 result[5] net62 0.041722f
C18184 _430_/a_1000_472# _091_ 0.025041f
C18185 net76 FILLER_0_5_206/a_124_375# 0.006974f
C18186 _176_ FILLER_0_11_78/a_36_472# 0.003603f
C18187 FILLER_0_15_142/a_124_375# fanout73/a_36_113# 0.00146f
C18188 net66 _440_/a_796_472# 0.002718f
C18189 net49 _440_/a_36_151# 0.021133f
C18190 net7 output16/a_224_472# 0.001321f
C18191 output42/a_224_472# net38 0.066219f
C18192 net19 net18 0.028285f
C18193 FILLER_0_7_146/a_124_375# net37 0.005315f
C18194 net35 _423_/a_2665_112# 0.019085f
C18195 net18 _418_/a_1204_472# 0.01349f
C18196 ctln[1] FILLER_0_3_221/a_124_375# 0.001391f
C18197 output8/a_224_472# FILLER_0_3_221/a_484_472# 0.001699f
C18198 _394_/a_728_93# net15 0.085551f
C18199 net65 _448_/a_36_151# 0.001983f
C18200 output10/a_224_472# vdd 0.107357f
C18201 net36 cal_count\[1\] 0.011481f
C18202 net68 _440_/a_36_151# 0.080854f
C18203 FILLER_0_5_54/a_124_375# FILLER_0_3_54/a_36_472# 0.001512f
C18204 net32 _419_/a_36_151# 0.006506f
C18205 _436_/a_2248_156# vdd 0.011151f
C18206 FILLER_0_14_123/a_36_472# vdd 0.088525f
C18207 FILLER_0_14_123/a_124_375# vss 0.004985f
C18208 fanout81/a_36_160# net81 0.025745f
C18209 _415_/a_796_472# net27 0.004502f
C18210 _415_/a_2248_156# output27/a_224_472# 0.001506f
C18211 ctlp[1] _420_/a_796_472# 0.001468f
C18212 mask\[5\] net35 0.003646f
C18213 _095_ _225_/a_36_160# 0.001084f
C18214 net65 output37/a_224_472# 0.096416f
C18215 vss _160_ 1.119894f
C18216 _430_/a_2248_156# mask\[2\] 0.009336f
C18217 _062_ _227_/a_36_160# 0.015411f
C18218 _072_ _250_/a_36_68# 0.007337f
C18219 FILLER_0_21_142/a_484_472# _098_ 0.001158f
C18220 net50 FILLER_0_3_54/a_124_375# 0.00189f
C18221 _154_ _153_ 0.719561f
C18222 _174_ _401_/a_244_472# 0.001957f
C18223 _423_/a_2560_156# vss 0.002241f
C18224 net54 FILLER_0_19_111/a_484_472# 0.00105f
C18225 net72 FILLER_0_17_56/a_572_375# 0.004473f
C18226 FILLER_0_2_101/a_36_472# net14 0.051153f
C18227 _412_/a_36_151# net9 0.005212f
C18228 FILLER_0_5_54/a_124_375# FILLER_0_6_47/a_932_472# 0.001597f
C18229 _255_/a_224_552# cal_itt\[3\] 0.003266f
C18230 net65 net5 0.004409f
C18231 _077_ _059_ 0.020736f
C18232 _093_ net14 0.11038f
C18233 trim_val\[4\] FILLER_0_2_165/a_36_472# 0.007765f
C18234 net20 _291_/a_36_160# 0.002375f
C18235 _116_ vss 0.235141f
C18236 FILLER_0_16_73/a_124_375# FILLER_0_17_72/a_124_375# 0.026339f
C18237 _341_/a_49_472# _141_ 0.006222f
C18238 _136_ FILLER_0_16_154/a_1380_472# 0.006517f
C18239 net74 _160_ 0.165289f
C18240 FILLER_0_20_169/a_36_472# vss 0.005112f
C18241 net39 _445_/a_36_151# 0.006056f
C18242 FILLER_0_1_266/a_36_472# net8 0.0138f
C18243 FILLER_0_5_117/a_36_472# _086_ 0.042352f
C18244 _008_ _418_/a_1000_472# 0.01006f
C18245 net16 _445_/a_2248_156# 0.003321f
C18246 net73 FILLER_0_18_139/a_484_472# 0.00131f
C18247 FILLER_0_11_101/a_124_375# _070_ 0.052406f
C18248 FILLER_0_12_136/a_1468_375# FILLER_0_13_142/a_932_472# 0.001684f
C18249 FILLER_0_9_270/a_36_472# vss 0.001642f
C18250 FILLER_0_9_270/a_484_472# vdd 0.006354f
C18251 FILLER_0_12_220/a_36_472# _090_ 0.023446f
C18252 net55 FILLER_0_13_80/a_36_472# 0.016536f
C18253 _004_ _094_ 0.213913f
C18254 net63 _275_/a_224_472# 0.002538f
C18255 _030_ vss 0.117034f
C18256 net49 vdd 0.872948f
C18257 FILLER_0_22_128/a_3172_472# _146_ 0.008065f
C18258 ctlp[1] _421_/a_1204_472# 0.003759f
C18259 _427_/a_2665_112# net23 0.032729f
C18260 state\[2\] FILLER_0_13_142/a_124_375# 0.010494f
C18261 net53 FILLER_0_13_142/a_1020_375# 0.001597f
C18262 _442_/a_2248_156# vdd 0.038702f
C18263 net72 _041_ 0.467856f
C18264 net15 FILLER_0_18_76/a_36_472# 0.001341f
C18265 _446_/a_1204_472# net17 0.003628f
C18266 net68 vdd 1.026897f
C18267 output20/a_224_472# _104_ 0.019295f
C18268 _316_/a_848_380# _123_ 0.0018f
C18269 _106_ _199_/a_36_160# 0.003376f
C18270 FILLER_0_4_144/a_124_375# _059_ 0.031451f
C18271 _076_ FILLER_0_8_239/a_124_375# 0.007237f
C18272 net15 _423_/a_2248_156# 0.048449f
C18273 _020_ vss 0.008954f
C18274 net72 _181_ 0.004503f
C18275 FILLER_0_9_28/a_484_472# net40 0.020293f
C18276 FILLER_0_5_117/a_36_472# _154_ 0.005034f
C18277 _424_/a_2248_156# FILLER_0_21_60/a_572_375# 0.030666f
C18278 _424_/a_2665_112# FILLER_0_21_60/a_124_375# 0.010688f
C18279 _070_ _081_ 0.00804f
C18280 FILLER_0_20_193/a_36_472# FILLER_0_19_187/a_572_375# 0.001543f
C18281 FILLER_0_15_290/a_36_472# result[3] 0.014709f
C18282 net4 calibrate 0.04302f
C18283 _187_ vss 0.080956f
C18284 _293_/a_36_472# output34/a_224_472# 0.001888f
C18285 _404_/a_36_472# _179_ 0.00141f
C18286 _086_ _321_/a_3662_472# 0.002598f
C18287 net73 FILLER_0_18_107/a_1020_375# 0.04487f
C18288 FILLER_0_3_54/a_36_472# _164_ 0.012512f
C18289 trim_val\[3\] FILLER_0_2_93/a_124_375# 0.001032f
C18290 _408_/a_728_93# net17 0.005494f
C18291 _077_ _453_/a_2248_156# 0.013877f
C18292 _131_ _134_ 0.887647f
C18293 _430_/a_36_151# vdd 0.112575f
C18294 _425_/a_796_472# vdd 0.002206f
C18295 vss FILLER_0_3_212/a_124_375# 0.009048f
C18296 vdd FILLER_0_3_212/a_36_472# 0.110132f
C18297 ctln[3] net19 0.003077f
C18298 mask\[7\] _435_/a_2248_156# 0.026974f
C18299 net15 net66 0.006618f
C18300 FILLER_0_4_177/a_124_375# _386_/a_848_380# 0.001277f
C18301 _056_ _055_ 0.155993f
C18302 net65 FILLER_0_1_266/a_572_375# 0.002969f
C18303 FILLER_0_5_117/a_124_375# _163_ 0.003096f
C18304 fanout56/a_36_113# _098_ 0.019463f
C18305 _070_ FILLER_0_10_94/a_572_375# 0.009837f
C18306 _164_ FILLER_0_6_47/a_932_472# 0.004272f
C18307 cal_count\[3\] FILLER_0_12_196/a_36_472# 0.079338f
C18308 _058_ net23 0.075446f
C18309 _114_ _134_ 0.015298f
C18310 fanout78/a_36_113# net18 0.001419f
C18311 fanout60/a_36_160# net18 0.004124f
C18312 FILLER_0_5_128/a_484_472# _160_ 0.003335f
C18313 net19 net62 0.352148f
C18314 _185_ _402_/a_1296_93# 0.001714f
C18315 _115_ _124_ 0.045023f
C18316 net45 net43 0.131763f
C18317 _315_/a_36_68# net23 0.030384f
C18318 _117_ vss 0.048946f
C18319 _333_/a_36_160# vdd 0.107883f
C18320 FILLER_0_4_107/a_484_472# _153_ 0.026082f
C18321 FILLER_0_4_107/a_1380_472# _154_ 0.005297f
C18322 _420_/a_36_151# FILLER_0_23_282/a_484_472# 0.001723f
C18323 _320_/a_36_472# vdd 0.086964f
C18324 _436_/a_2665_112# FILLER_0_22_128/a_124_375# 0.004834f
C18325 _436_/a_2248_156# FILLER_0_22_128/a_572_375# 0.006739f
C18326 _208_/a_36_160# vdd 0.014709f
C18327 mask\[5\] FILLER_0_18_177/a_2276_472# 0.001063f
C18328 FILLER_0_7_162/a_36_472# calibrate 0.014431f
C18329 _415_/a_448_472# _004_ 0.044374f
C18330 _408_/a_2215_68# _186_ 0.001205f
C18331 _026_ FILLER_0_20_87/a_124_375# 0.031902f
C18332 _072_ _162_ 0.090175f
C18333 net32 _421_/a_2560_156# 0.049213f
C18334 ctln[5] _037_ 0.19244f
C18335 _053_ FILLER_0_6_177/a_484_472# 0.015994f
C18336 _431_/a_36_151# FILLER_0_18_139/a_36_472# 0.002529f
C18337 net16 FILLER_0_6_37/a_124_375# 0.010358f
C18338 output28/a_224_472# net79 0.04262f
C18339 net41 net38 0.059214f
C18340 _449_/a_36_151# _038_ 0.019666f
C18341 FILLER_0_15_72/a_484_472# _451_/a_3129_107# 0.005866f
C18342 mask\[2\] net22 0.034216f
C18343 _414_/a_36_151# FILLER_0_7_195/a_36_472# 0.001723f
C18344 output45/a_224_472# vss 0.00543f
C18345 FILLER_0_16_57/a_572_375# _176_ 0.006422f
C18346 _267_/a_36_472# state\[1\] 0.001647f
C18347 result[6] vss 0.310169f
C18348 _143_ _091_ 0.007204f
C18349 _340_/a_36_160# mask\[6\] 0.010151f
C18350 _434_/a_1000_472# mask\[6\] 0.021582f
C18351 mask\[4\] FILLER_0_19_187/a_124_375# 0.006236f
C18352 FILLER_0_17_72/a_1916_375# _136_ 0.009573f
C18353 net15 _067_ 0.042278f
C18354 net81 mask\[2\] 0.002083f
C18355 _374_/a_36_68# _061_ 0.026111f
C18356 net79 _416_/a_796_472# 0.01137f
C18357 net36 _097_ 0.022089f
C18358 FILLER_0_8_247/a_1020_375# vdd -0.002559f
C18359 _421_/a_36_151# vss 0.021759f
C18360 _421_/a_448_472# vdd 0.030898f
C18361 net23 FILLER_0_22_128/a_1380_472# 0.0019f
C18362 output43/a_224_472# vdd -0.032713f
C18363 output12/a_224_472# _448_/a_36_151# 0.069748f
C18364 _277_/a_36_160# _094_ 0.007538f
C18365 FILLER_0_12_220/a_932_472# _070_ 0.001282f
C18366 _225_/a_36_160# vss 0.003244f
C18367 FILLER_0_20_193/a_484_472# vss 0.002439f
C18368 _091_ _136_ 0.075998f
C18369 FILLER_0_16_73/a_484_472# _175_ 0.036868f
C18370 _446_/a_448_472# net40 0.05302f
C18371 fanout54/a_36_160# _145_ 0.009257f
C18372 FILLER_0_17_72/a_3172_472# _131_ 0.003717f
C18373 _074_ _375_/a_1388_497# 0.005488f
C18374 _119_ _160_ 0.037232f
C18375 _281_/a_234_472# _098_ 0.003724f
C18376 _128_ _085_ 0.004532f
C18377 FILLER_0_5_198/a_484_472# net59 0.059394f
C18378 _210_/a_67_603# vdd 0.028101f
C18379 FILLER_0_4_91/a_484_472# _156_ 0.009828f
C18380 FILLER_0_17_104/a_1468_375# FILLER_0_16_115/a_124_375# 0.026339f
C18381 net53 _136_ 0.099584f
C18382 FILLER_0_18_139/a_1380_472# vss 0.009272f
C18383 net18 _193_/a_36_160# 0.114176f
C18384 net65 FILLER_0_3_172/a_2812_375# 0.003745f
C18385 net63 _435_/a_448_472# 0.009878f
C18386 output9/a_224_472# net59 0.051763f
C18387 FILLER_0_5_72/a_1468_375# _440_/a_2248_156# 0.030666f
C18388 FILLER_0_5_72/a_1020_375# _440_/a_2665_112# 0.010688f
C18389 FILLER_0_16_154/a_1468_375# vss 0.002071f
C18390 FILLER_0_16_154/a_36_472# vdd 0.00225f
C18391 _412_/a_796_472# cal_itt\[1\] 0.004226f
C18392 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_36_472# 0.086635f
C18393 _091_ _070_ 0.162632f
C18394 _056_ _058_ 0.988919f
C18395 FILLER_0_12_136/a_484_472# _076_ 0.001683f
C18396 fanout70/a_36_113# net70 0.073707f
C18397 net19 _420_/a_1000_472# 0.006558f
C18398 output9/a_224_472# net4 0.042449f
C18399 mask\[7\] FILLER_0_22_128/a_2276_472# 0.004398f
C18400 net44 FILLER_0_8_2/a_124_375# 0.083677f
C18401 net19 _109_ 0.005991f
C18402 _052_ FILLER_0_17_38/a_484_472# 0.001368f
C18403 FILLER_0_4_185/a_124_375# net76 0.053929f
C18404 net20 _073_ 0.437482f
C18405 FILLER_0_21_125/a_124_375# _140_ 0.031374f
C18406 _093_ FILLER_0_17_218/a_124_375# 0.003338f
C18407 FILLER_0_7_104/a_1468_375# vdd 0.026224f
C18408 mask\[0\] _138_ 0.22533f
C18409 mask\[5\] FILLER_0_21_206/a_36_472# 0.019416f
C18410 fanout78/a_36_113# net62 0.014177f
C18411 fanout60/a_36_160# net62 0.049222f
C18412 _068_ net47 0.001491f
C18413 FILLER_0_13_290/a_36_472# output30/a_224_472# 0.0323f
C18414 net20 _429_/a_2560_156# 0.002069f
C18415 FILLER_0_7_146/a_36_472# calibrate 0.060587f
C18416 _436_/a_1308_423# _050_ 0.022688f
C18417 vss _156_ 0.089339f
C18418 FILLER_0_18_107/a_2364_375# vdd 0.017472f
C18419 _434_/a_796_472# _023_ 0.002118f
C18420 _106_ net33 0.001049f
C18421 _413_/a_796_472# vdd 0.001569f
C18422 _365_/a_692_472# _156_ 0.001127f
C18423 net41 _233_/a_36_160# 0.053625f
C18424 _346_/a_49_472# _141_ 0.104653f
C18425 result[4] net20 0.001673f
C18426 net52 net55 0.016401f
C18427 _005_ _192_/a_67_603# 0.013886f
C18428 net54 FILLER_0_22_128/a_1916_375# 0.001933f
C18429 mask\[4\] vss 0.426009f
C18430 _448_/a_36_151# net12 0.133216f
C18431 _448_/a_1308_423# net22 0.045644f
C18432 FILLER_0_18_139/a_124_375# _145_ 0.00346f
C18433 _432_/a_2665_112# mask\[3\] 0.011428f
C18434 _108_ _107_ 0.018045f
C18435 net57 net14 0.05113f
C18436 _141_ FILLER_0_17_161/a_124_375# 0.040332f
C18437 net67 vss 0.435869f
C18438 _421_/a_2248_156# net19 0.016721f
C18439 fanout82/a_36_113# net82 0.003741f
C18440 FILLER_0_9_28/a_3172_472# net51 0.047897f
C18441 _010_ _419_/a_36_151# 0.002099f
C18442 _410_/a_36_68# _188_ 0.007731f
C18443 FILLER_0_24_274/a_484_472# vdd 0.004641f
C18444 FILLER_0_24_274/a_36_472# vss 0.001013f
C18445 output39/a_224_472# _054_ 0.002121f
C18446 _414_/a_1000_472# vdd 0.002568f
C18447 net39 _221_/a_36_160# 0.059979f
C18448 _422_/a_448_472# net19 0.003382f
C18449 net69 _168_ 0.035976f
C18450 _062_ net21 0.025648f
C18451 trim_mask\[1\] _154_ 0.004835f
C18452 FILLER_0_5_164/a_572_375# net37 0.014025f
C18453 FILLER_0_19_47/a_124_375# net26 0.008432f
C18454 ctln[3] cal_itt\[0\] 0.002081f
C18455 _077_ _134_ 0.043815f
C18456 _132_ _148_ 0.002873f
C18457 _077_ net48 0.142015f
C18458 _025_ FILLER_0_22_107/a_572_375# 0.090334f
C18459 _148_ FILLER_0_22_107/a_484_472# 0.004761f
C18460 _134_ FILLER_0_10_107/a_124_375# 0.009573f
C18461 net55 _216_/a_67_603# 0.071821f
C18462 _093_ FILLER_0_16_89/a_1020_375# 0.004133f
C18463 output13/a_224_472# net59 0.007733f
C18464 _415_/a_1204_472# vdd 0.00108f
C18465 net41 net55 0.033821f
C18466 FILLER_0_10_37/a_124_375# vss 0.006228f
C18467 FILLER_0_10_37/a_36_472# vdd 0.141896f
C18468 _408_/a_1936_472# vdd 0.022538f
C18469 _092_ FILLER_0_17_218/a_36_472# 0.033277f
C18470 _407_/a_36_472# _181_ 0.035594f
C18471 state\[1\] _113_ 0.107642f
C18472 _397_/a_244_68# net55 0.001173f
C18473 net16 FILLER_0_8_37/a_484_472# 0.004272f
C18474 mask\[0\] FILLER_0_15_212/a_1468_375# 0.001182f
C18475 _420_/a_1000_472# _009_ 0.019219f
C18476 _016_ _427_/a_448_472# 0.016416f
C18477 _450_/a_36_151# _039_ 0.018559f
C18478 net52 net23 0.093434f
C18479 _184_ vdd 0.202732f
C18480 _019_ net36 0.309649f
C18481 output14/a_224_472# _031_ 0.001077f
C18482 _379_/a_36_472# _166_ 0.038062f
C18483 _009_ _109_ 0.006736f
C18484 _101_ vdd 0.02756f
C18485 net18 _416_/a_448_472# 0.05521f
C18486 net50 net40 0.005105f
C18487 _443_/a_448_472# net13 0.002263f
C18488 _443_/a_796_472# net23 0.002306f
C18489 FILLER_0_9_28/a_36_472# output42/a_224_472# 0.010684f
C18490 _094_ net77 0.00405f
C18491 _250_/a_36_68# state\[2\] 0.038165f
C18492 output28/a_224_472# output29/a_224_472# 0.00289f
C18493 FILLER_0_3_78/a_36_472# _160_ 0.006564f
C18494 net50 _441_/a_1204_472# 0.006986f
C18495 net52 _441_/a_2665_112# 0.004975f
C18496 net50 trim_mask\[2\] 0.267074f
C18497 _440_/a_36_151# net47 0.013626f
C18498 FILLER_0_12_220/a_1020_375# vss 0.004698f
C18499 FILLER_0_12_220/a_1468_375# vdd 0.002801f
C18500 _188_ _120_ 0.046757f
C18501 FILLER_0_13_212/a_484_472# net79 0.00402f
C18502 _193_/a_36_160# net62 0.00227f
C18503 FILLER_0_4_49/a_124_375# net49 0.005427f
C18504 FILLER_0_4_49/a_484_472# net66 0.015555f
C18505 net55 _406_/a_36_159# 0.001219f
C18506 net72 FILLER_0_18_37/a_36_472# 0.043427f
C18507 net55 FILLER_0_18_37/a_572_375# 0.007169f
C18508 fanout50/a_36_160# _447_/a_2665_112# 0.002885f
C18509 FILLER_0_4_107/a_36_472# _160_ 0.009073f
C18510 _114_ _311_/a_66_473# 0.081048f
C18511 output44/a_224_472# net40 0.006489f
C18512 FILLER_0_17_72/a_572_375# vdd 0.002455f
C18513 FILLER_0_17_72/a_124_375# vss 0.048053f
C18514 FILLER_0_8_37/a_36_472# vdd 0.135405f
C18515 FILLER_0_8_37/a_572_375# vss 0.00282f
C18516 net52 fanout74/a_36_113# 0.001514f
C18517 FILLER_0_4_49/a_124_375# net68 0.008422f
C18518 net47 FILLER_0_4_91/a_36_472# 0.005186f
C18519 _274_/a_36_68# net4 0.037848f
C18520 FILLER_0_21_142/a_124_375# FILLER_0_21_133/a_124_375# 0.003228f
C18521 FILLER_0_9_28/a_124_375# FILLER_0_8_24/a_572_375# 0.05841f
C18522 _102_ _094_ 0.727442f
C18523 net74 _372_/a_786_69# 0.00149f
C18524 ctln[7] FILLER_0_0_130/a_124_375# 0.002726f
C18525 net50 _439_/a_1000_472# 0.005154f
C18526 net52 _439_/a_2248_156# 0.00258f
C18527 _072_ FILLER_0_10_214/a_124_375# 0.033245f
C18528 net82 _443_/a_36_151# 0.03565f
C18529 _070_ FILLER_0_11_109/a_36_472# 0.001091f
C18530 trimb[1] FILLER_0_18_2/a_1020_375# 0.01376f
C18531 _095_ FILLER_0_14_107/a_124_375# 0.01418f
C18532 _053_ FILLER_0_7_72/a_3172_472# 0.032946f
C18533 _425_/a_1204_472# net37 0.001403f
C18534 _013_ _183_ 0.00176f
C18535 _132_ _332_/a_36_472# 0.055537f
C18536 mask\[4\] FILLER_0_18_177/a_1828_472# 0.014226f
C18537 FILLER_0_13_100/a_124_375# vdd 0.039324f
C18538 _032_ trim_mask\[4\] 0.010578f
C18539 net38 _450_/a_448_472# 0.031891f
C18540 _010_ _420_/a_2248_156# 0.047408f
C18541 FILLER_0_18_209/a_36_472# _047_ 0.002672f
C18542 _131_ _331_/a_244_472# 0.002331f
C18543 _434_/a_2248_156# vdd 0.019386f
C18544 fanout79/a_36_160# _094_ 0.008308f
C18545 ctlp[1] FILLER_0_23_282/a_572_375# 0.009848f
C18546 mask\[8\] _437_/a_448_472# 0.008198f
C18547 _417_/a_1308_423# vss 0.002064f
C18548 FILLER_0_12_136/a_1468_375# vss 0.043987f
C18549 _030_ FILLER_0_3_78/a_36_472# 0.007376f
C18550 net49 FILLER_0_3_78/a_572_375# 0.066078f
C18551 _422_/a_448_472# _009_ 0.018984f
C18552 _012_ FILLER_0_23_60/a_36_472# 0.001572f
C18553 _277_/a_36_160# output34/a_224_472# 0.014508f
C18554 _031_ FILLER_0_2_111/a_484_472# 0.027347f
C18555 net69 FILLER_0_2_111/a_1380_472# 0.021896f
C18556 en clk 0.067072f
C18557 _379_/a_36_472# trim_mask\[1\] 0.003592f
C18558 _178_ _402_/a_1948_68# 0.00815f
C18559 _126_ FILLER_0_13_206/a_124_375# 0.002746f
C18560 net36 FILLER_0_18_76/a_124_375# 0.001741f
C18561 _065_ _447_/a_2248_156# 0.038629f
C18562 net23 _387_/a_36_113# 0.031688f
C18563 en_co_clk _171_ 0.003472f
C18564 _161_ _070_ 0.027757f
C18565 net70 vdd 0.858299f
C18566 FILLER_0_7_195/a_36_472# net21 0.005469f
C18567 _411_/a_36_151# net8 0.012319f
C18568 _141_ _098_ 0.0697f
C18569 net82 FILLER_0_2_177/a_124_375# 0.003837f
C18570 _140_ _354_/a_49_472# 0.004731f
C18571 _404_/a_36_472# _041_ 0.003068f
C18572 net78 _421_/a_448_472# 0.025808f
C18573 _077_ _229_/a_224_472# 0.001293f
C18574 net60 _421_/a_448_472# 0.052759f
C18575 net47 vdd 2.422992f
C18576 net61 fanout77/a_36_113# 0.080943f
C18577 _437_/a_448_472# vss 0.001524f
C18578 _437_/a_1308_423# vdd 0.005139f
C18579 _441_/a_2248_156# _164_ 0.040396f
C18580 trim_val\[2\] _164_ 0.005847f
C18581 net47 _365_/a_244_472# 0.001431f
C18582 FILLER_0_21_286/a_484_472# FILLER_0_23_290/a_124_375# 0.001404f
C18583 net31 net36 0.00943f
C18584 _074_ FILLER_0_3_221/a_1380_472# 0.001341f
C18585 _079_ FILLER_0_5_212/a_36_472# 0.005671f
C18586 _053_ _058_ 0.075418f
C18587 net55 FILLER_0_18_61/a_124_375# 0.040701f
C18588 _242_/a_36_160# FILLER_0_5_148/a_484_472# 0.003699f
C18589 FILLER_0_14_91/a_36_472# _095_ 0.014431f
C18590 FILLER_0_1_192/a_124_375# net21 0.067765f
C18591 net34 vss 0.481379f
C18592 _430_/a_36_151# _093_ 0.00184f
C18593 FILLER_0_14_81/a_36_472# _177_ 0.004294f
C18594 _086_ FILLER_0_7_104/a_572_375# 0.003137f
C18595 _063_ _445_/a_2248_156# 0.008121f
C18596 _326_/a_36_160# vss 0.002357f
C18597 output23/a_224_472# _049_ 0.001034f
C18598 net72 _012_ 0.002382f
C18599 mask\[5\] FILLER_0_19_195/a_36_472# 0.007596f
C18600 FILLER_0_7_72/a_2724_472# net50 0.007192f
C18601 FILLER_0_23_44/a_1468_375# vdd -0.013698f
C18602 result[7] FILLER_0_23_282/a_484_472# 0.013947f
C18603 net81 FILLER_0_15_212/a_1380_472# 0.003953f
C18604 en_co_clk _176_ 0.099475f
C18605 _017_ FILLER_0_14_107/a_932_472# 0.001941f
C18606 result[5] result[9] 0.064058f
C18607 _069_ net4 0.07542f
C18608 FILLER_0_18_107/a_932_472# FILLER_0_16_115/a_124_375# 0.001512f
C18609 cal_itt\[3\] calibrate 1.141592f
C18610 net15 FILLER_0_5_54/a_1380_472# 0.047774f
C18611 _067_ FILLER_0_12_20/a_572_375# 0.01186f
C18612 _147_ _208_/a_36_160# 0.006056f
C18613 fanout69/a_36_113# _032_ 0.003681f
C18614 _247_/a_36_160# _060_ 0.055366f
C18615 net72 FILLER_0_15_59/a_572_375# 0.00799f
C18616 net32 vdd 0.50705f
C18617 FILLER_0_4_152/a_36_472# net47 0.007541f
C18618 net52 trim_val\[4\] 0.21532f
C18619 mask\[3\] _094_ 0.00554f
C18620 _416_/a_448_472# net62 0.009111f
C18621 _094_ _283_/a_36_472# 0.004373f
C18622 _098_ _433_/a_2665_112# 0.01601f
C18623 FILLER_0_7_104/a_572_375# _154_ 0.020664f
C18624 output37/a_224_472# net64 0.110037f
C18625 _028_ FILLER_0_5_72/a_1020_375# 0.00123f
C18626 net17 _450_/a_2225_156# 0.033342f
C18627 FILLER_0_6_79/a_124_375# FILLER_0_6_47/a_3260_375# 0.012001f
C18628 _091_ FILLER_0_18_177/a_36_472# 0.012695f
C18629 output36/a_224_472# vdd 0.145046f
C18630 _077_ _439_/a_1308_423# 0.022235f
C18631 FILLER_0_9_60/a_124_375# vdd 0.005798f
C18632 net47 _452_/a_1040_527# 0.014695f
C18633 _096_ _113_ 0.650985f
C18634 mask\[9\] _438_/a_2665_112# 0.040085f
C18635 _183_ _179_ 0.017086f
C18636 FILLER_0_15_290/a_124_375# vdd 0.028723f
C18637 net64 net5 0.098088f
C18638 FILLER_0_17_226/a_124_375# fanout63/a_36_160# 0.008215f
C18639 _136_ FILLER_0_16_115/a_36_472# 0.013477f
C18640 FILLER_0_3_172/a_36_472# net22 0.012287f
C18641 FILLER_0_18_171/a_36_472# _141_ 0.002037f
C18642 _427_/a_448_472# _043_ 0.002896f
C18643 _226_/a_860_68# net21 0.00107f
C18644 _104_ result[8] 0.00201f
C18645 fanout66/a_36_113# _440_/a_36_151# 0.017895f
C18646 FILLER_0_8_127/a_124_375# _126_ 0.001799f
C18647 _285_/a_36_472# _045_ 0.00269f
C18648 _149_ _354_/a_49_472# 0.017453f
C18649 _424_/a_36_151# _012_ 0.005964f
C18650 _343_/a_665_69# mask\[3\] 0.001405f
C18651 ctln[0] net40 0.001334f
C18652 net65 en 0.001469f
C18653 _141_ FILLER_0_22_128/a_3172_472# 0.01947f
C18654 cal_count\[3\] _390_/a_36_68# 0.003074f
C18655 output8/a_224_472# net20 0.084627f
C18656 _257_/a_36_472# _122_ 0.007741f
C18657 _432_/a_36_151# FILLER_0_15_180/a_36_472# 0.002018f
C18658 _127_ _070_ 0.031272f
C18659 _282_/a_36_160# vdd 0.010099f
C18660 _075_ net59 0.01129f
C18661 trimb[1] _452_/a_2225_156# 0.004072f
C18662 output10/a_224_472# _411_/a_2665_112# 0.008469f
C18663 _112_ net37 0.070289f
C18664 _044_ FILLER_0_14_263/a_124_375# 0.001047f
C18665 FILLER_0_22_86/a_124_375# net71 0.002239f
C18666 _408_/a_1936_472# cal_count\[0\] 0.001434f
C18667 FILLER_0_5_128/a_36_472# net47 0.008459f
C18668 cal_count\[3\] _408_/a_718_524# 0.005968f
C18669 net27 fanout62/a_36_160# 0.005558f
C18670 _438_/a_2665_112# FILLER_0_19_111/a_36_472# 0.007491f
C18671 trim_val\[4\] _387_/a_36_113# 0.005339f
C18672 net76 _037_ 0.010891f
C18673 FILLER_0_17_282/a_124_375# vdd 0.004586f
C18674 _448_/a_448_472# vdd 0.02042f
C18675 _274_/a_36_68# net79 0.009814f
C18676 _087_ FILLER_0_5_181/a_124_375# 0.068f
C18677 cal_count\[3\] cal_count\[2\] 0.005307f
C18678 output44/a_224_472# net46 0.003211f
C18679 _359_/a_1044_488# _129_ 0.001111f
C18680 _077_ _311_/a_66_473# 0.002605f
C18681 _398_/a_36_113# _278_/a_36_160# 0.001636f
C18682 _088_ FILLER_0_3_172/a_2364_375# 0.002377f
C18683 _081_ _084_ 0.016804f
C18684 _431_/a_796_472# _137_ 0.002195f
C18685 FILLER_0_14_107/a_572_375# vdd 0.021509f
C18686 FILLER_0_14_107/a_124_375# vss 0.002674f
C18687 _059_ vss 0.714648f
C18688 _063_ FILLER_0_6_37/a_124_375# 0.012149f
C18689 output37/a_224_472# vss 0.026983f
C18690 _086_ FILLER_0_11_124/a_36_472# 0.010729f
C18691 FILLER_0_22_177/a_124_375# vss 0.002674f
C18692 FILLER_0_22_177/a_572_375# vdd -0.003694f
C18693 FILLER_0_1_98/a_124_375# trim_mask\[3\] 0.058544f
C18694 net69 _441_/a_796_472# 0.002057f
C18695 trim_val\[3\] _441_/a_2248_156# 0.027464f
C18696 cal_itt\[2\] FILLER_0_3_221/a_572_375# 0.060779f
C18697 net81 cal_itt\[1\] 0.387207f
C18698 FILLER_0_9_28/a_36_472# FILLER_0_10_28/a_36_472# 0.05841f
C18699 _328_/a_36_113# _114_ 0.058671f
C18700 net71 _437_/a_1000_472# 0.014459f
C18701 _447_/a_36_151# net69 0.001216f
C18702 _375_/a_36_68# vss 0.02182f
C18703 net5 vss 0.326032f
C18704 net63 FILLER_0_17_218/a_572_375# 0.006355f
C18705 _064_ _445_/a_2560_156# 0.005361f
C18706 cal_count\[3\] FILLER_0_11_124/a_36_472# 0.00702f
C18707 output34/a_224_472# _102_ 0.008577f
C18708 _261_/a_36_160# FILLER_0_5_148/a_36_472# 0.195478f
C18709 _070_ _071_ 0.001757f
C18710 FILLER_0_18_107/a_2364_375# _433_/a_36_151# 0.002106f
C18711 fanout66/a_36_113# vdd 0.049012f
C18712 _122_ FILLER_0_5_164/a_572_375# 0.001352f
C18713 net74 _059_ 0.004133f
C18714 _127_ FILLER_0_9_142/a_36_472# 0.004721f
C18715 _297_/a_36_472# mask\[6\] 0.02557f
C18716 _031_ _157_ 0.104339f
C18717 _273_/a_36_68# _070_ 0.013247f
C18718 _144_ _140_ 0.415736f
C18719 FILLER_0_8_127/a_124_375# _077_ 0.005095f
C18720 net20 FILLER_0_12_220/a_124_375# 0.003161f
C18721 net80 net36 0.036729f
C18722 FILLER_0_5_172/a_36_472# net47 0.0015f
C18723 _450_/a_36_151# clkc 0.033095f
C18724 _450_/a_1353_112# net6 0.054189f
C18725 net81 valid 0.11798f
C18726 _330_/a_224_472# _134_ 0.007508f
C18727 _308_/a_848_380# _114_ 0.005266f
C18728 FILLER_0_15_235/a_124_375# FILLER_0_14_235/a_124_375# 0.05841f
C18729 net75 net82 0.214597f
C18730 FILLER_0_12_136/a_932_472# FILLER_0_11_142/a_124_375# 0.001543f
C18731 _300_/a_224_472# _009_ 0.001405f
C18732 _439_/a_2665_112# trim_mask\[0\] 0.020363f
C18733 _415_/a_36_151# FILLER_0_11_282/a_124_375# 0.001822f
C18734 FILLER_0_10_78/a_932_472# net52 0.00207f
C18735 FILLER_0_12_136/a_1020_375# cal_count\[3\] 0.002916f
C18736 result[9] net19 0.540761f
C18737 _219_/a_36_160# net14 0.048037f
C18738 FILLER_0_18_177/a_1916_375# vdd 0.021f
C18739 _132_ _428_/a_1308_423# 0.027389f
C18740 FILLER_0_20_193/a_484_472# FILLER_0_19_195/a_124_375# 0.001543f
C18741 FILLER_0_4_107/a_36_472# _156_ 0.005297f
C18742 _428_/a_36_151# _131_ 0.00821f
C18743 result[7] FILLER_0_24_290/a_36_472# 0.005185f
C18744 ctln[1] FILLER_0_0_266/a_124_375# 0.01186f
C18745 _418_/a_1308_423# vss 0.001913f
C18746 _411_/a_2248_156# net75 0.032114f
C18747 _411_/a_1000_472# _000_ 0.023042f
C18748 _072_ _055_ 0.083351f
C18749 _419_/a_2560_156# vdd 0.003021f
C18750 _419_/a_2665_112# vss 0.004064f
C18751 _136_ _451_/a_2449_156# 0.004653f
C18752 net26 FILLER_0_21_28/a_1380_472# 0.035291f
C18753 FILLER_0_2_171/a_124_375# net22 0.009924f
C18754 FILLER_0_14_91/a_36_472# vss 0.001729f
C18755 FILLER_0_14_91/a_484_472# vdd 0.00605f
C18756 net48 _079_ 0.012855f
C18757 state\[1\] vdd 0.544231f
C18758 _155_ _163_ 0.296236f
C18759 _026_ _437_/a_448_472# 0.026072f
C18760 net41 _446_/a_36_151# 0.143017f
C18761 _453_/a_2248_156# vss 0.031525f
C18762 _453_/a_2665_112# vdd 0.005481f
C18763 _012_ FILLER_0_21_60/a_36_472# 0.017483f
C18764 _089_ FILLER_0_3_172/a_2276_472# 0.001522f
C18765 _114_ _428_/a_36_151# 0.008132f
C18766 net31 result[6] 0.002094f
C18767 _002_ _088_ 0.003969f
C18768 FILLER_0_10_214/a_36_472# _070_ 0.014734f
C18769 output35/a_224_472# net22 0.028095f
C18770 _069_ net79 0.045808f
C18771 _119_ _326_/a_36_160# 0.003944f
C18772 FILLER_0_15_212/a_484_472# mask\[1\] 0.007258f
C18773 FILLER_0_13_142/a_1020_375# net23 0.047331f
C18774 _425_/a_2248_156# calibrate 0.022237f
C18775 _003_ net37 0.046745f
C18776 output34/a_224_472# _198_/a_67_603# 0.00179f
C18777 FILLER_0_20_2/a_572_375# vss 0.001471f
C18778 FILLER_0_20_2/a_36_472# vdd 0.102471f
C18779 _053_ net52 0.042556f
C18780 FILLER_0_5_212/a_36_472# vss 0.00578f
C18781 FILLER_0_9_28/a_1916_375# _453_/a_36_151# 0.001543f
C18782 FILLER_0_18_177/a_3172_472# net21 0.010321f
C18783 _018_ FILLER_0_15_205/a_124_375# 0.002309f
C18784 trim_val\[4\] FILLER_0_5_164/a_484_472# 0.00172f
C18785 FILLER_0_16_57/a_1380_472# _175_ 0.002834f
C18786 FILLER_0_13_212/a_1468_375# net62 0.003327f
C18787 _341_/a_49_472# mask\[2\] 0.026222f
C18788 trim_val\[1\] vss 0.029927f
C18789 FILLER_0_1_266/a_36_472# vdd 0.008551f
C18790 FILLER_0_1_266/a_572_375# vss 0.001919f
C18791 net18 FILLER_0_9_282/a_124_375# 0.024657f
C18792 FILLER_0_8_107/a_124_375# _134_ 0.007753f
C18793 FILLER_0_2_165/a_124_375# net22 0.206491f
C18794 _151_ _153_ 0.027868f
C18795 mask\[5\] FILLER_0_20_193/a_124_375# 0.015793f
C18796 _236_/a_36_160# _444_/a_36_151# 0.034413f
C18797 FILLER_0_9_28/a_1828_472# net68 0.048468f
C18798 net80 FILLER_0_20_169/a_36_472# 0.024142f
C18799 FILLER_0_17_38/a_572_375# _182_ 0.035561f
C18800 _255_/a_224_552# _161_ 0.025424f
C18801 output34/a_224_472# mask\[3\] 0.002385f
C18802 _328_/a_36_113# _126_ 0.023932f
C18803 net56 fanout56/a_36_113# 0.015924f
C18804 cal_count\[2\] _278_/a_36_160# 0.023061f
C18805 FILLER_0_17_200/a_124_375# _432_/a_2665_112# 0.006271f
C18806 ctlp[9] FILLER_0_23_44/a_932_472# 0.001195f
C18807 _144_ _149_ 0.032178f
C18808 result[8] FILLER_0_24_274/a_932_472# 0.005458f
C18809 mask\[4\] FILLER_0_19_195/a_124_375# 0.006236f
C18810 _370_/a_124_24# _160_ 0.001126f
C18811 _205_/a_36_160# _048_ 0.040317f
C18812 result[9] _009_ 0.19745f
C18813 FILLER_0_6_47/a_36_472# vdd 0.090192f
C18814 FILLER_0_6_47/a_3260_375# vss 0.061766f
C18815 FILLER_0_15_212/a_932_472# vdd 0.001767f
C18816 FILLER_0_7_195/a_36_472# _062_ 0.0045f
C18817 _164_ _167_ 0.311625f
C18818 _093_ FILLER_0_17_72/a_572_375# 0.005609f
C18819 _402_/a_718_527# vdd 0.020893f
C18820 output32/a_224_472# net20 0.050019f
C18821 trim_mask\[4\] _386_/a_848_380# 0.001657f
C18822 net32 net78 0.055231f
C18823 net32 net60 0.509175f
C18824 result[5] net61 0.092275f
C18825 cal clk 0.033015f
C18826 FILLER_0_4_49/a_124_375# net47 0.006524f
C18827 _339_/a_36_160# _140_ 0.025058f
C18828 fanout52/a_36_160# _170_ 0.024724f
C18829 _009_ FILLER_0_23_282/a_36_472# 0.005974f
C18830 _304_/a_224_472# vss 0.001746f
C18831 FILLER_0_4_197/a_1020_375# net22 0.040565f
C18832 FILLER_0_8_247/a_484_472# calibrate 0.009318f
C18833 _152_ net23 0.001895f
C18834 _077_ FILLER_0_10_78/a_1020_375# 0.001131f
C18835 _070_ _246_/a_36_68# 0.056186f
C18836 _419_/a_1000_472# net77 0.001113f
C18837 FILLER_0_15_150/a_124_375# net36 0.005687f
C18838 _105_ vdd 0.565718f
C18839 _323_/a_36_113# _060_ 0.002584f
C18840 _422_/a_1308_423# mask\[7\] 0.045368f
C18841 net57 _333_/a_36_160# 0.008292f
C18842 _057_ state\[1\] 0.284428f
C18843 net52 _443_/a_1000_472# 0.016322f
C18844 output8/a_224_472# _073_ 0.043098f
C18845 FILLER_0_19_125/a_124_375# _145_ 0.006777f
C18846 cal_count\[2\] FILLER_0_15_2/a_124_375# 0.033559f
C18847 _072_ _058_ 0.029688f
C18848 _168_ vss 0.171346f
C18849 _426_/a_1308_423# calibrate 0.001708f
C18850 output26/a_224_472# vss 0.0137f
C18851 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1380_472# 0.013276f
C18852 fanout58/a_36_160# fanout59/a_36_160# 0.001216f
C18853 _119_ _059_ 0.039711f
C18854 FILLER_0_11_142/a_124_375# FILLER_0_11_135/a_124_375# 0.004426f
C18855 _077_ FILLER_0_9_72/a_932_472# 0.006408f
C18856 net15 FILLER_0_6_47/a_2364_375# 0.022624f
C18857 _028_ _077_ 0.017713f
C18858 _126_ _428_/a_36_151# 0.032026f
C18859 fanout74/a_36_113# _152_ 0.017267f
C18860 fanout76/a_36_160# net18 0.003319f
C18861 _453_/a_1204_472# _042_ 0.002408f
C18862 _113_ FILLER_0_15_180/a_124_375# 0.001512f
C18863 fanout53/a_36_160# _427_/a_2665_112# 0.00285f
C18864 net31 mask\[4\] 0.499009f
C18865 _346_/a_665_69# mask\[4\] 0.001125f
C18866 _093_ net70 0.001888f
C18867 _051_ vdd 0.036931f
C18868 _402_/a_728_93# _180_ 0.008035f
C18869 net7 _446_/a_36_151# 0.001237f
C18870 FILLER_0_18_53/a_484_472# vss 0.003579f
C18871 output38/a_224_472# vdd -0.006652f
C18872 FILLER_0_16_89/a_1468_375# _131_ 0.016581f
C18873 _119_ _375_/a_36_68# 0.007338f
C18874 _433_/a_1204_472# _022_ 0.005308f
C18875 _010_ vdd 0.121474f
C18876 _430_/a_448_472# net63 0.026599f
C18877 FILLER_0_4_107/a_1468_375# net47 0.012534f
C18878 FILLER_0_21_125/a_124_375# _098_ 0.006462f
C18879 _247_/a_36_160# vss 0.009308f
C18880 output23/a_224_472# ctlp[6] 0.024575f
C18881 fanout81/a_36_160# net82 0.027351f
C18882 FILLER_0_4_197/a_124_375# _079_ 0.004772f
C18883 FILLER_0_5_181/a_124_375# vdd 0.009553f
C18884 net4 _090_ 0.06324f
C18885 net23 _348_/a_49_472# 0.0037f
C18886 FILLER_0_21_28/a_572_375# vdd 0.013051f
C18887 FILLER_0_3_172/a_3260_375# vdd -0.013516f
C18888 FILLER_0_16_241/a_124_375# net30 0.028559f
C18889 FILLER_0_9_223/a_36_472# _070_ 0.006158f
C18890 FILLER_0_9_223/a_124_375# _076_ 0.004399f
C18891 ctln[0] trim[3] 0.216084f
C18892 _104_ net63 0.005363f
C18893 net4 FILLER_0_3_221/a_572_375# 0.030599f
C18894 _413_/a_1000_472# net82 0.002029f
C18895 _385_/a_36_68# vdd 0.01625f
C18896 net60 FILLER_0_17_282/a_124_375# 0.039003f
C18897 _029_ _156_ 0.018258f
C18898 mask\[7\] net22 0.275179f
C18899 FILLER_0_17_56/a_572_375# _183_ 0.002605f
C18900 _035_ net40 0.068572f
C18901 net50 FILLER_0_5_88/a_36_472# 0.00867f
C18902 _077_ _308_/a_848_380# 0.010515f
C18903 _173_ _450_/a_3129_107# 0.00264f
C18904 mask\[3\] net21 0.100738f
C18905 _446_/a_2665_112# net66 0.00195f
C18906 net22 net59 0.195226f
C18907 trim_mask\[2\] _035_ 0.004455f
C18908 FILLER_0_6_239/a_124_375# net76 0.001286f
C18909 FILLER_0_5_72/a_1468_375# net49 0.001276f
C18910 _112_ _122_ 0.120159f
C18911 _062_ _226_/a_860_68# 0.001842f
C18912 _096_ vdd 0.557569f
C18913 _136_ net23 0.031512f
C18914 _005_ _416_/a_796_472# 0.009162f
C18915 net52 _164_ 0.313379f
C18916 net4 net22 0.036966f
C18917 _443_/a_448_472# _170_ 0.056211f
C18918 net81 net59 0.074175f
C18919 FILLER_0_7_59/a_124_375# FILLER_0_6_47/a_1468_375# 0.05841f
C18920 _132_ FILLER_0_17_104/a_572_375# 0.003857f
C18921 _139_ mask\[2\] 0.035793f
C18922 net76 FILLER_0_3_172/a_572_375# 0.003315f
C18923 _415_/a_1308_423# FILLER_0_9_270/a_124_375# 0.001064f
C18924 FILLER_0_19_47/a_484_472# _052_ 0.01589f
C18925 ctln[1] _411_/a_1204_472# 0.031348f
C18926 FILLER_0_5_72/a_484_472# trim_mask\[1\] 0.012321f
C18927 net81 net4 0.003327f
C18928 FILLER_0_4_152/a_124_375# _386_/a_124_24# 0.010472f
C18929 _183_ _041_ 0.001931f
C18930 _431_/a_2665_112# _136_ 0.035394f
C18931 _412_/a_448_472# net18 0.049704f
C18932 net79 result[3] 0.138076f
C18933 ctln[3] FILLER_0_0_232/a_124_375# 0.012394f
C18934 _070_ net23 0.047632f
C18935 net65 cal 0.023638f
C18936 FILLER_0_7_233/a_124_375# vdd 0.03915f
C18937 net38 _452_/a_36_151# 0.010095f
C18938 FILLER_0_2_111/a_1380_472# vss 0.001679f
C18939 _317_/a_36_113# _123_ 0.037893f
C18940 _175_ _040_ 0.00133f
C18941 _188_ _453_/a_796_472# 0.00103f
C18942 FILLER_0_21_286/a_484_472# net18 0.001956f
C18943 result[7] result[8] 0.201281f
C18944 _114_ _085_ 0.056448f
C18945 trimb[2] trimb[3] 0.369908f
C18946 _134_ vss 0.088213f
C18947 _431_/a_448_472# net73 0.050964f
C18948 _414_/a_2248_156# _122_ 0.002838f
C18949 net48 vss 0.161385f
C18950 mask\[3\] FILLER_0_18_177/a_124_375# 0.002924f
C18951 _043_ FILLER_0_12_196/a_36_472# 0.001526f
C18952 _187_ _408_/a_728_93# 0.002598f
C18953 net35 FILLER_0_21_150/a_36_472# 0.004456f
C18954 fanout56/a_36_113# _095_ 0.004331f
C18955 output29/a_224_472# net29 0.038602f
C18956 _103_ _418_/a_1308_423# 0.004778f
C18957 _091_ _429_/a_1308_423# 0.031247f
C18958 net61 net19 0.132027f
C18959 net60 _418_/a_796_472# 0.008602f
C18960 net20 _419_/a_1204_472# 0.006482f
C18961 ctln[1] input1/a_36_113# 0.004419f
C18962 net60 _419_/a_2560_156# 0.006989f
C18963 _136_ FILLER_0_15_180/a_484_472# 0.002128f
C18964 _207_/a_67_603# mask\[6\] 0.072291f
C18965 vdd FILLER_0_13_72/a_124_375# -0.004549f
C18966 _141_ _137_ 0.40175f
C18967 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_124_375# 0.004426f
C18968 net34 _295_/a_36_472# 0.032003f
C18969 _146_ vss 0.078821f
C18970 net58 FILLER_0_9_282/a_572_375# 0.006142f
C18971 _111_ net71 0.002668f
C18972 result[4] _417_/a_36_151# 0.010571f
C18973 net80 FILLER_0_16_154/a_1468_375# 0.013593f
C18974 trim_mask\[4\] FILLER_0_2_165/a_36_472# 0.265591f
C18975 _432_/a_1308_423# _091_ 0.008903f
C18976 _046_ net30 0.006105f
C18977 FILLER_0_23_60/a_36_472# vdd 0.090554f
C18978 FILLER_0_23_60/a_124_375# vss 0.004081f
C18979 FILLER_0_6_177/a_124_375# vss 0.002362f
C18980 FILLER_0_6_177/a_572_375# vdd 0.02743f
C18981 ctlp[1] FILLER_0_23_290/a_36_472# 0.038596f
C18982 _141_ FILLER_0_19_171/a_36_472# 0.001292f
C18983 _052_ FILLER_0_21_60/a_124_375# 0.002308f
C18984 net65 FILLER_0_2_177/a_124_375# 0.018094f
C18985 _118_ _331_/a_448_472# 0.001166f
C18986 FILLER_0_9_28/a_124_375# net17 0.009179f
C18987 net55 FILLER_0_11_78/a_572_375# 0.002321f
C18988 FILLER_0_9_142/a_36_472# net23 0.001099f
C18989 net19 net37 0.030961f
C18990 _076_ net59 0.005449f
C18991 _099_ FILLER_0_15_235/a_484_472# 0.002657f
C18992 net21 FILLER_0_12_196/a_36_472# 0.001298f
C18993 FILLER_0_17_161/a_124_375# mask\[2\] 0.00227f
C18994 net4 _076_ 1.140706f
C18995 FILLER_0_21_142/a_36_472# net35 0.003079f
C18996 FILLER_0_24_96/a_36_472# net24 0.028193f
C18997 FILLER_0_16_255/a_124_375# _006_ 0.02007f
C18998 _057_ _096_ 0.001547f
C18999 _088_ net76 0.214494f
C19000 FILLER_0_5_109/a_36_472# FILLER_0_4_107/a_124_375# 0.001684f
C19001 _178_ _174_ 0.012157f
C19002 _423_/a_36_151# FILLER_0_23_44/a_932_472# 0.001723f
C19003 _075_ cal_itt\[3\] 0.731221f
C19004 _003_ _122_ 0.033778f
C19005 _068_ _311_/a_254_473# 0.002606f
C19006 mask\[4\] net80 0.034957f
C19007 net31 net34 0.080525f
C19008 _275_/a_224_472# vss 0.001498f
C19009 FILLER_0_15_116/a_484_472# net36 0.009319f
C19010 _427_/a_1000_472# _095_ 0.021594f
C19011 net68 FILLER_0_5_54/a_36_472# 0.012107f
C19012 _431_/a_2560_156# net53 0.002265f
C19013 _074_ _078_ 0.003088f
C19014 _396_/a_224_472# _176_ 0.008359f
C19015 _354_/a_49_472# _098_ 0.009677f
C19016 _133_ _313_/a_67_603# 0.002974f
C19017 FILLER_0_18_2/a_2276_472# net47 0.001369f
C19018 FILLER_0_18_139/a_124_375# FILLER_0_18_107/a_3260_375# 0.012552f
C19019 FILLER_0_4_99/a_36_472# vdd 0.094733f
C19020 FILLER_0_4_99/a_124_375# vss 0.017518f
C19021 FILLER_0_0_266/a_36_472# rstn 0.006108f
C19022 FILLER_0_5_54/a_932_472# trim_mask\[1\] 0.016187f
C19023 net72 vdd 1.425686f
C19024 _111_ _013_ 0.024203f
C19025 FILLER_0_13_65/a_124_375# net72 0.002341f
C19026 _118_ _315_/a_244_497# 0.003007f
C19027 FILLER_0_21_142/a_484_472# vss 0.034607f
C19028 _058_ FILLER_0_10_94/a_484_472# 0.002096f
C19029 mask\[4\] FILLER_0_18_139/a_1468_375# 0.023004f
C19030 net20 FILLER_0_15_212/a_1468_375# 0.006824f
C19031 _095_ _281_/a_234_472# 0.001467f
C19032 _034_ 0 0.304805f
C19033 _160_ 0 1.542665f
C19034 _166_ 0 0.299751f
C19035 trim[3] 0 1.777626f
C19036 output41/a_224_472# 0 2.38465f
C19037 clkc 0 0.763769f
C19038 net6 0 1.112469f
C19039 output6/a_224_472# 0 2.38465f
C19040 FILLER_0_12_196/a_36_472# 0 0.417394f
C19041 FILLER_0_12_196/a_124_375# 0 0.246306f
C19042 result[3] 0 0.50376f
C19043 net30 0 1.81422f
C19044 output30/a_224_472# 0 2.38465f
C19045 _047_ 0 0.374694f
C19046 _201_/a_67_603# 0 0.345683f
C19047 net62 0 4.932099f
C19048 _416_/a_2560_156# 0 0.016968f
C19049 _416_/a_2665_112# 0 0.62251f
C19050 _416_/a_2248_156# 0 0.371662f
C19051 _416_/a_1204_472# 0 0.012971f
C19052 _416_/a_1000_472# 0 0.291735f
C19053 _416_/a_796_472# 0 0.023206f
C19054 _416_/a_1308_423# 0 0.279043f
C19055 _416_/a_448_472# 0 0.684413f
C19056 _416_/a_36_151# 0 1.43589f
C19057 FILLER_0_13_290/a_36_472# 0 0.417394f
C19058 FILLER_0_13_290/a_124_375# 0 0.246306f
C19059 _278_/a_36_160# 0 0.696445f
C19060 _145_ 0 0.546455f
C19061 FILLER_0_13_72/a_484_472# 0 0.345058f
C19062 FILLER_0_13_72/a_36_472# 0 0.404746f
C19063 FILLER_0_13_72/a_572_375# 0 0.232991f
C19064 FILLER_0_13_72/a_124_375# 0 0.185089f
C19065 FILLER_0_14_235/a_484_472# 0 0.345058f
C19066 FILLER_0_14_235/a_36_472# 0 0.404746f
C19067 FILLER_0_14_235/a_572_375# 0 0.232991f
C19068 FILLER_0_14_235/a_124_375# 0 0.185089f
C19069 _156_ 0 0.593796f
C19070 _107_ 0 0.391583f
C19071 _295_/a_36_472# 0 0.031137f
C19072 _022_ 0 0.387773f
C19073 _433_/a_2560_156# 0 0.016968f
C19074 _433_/a_2665_112# 0 0.62251f
C19075 _433_/a_2248_156# 0 0.371662f
C19076 _433_/a_1204_472# 0 0.012971f
C19077 _433_/a_1000_472# 0 0.291735f
C19078 _433_/a_796_472# 0 0.023206f
C19079 _433_/a_1308_423# 0 0.279043f
C19080 _433_/a_448_472# 0 0.684413f
C19081 _433_/a_36_151# 0 1.43589f
C19082 FILLER_0_5_148/a_484_472# 0 0.345058f
C19083 FILLER_0_5_148/a_36_472# 0 0.404746f
C19084 FILLER_0_5_148/a_572_375# 0 0.232991f
C19085 FILLER_0_5_148/a_124_375# 0 0.185089f
C19086 _167_ 0 0.285904f
C19087 _381_/a_36_472# 0 0.031137f
C19088 trim[2] 0 0.79181f
C19089 net40 0 1.845219f
C19090 output40/a_224_472# 0 2.38465f
C19091 cal_count\[0\] 0 0.893784f
C19092 _039_ 0 0.412301f
C19093 _450_/a_2449_156# 0 0.049992f
C19094 _450_/a_2225_156# 0 0.434082f
C19095 _450_/a_3129_107# 0 0.58406f
C19096 _450_/a_836_156# 0 0.019766f
C19097 _450_/a_1040_527# 0 0.302082f
C19098 _450_/a_1353_112# 0 0.286513f
C19099 _450_/a_448_472# 0 1.21246f
C19100 _450_/a_36_151# 0 1.31409f
C19101 rstn 0 1.86494f
C19102 FILLER_0_8_156/a_484_472# 0 0.345058f
C19103 FILLER_0_8_156/a_36_472# 0 0.404746f
C19104 FILLER_0_8_156/a_572_375# 0 0.232991f
C19105 FILLER_0_8_156/a_124_375# 0 0.185089f
C19106 FILLER_0_6_37/a_36_472# 0 0.417394f
C19107 FILLER_0_6_37/a_124_375# 0 0.246306f
C19108 FILLER_0_21_60/a_484_472# 0 0.345058f
C19109 FILLER_0_21_60/a_36_472# 0 0.404746f
C19110 FILLER_0_21_60/a_572_375# 0 0.232991f
C19111 FILLER_0_21_60/a_124_375# 0 0.185089f
C19112 FILLER_0_22_107/a_484_472# 0 0.345058f
C19113 FILLER_0_22_107/a_36_472# 0 0.404746f
C19114 FILLER_0_22_107/a_572_375# 0 0.232991f
C19115 FILLER_0_22_107/a_124_375# 0 0.185089f
C19116 FILLER_0_16_115/a_36_472# 0 0.417394f
C19117 FILLER_0_16_115/a_124_375# 0 0.246306f
C19118 FILLER_0_19_134/a_36_472# 0 0.417394f
C19119 FILLER_0_19_134/a_124_375# 0 0.246306f
C19120 FILLER_0_3_212/a_36_472# 0 0.417394f
C19121 FILLER_0_3_212/a_124_375# 0 0.246306f
C19122 FILLER_0_10_94/a_484_472# 0 0.345058f
C19123 FILLER_0_10_94/a_36_472# 0 0.404746f
C19124 FILLER_0_10_94/a_572_375# 0 0.232991f
C19125 FILLER_0_10_94/a_124_375# 0 0.185089f
C19126 FILLER_0_4_91/a_484_472# 0 0.345058f
C19127 FILLER_0_4_91/a_36_472# 0 0.404746f
C19128 FILLER_0_4_91/a_572_375# 0 0.232991f
C19129 FILLER_0_4_91/a_124_375# 0 0.185089f
C19130 net14 0 1.508711f
C19131 _202_/a_36_160# 0 0.696445f
C19132 FILLER_0_6_231/a_484_472# 0 0.345058f
C19133 FILLER_0_6_231/a_36_472# 0 0.404746f
C19134 FILLER_0_6_231/a_572_375# 0 0.232991f
C19135 FILLER_0_6_231/a_124_375# 0 0.185089f
C19136 vss 0 65.60368f
C19137 vdd 0 1.086009p
C19138 _006_ 0 0.41456f
C19139 _417_/a_2560_156# 0 0.016968f
C19140 _417_/a_2665_112# 0 0.62251f
C19141 _417_/a_2248_156# 0 0.371662f
C19142 _417_/a_1204_472# 0 0.012971f
C19143 _417_/a_1000_472# 0 0.291735f
C19144 _417_/a_796_472# 0 0.023206f
C19145 _417_/a_1308_423# 0 0.279043f
C19146 _417_/a_448_472# 0 0.684413f
C19147 _417_/a_36_151# 0 1.43589f
C19148 _146_ 0 0.35443f
C19149 mask\[6\] 0 1.246962f
C19150 _348_/a_49_472# 0 0.054843f
C19151 _365_/a_36_68# 0 0.150048f
C19152 _023_ 0 0.345812f
C19153 _434_/a_2560_156# 0 0.016968f
C19154 _434_/a_2665_112# 0 0.62251f
C19155 _434_/a_2248_156# 0 0.371662f
C19156 _434_/a_1204_472# 0 0.012971f
C19157 _434_/a_1000_472# 0 0.291735f
C19158 _434_/a_796_472# 0 0.023206f
C19159 _434_/a_1308_423# 0 0.279043f
C19160 _434_/a_448_472# 0 0.684413f
C19161 _434_/a_36_151# 0 1.43589f
C19162 FILLER_0_5_136/a_36_472# 0 0.417394f
C19163 FILLER_0_5_136/a_124_375# 0 0.246306f
C19164 FILLER_0_18_209/a_484_472# 0 0.345058f
C19165 FILLER_0_18_209/a_36_472# 0 0.404746f
C19166 FILLER_0_18_209/a_572_375# 0 0.232991f
C19167 FILLER_0_18_209/a_124_375# 0 0.185089f
C19168 FILLER_0_12_28/a_36_472# 0 0.417394f
C19169 FILLER_0_12_28/a_124_375# 0 0.246306f
C19170 _040_ 0 0.355703f
C19171 _451_/a_2449_156# 0 0.049992f
C19172 _451_/a_2225_156# 0 0.434082f
C19173 _451_/a_3129_107# 0 0.58406f
C19174 _451_/a_836_156# 0 0.019766f
C19175 _451_/a_1040_527# 0 0.302082f
C19176 _451_/a_1353_112# 0 0.286513f
C19177 _451_/a_448_472# 0 1.21246f
C19178 _451_/a_36_151# 0 1.31409f
C19179 FILLER_0_6_47/a_3172_472# 0 0.345058f
C19180 FILLER_0_6_47/a_2724_472# 0 0.33241f
C19181 FILLER_0_6_47/a_2276_472# 0 0.33241f
C19182 FILLER_0_6_47/a_1828_472# 0 0.33241f
C19183 FILLER_0_6_47/a_1380_472# 0 0.33241f
C19184 FILLER_0_6_47/a_932_472# 0 0.33241f
C19185 FILLER_0_6_47/a_484_472# 0 0.33241f
C19186 FILLER_0_6_47/a_36_472# 0 0.404746f
C19187 FILLER_0_6_47/a_3260_375# 0 0.233093f
C19188 FILLER_0_6_47/a_2812_375# 0 0.17167f
C19189 FILLER_0_6_47/a_2364_375# 0 0.17167f
C19190 FILLER_0_6_47/a_1916_375# 0 0.17167f
C19191 FILLER_0_6_47/a_1468_375# 0 0.17167f
C19192 FILLER_0_6_47/a_1020_375# 0 0.17167f
C19193 FILLER_0_6_47/a_572_375# 0 0.17167f
C19194 FILLER_0_6_47/a_124_375# 0 0.185915f
C19195 FILLER_0_21_150/a_36_472# 0 0.417394f
C19196 FILLER_0_21_150/a_124_375# 0 0.246306f
C19197 FILLER_0_15_180/a_484_472# 0 0.345058f
C19198 FILLER_0_15_180/a_36_472# 0 0.404746f
C19199 FILLER_0_15_180/a_572_375# 0 0.232991f
C19200 FILLER_0_15_180/a_124_375# 0 0.185089f
C19201 FILLER_0_22_128/a_3172_472# 0 0.345058f
C19202 FILLER_0_22_128/a_2724_472# 0 0.33241f
C19203 FILLER_0_22_128/a_2276_472# 0 0.33241f
C19204 FILLER_0_22_128/a_1828_472# 0 0.33241f
C19205 FILLER_0_22_128/a_1380_472# 0 0.33241f
C19206 FILLER_0_22_128/a_932_472# 0 0.33241f
C19207 FILLER_0_22_128/a_484_472# 0 0.33241f
C19208 FILLER_0_22_128/a_36_472# 0 0.404746f
C19209 FILLER_0_22_128/a_3260_375# 0 0.233093f
C19210 FILLER_0_22_128/a_2812_375# 0 0.17167f
C19211 FILLER_0_22_128/a_2364_375# 0 0.17167f
C19212 FILLER_0_22_128/a_1916_375# 0 0.17167f
C19213 FILLER_0_22_128/a_1468_375# 0 0.17167f
C19214 FILLER_0_22_128/a_1020_375# 0 0.17167f
C19215 FILLER_0_22_128/a_572_375# 0 0.17167f
C19216 FILLER_0_22_128/a_124_375# 0 0.185915f
C19217 FILLER_0_19_111/a_484_472# 0 0.345058f
C19218 FILLER_0_19_111/a_36_472# 0 0.404746f
C19219 FILLER_0_19_111/a_572_375# 0 0.232991f
C19220 FILLER_0_19_111/a_124_375# 0 0.185089f
C19221 FILLER_0_19_155/a_484_472# 0 0.345058f
C19222 FILLER_0_19_155/a_36_472# 0 0.404746f
C19223 FILLER_0_19_155/a_572_375# 0 0.232991f
C19224 FILLER_0_19_155/a_124_375# 0 0.185089f
C19225 net11 0 1.328455f
C19226 net21 0 1.922829f
C19227 _007_ 0 0.309495f
C19228 net77 0 1.39077f
C19229 _418_/a_2560_156# 0 0.016968f
C19230 _418_/a_2665_112# 0 0.62251f
C19231 _418_/a_2248_156# 0 0.371662f
C19232 _418_/a_1204_472# 0 0.012971f
C19233 _418_/a_1000_472# 0 0.291735f
C19234 _418_/a_796_472# 0 0.023206f
C19235 _418_/a_1308_423# 0 0.279043f
C19236 _418_/a_448_472# 0 0.684413f
C19237 _418_/a_36_151# 0 1.43589f
C19238 _220_/a_67_603# 0 0.345683f
C19239 FILLER_0_9_282/a_484_472# 0 0.345058f
C19240 FILLER_0_9_282/a_36_472# 0 0.404746f
C19241 FILLER_0_9_282/a_572_375# 0 0.232991f
C19242 FILLER_0_9_282/a_124_375# 0 0.185089f
C19243 FILLER_0_18_37/a_1380_472# 0 0.345058f
C19244 FILLER_0_18_37/a_932_472# 0 0.33241f
C19245 FILLER_0_18_37/a_484_472# 0 0.33241f
C19246 FILLER_0_18_37/a_36_472# 0 0.404746f
C19247 FILLER_0_18_37/a_1468_375# 0 0.233029f
C19248 FILLER_0_18_37/a_1020_375# 0 0.171606f
C19249 FILLER_0_18_37/a_572_375# 0 0.171606f
C19250 FILLER_0_18_37/a_124_375# 0 0.185399f
C19251 FILLER_0_2_127/a_36_472# 0 0.417394f
C19252 FILLER_0_2_127/a_124_375# 0 0.246306f
C19253 _157_ 0 0.531763f
C19254 _435_/a_2560_156# 0 0.016968f
C19255 _435_/a_2665_112# 0 0.62251f
C19256 _435_/a_2248_156# 0 0.371662f
C19257 _435_/a_1204_472# 0 0.012971f
C19258 _435_/a_1000_472# 0 0.291735f
C19259 _435_/a_796_472# 0 0.023206f
C19260 _435_/a_1308_423# 0 0.279043f
C19261 _435_/a_448_472# 0 0.684413f
C19262 _435_/a_36_151# 0 1.43589f
C19263 _108_ 0 0.411979f
C19264 _297_/a_36_472# 0 0.031137f
C19265 trim_mask\[3\] 0 1.081535f
C19266 _164_ 0 1.3268f
C19267 _383_/a_36_472# 0 0.031137f
C19268 _041_ 0 0.299289f
C19269 _452_/a_2449_156# 0 0.049992f
C19270 _452_/a_2225_156# 0 0.434082f
C19271 _452_/a_3129_107# 0 0.58406f
C19272 _452_/a_836_156# 0 0.019766f
C19273 _452_/a_1040_527# 0 0.302082f
C19274 _452_/a_1353_112# 0 0.286513f
C19275 _452_/a_448_472# 0 1.21246f
C19276 _452_/a_36_151# 0 1.31409f
C19277 FILLER_0_6_79/a_36_472# 0 0.417394f
C19278 FILLER_0_6_79/a_124_375# 0 0.246306f
C19279 net59 0 5.044369f
C19280 FILLER_0_15_59/a_484_472# 0 0.345058f
C19281 FILLER_0_15_59/a_36_472# 0 0.404746f
C19282 FILLER_0_15_59/a_572_375# 0 0.232991f
C19283 FILLER_0_15_59/a_124_375# 0 0.185089f
C19284 FILLER_0_3_221/a_1380_472# 0 0.345058f
C19285 FILLER_0_3_221/a_932_472# 0 0.33241f
C19286 FILLER_0_3_221/a_484_472# 0 0.33241f
C19287 FILLER_0_3_221/a_36_472# 0 0.404746f
C19288 FILLER_0_3_221/a_1468_375# 0 0.233029f
C19289 FILLER_0_3_221/a_1020_375# 0 0.171606f
C19290 FILLER_0_3_221/a_572_375# 0 0.171606f
C19291 FILLER_0_3_221/a_124_375# 0 0.185399f
C19292 FILLER_0_19_187/a_484_472# 0 0.345058f
C19293 FILLER_0_19_187/a_36_472# 0 0.404746f
C19294 FILLER_0_19_187/a_572_375# 0 0.232991f
C19295 FILLER_0_19_187/a_124_375# 0 0.185089f
C19296 FILLER_0_20_15/a_1380_472# 0 0.345058f
C19297 FILLER_0_20_15/a_932_472# 0 0.33241f
C19298 FILLER_0_20_15/a_484_472# 0 0.33241f
C19299 FILLER_0_20_15/a_36_472# 0 0.404746f
C19300 FILLER_0_20_15/a_1468_375# 0 0.233029f
C19301 FILLER_0_20_15/a_1020_375# 0 0.171606f
C19302 FILLER_0_20_15/a_572_375# 0 0.171606f
C19303 FILLER_0_20_15/a_124_375# 0 0.185399f
C19304 _204_/a_67_603# 0 0.345683f
C19305 _419_/a_2560_156# 0 0.016968f
C19306 _419_/a_2665_112# 0 0.62251f
C19307 _419_/a_2248_156# 0 0.371662f
C19308 _419_/a_1204_472# 0 0.012971f
C19309 _419_/a_1000_472# 0 0.291735f
C19310 _419_/a_796_472# 0 0.023206f
C19311 _419_/a_1308_423# 0 0.279043f
C19312 _419_/a_448_472# 0 0.684413f
C19313 _419_/a_36_151# 0 1.43589f
C19314 _054_ 0 0.522819f
C19315 _221_/a_36_160# 0 0.386641f
C19316 FILLER_0_9_270/a_484_472# 0 0.345058f
C19317 FILLER_0_9_270/a_36_472# 0 0.404746f
C19318 FILLER_0_9_270/a_572_375# 0 0.232991f
C19319 FILLER_0_9_270/a_124_375# 0 0.185089f
C19320 FILLER_0_1_192/a_36_472# 0 0.417394f
C19321 FILLER_0_1_192/a_124_375# 0 0.246306f
C19322 FILLER_0_13_80/a_36_472# 0 0.417394f
C19323 FILLER_0_13_80/a_124_375# 0 0.246306f
C19324 _153_ 0 1.165862f
C19325 _154_ 0 1.167112f
C19326 _367_/a_36_68# 0 0.150048f
C19327 _436_/a_2560_156# 0 0.016968f
C19328 _436_/a_2665_112# 0 0.62251f
C19329 _436_/a_2248_156# 0 0.371662f
C19330 _436_/a_1204_472# 0 0.012971f
C19331 _436_/a_1000_472# 0 0.291735f
C19332 _436_/a_796_472# 0 0.023206f
C19333 _436_/a_1308_423# 0 0.279043f
C19334 _436_/a_448_472# 0 0.684413f
C19335 _436_/a_36_151# 0 1.43589f
C19336 FILLER_0_10_107/a_484_472# 0 0.345058f
C19337 FILLER_0_10_107/a_36_472# 0 0.404746f
C19338 FILLER_0_10_107/a_572_375# 0 0.232991f
C19339 FILLER_0_10_107/a_124_375# 0 0.185089f
C19340 _168_ 0 0.336537f
C19341 net51 0 2.105066f
C19342 _042_ 0 0.323587f
C19343 _453_/a_2560_156# 0 0.016968f
C19344 _453_/a_2665_112# 0 0.62251f
C19345 _453_/a_2248_156# 0 0.371662f
C19346 _453_/a_1204_472# 0 0.012971f
C19347 _453_/a_1000_472# 0 0.291735f
C19348 _453_/a_796_472# 0 0.023206f
C19349 _453_/a_1308_423# 0 0.279043f
C19350 _453_/a_448_472# 0 0.684413f
C19351 _453_/a_36_151# 0 1.43589f
C19352 FILLER_0_19_142/a_36_472# 0 0.417394f
C19353 FILLER_0_19_142/a_124_375# 0 0.246306f
C19354 _048_ 0 0.358805f
C19355 _205_/a_36_160# 0 0.696445f
C19356 net43 0 1.236377f
C19357 FILLER_0_3_78/a_484_472# 0 0.345058f
C19358 FILLER_0_3_78/a_36_472# 0 0.404746f
C19359 FILLER_0_3_78/a_572_375# 0 0.232991f
C19360 FILLER_0_3_78/a_124_375# 0 0.185089f
C19361 _437_/a_2560_156# 0 0.016968f
C19362 _437_/a_2665_112# 0 0.62251f
C19363 _437_/a_2248_156# 0 0.371662f
C19364 _437_/a_1204_472# 0 0.012971f
C19365 _437_/a_1000_472# 0 0.291735f
C19366 _437_/a_796_472# 0 0.023206f
C19367 _437_/a_1308_423# 0 0.279043f
C19368 _437_/a_448_472# 0 0.684413f
C19369 _437_/a_36_151# 0 1.43589f
C19370 _109_ 0 0.319326f
C19371 _299_/a_36_472# 0 0.031137f
C19372 net37 0 1.529713f
C19373 _385_/a_36_68# 0 0.112263f
C19374 FILLER_0_0_266/a_36_472# 0 0.417394f
C19375 FILLER_0_0_266/a_124_375# 0 0.246306f
C19376 net12 0 1.263595f
C19377 net22 0 2.108509f
C19378 FILLER_0_9_290/a_36_472# 0 0.417394f
C19379 FILLER_0_9_290/a_124_375# 0 0.246306f
C19380 _223_/a_36_160# 0 0.696445f
C19381 FILLER_0_14_263/a_36_472# 0 0.417394f
C19382 FILLER_0_14_263/a_124_375# 0 0.246306f
C19383 _158_ 0 0.309522f
C19384 _369_/a_36_68# 0 0.150048f
C19385 net71 0 1.420869f
C19386 _438_/a_2560_156# 0 0.016968f
C19387 _438_/a_2665_112# 0 0.62251f
C19388 _438_/a_2248_156# 0 0.371662f
C19389 _438_/a_1204_472# 0 0.012971f
C19390 _438_/a_1000_472# 0 0.291735f
C19391 _438_/a_796_472# 0 0.023206f
C19392 _438_/a_1308_423# 0 0.279043f
C19393 _438_/a_448_472# 0 0.684413f
C19394 _438_/a_36_151# 0 1.43589f
C19395 FILLER_0_23_274/a_36_472# 0 0.417394f
C19396 FILLER_0_23_274/a_124_375# 0 0.246306f
C19397 FILLER_0_17_282/a_36_472# 0 0.417394f
C19398 FILLER_0_17_282/a_124_375# 0 0.246306f
C19399 FILLER_0_5_198/a_484_472# 0 0.345058f
C19400 FILLER_0_5_198/a_36_472# 0 0.404746f
C19401 FILLER_0_5_198/a_572_375# 0 0.232991f
C19402 FILLER_0_5_198/a_124_375# 0 0.185089f
C19403 _163_ 0 1.03762f
C19404 _169_ 0 0.245383f
C19405 _386_/a_848_380# 0 0.40208f
C19406 _386_/a_124_24# 0 0.591898f
C19407 FILLER_0_20_2/a_484_472# 0 0.345058f
C19408 FILLER_0_20_2/a_36_472# 0 0.404746f
C19409 FILLER_0_20_2/a_572_375# 0 0.232991f
C19410 FILLER_0_20_2/a_124_375# 0 0.185089f
C19411 FILLER_0_16_154/a_1380_472# 0 0.345058f
C19412 FILLER_0_16_154/a_932_472# 0 0.33241f
C19413 FILLER_0_16_154/a_484_472# 0 0.33241f
C19414 FILLER_0_16_154/a_36_472# 0 0.404746f
C19415 FILLER_0_16_154/a_1468_375# 0 0.233029f
C19416 FILLER_0_16_154/a_1020_375# 0 0.171606f
C19417 FILLER_0_16_154/a_572_375# 0 0.171606f
C19418 FILLER_0_16_154/a_124_375# 0 0.185399f
C19419 FILLER_0_0_232/a_36_472# 0 0.417394f
C19420 FILLER_0_0_232/a_124_375# 0 0.246306f
C19421 FILLER_0_19_195/a_36_472# 0 0.417394f
C19422 FILLER_0_19_195/a_124_375# 0 0.246306f
C19423 _049_ 0 0.329957f
C19424 net33 0 1.934915f
C19425 _207_/a_67_603# 0 0.345683f
C19426 FILLER_0_3_54/a_36_472# 0 0.417394f
C19427 FILLER_0_3_54/a_124_375# 0 0.246306f
C19428 FILLER_0_2_101/a_36_472# 0 0.417394f
C19429 FILLER_0_2_101/a_124_375# 0 0.246306f
C19430 trim_mask\[0\] 0 0.605753f
C19431 _439_/a_2560_156# 0 0.016968f
C19432 _439_/a_2665_112# 0 0.62251f
C19433 _439_/a_2248_156# 0 0.371662f
C19434 _439_/a_1204_472# 0 0.012971f
C19435 _439_/a_1000_472# 0 0.291735f
C19436 _439_/a_796_472# 0 0.023206f
C19437 _439_/a_1308_423# 0 0.279043f
C19438 _439_/a_448_472# 0 0.684413f
C19439 _439_/a_36_151# 0 1.43589f
C19440 _066_ 0 0.333041f
C19441 FILLER_0_23_44/a_1380_472# 0 0.345058f
C19442 FILLER_0_23_44/a_932_472# 0 0.33241f
C19443 FILLER_0_23_44/a_484_472# 0 0.33241f
C19444 FILLER_0_23_44/a_36_472# 0 0.404746f
C19445 FILLER_0_23_44/a_1468_375# 0 0.233029f
C19446 FILLER_0_23_44/a_1020_375# 0 0.171606f
C19447 FILLER_0_23_44/a_572_375# 0 0.171606f
C19448 FILLER_0_23_44/a_124_375# 0 0.185399f
C19449 FILLER_0_23_88/a_36_472# 0 0.417394f
C19450 FILLER_0_23_88/a_124_375# 0 0.246306f
C19451 FILLER_0_5_164/a_484_472# 0 0.345058f
C19452 FILLER_0_5_164/a_36_472# 0 0.404746f
C19453 FILLER_0_5_164/a_572_375# 0 0.232991f
C19454 FILLER_0_5_164/a_124_375# 0 0.185089f
C19455 _060_ 0 2.485177f
C19456 _113_ 0 2.833205f
C19457 _090_ 0 2.629271f
C19458 _310_/a_49_472# 0 0.098072f
C19459 _037_ 0 0.467089f
C19460 _170_ 0 0.413995f
C19461 _387_/a_36_113# 0 0.418095f
C19462 _208_/a_36_160# 0 0.696445f
C19463 FILLER_0_18_76/a_484_472# 0 0.345058f
C19464 FILLER_0_18_76/a_36_472# 0 0.404746f
C19465 FILLER_0_18_76/a_572_375# 0 0.232991f
C19466 FILLER_0_18_76/a_124_375# 0 0.185089f
C19467 _225_/a_36_160# 0 0.386641f
C19468 FILLER_0_2_177/a_484_472# 0 0.345058f
C19469 FILLER_0_2_177/a_36_472# 0 0.404746f
C19470 FILLER_0_2_177/a_572_375# 0 0.232991f
C19471 FILLER_0_2_177/a_124_375# 0 0.185089f
C19472 FILLER_0_2_111/a_1380_472# 0 0.345058f
C19473 FILLER_0_2_111/a_932_472# 0 0.33241f
C19474 FILLER_0_2_111/a_484_472# 0 0.33241f
C19475 FILLER_0_2_111/a_36_472# 0 0.404746f
C19476 FILLER_0_2_111/a_1468_375# 0 0.233029f
C19477 FILLER_0_2_111/a_1020_375# 0 0.171606f
C19478 FILLER_0_2_111/a_572_375# 0 0.171606f
C19479 FILLER_0_2_111/a_124_375# 0 0.185399f
C19480 FILLER_0_15_228/a_36_472# 0 0.417394f
C19481 FILLER_0_15_228/a_124_375# 0 0.246306f
C19482 net47 0 2.314376f
C19483 _242_/a_36_160# 0 0.696445f
C19484 _117_ 0 1.266251f
C19485 _311_/a_66_473# 0 0.11665f
C19486 _043_ 0 0.487279f
C19487 _190_/a_36_160# 0 0.696445f
C19488 FILLER_0_9_105/a_484_472# 0 0.345058f
C19489 FILLER_0_9_105/a_36_472# 0 0.404746f
C19490 FILLER_0_9_105/a_572_375# 0 0.232991f
C19491 FILLER_0_9_105/a_124_375# 0 0.185089f
C19492 FILLER_0_13_100/a_36_472# 0 0.417394f
C19493 FILLER_0_13_100/a_124_375# 0 0.246306f
C19494 FILLER_0_22_177/a_1380_472# 0 0.345058f
C19495 FILLER_0_22_177/a_932_472# 0 0.33241f
C19496 FILLER_0_22_177/a_484_472# 0 0.33241f
C19497 FILLER_0_22_177/a_36_472# 0 0.404746f
C19498 FILLER_0_22_177/a_1468_375# 0 0.233029f
C19499 FILLER_0_22_177/a_1020_375# 0 0.171606f
C19500 FILLER_0_22_177/a_572_375# 0 0.171606f
C19501 FILLER_0_22_177/a_124_375# 0 0.185399f
C19502 FILLER_0_15_2/a_484_472# 0 0.345058f
C19503 FILLER_0_15_2/a_36_472# 0 0.404746f
C19504 FILLER_0_15_2/a_572_375# 0 0.232991f
C19505 FILLER_0_15_2/a_124_375# 0 0.185089f
C19506 FILLER_0_15_10/a_36_472# 0 0.417394f
C19507 FILLER_0_15_10/a_124_375# 0 0.246306f
C19508 FILLER_0_19_171/a_1380_472# 0 0.345058f
C19509 FILLER_0_19_171/a_932_472# 0 0.33241f
C19510 FILLER_0_19_171/a_484_472# 0 0.33241f
C19511 FILLER_0_19_171/a_36_472# 0 0.404746f
C19512 FILLER_0_19_171/a_1468_375# 0 0.233029f
C19513 FILLER_0_19_171/a_1020_375# 0 0.171606f
C19514 FILLER_0_19_171/a_572_375# 0 0.171606f
C19515 FILLER_0_19_171/a_124_375# 0 0.185399f
C19516 net13 0 1.176306f
C19517 net23 0 2.091399f
C19518 FILLER_0_20_87/a_36_472# 0 0.417394f
C19519 FILLER_0_20_87/a_124_375# 0 0.246306f
C19520 FILLER_0_20_98/a_36_472# 0 0.417394f
C19521 FILLER_0_20_98/a_124_375# 0 0.246306f
C19522 _055_ 0 1.782885f
C19523 FILLER_0_18_53/a_484_472# 0 0.345058f
C19524 FILLER_0_18_53/a_36_472# 0 0.404746f
C19525 FILLER_0_18_53/a_572_375# 0 0.232991f
C19526 FILLER_0_18_53/a_124_375# 0 0.185089f
C19527 FILLER_0_2_165/a_36_472# 0 0.417394f
C19528 FILLER_0_2_165/a_124_375# 0 0.246306f
C19529 FILLER_0_15_205/a_36_472# 0 0.417394f
C19530 FILLER_0_15_205/a_124_375# 0 0.246306f
C19531 FILLER_0_23_282/a_484_472# 0 0.345058f
C19532 FILLER_0_23_282/a_36_472# 0 0.404746f
C19533 FILLER_0_23_282/a_572_375# 0 0.232991f
C19534 FILLER_0_23_282/a_124_375# 0 0.185089f
C19535 net42 0 1.067446f
C19536 net17 0 2.210219f
C19537 _172_ 0 0.265782f
C19538 _171_ 0 0.300355f
C19539 _389_/a_36_148# 0 0.388358f
C19540 _080_ 0 0.328202f
C19541 _260_/a_36_68# 0 0.112263f
C19542 FILLER_0_0_96/a_36_472# 0 0.417394f
C19543 FILLER_0_0_96/a_124_375# 0 0.246306f
C19544 FILLER_0_9_72/a_1380_472# 0 0.345058f
C19545 FILLER_0_9_72/a_932_472# 0 0.33241f
C19546 FILLER_0_9_72/a_484_472# 0 0.33241f
C19547 FILLER_0_9_72/a_36_472# 0 0.404746f
C19548 FILLER_0_9_72/a_1468_375# 0 0.233029f
C19549 FILLER_0_9_72/a_1020_375# 0 0.171606f
C19550 FILLER_0_9_72/a_572_375# 0 0.171606f
C19551 FILLER_0_9_72/a_124_375# 0 0.185399f
C19552 FILLER_0_20_31/a_36_472# 0 0.417394f
C19553 FILLER_0_20_31/a_124_375# 0 0.246306f
C19554 _227_/a_36_160# 0 0.386641f
C19555 _120_ 0 1.533088f
C19556 _313_/a_67_603# 0 0.345683f
C19557 FILLER_0_5_172/a_36_472# 0 0.417394f
C19558 FILLER_0_5_172/a_124_375# 0 0.246306f
C19559 FILLER_0_12_20/a_484_472# 0 0.345058f
C19560 FILLER_0_12_20/a_36_472# 0 0.404746f
C19561 FILLER_0_12_20/a_572_375# 0 0.232991f
C19562 FILLER_0_12_20/a_124_375# 0 0.185089f
C19563 _134_ 0 0.365972f
C19564 _062_ 0 1.717773f
C19565 _059_ 0 1.686761f
C19566 _261_/a_36_160# 0 0.386641f
C19567 _044_ 0 0.388801f
C19568 mask\[1\] 0 1.295078f
C19569 _192_/a_67_603# 0 0.345683f
C19570 FILLER_0_13_142/a_1380_472# 0 0.345058f
C19571 FILLER_0_13_142/a_932_472# 0 0.33241f
C19572 FILLER_0_13_142/a_484_472# 0 0.33241f
C19573 FILLER_0_13_142/a_36_472# 0 0.404746f
C19574 FILLER_0_13_142/a_1468_375# 0 0.233029f
C19575 FILLER_0_13_142/a_1020_375# 0 0.171606f
C19576 FILLER_0_13_142/a_572_375# 0 0.171606f
C19577 FILLER_0_13_142/a_124_375# 0 0.185399f
C19578 FILLER_0_9_60/a_484_472# 0 0.345058f
C19579 FILLER_0_9_60/a_36_472# 0 0.404746f
C19580 FILLER_0_9_60/a_572_375# 0 0.232991f
C19581 FILLER_0_9_60/a_124_375# 0 0.185089f
C19582 FILLER_0_7_233/a_36_472# 0 0.417394f
C19583 FILLER_0_7_233/a_124_375# 0 0.246306f
C19584 _228_/a_36_68# 0 0.69549f
C19585 FILLER_0_21_206/a_36_472# 0 0.417394f
C19586 FILLER_0_21_206/a_124_375# 0 0.246306f
C19587 _067_ 0 0.851951f
C19588 _135_ 0 0.339478f
C19589 _193_/a_36_160# 0 0.696445f
C19590 _180_ 0 0.390598f
C19591 cal_count\[1\] 0 1.568289f
C19592 FILLER_0_4_213/a_484_472# 0 0.345058f
C19593 FILLER_0_4_213/a_36_472# 0 0.404746f
C19594 FILLER_0_4_213/a_572_375# 0 0.232991f
C19595 FILLER_0_4_213/a_124_375# 0 0.185089f
C19596 FILLER_0_11_282/a_36_472# 0 0.417394f
C19597 FILLER_0_11_282/a_124_375# 0 0.246306f
C19598 FILLER_0_18_61/a_36_472# 0 0.417394f
C19599 FILLER_0_18_61/a_124_375# 0 0.246306f
C19600 FILLER_0_15_235/a_484_472# 0 0.345058f
C19601 FILLER_0_15_235/a_36_472# 0 0.404746f
C19602 FILLER_0_15_235/a_572_375# 0 0.232991f
C19603 FILLER_0_15_235/a_124_375# 0 0.185089f
C19604 FILLER_0_23_290/a_36_472# 0 0.417394f
C19605 FILLER_0_23_290/a_124_375# 0 0.246306f
C19606 _121_ 0 0.532847f
C19607 _315_/a_36_68# 0 0.052951f
C19608 _246_/a_36_68# 0 0.69549f
C19609 FILLER_0_5_181/a_36_472# 0 0.417394f
C19610 FILLER_0_5_181/a_124_375# 0 0.246306f
C19611 _082_ 0 0.619901f
C19612 net8 0 1.163723f
C19613 net18 0 2.032159f
C19614 _332_/a_36_472# 0 0.031137f
C19615 _179_ 0 0.336984f
C19616 _401_/a_36_68# 0 0.112263f
C19617 FILLER_0_14_107/a_1380_472# 0 0.345058f
C19618 FILLER_0_14_107/a_932_472# 0 0.33241f
C19619 FILLER_0_14_107/a_484_472# 0 0.33241f
C19620 FILLER_0_14_107/a_36_472# 0 0.404746f
C19621 FILLER_0_14_107/a_1468_375# 0 0.233029f
C19622 FILLER_0_14_107/a_1020_375# 0 0.171606f
C19623 FILLER_0_14_107/a_572_375# 0 0.171606f
C19624 FILLER_0_14_107/a_124_375# 0 0.185399f
C19625 _097_ 0 0.592554f
C19626 FILLER_0_1_204/a_36_472# 0 0.417394f
C19627 FILLER_0_1_204/a_124_375# 0 0.246306f
C19628 FILLER_0_15_72/a_484_472# 0 0.345058f
C19629 FILLER_0_15_72/a_36_472# 0 0.404746f
C19630 FILLER_0_15_72/a_572_375# 0 0.232991f
C19631 FILLER_0_15_72/a_124_375# 0 0.185089f
C19632 FILLER_0_17_104/a_1380_472# 0 0.345058f
C19633 FILLER_0_17_104/a_932_472# 0 0.33241f
C19634 FILLER_0_17_104/a_484_472# 0 0.33241f
C19635 FILLER_0_17_104/a_36_472# 0 0.404746f
C19636 FILLER_0_17_104/a_1468_375# 0 0.233029f
C19637 FILLER_0_17_104/a_1020_375# 0 0.171606f
C19638 FILLER_0_17_104/a_572_375# 0 0.171606f
C19639 FILLER_0_17_104/a_124_375# 0 0.185399f
C19640 FILLER_0_8_37/a_484_472# 0 0.345058f
C19641 FILLER_0_8_37/a_36_472# 0 0.404746f
C19642 FILLER_0_8_37/a_572_375# 0 0.232991f
C19643 FILLER_0_8_37/a_124_375# 0 0.185089f
C19644 FILLER_0_15_212/a_1380_472# 0 0.345058f
C19645 FILLER_0_15_212/a_932_472# 0 0.33241f
C19646 FILLER_0_15_212/a_484_472# 0 0.33241f
C19647 FILLER_0_15_212/a_36_472# 0 0.404746f
C19648 FILLER_0_15_212/a_1468_375# 0 0.233029f
C19649 FILLER_0_15_212/a_1020_375# 0 0.171606f
C19650 FILLER_0_15_212/a_572_375# 0 0.171606f
C19651 FILLER_0_15_212/a_124_375# 0 0.185399f
C19652 FILLER_0_23_60/a_36_472# 0 0.417394f
C19653 FILLER_0_23_60/a_124_375# 0 0.246306f
C19654 _123_ 0 0.344874f
C19655 _122_ 0 0.600118f
C19656 calibrate 0 1.343796f
C19657 _316_/a_848_380# 0 0.40208f
C19658 _316_/a_124_24# 0 0.591898f
C19659 _247_/a_36_160# 0 0.696445f
C19660 FILLER_0_12_50/a_36_472# 0 0.417394f
C19661 FILLER_0_12_50/a_124_375# 0 0.246306f
C19662 _084_ 0 0.296163f
C19663 cal_itt\[0\] 0 1.831055f
C19664 cal_itt\[1\] 0 1.705665f
C19665 FILLER_0_11_109/a_36_472# 0 0.417394f
C19666 FILLER_0_11_109/a_124_375# 0 0.246306f
C19667 _182_ 0 0.34197f
C19668 _402_/a_1948_68# 0 0.022025f
C19669 _402_/a_718_527# 0 0.001795f
C19670 _402_/a_56_567# 0 0.424713f
C19671 _402_/a_728_93# 0 0.65929f
C19672 _402_/a_1296_93# 0 0.317801f
C19673 _045_ 0 0.349338f
C19674 mask\[2\] 0 1.335688f
C19675 _195_/a_67_603# 0 0.345683f
C19676 _333_/a_36_160# 0 0.386641f
C19677 _098_ 0 1.816151f
C19678 _147_ 0 0.322539f
C19679 _350_/a_49_472# 0 0.054843f
C19680 FILLER_0_12_236/a_484_472# 0 0.345058f
C19681 FILLER_0_12_236/a_36_472# 0 0.404746f
C19682 FILLER_0_12_236/a_572_375# 0 0.232991f
C19683 FILLER_0_12_236/a_124_375# 0 0.185089f
C19684 FILLER_0_2_171/a_36_472# 0 0.417394f
C19685 FILLER_0_2_171/a_124_375# 0 0.246306f
C19686 _014_ 0 0.363432f
C19687 _317_/a_36_113# 0 0.418095f
C19688 _248_/a_36_68# 0 0.69549f
C19689 FILLER_0_17_38/a_484_472# 0 0.345058f
C19690 FILLER_0_17_38/a_36_472# 0 0.404746f
C19691 FILLER_0_17_38/a_572_375# 0 0.232991f
C19692 FILLER_0_17_38/a_124_375# 0 0.185089f
C19693 _001_ 0 0.285216f
C19694 _265_/a_244_68# 0 0.138666f
C19695 _196_/a_36_160# 0 0.696445f
C19696 FILLER_0_6_90/a_484_472# 0 0.345058f
C19697 FILLER_0_6_90/a_36_472# 0 0.404746f
C19698 FILLER_0_6_90/a_572_375# 0 0.232991f
C19699 FILLER_0_6_90/a_124_375# 0 0.185089f
C19700 _183_ 0 0.356629f
C19701 _334_/a_36_160# 0 0.386641f
C19702 _282_/a_36_160# 0 0.386641f
C19703 _024_ 0 0.451815f
C19704 _009_ 0 0.397943f
C19705 _420_/a_2560_156# 0 0.016968f
C19706 _420_/a_2665_112# 0 0.62251f
C19707 _420_/a_2248_156# 0 0.371662f
C19708 _420_/a_1204_472# 0 0.012971f
C19709 _420_/a_1000_472# 0 0.291735f
C19710 _420_/a_796_472# 0 0.023206f
C19711 _420_/a_1308_423# 0 0.279043f
C19712 _420_/a_448_472# 0 0.684413f
C19713 _420_/a_36_151# 0 1.43589f
C19714 clk 0 1.162312f
C19715 FILLER_0_8_2/a_36_472# 0 0.417394f
C19716 FILLER_0_8_2/a_124_375# 0 0.246306f
C19717 FILLER_0_8_24/a_484_472# 0 0.345058f
C19718 FILLER_0_8_24/a_36_472# 0 0.404746f
C19719 FILLER_0_8_24/a_572_375# 0 0.232991f
C19720 FILLER_0_8_24/a_124_375# 0 0.185089f
C19721 _124_ 0 0.294081f
C19722 _118_ 0 1.378735f
C19723 _071_ 0 1.600488f
C19724 net9 0 1.13171f
C19725 net19 0 1.889339f
C19726 _138_ 0 0.33132f
C19727 _137_ 0 1.178616f
C19728 _335_/a_49_472# 0 0.054843f
C19729 _404_/a_36_472# 0 0.031137f
C19730 FILLER_0_20_107/a_36_472# 0 0.417394f
C19731 FILLER_0_20_107/a_124_375# 0 0.246306f
C19732 FILLER_0_9_142/a_36_472# 0 0.417394f
C19733 FILLER_0_9_142/a_124_375# 0 0.246306f
C19734 _099_ 0 1.152785f
C19735 _283_/a_36_472# 0 0.031137f
C19736 mask\[7\] 0 1.477838f
C19737 _352_/a_49_472# 0 0.054843f
C19738 _010_ 0 0.377779f
C19739 _421_/a_2560_156# 0 0.016968f
C19740 _421_/a_2665_112# 0 0.62251f
C19741 _421_/a_2248_156# 0 0.371662f
C19742 _421_/a_1204_472# 0 0.012971f
C19743 _421_/a_1000_472# 0 0.291735f
C19744 _421_/a_796_472# 0 0.023206f
C19745 _421_/a_1308_423# 0 0.279043f
C19746 _421_/a_448_472# 0 0.684413f
C19747 _421_/a_36_151# 0 1.43589f
C19748 FILLER_0_1_212/a_36_472# 0 0.417394f
C19749 FILLER_0_1_212/a_124_375# 0 0.246306f
C19750 FILLER_0_8_239/a_36_472# 0 0.417394f
C19751 FILLER_0_8_239/a_124_375# 0 0.246306f
C19752 _125_ 0 1.526603f
C19753 _058_ 0 1.483584f
C19754 FILLER_0_6_177/a_484_472# 0 0.345058f
C19755 FILLER_0_6_177/a_36_472# 0 0.404746f
C19756 FILLER_0_6_177/a_572_375# 0 0.232991f
C19757 FILLER_0_6_177/a_124_375# 0 0.185089f
C19758 state\[1\] 0 2.652405f
C19759 _267_/a_36_472# 0 0.137725f
C19760 _184_ 0 0.350066f
C19761 cal_count\[2\] 0 1.971854f
C19762 _405_/a_67_603# 0 0.345683f
C19763 _018_ 0 0.358633f
C19764 _046_ 0 0.361963f
C19765 _198_/a_67_603# 0 0.345683f
C19766 _094_ 0 1.263877f
C19767 _100_ 0 0.333135f
C19768 net36 0 2.262756f
C19769 FILLER_0_17_133/a_36_472# 0 0.417394f
C19770 FILLER_0_17_133/a_124_375# 0 0.246306f
C19771 _025_ 0 0.350324f
C19772 _148_ 0 0.325709f
C19773 _422_/a_2560_156# 0 0.016968f
C19774 _422_/a_2665_112# 0 0.62251f
C19775 _422_/a_2248_156# 0 0.371662f
C19776 _422_/a_1204_472# 0 0.012971f
C19777 _422_/a_1000_472# 0 0.291735f
C19778 _422_/a_796_472# 0 0.023206f
C19779 _422_/a_1308_423# 0 0.279043f
C19780 _422_/a_448_472# 0 0.684413f
C19781 _422_/a_36_151# 0 1.43589f
C19782 FILLER_0_1_266/a_484_472# 0 0.345058f
C19783 FILLER_0_1_266/a_36_472# 0 0.404746f
C19784 FILLER_0_1_266/a_572_375# 0 0.232991f
C19785 FILLER_0_1_266/a_124_375# 0 0.185089f
C19786 _152_ 0 0.918583f
C19787 _081_ 0 1.140656f
C19788 _370_/a_848_380# 0 0.40208f
C19789 _370_/a_124_24# 0 0.591898f
C19790 FILLER_0_24_274/a_1380_472# 0 0.345058f
C19791 FILLER_0_24_274/a_932_472# 0 0.33241f
C19792 FILLER_0_24_274/a_484_472# 0 0.33241f
C19793 FILLER_0_24_274/a_36_472# 0 0.404746f
C19794 FILLER_0_24_274/a_1468_375# 0 0.233029f
C19795 FILLER_0_24_274/a_1020_375# 0 0.171606f
C19796 FILLER_0_24_274/a_572_375# 0 0.171606f
C19797 FILLER_0_24_274/a_124_375# 0 0.185399f
C19798 _185_ 0 0.386917f
C19799 _406_/a_36_159# 0 0.374116f
C19800 _337_/a_49_472# 0 0.054843f
C19801 _199_/a_36_160# 0 0.696445f
C19802 _285_/a_36_472# 0 0.031137f
C19803 _354_/a_49_472# 0 0.054843f
C19804 _012_ 0 0.75195f
C19805 _423_/a_2560_156# 0 0.016968f
C19806 _423_/a_2665_112# 0 0.62251f
C19807 _423_/a_2248_156# 0 0.371662f
C19808 _423_/a_1204_472# 0 0.012971f
C19809 _423_/a_1000_472# 0 0.291735f
C19810 _423_/a_796_472# 0 0.023206f
C19811 _423_/a_1308_423# 0 0.279043f
C19812 _423_/a_448_472# 0 0.684413f
C19813 _423_/a_36_151# 0 1.43589f
C19814 FILLER_0_5_88/a_36_472# 0 0.417394f
C19815 FILLER_0_5_88/a_124_375# 0 0.246306f
C19816 trim_mask\[1\] 0 1.020743f
C19817 _029_ 0 0.308904f
C19818 _440_/a_2560_156# 0 0.016968f
C19819 _440_/a_2665_112# 0 0.62251f
C19820 _440_/a_2248_156# 0 0.371662f
C19821 _440_/a_1204_472# 0 0.012971f
C19822 _440_/a_1000_472# 0 0.291735f
C19823 _440_/a_796_472# 0 0.023206f
C19824 _440_/a_1308_423# 0 0.279043f
C19825 _440_/a_448_472# 0 0.684413f
C19826 _440_/a_36_151# 0 1.43589f
C19827 _159_ 0 0.351814f
C19828 _371_/a_36_113# 0 0.418095f
C19829 FILLER_0_17_56/a_484_472# 0 0.345058f
C19830 FILLER_0_17_56/a_36_472# 0 0.404746f
C19831 FILLER_0_17_56/a_572_375# 0 0.232991f
C19832 FILLER_0_17_56/a_124_375# 0 0.185089f
C19833 _083_ 0 0.527882f
C19834 _078_ 0 0.904554f
C19835 _269_/a_36_472# 0 0.031137f
C19836 _181_ 0 0.829168f
C19837 _407_/a_36_472# 0 0.031137f
C19838 _019_ 0 0.32907f
C19839 _139_ 0 0.346404f
C19840 FILLER_0_14_123/a_36_472# 0 0.417394f
C19841 FILLER_0_14_123/a_124_375# 0 0.246306f
C19842 _005_ 0 0.340993f
C19843 _101_ 0 0.280497f
C19844 _424_/a_2560_156# 0 0.016968f
C19845 _424_/a_2665_112# 0 0.62251f
C19846 _424_/a_2248_156# 0 0.371662f
C19847 _424_/a_1204_472# 0 0.012971f
C19848 _424_/a_1000_472# 0 0.291735f
C19849 _424_/a_796_472# 0 0.023206f
C19850 _424_/a_1308_423# 0 0.279043f
C19851 _424_/a_448_472# 0 0.684413f
C19852 _424_/a_36_151# 0 1.43589f
C19853 _026_ 0 0.320379f
C19854 _149_ 0 0.305496f
C19855 FILLER_0_5_54/a_1380_472# 0 0.345058f
C19856 FILLER_0_5_54/a_932_472# 0 0.33241f
C19857 FILLER_0_5_54/a_484_472# 0 0.33241f
C19858 FILLER_0_5_54/a_36_472# 0 0.404746f
C19859 FILLER_0_5_54/a_1468_375# 0 0.233029f
C19860 FILLER_0_5_54/a_1020_375# 0 0.171606f
C19861 FILLER_0_5_54/a_572_375# 0 0.171606f
C19862 FILLER_0_5_54/a_124_375# 0 0.185399f
C19863 FILLER_0_17_142/a_484_472# 0 0.345058f
C19864 FILLER_0_17_142/a_36_472# 0 0.404746f
C19865 FILLER_0_17_142/a_572_375# 0 0.232991f
C19866 FILLER_0_17_142/a_124_375# 0 0.185089f
C19867 _068_ 0 3.162692f
C19868 _076_ 0 3.812442f
C19869 _133_ 0 1.430901f
C19870 _070_ 0 3.115722f
C19871 _372_/a_170_472# 0 0.077257f
C19872 net49 0 5.140563f
C19873 _030_ 0 0.307083f
C19874 net66 0 1.472669f
C19875 _441_/a_2560_156# 0 0.016968f
C19876 _441_/a_2665_112# 0 0.62251f
C19877 _441_/a_2248_156# 0 0.371662f
C19878 _441_/a_1204_472# 0 0.012971f
C19879 _441_/a_1000_472# 0 0.291735f
C19880 _441_/a_796_472# 0 0.023206f
C19881 _441_/a_1308_423# 0 0.279043f
C19882 _441_/a_448_472# 0 0.684413f
C19883 _441_/a_36_151# 0 1.43589f
C19884 FILLER_0_5_206/a_36_472# 0 0.417394f
C19885 FILLER_0_5_206/a_124_375# 0 0.246306f
C19886 fanout49/a_36_160# 0 0.696445f
C19887 FILLER_0_8_247/a_1380_472# 0 0.345058f
C19888 FILLER_0_8_247/a_932_472# 0 0.33241f
C19889 FILLER_0_8_247/a_484_472# 0 0.33241f
C19890 FILLER_0_8_247/a_36_472# 0 0.404746f
C19891 FILLER_0_8_247/a_1468_375# 0 0.233029f
C19892 FILLER_0_8_247/a_1020_375# 0 0.171606f
C19893 FILLER_0_8_247/a_572_375# 0 0.171606f
C19894 FILLER_0_8_247/a_124_375# 0 0.185399f
C19895 FILLER_0_12_220/a_1380_472# 0 0.345058f
C19896 FILLER_0_12_220/a_932_472# 0 0.33241f
C19897 FILLER_0_12_220/a_484_472# 0 0.33241f
C19898 FILLER_0_12_220/a_36_472# 0 0.404746f
C19899 FILLER_0_12_220/a_1468_375# 0 0.233029f
C19900 FILLER_0_12_220/a_1020_375# 0 0.171606f
C19901 FILLER_0_12_220/a_572_375# 0 0.171606f
C19902 FILLER_0_12_220/a_124_375# 0 0.185399f
C19903 FILLER_0_21_286/a_484_472# 0 0.345058f
C19904 FILLER_0_21_286/a_36_472# 0 0.404746f
C19905 FILLER_0_21_286/a_572_375# 0 0.232991f
C19906 FILLER_0_21_286/a_124_375# 0 0.185089f
C19907 _140_ 0 1.276518f
C19908 _339_/a_36_160# 0 0.386641f
C19909 _095_ 0 2.689027f
C19910 _186_ 0 0.580923f
C19911 _408_/a_1936_472# 0 0.009918f
C19912 _408_/a_718_524# 0 0.005143f
C19913 _408_/a_56_524# 0 0.41096f
C19914 _408_/a_728_93# 0 0.654825f
C19915 _408_/a_1336_472# 0 0.316639f
C19916 FILLER_0_20_169/a_36_472# 0 0.417394f
C19917 FILLER_0_20_169/a_124_375# 0 0.246306f
C19918 _210_/a_67_603# 0 0.345683f
C19919 _425_/a_2560_156# 0 0.016968f
C19920 _425_/a_2665_112# 0 0.62251f
C19921 _425_/a_2248_156# 0 0.371662f
C19922 _425_/a_1204_472# 0 0.012971f
C19923 _425_/a_1000_472# 0 0.291735f
C19924 _425_/a_796_472# 0 0.023206f
C19925 _425_/a_1308_423# 0 0.279043f
C19926 _425_/a_448_472# 0 0.684413f
C19927 _425_/a_36_151# 0 1.43589f
C19928 net5 0 0.610761f
C19929 input5/a_36_113# 0 0.418095f
C19930 FILLER_0_11_78/a_484_472# 0 0.345058f
C19931 FILLER_0_11_78/a_36_472# 0 0.404746f
C19932 FILLER_0_11_78/a_572_375# 0 0.232991f
C19933 FILLER_0_11_78/a_124_375# 0 0.185089f
C19934 _102_ 0 0.335308f
C19935 _287_/a_36_472# 0 0.031137f
C19936 mask\[9\] 0 1.383606f
C19937 _356_/a_36_472# 0 0.031137f
C19938 _031_ 0 0.417351f
C19939 net69 0 1.020293f
C19940 _442_/a_2560_156# 0 0.016968f
C19941 _442_/a_2665_112# 0 0.62251f
C19942 _442_/a_2248_156# 0 0.371662f
C19943 _442_/a_1204_472# 0 0.012971f
C19944 _442_/a_1000_472# 0 0.291735f
C19945 _442_/a_796_472# 0 0.023206f
C19946 _442_/a_1308_423# 0 0.279043f
C19947 _442_/a_448_472# 0 0.684413f
C19948 _442_/a_36_151# 0 1.43589f
C19949 net64 0 2.598514f
C19950 fanout59/a_36_160# 0 0.696445f
C19951 FILLER_0_14_99/a_36_472# 0 0.417394f
C19952 FILLER_0_14_99/a_124_375# 0 0.246306f
C19953 _038_ 0 0.362839f
C19954 _136_ 0 1.345638f
C19955 _390_/a_36_68# 0 0.150048f
C19956 FILLER_0_15_282/a_484_472# 0 0.345058f
C19957 FILLER_0_15_282/a_36_472# 0 0.404746f
C19958 FILLER_0_15_282/a_572_375# 0 0.232991f
C19959 FILLER_0_15_282/a_124_375# 0 0.185089f
C19960 FILLER_0_11_124/a_36_472# 0 0.417394f
C19961 FILLER_0_11_124/a_124_375# 0 0.246306f
C19962 FILLER_0_11_135/a_36_472# 0 0.417394f
C19963 FILLER_0_11_135/a_124_375# 0 0.246306f
C19964 _188_ 0 0.349407f
C19965 cal_count\[3\] 0 1.862896f
C19966 _050_ 0 0.622354f
C19967 _211_/a_36_160# 0 0.386641f
C19968 net4 0 2.711508f
C19969 en 0 0.833743f
C19970 input4/a_36_68# 0 0.69549f
C19971 _426_/a_2560_156# 0 0.016968f
C19972 _426_/a_2665_112# 0 0.62251f
C19973 _426_/a_2248_156# 0 0.371662f
C19974 _426_/a_1204_472# 0 0.012971f
C19975 _426_/a_1000_472# 0 0.291735f
C19976 _426_/a_796_472# 0 0.023206f
C19977 _426_/a_1308_423# 0 0.279043f
C19978 _426_/a_448_472# 0 0.684413f
C19979 _426_/a_36_151# 0 1.43589f
C19980 _027_ 0 0.302949f
C19981 _150_ 0 0.320497f
C19982 FILLER_0_18_107/a_3172_472# 0 0.345058f
C19983 FILLER_0_18_107/a_2724_472# 0 0.33241f
C19984 FILLER_0_18_107/a_2276_472# 0 0.33241f
C19985 FILLER_0_18_107/a_1828_472# 0 0.33241f
C19986 FILLER_0_18_107/a_1380_472# 0 0.33241f
C19987 FILLER_0_18_107/a_932_472# 0 0.33241f
C19988 FILLER_0_18_107/a_484_472# 0 0.33241f
C19989 FILLER_0_18_107/a_36_472# 0 0.404746f
C19990 FILLER_0_18_107/a_3260_375# 0 0.233093f
C19991 FILLER_0_18_107/a_2812_375# 0 0.17167f
C19992 FILLER_0_18_107/a_2364_375# 0 0.17167f
C19993 FILLER_0_18_107/a_1916_375# 0 0.17167f
C19994 FILLER_0_18_107/a_1468_375# 0 0.17167f
C19995 FILLER_0_18_107/a_1020_375# 0 0.17167f
C19996 FILLER_0_18_107/a_572_375# 0 0.17167f
C19997 FILLER_0_18_107/a_124_375# 0 0.185915f
C19998 trim_mask\[4\] 0 0.987791f
C19999 _032_ 0 0.34876f
C20000 _443_/a_2560_156# 0 0.016968f
C20001 _443_/a_2665_112# 0 0.62251f
C20002 _443_/a_2248_156# 0 0.371662f
C20003 _443_/a_1204_472# 0 0.012971f
C20004 _443_/a_1000_472# 0 0.291735f
C20005 _443_/a_796_472# 0 0.023206f
C20006 _443_/a_1308_423# 0 0.279043f
C20007 _443_/a_448_472# 0 0.684413f
C20008 _443_/a_36_151# 0 1.43589f
C20009 _061_ 0 0.84986f
C20010 _056_ 0 2.393362f
C20011 _374_/a_36_68# 0 0.112263f
C20012 fanout58/a_36_160# 0 0.696445f
C20013 net74 0 1.237373f
C20014 fanout69/a_36_113# 0 0.418095f
C20015 _173_ 0 0.339446f
C20016 FILLER_0_3_142/a_36_472# 0 0.417394f
C20017 FILLER_0_3_142/a_124_375# 0 0.246306f
C20018 FILLER_0_17_64/a_36_472# 0 0.417394f
C20019 FILLER_0_17_64/a_124_375# 0 0.246306f
C20020 FILLER_0_11_101/a_484_472# 0 0.345058f
C20021 FILLER_0_11_101/a_36_472# 0 0.404746f
C20022 FILLER_0_11_101/a_572_375# 0 0.232991f
C20023 FILLER_0_11_101/a_124_375# 0 0.185089f
C20024 FILLER_0_22_86/a_1380_472# 0 0.345058f
C20025 FILLER_0_22_86/a_932_472# 0 0.33241f
C20026 FILLER_0_22_86/a_484_472# 0 0.33241f
C20027 FILLER_0_22_86/a_36_472# 0 0.404746f
C20028 FILLER_0_22_86/a_1468_375# 0 0.233029f
C20029 FILLER_0_22_86/a_1020_375# 0 0.171606f
C20030 FILLER_0_22_86/a_572_375# 0 0.171606f
C20031 FILLER_0_22_86/a_124_375# 0 0.185399f
C20032 net15 0 1.440851f
C20033 net24 0 1.61895f
C20034 net3 0 0.740676f
C20035 input3/a_36_113# 0 0.418095f
C20036 _103_ 0 0.350464f
C20037 _289_/a_36_472# 0 0.031137f
C20038 _151_ 0 0.300777f
C20039 _427_/a_2560_156# 0 0.016968f
C20040 _427_/a_2665_112# 0 0.91969f
C20041 _427_/a_2248_156# 0 0.30886f
C20042 _427_/a_1204_472# 0 0.012971f
C20043 _427_/a_1000_472# 0 0.291735f
C20044 _427_/a_796_472# 0 0.023206f
C20045 _427_/a_1308_423# 0 0.279043f
C20046 _427_/a_448_472# 0 0.684413f
C20047 _427_/a_36_151# 0 1.43587f
C20048 FILLER_0_17_161/a_36_472# 0 0.417394f
C20049 FILLER_0_17_161/a_124_375# 0 0.246306f
C20050 FILLER_0_18_139/a_1380_472# 0 0.345058f
C20051 FILLER_0_18_139/a_932_472# 0 0.33241f
C20052 FILLER_0_18_139/a_484_472# 0 0.33241f
C20053 FILLER_0_18_139/a_36_472# 0 0.404746f
C20054 FILLER_0_18_139/a_1468_375# 0 0.233029f
C20055 FILLER_0_18_139/a_1020_375# 0 0.171606f
C20056 FILLER_0_18_139/a_572_375# 0 0.171606f
C20057 FILLER_0_18_139/a_124_375# 0 0.185399f
C20058 _161_ 0 0.592909f
C20059 _162_ 0 0.597238f
C20060 _375_/a_36_68# 0 0.048026f
C20061 trim_val\[0\] 0 0.742779f
C20062 net67 0 1.662327f
C20063 _444_/a_2560_156# 0 0.016968f
C20064 _444_/a_2665_112# 0 0.62251f
C20065 _444_/a_2248_156# 0 0.371662f
C20066 _444_/a_1204_472# 0 0.012971f
C20067 _444_/a_1000_472# 0 0.291735f
C20068 _444_/a_796_472# 0 0.023206f
C20069 _444_/a_1308_423# 0 0.279043f
C20070 _444_/a_448_472# 0 0.684413f
C20071 _444_/a_36_151# 0 1.43589f
C20072 net65 0 0.804072f
C20073 fanout57/a_36_113# 0 0.418095f
C20074 fanout68/a_36_113# 0 0.418095f
C20075 FILLER_0_12_2/a_484_472# 0 0.345058f
C20076 FILLER_0_12_2/a_36_472# 0 0.404746f
C20077 FILLER_0_12_2/a_572_375# 0 0.232991f
C20078 FILLER_0_12_2/a_124_375# 0 0.185089f
C20079 net79 0 1.584979f
C20080 fanout79/a_36_160# 0 0.386641f
C20081 _392_/a_36_68# 0 0.112263f
C20082 FILLER_0_13_228/a_36_472# 0 0.417394f
C20083 FILLER_0_13_228/a_124_375# 0 0.246306f
C20084 FILLER_0_13_206/a_36_472# 0 0.417394f
C20085 FILLER_0_13_206/a_124_375# 0 0.246306f
C20086 FILLER_0_20_177/a_1380_472# 0 0.345058f
C20087 FILLER_0_20_177/a_932_472# 0 0.33241f
C20088 FILLER_0_20_177/a_484_472# 0 0.33241f
C20089 FILLER_0_20_177/a_36_472# 0 0.404746f
C20090 FILLER_0_20_177/a_1468_375# 0 0.233029f
C20091 FILLER_0_20_177/a_1020_375# 0 0.171606f
C20092 FILLER_0_20_177/a_572_375# 0 0.171606f
C20093 FILLER_0_20_177/a_124_375# 0 0.185399f
C20094 _051_ 0 0.349381f
C20095 _213_/a_67_603# 0 0.345683f
C20096 net2 0 0.461658f
C20097 input2/a_36_113# 0 0.418095f
C20098 _129_ 0 0.926508f
C20099 _131_ 0 1.734297f
C20100 _359_/a_36_488# 0 0.101145f
C20101 FILLER_0_11_64/a_36_472# 0 0.417394f
C20102 FILLER_0_11_64/a_124_375# 0 0.246306f
C20103 state\[2\] 0 0.607433f
C20104 net53 0 4.483899f
C20105 _017_ 0 0.334329f
C20106 net70 0 1.238296f
C20107 _428_/a_2560_156# 0 0.016968f
C20108 _428_/a_2665_112# 0 0.62251f
C20109 _428_/a_2248_156# 0 0.371662f
C20110 _428_/a_1204_472# 0 0.012971f
C20111 _428_/a_1000_472# 0 0.291735f
C20112 _428_/a_796_472# 0 0.023206f
C20113 _428_/a_1308_423# 0 0.279043f
C20114 _428_/a_448_472# 0 0.684413f
C20115 _428_/a_36_151# 0 1.43589f
C20116 FILLER_0_5_72/a_1380_472# 0 0.345058f
C20117 FILLER_0_5_72/a_932_472# 0 0.33241f
C20118 FILLER_0_5_72/a_484_472# 0 0.33241f
C20119 FILLER_0_5_72/a_36_472# 0 0.404746f
C20120 FILLER_0_5_72/a_1468_375# 0 0.233029f
C20121 FILLER_0_5_72/a_1020_375# 0 0.171606f
C20122 FILLER_0_5_72/a_572_375# 0 0.171606f
C20123 FILLER_0_5_72/a_124_375# 0 0.185399f
C20124 _376_/a_36_160# 0 0.386641f
C20125 trim_val\[1\] 0 0.683578f
C20126 _445_/a_2560_156# 0 0.016968f
C20127 _445_/a_2665_112# 0 0.62251f
C20128 _445_/a_2248_156# 0 0.371662f
C20129 _445_/a_1204_472# 0 0.012971f
C20130 _445_/a_1000_472# 0 0.291735f
C20131 _445_/a_796_472# 0 0.023206f
C20132 _445_/a_1308_423# 0 0.279043f
C20133 _445_/a_448_472# 0 0.684413f
C20134 _445_/a_36_151# 0 1.43589f
C20135 fanout67/a_36_160# 0 0.386641f
C20136 fanout56/a_36_113# 0 0.418095f
C20137 net78 0 0.686263f
C20138 fanout78/a_36_113# 0 0.418095f
C20139 _174_ 0 0.979741f
C20140 FILLER_0_0_198/a_36_472# 0 0.417394f
C20141 FILLER_0_0_198/a_124_375# 0 0.246306f
C20142 FILLER_0_15_290/a_36_472# 0 0.417394f
C20143 FILLER_0_15_290/a_124_375# 0 0.246306f
C20144 FILLER_0_24_290/a_36_472# 0 0.417394f
C20145 FILLER_0_24_290/a_124_375# 0 0.246306f
C20146 FILLER_0_4_107/a_1380_472# 0 0.345058f
C20147 FILLER_0_4_107/a_932_472# 0 0.33241f
C20148 FILLER_0_4_107/a_484_472# 0 0.33241f
C20149 FILLER_0_4_107/a_36_472# 0 0.404746f
C20150 FILLER_0_4_107/a_1468_375# 0 0.233029f
C20151 FILLER_0_4_107/a_1020_375# 0 0.171606f
C20152 FILLER_0_4_107/a_572_375# 0 0.171606f
C20153 FILLER_0_4_107/a_124_375# 0 0.185399f
C20154 FILLER_0_7_104/a_1380_472# 0 0.345058f
C20155 FILLER_0_7_104/a_932_472# 0 0.33241f
C20156 FILLER_0_7_104/a_484_472# 0 0.33241f
C20157 FILLER_0_7_104/a_36_472# 0 0.404746f
C20158 FILLER_0_7_104/a_1468_375# 0 0.233029f
C20159 FILLER_0_7_104/a_1020_375# 0 0.171606f
C20160 FILLER_0_7_104/a_572_375# 0 0.171606f
C20161 FILLER_0_7_104/a_124_375# 0 0.185399f
C20162 _214_/a_36_160# 0 0.386641f
C20163 net1 0 0.364811f
C20164 input1/a_36_113# 0 0.418095f
C20165 _429_/a_2560_156# 0 0.016968f
C20166 _429_/a_2665_112# 0 0.62251f
C20167 _429_/a_2248_156# 0 0.371662f
C20168 _429_/a_1204_472# 0 0.012971f
C20169 _429_/a_1000_472# 0 0.291735f
C20170 _429_/a_796_472# 0 0.023206f
C20171 _429_/a_1308_423# 0 0.279043f
C20172 _429_/a_448_472# 0 0.684413f
C20173 _429_/a_36_151# 0 1.43589f
C20174 _011_ 0 0.278979f
C20175 _377_/a_36_472# 0 0.031137f
C20176 fanout66/a_36_113# 0 0.418095f
C20177 _035_ 0 0.327801f
C20178 _446_/a_2560_156# 0 0.016968f
C20179 _446_/a_2665_112# 0 0.62251f
C20180 _446_/a_2248_156# 0 0.371662f
C20181 _446_/a_1204_472# 0 0.012971f
C20182 _446_/a_1000_472# 0 0.291735f
C20183 _446_/a_796_472# 0 0.023206f
C20184 _446_/a_1308_423# 0 0.279043f
C20185 _446_/a_448_472# 0 0.684413f
C20186 _446_/a_36_151# 0 1.43589f
C20187 fanout77/a_36_113# 0 0.418095f
C20188 FILLER_0_5_212/a_36_472# 0 0.417394f
C20189 FILLER_0_5_212/a_124_375# 0 0.246306f
C20190 fanout55/a_36_160# 0 0.696445f
C20191 _175_ 0 0.344159f
C20192 _394_/a_1936_472# 0 0.009918f
C20193 _394_/a_718_524# 0 0.005143f
C20194 _394_/a_56_524# 0 0.41096f
C20195 _394_/a_728_93# 0 0.654825f
C20196 _394_/a_1336_472# 0 0.316639f
C20197 FILLER_0_3_172/a_3172_472# 0 0.345058f
C20198 FILLER_0_3_172/a_2724_472# 0 0.33241f
C20199 FILLER_0_3_172/a_2276_472# 0 0.33241f
C20200 FILLER_0_3_172/a_1828_472# 0 0.33241f
C20201 FILLER_0_3_172/a_1380_472# 0 0.33241f
C20202 FILLER_0_3_172/a_932_472# 0 0.33241f
C20203 FILLER_0_3_172/a_484_472# 0 0.33241f
C20204 FILLER_0_3_172/a_36_472# 0 0.404746f
C20205 FILLER_0_3_172/a_3260_375# 0 0.233093f
C20206 FILLER_0_3_172/a_2812_375# 0 0.17167f
C20207 FILLER_0_3_172/a_2364_375# 0 0.17167f
C20208 FILLER_0_3_172/a_1916_375# 0 0.17167f
C20209 FILLER_0_3_172/a_1468_375# 0 0.17167f
C20210 FILLER_0_3_172/a_1020_375# 0 0.17167f
C20211 FILLER_0_3_172/a_572_375# 0 0.17167f
C20212 FILLER_0_3_172/a_124_375# 0 0.185915f
C20213 FILLER_0_17_72/a_3172_472# 0 0.345058f
C20214 FILLER_0_17_72/a_2724_472# 0 0.33241f
C20215 FILLER_0_17_72/a_2276_472# 0 0.33241f
C20216 FILLER_0_17_72/a_1828_472# 0 0.33241f
C20217 FILLER_0_17_72/a_1380_472# 0 0.33241f
C20218 FILLER_0_17_72/a_932_472# 0 0.33241f
C20219 FILLER_0_17_72/a_484_472# 0 0.33241f
C20220 FILLER_0_17_72/a_36_472# 0 0.404746f
C20221 FILLER_0_17_72/a_3260_375# 0 0.233093f
C20222 FILLER_0_17_72/a_2812_375# 0 0.17167f
C20223 FILLER_0_17_72/a_2364_375# 0 0.17167f
C20224 FILLER_0_17_72/a_1916_375# 0 0.17167f
C20225 FILLER_0_17_72/a_1468_375# 0 0.17167f
C20226 FILLER_0_17_72/a_1020_375# 0 0.17167f
C20227 FILLER_0_17_72/a_572_375# 0 0.17167f
C20228 FILLER_0_17_72/a_124_375# 0 0.185915f
C20229 FILLER_0_2_93/a_484_472# 0 0.345058f
C20230 FILLER_0_2_93/a_36_472# 0 0.404746f
C20231 FILLER_0_2_93/a_572_375# 0 0.232991f
C20232 FILLER_0_2_93/a_124_375# 0 0.185089f
C20233 FILLER_0_11_142/a_484_472# 0 0.345058f
C20234 FILLER_0_11_142/a_36_472# 0 0.404746f
C20235 FILLER_0_11_142/a_572_375# 0 0.232991f
C20236 FILLER_0_11_142/a_124_375# 0 0.185089f
C20237 net25 0 1.803174f
C20238 _232_/a_67_603# 0 0.345683f
C20239 net35 0 1.844415f
C20240 mask\[8\] 0 1.276111f
C20241 _301_/a_36_472# 0 0.031137f
C20242 _033_ 0 0.323682f
C20243 _165_ 0 0.331995f
C20244 FILLER_0_3_2/a_36_472# 0 0.417394f
C20245 FILLER_0_3_2/a_124_375# 0 0.246306f
C20246 trim_val\[3\] 0 0.719615f
C20247 _036_ 0 0.369206f
C20248 net68 0 1.735004f
C20249 _447_/a_2560_156# 0 0.016968f
C20250 _447_/a_2665_112# 0 0.62251f
C20251 _447_/a_2248_156# 0 0.371662f
C20252 _447_/a_1204_472# 0 0.012971f
C20253 _447_/a_1000_472# 0 0.291735f
C20254 _447_/a_796_472# 0 0.023206f
C20255 _447_/a_1308_423# 0 0.279043f
C20256 _447_/a_448_472# 0 0.684413f
C20257 _447_/a_36_151# 0 1.43589f
C20258 FILLER_0_19_28/a_484_472# 0 0.345058f
C20259 FILLER_0_19_28/a_36_472# 0 0.404746f
C20260 FILLER_0_19_28/a_572_375# 0 0.232991f
C20261 FILLER_0_19_28/a_124_375# 0 0.185089f
C20262 fanout65/a_36_113# 0 0.418095f
C20263 fanout76/a_36_160# 0 0.386641f
C20264 net54 0 5.456963f
C20265 fanout54/a_36_160# 0 0.696445f
C20266 FILLER_0_4_49/a_484_472# 0 0.345058f
C20267 FILLER_0_4_49/a_36_472# 0 0.404746f
C20268 FILLER_0_4_49/a_572_375# 0 0.232991f
C20269 FILLER_0_4_49/a_124_375# 0 0.185089f
C20270 _176_ 0 0.804011f
C20271 _085_ 0 2.280803f
C20272 _116_ 0 1.959915f
C20273 _395_/a_36_488# 0 0.101145f
C20274 FILLER_0_14_50/a_36_472# 0 0.417394f
C20275 FILLER_0_14_50/a_124_375# 0 0.246306f
C20276 FILLER_0_8_263/a_36_472# 0 0.417394f
C20277 FILLER_0_8_263/a_124_375# 0 0.246306f
C20278 FILLER_0_0_130/a_36_472# 0 0.417394f
C20279 FILLER_0_0_130/a_124_375# 0 0.246306f
C20280 FILLER_0_16_255/a_36_472# 0 0.417394f
C20281 FILLER_0_16_255/a_124_375# 0 0.246306f
C20282 FILLER_0_7_59/a_484_472# 0 0.345058f
C20283 FILLER_0_7_59/a_36_472# 0 0.404746f
C20284 FILLER_0_7_59/a_572_375# 0 0.232991f
C20285 FILLER_0_7_59/a_124_375# 0 0.185089f
C20286 ctlp[2] 0 0.17528f
C20287 output19/a_224_472# 0 2.38465f
C20288 FILLER_0_7_146/a_36_472# 0 0.417394f
C20289 FILLER_0_7_146/a_124_375# 0 0.246306f
C20290 _216_/a_67_603# 0 0.345683f
C20291 FILLER_0_15_116/a_484_472# 0 0.345058f
C20292 FILLER_0_15_116/a_36_472# 0 0.404746f
C20293 FILLER_0_15_116/a_572_375# 0 0.232991f
C20294 FILLER_0_15_116/a_124_375# 0 0.185089f
C20295 _063_ 0 0.370155f
C20296 _233_/a_36_160# 0 0.386641f
C20297 FILLER_0_21_28/a_3172_472# 0 0.345058f
C20298 FILLER_0_21_28/a_2724_472# 0 0.33241f
C20299 FILLER_0_21_28/a_2276_472# 0 0.33241f
C20300 FILLER_0_21_28/a_1828_472# 0 0.33241f
C20301 FILLER_0_21_28/a_1380_472# 0 0.33241f
C20302 FILLER_0_21_28/a_932_472# 0 0.33241f
C20303 FILLER_0_21_28/a_484_472# 0 0.33241f
C20304 FILLER_0_21_28/a_36_472# 0 0.404746f
C20305 FILLER_0_21_28/a_3260_375# 0 0.233093f
C20306 FILLER_0_21_28/a_2812_375# 0 0.17167f
C20307 FILLER_0_21_28/a_2364_375# 0 0.17167f
C20308 FILLER_0_21_28/a_1916_375# 0 0.17167f
C20309 FILLER_0_21_28/a_1468_375# 0 0.17167f
C20310 FILLER_0_21_28/a_1020_375# 0 0.17167f
C20311 FILLER_0_21_28/a_572_375# 0 0.17167f
C20312 FILLER_0_21_28/a_124_375# 0 0.185915f
C20313 _110_ 0 0.323912f
C20314 _379_/a_36_472# 0 0.031137f
C20315 trim_val\[4\] 0 0.662409f
C20316 net76 0 1.454269f
C20317 _448_/a_2560_156# 0 0.016968f
C20318 _448_/a_2665_112# 0 0.62251f
C20319 _448_/a_2248_156# 0 0.371662f
C20320 _448_/a_1204_472# 0 0.012971f
C20321 _448_/a_1000_472# 0 0.291735f
C20322 _448_/a_796_472# 0 0.023206f
C20323 _448_/a_1308_423# 0 0.279043f
C20324 _448_/a_448_472# 0 0.684413f
C20325 _448_/a_36_151# 0 1.43589f
C20326 fanout64/a_36_160# 0 0.386641f
C20327 fanout75/a_36_113# 0 0.418095f
C20328 _250_/a_36_68# 0 0.69549f
C20329 net56 0 0.843396f
C20330 fanout53/a_36_160# 0 0.696445f
C20331 _177_ 0 0.358286f
C20332 result[2] 0 0.230851f
C20333 net29 0 1.802718f
C20334 output29/a_224_472# 0 2.38465f
C20335 ctlp[1] 0 0.17418f
C20336 output18/a_224_472# 0 2.38465f
C20337 FILLER_0_14_181/a_36_472# 0 0.417394f
C20338 FILLER_0_14_181/a_124_375# 0 0.246306f
C20339 _052_ 0 0.569133f
C20340 _217_/a_36_160# 0 0.386641f
C20341 net44 0 1.407054f
C20342 _303_/a_36_472# 0 0.031137f
C20343 en_co_clk 0 0.346872f
C20344 net55 0 5.119958f
C20345 net72 0 1.366255f
C20346 _449_/a_2560_156# 0 0.016968f
C20347 _449_/a_2665_112# 0 0.62251f
C20348 _449_/a_2248_156# 0 0.371662f
C20349 _449_/a_1204_472# 0 0.012971f
C20350 _449_/a_1000_472# 0 0.291735f
C20351 _449_/a_796_472# 0 0.023206f
C20352 _449_/a_1308_423# 0 0.279043f
C20353 _449_/a_448_472# 0 0.684413f
C20354 _449_/a_36_151# 0 1.43589f
C20355 fanout52/a_36_160# 0 0.696445f
C20356 net82 0 0.706042f
C20357 fanout74/a_36_113# 0 0.418095f
C20358 FILLER_0_10_28/a_36_472# 0 0.417394f
C20359 FILLER_0_10_28/a_124_375# 0 0.246306f
C20360 mask\[0\] 0 2.242948f
C20361 _320_/a_36_472# 0 0.137725f
C20362 fanout63/a_36_160# 0 0.696445f
C20363 FILLER_0_14_81/a_36_472# 0 0.417394f
C20364 FILLER_0_14_81/a_124_375# 0 0.246306f
C20365 _397_/a_36_472# 0 0.031137f
C20366 FILLER_0_13_212/a_1380_472# 0 0.345058f
C20367 FILLER_0_13_212/a_932_472# 0 0.33241f
C20368 FILLER_0_13_212/a_484_472# 0 0.33241f
C20369 FILLER_0_13_212/a_36_472# 0 0.404746f
C20370 FILLER_0_13_212/a_1468_375# 0 0.233029f
C20371 FILLER_0_13_212/a_1020_375# 0 0.171606f
C20372 FILLER_0_13_212/a_572_375# 0 0.171606f
C20373 FILLER_0_13_212/a_124_375# 0 0.185399f
C20374 trim[1] 0 0.793787f
C20375 net39 0 1.445128f
C20376 output39/a_224_472# 0 2.38465f
C20377 result[1] 0 0.229507f
C20378 net28 0 1.759728f
C20379 output28/a_224_472# 0 2.38465f
C20380 ctlp[0] 0 1.002286f
C20381 output17/a_224_472# 0 2.38465f
C20382 FILLER_0_16_37/a_36_472# 0 0.417394f
C20383 FILLER_0_16_37/a_124_375# 0 0.246306f
C20384 net26 0 1.671545f
C20385 _064_ 0 0.581481f
C20386 trim_val\[2\] 0 0.65354f
C20387 trim_mask\[2\] 0 0.92551f
C20388 _235_/a_67_603# 0 0.345683f
C20389 _013_ 0 0.48783f
C20390 _111_ 0 0.369652f
C20391 FILLER_0_18_177/a_3172_472# 0 0.345058f
C20392 FILLER_0_18_177/a_2724_472# 0 0.33241f
C20393 FILLER_0_18_177/a_2276_472# 0 0.33241f
C20394 FILLER_0_18_177/a_1828_472# 0 0.33241f
C20395 FILLER_0_18_177/a_1380_472# 0 0.33241f
C20396 FILLER_0_18_177/a_932_472# 0 0.33241f
C20397 FILLER_0_18_177/a_484_472# 0 0.33241f
C20398 FILLER_0_18_177/a_36_472# 0 0.404746f
C20399 FILLER_0_18_177/a_3260_375# 0 0.233093f
C20400 FILLER_0_18_177/a_2812_375# 0 0.17167f
C20401 FILLER_0_18_177/a_2364_375# 0 0.17167f
C20402 FILLER_0_18_177/a_1916_375# 0 0.17167f
C20403 FILLER_0_18_177/a_1468_375# 0 0.17167f
C20404 FILLER_0_18_177/a_1020_375# 0 0.17167f
C20405 FILLER_0_18_177/a_572_375# 0 0.17167f
C20406 FILLER_0_18_177/a_124_375# 0 0.185915f
C20407 FILLER_0_18_100/a_36_472# 0 0.417394f
C20408 FILLER_0_18_100/a_124_375# 0 0.246306f
C20409 _073_ 0 0.953711f
C20410 _126_ 0 2.036767f
C20411 _069_ 0 2.034557f
C20412 _321_/a_170_472# 0 0.077257f
C20413 fanout51/a_36_113# 0 0.418095f
C20414 fanout62/a_36_160# 0 0.696445f
C20415 fanout73/a_36_113# 0 0.418095f
C20416 FILLER_0_19_47/a_484_472# 0 0.345058f
C20417 FILLER_0_19_47/a_36_472# 0 0.404746f
C20418 FILLER_0_19_47/a_572_375# 0 0.232991f
C20419 FILLER_0_19_47/a_124_375# 0 0.185089f
C20420 FILLER_0_14_91/a_484_472# 0 0.345058f
C20421 FILLER_0_14_91/a_36_472# 0 0.404746f
C20422 FILLER_0_14_91/a_572_375# 0 0.232991f
C20423 FILLER_0_14_91/a_124_375# 0 0.185089f
C20424 FILLER_0_10_214/a_36_472# 0 0.417394f
C20425 FILLER_0_10_214/a_124_375# 0 0.246306f
C20426 FILLER_0_10_247/a_36_472# 0 0.417394f
C20427 FILLER_0_10_247/a_124_375# 0 0.246306f
C20428 _178_ 0 1.252435f
C20429 _398_/a_36_113# 0 0.418095f
C20430 FILLER_0_16_241/a_36_472# 0 0.417394f
C20431 FILLER_0_16_241/a_124_375# 0 0.246306f
C20432 trim[0] 0 0.796081f
C20433 net38 0 1.529392f
C20434 output38/a_224_472# 0 2.38465f
C20435 ctln[9] 0 0.904836f
C20436 net16 0 1.295744f
C20437 output16/a_224_472# 0 2.38465f
C20438 result[0] 0 0.56622f
C20439 net27 0 2.023744f
C20440 output27/a_224_472# 0 2.38465f
C20441 _219_/a_36_160# 0 0.386641f
C20442 FILLER_0_20_193/a_484_472# 0 0.345058f
C20443 FILLER_0_20_193/a_36_472# 0 0.404746f
C20444 FILLER_0_20_193/a_572_375# 0 0.232991f
C20445 FILLER_0_20_193/a_124_375# 0 0.185089f
C20446 _236_/a_36_160# 0 0.696445f
C20447 _112_ 0 0.308886f
C20448 _305_/a_36_159# 0 0.374116f
C20449 _074_ 0 1.813232f
C20450 _253_/a_36_68# 0 0.061249f
C20451 net50 0 4.486121f
C20452 net52 0 3.536016f
C20453 fanout50/a_36_160# 0 0.696445f
C20454 FILLER_0_10_37/a_36_472# 0 0.417394f
C20455 FILLER_0_10_37/a_124_375# 0 0.246306f
C20456 fanout72/a_36_113# 0 0.418095f
C20457 fanout61/a_36_113# 0 0.418095f
C20458 _128_ 0 0.447252f
C20459 _127_ 0 1.291729f
C20460 _322_/a_848_380# 0 0.40208f
C20461 _322_/a_124_24# 0 0.591898f
C20462 _088_ 0 0.457961f
C20463 _079_ 0 1.114894f
C20464 _087_ 0 0.601674f
C20465 _270_/a_36_472# 0 0.031137f
C20466 FILLER_0_4_123/a_36_472# 0 0.417394f
C20467 FILLER_0_4_123/a_124_375# 0 0.246306f
C20468 FILLER_0_17_218/a_484_472# 0 0.345058f
C20469 FILLER_0_17_218/a_36_472# 0 0.404746f
C20470 FILLER_0_17_218/a_572_375# 0 0.232991f
C20471 FILLER_0_17_218/a_124_375# 0 0.185089f
C20472 valid 0 0.272072f
C20473 net48 0 1.219262f
C20474 output48/a_224_472# 0 2.38465f
C20475 sample 0 0.508149f
C20476 output37/a_224_472# 0 2.38465f
C20477 ctln[8] 0 1.547984f
C20478 output15/a_224_472# 0 2.38465f
C20479 ctlp[9] 0 0.73349f
C20480 output26/a_224_472# 0 2.38465f
C20481 FILLER_0_16_57/a_1380_472# 0 0.345058f
C20482 FILLER_0_16_57/a_932_472# 0 0.33241f
C20483 FILLER_0_16_57/a_484_472# 0 0.33241f
C20484 FILLER_0_16_57/a_36_472# 0 0.404746f
C20485 FILLER_0_16_57/a_1468_375# 0 0.233029f
C20486 FILLER_0_16_57/a_1020_375# 0 0.171606f
C20487 FILLER_0_16_57/a_572_375# 0 0.171606f
C20488 FILLER_0_16_57/a_124_375# 0 0.185399f
C20489 _306_/a_36_68# 0 0.69549f
C20490 _072_ 0 2.604301f
C20491 fanout82/a_36_113# 0 0.418095f
C20492 _015_ 0 0.406653f
C20493 _323_/a_36_113# 0 0.418095f
C20494 net60 0 5.024503f
C20495 net61 0 1.666523f
C20496 fanout60/a_36_160# 0 0.696445f
C20497 fanout71/a_36_113# 0 0.418095f
C20498 FILLER_0_6_239/a_36_472# 0 0.417394f
C20499 FILLER_0_6_239/a_124_375# 0 0.246306f
C20500 FILLER_0_4_99/a_36_472# 0 0.417394f
C20501 FILLER_0_4_99/a_124_375# 0 0.246306f
C20502 net57 0 1.383718f
C20503 FILLER_0_10_256/a_36_472# 0 0.417394f
C20504 FILLER_0_10_256/a_124_375# 0 0.246306f
C20505 cal_itt\[3\] 0 1.854962f
C20506 _340_/a_36_160# 0 0.386641f
C20507 FILLER_0_4_177/a_484_472# 0 0.345058f
C20508 FILLER_0_4_177/a_36_472# 0 0.404746f
C20509 FILLER_0_4_177/a_572_375# 0 0.232991f
C20510 FILLER_0_4_177/a_124_375# 0 0.185089f
C20511 FILLER_0_4_144/a_484_472# 0 0.345058f
C20512 FILLER_0_4_144/a_36_472# 0 0.404746f
C20513 FILLER_0_4_144/a_572_375# 0 0.232991f
C20514 FILLER_0_4_144/a_124_375# 0 0.185089f
C20515 ctln[7] 0 1.265946f
C20516 output14/a_224_472# 0 2.38465f
C20517 result[9] 0 0.8197f
C20518 output36/a_224_472# 0 2.38465f
C20519 trimb[4] 0 0.752332f
C20520 output47/a_224_472# 0 2.38465f
C20521 ctlp[8] 0 1.136333f
C20522 output25/a_224_472# 0 2.38465f
C20523 FILLER_0_12_136/a_1380_472# 0 0.345058f
C20524 FILLER_0_12_136/a_932_472# 0 0.33241f
C20525 FILLER_0_12_136/a_484_472# 0 0.33241f
C20526 FILLER_0_12_136/a_36_472# 0 0.404746f
C20527 FILLER_0_12_136/a_1468_375# 0 0.233029f
C20528 FILLER_0_12_136/a_1020_375# 0 0.171606f
C20529 FILLER_0_12_136/a_572_375# 0 0.171606f
C20530 FILLER_0_12_136/a_124_375# 0 0.185399f
C20531 FILLER_0_16_89/a_1380_472# 0 0.345058f
C20532 FILLER_0_16_89/a_932_472# 0 0.33241f
C20533 FILLER_0_16_89/a_484_472# 0 0.33241f
C20534 FILLER_0_16_89/a_36_472# 0 0.404746f
C20535 FILLER_0_16_89/a_1468_375# 0 0.233029f
C20536 FILLER_0_16_89/a_1020_375# 0 0.171606f
C20537 FILLER_0_16_89/a_572_375# 0 0.171606f
C20538 FILLER_0_16_89/a_124_375# 0 0.185399f
C20539 FILLER_0_21_125/a_484_472# 0 0.345058f
C20540 FILLER_0_21_125/a_36_472# 0 0.404746f
C20541 FILLER_0_21_125/a_572_375# 0 0.232991f
C20542 FILLER_0_21_125/a_124_375# 0 0.185089f
C20543 _238_/a_67_603# 0 0.345683f
C20544 _096_ 0 2.205532f
C20545 _093_ 0 1.893313f
C20546 FILLER_0_19_55/a_36_472# 0 0.417394f
C20547 FILLER_0_19_55/a_124_375# 0 0.246306f
C20548 net81 0 1.738987f
C20549 fanout81/a_36_160# 0 0.386641f
C20550 _057_ 0 1.600886f
C20551 _255_/a_224_552# 0 1.31114f
C20552 net73 0 1.058857f
C20553 fanout70/a_36_113# 0 0.418095f
C20554 _003_ 0 0.3064f
C20555 _089_ 0 0.36777f
C20556 _272_/a_36_472# 0 0.031137f
C20557 _187_ 0 0.311229f
C20558 _410_/a_36_68# 0 0.112263f
C20559 _141_ 0 1.249289f
C20560 mask\[3\] 0 1.26722f
C20561 _341_/a_49_472# 0 0.054843f
C20562 cal 0 0.793393f
C20563 FILLER_0_7_195/a_36_472# 0 0.417394f
C20564 FILLER_0_7_195/a_124_375# 0 0.246306f
C20565 FILLER_0_7_162/a_36_472# 0 0.417394f
C20566 FILLER_0_7_162/a_124_375# 0 0.246306f
C20567 ctln[6] 0 1.451644f
C20568 output13/a_224_472# 0 2.38465f
C20569 FILLER_0_18_2/a_3172_472# 0 0.345058f
C20570 FILLER_0_18_2/a_2724_472# 0 0.33241f
C20571 FILLER_0_18_2/a_2276_472# 0 0.33241f
C20572 FILLER_0_18_2/a_1828_472# 0 0.33241f
C20573 FILLER_0_18_2/a_1380_472# 0 0.33241f
C20574 FILLER_0_18_2/a_932_472# 0 0.33241f
C20575 FILLER_0_18_2/a_484_472# 0 0.33241f
C20576 FILLER_0_18_2/a_36_472# 0 0.404746f
C20577 FILLER_0_18_2/a_3260_375# 0 0.233093f
C20578 FILLER_0_18_2/a_2812_375# 0 0.17167f
C20579 FILLER_0_18_2/a_2364_375# 0 0.17167f
C20580 FILLER_0_18_2/a_1916_375# 0 0.17167f
C20581 FILLER_0_18_2/a_1468_375# 0 0.17167f
C20582 FILLER_0_18_2/a_1020_375# 0 0.17167f
C20583 FILLER_0_18_2/a_572_375# 0 0.17167f
C20584 FILLER_0_18_2/a_124_375# 0 0.185915f
C20585 trimb[3] 0 0.34698f
C20586 net46 0 1.13395f
C20587 output46/a_224_472# 0 2.38465f
C20588 result[8] 0 0.68837f
C20589 output35/a_224_472# 0 2.38465f
C20590 ctlp[7] 0 0.83567f
C20591 output24/a_224_472# 0 2.38465f
C20592 FILLER_0_8_107/a_36_472# 0 0.417394f
C20593 FILLER_0_8_107/a_124_375# 0 0.246306f
C20594 FILLER_0_12_124/a_36_472# 0 0.417394f
C20595 FILLER_0_12_124/a_124_375# 0 0.246306f
C20596 net41 0 1.746759f
C20597 _065_ 0 0.523724f
C20598 _239_/a_36_160# 0 0.696445f
C20599 FILLER_0_1_98/a_36_472# 0 0.417394f
C20600 FILLER_0_1_98/a_124_375# 0 0.246306f
C20601 _115_ 0 1.281516f
C20602 _114_ 0 2.293579f
C20603 _308_/a_848_380# 0 0.40208f
C20604 _308_/a_124_24# 0 0.591898f
C20605 _256_/a_36_68# 0 0.063181f
C20606 FILLER_0_10_78/a_1380_472# 0 0.345058f
C20607 FILLER_0_10_78/a_932_472# 0 0.33241f
C20608 FILLER_0_10_78/a_484_472# 0 0.33241f
C20609 FILLER_0_10_78/a_36_472# 0 0.404746f
C20610 FILLER_0_10_78/a_1468_375# 0 0.233029f
C20611 FILLER_0_10_78/a_1020_375# 0 0.171606f
C20612 FILLER_0_10_78/a_572_375# 0 0.171606f
C20613 FILLER_0_10_78/a_124_375# 0 0.185399f
C20614 _130_ 0 0.304085f
C20615 net80 0 1.375599f
C20616 fanout80/a_36_113# 0 0.418095f
C20617 net58 0 5.308423f
C20618 _000_ 0 0.382358f
C20619 net75 0 1.474299f
C20620 _411_/a_2560_156# 0 0.016968f
C20621 _411_/a_2665_112# 0 0.62251f
C20622 _411_/a_2248_156# 0 0.371662f
C20623 _411_/a_1204_472# 0 0.012971f
C20624 _411_/a_1000_472# 0 0.291735f
C20625 _411_/a_796_472# 0 0.023206f
C20626 _411_/a_1308_423# 0 0.279043f
C20627 _411_/a_448_472# 0 0.684413f
C20628 _411_/a_36_151# 0 1.43589f
C20629 state\[0\] 0 0.680109f
C20630 _273_/a_36_68# 0 0.69549f
C20631 _142_ 0 0.324372f
C20632 FILLER_0_9_223/a_484_472# 0 0.345058f
C20633 FILLER_0_9_223/a_36_472# 0 0.404746f
C20634 FILLER_0_9_223/a_572_375# 0 0.232991f
C20635 FILLER_0_9_223/a_124_375# 0 0.185089f
C20636 FILLER_0_4_197/a_1380_472# 0 0.345058f
C20637 FILLER_0_4_197/a_932_472# 0 0.33241f
C20638 FILLER_0_4_197/a_484_472# 0 0.33241f
C20639 FILLER_0_4_197/a_36_472# 0 0.404746f
C20640 FILLER_0_4_197/a_1468_375# 0 0.233029f
C20641 FILLER_0_4_197/a_1020_375# 0 0.171606f
C20642 FILLER_0_4_197/a_572_375# 0 0.171606f
C20643 FILLER_0_4_197/a_124_375# 0 0.185399f
C20644 FILLER_0_17_226/a_36_472# 0 0.417394f
C20645 FILLER_0_17_226/a_124_375# 0 0.246306f
C20646 FILLER_0_5_109/a_484_472# 0 0.345058f
C20647 FILLER_0_5_109/a_36_472# 0 0.404746f
C20648 FILLER_0_5_109/a_572_375# 0 0.232991f
C20649 FILLER_0_5_109/a_124_375# 0 0.185089f
C20650 ctln[5] 0 1.585113f
C20651 output12/a_224_472# 0 2.38465f
C20652 result[7] 0 0.24756f
C20653 net34 0 1.724665f
C20654 output34/a_224_472# 0 2.38465f
C20655 trimb[2] 0 0.839614f
C20656 net45 0 1.12041f
C20657 output45/a_224_472# 0 2.38465f
C20658 ctlp[6] 0 1.243017f
C20659 output23/a_224_472# 0 2.38465f
C20660 FILLER_0_15_142/a_484_472# 0 0.345058f
C20661 FILLER_0_15_142/a_36_472# 0 0.404746f
C20662 FILLER_0_15_142/a_572_375# 0 0.232991f
C20663 FILLER_0_15_142/a_124_375# 0 0.185089f
C20664 _077_ 0 1.645892f
C20665 _075_ 0 0.374516f
C20666 _257_/a_36_472# 0 0.031137f
C20667 _326_/a_36_160# 0 0.696445f
C20668 _412_/a_2560_156# 0 0.016968f
C20669 _412_/a_2665_112# 0 0.62251f
C20670 _412_/a_2248_156# 0 0.371662f
C20671 _412_/a_1204_472# 0 0.012971f
C20672 _412_/a_1000_472# 0 0.291735f
C20673 _412_/a_796_472# 0 0.023206f
C20674 _412_/a_1308_423# 0 0.279043f
C20675 _412_/a_448_472# 0 0.684413f
C20676 _412_/a_36_151# 0 1.43589f
C20677 _091_ 0 1.841339f
C20678 _274_/a_36_68# 0 0.063181f
C20679 _143_ 0 0.329289f
C20680 mask\[4\] 0 1.300438f
C20681 _343_/a_49_472# 0 0.054843f
C20682 FILLER_0_13_65/a_36_472# 0 0.417394f
C20683 FILLER_0_13_65/a_124_375# 0 0.246306f
C20684 _360_/a_36_160# 0 0.386641f
C20685 FILLER_0_4_185/a_36_472# 0 0.417394f
C20686 FILLER_0_4_185/a_124_375# 0 0.246306f
C20687 FILLER_0_4_152/a_36_472# 0 0.417394f
C20688 FILLER_0_4_152/a_124_375# 0 0.246306f
C20689 _291_/a_36_160# 0 0.386641f
C20690 ctln[2] 0 1.833091f
C20691 output9/a_224_472# 0 2.38465f
C20692 ctln[4] 0 1.461847f
C20693 output11/a_224_472# 0 2.38465f
C20694 trimb[1] 0 0.378532f
C20695 output44/a_224_472# 0 2.38465f
C20696 result[6] 0 0.19512f
C20697 output33/a_224_472# 0 2.38465f
C20698 ctlp[5] 0 1.282822f
C20699 output22/a_224_472# 0 2.38465f
C20700 FILLER_0_8_127/a_36_472# 0 0.417394f
C20701 FILLER_0_8_127/a_124_375# 0 0.246306f
C20702 FILLER_0_8_138/a_36_472# 0 0.417394f
C20703 FILLER_0_8_138/a_124_375# 0 0.246306f
C20704 FILLER_0_21_133/a_36_472# 0 0.417394f
C20705 FILLER_0_21_133/a_124_375# 0 0.246306f
C20706 FILLER_0_24_130/a_36_472# 0 0.417394f
C20707 FILLER_0_24_130/a_124_375# 0 0.246306f
C20708 FILLER_0_18_171/a_36_472# 0 0.417394f
C20709 FILLER_0_18_171/a_124_375# 0 0.246306f
C20710 _258_/a_36_160# 0 0.386641f
C20711 _016_ 0 0.314121f
C20712 _327_/a_36_472# 0 0.031137f
C20713 _189_/a_67_603# 0 0.345683f
C20714 FILLER_0_24_63/a_36_472# 0 0.417394f
C20715 FILLER_0_24_63/a_124_375# 0 0.246306f
C20716 FILLER_0_24_96/a_36_472# 0 0.417394f
C20717 FILLER_0_24_96/a_124_375# 0 0.246306f
C20718 cal_itt\[2\] 0 1.473514f
C20719 _002_ 0 0.289553f
C20720 _413_/a_2560_156# 0 0.016968f
C20721 _413_/a_2665_112# 0 0.62251f
C20722 _413_/a_2248_156# 0 0.371662f
C20723 _413_/a_1204_472# 0 0.012971f
C20724 _413_/a_1000_472# 0 0.291735f
C20725 _413_/a_796_472# 0 0.023206f
C20726 _413_/a_1308_423# 0 0.279043f
C20727 _413_/a_448_472# 0 0.684413f
C20728 _413_/a_36_151# 0 1.43589f
C20729 _092_ 0 0.680239f
C20730 FILLER_0_7_72/a_3172_472# 0 0.345058f
C20731 FILLER_0_7_72/a_2724_472# 0 0.33241f
C20732 FILLER_0_7_72/a_2276_472# 0 0.33241f
C20733 FILLER_0_7_72/a_1828_472# 0 0.33241f
C20734 FILLER_0_7_72/a_1380_472# 0 0.33241f
C20735 FILLER_0_7_72/a_932_472# 0 0.33241f
C20736 FILLER_0_7_72/a_484_472# 0 0.33241f
C20737 FILLER_0_7_72/a_36_472# 0 0.404746f
C20738 FILLER_0_7_72/a_3260_375# 0 0.233093f
C20739 FILLER_0_7_72/a_2812_375# 0 0.17167f
C20740 FILLER_0_7_72/a_2364_375# 0 0.17167f
C20741 FILLER_0_7_72/a_1916_375# 0 0.17167f
C20742 FILLER_0_7_72/a_1468_375# 0 0.17167f
C20743 FILLER_0_7_72/a_1020_375# 0 0.17167f
C20744 FILLER_0_7_72/a_572_375# 0 0.17167f
C20745 FILLER_0_7_72/a_124_375# 0 0.185915f
C20746 _086_ 0 2.45259f
C20747 _119_ 0 1.237181f
C20748 net63 0 5.362473f
C20749 _430_/a_2560_156# 0 0.016968f
C20750 _430_/a_2665_112# 0 0.62251f
C20751 _430_/a_2248_156# 0 0.371662f
C20752 _430_/a_1204_472# 0 0.012971f
C20753 _430_/a_1000_472# 0 0.291735f
C20754 _430_/a_796_472# 0 0.023206f
C20755 _430_/a_1308_423# 0 0.279043f
C20756 _430_/a_448_472# 0 0.684413f
C20757 _430_/a_36_151# 0 1.43589f
C20758 _292_/a_36_160# 0 0.386641f
C20759 comp 0 1.022965f
C20760 ctln[1] 0 1.11973f
C20761 output8/a_224_472# 0 2.38465f
C20762 ctln[3] 0 0.835391f
C20763 output10/a_224_472# 0 2.38465f
C20764 result[5] 0 0.206867f
C20765 net32 0 1.78884f
C20766 output32/a_224_472# 0 2.38465f
C20767 trimb[0] 0 0.847787f
C20768 output43/a_224_472# 0 2.38465f
C20769 ctlp[4] 0 0.37565f
C20770 output21/a_224_472# 0 2.38465f
C20771 _053_ 0 1.705161f
C20772 FILLER_0_16_107/a_484_472# 0 0.345058f
C20773 FILLER_0_16_107/a_36_472# 0 0.404746f
C20774 FILLER_0_16_107/a_572_375# 0 0.232991f
C20775 FILLER_0_16_107/a_124_375# 0 0.185089f
C20776 FILLER_0_3_204/a_36_472# 0 0.417394f
C20777 FILLER_0_3_204/a_124_375# 0 0.246306f
C20778 FILLER_0_9_28/a_3172_472# 0 0.345058f
C20779 FILLER_0_9_28/a_2724_472# 0 0.33241f
C20780 FILLER_0_9_28/a_2276_472# 0 0.33241f
C20781 FILLER_0_9_28/a_1828_472# 0 0.33241f
C20782 FILLER_0_9_28/a_1380_472# 0 0.33241f
C20783 FILLER_0_9_28/a_932_472# 0 0.33241f
C20784 FILLER_0_9_28/a_484_472# 0 0.33241f
C20785 FILLER_0_9_28/a_36_472# 0 0.404746f
C20786 FILLER_0_9_28/a_3260_375# 0 0.233093f
C20787 FILLER_0_9_28/a_2812_375# 0 0.17167f
C20788 FILLER_0_9_28/a_2364_375# 0 0.17167f
C20789 FILLER_0_9_28/a_1916_375# 0 0.17167f
C20790 FILLER_0_9_28/a_1468_375# 0 0.17167f
C20791 FILLER_0_9_28/a_1020_375# 0 0.17167f
C20792 FILLER_0_9_28/a_572_375# 0 0.17167f
C20793 FILLER_0_9_28/a_124_375# 0 0.185915f
C20794 _132_ 0 1.491425f
C20795 _328_/a_36_113# 0 0.418095f
C20796 _414_/a_2560_156# 0 0.016968f
C20797 _414_/a_2665_112# 0 0.62251f
C20798 _414_/a_2248_156# 0 0.371662f
C20799 _414_/a_1204_472# 0 0.012971f
C20800 _414_/a_1000_472# 0 0.291735f
C20801 _414_/a_796_472# 0 0.023206f
C20802 _414_/a_1308_423# 0 0.279043f
C20803 _414_/a_448_472# 0 0.684413f
C20804 _414_/a_36_151# 0 1.43589f
C20805 _276_/a_36_160# 0 0.386641f
C20806 _144_ 0 1.173846f
C20807 _345_/a_36_160# 0 0.386641f
C20808 _155_ 0 0.638535f
C20809 _020_ 0 0.316793f
C20810 _431_/a_2560_156# 0 0.016968f
C20811 _431_/a_2665_112# 0 0.62251f
C20812 _431_/a_2248_156# 0 0.371662f
C20813 _431_/a_1204_472# 0 0.012971f
C20814 _431_/a_1000_472# 0 0.291735f
C20815 _431_/a_796_472# 0 0.023206f
C20816 _431_/a_1308_423# 0 0.279043f
C20817 _431_/a_448_472# 0 0.684413f
C20818 _431_/a_36_151# 0 1.43589f
C20819 _105_ 0 1.21281f
C20820 _293_/a_36_472# 0 0.031137f
C20821 FILLER_0_5_128/a_484_472# 0 0.345058f
C20822 FILLER_0_5_128/a_36_472# 0 0.404746f
C20823 FILLER_0_5_128/a_572_375# 0 0.232991f
C20824 FILLER_0_5_128/a_124_375# 0 0.185089f
C20825 FILLER_0_5_117/a_36_472# 0 0.417394f
C20826 FILLER_0_5_117/a_124_375# 0 0.246306f
C20827 ctln[0] 0 1.423102f
C20828 net7 0 1.174913f
C20829 output7/a_224_472# 0 2.38465f
C20830 trim[4] 0 0.763069f
C20831 output42/a_224_472# 0 2.38465f
C20832 result[4] 0 0.038878f
C20833 net31 0 1.912935f
C20834 output31/a_224_472# 0 2.38465f
C20835 ctlp[3] 0 1.14968f
C20836 output20/a_224_472# 0 2.38465f
C20837 FILLER_0_16_73/a_484_472# 0 0.345058f
C20838 FILLER_0_16_73/a_36_472# 0 0.404746f
C20839 FILLER_0_16_73/a_572_375# 0 0.232991f
C20840 FILLER_0_16_73/a_124_375# 0 0.185089f
C20841 FILLER_0_21_142/a_484_472# 0 0.345058f
C20842 FILLER_0_21_142/a_36_472# 0 0.404746f
C20843 FILLER_0_21_142/a_572_375# 0 0.232991f
C20844 FILLER_0_21_142/a_124_375# 0 0.185089f
C20845 FILLER_0_15_150/a_36_472# 0 0.417394f
C20846 FILLER_0_15_150/a_124_375# 0 0.246306f
C20847 FILLER_0_19_125/a_36_472# 0 0.417394f
C20848 FILLER_0_19_125/a_124_375# 0 0.246306f
C20849 net10 0 1.480101f
C20850 net20 0 2.034189f
C20851 _277_/a_36_160# 0 0.386641f
C20852 _004_ 0 0.390107f
C20853 _415_/a_2560_156# 0 0.016968f
C20854 _415_/a_2665_112# 0 0.62251f
C20855 _415_/a_2248_156# 0 0.371662f
C20856 _415_/a_1204_472# 0 0.012971f
C20857 _415_/a_1000_472# 0 0.291735f
C20858 _415_/a_796_472# 0 0.023206f
C20859 _415_/a_1308_423# 0 0.279043f
C20860 _415_/a_448_472# 0 0.684413f
C20861 _415_/a_36_151# 0 1.43589f
C20862 mask\[5\] 0 1.334568f
C20863 _346_/a_49_472# 0 0.054843f
C20864 _028_ 0 0.386029f
C20865 _363_/a_36_68# 0 0.150048f
C20866 _021_ 0 0.316776f
C20867 _432_/a_2560_156# 0 0.016968f
C20868 _432_/a_2665_112# 0 0.62251f
C20869 _432_/a_2248_156# 0 0.371662f
C20870 _432_/a_1204_472# 0 0.012971f
C20871 _432_/a_1000_472# 0 0.291735f
C20872 _432_/a_796_472# 0 0.023206f
C20873 _432_/a_1308_423# 0 0.279043f
C20874 _432_/a_448_472# 0 0.684413f
C20875 _432_/a_36_151# 0 1.43589f
C20876 _008_ 0 0.423631f
C20877 _104_ 0 1.435764f
C20878 _106_ 0 0.378703f
C20879 FILLER_0_17_200/a_484_472# 0 0.345058f
C20880 FILLER_0_17_200/a_36_472# 0 0.404746f
C20881 FILLER_0_17_200/a_572_375# 0 0.232991f
C20882 FILLER_0_17_200/a_124_375# 0 0.185089f
.ends

