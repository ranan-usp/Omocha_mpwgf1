* NGSPICE file created from sarlogic.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VPW VNW VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VPW VNW VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VPW VNW VSUBS
X0 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN B1 a_257_69# VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VPW VNW VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VPW VNW VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VPW VNW VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VSUBS nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VPW VNW VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_455_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VPW VNW VSUBS
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VSUBS nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VSUBS nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VPW VNW VSUBS
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VSUBS nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VPW VNW VSUBS
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VSUBS nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VSUBS nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VPW VNW VSUBS
X0 VSS B a_36_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VPW VNW VSUBS
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VSUBS nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VSUBS nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VPW VNW VSUBS
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VSUBS nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VSUBS nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VSUBS nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VSUBS nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VSS B ZN VSUBS nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VSUBS nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VPW VNW VSUBS
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VPW VNW VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_1458_68# A3 a_1254_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VPW VNW VSUBS
X0 a_1229_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VSUBS nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VSUBS nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VSUBS nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VSUBS nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VSUBS nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VSS A2 a_1133_69# VSUBS nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VSUBS nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VSUBS nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VPW VNW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VPW VNW VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VSUBS nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VSUBS nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VSUBS nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VSUBS nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VSUBS nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VSUBS nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctln[8] ctln[9] 
+ ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8] ctlp[9] 
+ result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7] result[8] result[9] 
+ trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] 
+ rstn en cal clk comp clkc sample valid vdd vss 
XFILLER_0_17_200 vdd vss FILLER_0_17_200/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd ANTENNA_fanout56_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_432_ _021_ mask\[3\] net63 vss net80 vdd _432_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_294_ vdd vss _008_ _104_ _106_ _294_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ _363_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ _346_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd _415_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd _277_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 _200_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd _329_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss FILLER_0_19_125/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd ANTENNA__392__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss FILLER_0_15_150/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss FILLER_0_21_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss FILLER_0_16_73/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss output20/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss output31/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss output42/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss FILLER_0_5_117/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss FILLER_0_5_128/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput7 ctln[0] net7 vdd vss output7/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_431_ _020_ mask\[2\] net53 vss net70 vdd _431_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_293_ net31 vdd vss _106_ mask\[4\] _105_ _293_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_362_ vdd vss trim_mask\[1\] _155_ _362_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_276_ vss _093_ _092_ vdd _276_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_345_ vss _144_ _132_ vdd _345_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd _414_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd _328_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss FILLER_0_9_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_259_ _078_ vdd vss _080_ _073_ _076_ _259_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_204 vdd vss FILLER_0_3_204/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_107 vdd vss FILLER_0_16_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd ANTENNA_fanout79_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd ANTENNA__358__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss output21/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss output32/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss output43/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss output10/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss output8/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd ANTENNA_input3_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_430_ _019_ mask\[1\] net63 vss net80 vdd _430_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_292_ vss _105_ _098_ vdd _292_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_361_ vdd vss _154_ _086_ _119_ _361_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss FILLER_0_7_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ _344_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ _275_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd _413_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__191__I vss net17 vdd ANTENNA__191__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_96 vdd vss FILLER_0_24_96/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss FILLER_0_24_63/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_327_ _131_ vdd vss _016_ _127_ _130_ _327_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_189_ vdd vss _043_ net27 mask\[0\] _189_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_258_ vss _079_ _078_ vdd _258_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss FILLER_0_18_171/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss FILLER_0_24_130/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd ANTENNA__377__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss FILLER_0_21_133/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss FILLER_0_8_127/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss FILLER_0_8_138/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput33 result[6] net33 vdd vss output33/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput22 ctlp[5] net22 vdd vss output22/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss output44/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss output9/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss output11/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd ANTENNA__194__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd _291_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss FILLER_0_4_152/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss FILLER_0_4_185/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd _360_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss FILLER_0_13_65/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ _343_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd _412_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ _274_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__292__I vss _098_ vdd ANTENNA__292__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ _326_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ _257_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd _309_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd ANTENNA__197__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss FILLER_0_15_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__301__A2 vss _098_ vdd ANTENNA__301__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 ctlp[6] net23 vdd vss output23/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss output34/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss output45/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss output12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss FILLER_0_5_109/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss FILLER_0_17_226/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss FILLER_0_4_197/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ _290_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss FILLER_0_9_223/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ _342_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd _411_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_273_ vss _090_ state\[0\] vdd _273_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout80 vss net80 net81 vdd fanout80/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_78 vdd vss FILLER_0_10_78/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_325_ vdd vss _130_ _118_ _129_ _325_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ _256_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ _308_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss FILLER_0_1_98/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ _239_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss FILLER_0_12_124/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss FILLER_0_8_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 ctln[6] net13 vdd vss output13/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss output35/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss FILLER_0_18_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput24 ctlp[7] net24 vdd vss output24/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss output46/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss FILLER_0_7_162/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss FILLER_0_7_195/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd ANTENNA_input1_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd ANTENNA__414__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ _341_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss _410_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ _272_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd fanout70/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_324_ vdd vss _129_ calibrate _062_ _324_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout81 vss net81 net82 vdd fanout81/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_255_ _076_ vss vdd _057_ _255_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output40_I vss net40 vdd ANTENNA_output40_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__304__A1 vss _093_ vdd ANTENNA__304__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_55 vdd vss FILLER_0_19_55/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_307_ vdd vss _114_ _113_ _096_ _307_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] _238_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss FILLER_0_21_125/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss FILLER_0_16_89/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss FILLER_0_12_136/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput36 result[9] net36 vdd vss output36/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 ctlp[8] net25 vdd vss output25/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss output47/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss output14/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss FILLER_0_4_144/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss FILLER_0_4_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd _340_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ _271_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd ANTENNA__356__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__200__I vss net20 vdd ANTENNA__200__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd ANTENNA_fanout52_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss FILLER_0_10_256/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss FILLER_0_6_239/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_99 vdd vss FILLER_0_4_99/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout60 net60 vss vdd net61 fanout60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout71 vss net71 net73 vdd fanout71/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ _254_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_323_ vss _015_ _128_ vdd _323_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd fanout82/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_306_ vss _113_ _057_ vdd _306_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_237_ vdd vss net40 net45 _237_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_57 vdd vss FILLER_0_16_57/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss output26/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss output15/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss output48/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss output37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss FILLER_0_17_218/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss FILLER_0_4_123/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd ANTENNA__203__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ _270_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ _399_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ _322_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd fanout61/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd fanout72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout50 net50 vss vdd net52 fanout50/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_37 vdd vss FILLER_0_10_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] _253_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_236_ net40 vss vdd _064_ _236_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_305_ vdd vss _112_ net1 _081_ _305_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__206__I vss net22 vdd ANTENNA__206__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss FILLER_0_20_193/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd _219_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss output27/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss output16/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss output38/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss FILLER_0_16_241/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd _398_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_214 vdd vss FILLER_0_10_214/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vdd vss FILLER_0_10_247/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__209__I vss net23 vdd ANTENNA__209__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_91 vdd vss FILLER_0_14_91/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ _321_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_output19_I vss net19 vdd ANTENNA_output19_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss FILLER_0_19_47/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd fanout73/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout51 vss net51 net52 vdd fanout51/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_252_ vdd vss cal_itt\[0\] _073_ _252_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout62 net62 vss vdd net64 fanout62/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_100 vdd vss FILLER_0_18_100/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss FILLER_0_18_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ _304_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] _235_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd _218_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss FILLER_0_16_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss output17/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss output39/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss output28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss FILLER_0_13_212/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ _397_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss FILLER_0_14_81/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ _320_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xfanout63 net63 vss vdd net64 fanout63/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_28 vdd vss FILLER_0_10_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout52 net52 vss vdd net57 fanout52/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ _251_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout74 vss net74 net82 vdd fanout74/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_449_ _038_ en_co_clk net55 vss net72 vdd _449_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ _303_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd _234_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_181 vdd vss FILLER_0_14_181/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_217_ vss net26 _052_ vdd _217_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput18 ctlp[1] net18 vdd vss output18/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss output29/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd ANTENNA_fanout80_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ _396_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_250_ vss _072_ _071_ vdd _250_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout53 net53 vss vdd net56 fanout53/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout75 vss net75 net76 vdd fanout75/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd fanout64/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd _448_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ _379_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__216__A2 vss net36 vdd ANTENNA__216__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_302_ vdd vss _012_ _093_ _110_ _302_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss FILLER_0_21_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_233_ vss net39 _063_ vdd _233_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss FILLER_0_15_116/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd ANTENNA__373__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_146 vdd vss FILLER_0_7_146/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ vdd vss _052_ mask\[9\] net36 _216_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput19 ctlp[2] net19 vdd vss output19/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss FILLER_0_7_59/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss FILLER_0_16_255/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss FILLER_0_0_130/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss FILLER_0_8_263/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss FILLER_0_14_50/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ _395_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss FILLER_0_4_49/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 fanout54/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd fanout76/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd fanout65/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss FILLER_0_19_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_378_ vdd vss _033_ _160_ _165_ _378_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_2 vdd vss FILLER_0_3_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd _447_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ _301_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd ANTENNA_output17_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] _232_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd _215_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss FILLER_0_11_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss FILLER_0_2_93/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss FILLER_0_17_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss FILLER_0_3_172/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd ANTENNA_output47_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] _394_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 fanout55/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss FILLER_0_5_212/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd fanout77/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ _377_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout66 vss net66 net68 vdd fanout66/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd _446_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_300_ vdd vss _011_ _104_ _109_ _300_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ _231_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd _429_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd input1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd _214_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss FILLER_0_7_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss FILLER_0_4_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss FILLER_0_24_290/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss FILLER_0_15_290/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss FILLER_0_0_198/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ _393_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd fanout78/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd fanout56/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd fanout67/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_376_ vss _164_ _163_ vdd _376_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd _445_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_72 vdd vss FILLER_0_5_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_230_ vdd vss _062_ _060_ _061_ _230_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_428_ _017_ state\[2\] net53 vss net70 vdd _428_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ _359_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_11_64 vdd vss FILLER_0_11_64/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 vss net2 clk vdd input2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_177 vdd vss FILLER_0_20_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output22_I vss net22 vdd ANTENNA_output22_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 _213_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_206 vdd vss FILLER_0_13_206/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss FILLER_0_13_228/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss _392_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_2 vdd vss FILLER_0_12_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__282__I vss _098_ vdd ANTENNA__282__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout57 vss net57 net65 vdd fanout57/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout79 vss net79 net81 vdd fanout79/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout68 vss net68 net69 vdd fanout68/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd _444_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] _375_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_18_139 vdd vss FILLER_0_18_139/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__277__I vss _093_ vdd ANTENNA__277__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_427_ _016_ state\[1\] net53 vdd vss net70 _427_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_17_161 vdd vss FILLER_0_17_161/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_358_ vdd vss _053_ _151_ _358_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd ANTENNA__385__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ _289_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd input3/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd _212_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd ANTENNA_output15_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss FILLER_0_22_86/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss FILLER_0_11_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss FILLER_0_17_64/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss FILLER_0_3_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ _391_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout58 net58 vss vdd net59 fanout58/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout69 vss net69 net74 vdd fanout69/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd _443_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_374_ vdd _061_ _056_ _162_ calibrate vss _374_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_107 vdd vss FILLER_0_18_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd ANTENNA__394__A3/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ _288_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ _357_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 vss net4 en vdd input4/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_426_ _015_ state\[0\] net64 vss net81 vdd _426_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_211_ vss net24 _050_ vdd _211_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ _409_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_124 vdd vss FILLER_0_11_124/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_135 vdd vss FILLER_0_11_135/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss FILLER_0_15_282/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd ANTENNA__413__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ _390_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss FILLER_0_14_99/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 fanout59/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ _373_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd _442_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ _287_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ _356_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss FILLER_0_11_78/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd input5/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd _425_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 _210_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss FILLER_0_20_169/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] _408_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd _339_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd ANTENNA_output20_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss FILLER_0_21_286/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss FILLER_0_12_220/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss FILLER_0_8_247/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_206 vdd vss FILLER_0_5_206/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net49 vss vdd net50 fanout49/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ _372_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd _441_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_142 vdd vss FILLER_0_17_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__303__A2 vss _098_ vdd ANTENNA__303__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_54 vdd vss FILLER_0_5_54/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_286_ vdd vss _005_ _094_ _101_ _286_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_355_ vdd vss _149_ _026_ _355_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd _424_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_123 vdd vss FILLER_0_14_123/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ _338_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ _407_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ _269_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss FILLER_0_17_56/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd ANTENNA_input4_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd _440_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_371_ vss _032_ _159_ vdd _371_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_88 vdd vss FILLER_0_5_88/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_285_ net28 vdd vss _101_ mask\[1\] _099_ _285_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_423_ _012_ net35 net55 vss net72 vdd _423_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ _354_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_199_ net20 vss vdd _046_ _199_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ _337_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] _406_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ _268_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss FILLER_0_24_274/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ _370_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd ANTENNA_fanout55_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss FILLER_0_1_266/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_284_ vdd vss _004_ _094_ _100_ _284_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_422_ _011_ net34 net61 vss net78 vdd _422_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output36_I vss net36 vdd ANTENNA_output36_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_353_ vdd vss _148_ _025_ _353_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss FILLER_0_17_133/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_336_ vdd vss _138_ _018_ _336_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_198_ vdd vss _046_ mask\[3\] net30 _198_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] _405_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] _267_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss FILLER_0_6_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ _319_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss FILLER_0_8_239/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss FILLER_0_1_212/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd _421_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ _283_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ _352_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_142 vdd vss FILLER_0_9_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_266_ vdd vss _055_ _085_ _266_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ _335_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_107 vdd vss FILLER_0_20_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ _404_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_197_ vdd vss net19 net9 _197_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd _249_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_318_ vdd vss _124_ _115_ _118_ _318_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__409__A1 vss cal_count\[3\] vdd ANTENNA__409__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_24 vdd vss FILLER_0_8_24/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd ANTENNA__251__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss FILLER_0_8_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd ANTENNA_input2_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd _420_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ _351_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd _282_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd ANTENNA__390__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_403_ vdd vss _183_ cal_count\[2\] _176_ _403_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_334_ vss _137_ _132_ vdd _334_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_90 vdd vss FILLER_0_6_90/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output41_I vss net41 vdd ANTENNA_output41_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_196_ net19 vss vdd _045_ _196_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ _265_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd ANTENNA__395__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ vss _070_ _069_ vdd _248_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_38 vdd vss FILLER_0_17_38/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__409__A2 vss _077_ vdd ANTENNA__409__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd _317_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss FILLER_0_2_171/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss FILLER_0_12_236/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ _350_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ _281_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd ANTENNA__237__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd _333_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 _195_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] _402_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss FILLER_0_11_109/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] _264_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd ANTENNA__372__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss FILLER_0_12_50/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ _247_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate _316_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_212 vdd vss FILLER_0_15_212/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_60 vdd vss FILLER_0_23_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vss FILLER_0_8_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_72 vdd vss FILLER_0_15_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss FILLER_0_17_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_204 vdd vss FILLER_0_1_204/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ _280_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss FILLER_0_14_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_332_ _126_ vdd vss _017_ _127_ _135_ _332_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_401_ vdd _180_ _179_ _181_ _174_ vss _401_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_194_ vss net8 net18 vdd _194_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ _263_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss FILLER_0_5_181/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss _315_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_246_ vss _068_ _055_ vdd _246_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_290 vdd vss FILLER_0_23_290/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss FILLER_0_15_235/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ _229_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss FILLER_0_18_61/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss FILLER_0_11_282/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd ANTENNA_fanout76_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss FILLER_0_4_213/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_193_ net18 vss vdd _044_ _193_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_400_ vdd vss _180_ cal_count\[1\] _178_ _400_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_331_ _134_ vdd vss _135_ _086_ _132_ _331_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ _262_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd ANTENNA__303__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_245_ vdd vss net6 _067_ net67 _245_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_314_ vdd vss _121_ _085_ _069_ _314_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_206 vdd vss FILLER_0_21_206/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd _228_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss FILLER_0_7_233/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss FILLER_0_9_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_261_ vss _081_ _059_ vdd _261_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_192_ vdd vss _044_ mask\[1\] net28 _192_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_142 vdd vss FILLER_0_13_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_330_ vdd vss _134_ _133_ _062_ _330_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss FILLER_0_12_20/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss FILLER_0_5_172/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ vdd vss _120_ _059_ _119_ _313_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__190__I vss _043_ vdd ANTENNA__190__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_244_ vdd vss en_co_clk _067_ _244_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__257__A1 vss _053_ vdd ANTENNA__257__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd _227_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd ANTENNA__402__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss FILLER_0_20_31/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss FILLER_0_9_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss FILLER_0_0_96/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss _260_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ _389_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 _191_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_243_ vdd vss net47 net42 _243_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ _312_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_282 vdd vss FILLER_0_23_282/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss FILLER_0_15_205/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss FILLER_0_2_165/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss FILLER_0_18_53/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ _226_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd ANTENNA__426__CLK/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_87 vdd vss FILLER_0_20_87/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_98 vdd vss FILLER_0_20_98/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 _209_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss FILLER_0_19_171/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd ANTENNA__302__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss FILLER_0_15_10/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss FILLER_0_15_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss FILLER_0_22_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss FILLER_0_13_100/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss FILLER_0_9_105/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ _190_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ _388_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd ANTENNA_output18_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_242_ net47 vss vdd _066_ _242_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ _311_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_15_228 vdd vss FILLER_0_15_228/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss FILLER_0_2_111/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss FILLER_0_2_177/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd _225_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss FILLER_0_18_76/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ _208_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd _387_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_164 vdd vss FILLER_0_5_164/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_310_ _090_ vdd vss _117_ _060_ _113_ _310_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_88 vdd vss FILLER_0_23_88/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss FILLER_0_23_44/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd _439_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] _241_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_101 vdd vss FILLER_0_2_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss FILLER_0_3_54/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd _224_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd vss _049_ mask\[6\] net33 _207_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss FILLER_0_19_195/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss FILLER_0_0_232/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss FILLER_0_16_154/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd ANTENNA__257__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd ANTENNA__220__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss FILLER_0_20_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ _386_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss FILLER_0_5_198/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vdd vss FILLER_0_17_282/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_240_ vdd vss net41 net46 _240_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_274 vdd vss FILLER_0_23_274/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd _438_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ _369_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd ANTENNA_output23_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss FILLER_0_14_263/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] _223_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss FILLER_0_9_290/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 _206_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss FILLER_0_0_266/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss _385_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ _299_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd _437_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_368_ vdd vss trim_mask\[4\] _158_ _368_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_78 vdd vss FILLER_0_3_78/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_222_ vdd vss net38 net43 _222_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ _205_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss FILLER_0_19_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd _453_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ _384_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss FILLER_0_10_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ _298_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd _436_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd ANTENNA__408__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ _367_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss FILLER_0_13_80/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss FILLER_0_1_192/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_221_ vss net38 _054_ vdd _221_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_270 vdd vss FILLER_0_9_270/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_419_ _008_ net31 net60 vss net77 vdd _419_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 _204_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss FILLER_0_20_15/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss FILLER_0_19_187/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss FILLER_0_3_221/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss FILLER_0_15_59/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_79 vdd vss FILLER_0_6_79/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout58_I vss net59 vdd ANTENNA_fanout58_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 _452_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ _383_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd _435_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ _297_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__408__A2 vss cal_count\[3\] vdd ANTENNA__408__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_127 vdd vss FILLER_0_2_127/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_366_ vdd vss trim_mask\[3\] _157_ _366_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_37 vdd vss FILLER_0_18_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_220_ vdd vss _054_ trim_val\[0\] _053_ _220_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_282 vdd vss FILLER_0_9_282/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_418_ _007_ net30 net60 vss net77 vdd _418_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_349_ vdd vss _146_ _023_ _349_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output21_I vss net21 vdd ANTENNA_output21_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 _203_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss FILLER_0_19_155/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss FILLER_0_19_111/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss FILLER_0_22_128/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss FILLER_0_15_180/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss FILLER_0_21_150/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss FILLER_0_6_47/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_28 vdd vss FILLER_0_12_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 _451_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_382_ vdd vss _035_ _160_ _167_ _382_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss FILLER_0_18_209/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss FILLER_0_5_136/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ _296_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd _434_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ _365_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd ANTENNA__280__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd ANTENNA__240__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_279_ vdd vss _096_ _090_ state\[1\] _279_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ _348_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd _417_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_231 vdd vss FILLER_0_6_231/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ _202_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_91 vdd vss FILLER_0_4_91/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output14_I vss net14 vdd ANTENNA_output14_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_94 vdd vss FILLER_0_10_94/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss FILLER_0_3_212/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss FILLER_0_19_134/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss FILLER_0_16_115/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss FILLER_0_22_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss FILLER_0_21_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss FILLER_0_6_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__243__I vss net47 vdd ANTENNA__243__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I vss rstn vdd ANTENNA_input5_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_156 vdd vss FILLER_0_8_156/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 _450_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ _381_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput40 trim[2] net40 vdd vss output40/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_148 vdd vss FILLER_0_5_148/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd _433_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ _295_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ _364_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss FILLER_0_14_235/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss FILLER_0_13_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_416_ _005_ net28 net62 vss net79 vdd _416_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_13_290 vdd vss FILLER_0_13_290/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_347_ vdd vss _145_ _022_ _347_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 _278_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_201_ vdd vss _047_ mask\[4\] net31 _201_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd ANTENNA__448__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_196 vdd vss FILLER_0_12_196/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 result[3] net30 vdd vss output30/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput6 clkc net6 vdd vss output6/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss output41/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ _380_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
.ends

