magic
tech gf180mcuD
magscale 1 10
timestamp 1701760198
<< checkpaint >>
rect -2319 -2356 2319 2356
<< nwell >>
rect -319 -356 319 356
<< mvpmos >>
rect -55 -100 55 100
<< mvpdiff >>
rect -143 87 -55 100
rect -143 -87 -130 87
rect -84 -87 -55 87
rect -143 -100 -55 -87
rect 55 87 143 100
rect 55 -87 84 87
rect 130 -87 143 87
rect 55 -100 143 -87
<< mvpdiffc >>
rect -130 -87 -84 87
rect 84 -87 130 87
<< mvnsubdiff >>
rect -287 252 287 324
rect -287 -252 -215 252
rect 215 -252 287 252
rect -287 -265 287 -252
rect -287 -311 -171 -265
rect 171 -311 287 -265
rect -287 -324 287 -311
<< mvnsubdiffcont >>
rect -171 -311 171 -265
<< polysilicon >>
rect -55 179 55 192
rect -55 133 -42 179
rect 42 133 55 179
rect -55 100 55 133
rect -55 -183 55 -100
<< polycontact >>
rect -42 133 42 179
<< metal1 >>
rect -53 133 -42 179
rect 42 133 53 179
rect -130 87 -84 83
rect -130 -98 -84 -102
rect 84 87 130 83
rect 84 -98 130 -102
<< labels >>
flabel metal1 0 31 0 31 0 FreeSans 240 0 0 0 G
<< properties >>
string FIXED_BBOX -251 -288 251 288
<< end >>


