** sch_path: /home/oe23ranan/gf_analog/xschem/sar_10b/dac/dac.sch
**.subckt dac out sample vdd vss vin
*+ ctl[9],ctl[8],ctl[7],ctl[6],ctl[5],ctl[4],ctl[3],ctl[2],ctl[1],ctl[0] dum
*.ipin vin
*.ipin sample
*.opin out
*.ipin ctl[9],ctl[8],ctl[7],ctl[6],ctl[5],ctl[4],ctl[3],ctl[2],ctl[1],ctl[0]
*.ipin dum
*.iopin vdd
*.iopin vss
xca out n6 n0 n5 n4 n2 ndum n3 n1 n7 n8 n9 carray
xswt out sample vdd vin vss bootstrapped_sw_hv
xidum dum vss vss vdd vdd ndum sky130_fd_sc_hd__inv_2
xi0 ctl[0] vss vss vdd vdd n0 sky130_fd_sc_hd__inv_2
xi1 ctl[1] vss vss vdd vdd n1 sky130_fd_sc_hd__inv_2
xi2 ctl[2] vss vss vdd vdd n2 sky130_fd_sc_hd__inv_2
xi3 ctl[3] vss vss vdd vdd n3 sky130_fd_sc_hd__inv_2
xi4 ctl[4] vss vss vdd vdd n4 sky130_fd_sc_hd__inv_2
xi5 ctl[5] vss vss vdd vdd n5 sky130_fd_sc_hd__inv_2
xi6 ctl[6] vss vss vdd vdd n6 sky130_fd_sc_hd__inv_2
xi7 ctl[7] vss vss vdd vdd n7 sky130_fd_sc_hd__inv_2
xi8 ctl[8] vss vss vdd vdd n8 sky130_fd_sc_hd__inv_2
xi9 ctl[9] vss vss vdd vdd n9 sky130_fd_sc_hd__inv_2
**.ends

* expanding   symbol:  sar_10b/dac/carray.sym # of pins=12
** sym_path: /home/oe23ranan/gf_analog/xschem/sar_10b/dac/carray.sym
** sch_path: /home/oe23ranan/gf_analog/xschem/sar_10b/dac/carray.sch
.subckt carray top n6 n0 n5 n4 n2 ndum n3 n1 n7 n8 n9
*.iopin top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
*.iopin n8
*.iopin n9
xcdum top ndum unitcap
xc0 top n0 unitcap
xc1[1] top n1 unitcap
xc1[0] top n1 unitcap
xc2[3] top n2 unitcap
xc2[2] top n2 unitcap
xc2[1] top n2 unitcap
xc2[0] top n2 unitcap
xc3[7] top n3 unitcap
xc3[6] top n3 unitcap
xc3[5] top n3 unitcap
xc3[4] top n3 unitcap
xc3[3] top n3 unitcap
xc3[2] top n3 unitcap
xc3[1] top n3 unitcap
xc3[0] top n3 unitcap
xc4[15] top n4 unitcap
xc4[14] top n4 unitcap
xc4[13] top n4 unitcap
xc4[12] top n4 unitcap
xc4[11] top n4 unitcap
xc4[10] top n4 unitcap
xc4[9] top n4 unitcap
xc4[8] top n4 unitcap
xc4[7] top n4 unitcap
xc4[6] top n4 unitcap
xc4[5] top n4 unitcap
xc4[4] top n4 unitcap
xc4[3] top n4 unitcap
xc4[2] top n4 unitcap
xc4[1] top n4 unitcap
xc4[0] top n4 unitcap
xc5[31] top n5 unitcap
xc5[30] top n5 unitcap
xc5[29] top n5 unitcap
xc5[28] top n5 unitcap
xc5[27] top n5 unitcap
xc5[26] top n5 unitcap
xc5[25] top n5 unitcap
xc5[24] top n5 unitcap
xc5[23] top n5 unitcap
xc5[22] top n5 unitcap
xc5[21] top n5 unitcap
xc5[20] top n5 unitcap
xc5[19] top n5 unitcap
xc5[18] top n5 unitcap
xc5[17] top n5 unitcap
xc5[16] top n5 unitcap
xc5[15] top n5 unitcap
xc5[14] top n5 unitcap
xc5[13] top n5 unitcap
xc5[12] top n5 unitcap
xc5[11] top n5 unitcap
xc5[10] top n5 unitcap
xc5[9] top n5 unitcap
xc5[8] top n5 unitcap
xc5[7] top n5 unitcap
xc5[6] top n5 unitcap
xc5[5] top n5 unitcap
xc5[4] top n5 unitcap
xc5[3] top n5 unitcap
xc5[2] top n5 unitcap
xc5[1] top n5 unitcap
xc5[0] top n5 unitcap
xc6[63] top n6 unitcap
xc6[62] top n6 unitcap
xc6[61] top n6 unitcap
xc6[60] top n6 unitcap
xc6[59] top n6 unitcap
xc6[58] top n6 unitcap
xc6[57] top n6 unitcap
xc6[56] top n6 unitcap
xc6[55] top n6 unitcap
xc6[54] top n6 unitcap
xc6[53] top n6 unitcap
xc6[52] top n6 unitcap
xc6[51] top n6 unitcap
xc6[50] top n6 unitcap
xc6[49] top n6 unitcap
xc6[48] top n6 unitcap
xc6[47] top n6 unitcap
xc6[46] top n6 unitcap
xc6[45] top n6 unitcap
xc6[44] top n6 unitcap
xc6[43] top n6 unitcap
xc6[42] top n6 unitcap
xc6[41] top n6 unitcap
xc6[40] top n6 unitcap
xc6[39] top n6 unitcap
xc6[38] top n6 unitcap
xc6[37] top n6 unitcap
xc6[36] top n6 unitcap
xc6[35] top n6 unitcap
xc6[34] top n6 unitcap
xc6[33] top n6 unitcap
xc6[32] top n6 unitcap
xc6[31] top n6 unitcap
xc6[30] top n6 unitcap
xc6[29] top n6 unitcap
xc6[28] top n6 unitcap
xc6[27] top n6 unitcap
xc6[26] top n6 unitcap
xc6[25] top n6 unitcap
xc6[24] top n6 unitcap
xc6[23] top n6 unitcap
xc6[22] top n6 unitcap
xc6[21] top n6 unitcap
xc6[20] top n6 unitcap
xc6[19] top n6 unitcap
xc6[18] top n6 unitcap
xc6[17] top n6 unitcap
xc6[16] top n6 unitcap
xc6[15] top n6 unitcap
xc6[14] top n6 unitcap
xc6[13] top n6 unitcap
xc6[12] top n6 unitcap
xc6[11] top n6 unitcap
xc6[10] top n6 unitcap
xc6[9] top n6 unitcap
xc6[8] top n6 unitcap
xc6[7] top n6 unitcap
xc6[6] top n6 unitcap
xc6[5] top n6 unitcap
xc6[4] top n6 unitcap
xc6[3] top n6 unitcap
xc6[2] top n6 unitcap
xc6[1] top n6 unitcap
xc6[0] top n6 unitcap
xc7[127] top n7 unitcap
xc7[126] top n7 unitcap
xc7[125] top n7 unitcap
xc7[124] top n7 unitcap
xc7[123] top n7 unitcap
xc7[122] top n7 unitcap
xc7[121] top n7 unitcap
xc7[120] top n7 unitcap
xc7[119] top n7 unitcap
xc7[118] top n7 unitcap
xc7[117] top n7 unitcap
xc7[116] top n7 unitcap
xc7[115] top n7 unitcap
xc7[114] top n7 unitcap
xc7[113] top n7 unitcap
xc7[112] top n7 unitcap
xc7[111] top n7 unitcap
xc7[110] top n7 unitcap
xc7[109] top n7 unitcap
xc7[108] top n7 unitcap
xc7[107] top n7 unitcap
xc7[106] top n7 unitcap
xc7[105] top n7 unitcap
xc7[104] top n7 unitcap
xc7[103] top n7 unitcap
xc7[102] top n7 unitcap
xc7[101] top n7 unitcap
xc7[100] top n7 unitcap
xc7[99] top n7 unitcap
xc7[98] top n7 unitcap
xc7[97] top n7 unitcap
xc7[96] top n7 unitcap
xc7[95] top n7 unitcap
xc7[94] top n7 unitcap
xc7[93] top n7 unitcap
xc7[92] top n7 unitcap
xc7[91] top n7 unitcap
xc7[90] top n7 unitcap
xc7[89] top n7 unitcap
xc7[88] top n7 unitcap
xc7[87] top n7 unitcap
xc7[86] top n7 unitcap
xc7[85] top n7 unitcap
xc7[84] top n7 unitcap
xc7[83] top n7 unitcap
xc7[82] top n7 unitcap
xc7[81] top n7 unitcap
xc7[80] top n7 unitcap
xc7[79] top n7 unitcap
xc7[78] top n7 unitcap
xc7[77] top n7 unitcap
xc7[76] top n7 unitcap
xc7[75] top n7 unitcap
xc7[74] top n7 unitcap
xc7[73] top n7 unitcap
xc7[72] top n7 unitcap
xc7[71] top n7 unitcap
xc7[70] top n7 unitcap
xc7[69] top n7 unitcap
xc7[68] top n7 unitcap
xc7[67] top n7 unitcap
xc7[66] top n7 unitcap
xc7[65] top n7 unitcap
xc7[64] top n7 unitcap
xc7[63] top n7 unitcap
xc7[62] top n7 unitcap
xc7[61] top n7 unitcap
xc7[60] top n7 unitcap
xc7[59] top n7 unitcap
xc7[58] top n7 unitcap
xc7[57] top n7 unitcap
xc7[56] top n7 unitcap
xc7[55] top n7 unitcap
xc7[54] top n7 unitcap
xc7[53] top n7 unitcap
xc7[52] top n7 unitcap
xc7[51] top n7 unitcap
xc7[50] top n7 unitcap
xc7[49] top n7 unitcap
xc7[48] top n7 unitcap
xc7[47] top n7 unitcap
xc7[46] top n7 unitcap
xc7[45] top n7 unitcap
xc7[44] top n7 unitcap
xc7[43] top n7 unitcap
xc7[42] top n7 unitcap
xc7[41] top n7 unitcap
xc7[40] top n7 unitcap
xc7[39] top n7 unitcap
xc7[38] top n7 unitcap
xc7[37] top n7 unitcap
xc7[36] top n7 unitcap
xc7[35] top n7 unitcap
xc7[34] top n7 unitcap
xc7[33] top n7 unitcap
xc7[32] top n7 unitcap
xc7[31] top n7 unitcap
xc7[30] top n7 unitcap
xc7[29] top n7 unitcap
xc7[28] top n7 unitcap
xc7[27] top n7 unitcap
xc7[26] top n7 unitcap
xc7[25] top n7 unitcap
xc7[24] top n7 unitcap
xc7[23] top n7 unitcap
xc7[22] top n7 unitcap
xc7[21] top n7 unitcap
xc7[20] top n7 unitcap
xc7[19] top n7 unitcap
xc7[18] top n7 unitcap
xc7[17] top n7 unitcap
xc7[16] top n7 unitcap
xc7[15] top n7 unitcap
xc7[14] top n7 unitcap
xc7[13] top n7 unitcap
xc7[12] top n7 unitcap
xc7[11] top n7 unitcap
xc7[10] top n7 unitcap
xc7[9] top n7 unitcap
xc7[8] top n7 unitcap
xc7[7] top n7 unitcap
xc7[6] top n7 unitcap
xc7[5] top n7 unitcap
xc7[4] top n7 unitcap
xc7[3] top n7 unitcap
xc7[2] top n7 unitcap
xc7[1] top n7 unitcap
xc7[0] top n7 unitcap
xc8[255] top n8 unitcap
xc8[254] top n8 unitcap
xc8[253] top n8 unitcap
xc8[252] top n8 unitcap
xc8[251] top n8 unitcap
xc8[250] top n8 unitcap
xc8[249] top n8 unitcap
xc8[248] top n8 unitcap
xc8[247] top n8 unitcap
xc8[246] top n8 unitcap
xc8[245] top n8 unitcap
xc8[244] top n8 unitcap
xc8[243] top n8 unitcap
xc8[242] top n8 unitcap
xc8[241] top n8 unitcap
xc8[240] top n8 unitcap
xc8[239] top n8 unitcap
xc8[238] top n8 unitcap
xc8[237] top n8 unitcap
xc8[236] top n8 unitcap
xc8[235] top n8 unitcap
xc8[234] top n8 unitcap
xc8[233] top n8 unitcap
xc8[232] top n8 unitcap
xc8[231] top n8 unitcap
xc8[230] top n8 unitcap
xc8[229] top n8 unitcap
xc8[228] top n8 unitcap
xc8[227] top n8 unitcap
xc8[226] top n8 unitcap
xc8[225] top n8 unitcap
xc8[224] top n8 unitcap
xc8[223] top n8 unitcap
xc8[222] top n8 unitcap
xc8[221] top n8 unitcap
xc8[220] top n8 unitcap
xc8[219] top n8 unitcap
xc8[218] top n8 unitcap
xc8[217] top n8 unitcap
xc8[216] top n8 unitcap
xc8[215] top n8 unitcap
xc8[214] top n8 unitcap
xc8[213] top n8 unitcap
xc8[212] top n8 unitcap
xc8[211] top n8 unitcap
xc8[210] top n8 unitcap
xc8[209] top n8 unitcap
xc8[208] top n8 unitcap
xc8[207] top n8 unitcap
xc8[206] top n8 unitcap
xc8[205] top n8 unitcap
xc8[204] top n8 unitcap
xc8[203] top n8 unitcap
xc8[202] top n8 unitcap
xc8[201] top n8 unitcap
xc8[200] top n8 unitcap
xc8[199] top n8 unitcap
xc8[198] top n8 unitcap
xc8[197] top n8 unitcap
xc8[196] top n8 unitcap
xc8[195] top n8 unitcap
xc8[194] top n8 unitcap
xc8[193] top n8 unitcap
xc8[192] top n8 unitcap
xc8[191] top n8 unitcap
xc8[190] top n8 unitcap
xc8[189] top n8 unitcap
xc8[188] top n8 unitcap
xc8[187] top n8 unitcap
xc8[186] top n8 unitcap
xc8[185] top n8 unitcap
xc8[184] top n8 unitcap
xc8[183] top n8 unitcap
xc8[182] top n8 unitcap
xc8[181] top n8 unitcap
xc8[180] top n8 unitcap
xc8[179] top n8 unitcap
xc8[178] top n8 unitcap
xc8[177] top n8 unitcap
xc8[176] top n8 unitcap
xc8[175] top n8 unitcap
xc8[174] top n8 unitcap
xc8[173] top n8 unitcap
xc8[172] top n8 unitcap
xc8[171] top n8 unitcap
xc8[170] top n8 unitcap
xc8[169] top n8 unitcap
xc8[168] top n8 unitcap
xc8[167] top n8 unitcap
xc8[166] top n8 unitcap
xc8[165] top n8 unitcap
xc8[164] top n8 unitcap
xc8[163] top n8 unitcap
xc8[162] top n8 unitcap
xc8[161] top n8 unitcap
xc8[160] top n8 unitcap
xc8[159] top n8 unitcap
xc8[158] top n8 unitcap
xc8[157] top n8 unitcap
xc8[156] top n8 unitcap
xc8[155] top n8 unitcap
xc8[154] top n8 unitcap
xc8[153] top n8 unitcap
xc8[152] top n8 unitcap
xc8[151] top n8 unitcap
xc8[150] top n8 unitcap
xc8[149] top n8 unitcap
xc8[148] top n8 unitcap
xc8[147] top n8 unitcap
xc8[146] top n8 unitcap
xc8[145] top n8 unitcap
xc8[144] top n8 unitcap
xc8[143] top n8 unitcap
xc8[142] top n8 unitcap
xc8[141] top n8 unitcap
xc8[140] top n8 unitcap
xc8[139] top n8 unitcap
xc8[138] top n8 unitcap
xc8[137] top n8 unitcap
xc8[136] top n8 unitcap
xc8[135] top n8 unitcap
xc8[134] top n8 unitcap
xc8[133] top n8 unitcap
xc8[132] top n8 unitcap
xc8[131] top n8 unitcap
xc8[130] top n8 unitcap
xc8[129] top n8 unitcap
xc8[128] top n8 unitcap
xc8[127] top n8 unitcap
xc8[126] top n8 unitcap
xc8[125] top n8 unitcap
xc8[124] top n8 unitcap
xc8[123] top n8 unitcap
xc8[122] top n8 unitcap
xc8[121] top n8 unitcap
xc8[120] top n8 unitcap
xc8[119] top n8 unitcap
xc8[118] top n8 unitcap
xc8[117] top n8 unitcap
xc8[116] top n8 unitcap
xc8[115] top n8 unitcap
xc8[114] top n8 unitcap
xc8[113] top n8 unitcap
xc8[112] top n8 unitcap
xc8[111] top n8 unitcap
xc8[110] top n8 unitcap
xc8[109] top n8 unitcap
xc8[108] top n8 unitcap
xc8[107] top n8 unitcap
xc8[106] top n8 unitcap
xc8[105] top n8 unitcap
xc8[104] top n8 unitcap
xc8[103] top n8 unitcap
xc8[102] top n8 unitcap
xc8[101] top n8 unitcap
xc8[100] top n8 unitcap
xc8[99] top n8 unitcap
xc8[98] top n8 unitcap
xc8[97] top n8 unitcap
xc8[96] top n8 unitcap
xc8[95] top n8 unitcap
xc8[94] top n8 unitcap
xc8[93] top n8 unitcap
xc8[92] top n8 unitcap
xc8[91] top n8 unitcap
xc8[90] top n8 unitcap
xc8[89] top n8 unitcap
xc8[88] top n8 unitcap
xc8[87] top n8 unitcap
xc8[86] top n8 unitcap
xc8[85] top n8 unitcap
xc8[84] top n8 unitcap
xc8[83] top n8 unitcap
xc8[82] top n8 unitcap
xc8[81] top n8 unitcap
xc8[80] top n8 unitcap
xc8[79] top n8 unitcap
xc8[78] top n8 unitcap
xc8[77] top n8 unitcap
xc8[76] top n8 unitcap
xc8[75] top n8 unitcap
xc8[74] top n8 unitcap
xc8[73] top n8 unitcap
xc8[72] top n8 unitcap
xc8[71] top n8 unitcap
xc8[70] top n8 unitcap
xc8[69] top n8 unitcap
xc8[68] top n8 unitcap
xc8[67] top n8 unitcap
xc8[66] top n8 unitcap
xc8[65] top n8 unitcap
xc8[64] top n8 unitcap
xc8[63] top n8 unitcap
xc8[62] top n8 unitcap
xc8[61] top n8 unitcap
xc8[60] top n8 unitcap
xc8[59] top n8 unitcap
xc8[58] top n8 unitcap
xc8[57] top n8 unitcap
xc8[56] top n8 unitcap
xc8[55] top n8 unitcap
xc8[54] top n8 unitcap
xc8[53] top n8 unitcap
xc8[52] top n8 unitcap
xc8[51] top n8 unitcap
xc8[50] top n8 unitcap
xc8[49] top n8 unitcap
xc8[48] top n8 unitcap
xc8[47] top n8 unitcap
xc8[46] top n8 unitcap
xc8[45] top n8 unitcap
xc8[44] top n8 unitcap
xc8[43] top n8 unitcap
xc8[42] top n8 unitcap
xc8[41] top n8 unitcap
xc8[40] top n8 unitcap
xc8[39] top n8 unitcap
xc8[38] top n8 unitcap
xc8[37] top n8 unitcap
xc8[36] top n8 unitcap
xc8[35] top n8 unitcap
xc8[34] top n8 unitcap
xc8[33] top n8 unitcap
xc8[32] top n8 unitcap
xc8[31] top n8 unitcap
xc8[30] top n8 unitcap
xc8[29] top n8 unitcap
xc8[28] top n8 unitcap
xc8[27] top n8 unitcap
xc8[26] top n8 unitcap
xc8[25] top n8 unitcap
xc8[24] top n8 unitcap
xc8[23] top n8 unitcap
xc8[22] top n8 unitcap
xc8[21] top n8 unitcap
xc8[20] top n8 unitcap
xc8[19] top n8 unitcap
xc8[18] top n8 unitcap
xc8[17] top n8 unitcap
xc8[16] top n8 unitcap
xc8[15] top n8 unitcap
xc8[14] top n8 unitcap
xc8[13] top n8 unitcap
xc8[12] top n8 unitcap
xc8[11] top n8 unitcap
xc8[10] top n8 unitcap
xc8[9] top n8 unitcap
xc8[8] top n8 unitcap
xc8[7] top n8 unitcap
xc8[6] top n8 unitcap
xc8[5] top n8 unitcap
xc8[4] top n8 unitcap
xc8[3] top n8 unitcap
xc8[2] top n8 unitcap
xc8[1] top n8 unitcap
xc8[0] top n8 unitcap
xc9[511] top n9 unitcap
xc9[510] top n9 unitcap
xc9[509] top n9 unitcap
xc9[508] top n9 unitcap
xc9[507] top n9 unitcap
xc9[506] top n9 unitcap
xc9[505] top n9 unitcap
xc9[504] top n9 unitcap
xc9[503] top n9 unitcap
xc9[502] top n9 unitcap
xc9[501] top n9 unitcap
xc9[500] top n9 unitcap
xc9[499] top n9 unitcap
xc9[498] top n9 unitcap
xc9[497] top n9 unitcap
xc9[496] top n9 unitcap
xc9[495] top n9 unitcap
xc9[494] top n9 unitcap
xc9[493] top n9 unitcap
xc9[492] top n9 unitcap
xc9[491] top n9 unitcap
xc9[490] top n9 unitcap
xc9[489] top n9 unitcap
xc9[488] top n9 unitcap
xc9[487] top n9 unitcap
xc9[486] top n9 unitcap
xc9[485] top n9 unitcap
xc9[484] top n9 unitcap
xc9[483] top n9 unitcap
xc9[482] top n9 unitcap
xc9[481] top n9 unitcap
xc9[480] top n9 unitcap
xc9[479] top n9 unitcap
xc9[478] top n9 unitcap
xc9[477] top n9 unitcap
xc9[476] top n9 unitcap
xc9[475] top n9 unitcap
xc9[474] top n9 unitcap
xc9[473] top n9 unitcap
xc9[472] top n9 unitcap
xc9[471] top n9 unitcap
xc9[470] top n9 unitcap
xc9[469] top n9 unitcap
xc9[468] top n9 unitcap
xc9[467] top n9 unitcap
xc9[466] top n9 unitcap
xc9[465] top n9 unitcap
xc9[464] top n9 unitcap
xc9[463] top n9 unitcap
xc9[462] top n9 unitcap
xc9[461] top n9 unitcap
xc9[460] top n9 unitcap
xc9[459] top n9 unitcap
xc9[458] top n9 unitcap
xc9[457] top n9 unitcap
xc9[456] top n9 unitcap
xc9[455] top n9 unitcap
xc9[454] top n9 unitcap
xc9[453] top n9 unitcap
xc9[452] top n9 unitcap
xc9[451] top n9 unitcap
xc9[450] top n9 unitcap
xc9[449] top n9 unitcap
xc9[448] top n9 unitcap
xc9[447] top n9 unitcap
xc9[446] top n9 unitcap
xc9[445] top n9 unitcap
xc9[444] top n9 unitcap
xc9[443] top n9 unitcap
xc9[442] top n9 unitcap
xc9[441] top n9 unitcap
xc9[440] top n9 unitcap
xc9[439] top n9 unitcap
xc9[438] top n9 unitcap
xc9[437] top n9 unitcap
xc9[436] top n9 unitcap
xc9[435] top n9 unitcap
xc9[434] top n9 unitcap
xc9[433] top n9 unitcap
xc9[432] top n9 unitcap
xc9[431] top n9 unitcap
xc9[430] top n9 unitcap
xc9[429] top n9 unitcap
xc9[428] top n9 unitcap
xc9[427] top n9 unitcap
xc9[426] top n9 unitcap
xc9[425] top n9 unitcap
xc9[424] top n9 unitcap
xc9[423] top n9 unitcap
xc9[422] top n9 unitcap
xc9[421] top n9 unitcap
xc9[420] top n9 unitcap
xc9[419] top n9 unitcap
xc9[418] top n9 unitcap
xc9[417] top n9 unitcap
xc9[416] top n9 unitcap
xc9[415] top n9 unitcap
xc9[414] top n9 unitcap
xc9[413] top n9 unitcap
xc9[412] top n9 unitcap
xc9[411] top n9 unitcap
xc9[410] top n9 unitcap
xc9[409] top n9 unitcap
xc9[408] top n9 unitcap
xc9[407] top n9 unitcap
xc9[406] top n9 unitcap
xc9[405] top n9 unitcap
xc9[404] top n9 unitcap
xc9[403] top n9 unitcap
xc9[402] top n9 unitcap
xc9[401] top n9 unitcap
xc9[400] top n9 unitcap
xc9[399] top n9 unitcap
xc9[398] top n9 unitcap
xc9[397] top n9 unitcap
xc9[396] top n9 unitcap
xc9[395] top n9 unitcap
xc9[394] top n9 unitcap
xc9[393] top n9 unitcap
xc9[392] top n9 unitcap
xc9[391] top n9 unitcap
xc9[390] top n9 unitcap
xc9[389] top n9 unitcap
xc9[388] top n9 unitcap
xc9[387] top n9 unitcap
xc9[386] top n9 unitcap
xc9[385] top n9 unitcap
xc9[384] top n9 unitcap
xc9[383] top n9 unitcap
xc9[382] top n9 unitcap
xc9[381] top n9 unitcap
xc9[380] top n9 unitcap
xc9[379] top n9 unitcap
xc9[378] top n9 unitcap
xc9[377] top n9 unitcap
xc9[376] top n9 unitcap
xc9[375] top n9 unitcap
xc9[374] top n9 unitcap
xc9[373] top n9 unitcap
xc9[372] top n9 unitcap
xc9[371] top n9 unitcap
xc9[370] top n9 unitcap
xc9[369] top n9 unitcap
xc9[368] top n9 unitcap
xc9[367] top n9 unitcap
xc9[366] top n9 unitcap
xc9[365] top n9 unitcap
xc9[364] top n9 unitcap
xc9[363] top n9 unitcap
xc9[362] top n9 unitcap
xc9[361] top n9 unitcap
xc9[360] top n9 unitcap
xc9[359] top n9 unitcap
xc9[358] top n9 unitcap
xc9[357] top n9 unitcap
xc9[356] top n9 unitcap
xc9[355] top n9 unitcap
xc9[354] top n9 unitcap
xc9[353] top n9 unitcap
xc9[352] top n9 unitcap
xc9[351] top n9 unitcap
xc9[350] top n9 unitcap
xc9[349] top n9 unitcap
xc9[348] top n9 unitcap
xc9[347] top n9 unitcap
xc9[346] top n9 unitcap
xc9[345] top n9 unitcap
xc9[344] top n9 unitcap
xc9[343] top n9 unitcap
xc9[342] top n9 unitcap
xc9[341] top n9 unitcap
xc9[340] top n9 unitcap
xc9[339] top n9 unitcap
xc9[338] top n9 unitcap
xc9[337] top n9 unitcap
xc9[336] top n9 unitcap
xc9[335] top n9 unitcap
xc9[334] top n9 unitcap
xc9[333] top n9 unitcap
xc9[332] top n9 unitcap
xc9[331] top n9 unitcap
xc9[330] top n9 unitcap
xc9[329] top n9 unitcap
xc9[328] top n9 unitcap
xc9[327] top n9 unitcap
xc9[326] top n9 unitcap
xc9[325] top n9 unitcap
xc9[324] top n9 unitcap
xc9[323] top n9 unitcap
xc9[322] top n9 unitcap
xc9[321] top n9 unitcap
xc9[320] top n9 unitcap
xc9[319] top n9 unitcap
xc9[318] top n9 unitcap
xc9[317] top n9 unitcap
xc9[316] top n9 unitcap
xc9[315] top n9 unitcap
xc9[314] top n9 unitcap
xc9[313] top n9 unitcap
xc9[312] top n9 unitcap
xc9[311] top n9 unitcap
xc9[310] top n9 unitcap
xc9[309] top n9 unitcap
xc9[308] top n9 unitcap
xc9[307] top n9 unitcap
xc9[306] top n9 unitcap
xc9[305] top n9 unitcap
xc9[304] top n9 unitcap
xc9[303] top n9 unitcap
xc9[302] top n9 unitcap
xc9[301] top n9 unitcap
xc9[300] top n9 unitcap
xc9[299] top n9 unitcap
xc9[298] top n9 unitcap
xc9[297] top n9 unitcap
xc9[296] top n9 unitcap
xc9[295] top n9 unitcap
xc9[294] top n9 unitcap
xc9[293] top n9 unitcap
xc9[292] top n9 unitcap
xc9[291] top n9 unitcap
xc9[290] top n9 unitcap
xc9[289] top n9 unitcap
xc9[288] top n9 unitcap
xc9[287] top n9 unitcap
xc9[286] top n9 unitcap
xc9[285] top n9 unitcap
xc9[284] top n9 unitcap
xc9[283] top n9 unitcap
xc9[282] top n9 unitcap
xc9[281] top n9 unitcap
xc9[280] top n9 unitcap
xc9[279] top n9 unitcap
xc9[278] top n9 unitcap
xc9[277] top n9 unitcap
xc9[276] top n9 unitcap
xc9[275] top n9 unitcap
xc9[274] top n9 unitcap
xc9[273] top n9 unitcap
xc9[272] top n9 unitcap
xc9[271] top n9 unitcap
xc9[270] top n9 unitcap
xc9[269] top n9 unitcap
xc9[268] top n9 unitcap
xc9[267] top n9 unitcap
xc9[266] top n9 unitcap
xc9[265] top n9 unitcap
xc9[264] top n9 unitcap
xc9[263] top n9 unitcap
xc9[262] top n9 unitcap
xc9[261] top n9 unitcap
xc9[260] top n9 unitcap
xc9[259] top n9 unitcap
xc9[258] top n9 unitcap
xc9[257] top n9 unitcap
xc9[256] top n9 unitcap
xc9[255] top n9 unitcap
xc9[254] top n9 unitcap
xc9[253] top n9 unitcap
xc9[252] top n9 unitcap
xc9[251] top n9 unitcap
xc9[250] top n9 unitcap
xc9[249] top n9 unitcap
xc9[248] top n9 unitcap
xc9[247] top n9 unitcap
xc9[246] top n9 unitcap
xc9[245] top n9 unitcap
xc9[244] top n9 unitcap
xc9[243] top n9 unitcap
xc9[242] top n9 unitcap
xc9[241] top n9 unitcap
xc9[240] top n9 unitcap
xc9[239] top n9 unitcap
xc9[238] top n9 unitcap
xc9[237] top n9 unitcap
xc9[236] top n9 unitcap
xc9[235] top n9 unitcap
xc9[234] top n9 unitcap
xc9[233] top n9 unitcap
xc9[232] top n9 unitcap
xc9[231] top n9 unitcap
xc9[230] top n9 unitcap
xc9[229] top n9 unitcap
xc9[228] top n9 unitcap
xc9[227] top n9 unitcap
xc9[226] top n9 unitcap
xc9[225] top n9 unitcap
xc9[224] top n9 unitcap
xc9[223] top n9 unitcap
xc9[222] top n9 unitcap
xc9[221] top n9 unitcap
xc9[220] top n9 unitcap
xc9[219] top n9 unitcap
xc9[218] top n9 unitcap
xc9[217] top n9 unitcap
xc9[216] top n9 unitcap
xc9[215] top n9 unitcap
xc9[214] top n9 unitcap
xc9[213] top n9 unitcap
xc9[212] top n9 unitcap
xc9[211] top n9 unitcap
xc9[210] top n9 unitcap
xc9[209] top n9 unitcap
xc9[208] top n9 unitcap
xc9[207] top n9 unitcap
xc9[206] top n9 unitcap
xc9[205] top n9 unitcap
xc9[204] top n9 unitcap
xc9[203] top n9 unitcap
xc9[202] top n9 unitcap
xc9[201] top n9 unitcap
xc9[200] top n9 unitcap
xc9[199] top n9 unitcap
xc9[198] top n9 unitcap
xc9[197] top n9 unitcap
xc9[196] top n9 unitcap
xc9[195] top n9 unitcap
xc9[194] top n9 unitcap
xc9[193] top n9 unitcap
xc9[192] top n9 unitcap
xc9[191] top n9 unitcap
xc9[190] top n9 unitcap
xc9[189] top n9 unitcap
xc9[188] top n9 unitcap
xc9[187] top n9 unitcap
xc9[186] top n9 unitcap
xc9[185] top n9 unitcap
xc9[184] top n9 unitcap
xc9[183] top n9 unitcap
xc9[182] top n9 unitcap
xc9[181] top n9 unitcap
xc9[180] top n9 unitcap
xc9[179] top n9 unitcap
xc9[178] top n9 unitcap
xc9[177] top n9 unitcap
xc9[176] top n9 unitcap
xc9[175] top n9 unitcap
xc9[174] top n9 unitcap
xc9[173] top n9 unitcap
xc9[172] top n9 unitcap
xc9[171] top n9 unitcap
xc9[170] top n9 unitcap
xc9[169] top n9 unitcap
xc9[168] top n9 unitcap
xc9[167] top n9 unitcap
xc9[166] top n9 unitcap
xc9[165] top n9 unitcap
xc9[164] top n9 unitcap
xc9[163] top n9 unitcap
xc9[162] top n9 unitcap
xc9[161] top n9 unitcap
xc9[160] top n9 unitcap
xc9[159] top n9 unitcap
xc9[158] top n9 unitcap
xc9[157] top n9 unitcap
xc9[156] top n9 unitcap
xc9[155] top n9 unitcap
xc9[154] top n9 unitcap
xc9[153] top n9 unitcap
xc9[152] top n9 unitcap
xc9[151] top n9 unitcap
xc9[150] top n9 unitcap
xc9[149] top n9 unitcap
xc9[148] top n9 unitcap
xc9[147] top n9 unitcap
xc9[146] top n9 unitcap
xc9[145] top n9 unitcap
xc9[144] top n9 unitcap
xc9[143] top n9 unitcap
xc9[142] top n9 unitcap
xc9[141] top n9 unitcap
xc9[140] top n9 unitcap
xc9[139] top n9 unitcap
xc9[138] top n9 unitcap
xc9[137] top n9 unitcap
xc9[136] top n9 unitcap
xc9[135] top n9 unitcap
xc9[134] top n9 unitcap
xc9[133] top n9 unitcap
xc9[132] top n9 unitcap
xc9[131] top n9 unitcap
xc9[130] top n9 unitcap
xc9[129] top n9 unitcap
xc9[128] top n9 unitcap
xc9[127] top n9 unitcap
xc9[126] top n9 unitcap
xc9[125] top n9 unitcap
xc9[124] top n9 unitcap
xc9[123] top n9 unitcap
xc9[122] top n9 unitcap
xc9[121] top n9 unitcap
xc9[120] top n9 unitcap
xc9[119] top n9 unitcap
xc9[118] top n9 unitcap
xc9[117] top n9 unitcap
xc9[116] top n9 unitcap
xc9[115] top n9 unitcap
xc9[114] top n9 unitcap
xc9[113] top n9 unitcap
xc9[112] top n9 unitcap
xc9[111] top n9 unitcap
xc9[110] top n9 unitcap
xc9[109] top n9 unitcap
xc9[108] top n9 unitcap
xc9[107] top n9 unitcap
xc9[106] top n9 unitcap
xc9[105] top n9 unitcap
xc9[104] top n9 unitcap
xc9[103] top n9 unitcap
xc9[102] top n9 unitcap
xc9[101] top n9 unitcap
xc9[100] top n9 unitcap
xc9[99] top n9 unitcap
xc9[98] top n9 unitcap
xc9[97] top n9 unitcap
xc9[96] top n9 unitcap
xc9[95] top n9 unitcap
xc9[94] top n9 unitcap
xc9[93] top n9 unitcap
xc9[92] top n9 unitcap
xc9[91] top n9 unitcap
xc9[90] top n9 unitcap
xc9[89] top n9 unitcap
xc9[88] top n9 unitcap
xc9[87] top n9 unitcap
xc9[86] top n9 unitcap
xc9[85] top n9 unitcap
xc9[84] top n9 unitcap
xc9[83] top n9 unitcap
xc9[82] top n9 unitcap
xc9[81] top n9 unitcap
xc9[80] top n9 unitcap
xc9[79] top n9 unitcap
xc9[78] top n9 unitcap
xc9[77] top n9 unitcap
xc9[76] top n9 unitcap
xc9[75] top n9 unitcap
xc9[74] top n9 unitcap
xc9[73] top n9 unitcap
xc9[72] top n9 unitcap
xc9[71] top n9 unitcap
xc9[70] top n9 unitcap
xc9[69] top n9 unitcap
xc9[68] top n9 unitcap
xc9[67] top n9 unitcap
xc9[66] top n9 unitcap
xc9[65] top n9 unitcap
xc9[64] top n9 unitcap
xc9[63] top n9 unitcap
xc9[62] top n9 unitcap
xc9[61] top n9 unitcap
xc9[60] top n9 unitcap
xc9[59] top n9 unitcap
xc9[58] top n9 unitcap
xc9[57] top n9 unitcap
xc9[56] top n9 unitcap
xc9[55] top n9 unitcap
xc9[54] top n9 unitcap
xc9[53] top n9 unitcap
xc9[52] top n9 unitcap
xc9[51] top n9 unitcap
xc9[50] top n9 unitcap
xc9[49] top n9 unitcap
xc9[48] top n9 unitcap
xc9[47] top n9 unitcap
xc9[46] top n9 unitcap
xc9[45] top n9 unitcap
xc9[44] top n9 unitcap
xc9[43] top n9 unitcap
xc9[42] top n9 unitcap
xc9[41] top n9 unitcap
xc9[40] top n9 unitcap
xc9[39] top n9 unitcap
xc9[38] top n9 unitcap
xc9[37] top n9 unitcap
xc9[36] top n9 unitcap
xc9[35] top n9 unitcap
xc9[34] top n9 unitcap
xc9[33] top n9 unitcap
xc9[32] top n9 unitcap
xc9[31] top n9 unitcap
xc9[30] top n9 unitcap
xc9[29] top n9 unitcap
xc9[28] top n9 unitcap
xc9[27] top n9 unitcap
xc9[26] top n9 unitcap
xc9[25] top n9 unitcap
xc9[24] top n9 unitcap
xc9[23] top n9 unitcap
xc9[22] top n9 unitcap
xc9[21] top n9 unitcap
xc9[20] top n9 unitcap
xc9[19] top n9 unitcap
xc9[18] top n9 unitcap
xc9[17] top n9 unitcap
xc9[16] top n9 unitcap
xc9[15] top n9 unitcap
xc9[14] top n9 unitcap
xc9[13] top n9 unitcap
xc9[12] top n9 unitcap
xc9[11] top n9 unitcap
xc9[10] top n9 unitcap
xc9[9] top n9 unitcap
xc9[8] top n9 unitcap
xc9[7] top n9 unitcap
xc9[6] top n9 unitcap
xc9[5] top n9 unitcap
xc9[4] top n9 unitcap
xc9[3] top n9 unitcap
xc9[2] top n9 unitcap
xc9[1] top n9 unitcap
xc9[0] top n9 unitcap
.ends


* expanding   symbol:  switches/bootstrapped_sw_hv.sym # of pins=5
** sym_path: /home/oe23ranan/gf_analog/xschem/switches/bootstrapped_sw_hv.sym
** sch_path: /home/oe23ranan/gf_analog/xschem/switches/bootstrapped_sw_hv.sch
.subckt bootstrapped_sw_hv out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
xinv1 vdd en enb vss inv_lvt
XCbs[4] vbsh out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs[3] vbsh out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs[2] vbsh out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs[1] vbsh out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs[0] vbsh out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM3 vdd vss vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 vss enb vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMs out vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 out vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out enb out sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMs2 vss enb vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMs1 vss vdd vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar_10b/unitcap/unitcap.sym # of pins=2
** sym_path: /home/oe23ranan/gf_analog/xschem/sar_10b/unitcap/unitcap.sym
** sch_path: /home/oe23ranan/gf_analog/xschem/sar_10b/unitcap/unitcap.sch
.subckt unitcap cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2.6f m=1
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/gf_analog/xschem/logic/inv_lvt.sym
** sch_path: /home/oe23ranan/gf_analog/xschem/logic/inv_lvt.sch
.subckt inv_lvt vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
