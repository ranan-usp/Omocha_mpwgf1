* NGSPICE file created from dac.ext - technology: gf180mcuD

.subckt XM1_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM4_bs G D w_n319_n356# S
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XMs1_bs G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt bs_cap I1_1_1_R0_BOT I1_1_1_R0_TOP
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.339999u c_length=12.339999u
.ends

.subckt XM3_bs G D w_n319_n356# S
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_bs_inv G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_bs_inv G D w_n319_n356# S
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt bs_inv inv_in inv_out vdd vss
XXM1_bs_inv_0 inv_in inv_out vss vss XM1_bs_inv
XXM2_bs_inv_0 inv_in inv_out vdd vdd XM2_bs_inv
.ends

.subckt XMs_bs G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XMs2_bs G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt bootstrapped_sw vbsh vbsl vg vs vdd en enb bs_in bs_out vss
XXM1_bs_0 vg vbsl vss vss bs_in XM1_bs
XXM4_bs_0 vg vdd vbsh vbsh XM4_bs
XXMs1_bs_0 vdd vs vss vg XMs1_bs
Xbs_cap_0 vbsl vbsh bs_cap
Xbs_cap_1 vbsl vbsh bs_cap
XXM3_bs_0 enb vg vbsh vbsh XM3_bs
Xbs_cap_2 vbsl vbsh bs_cap
Xbs_cap_4 vbsl vbsh bs_cap
Xbs_cap_3 vbsl vbsh bs_cap
Xbs_inv_0 en enb vdd vss bs_inv
XXMs_bs_0 vg bs_out vss bs_in XMs_bs
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 enb vss vss vss vs XMs2_bs
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt inv_renketu inv$1_1/I inv$1_8/I inv$1_7/ZN inv$1_1/ZN inv$1_3/I inv$1_5/I
+ inv$1_7/I inv$1_9/ZN inv$1_9/I inv$1_3/ZN inv$1_6/ZN vdd inv$1_0/ZN inv$1_0/I inv$1_4/ZN
+ inv$1_2/I inv$1_10/I inv$1_4/I inv$1_10/ZN inv$1_8/ZN vss inv$1_6/I inv$1_2/ZN inv$1_5/ZN
Xinv$1_10 vss inv$1_10/ZN inv$1_10/I vdd vdd inv$1_10/VPW vss inv$1
Xinv$1_0 vss inv$1_0/ZN inv$1_0/I vdd vdd inv$1_0/VPW vss inv$1
Xinv$1_1 vss inv$1_1/ZN inv$1_1/I vdd vdd inv$1_1/VPW vss inv$1
Xinv$1_2 vss inv$1_2/ZN inv$1_2/I vdd vdd inv$1_2/VPW vss inv$1
Xinv$1_3 vss inv$1_3/ZN inv$1_3/I vdd vdd inv$1_3/VPW vss inv$1
Xinv$1_4 vss inv$1_4/ZN inv$1_4/I vdd vdd inv$1_4/VPW vss inv$1
Xinv$1_5 vss inv$1_5/ZN inv$1_5/I vdd vdd inv$1_5/VPW vss inv$1
Xinv$1_6 vss inv$1_6/ZN inv$1_6/I vdd vdd inv$1_6/VPW vss inv$1
Xinv$1_7 vss inv$1_7/ZN inv$1_7/I vdd vdd inv$1_7/VPW vss inv$1
Xinv$1_8 vss inv$1_8/ZN inv$1_8/I vdd vdd inv$1_8/VPW vss inv$1
Xinv$1_9 vss inv$1_9/ZN inv$1_9/I vdd vdd inv$1_9/VPW vss inv$1
.ends

.subckt dac vdd vss dac_in dac_out dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9
+ ctl10 sample
Xbootstrapped_sw_0 bootstrapped_sw_0/vbsh bootstrapped_sw_0/vbsl bootstrapped_sw_0/vg
+ bootstrapped_sw_0/vs vdd sample bootstrapped_sw_0/enb dac_in dac_out vss bootstrapped_sw
Xinv_renketu_0 ctl2 ctl7 carray_0/n6 carray_0/n2 ctl1 ctl4 ctl6 carray_0/n8 ctl8 carray_0/n1
+ carray_0/n5 vdd carray_0/ndum dum carray_0/n3 ctl10 ctl9 ctl3 carray_0/n9 carray_0/n7
+ vss ctl5 carray_0/n0 carray_0/n4 inv_renketu
.ends

