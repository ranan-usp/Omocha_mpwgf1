magic
tech gf180mcuD
magscale 1 10
timestamp 1701784929
<< checkpaint >>
rect -3188 -2356 3188 2356
<< pwell >>
rect -1188 -356 1188 356
<< mvnmos >>
rect -924 -100 -784 100
rect -680 -100 -540 100
rect -436 -100 -296 100
rect -192 -100 -52 100
rect 52 -100 192 100
rect 296 -100 436 100
rect 540 -100 680 100
rect 784 -100 924 100
<< mvndiff >>
rect -1012 87 -924 100
rect -1012 -87 -999 87
rect -953 -87 -924 87
rect -1012 -100 -924 -87
rect -784 87 -680 100
rect -784 -87 -755 87
rect -709 -87 -680 87
rect -784 -100 -680 -87
rect -540 87 -436 100
rect -540 -87 -511 87
rect -465 -87 -436 87
rect -540 -100 -436 -87
rect -296 87 -192 100
rect -296 -87 -267 87
rect -221 -87 -192 87
rect -296 -100 -192 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 192 87 296 100
rect 192 -87 221 87
rect 267 -87 296 87
rect 192 -100 296 -87
rect 436 87 540 100
rect 436 -87 465 87
rect 511 -87 540 87
rect 436 -100 540 -87
rect 680 87 784 100
rect 680 -87 709 87
rect 755 -87 784 87
rect 680 -100 784 -87
rect 924 87 1012 100
rect 924 -87 953 87
rect 999 -87 1012 87
rect 924 -100 1012 -87
<< mvndiffc >>
rect -999 -87 -953 87
rect -755 -87 -709 87
rect -511 -87 -465 87
rect -267 -87 -221 87
rect -23 -87 23 87
rect 221 -87 267 87
rect 465 -87 511 87
rect 709 -87 755 87
rect 953 -87 999 87
<< mvpsubdiff >>
rect -1156 252 1156 324
rect -1156 208 -1084 252
rect -1156 -208 -1143 208
rect -1097 -208 -1084 208
rect 1084 208 1156 252
rect -1156 -252 -1084 -208
rect 1084 -208 1097 208
rect 1143 -208 1156 208
rect 1084 -252 1156 -208
rect -1156 -324 1156 -252
<< mvpsubdiffcont >>
rect -1143 -208 -1097 208
rect 1097 -208 1143 208
<< polysilicon >>
rect -924 179 -784 192
rect -924 133 -911 179
rect -797 133 -784 179
rect -924 100 -784 133
rect -680 179 -540 192
rect -680 133 -667 179
rect -553 133 -540 179
rect -680 100 -540 133
rect -436 179 -296 192
rect -436 133 -423 179
rect -309 133 -296 179
rect -436 100 -296 133
rect -192 179 -52 192
rect -192 133 -179 179
rect -65 133 -52 179
rect -192 100 -52 133
rect 52 179 192 192
rect 52 133 65 179
rect 179 133 192 179
rect 52 100 192 133
rect 296 179 436 192
rect 296 133 309 179
rect 423 133 436 179
rect 296 100 436 133
rect 540 179 680 192
rect 540 133 553 179
rect 667 133 680 179
rect 540 100 680 133
rect 784 179 924 192
rect 784 133 797 179
rect 911 133 924 179
rect 784 100 924 133
rect -924 -183 -784 -100
rect -680 -183 -540 -100
rect -436 -183 -296 -100
rect -192 -183 -52 -100
rect 52 -183 192 -100
rect 296 -183 436 -100
rect 540 -183 680 -100
rect 784 -183 924 -100
<< polycontact >>
rect -911 133 -797 179
rect -667 133 -553 179
rect -423 133 -309 179
rect -179 133 -65 179
rect 65 133 179 179
rect 309 133 423 179
rect 553 133 667 179
rect 797 133 911 179
<< metal1 >>
rect -1143 208 -1097 204
rect 1097 208 1143 204
rect -922 133 -911 179
rect -797 133 -786 179
rect -678 133 -667 179
rect -553 133 -542 179
rect -434 133 -423 179
rect -309 133 -298 179
rect -190 133 -179 179
rect -65 133 -54 179
rect 54 133 65 179
rect 179 133 190 179
rect 298 133 309 179
rect 423 133 434 179
rect 542 133 553 179
rect 667 133 678 179
rect 786 133 797 179
rect 911 133 922 179
rect -999 87 -953 83
rect -999 -98 -953 -102
rect -755 87 -709 83
rect -755 -98 -709 -102
rect -511 87 -465 83
rect -511 -98 -465 -102
rect -267 87 -221 83
rect -267 -98 -221 -102
rect -23 87 23 83
rect -23 -98 23 -102
rect 221 87 267 83
rect 221 -98 267 -102
rect 465 87 511 83
rect 465 -98 511 -102
rect 709 87 755 83
rect 709 -98 755 -102
rect 953 87 999 83
rect 953 -98 999 -102
rect -1143 -219 -1097 -223
rect 1097 -219 1143 -223
<< labels >>
flabel metal1 -195 -1 -195 -1 0 FreeSans 240 0 0 0 D
flabel metal1 -170 31 -170 31 0 FreeSans 240 0 0 0 G
flabel metal1 -146 -1 -146 -1 0 FreeSans 240 0 0 0 S
flabel metal1 -122 31 -122 31 0 FreeSans 240 0 0 0 G
flabel metal1 -97 -1 -97 -1 0 FreeSans 240 0 0 0 D
flabel metal1 -73 31 -73 31 0 FreeSans 240 0 0 0 G
flabel metal1 -48 -1 -48 -1 0 FreeSans 240 0 0 0 S
flabel metal1 -24 31 -24 31 0 FreeSans 240 0 0 0 G
flabel metal1 0 -1 0 -1 0 FreeSans 240 0 0 0 D
flabel metal1 24 31 24 31 0 FreeSans 240 0 0 0 G
flabel metal1 48 -1 48 -1 0 FreeSans 240 0 0 0 S
flabel metal1 73 31 73 31 0 FreeSans 240 0 0 0 G
flabel metal1 97 -1 97 -1 0 FreeSans 240 0 0 0 D
flabel metal1 122 31 122 31 0 FreeSans 240 0 0 0 G
flabel metal1 146 -1 146 -1 0 FreeSans 240 0 0 0 S
flabel metal1 170 31 170 31 0 FreeSans 240 0 0 0 G
flabel metal1 195 -1 195 -1 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -1120 -288 1120 288
<< end >>


