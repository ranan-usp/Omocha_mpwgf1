* NGSPICE file created from carray_in.ext - technology: gf180mcuD

.subckt carray_in n1 n2 n3 n4 n5 n6 n7 n8 n9 n0 vss dac_out
C0 n6 n5 29.1995f
C1 n9 n8 87.65668f
C2 n4 dac_out 26.242765f
C3 dac_out n0 1.640173f
C4 n3 n7 0.894213f
C5 n1 n7 0.243006f
C6 n2 n7 0.487626f
C7 n4 n9 3.741774f
C8 n9 n0 0.825206f
C9 n7 n5 3.37237f
C10 n9 dac_out 0.846091p
C11 n8 n3 1.46349f
C12 n1 n8 0.333459f
C13 n8 n2 0.772498f
C14 n8 n5 5.6103f
C15 n6 n7 34.8991f
C16 n4 n3 26.505f
C17 n4 n1 0.145617f
C18 n1 n0 8.401715f
C19 n4 n2 0.215946f
C20 dac_out n3 13.12139f
C21 n1 dac_out 3.280347f
C22 dac_out n2 6.560692f
C23 n4 n5 28.093302f
C24 n6 n8 11.2197f
C25 n9 n3 1.912414f
C26 n9 n1 0.39415f
C27 dac_out n5 52.485596f
C28 n9 n2 0.997758f
C29 n9 n5 7.400846f
C30 n4 n6 0.617028f
C31 n6 dac_out 0.104976p
C32 n8 n7 50.741302f
C33 n1 n3 0.148119f
C34 n3 n2 23.4645f
C35 n9 n6 14.718489f
C36 n1 n2 15.5737f
C37 n3 n5 0.350346f
C38 n1 n5 0.145556f
C39 n2 n5 0.210974f
C40 n4 n7 1.70684f
C41 dac_out n7 0.209952p
C42 n6 n3 0.339322f
C43 n4 n8 2.84594f
C44 n1 n6 0.145088f
C45 n6 n2 0.210444f
C46 n9 n7 29.520088f
C47 n8 dac_out 0.420079p
C48 n0 vss 17.641516f
C49 n1 vss 26.92111f
C50 n4 vss 43.231865f
C51 n5 vss 54.41903f
C52 n2 vss 32.35876f
C53 n3 vss 35.924526f
C54 n9 vss 0.119661p
C55 dac_out vss 0.117131p
C56 n8 vss 91.1161f
C57 n7 vss 83.208f
C58 n6 vss 67.765594f
.ends

