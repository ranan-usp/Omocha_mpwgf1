* NGSPICE file created from saradc.ext - technology: gf180mcuD

.subckt XM2$3$1 a_n36_120# a_n116_n100# w_n460_n310#
X0 w_n460_n310# a_n36_120# a_n116_n100# w_n460_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$3$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt x4 out in vdd vss
XXM2$3$1_0 in out vdd XM2$3$1
XXM1$3$1_0 in vss out XM1$3$1
.ends

.subckt XM2$1$3 a_n36_120# a_n116_n100# w_n278_n310#
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$1$3 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt x2 out in vdd vss
XXM2$1$3_0 in out vdd XM2$1$3
XXM1$1$3_0 in vss out XM1$1$3
.ends

.subckt XM4$5 a_258_n1293# a_258_n1793# a_396_n1607# a_476_n1387#
X0 a_540_n1607# a_476_n1387# a_396_n1607# a_258_n1793# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM3$5 a_n67_n1582# a_n349_n1268# a_n131_n1362# a_n349_n1768#
X0 a_n67_n1582# a_n131_n1362# a_n211_n1582# a_n349_n1768# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2$2$1 a_n36_120# a_n116_n100# w_n460_n310#
X0 w_n460_n310# a_n36_120# a_n116_n100# w_n460_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$2$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt x3 out in vdd vss
XXM2$2$1_0 in out vdd XM2$2$1
XXM1$2$1_0 in vss out XM1$2$1
.ends

.subckt XM1$5 a_n36_20# a_n254_n386# a_n254_114# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2$5 a_n36_120# a_n116_n100# w_n278_n310#
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt x1 out in vdd XM1$5_0/a_n254_114# vss
XXM1$5_0 in vss XM1$5_0/a_n254_114# out XM1$5
XXM2$5_0 in out vdd XM2$5
.ends

.subckt latch Qn Q S R VSUBS
Xx4_0 x4_0/out S Q VSUBS x4
Xx2_0 Qn Q Q VSUBS x2
XXM4$5_0 VSUBS VSUBS Q x3_0/out XM4$5
XXM3$5_0 Qn VSUBS x4_0/out VSUBS XM3$5
Xx3_0 x3_0/out R Q VSUBS x3
Xx1_0 Q Qn Q VSUBS VSUBS x1
.ends

.subckt XM2$6 a_n36_120# a_n116_n100# w_n278_n310#
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$6 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt inv$2 out in vdd vss
XXM2$6_0 in out vdd XM2$6
XXM1$6_0 in vss out XM1$6
.ends

.subckt buffer in out inv$2_1/vdd VSUBS
Xinv$2_0 inv$2_1/in in inv$2_1/vdd VSUBS inv$2
Xinv$2_1 out inv$2_1/in inv$2_1/vdd VSUBS inv$2
.ends

.subckt XM3 a_n3152_1140# a_n3064_1048# w_n3314_932# a_n2964_1140#
X0 a_n2964_1140# a_n3064_1048# a_n3152_1140# w_n3314_932# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM1 a_912_4129# a_995_4229# a_811_3903# a_1507_3903# a_995_4041#
X0 a_995_4229# a_912_4129# a_995_4041# a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs a_1030_4680# a_1030_4868# a_947_4768# a_846_4542#
X0 a_1030_4868# a_947_4768# a_1030_4680# a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668#
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0_m4m5_noshield c_width=8u c_length=8u
.ends

.subckt sw_cap_unit in out
Xcap_mim_2p0fF_8JNR63_0 out in cap_mim_2p0fF_8JNR63
.ends

.subckt sw_cap out in
Xsw_cap_unit_0 in out sw_cap_unit
Xsw_cap_unit_1 in out sw_cap_unit
Xsw_cap_unit_2 in out sw_cap_unit
Xsw_cap_unit_3 in out sw_cap_unit
Xsw_cap_unit_4 in out sw_cap_unit
.ends

.subckt XMs1 a_n2529_n616# a_n2717_n616# a_n2629_n699# a_n2855_n800#
X0 a_n2529_n616# a_n2629_n699# a_n2717_n616# a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM4 a_n2550_442# a_n2362_442# w_n2712_234# a_n2462_359#
X0 a_n2362_442# a_n2462_359# a_n2550_442# w_n2712_234# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM2_inv a_n36_120# a_n116_n100# w_n278_n310#
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1_inv a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt inv out in vdd vss
XXM2_inv_0 in out vdd XM2_inv
XXM1_inv_0 in vss out XM1_inv
.ends

.subckt XM2 a_912_3686# a_811_3460# a_995_3786# a_1507_3460# a_995_3598#
X0 a_995_3786# a_912_3686# a_995_3598# a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs2 a_n3762_561# a_n3988_469# a_n3662_653# a_n3850_653# a_n3988_1165#
X0 a_n3662_653# a_n3762_561# a_n3850_653# a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt bootstrapped_sw vbsl vbsh in vdd vss en enb out vs vg
XXM3_0 vbsh vg XM4_0/w_n2712_234# vdd XM3
XXM1_0 vg vbsl vss vss in XM1
XXMs_0 out in vg vss XMs
Xsw_cap_0 vbsh vbsl sw_cap
XXMs1_0 vs vg vdd vss XMs1
XXM4_0 vg vbsh XM4_0/w_n2712_234# enb XM4
Xinv_0 enb en vdd vss inv
XXM2_0 enb vss vss vss vbsl XM2
XXMs2_0 enb vss vss vs vss XMs2
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt dummy VSS ZN I VDD VNW VPW
X0 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt inv_renketu inv$1_8/I inv$1_1/I inv$1_3/I inv$1_5/I inv$1_7/I inv$1_9/ZN inv$1_6/ZN
+ inv$1_0/ZN inv$1_0/I inv$1_4/ZN inv$1_9/I inv$1_2/I inv$1_10/I inv$1_7/ZN inv$1_1/ZN
+ inv$1_3/ZN inv$1_4/I inv$1_8/ZN inv$1_10/ZN VSUBS inv$1_6/I inv$1_2/ZN inv$1_5/ZN
Xinv$1_10 inv$1_9/VSS inv$1_10/ZN inv$1_10/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_0 inv$1_9/VSS inv$1_0/ZN inv$1_0/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_1 inv$1_9/VSS inv$1_1/ZN inv$1_1/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_2 inv$1_9/VSS inv$1_2/ZN inv$1_2/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_3 inv$1_9/VSS inv$1_3/ZN inv$1_3/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_4 inv$1_9/VSS inv$1_4/ZN inv$1_4/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_5 inv$1_9/VSS inv$1_5/ZN inv$1_5/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_6 inv$1_9/VSS inv$1_6/ZN inv$1_6/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_7 inv$1_9/VSS inv$1_7/ZN inv$1_7/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_8 inv$1_9/VSS inv$1_8/ZN inv$1_8/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_9 inv$1_9/VSS inv$1_9/ZN inv$1_9/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xdummy_0 inv$1_9/VSS dummy_0/ZN dummy_0/I inv$1_9/VDD inv$1_9/VNW VSUBS dummy
Xdummy_1 inv$1_9/VSS dummy_1/ZN dummy_1/I inv$1_9/VDD inv$1_9/VNW VSUBS dummy
.ends

.subckt dacp ctl0 in dum ctl2 ctl1 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 out ndum n1
+ n2 n3 n4 n5 n6 n7 n8 n9 n0 sample bootstrapped_sw_0/vbsh vdd vss
Xbootstrapped_sw_0 bootstrapped_sw_0/vbsl bootstrapped_sw_0/vbsh in vdd vss sample
+ bootstrapped_sw_0/enb out bootstrapped_sw_0/vs bootstrapped_sw_0/vg bootstrapped_sw
Xinv_renketu_0 ctl7 ctl2 ctl1 ctl4 ctl6 n8 n5 ndum dum n3 ctl8 ctl0 ctl9 n6 n2 n1
+ ctl3 n7 n9 vss ctl5 n0 n4 inv_renketu
.ends

.subckt inv$1$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt dummy$1 VSS ZN I VDD VNW VPW
X0 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt inv_renketu$1 inv$1$1_7/I inv$1$1_6/ZN inv$1$1_9/ZN inv$1$1_0/I inv$1$1_10/I
+ inv$1$1_0/ZN inv$1$1_4/I inv$1$1_6/I inv$1$1_8/ZN inv$1$1_5/ZN inv$1$1_8/I inv$1$1_2/I
+ inv$1$1_2/ZN inv$1$1_1/I inv$1$1_9/I inv$1$1_7/ZN inv$1$1_3/ZN inv$1$1_3/I inv$1$1_4/ZN
+ inv$1$1_1/ZN inv$1$1_5/I inv$1$1_10/ZN VSUBS
Xinv$1$1_0 inv$1$1_9/VSS inv$1$1_0/ZN inv$1$1_0/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_1 inv$1$1_9/VSS inv$1$1_1/ZN inv$1$1_1/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_2 inv$1$1_9/VSS inv$1$1_2/ZN inv$1$1_2/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_3 inv$1$1_9/VSS inv$1$1_3/ZN inv$1$1_3/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_4 inv$1$1_9/VSS inv$1$1_4/ZN inv$1$1_4/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_5 inv$1$1_9/VSS inv$1$1_5/ZN inv$1$1_5/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_6 inv$1$1_9/VSS inv$1$1_6/ZN inv$1$1_6/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_7 inv$1$1_9/VSS inv$1$1_7/ZN inv$1$1_7/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_8 inv$1$1_9/VSS inv$1$1_8/ZN inv$1$1_8/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xdummy$1_0 inv$1$1_9/VSS dummy$1_0/ZN dummy$1_0/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ dummy$1
Xinv$1$1_9 inv$1$1_9/VSS inv$1$1_9/ZN inv$1$1_9/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xdummy$1_1 inv$1$1_9/VSS dummy$1_1/ZN dummy$1_1/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ dummy$1
Xinv$1$1_10 inv$1$1_9/VSS inv$1$1_10/ZN inv$1$1_10/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
.ends

.subckt XMs$1 a_1030_4680# a_1030_4868# a_947_4768# a_846_4542#
X0 a_1030_4868# a_947_4768# a_1030_4680# a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM3$4 a_n3152_1140# a_n3064_1048# w_n3314_932# a_n2964_1140#
X0 a_n2964_1140# a_n3064_1048# a_n3152_1140# w_n3314_932# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM2_inv$1 a_n36_120# a_n116_n100# w_n278_n310#
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1_inv$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt inv$3 out in vdd vss
XXM2_inv$1_0 in out vdd XM2_inv$1
XXM1_inv$1_0 in vss out XM1_inv$1
.ends

.subckt XMs2$1 a_n3762_561# a_n3988_469# a_n3662_653# a_n3850_653# a_n3988_1165#
X0 a_n3662_653# a_n3762_561# a_n3850_653# a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM2$4 a_912_3686# a_811_3460# a_995_3786# a_1507_3460# a_995_3598#
X0 a_995_3786# a_912_3686# a_995_3598# a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt cap_mim_2p0fF_8JNR63$1 m4_n3440_n548# m4_n3800_n668#
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0_m4m5_noshield c_width=8u c_length=8u
.ends

.subckt sw_cap_unit$1 in out
Xcap_mim_2p0fF_8JNR63_0 out in cap_mim_2p0fF_8JNR63$1
.ends

.subckt sw_cap$1 out in
Xsw_cap_unit$1_0 in out sw_cap_unit$1
Xsw_cap_unit$1_1 in out sw_cap_unit$1
Xsw_cap_unit$1_2 in out sw_cap_unit$1
Xsw_cap_unit$1_3 in out sw_cap_unit$1
Xsw_cap_unit$1_4 in out sw_cap_unit$1
.ends

.subckt XMs1$1 a_n2529_n616# a_n2717_n616# a_n2629_n699# a_n2855_n800#
X0 a_n2529_n616# a_n2629_n699# a_n2717_n616# a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM1$4 a_912_4129# a_995_4229# a_811_3903# a_1507_3903# a_995_4041#
X0 a_995_4229# a_912_4129# a_995_4041# a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM4$4 a_n2550_442# a_n2362_442# w_n2712_234# a_n2462_359#
X0 a_n2362_442# a_n2462_359# a_n2550_442# w_n2712_234# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt bootstrapped_sw$1 vbsl vbsh in vdd vss en enb out vs vg
XXMs$1_0 out in vg vss XMs$1
XXM3$4_0 vbsh vg XM4$4_0/w_n2712_234# vdd XM3$4
Xinv$3_0 enb en vdd vss inv$3
XXMs2$1_0 enb vss vss vs vss XMs2$1
XXM2$4_0 enb vss vss vss vbsl XM2$4
Xsw_cap$1_0 vbsh vbsl sw_cap$1
XXMs1$1_0 vs vg vdd vss XMs1$1
XXM1$4_0 vg vbsl vss vss in XM1$4
XXM4$4_0 vg vbsh XM4$4_0/w_n2712_234# enb XM4$4
.ends

.subckt dacn in dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl0 out ndum n1
+ n2 n3 n4 n5 n6 n7 n8 n9 n0 sample vdd bootstrapped_sw$1_0/vbsh vss
Xinv_renketu$1_0 ctl6 n5 n8 dum ctl9 ndum ctl3 ctl5 n7 n4 ctl7 ctl0 n0 ctl2 ctl8 n6
+ n1 ctl1 n3 n2 ctl4 n9 vss inv_renketu$1
Xbootstrapped_sw$1_0 bootstrapped_sw$1_0/vbsl bootstrapped_sw$1_0/vbsh in vdd vss
+ sample bootstrapped_sw$1_0/enb out bootstrapped_sw$1_0/vs bootstrapped_sw$1_0/vg
+ bootstrapped_sw$1
.ends

.subckt XMinn a_719_n1284# a_937_n880# a_857_n1100# a_719_n788# a_1001_n1100#
X0 a_1001_n1100# a_937_n880# a_857_n1100# a_719_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$3 a_n1416_1000# a_n1336_908# a_n1272_1000# w_n1578_790#
X0 a_n1272_1000# a_n1336_908# a_n1416_1000# w_n1578_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM3$2 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2$2 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM0$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$2 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM4$2 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt trim_switch$1 m1_n149_n1117# m1_n1378_n1819# m1_711_n1117# m1_n2738_n1819#
+ m1_n447_n1117# m1_n2669_n1117# XM1$2_0/a_n202_583# XM0$1_0/a_n346_583# m1_n1309_n1117#
+ m1_802_n1819# VSUBS
XXM3$2_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$2
XXM2$2_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$2
XXM0$1_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0$1_0/a_n346_583# XM0$1
XXM1$2_0 VSUBS XM1$2_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$2
XXM4$2_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$2
.ends

.subckt trim drain d_4 d_1 d_0 d_2 d_3 n4 n1 n0 n2 n3 VSUBS
Xtrim_switch$1_0 d_1 n2 d_4 n3 d_0 d_3 n1 n0 d_2 n4 VSUBS trim_switch$1
.ends

.subckt XMl4 a_44_908# a_108_1000# a_n36_1000# w_n198_790#
X0 a_108_1000# a_44_908# a_n36_1000# w_n198_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM4$3 a_1264_908# a_1328_1000# w_1022_790# a_1184_1000#
X0 a_1328_1000# a_1264_908# a_1184_1000# w_1022_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XMl2 a_33_n1100# a_n111_n1100# a_n31_n880# a_n249_n1284#
X0 a_33_n1100# a_n31_n880# a_n111_n1100# a_n249_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM3$3 a_n71_n882# a_73_n882# a_9_n662# w_n509_n1092#
X0 a_73_n882# a_9_n662# a_n71_n882# w_n509_n1092# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XMdiff a_721_n1097# a_817_n1189# a_439_n1281# a_657_n1189# a_577_n1097# a_881_n1097#
X0 a_721_n1097# a_657_n1189# a_577_n1097# a_439_n1281# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_881_n1097# a_817_n1189# a_721_n1097# a_439_n1281# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt XMl3 a_n116_908# w_n634_790# a_n196_1000# a_n52_1000#
X0 a_n52_1000# a_n116_908# a_n196_1000# w_n634_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM4$1 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt XM2$1$1 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1$1$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM3$1 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM0 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt trim_switch m1_n149_n1117# XM0_0/a_n346_583# m1_711_n1117# m1_n447_n1117#
+ m1_n2669_n1117# m1_n1378_n1819# m1_802_n1819# m1_n1309_n1117# XM1$1$1_0/a_n202_583#
+ m1_n2738_n1819# VSUBS
XXM4$1_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$1
XXM2$1$1_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$1$1
XXM1$1$1_0 VSUBS XM1$1$1_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$1$1
XXM3$1_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$1
XXM0_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0_0/a_n346_583# XM0
.ends

.subckt trimb d_4 d_1 d_0 d_2 d_3 n4 n1 n0 n2 n3 drain VSUBS
Xtrim_switch_0 d_1 n0 d_4 d_0 d_3 n2 n4 d_2 n1 n3 VSUBS trim_switch
.ends

.subckt XMl1 a_1362_n1100# a_1442_n880# a_1506_n1100# a_1224_n1284#
X0 a_1506_n1100# a_1442_n880# a_1362_n1100# a_1224_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2$3 a_69_n911# w_n237_n1121# a_5_n691# a_n75_n911#
X0 a_69_n911# a_5_n691# a_n75_n911# w_n237_n1121# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XMinp a_251_n1284# a_389_n1100# a_251_n788# a_469_n880# a_533_n1100#
X0 a_533_n1100# a_469_n880# a_389_n1100# a_251_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt comparator vdd outp outn vp vn trim3 trimb0 trimb3 diff ip in clkc trim4 trim2
+ trim1 trim0 trimb4 trimb2 vss trimb1
XXMinn_0 vss vn in vss diff XMinn
XXM1$3_0 in clkc vdd vdd XM1$3
Xtrim_0 in trim4 trim1 trim0 trim2 trim3 trim_0/n4 trim_0/n1 trim_0/n0 trim_0/n2 trim_0/n3
+ vss trim
XXMl4_0 outn outp vdd vdd XMl4
XXM4$3_0 clkc ip vdd vdd XM4$3
XXMl2_0 outp ip outn vss XMl2
XXM3$3_0 outp vdd clkc vdd XM3$3
XXMdiff_0 diff clkc vss clkc vss vss XMdiff
XXMl3_0 outp vdd outn vdd XMl3
Xtrimb_0 trimb4 trimb1 trimb0 trimb2 trimb3 trimb_0/n4 trimb_0/n1 trimb_0/n0 trimb_0/n2
+ trimb_0/n3 ip vss trimb
XXMl1_0 outn outp in vss XMl1
XXM2$3_0 outn vdd clkc vdd XM2$3
XXMinp_0 vss diff vss vp ip XMinp
.ends

.subckt cap_mim_2p0fF_RCWXT2$1 m4_n3120_n3000# m4_n3240_n3120#
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30_flip cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ cap_mim_2p0fF_RCWXT2$1
.ends

.subckt cap_mim_2p0fF_RCWXT2 m4_n3120_n3000# m4_n3240_n3120#
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ cap_mim_2p0fF_RCWXT2
.ends

.subckt mim_cap1 m5_n86730_51500# m5_n11730_51500# m5_n33870_51500# m5_86130_51500#
+ m5_14520_n66196# m5_n18870_51500# m5_44520_n66196# m5_n30480_n66196# m5_74520_n66196#
+ m5_33270_51500# m5_11130_51500# m5_n480_n66196# m5_n60480_n66196# m5_18270_51500#
+ m5_n90480_n66196# m5_104520_n66196# m5_n41730_51500# m5_n63870_51500# m5_n26730_51500#
+ m5_n48870_51500# m5_n3870_51500# m5_n105480_n66196# m5_n101730_51500# m5_63270_51500#
+ m5_n108870_51500# m5_48270_51500# m5_41130_51500# m5_29520_n66196# m5_26130_51500#
+ m5_n15480_n66196# m5_n93870_51500# m5_59520_n66196# m5_3270_51500# m5_n71730_51500#
+ m5_n78870_51500# m5_n45480_n66196# m5_n56730_51500# m5_89520_n66196# m5_n75480_n66196#
+ m5_93270_51500# m5_71130_51500# m5_101130_51500# m5_78270_51500# m5_56130_51500#
+ m5_108270_51500#
Xmim_cap_30_30_flip_233 m5_89520_n66196# mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_222 m5_14520_n66196# mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_200 m5_44520_n66196# mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_211 m5_n480_n66196# mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_68 m5_n45480_n66196# mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_57 m5_n15480_n66196# mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_79 m5_n75480_n66196# mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_13 m5_44520_n66196# mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_24 m5_44520_n66196# mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_46 m5_89520_n66196# mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_35 m5_29520_n66196# mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_213 m5_29520_n66196# m5_26130_51500# mim_cap_30_30
Xmim_cap_30_30_224 m5_104520_n66196# mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_202 m5_29520_n66196# mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_235 m5_59520_n66196# mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_212 m5_44520_n66196# m5_48270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_234 m5_74520_n66196# mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_223 m5_n480_n66196# mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_201 m5_29520_n66196# mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_58 m5_n30480_n66196# mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_69 m5_n30480_n66196# mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_14 m5_29520_n66196# mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_25 m5_29520_n66196# mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_47 m5_74520_n66196# mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_36 m5_104520_n66196# mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_214 m5_14520_n66196# m5_11130_51500# mim_cap_30_30
Xmim_cap_30_30_225 m5_89520_n66196# mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_203 m5_14520_n66196# mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_236 m5_59520_n66196# mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_224 m5_104520_n66196# m5_108270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_213 m5_29520_n66196# m5_33270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_235 m5_59520_n66196# mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_202 m5_14520_n66196# mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_59 m5_n45480_n66196# mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_15 m5_14520_n66196# mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_48 m5_59520_n66196# mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_26 m5_14520_n66196# mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_37 m5_104520_n66196# mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_226 m5_74520_n66196# mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_204 m5_14520_n66196# mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_237 m5_59520_n66196# mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_215 m5_44520_n66196# mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_225 m5_89520_n66196# m5_93270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_214 m5_14520_n66196# m5_18270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_236 m5_104520_n66196# mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_203 m5_n480_n66196# mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_16 m5_29520_n66196# mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_49 m5_59520_n66196# mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_38 m5_89520_n66196# mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_27 m5_14520_n66196# mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_227 m5_89520_n66196# mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_238 m5_59520_n66196# mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_205 m5_44520_n66196# mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_216 m5_29520_n66196# mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_226 m5_74520_n66196# m5_78270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_215 m5_n480_n66196# m5_3270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_237 m5_89520_n66196# mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_204 m5_44520_n66196# mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_17 m5_44520_n66196# mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_28 m5_44520_n66196# mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_39 m5_74520_n66196# mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_228 m5_104520_n66196# mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_217 m5_44520_n66196# mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_239 m5_59520_n66196# mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_206 m5_29520_n66196# mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_227 m5_59520_n66196# m5_63270_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_216 m5_44520_n66196# mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_238 m5_74520_n66196# mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_205 m5_29520_n66196# mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_18 m5_29520_n66196# mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_29 m5_29520_n66196# mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_229 m5_89520_n66196# mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_218 m5_29520_n66196# mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_207 m5_14520_n66196# mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_228 m5_104520_n66196# mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_217 m5_29520_n66196# mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_206 m5_14520_n66196# mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_239 m5_59520_n66196# mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_19 m5_14520_n66196# mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_219 m5_44520_n66196# mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_208 m5_29520_n66196# mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_229 m5_89520_n66196# mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_218 m5_14520_n66196# mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_207 m5_n480_n66196# mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_209 m5_14520_n66196# mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_219 m5_n480_n66196# mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_208 m5_44520_n66196# mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_190 m5_74520_n66196# mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_209 m5_29520_n66196# mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_90 m5_n90480_n66196# mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_180 m5_n30480_n66196# mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_191 m5_74520_n66196# mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_80 m5_n75480_n66196# mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_91 m5_n90480_n66196# mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_190 m5_74520_n66196# mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_170 m5_n45480_n66196# m5_n48870_51500# mim_cap_30_30
Xmim_cap_30_30_181 m5_n45480_n66196# mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_192 m5_104520_n66196# mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_81 m5_n90480_n66196# mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_70 m5_n15480_n66196# mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_92 m5_n75480_n66196# mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_0 m5_59520_n66196# mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_191 m5_59520_n66196# mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_180 m5_104520_n66196# mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_0 m5_89520_n66196# mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_160 m5_n105480_n66196# mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_193 m5_89520_n66196# mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_182 m5_n45480_n66196# mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_171 m5_n480_n66196# mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_60 m5_59520_n66196# mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_82 m5_n75480_n66196# mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_71 m5_n30480_n66196# mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_93 m5_n90480_n66196# mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_1 m5_104520_n66196# mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_170 m5_n60480_n66196# mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_192 m5_44520_n66196# mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_181 m5_89520_n66196# mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_1 m5_74520_n66196# mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_183 m5_n480_n66196# m5_n3870_51500# mim_cap_30_30
Xmim_cap_30_30_172 m5_n480_n66196# mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_150 m5_n60480_n66196# mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_194 m5_74520_n66196# mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_161 m5_n90480_n66196# mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_83 m5_n90480_n66196# mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_72 m5_n45480_n66196# mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_94 m5_n75480_n66196# mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_50 m5_74520_n66196# mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_61 m5_104520_n66196# mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_2 m5_89520_n66196# mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_160 m5_n30480_n66196# mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_193 m5_29520_n66196# mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_182 m5_74520_n66196# mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_171 m5_n60480_n66196# mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_2 m5_104520_n66196# mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_173 m5_n15480_n66196# mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_162 m5_n60480_n66196# mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_184 m5_89520_n66196# mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_195 m5_104520_n66196# mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_140 m5_n105480_n66196# mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_151 m5_n105480_n66196# mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_73 m5_n15480_n66196# mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_84 m5_n75480_n66196# mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_95 m5_n90480_n66196# mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_51 m5_59520_n66196# mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_40 m5_44520_n66196# mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_62 m5_89520_n66196# mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_3 m5_104520_n66196# mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_161 m5_n45480_n66196# mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_172 m5_n60480_n66196# mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_194 m5_14520_n66196# mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_183 m5_59520_n66196# mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_150 m5_n105480_n66196# mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_3 m5_89520_n66196# mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_174 m5_n30480_n66196# mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_152 m5_n75480_n66196# mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_141 m5_n105480_n66196# mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_196 m5_44520_n66196# mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_130 m5_n15480_n66196# mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_185 m5_104520_n66196# mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_163 m5_n105480_n66196# mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_30 m5_29520_n66196# mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_74 m5_n30480_n66196# mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_85 m5_n90480_n66196# mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_52 m5_104520_n66196# mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_96 m5_n105480_n66196# mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_41 m5_29520_n66196# mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_63 m5_74520_n66196# mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_4 m5_89520_n66196# mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_151 m5_n105480_n66196# mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_162 m5_n15480_n66196# mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_140 m5_n75480_n66196# mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_173 m5_n60480_n66196# mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_184 m5_104520_n66196# mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_195 m5_n480_n66196# mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_4 m5_74520_n66196# mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_131 m5_n30480_n66196# mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_120 m5_n30480_n66196# mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_153 m5_n90480_n66196# mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_186 m5_89520_n66196# mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_142 m5_n60480_n66196# mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_197 m5_44520_n66196# mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_164 m5_n60480_n66196# mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_175 m5_n15480_n66196# mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_31 m5_14520_n66196# mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_75 m5_n45480_n66196# mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_20 m5_29520_n66196# mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_64 m5_n15480_n66196# mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_86 m5_n75480_n66196# mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_42 m5_44520_n66196# mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_53 m5_89520_n66196# mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_97 m5_n105480_n66196# mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_5 m5_74520_n66196# mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_152 m5_n105480_n66196# m5_n101730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_163 m5_n30480_n66196# mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_141 m5_n90480_n66196# mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_174 m5_n60480_n66196# mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_130 m5_n45480_n66196# mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_196 m5_44520_n66196# mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_185 m5_89520_n66196# mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_5 m5_104520_n66196# mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_154 m5_n60480_n66196# m5_n63870_51500# mim_cap_30_30
Xmim_cap_30_30_176 m5_n45480_n66196# mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_165 m5_n60480_n66196# mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_110 m5_n480_n66196# mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_132 m5_n480_n66196# mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_121 m5_n45480_n66196# mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_143 m5_n75480_n66196# mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_198 m5_29520_n66196# mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_187 m5_104520_n66196# mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_76 m5_n105480_n66196# mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_21 m5_14520_n66196# mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_65 m5_n30480_n66196# mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_10 m5_104520_n66196# mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_32 m5_44520_n66196# mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_43 m5_29520_n66196# mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_54 m5_74520_n66196# mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_87 m5_n90480_n66196# mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_98 m5_n105480_n66196# mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_6 m5_59520_n66196# mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_153 m5_n75480_n66196# mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_164 m5_n45480_n66196# mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_175 m5_n60480_n66196# mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_131 m5_n15480_n66196# mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_142 m5_n75480_n66196# mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_120 m5_n15480_n66196# mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_197 m5_29520_n66196# mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_186 m5_74520_n66196# mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_6 m5_89520_n66196# mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_155 m5_n75480_n66196# m5_n78870_51500# mim_cap_30_30
Xmim_cap_30_30_166 m5_n75480_n66196# mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_111 m5_n15480_n66196# mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_100 m5_n105480_n66196# mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_133 m5_n15480_n66196# mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_144 m5_n90480_n66196# mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_122 m5_n30480_n66196# mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_199 m5_14520_n66196# mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_188 m5_89520_n66196# mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_177 m5_n30480_n66196# mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_77 m5_n105480_n66196# mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_22 m5_n480_n66196# mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_66 m5_n45480_n66196# mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_11 m5_89520_n66196# mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_99 m5_n105480_n66196# mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_33 m5_29520_n66196# mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_44 m5_14520_n66196# mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_55 m5_59520_n66196# mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_88 m5_n75480_n66196# mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_7 m5_74520_n66196# mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_110 m5_n30480_n66196# mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_121 m5_n30480_n66196# mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_154 m5_n90480_n66196# mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_176 m5_104520_n66196# mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_143 m5_n90480_n66196# mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_198 m5_14520_n66196# mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_187 m5_59520_n66196# mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_132 m5_n105480_n66196# mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_165 m5_n15480_n66196# mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_7 m5_104520_n66196# mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_156 m5_n90480_n66196# m5_n93870_51500# mim_cap_30_30
Xmim_cap_30_30_167 m5_n90480_n66196# mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_178 m5_n480_n66196# mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_101 m5_n105480_n66196# mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_112 m5_n30480_n66196# mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_145 m5_n75480_n66196# mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_123 m5_n45480_n66196# mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_189 m5_74520_n66196# mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_134 m5_n480_n66196# mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_23 m5_14520_n66196# mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_67 m5_n15480_n66196# mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_78 m5_n105480_n66196# mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_12 m5_74520_n66196# mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_34 m5_14520_n66196# mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_56 m5_104520_n66196# mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_45 m5_n480_n66196# mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_89 m5_n75480_n66196# mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_8 m5_59520_n66196# mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_100 m5_n45480_n66196# mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_111 m5_n15480_n66196# mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_177 m5_89520_n66196# mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_188 m5_104520_n66196# mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_133 m5_n105480_n66196# mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_122 m5_n45480_n66196# mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_199 m5_n480_n66196# mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_144 m5_n90480_n66196# mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_155 m5_n75480_n66196# mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_166 m5_n30480_n66196# mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_8 m5_89520_n66196# mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_168 m5_n15480_n66196# m5_n18870_51500# mim_cap_30_30
Xmim_cap_30_30_157 m5_n105480_n66196# m5_n108870_51500# mim_cap_30_30
Xmim_cap_30_30_179 m5_n15480_n66196# mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_102 m5_n105480_n66196# mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_113 m5_n45480_n66196# mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_135 m5_n45480_n66196# mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_146 m5_n60480_n66196# mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_124 m5_n15480_n66196# mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_68 m5_n30480_n66196# mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_79 m5_n105480_n66196# mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_24 m5_44520_n66196# mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_13 m5_59520_n66196# mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_35 m5_n480_n66196# mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_57 m5_89520_n66196# mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_46 m5_14520_n66196# mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_9 m5_104520_n66196# mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_156 m5_n15480_n66196# m5_n11730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_145 m5_n75480_n66196# mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_101 m5_n15480_n66196# mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_112 m5_n60480_n66196# mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_123 m5_n30480_n66196# mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_178 m5_74520_n66196# mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_134 m5_n105480_n66196# mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_189 m5_89520_n66196# mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_167 m5_n45480_n66196# mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_9 m5_74520_n66196# mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_103 m5_n105480_n66196# mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_114 m5_n480_n66196# mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_136 m5_n105480_n66196# mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_147 m5_n75480_n66196# mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_125 m5_n30480_n66196# mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_169 m5_n30480_n66196# m5_n33870_51500# mim_cap_30_30
Xmim_cap_30_30_158 m5_n105480_n66196# mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_14 m5_89520_n66196# mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_69 m5_n45480_n66196# mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_25 m5_29520_n66196# mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_58 m5_74520_n66196# mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_36 m5_44520_n66196# mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_47 m5_n480_n66196# mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_157 m5_n30480_n66196# m5_n26730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_168 m5_n60480_n66196# m5_n56730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_146 m5_n90480_n66196# mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_113 m5_n60480_n66196# mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_102 m5_n30480_n66196# mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_135 m5_n105480_n66196# mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_124 m5_n45480_n66196# mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_179 m5_59520_n66196# mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_104 m5_n30480_n66196# mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_115 m5_n15480_n66196# mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_137 m5_n60480_n66196# mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_148 m5_n90480_n66196# mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_126 m5_n45480_n66196# mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_159 m5_n75480_n66196# mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_15 m5_74520_n66196# mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_26 m5_14520_n66196# mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_59 m5_59520_n66196# mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_37 m5_29520_n66196# mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_48 m5_104520_n66196# mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_158 m5_n45480_n66196# m5_n41730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_147 m5_n75480_n66196# m5_n71730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_169 m5_n60480_n66196# mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_114 m5_n60480_n66196# mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_103 m5_n45480_n66196# mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_136 m5_n75480_n66196# mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_125 m5_n15480_n66196# mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_105 m5_n45480_n66196# mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_116 m5_n30480_n66196# mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_149 m5_n90480_n66196# mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_138 m5_n75480_n66196# mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_127 m5_n480_n66196# mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_16 m5_n480_n66196# mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_27 m5_n480_n66196# mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_38 m5_14520_n66196# mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_49 m5_89520_n66196# mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_115 m5_n60480_n66196# mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_104 m5_n15480_n66196# mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_137 m5_n90480_n66196# mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_126 m5_n30480_n66196# mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_148 m5_n90480_n66196# m5_n86730_51500# mim_cap_30_30_flip
Xmim_cap_30_30_flip_159 m5_n15480_n66196# mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_117 m5_n45480_n66196# mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_106 m5_n480_n66196# mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_139 m5_n90480_n66196# mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_128 m5_n15480_n66196# mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_17 m5_44520_n66196# mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_28 m5_n480_n66196# mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_39 m5_n480_n66196# mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_149 m5_n105480_n66196# mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_116 m5_n60480_n66196# mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_105 m5_n30480_n66196# mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_138 m5_n75480_n66196# mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_127 m5_n45480_n66196# mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_118 m5_n480_n66196# mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_107 m5_n15480_n66196# mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_129 m5_n480_n66196# mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_90 m5_n60480_n66196# mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_29 m5_44520_n66196# mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_18 m5_29520_n66196# mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_117 m5_n60480_n66196# mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_106 m5_n45480_n66196# mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_139 m5_n90480_n66196# mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_128 m5_n15480_n66196# mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_119 m5_n15480_n66196# mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_108 m5_n30480_n66196# mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_80 m5_n90480_n66196# mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_91 m5_n75480_n66196# mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_19 m5_44520_n66196# mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_118 m5_n60480_n66196# mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_107 m5_n15480_n66196# mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_129 m5_n30480_n66196# mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_109 m5_n45480_n66196# mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_70 m5_n45480_n66196# mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_81 m5_n60480_n66196# mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_92 m5_n90480_n66196# mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_119 m5_n60480_n66196# mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_108 m5_n30480_n66196# mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_82 m5_n75480_n66196# mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_60 m5_n30480_n66196# mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_71 m5_n15480_n66196# mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_93 m5_n60480_n66196# mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_109 m5_n45480_n66196# mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_50 m5_59520_n66196# mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_83 m5_n90480_n66196# mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_72 m5_n60480_n66196# mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_61 m5_n45480_n66196# mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_94 m5_n75480_n66196# mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_73 m5_n75480_n66196# mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_84 m5_n105480_n66196# mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_62 m5_n480_n66196# mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_95 m5_n90480_n66196# mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_51 m5_59520_n66196# mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_40 m5_89520_n66196# mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_74 m5_n90480_n66196# mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_52 m5_59520_n66196# mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_85 m5_n105480_n66196# mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_63 m5_n480_n66196# mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_96 m5_n75480_n66196# mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_30 m5_44520_n66196# mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_41 m5_74520_n66196# mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_230 m5_74520_n66196# mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_75 m5_n60480_n66196# mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_20 m5_29520_n66196# mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_64 m5_n15480_n66196# mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_86 m5_n105480_n66196# mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_53 m5_59520_n66196# mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_31 m5_29520_n66196# mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_42 m5_104520_n66196# mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_97 m5_n60480_n66196# mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_220 m5_104520_n66196# m5_101130_51500# mim_cap_30_30
Xmim_cap_30_30_231 m5_74520_n66196# mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_230 m5_74520_n66196# mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_65 m5_n480_n66196# mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_76 m5_n75480_n66196# mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_10 m5_74520_n66196# mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_54 m5_59520_n66196# mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_21 m5_14520_n66196# mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_87 m5_n105480_n66196# mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_32 m5_14520_n66196# mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_43 m5_89520_n66196# mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_98 m5_n75480_n66196# mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_221 m5_89520_n66196# m5_86130_51500# mim_cap_30_30
Xmim_cap_30_30_232 m5_59520_n66196# m5_56130_51500# mim_cap_30_30
Xmim_cap_30_30_210 m5_14520_n66196# mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_231 m5_59520_n66196# mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_220 m5_44520_n66196# mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_66 m5_n15480_n66196# mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_77 m5_n90480_n66196# mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_11 m5_104520_n66196# mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_22 m5_14520_n66196# mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_88 m5_n90480_n66196# mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_44 m5_74520_n66196# mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_99 m5_n90480_n66196# mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_33 m5_14520_n66196# mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_55 m5_59520_n66196# mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_222 m5_74520_n66196# m5_71130_51500# mim_cap_30_30
Xmim_cap_30_30_233 m5_59520_n66196# mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_200 m5_29520_n66196# mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_211 m5_14520_n66196# mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_flip_232 m5_104520_n66196# mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_221 m5_29520_n66196# mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_flip_210 m5_14520_n66196# mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30_flip
Xmim_cap_30_30_67 m5_n30480_n66196# mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_12 m5_44520_n66196# mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_23 m5_44520_n66196# mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_56 m5_n480_n66196# mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_78 m5_n60480_n66196# mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_89 m5_n60480_n66196# mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_45 m5_104520_n66196# mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_34 m5_44520_n66196# mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_212 m5_44520_n66196# m5_41130_51500# mim_cap_30_30
Xmim_cap_30_30_234 m5_59520_n66196# mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_223 m5_104520_n66196# mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
Xmim_cap_30_30_201 m5_44520_n66196# mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ mim_cap_30_30
.ends

.subckt cap_mim_2p0fF_DMYL6H m4_n114303_n17580# m4_n114183_n17460#
X0 m4_n114183_n17460# m4_n114303_n17580# cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
.ends

.subckt mim_cap_100_100 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ cap_mim_2p0fF_DMYL6H
.ends

.subckt cap_mim_2p0fF_RCWXT2$2 m4_n3148_n3000# m4_n3268_n3120#
X0 m4_n3148_n3000# m4_n3268_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30$1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120#
+ cap_mim_2p0fF_RCWXT2$2
.ends

.subckt cap_mim_2p0fF_DMYL6H$1 m4_93823_n2660# m4_93943_n2540#
X0 m4_93943_n2540# m4_93823_n2660# cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
.ends

.subckt mim_cap_100_100$1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ cap_mim_2p0fF_DMYL6H$1
.ends

.subckt mim_cap2 vdd vss
Xmim_cap_100_100_1 vss vdd mim_cap_100_100
Xmim_cap_100_100_0 vss vdd mim_cap_100_100
Xmim_cap_100_100_2 vss vdd mim_cap_100_100
Xmim_cap_100_100_3 vss vdd mim_cap_100_100
Xmim_cap_30_30$1_20 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_0 vss vdd mim_cap_30_30$1
Xmim_cap_100_100_4 vss vdd mim_cap_100_100
Xmim_cap_30_30$1_22 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_21 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_11 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_10 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_1 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_23 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_12 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_2 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_24 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_13 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_3 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_14 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_4 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_15 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_6 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_5 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_16 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_7 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_17 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_8 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_18 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_9 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_19 vss vdd mim_cap_30_30$1
Xmim_cap_100_100$1_0 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_1 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_2 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_4 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_3 vss vdd mim_cap_100_100$1
.ends

.subckt mim_cap_boss vss vdd
Xmim_cap1_0 vdd vdd vdd vdd vss vdd vss vss vss vdd vdd vss vss vdd vss vss vdd vdd
+ vdd vdd vdd vss vdd vdd vdd vdd vdd vss vdd vss vdd vss vdd vdd vdd vss vdd vss
+ vss vdd vdd vdd vdd vdd vdd mim_cap1
Xmim_cap2_0 vdd vss mim_cap2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VNW VPW
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VPW nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VNW VPW
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VNW VPW
X0 Z a_36_160# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VPW nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VNW VPW
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VNW VPW
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VNW VPW
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VPW nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VPW nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VPW nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VNW VPW
X0 VSS B ZN VPW nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VPW nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VNW VPW
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VPW nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VNW VPW
X0 a_1229_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VPW nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VNW VPW
X0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VPW nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VPW nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VPW nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VPW nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VPW nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VPW nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VPW nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VPW nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctln[8]
+ ctln[9] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8]
+ ctlp[9] cal clk clkc comp en result[0] result[1] result[2] result[3] result[4] result[5]
+ result[6] result[7] result[8] result[9] rstn sample trim[0] trim[1] trim[2] trim[3]
+ trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] valid vdd vss
XFILLER_0_17_200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_432_ _021_ mask\[3\] net63 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_294_ vdd vss _008_ _104_ _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput7 ctln[0] net7 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_431_ _020_ mask\[2\] net53 vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_293_ net31 vdd vss _106_ mask\[4\] _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_362_ vdd vss trim_mask\[1\] _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_276_ vss _093_ _092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_345_ vss _144_ _132_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_259_ _078_ vdd vss _080_ _073_ _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_430_ _019_ mask\[1\] net63 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_292_ vss _105_ _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_361_ vdd vss _154_ _086_ _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__191__I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_327_ _131_ vdd vss _016_ _127_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_189_ vdd vss _043_ net27 mask\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_258_ vss _079_ _078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput33 result[6] net33 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput22 ctlp[5] net22 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__292__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__301__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 ctlp[6] net23 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_273_ vss _090_ state\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout80 vss net80 net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_78 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_325_ vdd vss _130_ _118_ _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 ctln[6] net13 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput24 ctlp[7] net24 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_324_ vdd vss _129_ calibrate _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout81 vss net81 net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_255_ _076_ vss vdd _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output40_I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__304__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_55 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_307_ vdd vss _114_ _113_ _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput36 result[9] net36 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 ctlp[8] net25 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__200__I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_99 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout60 net60 vss vdd net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout71 vss net71 net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_323_ vss _015_ _128_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_306_ vss _113_ _057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_237_ vdd vss net40 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_57 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout50 net50 vss vdd net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_236_ net40 vss vdd _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_305_ vdd vss _112_ net1 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__206__I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__209__I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_output19_I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout51 vss net51 net52 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_252_ vdd vss cal_itt\[0\] _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout62 net62 vss vdd net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xfanout63 net63 vss vdd net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout52 net52 vss vdd net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout74 vss net74 net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_449_ _038_ en_co_clk net55 vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_217_ vss net26 _052_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput18 ctlp[1] net18 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_250_ vss _072_ _071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout53 net53 vss vdd net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout75 vss net75 net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__216__A2 vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_302_ vdd vss _012_ _093_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_233_ vss net39 _063_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ vdd vss _052_ mask\[9\] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput19 ctlp[2] net19 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_378_ vdd vss _033_ _160_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout66 vss net66 net68 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_300_ vdd vss _011_ _104_ _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_376_ vss _164_ _163_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_230_ vdd vss _062_ _060_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_428_ _017_ state\[2\] net53 vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_11_64 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 vss net2 clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output22_I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__282__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout57 vss net57 net65 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout79 vss net79 net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout68 vss net68 net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_18_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__277__I vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_427_ _016_ state\[1\] net53 vdd vss net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_17_161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_358_ vdd vss _053_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout58 net58 vss vdd net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout69 vss net69 net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_374_ vdd _061_ _056_ _162_ calibrate vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 vss net4 en vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_426_ _015_ state\[0\] net64 vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_211_ vss net24 _050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net49 vss vdd net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__303__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_54 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_286_ vdd vss _005_ _094_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_355_ vdd vss _149_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_371_ vss _032_ _159_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_285_ net28 vdd vss _101_ mask\[1\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_423_ _012_ net35 net55 vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_199_ net20 vss vdd _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_284_ vdd vss _004_ _094_ _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_422_ _011_ net34 net61 vss net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output36_I vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_353_ vdd vss _148_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_336_ vdd vss _138_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_198_ vdd vss _046_ mask\[3\] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_266_ vdd vss _055_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_197_ vdd vss net19 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_318_ vdd vss _124_ _115_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__409__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_24 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_403_ vdd vss _183_ cal_count\[2\] _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_334_ vss _137_ _132_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_90 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output41_I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_196_ net19 vss vdd _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ vss _070_ _069_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_38 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__409__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_60 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_332_ _126_ vdd vss _017_ _127_ _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_401_ vdd _180_ _179_ _181_ _174_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_194_ vss net8 net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_246_ vss _068_ _055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_193_ net18 vss vdd _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_400_ vdd vss _180_ cal_count\[1\] _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_331_ _134_ vdd vss _135_ _086_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_245_ vdd vss net6 _067_ net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_314_ vdd vss _121_ _085_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_261_ vss _081_ _059_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_192_ vdd vss _044_ mask\[1\] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_330_ vdd vss _134_ _133_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ vdd vss _120_ _059_ _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__190__I vss _043_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_244_ vdd vss en_co_clk _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__257__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_243_ vdd vss net47 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_87 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_98 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_242_ net47 vss vdd _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_15_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_310_ _090_ vdd vss _117_ _060_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2$1
X_207_ vdd vss _049_ mask\[6\] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_240_ vdd vss net41 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_368_ vdd vss trim_mask\[4\] _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_78 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_222_ vdd vss net38 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_221_ vss net38 _054_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_270 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_419_ _008_ net31 net60 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_79 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout58_I vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__408__A2 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_366_ vdd vss trim_mask\[3\] _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_220_ vdd vss _054_ trim_val\[0\] _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_418_ _007_ net30 net60 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_349_ vdd vss _146_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output21_I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_28 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_382_ vdd vss _035_ _160_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_279_ vdd vss _096_ _090_ state\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output14_I vss net14 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_94 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__243__I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I vss rstn vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput40 trim[2] net40 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_416_ _005_ net28 net62 vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_13_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_347_ vdd vss _145_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_201_ vdd vss _047_ mask\[4\] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 result[3] net30 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput6 clkc net6 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
.ends

.subckt saradc trim3 trim2 trim0 trim1 trim4 trimb3 trimb2 trimb0 trimb1 trimb4 cmp_outn
+ cmp_outp cmp_vinn cmp_vinp vss ctlp2 ctlp1 ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9
+ ctlp0 vdd ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctln8 ctln9 ctln0 cmp_clkc sample
+ vinn rstn clk en cal valid vinp result0 result1 result2 result3 result4 result5
+ result6 result7 result8 result9
Xlatch_0 latch_0/Qn vdd cmp_outp cmp_outn vss latch
Xbuffer_0 buffer_0/in cmp_clkc vdd vss buffer
Xdacp_0 ctlp0 vinp vdd ctlp2 ctlp1 ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9 cmp_vinp
+ dacp_0/ndum dacp_0/n1 dacp_0/n2 dacp_0/n3 dacp_0/n4 dacp_0/n5 dacp_0/n6 dacp_0/n7
+ dacp_0/n8 dacp_0/n9 dacp_0/n0 sample dacp_0/bootstrapped_sw_0/vbsh vdd vss dacp
Xdacn_0 vinn vdd ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctln8 ctln9 ctln0 cmp_vinn
+ dacn_0/ndum dacn_0/n1 dacn_0/n2 dacn_0/n3 dacn_0/n4 dacn_0/n5 dacn_0/n6 dacn_0/n7
+ dacn_0/n8 dacn_0/n9 dacn_0/n0 sample vdd dacn_0/bootstrapped_sw$1_0/vbsh vss dacn
Xcomparator_0 vdd cmp_outp cmp_outn cmp_vinp cmp_vinn trim3 trimb0 trimb3 comparator_0/diff
+ comparator_0/ip comparator_0/in cmp_clkc trim4 trim2 trim1 trim0 trimb4 trimb2 vss
+ trimb1 comparator
Xmim_cap_boss_0 vss vdd mim_cap_boss
Xmim_cap_boss_1 vss vdd mim_cap_boss
Xsarlogic_0 ctln0 ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctln8 ctln9 ctlp0 ctlp1
+ ctlp2 ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9 cal clk buffer_0/in vdd en result0
+ result1 result2 result3 result4 result5 result6 result7 result8 result9 rstn sample
+ trim0 trim1 trim2 trim3 trim4 trimb0 trimb1 trimb2 trimb3 trimb4 valid vdd vss sarlogic
.ends

