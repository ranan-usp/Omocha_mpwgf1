* NGSPICE file created from carray_in.ext - technology: gf180mcuD

.subckt carray_in n1 n2 n3 n4 n5 n6 n7 n8 n9 n0 dac_out
.ends

