* NGSPICE file created from comparator.ext - technology: gf180mcuD

.subckt XMdiff_cmp G D S a_n424_n324#
X0 S G D a_n424_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X1 D G S a_n424_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.062705f
C1 S G 0.005736f
C2 S D 0.076395f
C3 S a_n424_n324# 0.226354f
C4 D a_n424_n324# 0.027968f
C5 G a_n424_n324# 0.714768f
.ends

.subckt XM3_trims a_n2052_n100# a_n2668_n324# a_n1808_n100# a_n1948_n183# a_n1564_n100#
+ a_n2524_n100# a_n1704_n183# a_n2296_n100# a_n2192_n183# a_n2436_n183#
X0 a_n2052_n100# a_n2192_n183# a_n2296_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n1564_n100# a_n1704_n183# a_n1808_n100# a_n2668_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X2 a_n1808_n100# a_n1948_n183# a_n2052_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_n2296_n100# a_n2436_n183# a_n2524_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
C0 a_n1564_n100# a_n1704_n183# 0.002868f
C1 a_n2052_n100# a_n2296_n100# 0.038197f
C2 a_n2436_n183# a_n2192_n183# 0.039785f
C3 a_n2296_n100# a_n2436_n183# 0.002868f
C4 a_n2296_n100# a_n2524_n100# 0.038197f
C5 a_n1808_n100# a_n1948_n183# 0.002868f
C6 a_n1948_n183# a_n2192_n183# 0.039785f
C7 a_n1564_n100# a_n1808_n100# 0.038197f
C8 a_n2296_n100# a_n2192_n183# 0.002868f
C9 a_n1808_n100# a_n1704_n183# 0.002868f
C10 a_n1808_n100# a_n2052_n100# 0.038197f
C11 a_n1704_n183# a_n1948_n183# 0.039785f
C12 a_n2524_n100# a_n2436_n183# 0.002868f
C13 a_n2052_n100# a_n2192_n183# 0.002868f
C14 a_n2052_n100# a_n1948_n183# 0.002868f
C15 a_n1564_n100# a_n2668_n324# 0.061257f
C16 a_n1808_n100# a_n2668_n324# 0.036353f
C17 a_n2052_n100# a_n2668_n324# 0.036353f
C18 a_n2296_n100# a_n2668_n324# 0.036353f
C19 a_n2524_n100# a_n2668_n324# 0.113177f
C20 a_n1704_n183# a_n2668_n324# 0.334286f
C21 a_n1948_n183# a_n2668_n324# 0.306841f
C22 a_n2192_n183# a_n2668_n324# 0.30709f
C23 a_n2436_n183# a_n2668_n324# 0.34169f
.ends

.subckt XM2_trims a_n4456_n324# a_n3948_n183# a_n3808_n100# a_n4280_n100# a_n4052_n100#
+ a_n4192_n183# a_n4456_252#
X0 a_n4052_n100# a_n4192_n183# a_n4280_n100# a_n4456_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X1 a_n3808_n100# a_n3948_n183# a_n4052_n100# a_n4456_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_n4052_n100# a_n4192_n183# 0.002868f
C1 a_n3948_n183# a_n4192_n183# 0.039785f
C2 a_n4052_n100# a_n3948_n183# 0.002868f
C3 a_n3808_n100# a_n4052_n100# 0.038197f
C4 a_n4280_n100# a_n4192_n183# 0.002868f
C5 a_n3808_n100# a_n3948_n183# 0.002868f
C6 a_n4052_n100# a_n4280_n100# 0.038197f
C7 a_n3808_n100# a_n4456_n324# 0.061257f
C8 a_n4052_n100# a_n4456_n324# 0.036353f
C9 a_n4280_n100# a_n4456_n324# 0.061257f
C10 a_n3948_n183# a_n4456_n324# 0.334154f
C11 a_n4192_n183# a_n4456_n324# 0.334154f
.ends

.subckt XM1_trims G D a_n5302_n324# S a_n5302_252#
X0 D G S a_n5302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 S G 0.002868f
C2 D G 0.002868f
C3 D a_n5302_n324# 0.061257f
C4 S a_n5302_n324# 0.061257f
C5 G a_n5302_n324# 0.361695f
.ends

.subckt XM4_trims a_436_n100# a_192_n100# a_n1188_n324# a_n296_n100# a_784_n183# a_n192_n183#
+ a_n436_n183# a_540_n183# a_n52_n100# a_924_n100# a_680_n100# a_n1012_n100# a_n784_n100#
+ a_n924_n183# a_n680_n183# a_n540_n100# a_296_n183# a_52_n183#
X0 a_436_n100# a_296_n183# a_192_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n784_n100# a_n924_n183# a_n1012_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X2 a_192_n100# a_52_n183# a_n52_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_680_n100# a_540_n183# a_436_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X4 a_924_n100# a_784_n183# a_680_n100# a_n1188_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X5 a_n52_n100# a_n192_n183# a_n296_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X6 a_n296_n100# a_n436_n183# a_n540_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X7 a_n540_n100# a_n680_n183# a_n784_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_924_n100# a_784_n183# 0.002868f
C1 a_n52_n100# a_52_n183# 0.002868f
C2 a_n192_n183# a_n436_n183# 0.039785f
C3 a_n784_n100# a_n540_n100# 0.038197f
C4 a_n1012_n100# a_n924_n183# 0.002868f
C5 a_n540_n100# a_n296_n100# 0.038197f
C6 a_n436_n183# a_n296_n100# 0.002868f
C7 a_192_n100# a_296_n183# 0.002868f
C8 a_540_n183# a_296_n183# 0.039785f
C9 a_n784_n100# a_n1012_n100# 0.038197f
C10 a_n680_n183# a_n540_n100# 0.002868f
C11 a_n436_n183# a_n680_n183# 0.039785f
C12 a_680_n100# a_540_n183# 0.002868f
C13 a_n784_n100# a_n924_n183# 0.002868f
C14 a_680_n100# a_924_n100# 0.038197f
C15 a_296_n183# a_52_n183# 0.039785f
C16 a_n680_n183# a_n924_n183# 0.039785f
C17 a_n192_n183# a_n296_n100# 0.002868f
C18 a_436_n100# a_296_n183# 0.002868f
C19 a_n436_n183# a_n540_n100# 0.002868f
C20 a_n52_n100# a_n192_n183# 0.002868f
C21 a_680_n100# a_784_n183# 0.002868f
C22 a_680_n100# a_436_n100# 0.038197f
C23 a_n784_n100# a_n680_n183# 0.002868f
C24 a_192_n100# a_n52_n100# 0.038197f
C25 a_52_n183# a_n192_n183# 0.039785f
C26 a_n52_n100# a_n296_n100# 0.038197f
C27 a_192_n100# a_52_n183# 0.002868f
C28 a_784_n183# a_540_n183# 0.039785f
C29 a_436_n100# a_540_n183# 0.002868f
C30 a_436_n100# a_192_n100# 0.038197f
C31 a_924_n100# a_n1188_n324# 0.113177f
C32 a_680_n100# a_n1188_n324# 0.036353f
C33 a_436_n100# a_n1188_n324# 0.036353f
C34 a_192_n100# a_n1188_n324# 0.036353f
C35 a_n52_n100# a_n1188_n324# 0.036353f
C36 a_n296_n100# a_n1188_n324# 0.036353f
C37 a_n540_n100# a_n1188_n324# 0.036353f
C38 a_n784_n100# a_n1188_n324# 0.036353f
C39 a_n1012_n100# a_n1188_n324# 0.061257f
C40 a_784_n183# a_n1188_n324# 0.34169f
C41 a_540_n183# a_n1188_n324# 0.30709f
C42 a_296_n183# a_n1188_n324# 0.306841f
C43 a_52_n183# a_n1188_n324# 0.306744f
C44 a_n192_n183# a_n1188_n324# 0.306698f
C45 a_n436_n183# a_n1188_n324# 0.306672f
C46 a_n680_n183# a_n1188_n324# 0.306613f
C47 a_n924_n183# a_n1188_n324# 0.334154f
.ends

.subckt XM0_trims G D a_n5334_252# a_n5334_n324# S
X0 S G D a_n5334_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S G 0.002868f
C1 D G 0.002868f
C2 S D 0.038197f
C3 S a_n5334_n324# 0.061257f
C4 D a_n5334_n324# 0.061257f
C5 G a_n5334_n324# 0.361695f
.ends

.subckt trim_switch d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 temp
XXM3_trims_0 n3 temp temp d_3 n3 n3 d_3 temp d_3 d_3 XM3_trims
XXM2_trims_0 temp d_2 n2 n2 temp d_2 temp XM2_trims
XXM1_trims_0 d_1 n1 temp temp temp XM1_trims
XXM4_trims_0 n4 temp temp temp d_4 d_4 d_4 d_4 n4 n4 temp n4 temp d_4 d_4 n4 d_4 d_4
+ XM4_trims
XXM0_trims_0 d_0 n0 temp temp temp XM0_trims
C0 n2 temp 0.250074f
C1 n1 n0 0.025226f
C2 d_2 d_3 0.03061f
C3 d_2 temp 0.167792f
C4 n4 n1 0.068796f
C5 d_2 d_0 0.047211f
C6 n3 d_3 0.171874f
C7 n3 temp 0.525466f
C8 temp n0 0.099633f
C9 n2 d_2 0.052339f
C10 n4 temp 0.911975f
C11 n0 d_0 0.05352f
C12 n1 temp 0.099633f
C13 n1 d_1 0.05352f
C14 n2 n3 0.068796f
C15 n2 n0 0.068796f
C16 n4 d_4 0.398929f
C17 temp d_3 0.296319f
C18 d_1 temp 0.066702f
C19 temp d_0 0.061234f
C20 d_1 d_0 0.106626f
C21 d_4 temp 0.548654f
C22 d_4 d_1 0.02706f
C23 temp 0 2.446552f
C24 n0 0 0.124932f
C25 d_0 0 0.439168f
C26 n4 0 1.16294f
C27 d_4 0 2.753248f
C28 n1 0 0.124932f
C29 d_1 0 0.45424f
C30 n2 0 0.387627f
C31 d_2 0 0.774668f
C32 n3 0 0.70735f
C33 d_3 0 1.473152f
.ends

.subckt trim d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n3 drain n2 vss
Xtrim_switch_0 d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 vss trim_switch
C0 d_0 n0 0.010314f
C1 n4 n2 0.616308f
C2 n3 n2 0.584482f
C3 drain n2 3.213024f
C4 n1 n2 0.092902f
C5 n4 vss 0.206884f
C6 n0 n2 0.116341f
C7 n3 vss 0.139026f
C8 drain vss 3.229077f
C9 n1 vss 0.017014f
C10 vss n0 0.017474f
C11 n1 d_1 0.009441f
C12 n4 n3 1.599582f
C13 n4 drain 12.877382f
C14 n4 n1 0.166777f
C15 n3 drain 6.427484f
C16 n3 n1 0.087807f
C17 n1 drain 1.60623f
C18 n4 n0 0.166348f
C19 n3 n0 0.087807f
C20 drain n0 1.60623f
C21 n1 n0 0.506269f
C22 n4 d_4 0.001311f
C23 vss n2 0.024554f
C24 d_1 n2 0.00105f
C25 n0 0 0.627477f
C26 n1 0 0.643951f
C27 n4 0 4.635427f
C28 drain 0 -9.135383f
C29 n2 0 1.998525f
C30 n3 0 3.342805f
C31 vss 0 4.401155f
C32 d_0 0 0.431586f
C33 d_4 0 2.753248f
C34 d_1 0 0.446833f
C35 d_2 0 0.774668f
C36 d_3 0 1.473152f
.ends

.subckt XMinp_cmp G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 S D 0.038197f
C2 S G 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM4_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.019807f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMl4_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.021497f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12132f
.ends

.subckt XMl3_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.021497f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XM3_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.021497f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XMinn_cmp G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 S D 0.038197f
C2 S G 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM2_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.021497f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XMl2_cmp G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.368221f
.ends

.subckt XM1_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 S w_n319_n356# 0.021189f
C2 G D 0.002389f
C3 S D 0.045397f
C4 S G 0.002389f
C5 w_n319_n356# D 0.019807f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMl1_cmp G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.368221f
.ends

.subckt comparator trim1 trim0 trim2 trim3 trim4 trimb4 trimb1 trimb0 trimb2 trimb3
+ vp vn outp outn clkc vss vdd
XXMdiff_cmp_0 clkc diff vss vss XMdiff_cmp
Xtrim_0 trimb0 trimb4 trimb1 trimb2 trimb3 trim_0/n1 trim_0/n4 trim_0/n0 trim_0/n3
+ ip trim_0/n2 vss trim
Xtrim_1 trim0 trim4 trim1 trim2 trim3 trim_1/n1 trim_1/n4 trim_1/n0 trim_1/n3 in trim_1/n2
+ vss trim
XXMinp_cmp_0 vp ip vss vss diff XMinp_cmp
XXM4_cmp_0 clkc ip vdd vdd vss XM4_cmp
XXMl4_cmp_0 outn outp vdd vdd vss XMl4_cmp
XXMl3_cmp_0 outp outn vdd vdd vss XMl3_cmp
XXM3_cmp_0 clkc outp vdd vdd vss XM3_cmp
XXMinn_cmp_0 vn in vss vss diff XMinn_cmp
XXM2_cmp_0 clkc outn vdd vdd vss XM2_cmp
XXMl2_cmp_0 outn outp vss ip XMl2_cmp
XXM1_cmp_0 clkc in vdd vdd vss XM1_cmp
XXMl1_cmp_0 outp outn vss in XMl1_cmp
C0 trimb4 trim_0/n4 0.002904f
C1 clkc diff 0.019234f
C2 trimb2 vss 0.037673f
C3 trim2 trim4 0.001666f
C4 vp vss 0.026857f
C5 trim4 vss 0.154051f
C6 diff ip 0.098316f
C7 trim_1/n0 in 1.606869f
C8 clkc outp 0.295692f
C9 clkc vdd 0.289807f
C10 outp ip 0.10316f
C11 diff vn 0.009142f
C12 ip vdd 0.108547f
C13 trim1 trim_1/n4 0.001799f
C14 trim_1/n4 trim_1/n3 0.241184f
C15 trim_0/n4 ip 12.853152f
C16 trim0 trim1 0.713549f
C17 outp vn 0.19705f
C18 vn vdd 0.069074f
C19 trim_0/n0 trim_0/n4 0.032158f
C20 in trim_1/n3 6.426837f
C21 outn in 0.103141f
C22 trimb4 trimb1 0.397758f
C23 outn clkc 0.29566f
C24 trim_1/n4 trim_1/n1 0.032158f
C25 outn ip 0.018487f
C26 diff vss 0.080305f
C27 trim_1/n1 in 1.606869f
C28 trimb1 trimb0 0.713549f
C29 outn vn 0.199287f
C30 vp diff 0.009142f
C31 trim_1/n4 in 12.853152f
C32 trim_0/n3 trim_0/n4 0.241184f
C33 outp vss 0.458491f
C34 vp outp 0.256864f
C35 vp vdd 0.069074f
C36 trim_0/n4 vss 0.083236f
C37 clkc in 0.528032f
C38 trimb4 trimb0 0.002527f
C39 trim_0/n2 trim_0/n4 0.128631f
C40 trim2 trim3 0.902342f
C41 vss trim3 0.039536f
C42 trim1 vss 0.091365f
C43 trim_1/n4 trim_1/n2 0.128631f
C44 outn vss 0.457585f
C45 in vn 0.448228f
C46 trim1 trim4 0.397758f
C47 trim_0/n1 trim_0/n4 0.032158f
C48 clkc ip 0.528032f
C49 vp outn 0.159375f
C50 in trim_1/n2 3.218424f
C51 trimb1 vss 0.091365f
C52 clkc vn 0.133362f
C53 trim_0/n0 ip 1.606869f
C54 diff outp 0.005373f
C55 outp vdd 0.454873f
C56 trim_1/n4 vss 0.083236f
C57 trim0 trim2 0.786004f
C58 trim0 vss 0.040411f
C59 trimb4 vss 0.154051f
C60 trim_1/n4 trim4 0.002904f
C61 trimb4 trimb2 0.001666f
C62 in vss 3.44372f
C63 trim0 trim4 0.002527f
C64 trim_0/n3 ip 6.426837f
C65 clkc vss 0.615121f
C66 outn diff 0.002551f
C67 trimb0 vss 0.040411f
C68 vp clkc 0.133362f
C69 trimb2 trimb0 0.786004f
C70 vss ip 3.443847f
C71 outn outp 1.39519f
C72 vp ip 0.448228f
C73 outn vdd 0.503383f
C74 vn vss 0.026857f
C75 vp vn 0.125877f
C76 trim_0/n2 ip 3.218424f
C77 trimb1 trim_0/n4 0.001799f
C78 trim_0/n1 ip 1.606869f
C79 trimb3 vss 0.039536f
C80 trimb2 trimb3 0.902342f
C81 diff in 0.098316f
C82 trim_0/n1 trim_0/n0 0.032158f
C83 trim_1/n0 trim_1/n1 0.032158f
C84 outp in 0.018491f
C85 trim2 vss 0.037673f
C86 in vdd 0.108547f
C87 trim_1/n4 trim_1/n0 0.032158f
C88 outp 0 2.271068f
C89 outn 0 2.225997f
C90 vdd 0 9.215822f
C91 vn 0 1.207921f
C92 vp 0 1.193091f
C93 trim_1/n0 0 0.627477f
C94 trim_1/n1 0 0.643951f
C95 trim_1/n4 0 4.635427f
C96 in 0 -7.798843f
C97 trim_1/n2 0 1.998525f
C98 trim_1/n3 0 3.342805f
C99 vss 0 12.362443f
C100 trim0 0 1.018331f
C101 trim4 0 3.13965f
C102 trim1 0 1.001356f
C103 trim2 0 1.580338f
C104 trim3 0 3.420755f
C105 trim_0/n0 0 0.627477f
C106 trim_0/n1 0 0.643951f
C107 trim_0/n4 0 4.635427f
C108 ip 0 -7.798843f
C109 trim_0/n2 0 1.998525f
C110 trim_0/n3 0 3.342805f
C111 trimb0 0 1.018331f
C112 trimb4 0 3.13965f
C113 trimb1 0 1.001356f
C114 trimb2 0 1.580338f
C115 trimb3 0 3.420755f
C116 diff 0 0.21132f
C117 clkc 0 4.576592f
.ends

