** sch_path: /home/oe23ranan/gf_analog/xschem/sar_10b/dac/carray.sch
**.subckt carray top n6 n0 n5 n4 n2 ndum n3 n1 n7 n8 n9
*.iopin carray_top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
*.iopin n8
*.iopin n9
*.iopin vss
xcdum carray_top ndum unitcap
xc0 carray_top n0 unitcap
xc1[1] carray_top n1 unitcap
xc1[0] carray_top n1 unitcap
xc2[3] carray_top n2 unitcap
xc2[2] carray_top n2 unitcap
xc2[1] carray_top n2 unitcap
xc2[0] carray_top n2 unitcap
xc3[7] carray_top n3 unitcap
xc3[6] carray_top n3 unitcap
xc3[5] carray_top n3 unitcap
xc3[4] carray_top n3 unitcap
xc3[3] carray_top n3 unitcap
xc3[2] carray_top n3 unitcap
xc3[1] carray_top n3 unitcap
xc3[0] carray_top n3 unitcap
xc4[15] carray_top n4 unitcap
xc4[14] carray_top n4 unitcap
xc4[13] carray_top n4 unitcap
xc4[12] carray_top n4 unitcap
xc4[11] carray_top n4 unitcap
xc4[10] carray_top n4 unitcap
xc4[9] carray_top n4 unitcap
xc4[8] carray_top n4 unitcap
xc4[7] carray_top n4 unitcap
xc4[6] carray_top n4 unitcap
xc4[5] carray_top n4 unitcap
xc4[4] carray_top n4 unitcap
xc4[3] carray_top n4 unitcap
xc4[2] carray_top n4 unitcap
xc4[1] carray_top n4 unitcap
xc4[0] carray_top n4 unitcap
xc5[31] carray_top n5 unitcap
xc5[30] carray_top n5 unitcap
xc5[29] carray_top n5 unitcap
xc5[28] carray_top n5 unitcap
xc5[27] carray_top n5 unitcap
xc5[26] carray_top n5 unitcap
xc5[25] carray_top n5 unitcap
xc5[24] carray_top n5 unitcap
xc5[23] carray_top n5 unitcap
xc5[22] carray_top n5 unitcap
xc5[21] carray_top n5 unitcap
xc5[20] carray_top n5 unitcap
xc5[19] carray_top n5 unitcap
xc5[18] carray_top n5 unitcap
xc5[17] carray_top n5 unitcap
xc5[16] carray_top n5 unitcap
xc5[15] carray_top n5 unitcap
xc5[14] carray_top n5 unitcap
xc5[13] carray_top n5 unitcap
xc5[12] carray_top n5 unitcap
xc5[11] carray_top n5 unitcap
xc5[10] carray_top n5 unitcap
xc5[9] carray_top n5 unitcap
xc5[8] carray_top n5 unitcap
xc5[7] carray_top n5 unitcap
xc5[6] carray_top n5 unitcap
xc5[5] carray_top n5 unitcap
xc5[4] carray_top n5 unitcap
xc5[3] carray_top n5 unitcap
xc5[2] carray_top n5 unitcap
xc5[1] carray_top n5 unitcap
xc5[0] carray_top n5 unitcap
xc6[63] carray_top n6 unitcap
xc6[62] carray_top n6 unitcap
xc6[61] carray_top n6 unitcap
xc6[60] carray_top n6 unitcap
xc6[59] carray_top n6 unitcap
xc6[58] carray_top n6 unitcap
xc6[57] carray_top n6 unitcap
xc6[56] carray_top n6 unitcap
xc6[55] carray_top n6 unitcap
xc6[54] carray_top n6 unitcap
xc6[53] carray_top n6 unitcap
xc6[52] carray_top n6 unitcap
xc6[51] carray_top n6 unitcap
xc6[50] carray_top n6 unitcap
xc6[49] carray_top n6 unitcap
xc6[48] carray_top n6 unitcap
xc6[47] carray_top n6 unitcap
xc6[46] carray_top n6 unitcap
xc6[45] carray_top n6 unitcap
xc6[44] carray_top n6 unitcap
xc6[43] carray_top n6 unitcap
xc6[42] carray_top n6 unitcap
xc6[41] carray_top n6 unitcap
xc6[40] carray_top n6 unitcap
xc6[39] carray_top n6 unitcap
xc6[38] carray_top n6 unitcap
xc6[37] carray_top n6 unitcap
xc6[36] carray_top n6 unitcap
xc6[35] carray_top n6 unitcap
xc6[34] carray_top n6 unitcap
xc6[33] carray_top n6 unitcap
xc6[32] carray_top n6 unitcap
xc6[31] carray_top n6 unitcap
xc6[30] carray_top n6 unitcap
xc6[29] carray_top n6 unitcap
xc6[28] carray_top n6 unitcap
xc6[27] carray_top n6 unitcap
xc6[26] carray_top n6 unitcap
xc6[25] carray_top n6 unitcap
xc6[24] carray_top n6 unitcap
xc6[23] carray_top n6 unitcap
xc6[22] carray_top n6 unitcap
xc6[21] carray_top n6 unitcap
xc6[20] carray_top n6 unitcap
xc6[19] carray_top n6 unitcap
xc6[18] carray_top n6 unitcap
xc6[17] carray_top n6 unitcap
xc6[16] carray_top n6 unitcap
xc6[15] carray_top n6 unitcap
xc6[14] carray_top n6 unitcap
xc6[13] carray_top n6 unitcap
xc6[12] carray_top n6 unitcap
xc6[11] carray_top n6 unitcap
xc6[10] carray_top n6 unitcap
xc6[9] carray_top n6 unitcap
xc6[8] carray_top n6 unitcap
xc6[7] carray_top n6 unitcap
xc6[6] carray_top n6 unitcap
xc6[5] carray_top n6 unitcap
xc6[4] carray_top n6 unitcap
xc6[3] carray_top n6 unitcap
xc6[2] carray_top n6 unitcap
xc6[1] carray_top n6 unitcap
xc6[0] carray_top n6 unitcap
xc7[127] carray_top n7 unitcap
xc7[126] carray_top n7 unitcap
xc7[125] carray_top n7 unitcap
xc7[124] carray_top n7 unitcap
xc7[123] carray_top n7 unitcap
xc7[122] carray_top n7 unitcap
xc7[121] carray_top n7 unitcap
xc7[120] carray_top n7 unitcap
xc7[119] carray_top n7 unitcap
xc7[118] carray_top n7 unitcap
xc7[117] carray_top n7 unitcap
xc7[116] carray_top n7 unitcap
xc7[115] carray_top n7 unitcap
xc7[114] carray_top n7 unitcap
xc7[113] carray_top n7 unitcap
xc7[112] carray_top n7 unitcap
xc7[111] carray_top n7 unitcap
xc7[110] carray_top n7 unitcap
xc7[109] carray_top n7 unitcap
xc7[108] carray_top n7 unitcap
xc7[107] carray_top n7 unitcap
xc7[106] carray_top n7 unitcap
xc7[105] carray_top n7 unitcap
xc7[104] carray_top n7 unitcap
xc7[103] carray_top n7 unitcap
xc7[102] carray_top n7 unitcap
xc7[101] carray_top n7 unitcap
xc7[100] carray_top n7 unitcap
xc7[99] carray_top n7 unitcap
xc7[98] carray_top n7 unitcap
xc7[97] carray_top n7 unitcap
xc7[96] carray_top n7 unitcap
xc7[95] carray_top n7 unitcap
xc7[94] carray_top n7 unitcap
xc7[93] carray_top n7 unitcap
xc7[92] carray_top n7 unitcap
xc7[91] carray_top n7 unitcap
xc7[90] carray_top n7 unitcap
xc7[89] carray_top n7 unitcap
xc7[88] carray_top n7 unitcap
xc7[87] carray_top n7 unitcap
xc7[86] carray_top n7 unitcap
xc7[85] carray_top n7 unitcap
xc7[84] carray_top n7 unitcap
xc7[83] carray_top n7 unitcap
xc7[82] carray_top n7 unitcap
xc7[81] carray_top n7 unitcap
xc7[80] carray_top n7 unitcap
xc7[79] carray_top n7 unitcap
xc7[78] carray_top n7 unitcap
xc7[77] carray_top n7 unitcap
xc7[76] carray_top n7 unitcap
xc7[75] carray_top n7 unitcap
xc7[74] carray_top n7 unitcap
xc7[73] carray_top n7 unitcap
xc7[72] carray_top n7 unitcap
xc7[71] carray_top n7 unitcap
xc7[70] carray_top n7 unitcap
xc7[69] carray_top n7 unitcap
xc7[68] carray_top n7 unitcap
xc7[67] carray_top n7 unitcap
xc7[66] carray_top n7 unitcap
xc7[65] carray_top n7 unitcap
xc7[64] carray_top n7 unitcap
xc7[63] carray_top n7 unitcap
xc7[62] carray_top n7 unitcap
xc7[61] carray_top n7 unitcap
xc7[60] carray_top n7 unitcap
xc7[59] carray_top n7 unitcap
xc7[58] carray_top n7 unitcap
xc7[57] carray_top n7 unitcap
xc7[56] carray_top n7 unitcap
xc7[55] carray_top n7 unitcap
xc7[54] carray_top n7 unitcap
xc7[53] carray_top n7 unitcap
xc7[52] carray_top n7 unitcap
xc7[51] carray_top n7 unitcap
xc7[50] carray_top n7 unitcap
xc7[49] carray_top n7 unitcap
xc7[48] carray_top n7 unitcap
xc7[47] carray_top n7 unitcap
xc7[46] carray_top n7 unitcap
xc7[45] carray_top n7 unitcap
xc7[44] carray_top n7 unitcap
xc7[43] carray_top n7 unitcap
xc7[42] carray_top n7 unitcap
xc7[41] carray_top n7 unitcap
xc7[40] carray_top n7 unitcap
xc7[39] carray_top n7 unitcap
xc7[38] carray_top n7 unitcap
xc7[37] carray_top n7 unitcap
xc7[36] carray_top n7 unitcap
xc7[35] carray_top n7 unitcap
xc7[34] carray_top n7 unitcap
xc7[33] carray_top n7 unitcap
xc7[32] carray_top n7 unitcap
xc7[31] carray_top n7 unitcap
xc7[30] carray_top n7 unitcap
xc7[29] carray_top n7 unitcap
xc7[28] carray_top n7 unitcap
xc7[27] carray_top n7 unitcap
xc7[26] carray_top n7 unitcap
xc7[25] carray_top n7 unitcap
xc7[24] carray_top n7 unitcap
xc7[23] carray_top n7 unitcap
xc7[22] carray_top n7 unitcap
xc7[21] carray_top n7 unitcap
xc7[20] carray_top n7 unitcap
xc7[19] carray_top n7 unitcap
xc7[18] carray_top n7 unitcap
xc7[17] carray_top n7 unitcap
xc7[16] carray_top n7 unitcap
xc7[15] carray_top n7 unitcap
xc7[14] carray_top n7 unitcap
xc7[13] carray_top n7 unitcap
xc7[12] carray_top n7 unitcap
xc7[11] carray_top n7 unitcap
xc7[10] carray_top n7 unitcap
xc7[9] carray_top n7 unitcap
xc7[8] carray_top n7 unitcap
xc7[7] carray_top n7 unitcap
xc7[6] carray_top n7 unitcap
xc7[5] carray_top n7 unitcap
xc7[4] carray_top n7 unitcap
xc7[3] carray_top n7 unitcap
xc7[2] carray_top n7 unitcap
xc7[1] carray_top n7 unitcap
xc7[0] carray_top n7 unitcap
xc8[255] carray_top n8 unitcap
xc8[254] carray_top n8 unitcap
xc8[253] carray_top n8 unitcap
xc8[252] carray_top n8 unitcap
xc8[251] carray_top n8 unitcap
xc8[250] carray_top n8 unitcap
xc8[249] carray_top n8 unitcap
xc8[248] carray_top n8 unitcap
xc8[247] carray_top n8 unitcap
xc8[246] carray_top n8 unitcap
xc8[245] carray_top n8 unitcap
xc8[244] carray_top n8 unitcap
xc8[243] carray_top n8 unitcap
xc8[242] carray_top n8 unitcap
xc8[241] carray_top n8 unitcap
xc8[240] carray_top n8 unitcap
xc8[239] carray_top n8 unitcap
xc8[238] carray_top n8 unitcap
xc8[237] carray_top n8 unitcap
xc8[236] carray_top n8 unitcap
xc8[235] carray_top n8 unitcap
xc8[234] carray_top n8 unitcap
xc8[233] carray_top n8 unitcap
xc8[232] carray_top n8 unitcap
xc8[231] carray_top n8 unitcap
xc8[230] carray_top n8 unitcap
xc8[229] carray_top n8 unitcap
xc8[228] carray_top n8 unitcap
xc8[227] carray_top n8 unitcap
xc8[226] carray_top n8 unitcap
xc8[225] carray_top n8 unitcap
xc8[224] carray_top n8 unitcap
xc8[223] carray_top n8 unitcap
xc8[222] carray_top n8 unitcap
xc8[221] carray_top n8 unitcap
xc8[220] carray_top n8 unitcap
xc8[219] carray_top n8 unitcap
xc8[218] carray_top n8 unitcap
xc8[217] carray_top n8 unitcap
xc8[216] carray_top n8 unitcap
xc8[215] carray_top n8 unitcap
xc8[214] carray_top n8 unitcap
xc8[213] carray_top n8 unitcap
xc8[212] carray_top n8 unitcap
xc8[211] carray_top n8 unitcap
xc8[210] carray_top n8 unitcap
xc8[209] carray_top n8 unitcap
xc8[208] carray_top n8 unitcap
xc8[207] carray_top n8 unitcap
xc8[206] carray_top n8 unitcap
xc8[205] carray_top n8 unitcap
xc8[204] carray_top n8 unitcap
xc8[203] carray_top n8 unitcap
xc8[202] carray_top n8 unitcap
xc8[201] carray_top n8 unitcap
xc8[200] carray_top n8 unitcap
xc8[199] carray_top n8 unitcap
xc8[198] carray_top n8 unitcap
xc8[197] carray_top n8 unitcap
xc8[196] carray_top n8 unitcap
xc8[195] carray_top n8 unitcap
xc8[194] carray_top n8 unitcap
xc8[193] carray_top n8 unitcap
xc8[192] carray_top n8 unitcap
xc8[191] carray_top n8 unitcap
xc8[190] carray_top n8 unitcap
xc8[189] carray_top n8 unitcap
xc8[188] carray_top n8 unitcap
xc8[187] carray_top n8 unitcap
xc8[186] carray_top n8 unitcap
xc8[185] carray_top n8 unitcap
xc8[184] carray_top n8 unitcap
xc8[183] carray_top n8 unitcap
xc8[182] carray_top n8 unitcap
xc8[181] carray_top n8 unitcap
xc8[180] carray_top n8 unitcap
xc8[179] carray_top n8 unitcap
xc8[178] carray_top n8 unitcap
xc8[177] carray_top n8 unitcap
xc8[176] carray_top n8 unitcap
xc8[175] carray_top n8 unitcap
xc8[174] carray_top n8 unitcap
xc8[173] carray_top n8 unitcap
xc8[172] carray_top n8 unitcap
xc8[171] carray_top n8 unitcap
xc8[170] carray_top n8 unitcap
xc8[169] carray_top n8 unitcap
xc8[168] carray_top n8 unitcap
xc8[167] carray_top n8 unitcap
xc8[166] carray_top n8 unitcap
xc8[165] carray_top n8 unitcap
xc8[164] carray_top n8 unitcap
xc8[163] carray_top n8 unitcap
xc8[162] carray_top n8 unitcap
xc8[161] carray_top n8 unitcap
xc8[160] carray_top n8 unitcap
xc8[159] carray_top n8 unitcap
xc8[158] carray_top n8 unitcap
xc8[157] carray_top n8 unitcap
xc8[156] carray_top n8 unitcap
xc8[155] carray_top n8 unitcap
xc8[154] carray_top n8 unitcap
xc8[153] carray_top n8 unitcap
xc8[152] carray_top n8 unitcap
xc8[151] carray_top n8 unitcap
xc8[150] carray_top n8 unitcap
xc8[149] carray_top n8 unitcap
xc8[148] carray_top n8 unitcap
xc8[147] carray_top n8 unitcap
xc8[146] carray_top n8 unitcap
xc8[145] carray_top n8 unitcap
xc8[144] carray_top n8 unitcap
xc8[143] carray_top n8 unitcap
xc8[142] carray_top n8 unitcap
xc8[141] carray_top n8 unitcap
xc8[140] carray_top n8 unitcap
xc8[139] carray_top n8 unitcap
xc8[138] carray_top n8 unitcap
xc8[137] carray_top n8 unitcap
xc8[136] carray_top n8 unitcap
xc8[135] carray_top n8 unitcap
xc8[134] carray_top n8 unitcap
xc8[133] carray_top n8 unitcap
xc8[132] carray_top n8 unitcap
xc8[131] carray_top n8 unitcap
xc8[130] carray_top n8 unitcap
xc8[129] carray_top n8 unitcap
xc8[128] carray_top n8 unitcap
xc8[127] carray_top n8 unitcap
xc8[126] carray_top n8 unitcap
xc8[125] carray_top n8 unitcap
xc8[124] carray_top n8 unitcap
xc8[123] carray_top n8 unitcap
xc8[122] carray_top n8 unitcap
xc8[121] carray_top n8 unitcap
xc8[120] carray_top n8 unitcap
xc8[119] carray_top n8 unitcap
xc8[118] carray_top n8 unitcap
xc8[117] carray_top n8 unitcap
xc8[116] carray_top n8 unitcap
xc8[115] carray_top n8 unitcap
xc8[114] carray_top n8 unitcap
xc8[113] carray_top n8 unitcap
xc8[112] carray_top n8 unitcap
xc8[111] carray_top n8 unitcap
xc8[110] carray_top n8 unitcap
xc8[109] carray_top n8 unitcap
xc8[108] carray_top n8 unitcap
xc8[107] carray_top n8 unitcap
xc8[106] carray_top n8 unitcap
xc8[105] carray_top n8 unitcap
xc8[104] carray_top n8 unitcap
xc8[103] carray_top n8 unitcap
xc8[102] carray_top n8 unitcap
xc8[101] carray_top n8 unitcap
xc8[100] carray_top n8 unitcap
xc8[99] carray_top n8 unitcap
xc8[98] carray_top n8 unitcap
xc8[97] carray_top n8 unitcap
xc8[96] carray_top n8 unitcap
xc8[95] carray_top n8 unitcap
xc8[94] carray_top n8 unitcap
xc8[93] carray_top n8 unitcap
xc8[92] carray_top n8 unitcap
xc8[91] carray_top n8 unitcap
xc8[90] carray_top n8 unitcap
xc8[89] carray_top n8 unitcap
xc8[88] carray_top n8 unitcap
xc8[87] carray_top n8 unitcap
xc8[86] carray_top n8 unitcap
xc8[85] carray_top n8 unitcap
xc8[84] carray_top n8 unitcap
xc8[83] carray_top n8 unitcap
xc8[82] carray_top n8 unitcap
xc8[81] carray_top n8 unitcap
xc8[80] carray_top n8 unitcap
xc8[79] carray_top n8 unitcap
xc8[78] carray_top n8 unitcap
xc8[77] carray_top n8 unitcap
xc8[76] carray_top n8 unitcap
xc8[75] carray_top n8 unitcap
xc8[74] carray_top n8 unitcap
xc8[73] carray_top n8 unitcap
xc8[72] carray_top n8 unitcap
xc8[71] carray_top n8 unitcap
xc8[70] carray_top n8 unitcap
xc8[69] carray_top n8 unitcap
xc8[68] carray_top n8 unitcap
xc8[67] carray_top n8 unitcap
xc8[66] carray_top n8 unitcap
xc8[65] carray_top n8 unitcap
xc8[64] carray_top n8 unitcap
xc8[63] carray_top n8 unitcap
xc8[62] carray_top n8 unitcap
xc8[61] carray_top n8 unitcap
xc8[60] carray_top n8 unitcap
xc8[59] carray_top n8 unitcap
xc8[58] carray_top n8 unitcap
xc8[57] carray_top n8 unitcap
xc8[56] carray_top n8 unitcap
xc8[55] carray_top n8 unitcap
xc8[54] carray_top n8 unitcap
xc8[53] carray_top n8 unitcap
xc8[52] carray_top n8 unitcap
xc8[51] carray_top n8 unitcap
xc8[50] carray_top n8 unitcap
xc8[49] carray_top n8 unitcap
xc8[48] carray_top n8 unitcap
xc8[47] carray_top n8 unitcap
xc8[46] carray_top n8 unitcap
xc8[45] carray_top n8 unitcap
xc8[44] carray_top n8 unitcap
xc8[43] carray_top n8 unitcap
xc8[42] carray_top n8 unitcap
xc8[41] carray_top n8 unitcap
xc8[40] carray_top n8 unitcap
xc8[39] carray_top n8 unitcap
xc8[38] carray_top n8 unitcap
xc8[37] carray_top n8 unitcap
xc8[36] carray_top n8 unitcap
xc8[35] carray_top n8 unitcap
xc8[34] carray_top n8 unitcap
xc8[33] carray_top n8 unitcap
xc8[32] carray_top n8 unitcap
xc8[31] carray_top n8 unitcap
xc8[30] carray_top n8 unitcap
xc8[29] carray_top n8 unitcap
xc8[28] carray_top n8 unitcap
xc8[27] carray_top n8 unitcap
xc8[26] carray_top n8 unitcap
xc8[25] carray_top n8 unitcap
xc8[24] carray_top n8 unitcap
xc8[23] carray_top n8 unitcap
xc8[22] carray_top n8 unitcap
xc8[21] carray_top n8 unitcap
xc8[20] carray_top n8 unitcap
xc8[19] carray_top n8 unitcap
xc8[18] carray_top n8 unitcap
xc8[17] carray_top n8 unitcap
xc8[16] carray_top n8 unitcap
xc8[15] carray_top n8 unitcap
xc8[14] carray_top n8 unitcap
xc8[13] carray_top n8 unitcap
xc8[12] carray_top n8 unitcap
xc8[11] carray_top n8 unitcap
xc8[10] carray_top n8 unitcap
xc8[9] carray_top n8 unitcap
xc8[8] carray_top n8 unitcap
xc8[7] carray_top n8 unitcap
xc8[6] carray_top n8 unitcap
xc8[5] carray_top n8 unitcap
xc8[4] carray_top n8 unitcap
xc8[3] carray_top n8 unitcap
xc8[2] carray_top n8 unitcap
xc8[1] carray_top n8 unitcap
xc8[0] carray_top n8 unitcap
xc9[511] carray_top n9 unitcap
xc9[510] carray_top n9 unitcap
xc9[509] carray_top n9 unitcap
xc9[508] carray_top n9 unitcap
xc9[507] carray_top n9 unitcap
xc9[506] carray_top n9 unitcap
xc9[505] carray_top n9 unitcap
xc9[504] carray_top n9 unitcap
xc9[503] carray_top n9 unitcap
xc9[502] carray_top n9 unitcap
xc9[501] carray_top n9 unitcap
xc9[500] carray_top n9 unitcap
xc9[499] carray_top n9 unitcap
xc9[498] carray_top n9 unitcap
xc9[497] carray_top n9 unitcap
xc9[496] carray_top n9 unitcap
xc9[495] carray_top n9 unitcap
xc9[494] carray_top n9 unitcap
xc9[493] carray_top n9 unitcap
xc9[492] carray_top n9 unitcap
xc9[491] carray_top n9 unitcap
xc9[490] carray_top n9 unitcap
xc9[489] carray_top n9 unitcap
xc9[488] carray_top n9 unitcap
xc9[487] carray_top n9 unitcap
xc9[486] carray_top n9 unitcap
xc9[485] carray_top n9 unitcap
xc9[484] carray_top n9 unitcap
xc9[483] carray_top n9 unitcap
xc9[482] carray_top n9 unitcap
xc9[481] carray_top n9 unitcap
xc9[480] carray_top n9 unitcap
xc9[479] carray_top n9 unitcap
xc9[478] carray_top n9 unitcap
xc9[477] carray_top n9 unitcap
xc9[476] carray_top n9 unitcap
xc9[475] carray_top n9 unitcap
xc9[474] carray_top n9 unitcap
xc9[473] carray_top n9 unitcap
xc9[472] carray_top n9 unitcap
xc9[471] carray_top n9 unitcap
xc9[470] carray_top n9 unitcap
xc9[469] carray_top n9 unitcap
xc9[468] carray_top n9 unitcap
xc9[467] carray_top n9 unitcap
xc9[466] carray_top n9 unitcap
xc9[465] carray_top n9 unitcap
xc9[464] carray_top n9 unitcap
xc9[463] carray_top n9 unitcap
xc9[462] carray_top n9 unitcap
xc9[461] carray_top n9 unitcap
xc9[460] carray_top n9 unitcap
xc9[459] carray_top n9 unitcap
xc9[458] carray_top n9 unitcap
xc9[457] carray_top n9 unitcap
xc9[456] carray_top n9 unitcap
xc9[455] carray_top n9 unitcap
xc9[454] carray_top n9 unitcap
xc9[453] carray_top n9 unitcap
xc9[452] carray_top n9 unitcap
xc9[451] carray_top n9 unitcap
xc9[450] carray_top n9 unitcap
xc9[449] carray_top n9 unitcap
xc9[448] carray_top n9 unitcap
xc9[447] carray_top n9 unitcap
xc9[446] carray_top n9 unitcap
xc9[445] carray_top n9 unitcap
xc9[444] carray_top n9 unitcap
xc9[443] carray_top n9 unitcap
xc9[442] carray_top n9 unitcap
xc9[441] carray_top n9 unitcap
xc9[440] carray_top n9 unitcap
xc9[439] carray_top n9 unitcap
xc9[438] carray_top n9 unitcap
xc9[437] carray_top n9 unitcap
xc9[436] carray_top n9 unitcap
xc9[435] carray_top n9 unitcap
xc9[434] carray_top n9 unitcap
xc9[433] carray_top n9 unitcap
xc9[432] carray_top n9 unitcap
xc9[431] carray_top n9 unitcap
xc9[430] carray_top n9 unitcap
xc9[429] carray_top n9 unitcap
xc9[428] carray_top n9 unitcap
xc9[427] carray_top n9 unitcap
xc9[426] carray_top n9 unitcap
xc9[425] carray_top n9 unitcap
xc9[424] carray_top n9 unitcap
xc9[423] carray_top n9 unitcap
xc9[422] carray_top n9 unitcap
xc9[421] carray_top n9 unitcap
xc9[420] carray_top n9 unitcap
xc9[419] carray_top n9 unitcap
xc9[418] carray_top n9 unitcap
xc9[417] carray_top n9 unitcap
xc9[416] carray_top n9 unitcap
xc9[415] carray_top n9 unitcap
xc9[414] carray_top n9 unitcap
xc9[413] carray_top n9 unitcap
xc9[412] carray_top n9 unitcap
xc9[411] carray_top n9 unitcap
xc9[410] carray_top n9 unitcap
xc9[409] carray_top n9 unitcap
xc9[408] carray_top n9 unitcap
xc9[407] carray_top n9 unitcap
xc9[406] carray_top n9 unitcap
xc9[405] carray_top n9 unitcap
xc9[404] carray_top n9 unitcap
xc9[403] carray_top n9 unitcap
xc9[402] carray_top n9 unitcap
xc9[401] carray_top n9 unitcap
xc9[400] carray_top n9 unitcap
xc9[399] carray_top n9 unitcap
xc9[398] carray_top n9 unitcap
xc9[397] carray_top n9 unitcap
xc9[396] carray_top n9 unitcap
xc9[395] carray_top n9 unitcap
xc9[394] carray_top n9 unitcap
xc9[393] carray_top n9 unitcap
xc9[392] carray_top n9 unitcap
xc9[391] carray_top n9 unitcap
xc9[390] carray_top n9 unitcap
xc9[389] carray_top n9 unitcap
xc9[388] carray_top n9 unitcap
xc9[387] carray_top n9 unitcap
xc9[386] carray_top n9 unitcap
xc9[385] carray_top n9 unitcap
xc9[384] carray_top n9 unitcap
xc9[383] carray_top n9 unitcap
xc9[382] carray_top n9 unitcap
xc9[381] carray_top n9 unitcap
xc9[380] carray_top n9 unitcap
xc9[379] carray_top n9 unitcap
xc9[378] carray_top n9 unitcap
xc9[377] carray_top n9 unitcap
xc9[376] carray_top n9 unitcap
xc9[375] carray_top n9 unitcap
xc9[374] carray_top n9 unitcap
xc9[373] carray_top n9 unitcap
xc9[372] carray_top n9 unitcap
xc9[371] carray_top n9 unitcap
xc9[370] carray_top n9 unitcap
xc9[369] carray_top n9 unitcap
xc9[368] carray_top n9 unitcap
xc9[367] carray_top n9 unitcap
xc9[366] carray_top n9 unitcap
xc9[365] carray_top n9 unitcap
xc9[364] carray_top n9 unitcap
xc9[363] carray_top n9 unitcap
xc9[362] carray_top n9 unitcap
xc9[361] carray_top n9 unitcap
xc9[360] carray_top n9 unitcap
xc9[359] carray_top n9 unitcap
xc9[358] carray_top n9 unitcap
xc9[357] carray_top n9 unitcap
xc9[356] carray_top n9 unitcap
xc9[355] carray_top n9 unitcap
xc9[354] carray_top n9 unitcap
xc9[353] carray_top n9 unitcap
xc9[352] carray_top n9 unitcap
xc9[351] carray_top n9 unitcap
xc9[350] carray_top n9 unitcap
xc9[349] carray_top n9 unitcap
xc9[348] carray_top n9 unitcap
xc9[347] carray_top n9 unitcap
xc9[346] carray_top n9 unitcap
xc9[345] carray_top n9 unitcap
xc9[344] carray_top n9 unitcap
xc9[343] carray_top n9 unitcap
xc9[342] carray_top n9 unitcap
xc9[341] carray_top n9 unitcap
xc9[340] carray_top n9 unitcap
xc9[339] carray_top n9 unitcap
xc9[338] carray_top n9 unitcap
xc9[337] carray_top n9 unitcap
xc9[336] carray_top n9 unitcap
xc9[335] carray_top n9 unitcap
xc9[334] carray_top n9 unitcap
xc9[333] carray_top n9 unitcap
xc9[332] carray_top n9 unitcap
xc9[331] carray_top n9 unitcap
xc9[330] carray_top n9 unitcap
xc9[329] carray_top n9 unitcap
xc9[328] carray_top n9 unitcap
xc9[327] carray_top n9 unitcap
xc9[326] carray_top n9 unitcap
xc9[325] carray_top n9 unitcap
xc9[324] carray_top n9 unitcap
xc9[323] carray_top n9 unitcap
xc9[322] carray_top n9 unitcap
xc9[321] carray_top n9 unitcap
xc9[320] carray_top n9 unitcap
xc9[319] carray_top n9 unitcap
xc9[318] carray_top n9 unitcap
xc9[317] carray_top n9 unitcap
xc9[316] carray_top n9 unitcap
xc9[315] carray_top n9 unitcap
xc9[314] carray_top n9 unitcap
xc9[313] carray_top n9 unitcap
xc9[312] carray_top n9 unitcap
xc9[311] carray_top n9 unitcap
xc9[310] carray_top n9 unitcap
xc9[309] carray_top n9 unitcap
xc9[308] carray_top n9 unitcap
xc9[307] carray_top n9 unitcap
xc9[306] carray_top n9 unitcap
xc9[305] carray_top n9 unitcap
xc9[304] carray_top n9 unitcap
xc9[303] carray_top n9 unitcap
xc9[302] carray_top n9 unitcap
xc9[301] carray_top n9 unitcap
xc9[300] carray_top n9 unitcap
xc9[299] carray_top n9 unitcap
xc9[298] carray_top n9 unitcap
xc9[297] carray_top n9 unitcap
xc9[296] carray_top n9 unitcap
xc9[295] carray_top n9 unitcap
xc9[294] carray_top n9 unitcap
xc9[293] carray_top n9 unitcap
xc9[292] carray_top n9 unitcap
xc9[291] carray_top n9 unitcap
xc9[290] carray_top n9 unitcap
xc9[289] carray_top n9 unitcap
xc9[288] carray_top n9 unitcap
xc9[287] carray_top n9 unitcap
xc9[286] carray_top n9 unitcap
xc9[285] carray_top n9 unitcap
xc9[284] carray_top n9 unitcap
xc9[283] carray_top n9 unitcap
xc9[282] carray_top n9 unitcap
xc9[281] carray_top n9 unitcap
xc9[280] carray_top n9 unitcap
xc9[279] carray_top n9 unitcap
xc9[278] carray_top n9 unitcap
xc9[277] carray_top n9 unitcap
xc9[276] carray_top n9 unitcap
xc9[275] carray_top n9 unitcap
xc9[274] carray_top n9 unitcap
xc9[273] carray_top n9 unitcap
xc9[272] carray_top n9 unitcap
xc9[271] carray_top n9 unitcap
xc9[270] carray_top n9 unitcap
xc9[269] carray_top n9 unitcap
xc9[268] carray_top n9 unitcap
xc9[267] carray_top n9 unitcap
xc9[266] carray_top n9 unitcap
xc9[265] carray_top n9 unitcap
xc9[264] carray_top n9 unitcap
xc9[263] carray_top n9 unitcap
xc9[262] carray_top n9 unitcap
xc9[261] carray_top n9 unitcap
xc9[260] carray_top n9 unitcap
xc9[259] carray_top n9 unitcap
xc9[258] carray_top n9 unitcap
xc9[257] carray_top n9 unitcap
xc9[256] carray_top n9 unitcap
xc9[255] carray_top n9 unitcap
xc9[254] carray_top n9 unitcap
xc9[253] carray_top n9 unitcap
xc9[252] carray_top n9 unitcap
xc9[251] carray_top n9 unitcap
xc9[250] carray_top n9 unitcap
xc9[249] carray_top n9 unitcap
xc9[248] carray_top n9 unitcap
xc9[247] carray_top n9 unitcap
xc9[246] carray_top n9 unitcap
xc9[245] carray_top n9 unitcap
xc9[244] carray_top n9 unitcap
xc9[243] carray_top n9 unitcap
xc9[242] carray_top n9 unitcap
xc9[241] carray_top n9 unitcap
xc9[240] carray_top n9 unitcap
xc9[239] carray_top n9 unitcap
xc9[238] carray_top n9 unitcap
xc9[237] carray_top n9 unitcap
xc9[236] carray_top n9 unitcap
xc9[235] carray_top n9 unitcap
xc9[234] carray_top n9 unitcap
xc9[233] carray_top n9 unitcap
xc9[232] carray_top n9 unitcap
xc9[231] carray_top n9 unitcap
xc9[230] carray_top n9 unitcap
xc9[229] carray_top n9 unitcap
xc9[228] carray_top n9 unitcap
xc9[227] carray_top n9 unitcap
xc9[226] carray_top n9 unitcap
xc9[225] carray_top n9 unitcap
xc9[224] carray_top n9 unitcap
xc9[223] carray_top n9 unitcap
xc9[222] carray_top n9 unitcap
xc9[221] carray_top n9 unitcap
xc9[220] carray_top n9 unitcap
xc9[219] carray_top n9 unitcap
xc9[218] carray_top n9 unitcap
xc9[217] carray_top n9 unitcap
xc9[216] carray_top n9 unitcap
xc9[215] carray_top n9 unitcap
xc9[214] carray_top n9 unitcap
xc9[213] carray_top n9 unitcap
xc9[212] carray_top n9 unitcap
xc9[211] carray_top n9 unitcap
xc9[210] carray_top n9 unitcap
xc9[209] carray_top n9 unitcap
xc9[208] carray_top n9 unitcap
xc9[207] carray_top n9 unitcap
xc9[206] carray_top n9 unitcap
xc9[205] carray_top n9 unitcap
xc9[204] carray_top n9 unitcap
xc9[203] carray_top n9 unitcap
xc9[202] carray_top n9 unitcap
xc9[201] carray_top n9 unitcap
xc9[200] carray_top n9 unitcap
xc9[199] carray_top n9 unitcap
xc9[198] carray_top n9 unitcap
xc9[197] carray_top n9 unitcap
xc9[196] carray_top n9 unitcap
xc9[195] carray_top n9 unitcap
xc9[194] carray_top n9 unitcap
xc9[193] carray_top n9 unitcap
xc9[192] carray_top n9 unitcap
xc9[191] carray_top n9 unitcap
xc9[190] carray_top n9 unitcap
xc9[189] carray_top n9 unitcap
xc9[188] carray_top n9 unitcap
xc9[187] carray_top n9 unitcap
xc9[186] carray_top n9 unitcap
xc9[185] carray_top n9 unitcap
xc9[184] carray_top n9 unitcap
xc9[183] carray_top n9 unitcap
xc9[182] carray_top n9 unitcap
xc9[181] carray_top n9 unitcap
xc9[180] carray_top n9 unitcap
xc9[179] carray_top n9 unitcap
xc9[178] carray_top n9 unitcap
xc9[177] carray_top n9 unitcap
xc9[176] carray_top n9 unitcap
xc9[175] carray_top n9 unitcap
xc9[174] carray_top n9 unitcap
xc9[173] carray_top n9 unitcap
xc9[172] carray_top n9 unitcap
xc9[171] carray_top n9 unitcap
xc9[170] carray_top n9 unitcap
xc9[169] carray_top n9 unitcap
xc9[168] carray_top n9 unitcap
xc9[167] carray_top n9 unitcap
xc9[166] carray_top n9 unitcap
xc9[165] carray_top n9 unitcap
xc9[164] carray_top n9 unitcap
xc9[163] carray_top n9 unitcap
xc9[162] carray_top n9 unitcap
xc9[161] carray_top n9 unitcap
xc9[160] carray_top n9 unitcap
xc9[159] carray_top n9 unitcap
xc9[158] carray_top n9 unitcap
xc9[157] carray_top n9 unitcap
xc9[156] carray_top n9 unitcap
xc9[155] carray_top n9 unitcap
xc9[154] carray_top n9 unitcap
xc9[153] carray_top n9 unitcap
xc9[152] carray_top n9 unitcap
xc9[151] carray_top n9 unitcap
xc9[150] carray_top n9 unitcap
xc9[149] carray_top n9 unitcap
xc9[148] carray_top n9 unitcap
xc9[147] carray_top n9 unitcap
xc9[146] carray_top n9 unitcap
xc9[145] carray_top n9 unitcap
xc9[144] carray_top n9 unitcap
xc9[143] carray_top n9 unitcap
xc9[142] carray_top n9 unitcap
xc9[141] carray_top n9 unitcap
xc9[140] carray_top n9 unitcap
xc9[139] carray_top n9 unitcap
xc9[138] carray_top n9 unitcap
xc9[137] carray_top n9 unitcap
xc9[136] carray_top n9 unitcap
xc9[135] carray_top n9 unitcap
xc9[134] carray_top n9 unitcap
xc9[133] carray_top n9 unitcap
xc9[132] carray_top n9 unitcap
xc9[131] carray_top n9 unitcap
xc9[130] carray_top n9 unitcap
xc9[129] carray_top n9 unitcap
xc9[128] carray_top n9 unitcap
xc9[127] carray_top n9 unitcap
xc9[126] carray_top n9 unitcap
xc9[125] carray_top n9 unitcap
xc9[124] carray_top n9 unitcap
xc9[123] carray_top n9 unitcap
xc9[122] carray_top n9 unitcap
xc9[121] carray_top n9 unitcap
xc9[120] carray_top n9 unitcap
xc9[119] carray_top n9 unitcap
xc9[118] carray_top n9 unitcap
xc9[117] carray_top n9 unitcap
xc9[116] carray_top n9 unitcap
xc9[115] carray_top n9 unitcap
xc9[114] carray_top n9 unitcap
xc9[113] carray_top n9 unitcap
xc9[112] carray_top n9 unitcap
xc9[111] carray_top n9 unitcap
xc9[110] carray_top n9 unitcap
xc9[109] carray_top n9 unitcap
xc9[108] carray_top n9 unitcap
xc9[107] carray_top n9 unitcap
xc9[106] carray_top n9 unitcap
xc9[105] carray_top n9 unitcap
xc9[104] carray_top n9 unitcap
xc9[103] carray_top n9 unitcap
xc9[102] carray_top n9 unitcap
xc9[101] carray_top n9 unitcap
xc9[100] carray_top n9 unitcap
xc9[99] carray_top n9 unitcap
xc9[98] carray_top n9 unitcap
xc9[97] carray_top n9 unitcap
xc9[96] carray_top n9 unitcap
xc9[95] carray_top n9 unitcap
xc9[94] carray_top n9 unitcap
xc9[93] carray_top n9 unitcap
xc9[92] carray_top n9 unitcap
xc9[91] carray_top n9 unitcap
xc9[90] carray_top n9 unitcap
xc9[89] carray_top n9 unitcap
xc9[88] carray_top n9 unitcap
xc9[87] carray_top n9 unitcap
xc9[86] carray_top n9 unitcap
xc9[85] carray_top n9 unitcap
xc9[84] carray_top n9 unitcap
xc9[83] carray_top n9 unitcap
xc9[82] carray_top n9 unitcap
xc9[81] carray_top n9 unitcap
xc9[80] carray_top n9 unitcap
xc9[79] carray_top n9 unitcap
xc9[78] carray_top n9 unitcap
xc9[77] carray_top n9 unitcap
xc9[76] carray_top n9 unitcap
xc9[75] carray_top n9 unitcap
xc9[74] carray_top n9 unitcap
xc9[73] carray_top n9 unitcap
xc9[72] carray_top n9 unitcap
xc9[71] carray_top n9 unitcap
xc9[70] carray_top n9 unitcap
xc9[69] carray_top n9 unitcap
xc9[68] carray_top n9 unitcap
xc9[67] carray_top n9 unitcap
xc9[66] carray_top n9 unitcap
xc9[65] carray_top n9 unitcap
xc9[64] carray_top n9 unitcap
xc9[63] carray_top n9 unitcap
xc9[62] carray_top n9 unitcap
xc9[61] carray_top n9 unitcap
xc9[60] carray_top n9 unitcap
xc9[59] carray_top n9 unitcap
xc9[58] carray_top n9 unitcap
xc9[57] carray_top n9 unitcap
xc9[56] carray_top n9 unitcap
xc9[55] carray_top n9 unitcap
xc9[54] carray_top n9 unitcap
xc9[53] carray_top n9 unitcap
xc9[52] carray_top n9 unitcap
xc9[51] carray_top n9 unitcap
xc9[50] carray_top n9 unitcap
xc9[49] carray_top n9 unitcap
xc9[48] carray_top n9 unitcap
xc9[47] carray_top n9 unitcap
xc9[46] carray_top n9 unitcap
xc9[45] carray_top n9 unitcap
xc9[44] carray_top n9 unitcap
xc9[43] carray_top n9 unitcap
xc9[42] carray_top n9 unitcap
xc9[41] carray_top n9 unitcap
xc9[40] carray_top n9 unitcap
xc9[39] carray_top n9 unitcap
xc9[38] carray_top n9 unitcap
xc9[37] carray_top n9 unitcap
xc9[36] carray_top n9 unitcap
xc9[35] carray_top n9 unitcap
xc9[34] carray_top n9 unitcap
xc9[33] carray_top n9 unitcap
xc9[32] carray_top n9 unitcap
xc9[31] carray_top n9 unitcap
xc9[30] carray_top n9 unitcap
xc9[29] carray_top n9 unitcap
xc9[28] carray_top n9 unitcap
xc9[27] carray_top n9 unitcap
xc9[26] carray_top n9 unitcap
xc9[25] carray_top n9 unitcap
xc9[24] carray_top n9 unitcap
xc9[23] carray_top n9 unitcap
xc9[22] carray_top n9 unitcap
xc9[21] carray_top n9 unitcap
xc9[20] carray_top n9 unitcap
xc9[19] carray_top n9 unitcap
xc9[18] carray_top n9 unitcap
xc9[17] carray_top n9 unitcap
xc9[16] carray_top n9 unitcap
xc9[15] carray_top n9 unitcap
xc9[14] carray_top n9 unitcap
xc9[13] carray_top n9 unitcap
xc9[12] carray_top n9 unitcap
xc9[11] carray_top n9 unitcap
xc9[10] carray_top n9 unitcap
xc9[9] carray_top n9 unitcap
xc9[8] carray_top n9 unitcap
xc9[7] carray_top n9 unitcap
xc9[6] carray_top n9 unitcap
xc9[5] carray_top n9 unitcap
xc9[4] carray_top n9 unitcap
xc9[3] carray_top n9 unitcap
xc9[2] carray_top n9 unitcap
xc9[1] carray_top n9 unitcap
xc9[0] carray_top n9 unitcap
**.ends

* expanding   symbol:  sar_10b/unitcap/unitcap.sym # of pins=2
** sym_path: /home/oe23ranan/gf_analog/xschem/sar_10b/unitcap/unitcap.sym
** sch_path: /home/oe23ranan/gf_analog/xschem/sar_10b/unitcap/unitcap.sch
.subckt unitcap cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2.6f m=1
.ends

.end
