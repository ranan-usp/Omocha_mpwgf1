module saradc(
	inout vdd,
	inout vss,
	input [9:0] user_input,
	input cal,
	input en,
	input clk,
	input rstn,
	output valid,
	output [9:0] result
);
endmodule