* NGSPICE file created from latch.ext - technology: gf180mcuD

.subckt XM2_latch_x4 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G S 0.143803f
C1 D G 0.001764f
C2 D S 0.09188f
C3 D VSUBS 0.04225f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.56551f
.ends

.subckt XM1_latch_x4 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134096f
C2 G S 0.226575f
.ends

.subckt x4_latch in out XM2_latch_x4_0/S VSUBS
XXM2_latch_x4_0 in out XM2_latch_x4_0/S VSUBS XM2_latch_x4
XXM1_latch_x4_0 in out VSUBS XM1_latch_x4
C0 in XM2_latch_x4_0/S 0.039699f
C1 out in 0.057341f
C2 out XM2_latch_x4_0/S 0.102755f
C3 out VSUBS 0.49906f
C4 in VSUBS 0.450066f
C5 XM2_latch_x4_0/S VSUBS 1.7619f
.ends

.subckt XM2_latch_x3 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 S D 0.09188f
C2 S G 0.143803f
C3 D VSUBS 0.04225f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.56551f
.ends

.subckt XM1_latch_x3 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.226575f
.ends

.subckt x3_latch in out XM2_latch_x3_0/S VSUBS
XXM2_latch_x3_0 in out XM2_latch_x3_0/S VSUBS XM2_latch_x3
XXM1_latch_x3_0 in out VSUBS XM1_latch_x3
C0 in out 0.057341f
C1 XM2_latch_x3_0/S out 0.102755f
C2 XM2_latch_x3_0/S in 0.039699f
C3 out VSUBS 0.49906f
C4 in VSUBS 0.450066f
C5 XM2_latch_x3_0/S VSUBS 1.761853f
.ends

.subckt XM4_latch G D a_258_n1293# S
X0 S G D S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt XM2_latch_x2 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 S G 0.143685f
C2 S D 0.091354f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.5328f
.ends

.subckt XM1_latch_x2 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt x2_latch in out XM2_latch_x2_0/S VSUBS
XXM2_latch_x2_0 in out XM2_latch_x2_0/S VSUBS XM2_latch_x2
XXM1_latch_x2_0 in out VSUBS XM1_latch_x2
C0 out in 0.057341f
C1 XM2_latch_x2_0/S in 0.039609f
C2 XM2_latch_x2_0/S out 0.088354f
C3 out VSUBS 0.511014f
C4 in VSUBS 0.449897f
C5 XM2_latch_x2_0/S VSUBS 1.73873f
.ends

.subckt XM3_latch G D a_n349_n1268# S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt XM2_latch_x1 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S G 0.143685f
C1 S D 0.091354f
C2 D G 0.001764f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.5328f
.ends

.subckt XM1_latch_x1 G D S a_n254_114#
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt x1_latch in out XM1_latch_x1_0/a_n254_114# XM2_latch_x1_0/S VSUBS
XXM2_latch_x1_0 in out XM2_latch_x1_0/S VSUBS XM2_latch_x1
XXM1_latch_x1_0 in out VSUBS XM1_latch_x1_0/a_n254_114# XM1_latch_x1
C0 XM2_latch_x1_0/S in 0.039609f
C1 XM2_latch_x1_0/S out 0.088354f
C2 out in 0.057341f
C3 out VSUBS 0.511014f
C4 in VSUBS 0.449897f
C5 XM2_latch_x1_0/S VSUBS 1.738608f
.ends

.subckt latch tutyuu1 tutyuu2 Qn Q S R vss vdd
Xx4_latch_0 S tutyuu1 vdd vss x4_latch
Xx3_latch_0 R tutyuu2 vdd vss x3_latch
XXM4_latch_0 tutyuu2 Q vss vss XM4_latch
Xx2_latch_0 Q Qn vdd vss x2_latch
XXM3_latch_0 tutyuu1 Qn vss vss XM3_latch
Xx1_latch_0 Qn Q vss vdd vss x1_latch
C0 tutyuu2 Q 0.109341f
C1 tutyuu1 Q 0.060871f
C2 vdd R 0.053607f
C3 Qn tutyuu2 0.060761f
C4 tutyuu1 Qn 0.109231f
C5 tutyuu1 S 0.115854f
C6 Qn Q 1.472762f
C7 vdd tutyuu2 0.101384f
C8 tutyuu1 vdd 0.101448f
C9 vdd Q 0.35434f
C10 S Qn 0.011276f
C11 Qn vdd 0.059024f
C12 S vdd 0.053607f
C13 tutyuu2 R 0.115854f
C14 R Q 0.011346f
C15 vdd vss 5.959083f
C16 Qn vss 0.913293f
C17 Q vss 0.942836f
C18 tutyuu2 vss 0.702253f
C19 R vss 0.476811f
C20 tutyuu1 vss 0.702189f
C21 S vss 0.476811f
.ends

