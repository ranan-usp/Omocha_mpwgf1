VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sarlogic
  CLASS BLOCK ;
  FOREIGN sarlogic ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 130.000 ;
  PIN cal
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 29.120 180.000 29.680 ;
    END
  END cal
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 13.440 180.000 14.000 ;
    END
  END clk
  PIN clkc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END clkc
  PIN comp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 4.000 70.000 ;
    END
  END comp
  PIN ctln[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 0.000 9.520 4.000 ;
    END
  END ctln[0]
  PIN ctln[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 4.000 ;
    END
  END ctln[1]
  PIN ctln[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END ctln[2]
  PIN ctln[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END ctln[3]
  PIN ctln[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END ctln[4]
  PIN ctln[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END ctln[5]
  PIN ctln[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END ctln[6]
  PIN ctln[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END ctln[7]
  PIN ctln[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END ctln[8]
  PIN ctln[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END ctln[9]
  PIN ctlp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 126.000 9.520 130.000 ;
    END
  END ctlp[0]
  PIN ctlp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 126.000 170.800 130.000 ;
    END
  END ctlp[1]
  PIN ctlp[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 126.000 152.880 130.000 ;
    END
  END ctlp[2]
  PIN ctlp[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 126.000 134.960 130.000 ;
    END
  END ctlp[3]
  PIN ctlp[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 126.000 117.040 130.000 ;
    END
  END ctlp[4]
  PIN ctlp[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 126.000 99.120 130.000 ;
    END
  END ctlp[5]
  PIN ctlp[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 126.000 81.200 130.000 ;
    END
  END ctlp[6]
  PIN ctlp[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 126.000 63.280 130.000 ;
    END
  END ctlp[7]
  PIN ctlp[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 126.000 45.360 130.000 ;
    END
  END ctlp[8]
  PIN ctlp[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 126.000 27.440 130.000 ;
    END
  END ctlp[9]
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 21.280 180.000 21.840 ;
    END
  END en
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 52.640 180.000 53.200 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 60.480 180.000 61.040 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 68.320 180.000 68.880 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 76.160 180.000 76.720 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 84.000 180.000 84.560 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 91.840 180.000 92.400 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 99.680 180.000 100.240 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 107.520 180.000 108.080 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 115.360 180.000 115.920 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 123.200 180.000 123.760 ;
    END
  END result[9]
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 5.600 180.000 6.160 ;
    END
  END rstn
  PIN sample
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 44.800 180.000 45.360 ;
    END
  END sample
  PIN trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END trim[0]
  PIN trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END trim[1]
  PIN trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END trim[2]
  PIN trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.960 4.000 9.520 ;
    END
  END trim[3]
  PIN trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.280 4.000 49.840 ;
    END
  END trim[4]
  PIN trimb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END trimb[0]
  PIN trimb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.600 4.000 90.160 ;
    END
  END trimb[1]
  PIN trimb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 4.000 110.320 ;
    END
  END trimb[2]
  PIN trimb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 4.000 120.400 ;
    END
  END trimb[3]
  PIN trimb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 4.000 80.080 ;
    END
  END trimb[4]
  PIN valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 176.000 36.960 180.000 37.520 ;
    END
  END valid
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 26.710 15.380 28.310 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.290 15.380 69.890 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.870 15.380 111.470 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.450 15.380 153.050 113.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 47.500 15.380 49.100 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 89.080 15.380 90.680 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 130.660 15.380 132.260 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.240 15.380 173.840 113.980 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 173.840 113.980 ;
      LAYER Metal2 ;
        RECT 8.540 125.700 8.660 126.420 ;
        RECT 9.820 125.700 26.580 126.420 ;
        RECT 27.740 125.700 44.500 126.420 ;
        RECT 45.660 125.700 62.420 126.420 ;
        RECT 63.580 125.700 80.340 126.420 ;
        RECT 81.500 125.700 98.260 126.420 ;
        RECT 99.420 125.700 116.180 126.420 ;
        RECT 117.340 125.700 134.100 126.420 ;
        RECT 135.260 125.700 152.020 126.420 ;
        RECT 153.180 125.700 169.940 126.420 ;
        RECT 171.100 125.700 173.700 126.420 ;
        RECT 8.540 4.300 173.700 125.700 ;
        RECT 8.540 3.500 8.660 4.300 ;
        RECT 9.820 3.500 26.580 4.300 ;
        RECT 27.740 3.500 44.500 4.300 ;
        RECT 45.660 3.500 62.420 4.300 ;
        RECT 63.580 3.500 80.340 4.300 ;
        RECT 81.500 3.500 98.260 4.300 ;
        RECT 99.420 3.500 116.180 4.300 ;
        RECT 117.340 3.500 134.100 4.300 ;
        RECT 135.260 3.500 152.020 4.300 ;
        RECT 153.180 3.500 169.940 4.300 ;
        RECT 171.100 3.500 173.700 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 122.900 175.700 123.620 ;
        RECT 4.000 120.700 176.000 122.900 ;
        RECT 4.300 119.540 176.000 120.700 ;
        RECT 4.000 116.220 176.000 119.540 ;
        RECT 4.000 115.060 175.700 116.220 ;
        RECT 4.000 110.620 176.000 115.060 ;
        RECT 4.300 109.460 176.000 110.620 ;
        RECT 4.000 108.380 176.000 109.460 ;
        RECT 4.000 107.220 175.700 108.380 ;
        RECT 4.000 100.540 176.000 107.220 ;
        RECT 4.300 99.380 175.700 100.540 ;
        RECT 4.000 92.700 176.000 99.380 ;
        RECT 4.000 91.540 175.700 92.700 ;
        RECT 4.000 90.460 176.000 91.540 ;
        RECT 4.300 89.300 176.000 90.460 ;
        RECT 4.000 84.860 176.000 89.300 ;
        RECT 4.000 83.700 175.700 84.860 ;
        RECT 4.000 80.380 176.000 83.700 ;
        RECT 4.300 79.220 176.000 80.380 ;
        RECT 4.000 77.020 176.000 79.220 ;
        RECT 4.000 75.860 175.700 77.020 ;
        RECT 4.000 70.300 176.000 75.860 ;
        RECT 4.300 69.180 176.000 70.300 ;
        RECT 4.300 69.140 175.700 69.180 ;
        RECT 4.000 68.020 175.700 69.140 ;
        RECT 4.000 61.340 176.000 68.020 ;
        RECT 4.000 60.220 175.700 61.340 ;
        RECT 4.300 60.180 175.700 60.220 ;
        RECT 4.300 59.060 176.000 60.180 ;
        RECT 4.000 53.500 176.000 59.060 ;
        RECT 4.000 52.340 175.700 53.500 ;
        RECT 4.000 50.140 176.000 52.340 ;
        RECT 4.300 48.980 176.000 50.140 ;
        RECT 4.000 45.660 176.000 48.980 ;
        RECT 4.000 44.500 175.700 45.660 ;
        RECT 4.000 40.060 176.000 44.500 ;
        RECT 4.300 38.900 176.000 40.060 ;
        RECT 4.000 37.820 176.000 38.900 ;
        RECT 4.000 36.660 175.700 37.820 ;
        RECT 4.000 29.980 176.000 36.660 ;
        RECT 4.300 28.820 175.700 29.980 ;
        RECT 4.000 22.140 176.000 28.820 ;
        RECT 4.000 20.980 175.700 22.140 ;
        RECT 4.000 19.900 176.000 20.980 ;
        RECT 4.300 18.740 176.000 19.900 ;
        RECT 4.000 14.300 176.000 18.740 ;
        RECT 4.000 13.140 175.700 14.300 ;
        RECT 4.000 9.820 176.000 13.140 ;
        RECT 4.300 8.660 176.000 9.820 ;
        RECT 4.000 6.460 176.000 8.660 ;
        RECT 4.000 5.740 175.700 6.460 ;
      LAYER Metal4 ;
        RECT 96.460 47.690 100.660 65.990 ;
  END
END sarlogic
END LIBRARY

