* NGSPICE file created from carray.ext - technology: gf180mcuD

.subckt carray n9 n0 n8 n7 n6 n5 n4 n3 n2 n1 ndum carray_out
C0 n3 n7 0.891504f
C1 n5 n4 27.491999f
C2 n3 n1 0.137399f
C3 n2 n8 0.770114f
C4 n5 n9 7.399346f
C5 n6 n7 34.326103f
C6 n5 carray_out 52.565514f
C7 n1 n6 0.134562f
C8 n4 n8 2.84323f
C9 n9 n8 87.10268f
C10 n3 n2 22.8406f
C11 n8 carray_out 0.420151p
C12 n6 n2 0.207877f
C13 n3 n4 25.8929f
C14 n3 n9 1.911224f
C15 n3 carray_out 13.201303f
C16 n6 n4 0.614078f
C17 n1 n7 0.205173f
C18 n9 n6 14.716789f
C19 n5 n8 5.60732f
C20 n6 carray_out 0.105055p
C21 n7 n2 0.485242f
C22 n0 n1 8.469266f
C23 n3 n5 0.346757f
C24 n1 n2 16.597801f
C25 n7 n4 1.70387f
C26 n9 n7 29.516087f
C27 n5 n6 28.589401f
C28 n3 n8 1.46111f
C29 n1 n4 0.134826f
C30 n1 n9 0.342393f
C31 n7 carray_out 0.210031p
C32 n1 carray_out 3.365891f
C33 n6 n8 11.2161f
C34 n1 ndum 8.161697f
C35 n0 n9 0.184985f
C36 n4 n2 0.213096f
C37 n9 n2 0.996568f
C38 n0 carray_out 1.684219f
C39 n2 carray_out 6.640605f
C40 n3 n6 0.336612f
C41 n5 n7 3.36878f
C42 n9 n4 3.740573f
C43 n5 n1 0.134705f
C44 n4 carray_out 26.32268f
C45 n9 carray_out 0.846153p
C46 n7 n8 50.178104f
C47 n9 ndum 0.127951f
C48 n1 n8 0.278221f
C49 ndum carray_out 1.640173f
C50 n5 n2 0.207999f
C51 n4 VSUBS 42.229664f
C52 ndum VSUBS 13.717415f
C53 n5 VSUBS 53.39593f
C54 n9 VSUBS 0.118604p
C55 carray_out VSUBS 0.118526p
C56 n8 VSUBS 90.036354f
C57 n7 VSUBS 82.1809f
C58 n6 VSUBS 66.84599f
C59 n0 VSUBS 16.513115f
C60 n2 VSUBS 30.672361f
C61 n1 VSUBS 17.314531f
C62 n3 VSUBS 34.940525f
.ends

