magic
tech gf180mcuD
magscale 1 5
timestamp 1702006702
<< metal1 >>
rect 672 8245 9296 8262
rect 672 8219 1685 8245
rect 1711 8219 1737 8245
rect 1763 8219 1789 8245
rect 1815 8219 3841 8245
rect 3867 8219 3893 8245
rect 3919 8219 3945 8245
rect 3971 8219 5997 8245
rect 6023 8219 6049 8245
rect 6075 8219 6101 8245
rect 6127 8219 8153 8245
rect 8179 8219 8205 8245
rect 8231 8219 8257 8245
rect 8283 8219 9296 8245
rect 672 8202 9296 8219
rect 5783 8161 5809 8167
rect 7457 8135 7463 8161
rect 7489 8135 7495 8161
rect 5783 8129 5809 8135
rect 855 8049 881 8055
rect 855 8017 881 8023
rect 1191 8049 1217 8055
rect 1191 8017 1217 8023
rect 1583 8049 1609 8055
rect 6281 8023 6287 8049
rect 6313 8023 6319 8049
rect 7961 8023 7967 8049
rect 7993 8023 7999 8049
rect 8577 8023 8583 8049
rect 8609 8023 8615 8049
rect 8913 8023 8919 8049
rect 8945 8023 8951 8049
rect 1583 8017 1609 8023
rect 8807 7993 8833 7999
rect 8807 7961 8833 7967
rect 1023 7937 1049 7943
rect 1023 7905 1049 7911
rect 1359 7937 1385 7943
rect 1359 7905 1385 7911
rect 8471 7937 8497 7943
rect 8471 7905 8497 7911
rect 672 7853 9376 7870
rect 672 7827 2763 7853
rect 2789 7827 2815 7853
rect 2841 7827 2867 7853
rect 2893 7827 4919 7853
rect 4945 7827 4971 7853
rect 4997 7827 5023 7853
rect 5049 7827 7075 7853
rect 7101 7827 7127 7853
rect 7153 7827 7179 7853
rect 7205 7827 9231 7853
rect 9257 7827 9283 7853
rect 9309 7827 9335 7853
rect 9361 7827 9376 7853
rect 672 7810 9376 7827
rect 1079 7769 1105 7775
rect 1079 7737 1105 7743
rect 6455 7769 6481 7775
rect 6455 7737 6481 7743
rect 8695 7713 8721 7719
rect 8695 7681 8721 7687
rect 9087 7713 9113 7719
rect 9087 7681 9113 7687
rect 6953 7631 6959 7657
rect 6985 7631 6991 7657
rect 8409 7631 8415 7657
rect 8441 7631 8447 7657
rect 8801 7631 8807 7657
rect 8833 7631 8839 7657
rect 7911 7601 7937 7607
rect 7911 7569 7937 7575
rect 9031 7545 9057 7551
rect 9031 7513 9057 7519
rect 672 7461 9296 7478
rect 672 7435 1685 7461
rect 1711 7435 1737 7461
rect 1763 7435 1789 7461
rect 1815 7435 3841 7461
rect 3867 7435 3893 7461
rect 3919 7435 3945 7461
rect 3971 7435 5997 7461
rect 6023 7435 6049 7461
rect 6075 7435 6101 7461
rect 6127 7435 8153 7461
rect 8179 7435 8205 7461
rect 8231 7435 8257 7461
rect 8283 7435 9296 7461
rect 672 7418 9296 7435
rect 7631 7265 7657 7271
rect 8913 7239 8919 7265
rect 8945 7239 8951 7265
rect 7631 7233 7657 7239
rect 855 7209 881 7215
rect 855 7177 881 7183
rect 1023 7209 1049 7215
rect 1023 7177 1049 7183
rect 1247 7209 1273 7215
rect 1247 7177 1273 7183
rect 7575 7153 7601 7159
rect 7575 7121 7601 7127
rect 8583 7153 8609 7159
rect 8583 7121 8609 7127
rect 672 7069 9376 7086
rect 672 7043 2763 7069
rect 2789 7043 2815 7069
rect 2841 7043 2867 7069
rect 2893 7043 4919 7069
rect 4945 7043 4971 7069
rect 4997 7043 5023 7069
rect 5049 7043 7075 7069
rect 7101 7043 7127 7069
rect 7153 7043 7179 7069
rect 7205 7043 9231 7069
rect 9257 7043 9283 7069
rect 9309 7043 9335 7069
rect 9361 7043 9376 7069
rect 672 7026 9376 7043
rect 8695 6985 8721 6991
rect 8695 6953 8721 6959
rect 9087 6929 9113 6935
rect 9087 6897 9113 6903
rect 8353 6847 8359 6873
rect 8385 6847 8391 6873
rect 8801 6847 8807 6873
rect 8833 6847 8839 6873
rect 7793 6791 7799 6817
rect 7825 6791 7831 6817
rect 9031 6761 9057 6767
rect 9031 6729 9057 6735
rect 672 6677 9296 6694
rect 672 6651 1685 6677
rect 1711 6651 1737 6677
rect 1763 6651 1789 6677
rect 1815 6651 3841 6677
rect 3867 6651 3893 6677
rect 3919 6651 3945 6677
rect 3971 6651 5997 6677
rect 6023 6651 6049 6677
rect 6075 6651 6101 6677
rect 6127 6651 8153 6677
rect 8179 6651 8205 6677
rect 8231 6651 8257 6677
rect 8283 6651 9296 6677
rect 672 6634 9296 6651
rect 8583 6537 8609 6543
rect 8583 6505 8609 6511
rect 8857 6455 8863 6481
rect 8889 6455 8895 6481
rect 855 6425 881 6431
rect 855 6393 881 6399
rect 1023 6425 1049 6431
rect 1023 6393 1049 6399
rect 1247 6369 1273 6375
rect 1247 6337 1273 6343
rect 672 6285 9376 6302
rect 672 6259 2763 6285
rect 2789 6259 2815 6285
rect 2841 6259 2867 6285
rect 2893 6259 4919 6285
rect 4945 6259 4971 6285
rect 4997 6259 5023 6285
rect 5049 6259 7075 6285
rect 7101 6259 7127 6285
rect 7153 6259 7179 6285
rect 7205 6259 9231 6285
rect 9257 6259 9283 6285
rect 9309 6259 9335 6285
rect 9361 6259 9376 6285
rect 672 6242 9376 6259
rect 8751 6145 8777 6151
rect 8751 6113 8777 6119
rect 9031 6033 9057 6039
rect 9031 6001 9057 6007
rect 8695 5977 8721 5983
rect 8695 5945 8721 5951
rect 672 5893 9296 5910
rect 672 5867 1685 5893
rect 1711 5867 1737 5893
rect 1763 5867 1789 5893
rect 1815 5867 3841 5893
rect 3867 5867 3893 5893
rect 3919 5867 3945 5893
rect 3971 5867 5997 5893
rect 6023 5867 6049 5893
rect 6075 5867 6101 5893
rect 6127 5867 8153 5893
rect 8179 5867 8205 5893
rect 8231 5867 8257 5893
rect 8283 5867 9296 5893
rect 672 5850 9296 5867
rect 8975 5809 9001 5815
rect 8975 5777 9001 5783
rect 7793 5671 7799 5697
rect 7825 5671 7831 5697
rect 855 5641 881 5647
rect 855 5609 881 5615
rect 1023 5641 1049 5647
rect 1023 5609 1049 5615
rect 1247 5585 1273 5591
rect 1247 5553 1273 5559
rect 672 5501 9376 5518
rect 672 5475 2763 5501
rect 2789 5475 2815 5501
rect 2841 5475 2867 5501
rect 2893 5475 4919 5501
rect 4945 5475 4971 5501
rect 4997 5475 5023 5501
rect 5049 5475 7075 5501
rect 7101 5475 7127 5501
rect 7153 5475 7179 5501
rect 7205 5475 9231 5501
rect 9257 5475 9283 5501
rect 9309 5475 9335 5501
rect 9361 5475 9376 5501
rect 672 5458 9376 5475
rect 8863 5417 8889 5423
rect 8863 5385 8889 5391
rect 8695 5361 8721 5367
rect 8695 5329 8721 5335
rect 9087 5361 9113 5367
rect 9087 5329 9113 5335
rect 7345 5279 7351 5305
rect 7377 5279 7383 5305
rect 8303 5193 8329 5199
rect 8303 5161 8329 5167
rect 672 5109 9296 5126
rect 672 5083 1685 5109
rect 1711 5083 1737 5109
rect 1763 5083 1789 5109
rect 1815 5083 3841 5109
rect 3867 5083 3893 5109
rect 3919 5083 3945 5109
rect 3971 5083 5997 5109
rect 6023 5083 6049 5109
rect 6075 5083 6101 5109
rect 6127 5083 8153 5109
rect 8179 5083 8205 5109
rect 8231 5083 8257 5109
rect 8283 5083 9296 5109
rect 672 5066 9296 5083
rect 8583 5025 8609 5031
rect 8583 4993 8609 4999
rect 7569 4887 7575 4913
rect 7601 4887 7607 4913
rect 8857 4887 8863 4913
rect 8889 4887 8895 4913
rect 855 4857 881 4863
rect 855 4825 881 4831
rect 1247 4857 1273 4863
rect 1247 4825 1273 4831
rect 7463 4857 7489 4863
rect 7463 4825 7489 4831
rect 1023 4801 1049 4807
rect 1023 4769 1049 4775
rect 7351 4801 7377 4807
rect 7351 4769 7377 4775
rect 672 4717 9376 4734
rect 672 4691 2763 4717
rect 2789 4691 2815 4717
rect 2841 4691 2867 4717
rect 2893 4691 4919 4717
rect 4945 4691 4971 4717
rect 4997 4691 5023 4717
rect 5049 4691 7075 4717
rect 7101 4691 7127 4717
rect 7153 4691 7179 4717
rect 7205 4691 9231 4717
rect 9257 4691 9283 4717
rect 9309 4691 9335 4717
rect 9361 4691 9376 4717
rect 672 4674 9376 4691
rect 6959 4633 6985 4639
rect 6959 4601 6985 4607
rect 8695 4633 8721 4639
rect 8695 4601 8721 4607
rect 8863 4577 8889 4583
rect 8863 4545 8889 4551
rect 9087 4577 9113 4583
rect 9087 4545 9113 4551
rect 7233 4495 7239 4521
rect 7265 4495 7271 4521
rect 8303 4409 8329 4415
rect 8303 4377 8329 4383
rect 9031 4409 9057 4415
rect 9031 4377 9057 4383
rect 672 4325 9296 4342
rect 672 4299 1685 4325
rect 1711 4299 1737 4325
rect 1763 4299 1789 4325
rect 1815 4299 3841 4325
rect 3867 4299 3893 4325
rect 3919 4299 3945 4325
rect 3971 4299 5997 4325
rect 6023 4299 6049 4325
rect 6075 4299 6101 4325
rect 6127 4299 8153 4325
rect 8179 4299 8205 4325
rect 8231 4299 8257 4325
rect 8283 4299 9296 4325
rect 672 4282 9296 4299
rect 7239 4241 7265 4247
rect 7239 4209 7265 4215
rect 8583 4241 8609 4247
rect 8583 4209 8609 4215
rect 9025 4103 9031 4129
rect 9057 4103 9063 4129
rect 7295 4073 7321 4079
rect 7295 4041 7321 4047
rect 7463 4073 7489 4079
rect 7463 4041 7489 4047
rect 7631 4073 7657 4079
rect 7631 4041 7657 4047
rect 7127 4017 7153 4023
rect 7127 3985 7153 3991
rect 672 3933 9376 3950
rect 672 3907 2763 3933
rect 2789 3907 2815 3933
rect 2841 3907 2867 3933
rect 2893 3907 4919 3933
rect 4945 3907 4971 3933
rect 4997 3907 5023 3933
rect 5049 3907 7075 3933
rect 7101 3907 7127 3933
rect 7153 3907 7179 3933
rect 7205 3907 9231 3933
rect 9257 3907 9283 3933
rect 9309 3907 9335 3933
rect 9361 3907 9376 3933
rect 672 3890 9376 3907
rect 8695 3849 8721 3855
rect 8695 3817 8721 3823
rect 9031 3849 9057 3855
rect 9031 3817 9057 3823
rect 1023 3793 1049 3799
rect 1023 3761 1049 3767
rect 855 3737 881 3743
rect 8353 3711 8359 3737
rect 8385 3711 8391 3737
rect 8801 3711 8807 3737
rect 8833 3711 8839 3737
rect 855 3705 881 3711
rect 1247 3681 1273 3687
rect 1247 3649 1273 3655
rect 9087 3681 9113 3687
rect 9087 3649 9113 3655
rect 7911 3625 7937 3631
rect 7911 3593 7937 3599
rect 672 3541 9296 3558
rect 672 3515 1685 3541
rect 1711 3515 1737 3541
rect 1763 3515 1789 3541
rect 1815 3515 3841 3541
rect 3867 3515 3893 3541
rect 3919 3515 3945 3541
rect 3971 3515 5997 3541
rect 6023 3515 6049 3541
rect 6075 3515 6101 3541
rect 6127 3515 8153 3541
rect 8179 3515 8205 3541
rect 8231 3515 8257 3541
rect 8283 3515 9296 3541
rect 672 3498 9296 3515
rect 8583 3457 8609 3463
rect 8583 3425 8609 3431
rect 8969 3319 8975 3345
rect 9001 3319 9007 3345
rect 7631 3233 7657 3239
rect 7631 3201 7657 3207
rect 672 3149 9376 3166
rect 672 3123 2763 3149
rect 2789 3123 2815 3149
rect 2841 3123 2867 3149
rect 2893 3123 4919 3149
rect 4945 3123 4971 3149
rect 4997 3123 5023 3149
rect 5049 3123 7075 3149
rect 7101 3123 7127 3149
rect 7153 3123 7179 3149
rect 7205 3123 9231 3149
rect 9257 3123 9283 3149
rect 9309 3123 9335 3149
rect 9361 3123 9376 3149
rect 672 3106 9376 3123
rect 1023 3065 1049 3071
rect 1023 3033 1049 3039
rect 8695 3065 8721 3071
rect 8695 3033 8721 3039
rect 8975 3065 9001 3071
rect 8975 3033 9001 3039
rect 8751 3009 8777 3015
rect 8751 2977 8777 2983
rect 8919 3009 8945 3015
rect 8919 2977 8945 2983
rect 855 2953 881 2959
rect 7345 2927 7351 2953
rect 7377 2927 7383 2953
rect 855 2921 881 2927
rect 1247 2897 1273 2903
rect 1247 2865 1273 2871
rect 7631 2841 7657 2847
rect 7631 2809 7657 2815
rect 672 2757 9296 2774
rect 672 2731 1685 2757
rect 1711 2731 1737 2757
rect 1763 2731 1789 2757
rect 1815 2731 3841 2757
rect 3867 2731 3893 2757
rect 3919 2731 3945 2757
rect 3971 2731 5997 2757
rect 6023 2731 6049 2757
rect 6075 2731 6101 2757
rect 6127 2731 8153 2757
rect 8179 2731 8205 2757
rect 8231 2731 8257 2757
rect 8283 2731 9296 2757
rect 672 2714 9296 2731
rect 8353 2647 8359 2673
rect 8385 2647 8391 2673
rect 7687 2617 7713 2623
rect 7687 2585 7713 2591
rect 8969 2535 8975 2561
rect 9001 2535 9007 2561
rect 672 2365 9376 2382
rect 672 2339 2763 2365
rect 2789 2339 2815 2365
rect 2841 2339 2867 2365
rect 2893 2339 4919 2365
rect 4945 2339 4971 2365
rect 4997 2339 5023 2365
rect 5049 2339 7075 2365
rect 7101 2339 7127 2365
rect 7153 2339 7179 2365
rect 7205 2339 9231 2365
rect 9257 2339 9283 2365
rect 9309 2339 9335 2365
rect 9361 2339 9376 2365
rect 672 2322 9376 2339
rect 1023 2281 1049 2287
rect 1023 2249 1049 2255
rect 7911 2281 7937 2287
rect 9087 2281 9113 2287
rect 8689 2255 8695 2281
rect 8721 2255 8727 2281
rect 7911 2249 7937 2255
rect 9087 2249 9113 2255
rect 855 2169 881 2175
rect 6953 2143 6959 2169
rect 6985 2143 6991 2169
rect 8185 2143 8191 2169
rect 8217 2143 8223 2169
rect 8801 2143 8807 2169
rect 8833 2143 8839 2169
rect 855 2137 881 2143
rect 1247 2113 1273 2119
rect 1247 2081 1273 2087
rect 6455 2057 6481 2063
rect 6455 2025 6481 2031
rect 672 1973 9296 1990
rect 672 1947 1685 1973
rect 1711 1947 1737 1973
rect 1763 1947 1789 1973
rect 1815 1947 3841 1973
rect 3867 1947 3893 1973
rect 3919 1947 3945 1973
rect 3971 1947 5997 1973
rect 6023 1947 6049 1973
rect 6075 1947 6101 1973
rect 6127 1947 8153 1973
rect 8179 1947 8205 1973
rect 8231 1947 8257 1973
rect 8283 1947 9296 1973
rect 672 1930 9296 1947
rect 8471 1889 8497 1895
rect 8471 1857 8497 1863
rect 8527 1833 8553 1839
rect 7513 1807 7519 1833
rect 7545 1807 7551 1833
rect 8527 1801 8553 1807
rect 6281 1751 6287 1777
rect 6313 1751 6319 1777
rect 8185 1751 8191 1777
rect 8217 1751 8223 1777
rect 855 1721 881 1727
rect 855 1689 881 1695
rect 1023 1721 1049 1727
rect 1023 1689 1049 1695
rect 1247 1721 1273 1727
rect 1247 1689 1273 1695
rect 5783 1665 5809 1671
rect 5783 1633 5809 1639
rect 672 1581 9376 1598
rect 672 1555 2763 1581
rect 2789 1555 2815 1581
rect 2841 1555 2867 1581
rect 2893 1555 4919 1581
rect 4945 1555 4971 1581
rect 4997 1555 5023 1581
rect 5049 1555 7075 1581
rect 7101 1555 7127 1581
rect 7153 1555 7179 1581
rect 7205 1555 9231 1581
rect 9257 1555 9283 1581
rect 9309 1555 9335 1581
rect 9361 1555 9376 1581
rect 672 1538 9376 1555
<< via1 >>
rect 1685 8219 1711 8245
rect 1737 8219 1763 8245
rect 1789 8219 1815 8245
rect 3841 8219 3867 8245
rect 3893 8219 3919 8245
rect 3945 8219 3971 8245
rect 5997 8219 6023 8245
rect 6049 8219 6075 8245
rect 6101 8219 6127 8245
rect 8153 8219 8179 8245
rect 8205 8219 8231 8245
rect 8257 8219 8283 8245
rect 5783 8135 5809 8161
rect 7463 8135 7489 8161
rect 855 8023 881 8049
rect 1191 8023 1217 8049
rect 1583 8023 1609 8049
rect 6287 8023 6313 8049
rect 7967 8023 7993 8049
rect 8583 8023 8609 8049
rect 8919 8023 8945 8049
rect 8807 7967 8833 7993
rect 1023 7911 1049 7937
rect 1359 7911 1385 7937
rect 8471 7911 8497 7937
rect 2763 7827 2789 7853
rect 2815 7827 2841 7853
rect 2867 7827 2893 7853
rect 4919 7827 4945 7853
rect 4971 7827 4997 7853
rect 5023 7827 5049 7853
rect 7075 7827 7101 7853
rect 7127 7827 7153 7853
rect 7179 7827 7205 7853
rect 9231 7827 9257 7853
rect 9283 7827 9309 7853
rect 9335 7827 9361 7853
rect 1079 7743 1105 7769
rect 6455 7743 6481 7769
rect 8695 7687 8721 7713
rect 9087 7687 9113 7713
rect 6959 7631 6985 7657
rect 8415 7631 8441 7657
rect 8807 7631 8833 7657
rect 7911 7575 7937 7601
rect 9031 7519 9057 7545
rect 1685 7435 1711 7461
rect 1737 7435 1763 7461
rect 1789 7435 1815 7461
rect 3841 7435 3867 7461
rect 3893 7435 3919 7461
rect 3945 7435 3971 7461
rect 5997 7435 6023 7461
rect 6049 7435 6075 7461
rect 6101 7435 6127 7461
rect 8153 7435 8179 7461
rect 8205 7435 8231 7461
rect 8257 7435 8283 7461
rect 7631 7239 7657 7265
rect 8919 7239 8945 7265
rect 855 7183 881 7209
rect 1023 7183 1049 7209
rect 1247 7183 1273 7209
rect 7575 7127 7601 7153
rect 8583 7127 8609 7153
rect 2763 7043 2789 7069
rect 2815 7043 2841 7069
rect 2867 7043 2893 7069
rect 4919 7043 4945 7069
rect 4971 7043 4997 7069
rect 5023 7043 5049 7069
rect 7075 7043 7101 7069
rect 7127 7043 7153 7069
rect 7179 7043 7205 7069
rect 9231 7043 9257 7069
rect 9283 7043 9309 7069
rect 9335 7043 9361 7069
rect 8695 6959 8721 6985
rect 9087 6903 9113 6929
rect 8359 6847 8385 6873
rect 8807 6847 8833 6873
rect 7799 6791 7825 6817
rect 9031 6735 9057 6761
rect 1685 6651 1711 6677
rect 1737 6651 1763 6677
rect 1789 6651 1815 6677
rect 3841 6651 3867 6677
rect 3893 6651 3919 6677
rect 3945 6651 3971 6677
rect 5997 6651 6023 6677
rect 6049 6651 6075 6677
rect 6101 6651 6127 6677
rect 8153 6651 8179 6677
rect 8205 6651 8231 6677
rect 8257 6651 8283 6677
rect 8583 6511 8609 6537
rect 8863 6455 8889 6481
rect 855 6399 881 6425
rect 1023 6399 1049 6425
rect 1247 6343 1273 6369
rect 2763 6259 2789 6285
rect 2815 6259 2841 6285
rect 2867 6259 2893 6285
rect 4919 6259 4945 6285
rect 4971 6259 4997 6285
rect 5023 6259 5049 6285
rect 7075 6259 7101 6285
rect 7127 6259 7153 6285
rect 7179 6259 7205 6285
rect 9231 6259 9257 6285
rect 9283 6259 9309 6285
rect 9335 6259 9361 6285
rect 8751 6119 8777 6145
rect 9031 6007 9057 6033
rect 8695 5951 8721 5977
rect 1685 5867 1711 5893
rect 1737 5867 1763 5893
rect 1789 5867 1815 5893
rect 3841 5867 3867 5893
rect 3893 5867 3919 5893
rect 3945 5867 3971 5893
rect 5997 5867 6023 5893
rect 6049 5867 6075 5893
rect 6101 5867 6127 5893
rect 8153 5867 8179 5893
rect 8205 5867 8231 5893
rect 8257 5867 8283 5893
rect 8975 5783 9001 5809
rect 7799 5671 7825 5697
rect 855 5615 881 5641
rect 1023 5615 1049 5641
rect 1247 5559 1273 5585
rect 2763 5475 2789 5501
rect 2815 5475 2841 5501
rect 2867 5475 2893 5501
rect 4919 5475 4945 5501
rect 4971 5475 4997 5501
rect 5023 5475 5049 5501
rect 7075 5475 7101 5501
rect 7127 5475 7153 5501
rect 7179 5475 7205 5501
rect 9231 5475 9257 5501
rect 9283 5475 9309 5501
rect 9335 5475 9361 5501
rect 8863 5391 8889 5417
rect 8695 5335 8721 5361
rect 9087 5335 9113 5361
rect 7351 5279 7377 5305
rect 8303 5167 8329 5193
rect 1685 5083 1711 5109
rect 1737 5083 1763 5109
rect 1789 5083 1815 5109
rect 3841 5083 3867 5109
rect 3893 5083 3919 5109
rect 3945 5083 3971 5109
rect 5997 5083 6023 5109
rect 6049 5083 6075 5109
rect 6101 5083 6127 5109
rect 8153 5083 8179 5109
rect 8205 5083 8231 5109
rect 8257 5083 8283 5109
rect 8583 4999 8609 5025
rect 7575 4887 7601 4913
rect 8863 4887 8889 4913
rect 855 4831 881 4857
rect 1247 4831 1273 4857
rect 7463 4831 7489 4857
rect 1023 4775 1049 4801
rect 7351 4775 7377 4801
rect 2763 4691 2789 4717
rect 2815 4691 2841 4717
rect 2867 4691 2893 4717
rect 4919 4691 4945 4717
rect 4971 4691 4997 4717
rect 5023 4691 5049 4717
rect 7075 4691 7101 4717
rect 7127 4691 7153 4717
rect 7179 4691 7205 4717
rect 9231 4691 9257 4717
rect 9283 4691 9309 4717
rect 9335 4691 9361 4717
rect 6959 4607 6985 4633
rect 8695 4607 8721 4633
rect 8863 4551 8889 4577
rect 9087 4551 9113 4577
rect 7239 4495 7265 4521
rect 8303 4383 8329 4409
rect 9031 4383 9057 4409
rect 1685 4299 1711 4325
rect 1737 4299 1763 4325
rect 1789 4299 1815 4325
rect 3841 4299 3867 4325
rect 3893 4299 3919 4325
rect 3945 4299 3971 4325
rect 5997 4299 6023 4325
rect 6049 4299 6075 4325
rect 6101 4299 6127 4325
rect 8153 4299 8179 4325
rect 8205 4299 8231 4325
rect 8257 4299 8283 4325
rect 7239 4215 7265 4241
rect 8583 4215 8609 4241
rect 9031 4103 9057 4129
rect 7295 4047 7321 4073
rect 7463 4047 7489 4073
rect 7631 4047 7657 4073
rect 7127 3991 7153 4017
rect 2763 3907 2789 3933
rect 2815 3907 2841 3933
rect 2867 3907 2893 3933
rect 4919 3907 4945 3933
rect 4971 3907 4997 3933
rect 5023 3907 5049 3933
rect 7075 3907 7101 3933
rect 7127 3907 7153 3933
rect 7179 3907 7205 3933
rect 9231 3907 9257 3933
rect 9283 3907 9309 3933
rect 9335 3907 9361 3933
rect 8695 3823 8721 3849
rect 9031 3823 9057 3849
rect 1023 3767 1049 3793
rect 855 3711 881 3737
rect 8359 3711 8385 3737
rect 8807 3711 8833 3737
rect 1247 3655 1273 3681
rect 9087 3655 9113 3681
rect 7911 3599 7937 3625
rect 1685 3515 1711 3541
rect 1737 3515 1763 3541
rect 1789 3515 1815 3541
rect 3841 3515 3867 3541
rect 3893 3515 3919 3541
rect 3945 3515 3971 3541
rect 5997 3515 6023 3541
rect 6049 3515 6075 3541
rect 6101 3515 6127 3541
rect 8153 3515 8179 3541
rect 8205 3515 8231 3541
rect 8257 3515 8283 3541
rect 8583 3431 8609 3457
rect 8975 3319 9001 3345
rect 7631 3207 7657 3233
rect 2763 3123 2789 3149
rect 2815 3123 2841 3149
rect 2867 3123 2893 3149
rect 4919 3123 4945 3149
rect 4971 3123 4997 3149
rect 5023 3123 5049 3149
rect 7075 3123 7101 3149
rect 7127 3123 7153 3149
rect 7179 3123 7205 3149
rect 9231 3123 9257 3149
rect 9283 3123 9309 3149
rect 9335 3123 9361 3149
rect 1023 3039 1049 3065
rect 8695 3039 8721 3065
rect 8975 3039 9001 3065
rect 8751 2983 8777 3009
rect 8919 2983 8945 3009
rect 855 2927 881 2953
rect 7351 2927 7377 2953
rect 1247 2871 1273 2897
rect 7631 2815 7657 2841
rect 1685 2731 1711 2757
rect 1737 2731 1763 2757
rect 1789 2731 1815 2757
rect 3841 2731 3867 2757
rect 3893 2731 3919 2757
rect 3945 2731 3971 2757
rect 5997 2731 6023 2757
rect 6049 2731 6075 2757
rect 6101 2731 6127 2757
rect 8153 2731 8179 2757
rect 8205 2731 8231 2757
rect 8257 2731 8283 2757
rect 8359 2647 8385 2673
rect 7687 2591 7713 2617
rect 8975 2535 9001 2561
rect 2763 2339 2789 2365
rect 2815 2339 2841 2365
rect 2867 2339 2893 2365
rect 4919 2339 4945 2365
rect 4971 2339 4997 2365
rect 5023 2339 5049 2365
rect 7075 2339 7101 2365
rect 7127 2339 7153 2365
rect 7179 2339 7205 2365
rect 9231 2339 9257 2365
rect 9283 2339 9309 2365
rect 9335 2339 9361 2365
rect 1023 2255 1049 2281
rect 7911 2255 7937 2281
rect 8695 2255 8721 2281
rect 9087 2255 9113 2281
rect 855 2143 881 2169
rect 6959 2143 6985 2169
rect 8191 2143 8217 2169
rect 8807 2143 8833 2169
rect 1247 2087 1273 2113
rect 6455 2031 6481 2057
rect 1685 1947 1711 1973
rect 1737 1947 1763 1973
rect 1789 1947 1815 1973
rect 3841 1947 3867 1973
rect 3893 1947 3919 1973
rect 3945 1947 3971 1973
rect 5997 1947 6023 1973
rect 6049 1947 6075 1973
rect 6101 1947 6127 1973
rect 8153 1947 8179 1973
rect 8205 1947 8231 1973
rect 8257 1947 8283 1973
rect 8471 1863 8497 1889
rect 7519 1807 7545 1833
rect 8527 1807 8553 1833
rect 6287 1751 6313 1777
rect 8191 1751 8217 1777
rect 855 1695 881 1721
rect 1023 1695 1049 1721
rect 1247 1695 1273 1721
rect 5783 1639 5809 1665
rect 2763 1555 2789 1581
rect 2815 1555 2841 1581
rect 2867 1555 2893 1581
rect 4919 1555 4945 1581
rect 4971 1555 4997 1581
rect 5023 1555 5049 1581
rect 7075 1555 7101 1581
rect 7127 1555 7153 1581
rect 7179 1555 7205 1581
rect 9231 1555 9257 1581
rect 9283 1555 9309 1581
rect 9335 1555 9361 1581
<< metal2 >>
rect 7462 9226 7490 9231
rect 854 9002 882 9007
rect 854 8050 882 8974
rect 5782 8778 5810 8783
rect 1684 8246 1816 8251
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1684 8213 1816 8218
rect 3840 8246 3972 8251
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3840 8213 3972 8218
rect 5782 8161 5810 8750
rect 6454 8330 6482 8335
rect 5996 8246 6128 8251
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 5996 8213 6128 8218
rect 5782 8135 5783 8161
rect 5809 8135 5810 8161
rect 5782 8129 5810 8135
rect 1190 8106 1218 8111
rect 1190 8050 1218 8078
rect 854 8003 882 8022
rect 1078 8049 1218 8050
rect 1078 8023 1191 8049
rect 1217 8023 1218 8049
rect 1078 8022 1218 8023
rect 1022 7938 1050 7943
rect 1022 7891 1050 7910
rect 1078 7769 1106 8022
rect 1190 8017 1218 8022
rect 1582 8050 1610 8055
rect 1582 8003 1610 8022
rect 6286 8050 6314 8055
rect 6286 8003 6314 8022
rect 1078 7743 1079 7769
rect 1105 7743 1106 7769
rect 1078 7737 1106 7743
rect 1358 7937 1386 7943
rect 1358 7911 1359 7937
rect 1385 7911 1386 7937
rect 1358 7770 1386 7911
rect 2762 7854 2894 7859
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2762 7821 2894 7826
rect 4918 7854 5050 7859
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 4918 7821 5050 7826
rect 1358 7737 1386 7742
rect 6454 7769 6482 8302
rect 7462 8161 7490 9198
rect 8152 8246 8284 8251
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8152 8213 8284 8218
rect 7462 8135 7463 8161
rect 7489 8135 7490 8161
rect 7462 8129 7490 8135
rect 7966 8049 7994 8055
rect 7966 8023 7967 8049
rect 7993 8023 7994 8049
rect 6454 7743 6455 7769
rect 6481 7743 6482 7769
rect 6454 7737 6482 7743
rect 6958 7938 6986 7943
rect 6958 7657 6986 7910
rect 7798 7882 7826 7887
rect 7074 7854 7206 7859
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7074 7821 7206 7826
rect 6958 7631 6959 7657
rect 6985 7631 6986 7657
rect 6958 7625 6986 7631
rect 7630 7770 7658 7775
rect 1684 7462 1816 7467
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1684 7429 1816 7434
rect 3840 7462 3972 7467
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3840 7429 3972 7434
rect 5996 7462 6128 7467
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 5996 7429 6128 7434
rect 1022 7266 1050 7271
rect 854 7210 882 7215
rect 854 7163 882 7182
rect 1022 7209 1050 7238
rect 7630 7265 7658 7742
rect 7630 7239 7631 7265
rect 7657 7239 7658 7265
rect 7630 7233 7658 7239
rect 1022 7183 1023 7209
rect 1049 7183 1050 7209
rect 1022 7177 1050 7183
rect 1246 7210 1274 7215
rect 1246 7163 1274 7182
rect 7574 7154 7602 7159
rect 7518 7153 7602 7154
rect 7518 7127 7575 7153
rect 7601 7127 7602 7153
rect 7518 7126 7602 7127
rect 2762 7070 2894 7075
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2762 7037 2894 7042
rect 4918 7070 5050 7075
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 4918 7037 5050 7042
rect 7074 7070 7206 7075
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7074 7037 7206 7042
rect 1684 6678 1816 6683
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1684 6645 1816 6650
rect 3840 6678 3972 6683
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3840 6645 3972 6650
rect 5996 6678 6128 6683
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 5996 6645 6128 6650
rect 854 6425 882 6431
rect 854 6399 855 6425
rect 881 6399 882 6425
rect 854 6314 882 6399
rect 1022 6426 1050 6431
rect 1022 6379 1050 6398
rect 854 6281 882 6286
rect 1246 6369 1274 6375
rect 1246 6343 1247 6369
rect 1273 6343 1274 6369
rect 1246 6314 1274 6343
rect 1246 6281 1274 6286
rect 2762 6286 2894 6291
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2762 6253 2894 6258
rect 4918 6286 5050 6291
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 4918 6253 5050 6258
rect 7074 6286 7206 6291
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7074 6253 7206 6258
rect 1684 5894 1816 5899
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1684 5861 1816 5866
rect 3840 5894 3972 5899
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3840 5861 3972 5866
rect 5996 5894 6128 5899
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 5996 5861 6128 5866
rect 1022 5698 1050 5703
rect 854 5641 882 5647
rect 854 5615 855 5641
rect 881 5615 882 5641
rect 854 5418 882 5615
rect 1022 5641 1050 5670
rect 1022 5615 1023 5641
rect 1049 5615 1050 5641
rect 1022 5609 1050 5615
rect 854 5385 882 5390
rect 1246 5585 1274 5591
rect 1246 5559 1247 5585
rect 1273 5559 1274 5585
rect 1246 5418 1274 5559
rect 2762 5502 2894 5507
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2762 5469 2894 5474
rect 4918 5502 5050 5507
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 4918 5469 5050 5474
rect 7074 5502 7206 5507
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7074 5469 7206 5474
rect 1246 5385 1274 5390
rect 7350 5306 7378 5311
rect 7350 5305 7490 5306
rect 7350 5279 7351 5305
rect 7377 5279 7490 5305
rect 7350 5278 7490 5279
rect 7350 5273 7378 5278
rect 1684 5110 1816 5115
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1684 5077 1816 5082
rect 3840 5110 3972 5115
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3840 5077 3972 5082
rect 5996 5110 6128 5115
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 5996 5077 6128 5082
rect 854 4858 882 4863
rect 854 4522 882 4830
rect 1246 4858 1274 4863
rect 1246 4811 1274 4830
rect 7462 4857 7490 5278
rect 7462 4831 7463 4857
rect 7489 4831 7490 4857
rect 7462 4825 7490 4831
rect 1022 4802 1050 4807
rect 1022 4755 1050 4774
rect 6958 4802 6986 4807
rect 2762 4718 2894 4723
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2762 4685 2894 4690
rect 4918 4718 5050 4723
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 4918 4685 5050 4690
rect 6958 4633 6986 4774
rect 7350 4802 7378 4807
rect 7350 4755 7378 4774
rect 7074 4718 7206 4723
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7074 4685 7206 4690
rect 6958 4607 6959 4633
rect 6985 4607 6986 4633
rect 6958 4578 6986 4607
rect 6958 4545 6986 4550
rect 854 4489 882 4494
rect 7238 4521 7266 4527
rect 7238 4495 7239 4521
rect 7265 4495 7266 4521
rect 1684 4326 1816 4331
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1684 4293 1816 4298
rect 3840 4326 3972 4331
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3840 4293 3972 4298
rect 5996 4326 6128 4331
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 5996 4293 6128 4298
rect 7238 4241 7266 4495
rect 7238 4215 7239 4241
rect 7265 4215 7266 4241
rect 7238 4209 7266 4215
rect 7518 4214 7546 7126
rect 7574 7121 7602 7126
rect 7798 6817 7826 7854
rect 7910 7602 7938 7607
rect 7910 7555 7938 7574
rect 7798 6791 7799 6817
rect 7825 6791 7826 6817
rect 7798 6785 7826 6791
rect 7798 5697 7826 5703
rect 7798 5671 7799 5697
rect 7825 5671 7826 5697
rect 7350 4186 7546 4214
rect 7574 4913 7602 4919
rect 7574 4887 7575 4913
rect 7601 4887 7602 4913
rect 7574 4802 7602 4887
rect 1078 4074 1106 4079
rect 1022 3794 1050 3799
rect 1022 3747 1050 3766
rect 854 3737 882 3743
rect 854 3711 855 3737
rect 881 3711 882 3737
rect 854 3626 882 3711
rect 854 3593 882 3598
rect 1078 3514 1106 4046
rect 7294 4074 7322 4079
rect 7126 4018 7154 4037
rect 7294 4027 7322 4046
rect 7014 3990 7126 4018
rect 2762 3934 2894 3939
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2762 3901 2894 3906
rect 4918 3934 5050 3939
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 4918 3901 5050 3906
rect 7014 3794 7042 3990
rect 7126 3985 7154 3990
rect 7074 3934 7206 3939
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7074 3901 7206 3906
rect 7014 3761 7042 3766
rect 1246 3681 1274 3687
rect 1246 3655 1247 3681
rect 1273 3655 1274 3681
rect 1246 3626 1274 3655
rect 1246 3593 1274 3598
rect 1022 3486 1106 3514
rect 1684 3542 1816 3547
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1684 3509 1816 3514
rect 3840 3542 3972 3547
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3840 3509 3972 3514
rect 5996 3542 6128 3547
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 5996 3509 6128 3514
rect 1022 3065 1050 3486
rect 1022 3039 1023 3065
rect 1049 3039 1050 3065
rect 1022 3033 1050 3039
rect 1078 3234 1106 3239
rect 854 2953 882 2959
rect 854 2927 855 2953
rect 881 2927 882 2953
rect 854 2730 882 2927
rect 854 2697 882 2702
rect 1022 2282 1050 2287
rect 1078 2282 1106 3206
rect 2762 3150 2894 3155
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2762 3117 2894 3122
rect 4918 3150 5050 3155
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 4918 3117 5050 3122
rect 7074 3150 7206 3155
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7074 3117 7206 3122
rect 7350 2953 7378 4186
rect 7462 4073 7490 4079
rect 7462 4047 7463 4073
rect 7489 4047 7490 4073
rect 7462 4018 7490 4047
rect 7462 3985 7490 3990
rect 7574 3234 7602 4774
rect 7798 4214 7826 5671
rect 7686 4186 7826 4214
rect 7630 4074 7658 4079
rect 7686 4074 7714 4186
rect 7630 4073 7714 4074
rect 7630 4047 7631 4073
rect 7657 4047 7714 4073
rect 7630 4046 7714 4047
rect 7630 4041 7658 4046
rect 7910 3625 7938 3631
rect 7910 3599 7911 3625
rect 7937 3599 7938 3625
rect 7910 3402 7938 3599
rect 7910 3369 7938 3374
rect 7630 3234 7658 3239
rect 7574 3206 7630 3234
rect 7630 3187 7658 3206
rect 7350 2927 7351 2953
rect 7377 2927 7378 2953
rect 7350 2921 7378 2927
rect 7686 3010 7714 3015
rect 1246 2897 1274 2903
rect 1246 2871 1247 2897
rect 1273 2871 1274 2897
rect 1246 2730 1274 2871
rect 7630 2841 7658 2847
rect 7630 2815 7631 2841
rect 7657 2815 7658 2841
rect 1684 2758 1816 2763
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1684 2725 1816 2730
rect 3840 2758 3972 2763
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3840 2725 3972 2730
rect 5996 2758 6128 2763
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 5996 2725 6128 2730
rect 1246 2697 1274 2702
rect 7630 2562 7658 2815
rect 7686 2617 7714 2982
rect 7686 2591 7687 2617
rect 7713 2591 7714 2617
rect 7686 2585 7714 2591
rect 7462 2534 7658 2562
rect 2762 2366 2894 2371
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2762 2333 2894 2338
rect 4918 2366 5050 2371
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 4918 2333 5050 2338
rect 7074 2366 7206 2371
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7074 2333 7206 2338
rect 1022 2281 1106 2282
rect 1022 2255 1023 2281
rect 1049 2255 1106 2281
rect 1022 2254 1106 2255
rect 1022 2249 1050 2254
rect 854 2169 882 2175
rect 854 2143 855 2169
rect 881 2143 882 2169
rect 854 2114 882 2143
rect 6958 2170 6986 2175
rect 6958 2123 6986 2142
rect 854 1834 882 2086
rect 1246 2114 1274 2119
rect 1246 2067 1274 2086
rect 6454 2057 6482 2063
rect 6454 2031 6455 2057
rect 6481 2031 6482 2057
rect 1684 1974 1816 1979
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1684 1941 1816 1946
rect 3840 1974 3972 1979
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3840 1941 3972 1946
rect 5996 1974 6128 1979
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 5996 1941 6128 1946
rect 854 1801 882 1806
rect 1022 1834 1050 1839
rect 854 1721 882 1727
rect 854 1695 855 1721
rect 881 1695 882 1721
rect 854 1666 882 1695
rect 1022 1721 1050 1806
rect 6286 1778 6314 1783
rect 6286 1731 6314 1750
rect 1022 1695 1023 1721
rect 1049 1695 1050 1721
rect 1022 1689 1050 1695
rect 1246 1721 1274 1727
rect 1246 1695 1247 1721
rect 1273 1695 1274 1721
rect 854 938 882 1638
rect 1246 1666 1274 1695
rect 1246 1633 1274 1638
rect 5782 1665 5810 1671
rect 5782 1639 5783 1665
rect 5809 1639 5810 1665
rect 2762 1582 2894 1587
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2762 1549 2894 1554
rect 4918 1582 5050 1587
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 4918 1549 5050 1554
rect 5782 1162 5810 1639
rect 5782 1129 5810 1134
rect 854 905 882 910
rect 6454 882 6482 2031
rect 7462 1666 7490 2534
rect 7910 2506 7938 2511
rect 7910 2281 7938 2478
rect 7910 2255 7911 2281
rect 7937 2255 7938 2281
rect 7910 2249 7938 2255
rect 7966 2282 7994 8023
rect 8582 8049 8610 8055
rect 8582 8023 8583 8049
rect 8609 8023 8610 8049
rect 8470 7938 8498 7943
rect 8470 7891 8498 7910
rect 8582 7770 8610 8023
rect 8806 8050 8834 8055
rect 8806 7993 8834 8022
rect 8806 7967 8807 7993
rect 8833 7967 8834 7993
rect 8806 7961 8834 7967
rect 8918 8049 8946 8055
rect 8918 8023 8919 8049
rect 8945 8023 8946 8049
rect 8918 7994 8946 8023
rect 8946 7966 9114 7994
rect 8918 7961 8946 7966
rect 8582 7737 8610 7742
rect 8358 7714 8386 7719
rect 8152 7462 8284 7467
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8152 7429 8284 7434
rect 8358 6873 8386 7686
rect 8694 7714 8722 7719
rect 8694 7667 8722 7686
rect 9086 7713 9114 7966
rect 9230 7854 9362 7859
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9230 7821 9362 7826
rect 9086 7687 9087 7713
rect 9113 7687 9114 7713
rect 9086 7681 9114 7687
rect 8414 7658 8442 7663
rect 8414 7657 8666 7658
rect 8414 7631 8415 7657
rect 8441 7631 8666 7657
rect 8414 7630 8666 7631
rect 8414 7625 8442 7630
rect 8582 7154 8610 7159
rect 8582 7107 8610 7126
rect 8638 6986 8666 7630
rect 8806 7657 8834 7663
rect 8806 7631 8807 7657
rect 8833 7631 8834 7657
rect 8806 7266 8834 7631
rect 9030 7546 9058 7551
rect 9030 7545 9170 7546
rect 9030 7519 9031 7545
rect 9057 7519 9170 7545
rect 9030 7518 9170 7519
rect 9030 7513 9058 7518
rect 8806 7233 8834 7238
rect 8918 7265 8946 7271
rect 8918 7239 8919 7265
rect 8945 7239 8946 7265
rect 8694 6986 8722 6991
rect 8638 6985 8722 6986
rect 8638 6959 8695 6985
rect 8721 6959 8722 6985
rect 8638 6958 8722 6959
rect 8694 6953 8722 6958
rect 8806 6874 8834 6879
rect 8358 6847 8359 6873
rect 8385 6847 8386 6873
rect 8358 6841 8386 6847
rect 8750 6873 8834 6874
rect 8750 6847 8807 6873
rect 8833 6847 8834 6873
rect 8750 6846 8834 6847
rect 8470 6762 8498 6767
rect 8152 6678 8284 6683
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8152 6645 8284 6650
rect 7966 2249 7994 2254
rect 8078 5978 8106 5983
rect 8078 2170 8106 5950
rect 8152 5894 8284 5899
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8152 5861 8284 5866
rect 8302 5194 8330 5213
rect 8302 5161 8330 5166
rect 8152 5110 8284 5115
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8152 5077 8284 5082
rect 8302 4410 8330 4415
rect 8302 4409 8386 4410
rect 8302 4383 8303 4409
rect 8329 4383 8386 4409
rect 8302 4382 8386 4383
rect 8302 4377 8330 4382
rect 8152 4326 8284 4331
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8152 4293 8284 4298
rect 8358 4298 8386 4382
rect 8358 4265 8386 4270
rect 8470 4214 8498 6734
rect 8582 6538 8610 6543
rect 8582 6491 8610 6510
rect 8750 6426 8778 6846
rect 8806 6841 8834 6846
rect 8862 6482 8890 6487
rect 8750 6145 8778 6398
rect 8750 6119 8751 6145
rect 8777 6119 8778 6145
rect 8750 6113 8778 6119
rect 8806 6481 8890 6482
rect 8806 6455 8863 6481
rect 8889 6455 8890 6481
rect 8806 6454 8890 6455
rect 8694 5978 8722 5983
rect 8694 5931 8722 5950
rect 8694 5698 8722 5703
rect 8582 5474 8610 5479
rect 8582 5025 8610 5446
rect 8694 5362 8722 5670
rect 8694 5315 8722 5334
rect 8806 5194 8834 6454
rect 8862 6449 8890 6454
rect 8862 5418 8890 5423
rect 8918 5418 8946 7239
rect 9086 7266 9114 7271
rect 9086 6929 9114 7238
rect 9086 6903 9087 6929
rect 9113 6903 9114 6929
rect 9086 6897 9114 6903
rect 9030 6762 9058 6767
rect 9030 6715 9058 6734
rect 8974 6090 9002 6095
rect 8974 5809 9002 6062
rect 8974 5783 8975 5809
rect 9001 5783 9002 5809
rect 8974 5777 9002 5783
rect 9030 6033 9058 6039
rect 9030 6007 9031 6033
rect 9057 6007 9058 6033
rect 8862 5417 8946 5418
rect 8862 5391 8863 5417
rect 8889 5391 8946 5417
rect 8862 5390 8946 5391
rect 8862 5385 8890 5390
rect 9030 5362 9058 6007
rect 9086 5362 9114 5367
rect 9030 5334 9086 5362
rect 8582 4999 8583 5025
rect 8609 4999 8610 5025
rect 8582 4993 8610 4999
rect 8694 5166 8834 5194
rect 8414 4186 8498 4214
rect 8582 4634 8610 4639
rect 8582 4241 8610 4606
rect 8694 4633 8722 5166
rect 8862 4914 8890 4919
rect 8694 4607 8695 4633
rect 8721 4607 8722 4633
rect 8694 4601 8722 4607
rect 8806 4913 8890 4914
rect 8806 4887 8863 4913
rect 8889 4887 8890 4913
rect 8806 4886 8890 4887
rect 8582 4215 8583 4241
rect 8609 4215 8610 4241
rect 8582 4209 8610 4215
rect 8806 4214 8834 4886
rect 8862 4881 8890 4886
rect 8694 4186 8834 4214
rect 8862 4578 8890 4583
rect 8358 3737 8386 3743
rect 8358 3711 8359 3737
rect 8385 3711 8386 3737
rect 8152 3542 8284 3547
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8152 3509 8284 3514
rect 8358 3066 8386 3711
rect 8358 3033 8386 3038
rect 8358 2954 8386 2959
rect 8152 2758 8284 2763
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8152 2725 8284 2730
rect 8358 2673 8386 2926
rect 8358 2647 8359 2673
rect 8385 2647 8386 2673
rect 8358 2641 8386 2647
rect 8190 2170 8218 2175
rect 8078 2169 8218 2170
rect 8078 2143 8191 2169
rect 8217 2143 8218 2169
rect 8078 2142 8218 2143
rect 8190 2137 8218 2142
rect 7518 2058 7546 2063
rect 7518 1833 7546 2030
rect 8152 1974 8284 1979
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8152 1941 8284 1946
rect 8414 1890 8442 4186
rect 8694 3849 8722 4186
rect 8694 3823 8695 3849
rect 8721 3823 8722 3849
rect 8694 3817 8722 3823
rect 8806 4074 8834 4079
rect 8582 3738 8610 3743
rect 8582 3457 8610 3710
rect 8806 3737 8834 4046
rect 8806 3711 8807 3737
rect 8833 3711 8834 3737
rect 8806 3705 8834 3711
rect 8862 3514 8890 4550
rect 9086 4577 9114 5334
rect 9086 4551 9087 4577
rect 9113 4551 9114 4577
rect 9086 4545 9114 4551
rect 9030 4409 9058 4415
rect 9030 4383 9031 4409
rect 9057 4383 9058 4409
rect 9030 4214 9058 4383
rect 8974 4186 9058 4214
rect 8582 3431 8583 3457
rect 8609 3431 8610 3457
rect 8582 3425 8610 3431
rect 8750 3486 8890 3514
rect 8918 4018 8946 4023
rect 8694 3066 8722 3071
rect 8694 3019 8722 3038
rect 8750 3010 8778 3486
rect 8750 2963 8778 2982
rect 8918 3009 8946 3990
rect 8974 3514 9002 4186
rect 9030 4129 9058 4135
rect 9030 4103 9031 4129
rect 9057 4103 9058 4129
rect 9030 3849 9058 4103
rect 9030 3823 9031 3849
rect 9057 3823 9058 3849
rect 9030 3817 9058 3823
rect 9086 3681 9114 3687
rect 9086 3655 9087 3681
rect 9113 3655 9114 3681
rect 8974 3486 9058 3514
rect 8974 3345 9002 3351
rect 8974 3319 8975 3345
rect 9001 3319 9002 3345
rect 8974 3065 9002 3319
rect 8974 3039 8975 3065
rect 9001 3039 9002 3065
rect 8974 3033 9002 3039
rect 8918 2983 8919 3009
rect 8945 2983 8946 3009
rect 8918 2394 8946 2983
rect 8974 2562 9002 2567
rect 9030 2562 9058 3486
rect 9086 3234 9114 3655
rect 9086 3201 9114 3206
rect 8974 2561 9058 2562
rect 8974 2535 8975 2561
rect 9001 2535 9058 2561
rect 8974 2534 9058 2535
rect 8974 2529 9002 2534
rect 8918 2366 9114 2394
rect 8694 2282 8722 2287
rect 8694 2235 8722 2254
rect 9086 2281 9114 2366
rect 9086 2255 9087 2281
rect 9113 2255 9114 2281
rect 9086 2249 9114 2255
rect 7518 1807 7519 1833
rect 7545 1807 7546 1833
rect 7518 1801 7546 1807
rect 8190 1862 8442 1890
rect 8470 2170 8498 2175
rect 8470 1889 8498 2142
rect 8470 1863 8471 1889
rect 8497 1863 8498 1889
rect 8190 1777 8218 1862
rect 8470 1857 8498 1863
rect 8806 2169 8834 2175
rect 8806 2143 8807 2169
rect 8833 2143 8834 2169
rect 8526 1834 8554 1839
rect 8526 1787 8554 1806
rect 8806 1834 8834 2143
rect 8806 1801 8834 1806
rect 8190 1751 8191 1777
rect 8217 1751 8218 1777
rect 8190 1745 8218 1751
rect 9142 1778 9170 7518
rect 9230 7070 9362 7075
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9230 7037 9362 7042
rect 9230 6286 9362 6291
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9230 6253 9362 6258
rect 9230 5502 9362 5507
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9230 5469 9362 5474
rect 9230 4718 9362 4723
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9230 4685 9362 4690
rect 9230 3934 9362 3939
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9230 3901 9362 3906
rect 9230 3150 9362 3155
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9230 3117 9362 3122
rect 9230 2366 9362 2371
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9230 2333 9362 2338
rect 9142 1745 9170 1750
rect 7518 1666 7546 1671
rect 7462 1638 7518 1666
rect 7518 1633 7546 1638
rect 7074 1582 7206 1587
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7074 1549 7206 1554
rect 9230 1582 9362 1587
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9230 1549 9362 1554
rect 6454 849 6482 854
<< via2 >>
rect 7462 9198 7490 9226
rect 854 8974 882 9002
rect 5782 8750 5810 8778
rect 1684 8245 1712 8246
rect 1684 8219 1685 8245
rect 1685 8219 1711 8245
rect 1711 8219 1712 8245
rect 1684 8218 1712 8219
rect 1736 8245 1764 8246
rect 1736 8219 1737 8245
rect 1737 8219 1763 8245
rect 1763 8219 1764 8245
rect 1736 8218 1764 8219
rect 1788 8245 1816 8246
rect 1788 8219 1789 8245
rect 1789 8219 1815 8245
rect 1815 8219 1816 8245
rect 1788 8218 1816 8219
rect 3840 8245 3868 8246
rect 3840 8219 3841 8245
rect 3841 8219 3867 8245
rect 3867 8219 3868 8245
rect 3840 8218 3868 8219
rect 3892 8245 3920 8246
rect 3892 8219 3893 8245
rect 3893 8219 3919 8245
rect 3919 8219 3920 8245
rect 3892 8218 3920 8219
rect 3944 8245 3972 8246
rect 3944 8219 3945 8245
rect 3945 8219 3971 8245
rect 3971 8219 3972 8245
rect 3944 8218 3972 8219
rect 6454 8302 6482 8330
rect 5996 8245 6024 8246
rect 5996 8219 5997 8245
rect 5997 8219 6023 8245
rect 6023 8219 6024 8245
rect 5996 8218 6024 8219
rect 6048 8245 6076 8246
rect 6048 8219 6049 8245
rect 6049 8219 6075 8245
rect 6075 8219 6076 8245
rect 6048 8218 6076 8219
rect 6100 8245 6128 8246
rect 6100 8219 6101 8245
rect 6101 8219 6127 8245
rect 6127 8219 6128 8245
rect 6100 8218 6128 8219
rect 1190 8078 1218 8106
rect 854 8049 882 8050
rect 854 8023 855 8049
rect 855 8023 881 8049
rect 881 8023 882 8049
rect 854 8022 882 8023
rect 1022 7937 1050 7938
rect 1022 7911 1023 7937
rect 1023 7911 1049 7937
rect 1049 7911 1050 7937
rect 1022 7910 1050 7911
rect 1582 8049 1610 8050
rect 1582 8023 1583 8049
rect 1583 8023 1609 8049
rect 1609 8023 1610 8049
rect 1582 8022 1610 8023
rect 6286 8049 6314 8050
rect 6286 8023 6287 8049
rect 6287 8023 6313 8049
rect 6313 8023 6314 8049
rect 6286 8022 6314 8023
rect 2762 7853 2790 7854
rect 2762 7827 2763 7853
rect 2763 7827 2789 7853
rect 2789 7827 2790 7853
rect 2762 7826 2790 7827
rect 2814 7853 2842 7854
rect 2814 7827 2815 7853
rect 2815 7827 2841 7853
rect 2841 7827 2842 7853
rect 2814 7826 2842 7827
rect 2866 7853 2894 7854
rect 2866 7827 2867 7853
rect 2867 7827 2893 7853
rect 2893 7827 2894 7853
rect 2866 7826 2894 7827
rect 4918 7853 4946 7854
rect 4918 7827 4919 7853
rect 4919 7827 4945 7853
rect 4945 7827 4946 7853
rect 4918 7826 4946 7827
rect 4970 7853 4998 7854
rect 4970 7827 4971 7853
rect 4971 7827 4997 7853
rect 4997 7827 4998 7853
rect 4970 7826 4998 7827
rect 5022 7853 5050 7854
rect 5022 7827 5023 7853
rect 5023 7827 5049 7853
rect 5049 7827 5050 7853
rect 5022 7826 5050 7827
rect 1358 7742 1386 7770
rect 8152 8245 8180 8246
rect 8152 8219 8153 8245
rect 8153 8219 8179 8245
rect 8179 8219 8180 8245
rect 8152 8218 8180 8219
rect 8204 8245 8232 8246
rect 8204 8219 8205 8245
rect 8205 8219 8231 8245
rect 8231 8219 8232 8245
rect 8204 8218 8232 8219
rect 8256 8245 8284 8246
rect 8256 8219 8257 8245
rect 8257 8219 8283 8245
rect 8283 8219 8284 8245
rect 8256 8218 8284 8219
rect 6958 7910 6986 7938
rect 7074 7853 7102 7854
rect 7074 7827 7075 7853
rect 7075 7827 7101 7853
rect 7101 7827 7102 7853
rect 7074 7826 7102 7827
rect 7126 7853 7154 7854
rect 7126 7827 7127 7853
rect 7127 7827 7153 7853
rect 7153 7827 7154 7853
rect 7126 7826 7154 7827
rect 7178 7853 7206 7854
rect 7178 7827 7179 7853
rect 7179 7827 7205 7853
rect 7205 7827 7206 7853
rect 7178 7826 7206 7827
rect 7798 7854 7826 7882
rect 7630 7742 7658 7770
rect 1684 7461 1712 7462
rect 1684 7435 1685 7461
rect 1685 7435 1711 7461
rect 1711 7435 1712 7461
rect 1684 7434 1712 7435
rect 1736 7461 1764 7462
rect 1736 7435 1737 7461
rect 1737 7435 1763 7461
rect 1763 7435 1764 7461
rect 1736 7434 1764 7435
rect 1788 7461 1816 7462
rect 1788 7435 1789 7461
rect 1789 7435 1815 7461
rect 1815 7435 1816 7461
rect 1788 7434 1816 7435
rect 3840 7461 3868 7462
rect 3840 7435 3841 7461
rect 3841 7435 3867 7461
rect 3867 7435 3868 7461
rect 3840 7434 3868 7435
rect 3892 7461 3920 7462
rect 3892 7435 3893 7461
rect 3893 7435 3919 7461
rect 3919 7435 3920 7461
rect 3892 7434 3920 7435
rect 3944 7461 3972 7462
rect 3944 7435 3945 7461
rect 3945 7435 3971 7461
rect 3971 7435 3972 7461
rect 3944 7434 3972 7435
rect 5996 7461 6024 7462
rect 5996 7435 5997 7461
rect 5997 7435 6023 7461
rect 6023 7435 6024 7461
rect 5996 7434 6024 7435
rect 6048 7461 6076 7462
rect 6048 7435 6049 7461
rect 6049 7435 6075 7461
rect 6075 7435 6076 7461
rect 6048 7434 6076 7435
rect 6100 7461 6128 7462
rect 6100 7435 6101 7461
rect 6101 7435 6127 7461
rect 6127 7435 6128 7461
rect 6100 7434 6128 7435
rect 1022 7238 1050 7266
rect 854 7209 882 7210
rect 854 7183 855 7209
rect 855 7183 881 7209
rect 881 7183 882 7209
rect 854 7182 882 7183
rect 1246 7209 1274 7210
rect 1246 7183 1247 7209
rect 1247 7183 1273 7209
rect 1273 7183 1274 7209
rect 1246 7182 1274 7183
rect 2762 7069 2790 7070
rect 2762 7043 2763 7069
rect 2763 7043 2789 7069
rect 2789 7043 2790 7069
rect 2762 7042 2790 7043
rect 2814 7069 2842 7070
rect 2814 7043 2815 7069
rect 2815 7043 2841 7069
rect 2841 7043 2842 7069
rect 2814 7042 2842 7043
rect 2866 7069 2894 7070
rect 2866 7043 2867 7069
rect 2867 7043 2893 7069
rect 2893 7043 2894 7069
rect 2866 7042 2894 7043
rect 4918 7069 4946 7070
rect 4918 7043 4919 7069
rect 4919 7043 4945 7069
rect 4945 7043 4946 7069
rect 4918 7042 4946 7043
rect 4970 7069 4998 7070
rect 4970 7043 4971 7069
rect 4971 7043 4997 7069
rect 4997 7043 4998 7069
rect 4970 7042 4998 7043
rect 5022 7069 5050 7070
rect 5022 7043 5023 7069
rect 5023 7043 5049 7069
rect 5049 7043 5050 7069
rect 5022 7042 5050 7043
rect 7074 7069 7102 7070
rect 7074 7043 7075 7069
rect 7075 7043 7101 7069
rect 7101 7043 7102 7069
rect 7074 7042 7102 7043
rect 7126 7069 7154 7070
rect 7126 7043 7127 7069
rect 7127 7043 7153 7069
rect 7153 7043 7154 7069
rect 7126 7042 7154 7043
rect 7178 7069 7206 7070
rect 7178 7043 7179 7069
rect 7179 7043 7205 7069
rect 7205 7043 7206 7069
rect 7178 7042 7206 7043
rect 1684 6677 1712 6678
rect 1684 6651 1685 6677
rect 1685 6651 1711 6677
rect 1711 6651 1712 6677
rect 1684 6650 1712 6651
rect 1736 6677 1764 6678
rect 1736 6651 1737 6677
rect 1737 6651 1763 6677
rect 1763 6651 1764 6677
rect 1736 6650 1764 6651
rect 1788 6677 1816 6678
rect 1788 6651 1789 6677
rect 1789 6651 1815 6677
rect 1815 6651 1816 6677
rect 1788 6650 1816 6651
rect 3840 6677 3868 6678
rect 3840 6651 3841 6677
rect 3841 6651 3867 6677
rect 3867 6651 3868 6677
rect 3840 6650 3868 6651
rect 3892 6677 3920 6678
rect 3892 6651 3893 6677
rect 3893 6651 3919 6677
rect 3919 6651 3920 6677
rect 3892 6650 3920 6651
rect 3944 6677 3972 6678
rect 3944 6651 3945 6677
rect 3945 6651 3971 6677
rect 3971 6651 3972 6677
rect 3944 6650 3972 6651
rect 5996 6677 6024 6678
rect 5996 6651 5997 6677
rect 5997 6651 6023 6677
rect 6023 6651 6024 6677
rect 5996 6650 6024 6651
rect 6048 6677 6076 6678
rect 6048 6651 6049 6677
rect 6049 6651 6075 6677
rect 6075 6651 6076 6677
rect 6048 6650 6076 6651
rect 6100 6677 6128 6678
rect 6100 6651 6101 6677
rect 6101 6651 6127 6677
rect 6127 6651 6128 6677
rect 6100 6650 6128 6651
rect 1022 6425 1050 6426
rect 1022 6399 1023 6425
rect 1023 6399 1049 6425
rect 1049 6399 1050 6425
rect 1022 6398 1050 6399
rect 854 6286 882 6314
rect 1246 6286 1274 6314
rect 2762 6285 2790 6286
rect 2762 6259 2763 6285
rect 2763 6259 2789 6285
rect 2789 6259 2790 6285
rect 2762 6258 2790 6259
rect 2814 6285 2842 6286
rect 2814 6259 2815 6285
rect 2815 6259 2841 6285
rect 2841 6259 2842 6285
rect 2814 6258 2842 6259
rect 2866 6285 2894 6286
rect 2866 6259 2867 6285
rect 2867 6259 2893 6285
rect 2893 6259 2894 6285
rect 2866 6258 2894 6259
rect 4918 6285 4946 6286
rect 4918 6259 4919 6285
rect 4919 6259 4945 6285
rect 4945 6259 4946 6285
rect 4918 6258 4946 6259
rect 4970 6285 4998 6286
rect 4970 6259 4971 6285
rect 4971 6259 4997 6285
rect 4997 6259 4998 6285
rect 4970 6258 4998 6259
rect 5022 6285 5050 6286
rect 5022 6259 5023 6285
rect 5023 6259 5049 6285
rect 5049 6259 5050 6285
rect 5022 6258 5050 6259
rect 7074 6285 7102 6286
rect 7074 6259 7075 6285
rect 7075 6259 7101 6285
rect 7101 6259 7102 6285
rect 7074 6258 7102 6259
rect 7126 6285 7154 6286
rect 7126 6259 7127 6285
rect 7127 6259 7153 6285
rect 7153 6259 7154 6285
rect 7126 6258 7154 6259
rect 7178 6285 7206 6286
rect 7178 6259 7179 6285
rect 7179 6259 7205 6285
rect 7205 6259 7206 6285
rect 7178 6258 7206 6259
rect 1684 5893 1712 5894
rect 1684 5867 1685 5893
rect 1685 5867 1711 5893
rect 1711 5867 1712 5893
rect 1684 5866 1712 5867
rect 1736 5893 1764 5894
rect 1736 5867 1737 5893
rect 1737 5867 1763 5893
rect 1763 5867 1764 5893
rect 1736 5866 1764 5867
rect 1788 5893 1816 5894
rect 1788 5867 1789 5893
rect 1789 5867 1815 5893
rect 1815 5867 1816 5893
rect 1788 5866 1816 5867
rect 3840 5893 3868 5894
rect 3840 5867 3841 5893
rect 3841 5867 3867 5893
rect 3867 5867 3868 5893
rect 3840 5866 3868 5867
rect 3892 5893 3920 5894
rect 3892 5867 3893 5893
rect 3893 5867 3919 5893
rect 3919 5867 3920 5893
rect 3892 5866 3920 5867
rect 3944 5893 3972 5894
rect 3944 5867 3945 5893
rect 3945 5867 3971 5893
rect 3971 5867 3972 5893
rect 3944 5866 3972 5867
rect 5996 5893 6024 5894
rect 5996 5867 5997 5893
rect 5997 5867 6023 5893
rect 6023 5867 6024 5893
rect 5996 5866 6024 5867
rect 6048 5893 6076 5894
rect 6048 5867 6049 5893
rect 6049 5867 6075 5893
rect 6075 5867 6076 5893
rect 6048 5866 6076 5867
rect 6100 5893 6128 5894
rect 6100 5867 6101 5893
rect 6101 5867 6127 5893
rect 6127 5867 6128 5893
rect 6100 5866 6128 5867
rect 1022 5670 1050 5698
rect 854 5390 882 5418
rect 2762 5501 2790 5502
rect 2762 5475 2763 5501
rect 2763 5475 2789 5501
rect 2789 5475 2790 5501
rect 2762 5474 2790 5475
rect 2814 5501 2842 5502
rect 2814 5475 2815 5501
rect 2815 5475 2841 5501
rect 2841 5475 2842 5501
rect 2814 5474 2842 5475
rect 2866 5501 2894 5502
rect 2866 5475 2867 5501
rect 2867 5475 2893 5501
rect 2893 5475 2894 5501
rect 2866 5474 2894 5475
rect 4918 5501 4946 5502
rect 4918 5475 4919 5501
rect 4919 5475 4945 5501
rect 4945 5475 4946 5501
rect 4918 5474 4946 5475
rect 4970 5501 4998 5502
rect 4970 5475 4971 5501
rect 4971 5475 4997 5501
rect 4997 5475 4998 5501
rect 4970 5474 4998 5475
rect 5022 5501 5050 5502
rect 5022 5475 5023 5501
rect 5023 5475 5049 5501
rect 5049 5475 5050 5501
rect 5022 5474 5050 5475
rect 7074 5501 7102 5502
rect 7074 5475 7075 5501
rect 7075 5475 7101 5501
rect 7101 5475 7102 5501
rect 7074 5474 7102 5475
rect 7126 5501 7154 5502
rect 7126 5475 7127 5501
rect 7127 5475 7153 5501
rect 7153 5475 7154 5501
rect 7126 5474 7154 5475
rect 7178 5501 7206 5502
rect 7178 5475 7179 5501
rect 7179 5475 7205 5501
rect 7205 5475 7206 5501
rect 7178 5474 7206 5475
rect 1246 5390 1274 5418
rect 1684 5109 1712 5110
rect 1684 5083 1685 5109
rect 1685 5083 1711 5109
rect 1711 5083 1712 5109
rect 1684 5082 1712 5083
rect 1736 5109 1764 5110
rect 1736 5083 1737 5109
rect 1737 5083 1763 5109
rect 1763 5083 1764 5109
rect 1736 5082 1764 5083
rect 1788 5109 1816 5110
rect 1788 5083 1789 5109
rect 1789 5083 1815 5109
rect 1815 5083 1816 5109
rect 1788 5082 1816 5083
rect 3840 5109 3868 5110
rect 3840 5083 3841 5109
rect 3841 5083 3867 5109
rect 3867 5083 3868 5109
rect 3840 5082 3868 5083
rect 3892 5109 3920 5110
rect 3892 5083 3893 5109
rect 3893 5083 3919 5109
rect 3919 5083 3920 5109
rect 3892 5082 3920 5083
rect 3944 5109 3972 5110
rect 3944 5083 3945 5109
rect 3945 5083 3971 5109
rect 3971 5083 3972 5109
rect 3944 5082 3972 5083
rect 5996 5109 6024 5110
rect 5996 5083 5997 5109
rect 5997 5083 6023 5109
rect 6023 5083 6024 5109
rect 5996 5082 6024 5083
rect 6048 5109 6076 5110
rect 6048 5083 6049 5109
rect 6049 5083 6075 5109
rect 6075 5083 6076 5109
rect 6048 5082 6076 5083
rect 6100 5109 6128 5110
rect 6100 5083 6101 5109
rect 6101 5083 6127 5109
rect 6127 5083 6128 5109
rect 6100 5082 6128 5083
rect 854 4857 882 4858
rect 854 4831 855 4857
rect 855 4831 881 4857
rect 881 4831 882 4857
rect 854 4830 882 4831
rect 1246 4857 1274 4858
rect 1246 4831 1247 4857
rect 1247 4831 1273 4857
rect 1273 4831 1274 4857
rect 1246 4830 1274 4831
rect 1022 4801 1050 4802
rect 1022 4775 1023 4801
rect 1023 4775 1049 4801
rect 1049 4775 1050 4801
rect 1022 4774 1050 4775
rect 6958 4774 6986 4802
rect 2762 4717 2790 4718
rect 2762 4691 2763 4717
rect 2763 4691 2789 4717
rect 2789 4691 2790 4717
rect 2762 4690 2790 4691
rect 2814 4717 2842 4718
rect 2814 4691 2815 4717
rect 2815 4691 2841 4717
rect 2841 4691 2842 4717
rect 2814 4690 2842 4691
rect 2866 4717 2894 4718
rect 2866 4691 2867 4717
rect 2867 4691 2893 4717
rect 2893 4691 2894 4717
rect 2866 4690 2894 4691
rect 4918 4717 4946 4718
rect 4918 4691 4919 4717
rect 4919 4691 4945 4717
rect 4945 4691 4946 4717
rect 4918 4690 4946 4691
rect 4970 4717 4998 4718
rect 4970 4691 4971 4717
rect 4971 4691 4997 4717
rect 4997 4691 4998 4717
rect 4970 4690 4998 4691
rect 5022 4717 5050 4718
rect 5022 4691 5023 4717
rect 5023 4691 5049 4717
rect 5049 4691 5050 4717
rect 5022 4690 5050 4691
rect 7350 4801 7378 4802
rect 7350 4775 7351 4801
rect 7351 4775 7377 4801
rect 7377 4775 7378 4801
rect 7350 4774 7378 4775
rect 7074 4717 7102 4718
rect 7074 4691 7075 4717
rect 7075 4691 7101 4717
rect 7101 4691 7102 4717
rect 7074 4690 7102 4691
rect 7126 4717 7154 4718
rect 7126 4691 7127 4717
rect 7127 4691 7153 4717
rect 7153 4691 7154 4717
rect 7126 4690 7154 4691
rect 7178 4717 7206 4718
rect 7178 4691 7179 4717
rect 7179 4691 7205 4717
rect 7205 4691 7206 4717
rect 7178 4690 7206 4691
rect 6958 4550 6986 4578
rect 854 4494 882 4522
rect 1684 4325 1712 4326
rect 1684 4299 1685 4325
rect 1685 4299 1711 4325
rect 1711 4299 1712 4325
rect 1684 4298 1712 4299
rect 1736 4325 1764 4326
rect 1736 4299 1737 4325
rect 1737 4299 1763 4325
rect 1763 4299 1764 4325
rect 1736 4298 1764 4299
rect 1788 4325 1816 4326
rect 1788 4299 1789 4325
rect 1789 4299 1815 4325
rect 1815 4299 1816 4325
rect 1788 4298 1816 4299
rect 3840 4325 3868 4326
rect 3840 4299 3841 4325
rect 3841 4299 3867 4325
rect 3867 4299 3868 4325
rect 3840 4298 3868 4299
rect 3892 4325 3920 4326
rect 3892 4299 3893 4325
rect 3893 4299 3919 4325
rect 3919 4299 3920 4325
rect 3892 4298 3920 4299
rect 3944 4325 3972 4326
rect 3944 4299 3945 4325
rect 3945 4299 3971 4325
rect 3971 4299 3972 4325
rect 3944 4298 3972 4299
rect 5996 4325 6024 4326
rect 5996 4299 5997 4325
rect 5997 4299 6023 4325
rect 6023 4299 6024 4325
rect 5996 4298 6024 4299
rect 6048 4325 6076 4326
rect 6048 4299 6049 4325
rect 6049 4299 6075 4325
rect 6075 4299 6076 4325
rect 6048 4298 6076 4299
rect 6100 4325 6128 4326
rect 6100 4299 6101 4325
rect 6101 4299 6127 4325
rect 6127 4299 6128 4325
rect 6100 4298 6128 4299
rect 7910 7601 7938 7602
rect 7910 7575 7911 7601
rect 7911 7575 7937 7601
rect 7937 7575 7938 7601
rect 7910 7574 7938 7575
rect 7574 4774 7602 4802
rect 1078 4046 1106 4074
rect 1022 3793 1050 3794
rect 1022 3767 1023 3793
rect 1023 3767 1049 3793
rect 1049 3767 1050 3793
rect 1022 3766 1050 3767
rect 854 3598 882 3626
rect 7294 4073 7322 4074
rect 7294 4047 7295 4073
rect 7295 4047 7321 4073
rect 7321 4047 7322 4073
rect 7294 4046 7322 4047
rect 7126 4017 7154 4018
rect 7126 3991 7127 4017
rect 7127 3991 7153 4017
rect 7153 3991 7154 4017
rect 7126 3990 7154 3991
rect 2762 3933 2790 3934
rect 2762 3907 2763 3933
rect 2763 3907 2789 3933
rect 2789 3907 2790 3933
rect 2762 3906 2790 3907
rect 2814 3933 2842 3934
rect 2814 3907 2815 3933
rect 2815 3907 2841 3933
rect 2841 3907 2842 3933
rect 2814 3906 2842 3907
rect 2866 3933 2894 3934
rect 2866 3907 2867 3933
rect 2867 3907 2893 3933
rect 2893 3907 2894 3933
rect 2866 3906 2894 3907
rect 4918 3933 4946 3934
rect 4918 3907 4919 3933
rect 4919 3907 4945 3933
rect 4945 3907 4946 3933
rect 4918 3906 4946 3907
rect 4970 3933 4998 3934
rect 4970 3907 4971 3933
rect 4971 3907 4997 3933
rect 4997 3907 4998 3933
rect 4970 3906 4998 3907
rect 5022 3933 5050 3934
rect 5022 3907 5023 3933
rect 5023 3907 5049 3933
rect 5049 3907 5050 3933
rect 5022 3906 5050 3907
rect 7074 3933 7102 3934
rect 7074 3907 7075 3933
rect 7075 3907 7101 3933
rect 7101 3907 7102 3933
rect 7074 3906 7102 3907
rect 7126 3933 7154 3934
rect 7126 3907 7127 3933
rect 7127 3907 7153 3933
rect 7153 3907 7154 3933
rect 7126 3906 7154 3907
rect 7178 3933 7206 3934
rect 7178 3907 7179 3933
rect 7179 3907 7205 3933
rect 7205 3907 7206 3933
rect 7178 3906 7206 3907
rect 7014 3766 7042 3794
rect 1246 3598 1274 3626
rect 1684 3541 1712 3542
rect 1684 3515 1685 3541
rect 1685 3515 1711 3541
rect 1711 3515 1712 3541
rect 1684 3514 1712 3515
rect 1736 3541 1764 3542
rect 1736 3515 1737 3541
rect 1737 3515 1763 3541
rect 1763 3515 1764 3541
rect 1736 3514 1764 3515
rect 1788 3541 1816 3542
rect 1788 3515 1789 3541
rect 1789 3515 1815 3541
rect 1815 3515 1816 3541
rect 1788 3514 1816 3515
rect 3840 3541 3868 3542
rect 3840 3515 3841 3541
rect 3841 3515 3867 3541
rect 3867 3515 3868 3541
rect 3840 3514 3868 3515
rect 3892 3541 3920 3542
rect 3892 3515 3893 3541
rect 3893 3515 3919 3541
rect 3919 3515 3920 3541
rect 3892 3514 3920 3515
rect 3944 3541 3972 3542
rect 3944 3515 3945 3541
rect 3945 3515 3971 3541
rect 3971 3515 3972 3541
rect 3944 3514 3972 3515
rect 5996 3541 6024 3542
rect 5996 3515 5997 3541
rect 5997 3515 6023 3541
rect 6023 3515 6024 3541
rect 5996 3514 6024 3515
rect 6048 3541 6076 3542
rect 6048 3515 6049 3541
rect 6049 3515 6075 3541
rect 6075 3515 6076 3541
rect 6048 3514 6076 3515
rect 6100 3541 6128 3542
rect 6100 3515 6101 3541
rect 6101 3515 6127 3541
rect 6127 3515 6128 3541
rect 6100 3514 6128 3515
rect 1078 3206 1106 3234
rect 854 2702 882 2730
rect 2762 3149 2790 3150
rect 2762 3123 2763 3149
rect 2763 3123 2789 3149
rect 2789 3123 2790 3149
rect 2762 3122 2790 3123
rect 2814 3149 2842 3150
rect 2814 3123 2815 3149
rect 2815 3123 2841 3149
rect 2841 3123 2842 3149
rect 2814 3122 2842 3123
rect 2866 3149 2894 3150
rect 2866 3123 2867 3149
rect 2867 3123 2893 3149
rect 2893 3123 2894 3149
rect 2866 3122 2894 3123
rect 4918 3149 4946 3150
rect 4918 3123 4919 3149
rect 4919 3123 4945 3149
rect 4945 3123 4946 3149
rect 4918 3122 4946 3123
rect 4970 3149 4998 3150
rect 4970 3123 4971 3149
rect 4971 3123 4997 3149
rect 4997 3123 4998 3149
rect 4970 3122 4998 3123
rect 5022 3149 5050 3150
rect 5022 3123 5023 3149
rect 5023 3123 5049 3149
rect 5049 3123 5050 3149
rect 5022 3122 5050 3123
rect 7074 3149 7102 3150
rect 7074 3123 7075 3149
rect 7075 3123 7101 3149
rect 7101 3123 7102 3149
rect 7074 3122 7102 3123
rect 7126 3149 7154 3150
rect 7126 3123 7127 3149
rect 7127 3123 7153 3149
rect 7153 3123 7154 3149
rect 7126 3122 7154 3123
rect 7178 3149 7206 3150
rect 7178 3123 7179 3149
rect 7179 3123 7205 3149
rect 7205 3123 7206 3149
rect 7178 3122 7206 3123
rect 7462 3990 7490 4018
rect 7910 3374 7938 3402
rect 7630 3233 7658 3234
rect 7630 3207 7631 3233
rect 7631 3207 7657 3233
rect 7657 3207 7658 3233
rect 7630 3206 7658 3207
rect 7686 2982 7714 3010
rect 1246 2702 1274 2730
rect 1684 2757 1712 2758
rect 1684 2731 1685 2757
rect 1685 2731 1711 2757
rect 1711 2731 1712 2757
rect 1684 2730 1712 2731
rect 1736 2757 1764 2758
rect 1736 2731 1737 2757
rect 1737 2731 1763 2757
rect 1763 2731 1764 2757
rect 1736 2730 1764 2731
rect 1788 2757 1816 2758
rect 1788 2731 1789 2757
rect 1789 2731 1815 2757
rect 1815 2731 1816 2757
rect 1788 2730 1816 2731
rect 3840 2757 3868 2758
rect 3840 2731 3841 2757
rect 3841 2731 3867 2757
rect 3867 2731 3868 2757
rect 3840 2730 3868 2731
rect 3892 2757 3920 2758
rect 3892 2731 3893 2757
rect 3893 2731 3919 2757
rect 3919 2731 3920 2757
rect 3892 2730 3920 2731
rect 3944 2757 3972 2758
rect 3944 2731 3945 2757
rect 3945 2731 3971 2757
rect 3971 2731 3972 2757
rect 3944 2730 3972 2731
rect 5996 2757 6024 2758
rect 5996 2731 5997 2757
rect 5997 2731 6023 2757
rect 6023 2731 6024 2757
rect 5996 2730 6024 2731
rect 6048 2757 6076 2758
rect 6048 2731 6049 2757
rect 6049 2731 6075 2757
rect 6075 2731 6076 2757
rect 6048 2730 6076 2731
rect 6100 2757 6128 2758
rect 6100 2731 6101 2757
rect 6101 2731 6127 2757
rect 6127 2731 6128 2757
rect 6100 2730 6128 2731
rect 2762 2365 2790 2366
rect 2762 2339 2763 2365
rect 2763 2339 2789 2365
rect 2789 2339 2790 2365
rect 2762 2338 2790 2339
rect 2814 2365 2842 2366
rect 2814 2339 2815 2365
rect 2815 2339 2841 2365
rect 2841 2339 2842 2365
rect 2814 2338 2842 2339
rect 2866 2365 2894 2366
rect 2866 2339 2867 2365
rect 2867 2339 2893 2365
rect 2893 2339 2894 2365
rect 2866 2338 2894 2339
rect 4918 2365 4946 2366
rect 4918 2339 4919 2365
rect 4919 2339 4945 2365
rect 4945 2339 4946 2365
rect 4918 2338 4946 2339
rect 4970 2365 4998 2366
rect 4970 2339 4971 2365
rect 4971 2339 4997 2365
rect 4997 2339 4998 2365
rect 4970 2338 4998 2339
rect 5022 2365 5050 2366
rect 5022 2339 5023 2365
rect 5023 2339 5049 2365
rect 5049 2339 5050 2365
rect 5022 2338 5050 2339
rect 7074 2365 7102 2366
rect 7074 2339 7075 2365
rect 7075 2339 7101 2365
rect 7101 2339 7102 2365
rect 7074 2338 7102 2339
rect 7126 2365 7154 2366
rect 7126 2339 7127 2365
rect 7127 2339 7153 2365
rect 7153 2339 7154 2365
rect 7126 2338 7154 2339
rect 7178 2365 7206 2366
rect 7178 2339 7179 2365
rect 7179 2339 7205 2365
rect 7205 2339 7206 2365
rect 7178 2338 7206 2339
rect 6958 2169 6986 2170
rect 6958 2143 6959 2169
rect 6959 2143 6985 2169
rect 6985 2143 6986 2169
rect 6958 2142 6986 2143
rect 854 2086 882 2114
rect 1246 2113 1274 2114
rect 1246 2087 1247 2113
rect 1247 2087 1273 2113
rect 1273 2087 1274 2113
rect 1246 2086 1274 2087
rect 1684 1973 1712 1974
rect 1684 1947 1685 1973
rect 1685 1947 1711 1973
rect 1711 1947 1712 1973
rect 1684 1946 1712 1947
rect 1736 1973 1764 1974
rect 1736 1947 1737 1973
rect 1737 1947 1763 1973
rect 1763 1947 1764 1973
rect 1736 1946 1764 1947
rect 1788 1973 1816 1974
rect 1788 1947 1789 1973
rect 1789 1947 1815 1973
rect 1815 1947 1816 1973
rect 1788 1946 1816 1947
rect 3840 1973 3868 1974
rect 3840 1947 3841 1973
rect 3841 1947 3867 1973
rect 3867 1947 3868 1973
rect 3840 1946 3868 1947
rect 3892 1973 3920 1974
rect 3892 1947 3893 1973
rect 3893 1947 3919 1973
rect 3919 1947 3920 1973
rect 3892 1946 3920 1947
rect 3944 1973 3972 1974
rect 3944 1947 3945 1973
rect 3945 1947 3971 1973
rect 3971 1947 3972 1973
rect 3944 1946 3972 1947
rect 5996 1973 6024 1974
rect 5996 1947 5997 1973
rect 5997 1947 6023 1973
rect 6023 1947 6024 1973
rect 5996 1946 6024 1947
rect 6048 1973 6076 1974
rect 6048 1947 6049 1973
rect 6049 1947 6075 1973
rect 6075 1947 6076 1973
rect 6048 1946 6076 1947
rect 6100 1973 6128 1974
rect 6100 1947 6101 1973
rect 6101 1947 6127 1973
rect 6127 1947 6128 1973
rect 6100 1946 6128 1947
rect 854 1806 882 1834
rect 1022 1806 1050 1834
rect 6286 1777 6314 1778
rect 6286 1751 6287 1777
rect 6287 1751 6313 1777
rect 6313 1751 6314 1777
rect 6286 1750 6314 1751
rect 854 1638 882 1666
rect 1246 1638 1274 1666
rect 2762 1581 2790 1582
rect 2762 1555 2763 1581
rect 2763 1555 2789 1581
rect 2789 1555 2790 1581
rect 2762 1554 2790 1555
rect 2814 1581 2842 1582
rect 2814 1555 2815 1581
rect 2815 1555 2841 1581
rect 2841 1555 2842 1581
rect 2814 1554 2842 1555
rect 2866 1581 2894 1582
rect 2866 1555 2867 1581
rect 2867 1555 2893 1581
rect 2893 1555 2894 1581
rect 2866 1554 2894 1555
rect 4918 1581 4946 1582
rect 4918 1555 4919 1581
rect 4919 1555 4945 1581
rect 4945 1555 4946 1581
rect 4918 1554 4946 1555
rect 4970 1581 4998 1582
rect 4970 1555 4971 1581
rect 4971 1555 4997 1581
rect 4997 1555 4998 1581
rect 4970 1554 4998 1555
rect 5022 1581 5050 1582
rect 5022 1555 5023 1581
rect 5023 1555 5049 1581
rect 5049 1555 5050 1581
rect 5022 1554 5050 1555
rect 5782 1134 5810 1162
rect 854 910 882 938
rect 7910 2478 7938 2506
rect 8470 7937 8498 7938
rect 8470 7911 8471 7937
rect 8471 7911 8497 7937
rect 8497 7911 8498 7937
rect 8470 7910 8498 7911
rect 8806 8022 8834 8050
rect 8918 7966 8946 7994
rect 8582 7742 8610 7770
rect 8358 7686 8386 7714
rect 8152 7461 8180 7462
rect 8152 7435 8153 7461
rect 8153 7435 8179 7461
rect 8179 7435 8180 7461
rect 8152 7434 8180 7435
rect 8204 7461 8232 7462
rect 8204 7435 8205 7461
rect 8205 7435 8231 7461
rect 8231 7435 8232 7461
rect 8204 7434 8232 7435
rect 8256 7461 8284 7462
rect 8256 7435 8257 7461
rect 8257 7435 8283 7461
rect 8283 7435 8284 7461
rect 8256 7434 8284 7435
rect 8694 7713 8722 7714
rect 8694 7687 8695 7713
rect 8695 7687 8721 7713
rect 8721 7687 8722 7713
rect 8694 7686 8722 7687
rect 9230 7853 9258 7854
rect 9230 7827 9231 7853
rect 9231 7827 9257 7853
rect 9257 7827 9258 7853
rect 9230 7826 9258 7827
rect 9282 7853 9310 7854
rect 9282 7827 9283 7853
rect 9283 7827 9309 7853
rect 9309 7827 9310 7853
rect 9282 7826 9310 7827
rect 9334 7853 9362 7854
rect 9334 7827 9335 7853
rect 9335 7827 9361 7853
rect 9361 7827 9362 7853
rect 9334 7826 9362 7827
rect 8582 7153 8610 7154
rect 8582 7127 8583 7153
rect 8583 7127 8609 7153
rect 8609 7127 8610 7153
rect 8582 7126 8610 7127
rect 8806 7238 8834 7266
rect 8470 6734 8498 6762
rect 8152 6677 8180 6678
rect 8152 6651 8153 6677
rect 8153 6651 8179 6677
rect 8179 6651 8180 6677
rect 8152 6650 8180 6651
rect 8204 6677 8232 6678
rect 8204 6651 8205 6677
rect 8205 6651 8231 6677
rect 8231 6651 8232 6677
rect 8204 6650 8232 6651
rect 8256 6677 8284 6678
rect 8256 6651 8257 6677
rect 8257 6651 8283 6677
rect 8283 6651 8284 6677
rect 8256 6650 8284 6651
rect 7966 2254 7994 2282
rect 8078 5950 8106 5978
rect 8152 5893 8180 5894
rect 8152 5867 8153 5893
rect 8153 5867 8179 5893
rect 8179 5867 8180 5893
rect 8152 5866 8180 5867
rect 8204 5893 8232 5894
rect 8204 5867 8205 5893
rect 8205 5867 8231 5893
rect 8231 5867 8232 5893
rect 8204 5866 8232 5867
rect 8256 5893 8284 5894
rect 8256 5867 8257 5893
rect 8257 5867 8283 5893
rect 8283 5867 8284 5893
rect 8256 5866 8284 5867
rect 8302 5193 8330 5194
rect 8302 5167 8303 5193
rect 8303 5167 8329 5193
rect 8329 5167 8330 5193
rect 8302 5166 8330 5167
rect 8152 5109 8180 5110
rect 8152 5083 8153 5109
rect 8153 5083 8179 5109
rect 8179 5083 8180 5109
rect 8152 5082 8180 5083
rect 8204 5109 8232 5110
rect 8204 5083 8205 5109
rect 8205 5083 8231 5109
rect 8231 5083 8232 5109
rect 8204 5082 8232 5083
rect 8256 5109 8284 5110
rect 8256 5083 8257 5109
rect 8257 5083 8283 5109
rect 8283 5083 8284 5109
rect 8256 5082 8284 5083
rect 8152 4325 8180 4326
rect 8152 4299 8153 4325
rect 8153 4299 8179 4325
rect 8179 4299 8180 4325
rect 8152 4298 8180 4299
rect 8204 4325 8232 4326
rect 8204 4299 8205 4325
rect 8205 4299 8231 4325
rect 8231 4299 8232 4325
rect 8204 4298 8232 4299
rect 8256 4325 8284 4326
rect 8256 4299 8257 4325
rect 8257 4299 8283 4325
rect 8283 4299 8284 4325
rect 8256 4298 8284 4299
rect 8358 4270 8386 4298
rect 8582 6537 8610 6538
rect 8582 6511 8583 6537
rect 8583 6511 8609 6537
rect 8609 6511 8610 6537
rect 8582 6510 8610 6511
rect 8750 6398 8778 6426
rect 8694 5977 8722 5978
rect 8694 5951 8695 5977
rect 8695 5951 8721 5977
rect 8721 5951 8722 5977
rect 8694 5950 8722 5951
rect 8694 5670 8722 5698
rect 8582 5446 8610 5474
rect 8694 5361 8722 5362
rect 8694 5335 8695 5361
rect 8695 5335 8721 5361
rect 8721 5335 8722 5361
rect 8694 5334 8722 5335
rect 9086 7238 9114 7266
rect 9030 6761 9058 6762
rect 9030 6735 9031 6761
rect 9031 6735 9057 6761
rect 9057 6735 9058 6761
rect 9030 6734 9058 6735
rect 8974 6062 9002 6090
rect 9086 5361 9114 5362
rect 9086 5335 9087 5361
rect 9087 5335 9113 5361
rect 9113 5335 9114 5361
rect 9086 5334 9114 5335
rect 8582 4606 8610 4634
rect 8862 4577 8890 4578
rect 8862 4551 8863 4577
rect 8863 4551 8889 4577
rect 8889 4551 8890 4577
rect 8862 4550 8890 4551
rect 8152 3541 8180 3542
rect 8152 3515 8153 3541
rect 8153 3515 8179 3541
rect 8179 3515 8180 3541
rect 8152 3514 8180 3515
rect 8204 3541 8232 3542
rect 8204 3515 8205 3541
rect 8205 3515 8231 3541
rect 8231 3515 8232 3541
rect 8204 3514 8232 3515
rect 8256 3541 8284 3542
rect 8256 3515 8257 3541
rect 8257 3515 8283 3541
rect 8283 3515 8284 3541
rect 8256 3514 8284 3515
rect 8358 3038 8386 3066
rect 8358 2926 8386 2954
rect 8152 2757 8180 2758
rect 8152 2731 8153 2757
rect 8153 2731 8179 2757
rect 8179 2731 8180 2757
rect 8152 2730 8180 2731
rect 8204 2757 8232 2758
rect 8204 2731 8205 2757
rect 8205 2731 8231 2757
rect 8231 2731 8232 2757
rect 8204 2730 8232 2731
rect 8256 2757 8284 2758
rect 8256 2731 8257 2757
rect 8257 2731 8283 2757
rect 8283 2731 8284 2757
rect 8256 2730 8284 2731
rect 7518 2030 7546 2058
rect 8152 1973 8180 1974
rect 8152 1947 8153 1973
rect 8153 1947 8179 1973
rect 8179 1947 8180 1973
rect 8152 1946 8180 1947
rect 8204 1973 8232 1974
rect 8204 1947 8205 1973
rect 8205 1947 8231 1973
rect 8231 1947 8232 1973
rect 8204 1946 8232 1947
rect 8256 1973 8284 1974
rect 8256 1947 8257 1973
rect 8257 1947 8283 1973
rect 8283 1947 8284 1973
rect 8256 1946 8284 1947
rect 8806 4046 8834 4074
rect 8582 3710 8610 3738
rect 8918 3990 8946 4018
rect 8694 3065 8722 3066
rect 8694 3039 8695 3065
rect 8695 3039 8721 3065
rect 8721 3039 8722 3065
rect 8694 3038 8722 3039
rect 8750 3009 8778 3010
rect 8750 2983 8751 3009
rect 8751 2983 8777 3009
rect 8777 2983 8778 3009
rect 8750 2982 8778 2983
rect 9086 3206 9114 3234
rect 8694 2281 8722 2282
rect 8694 2255 8695 2281
rect 8695 2255 8721 2281
rect 8721 2255 8722 2281
rect 8694 2254 8722 2255
rect 8470 2142 8498 2170
rect 8526 1833 8554 1834
rect 8526 1807 8527 1833
rect 8527 1807 8553 1833
rect 8553 1807 8554 1833
rect 8526 1806 8554 1807
rect 8806 1806 8834 1834
rect 9230 7069 9258 7070
rect 9230 7043 9231 7069
rect 9231 7043 9257 7069
rect 9257 7043 9258 7069
rect 9230 7042 9258 7043
rect 9282 7069 9310 7070
rect 9282 7043 9283 7069
rect 9283 7043 9309 7069
rect 9309 7043 9310 7069
rect 9282 7042 9310 7043
rect 9334 7069 9362 7070
rect 9334 7043 9335 7069
rect 9335 7043 9361 7069
rect 9361 7043 9362 7069
rect 9334 7042 9362 7043
rect 9230 6285 9258 6286
rect 9230 6259 9231 6285
rect 9231 6259 9257 6285
rect 9257 6259 9258 6285
rect 9230 6258 9258 6259
rect 9282 6285 9310 6286
rect 9282 6259 9283 6285
rect 9283 6259 9309 6285
rect 9309 6259 9310 6285
rect 9282 6258 9310 6259
rect 9334 6285 9362 6286
rect 9334 6259 9335 6285
rect 9335 6259 9361 6285
rect 9361 6259 9362 6285
rect 9334 6258 9362 6259
rect 9230 5501 9258 5502
rect 9230 5475 9231 5501
rect 9231 5475 9257 5501
rect 9257 5475 9258 5501
rect 9230 5474 9258 5475
rect 9282 5501 9310 5502
rect 9282 5475 9283 5501
rect 9283 5475 9309 5501
rect 9309 5475 9310 5501
rect 9282 5474 9310 5475
rect 9334 5501 9362 5502
rect 9334 5475 9335 5501
rect 9335 5475 9361 5501
rect 9361 5475 9362 5501
rect 9334 5474 9362 5475
rect 9230 4717 9258 4718
rect 9230 4691 9231 4717
rect 9231 4691 9257 4717
rect 9257 4691 9258 4717
rect 9230 4690 9258 4691
rect 9282 4717 9310 4718
rect 9282 4691 9283 4717
rect 9283 4691 9309 4717
rect 9309 4691 9310 4717
rect 9282 4690 9310 4691
rect 9334 4717 9362 4718
rect 9334 4691 9335 4717
rect 9335 4691 9361 4717
rect 9361 4691 9362 4717
rect 9334 4690 9362 4691
rect 9230 3933 9258 3934
rect 9230 3907 9231 3933
rect 9231 3907 9257 3933
rect 9257 3907 9258 3933
rect 9230 3906 9258 3907
rect 9282 3933 9310 3934
rect 9282 3907 9283 3933
rect 9283 3907 9309 3933
rect 9309 3907 9310 3933
rect 9282 3906 9310 3907
rect 9334 3933 9362 3934
rect 9334 3907 9335 3933
rect 9335 3907 9361 3933
rect 9361 3907 9362 3933
rect 9334 3906 9362 3907
rect 9230 3149 9258 3150
rect 9230 3123 9231 3149
rect 9231 3123 9257 3149
rect 9257 3123 9258 3149
rect 9230 3122 9258 3123
rect 9282 3149 9310 3150
rect 9282 3123 9283 3149
rect 9283 3123 9309 3149
rect 9309 3123 9310 3149
rect 9282 3122 9310 3123
rect 9334 3149 9362 3150
rect 9334 3123 9335 3149
rect 9335 3123 9361 3149
rect 9361 3123 9362 3149
rect 9334 3122 9362 3123
rect 9230 2365 9258 2366
rect 9230 2339 9231 2365
rect 9231 2339 9257 2365
rect 9257 2339 9258 2365
rect 9230 2338 9258 2339
rect 9282 2365 9310 2366
rect 9282 2339 9283 2365
rect 9283 2339 9309 2365
rect 9309 2339 9310 2365
rect 9282 2338 9310 2339
rect 9334 2365 9362 2366
rect 9334 2339 9335 2365
rect 9335 2339 9361 2365
rect 9361 2339 9362 2365
rect 9334 2338 9362 2339
rect 9142 1750 9170 1778
rect 7518 1638 7546 1666
rect 7074 1581 7102 1582
rect 7074 1555 7075 1581
rect 7075 1555 7101 1581
rect 7101 1555 7102 1581
rect 7074 1554 7102 1555
rect 7126 1581 7154 1582
rect 7126 1555 7127 1581
rect 7127 1555 7153 1581
rect 7153 1555 7154 1581
rect 7126 1554 7154 1555
rect 7178 1581 7206 1582
rect 7178 1555 7179 1581
rect 7179 1555 7205 1581
rect 7205 1555 7206 1581
rect 7178 1554 7206 1555
rect 9230 1581 9258 1582
rect 9230 1555 9231 1581
rect 9231 1555 9257 1581
rect 9257 1555 9258 1581
rect 9230 1554 9258 1555
rect 9282 1581 9310 1582
rect 9282 1555 9283 1581
rect 9283 1555 9309 1581
rect 9309 1555 9310 1581
rect 9282 1554 9310 1555
rect 9334 1581 9362 1582
rect 9334 1555 9335 1581
rect 9335 1555 9361 1581
rect 9361 1555 9362 1581
rect 9334 1554 9362 1555
rect 6454 854 6482 882
<< metal3 >>
rect 9600 9226 10000 9240
rect 7457 9198 7462 9226
rect 7490 9198 10000 9226
rect 9600 9184 10000 9198
rect 0 9002 400 9016
rect 0 8974 854 9002
rect 882 8974 887 9002
rect 0 8960 400 8974
rect 9600 8778 10000 8792
rect 5777 8750 5782 8778
rect 5810 8750 10000 8778
rect 9600 8736 10000 8750
rect 9600 8330 10000 8344
rect 6449 8302 6454 8330
rect 6482 8302 10000 8330
rect 9600 8288 10000 8302
rect 1679 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1821 8246
rect 3835 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3977 8246
rect 5991 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6133 8246
rect 8147 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8289 8246
rect 0 8106 400 8120
rect 0 8078 1190 8106
rect 1218 8078 1223 8106
rect 0 8064 400 8078
rect 849 8022 854 8050
rect 882 8022 1582 8050
rect 1610 8022 1615 8050
rect 6281 8022 6286 8050
rect 6314 8022 8806 8050
rect 8834 8022 8839 8050
rect 4186 7966 8918 7994
rect 8946 7966 8951 7994
rect 4186 7938 4214 7966
rect 1017 7910 1022 7938
rect 1050 7910 4214 7938
rect 6953 7910 6958 7938
rect 6986 7910 8470 7938
rect 8498 7910 8503 7938
rect 8582 7910 9450 7938
rect 8582 7882 8610 7910
rect 7793 7854 7798 7882
rect 7826 7854 8610 7882
rect 9422 7882 9450 7910
rect 9600 7882 10000 7896
rect 9422 7854 10000 7882
rect 2757 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2899 7854
rect 4913 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5055 7854
rect 7069 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7211 7854
rect 9225 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9367 7854
rect 9600 7840 10000 7854
rect 1353 7742 1358 7770
rect 1386 7742 7630 7770
rect 7658 7742 8582 7770
rect 8610 7742 8615 7770
rect 8353 7686 8358 7714
rect 8386 7686 8694 7714
rect 8722 7686 8727 7714
rect 7905 7574 7910 7602
rect 7938 7574 7943 7602
rect 7910 7546 7938 7574
rect 7910 7518 8442 7546
rect 1679 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1821 7462
rect 3835 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3977 7462
rect 5991 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6133 7462
rect 8147 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8289 7462
rect 8414 7434 8442 7518
rect 9600 7434 10000 7448
rect 8414 7406 10000 7434
rect 9600 7392 10000 7406
rect 1017 7238 1022 7266
rect 1050 7238 8806 7266
rect 8834 7238 9086 7266
rect 9114 7238 9119 7266
rect 0 7210 400 7224
rect 0 7182 854 7210
rect 882 7182 1246 7210
rect 1274 7182 1279 7210
rect 0 7168 400 7182
rect 8577 7126 8582 7154
rect 8610 7126 8615 7154
rect 2757 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2899 7070
rect 4913 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5055 7070
rect 7069 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7211 7070
rect 8582 6986 8610 7126
rect 9225 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9367 7070
rect 9600 6986 10000 7000
rect 8582 6958 10000 6986
rect 9600 6944 10000 6958
rect 8465 6734 8470 6762
rect 8498 6734 9030 6762
rect 9058 6734 9063 6762
rect 1679 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1821 6678
rect 3835 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3977 6678
rect 5991 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6133 6678
rect 8147 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8289 6678
rect 9600 6538 10000 6552
rect 8577 6510 8582 6538
rect 8610 6510 10000 6538
rect 9600 6496 10000 6510
rect 1017 6398 1022 6426
rect 1050 6398 8750 6426
rect 8778 6398 8783 6426
rect 0 6314 400 6328
rect 0 6286 854 6314
rect 882 6286 1246 6314
rect 1274 6286 1279 6314
rect 0 6272 400 6286
rect 2757 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2899 6286
rect 4913 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5055 6286
rect 7069 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7211 6286
rect 9225 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9367 6286
rect 9600 6090 10000 6104
rect 8969 6062 8974 6090
rect 9002 6062 10000 6090
rect 9600 6048 10000 6062
rect 8073 5950 8078 5978
rect 8106 5950 8694 5978
rect 8722 5950 8727 5978
rect 1679 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1821 5894
rect 3835 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3977 5894
rect 5991 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6133 5894
rect 8147 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8289 5894
rect 1017 5670 1022 5698
rect 1050 5670 8694 5698
rect 8722 5670 8727 5698
rect 9600 5642 10000 5656
rect 8582 5614 10000 5642
rect 2757 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2899 5502
rect 4913 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5055 5502
rect 7069 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7211 5502
rect 8582 5474 8610 5614
rect 9600 5600 10000 5614
rect 9225 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9367 5502
rect 8577 5446 8582 5474
rect 8610 5446 8615 5474
rect 0 5418 400 5432
rect 0 5390 854 5418
rect 882 5390 1246 5418
rect 1274 5390 1279 5418
rect 0 5376 400 5390
rect 8689 5334 8694 5362
rect 8722 5334 9086 5362
rect 9114 5334 9119 5362
rect 9600 5194 10000 5208
rect 8297 5166 8302 5194
rect 8330 5166 10000 5194
rect 9600 5152 10000 5166
rect 1679 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1821 5110
rect 3835 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3977 5110
rect 5991 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6133 5110
rect 8147 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8289 5110
rect 849 4830 854 4858
rect 882 4830 1246 4858
rect 1274 4830 1279 4858
rect 1017 4774 1022 4802
rect 1050 4774 6958 4802
rect 6986 4774 6991 4802
rect 7345 4774 7350 4802
rect 7378 4774 7574 4802
rect 7602 4774 7607 4802
rect 9600 4746 10000 4760
rect 9422 4718 10000 4746
rect 2757 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2899 4718
rect 4913 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5055 4718
rect 7069 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7211 4718
rect 9225 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9367 4718
rect 9422 4634 9450 4718
rect 9600 4704 10000 4718
rect 8577 4606 8582 4634
rect 8610 4606 9450 4634
rect 6953 4550 6958 4578
rect 6986 4550 8862 4578
rect 8890 4550 8895 4578
rect 0 4522 400 4536
rect 0 4494 854 4522
rect 882 4494 887 4522
rect 0 4480 400 4494
rect 1679 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1821 4326
rect 3835 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3977 4326
rect 5991 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6133 4326
rect 8147 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8289 4326
rect 9600 4298 10000 4312
rect 8353 4270 8358 4298
rect 8386 4270 10000 4298
rect 9600 4256 10000 4270
rect 1073 4046 1078 4074
rect 1106 4046 7294 4074
rect 7322 4046 8806 4074
rect 8834 4046 8839 4074
rect 7121 3990 7126 4018
rect 7154 3990 7462 4018
rect 7490 3990 8918 4018
rect 8946 3990 8951 4018
rect 2757 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2899 3934
rect 4913 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5055 3934
rect 7069 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7211 3934
rect 9225 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9367 3934
rect 9600 3850 10000 3864
rect 8582 3822 10000 3850
rect 1017 3766 1022 3794
rect 1050 3766 7014 3794
rect 7042 3766 7047 3794
rect 8582 3738 8610 3822
rect 9600 3808 10000 3822
rect 8577 3710 8582 3738
rect 8610 3710 8615 3738
rect 0 3626 400 3640
rect 0 3598 854 3626
rect 882 3598 1246 3626
rect 1274 3598 1279 3626
rect 0 3584 400 3598
rect 1679 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1821 3542
rect 3835 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3977 3542
rect 5991 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6133 3542
rect 8147 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8289 3542
rect 9600 3402 10000 3416
rect 7905 3374 7910 3402
rect 7938 3374 10000 3402
rect 9600 3360 10000 3374
rect 1073 3206 1078 3234
rect 1106 3206 7630 3234
rect 7658 3206 9086 3234
rect 9114 3206 9119 3234
rect 2757 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2899 3150
rect 4913 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5055 3150
rect 7069 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7211 3150
rect 9225 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9367 3150
rect 8353 3038 8358 3066
rect 8386 3038 8694 3066
rect 8722 3038 8727 3066
rect 7681 2982 7686 3010
rect 7714 2982 8750 3010
rect 8778 2982 8783 3010
rect 9600 2954 10000 2968
rect 8353 2926 8358 2954
rect 8386 2926 10000 2954
rect 9600 2912 10000 2926
rect 0 2730 400 2744
rect 1679 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1821 2758
rect 3835 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3977 2758
rect 5991 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6133 2758
rect 8147 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8289 2758
rect 0 2702 854 2730
rect 882 2702 1246 2730
rect 1274 2702 1279 2730
rect 0 2688 400 2702
rect 9600 2506 10000 2520
rect 7905 2478 7910 2506
rect 7938 2478 10000 2506
rect 9600 2464 10000 2478
rect 2757 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2899 2366
rect 4913 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5055 2366
rect 7069 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7211 2366
rect 9225 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9367 2366
rect 7961 2254 7966 2282
rect 7994 2254 8694 2282
rect 8722 2254 8727 2282
rect 6953 2142 6958 2170
rect 6986 2142 8470 2170
rect 8498 2142 8503 2170
rect 849 2086 854 2114
rect 882 2086 1246 2114
rect 1274 2086 1279 2114
rect 9600 2058 10000 2072
rect 7513 2030 7518 2058
rect 7546 2030 10000 2058
rect 9600 2016 10000 2030
rect 1679 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1821 1974
rect 3835 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3977 1974
rect 5991 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6133 1974
rect 8147 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8289 1974
rect 0 1834 400 1848
rect 0 1806 854 1834
rect 882 1806 887 1834
rect 1017 1806 1022 1834
rect 1050 1806 8526 1834
rect 8554 1806 8806 1834
rect 8834 1806 8839 1834
rect 0 1792 400 1806
rect 6281 1750 6286 1778
rect 6314 1750 9142 1778
rect 9170 1750 9175 1778
rect 849 1638 854 1666
rect 882 1638 1246 1666
rect 1274 1638 1279 1666
rect 7513 1638 7518 1666
rect 7546 1638 9450 1666
rect 9422 1610 9450 1638
rect 9600 1610 10000 1624
rect 9422 1582 10000 1610
rect 2757 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2899 1582
rect 4913 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5055 1582
rect 7069 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7211 1582
rect 9225 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9367 1582
rect 9600 1568 10000 1582
rect 9600 1162 10000 1176
rect 5777 1134 5782 1162
rect 5810 1134 10000 1162
rect 9600 1120 10000 1134
rect 0 938 400 952
rect 0 910 854 938
rect 882 910 887 938
rect 0 896 400 910
rect 6449 854 6454 882
rect 6482 854 6762 882
rect 6734 714 6762 854
rect 9600 714 10000 728
rect 6734 686 10000 714
rect 9600 672 10000 686
<< via3 >>
rect 1684 8218 1712 8246
rect 1736 8218 1764 8246
rect 1788 8218 1816 8246
rect 3840 8218 3868 8246
rect 3892 8218 3920 8246
rect 3944 8218 3972 8246
rect 5996 8218 6024 8246
rect 6048 8218 6076 8246
rect 6100 8218 6128 8246
rect 8152 8218 8180 8246
rect 8204 8218 8232 8246
rect 8256 8218 8284 8246
rect 2762 7826 2790 7854
rect 2814 7826 2842 7854
rect 2866 7826 2894 7854
rect 4918 7826 4946 7854
rect 4970 7826 4998 7854
rect 5022 7826 5050 7854
rect 7074 7826 7102 7854
rect 7126 7826 7154 7854
rect 7178 7826 7206 7854
rect 9230 7826 9258 7854
rect 9282 7826 9310 7854
rect 9334 7826 9362 7854
rect 1684 7434 1712 7462
rect 1736 7434 1764 7462
rect 1788 7434 1816 7462
rect 3840 7434 3868 7462
rect 3892 7434 3920 7462
rect 3944 7434 3972 7462
rect 5996 7434 6024 7462
rect 6048 7434 6076 7462
rect 6100 7434 6128 7462
rect 8152 7434 8180 7462
rect 8204 7434 8232 7462
rect 8256 7434 8284 7462
rect 2762 7042 2790 7070
rect 2814 7042 2842 7070
rect 2866 7042 2894 7070
rect 4918 7042 4946 7070
rect 4970 7042 4998 7070
rect 5022 7042 5050 7070
rect 7074 7042 7102 7070
rect 7126 7042 7154 7070
rect 7178 7042 7206 7070
rect 9230 7042 9258 7070
rect 9282 7042 9310 7070
rect 9334 7042 9362 7070
rect 1684 6650 1712 6678
rect 1736 6650 1764 6678
rect 1788 6650 1816 6678
rect 3840 6650 3868 6678
rect 3892 6650 3920 6678
rect 3944 6650 3972 6678
rect 5996 6650 6024 6678
rect 6048 6650 6076 6678
rect 6100 6650 6128 6678
rect 8152 6650 8180 6678
rect 8204 6650 8232 6678
rect 8256 6650 8284 6678
rect 2762 6258 2790 6286
rect 2814 6258 2842 6286
rect 2866 6258 2894 6286
rect 4918 6258 4946 6286
rect 4970 6258 4998 6286
rect 5022 6258 5050 6286
rect 7074 6258 7102 6286
rect 7126 6258 7154 6286
rect 7178 6258 7206 6286
rect 9230 6258 9258 6286
rect 9282 6258 9310 6286
rect 9334 6258 9362 6286
rect 1684 5866 1712 5894
rect 1736 5866 1764 5894
rect 1788 5866 1816 5894
rect 3840 5866 3868 5894
rect 3892 5866 3920 5894
rect 3944 5866 3972 5894
rect 5996 5866 6024 5894
rect 6048 5866 6076 5894
rect 6100 5866 6128 5894
rect 8152 5866 8180 5894
rect 8204 5866 8232 5894
rect 8256 5866 8284 5894
rect 2762 5474 2790 5502
rect 2814 5474 2842 5502
rect 2866 5474 2894 5502
rect 4918 5474 4946 5502
rect 4970 5474 4998 5502
rect 5022 5474 5050 5502
rect 7074 5474 7102 5502
rect 7126 5474 7154 5502
rect 7178 5474 7206 5502
rect 9230 5474 9258 5502
rect 9282 5474 9310 5502
rect 9334 5474 9362 5502
rect 1684 5082 1712 5110
rect 1736 5082 1764 5110
rect 1788 5082 1816 5110
rect 3840 5082 3868 5110
rect 3892 5082 3920 5110
rect 3944 5082 3972 5110
rect 5996 5082 6024 5110
rect 6048 5082 6076 5110
rect 6100 5082 6128 5110
rect 8152 5082 8180 5110
rect 8204 5082 8232 5110
rect 8256 5082 8284 5110
rect 2762 4690 2790 4718
rect 2814 4690 2842 4718
rect 2866 4690 2894 4718
rect 4918 4690 4946 4718
rect 4970 4690 4998 4718
rect 5022 4690 5050 4718
rect 7074 4690 7102 4718
rect 7126 4690 7154 4718
rect 7178 4690 7206 4718
rect 9230 4690 9258 4718
rect 9282 4690 9310 4718
rect 9334 4690 9362 4718
rect 1684 4298 1712 4326
rect 1736 4298 1764 4326
rect 1788 4298 1816 4326
rect 3840 4298 3868 4326
rect 3892 4298 3920 4326
rect 3944 4298 3972 4326
rect 5996 4298 6024 4326
rect 6048 4298 6076 4326
rect 6100 4298 6128 4326
rect 8152 4298 8180 4326
rect 8204 4298 8232 4326
rect 8256 4298 8284 4326
rect 2762 3906 2790 3934
rect 2814 3906 2842 3934
rect 2866 3906 2894 3934
rect 4918 3906 4946 3934
rect 4970 3906 4998 3934
rect 5022 3906 5050 3934
rect 7074 3906 7102 3934
rect 7126 3906 7154 3934
rect 7178 3906 7206 3934
rect 9230 3906 9258 3934
rect 9282 3906 9310 3934
rect 9334 3906 9362 3934
rect 1684 3514 1712 3542
rect 1736 3514 1764 3542
rect 1788 3514 1816 3542
rect 3840 3514 3868 3542
rect 3892 3514 3920 3542
rect 3944 3514 3972 3542
rect 5996 3514 6024 3542
rect 6048 3514 6076 3542
rect 6100 3514 6128 3542
rect 8152 3514 8180 3542
rect 8204 3514 8232 3542
rect 8256 3514 8284 3542
rect 2762 3122 2790 3150
rect 2814 3122 2842 3150
rect 2866 3122 2894 3150
rect 4918 3122 4946 3150
rect 4970 3122 4998 3150
rect 5022 3122 5050 3150
rect 7074 3122 7102 3150
rect 7126 3122 7154 3150
rect 7178 3122 7206 3150
rect 9230 3122 9258 3150
rect 9282 3122 9310 3150
rect 9334 3122 9362 3150
rect 1684 2730 1712 2758
rect 1736 2730 1764 2758
rect 1788 2730 1816 2758
rect 3840 2730 3868 2758
rect 3892 2730 3920 2758
rect 3944 2730 3972 2758
rect 5996 2730 6024 2758
rect 6048 2730 6076 2758
rect 6100 2730 6128 2758
rect 8152 2730 8180 2758
rect 8204 2730 8232 2758
rect 8256 2730 8284 2758
rect 2762 2338 2790 2366
rect 2814 2338 2842 2366
rect 2866 2338 2894 2366
rect 4918 2338 4946 2366
rect 4970 2338 4998 2366
rect 5022 2338 5050 2366
rect 7074 2338 7102 2366
rect 7126 2338 7154 2366
rect 7178 2338 7206 2366
rect 9230 2338 9258 2366
rect 9282 2338 9310 2366
rect 9334 2338 9362 2366
rect 1684 1946 1712 1974
rect 1736 1946 1764 1974
rect 1788 1946 1816 1974
rect 3840 1946 3868 1974
rect 3892 1946 3920 1974
rect 3944 1946 3972 1974
rect 5996 1946 6024 1974
rect 6048 1946 6076 1974
rect 6100 1946 6128 1974
rect 8152 1946 8180 1974
rect 8204 1946 8232 1974
rect 8256 1946 8284 1974
rect 2762 1554 2790 1582
rect 2814 1554 2842 1582
rect 2866 1554 2894 1582
rect 4918 1554 4946 1582
rect 4970 1554 4998 1582
rect 5022 1554 5050 1582
rect 7074 1554 7102 1582
rect 7126 1554 7154 1582
rect 7178 1554 7206 1582
rect 9230 1554 9258 1582
rect 9282 1554 9310 1582
rect 9334 1554 9362 1582
<< metal4 >>
rect 1670 8246 1830 8262
rect 1670 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1830 8246
rect 1670 7462 1830 8218
rect 1670 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1830 7462
rect 1670 6678 1830 7434
rect 1670 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1830 6678
rect 1670 5894 1830 6650
rect 1670 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1830 5894
rect 1670 5110 1830 5866
rect 1670 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1830 5110
rect 1670 4326 1830 5082
rect 1670 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1830 4326
rect 1670 3542 1830 4298
rect 1670 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1830 3542
rect 1670 2758 1830 3514
rect 1670 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1830 2758
rect 1670 1974 1830 2730
rect 1670 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1830 1974
rect 1670 1538 1830 1946
rect 2748 7854 2908 8262
rect 2748 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2908 7854
rect 2748 7070 2908 7826
rect 2748 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2908 7070
rect 2748 6286 2908 7042
rect 2748 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2908 6286
rect 2748 5502 2908 6258
rect 2748 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2908 5502
rect 2748 4718 2908 5474
rect 2748 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2908 4718
rect 2748 3934 2908 4690
rect 2748 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2908 3934
rect 2748 3150 2908 3906
rect 2748 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2908 3150
rect 2748 2366 2908 3122
rect 2748 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2908 2366
rect 2748 1582 2908 2338
rect 2748 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2908 1582
rect 2748 1538 2908 1554
rect 3826 8246 3986 8262
rect 3826 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3986 8246
rect 3826 7462 3986 8218
rect 3826 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3986 7462
rect 3826 6678 3986 7434
rect 3826 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3986 6678
rect 3826 5894 3986 6650
rect 3826 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3986 5894
rect 3826 5110 3986 5866
rect 3826 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3986 5110
rect 3826 4326 3986 5082
rect 3826 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3986 4326
rect 3826 3542 3986 4298
rect 3826 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3986 3542
rect 3826 2758 3986 3514
rect 3826 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3986 2758
rect 3826 1974 3986 2730
rect 3826 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3986 1974
rect 3826 1538 3986 1946
rect 4904 7854 5064 8262
rect 4904 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5064 7854
rect 4904 7070 5064 7826
rect 4904 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5064 7070
rect 4904 6286 5064 7042
rect 4904 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5064 6286
rect 4904 5502 5064 6258
rect 4904 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5064 5502
rect 4904 4718 5064 5474
rect 4904 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5064 4718
rect 4904 3934 5064 4690
rect 4904 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5064 3934
rect 4904 3150 5064 3906
rect 4904 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5064 3150
rect 4904 2366 5064 3122
rect 4904 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5064 2366
rect 4904 1582 5064 2338
rect 4904 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5064 1582
rect 4904 1538 5064 1554
rect 5982 8246 6142 8262
rect 5982 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6142 8246
rect 5982 7462 6142 8218
rect 5982 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6142 7462
rect 5982 6678 6142 7434
rect 5982 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6142 6678
rect 5982 5894 6142 6650
rect 5982 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6142 5894
rect 5982 5110 6142 5866
rect 5982 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6142 5110
rect 5982 4326 6142 5082
rect 5982 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6142 4326
rect 5982 3542 6142 4298
rect 5982 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6142 3542
rect 5982 2758 6142 3514
rect 5982 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6142 2758
rect 5982 1974 6142 2730
rect 5982 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6142 1974
rect 5982 1538 6142 1946
rect 7060 7854 7220 8262
rect 7060 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7220 7854
rect 7060 7070 7220 7826
rect 7060 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7220 7070
rect 7060 6286 7220 7042
rect 7060 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7220 6286
rect 7060 5502 7220 6258
rect 7060 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7220 5502
rect 7060 4718 7220 5474
rect 7060 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7220 4718
rect 7060 3934 7220 4690
rect 7060 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7220 3934
rect 7060 3150 7220 3906
rect 7060 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7220 3150
rect 7060 2366 7220 3122
rect 7060 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7220 2366
rect 7060 1582 7220 2338
rect 7060 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7220 1582
rect 7060 1538 7220 1554
rect 8138 8246 8298 8262
rect 8138 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8298 8246
rect 8138 7462 8298 8218
rect 8138 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8298 7462
rect 8138 6678 8298 7434
rect 8138 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8298 6678
rect 8138 5894 8298 6650
rect 8138 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8298 5894
rect 8138 5110 8298 5866
rect 8138 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8298 5110
rect 8138 4326 8298 5082
rect 8138 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8298 4326
rect 8138 3542 8298 4298
rect 8138 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8298 3542
rect 8138 2758 8298 3514
rect 8138 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8298 2758
rect 8138 1974 8298 2730
rect 8138 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8298 1974
rect 8138 1538 8298 1946
rect 9216 7854 9376 8262
rect 9216 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9376 7854
rect 9216 7070 9376 7826
rect 9216 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9376 7070
rect 9216 6286 9376 7042
rect 9216 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9376 6286
rect 9216 5502 9376 6258
rect 9216 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9376 5502
rect 9216 4718 9376 5474
rect 9216 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9376 4718
rect 9216 3934 9376 4690
rect 9216 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9376 3934
rect 9216 3150 9376 3906
rect 9216 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9376 3150
rect 9216 2366 9376 3122
rect 9216 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9376 2366
rect 9216 1582 9376 2338
rect 9216 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9376 1582
rect 9216 1538 9376 1554
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _00_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 9184 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _01_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 8624 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _02_
timestamp 1694700623
transform -1 0 9184 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _03_
timestamp 1694700623
transform -1 0 7392 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _04_
timestamp 1694700623
transform 1 0 8848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _05_
timestamp 1694700623
transform -1 0 8848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _06_
timestamp 1694700623
transform -1 0 9184 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _07_
timestamp 1694700623
transform -1 0 8848 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _08_
timestamp 1694700623
transform -1 0 9184 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _09_
timestamp 1694700623
transform -1 0 7728 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _10_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 8960 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _11_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 7728 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _12_
timestamp 1694700623
transform -1 0 8960 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _13_
timestamp 1694700623
transform 1 0 7392 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _14_
timestamp 1694700623
transform -1 0 8960 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _15_
timestamp 1694700623
transform 1 0 8624 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _16_
timestamp 1694700623
transform -1 0 8960 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _17_
timestamp 1694700623
transform -1 0 8960 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _18_
timestamp 1694700623
transform -1 0 8736 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _19_
timestamp 1694700623
transform -1 0 9072 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__02__I pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 7616 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__04__I
timestamp 1694700623
transform 1 0 9072 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__05__I
timestamp 1694700623
transform -1 0 7728 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__06__I
timestamp 1694700623
transform -1 0 9072 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__11__I
timestamp 1694700623
transform -1 0 7392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__13__I
timestamp 1694700623
transform -1 0 7168 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__14__I
timestamp 1694700623
transform 1 0 6944 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__15__I
timestamp 1694700623
transform 1 0 9072 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1694700623
transform 1 0 1232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1694700623
transform 1 0 1232 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1694700623
transform 1 0 1232 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1694700623
transform 1 0 1232 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1694700623
transform 1 0 1232 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1694700623
transform 1 0 1232 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1694700623
transform 1 0 1232 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1694700623
transform 1 0 1232 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1694700623
transform -1 0 1120 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1694700623
transform 1 0 1568 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_8 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1120 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_12 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1344 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_28 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2240 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32
timestamp 1694700623
transform 1 0 2464 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1694700623
transform 1 0 4592 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1694700623
transform 1 0 4816 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104
timestamp 1694700623
transform 1 0 6496 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1694700623
transform 1 0 6720 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_142 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 8624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_150
timestamp 1694700623
transform 1 0 9072 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1694700623
transform 1 0 1120 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_12
timestamp 1694700623
transform 1 0 1344 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_44
timestamp 1694700623
transform 1 0 3136 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_60
timestamp 1694700623
transform 1 0 4032 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1694700623
transform 1 0 4480 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1694700623
transform 1 0 4704 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_148
timestamp 1694700623
transform 1 0 8960 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1694700623
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1694700623
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1694700623
transform 1 0 6664 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_123
timestamp 1694700623
transform 1 0 7560 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1694700623
transform 1 0 1120 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_12
timestamp 1694700623
transform 1 0 1344 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_44
timestamp 1694700623
transform 1 0 3136 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_60
timestamp 1694700623
transform 1 0 4032 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1694700623
transform 1 0 4480 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1694700623
transform 1 0 4704 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_104
timestamp 1694700623
transform 1 0 6496 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_112
timestamp 1694700623
transform 1 0 6944 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1694700623
transform 1 0 9072 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1694700623
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1694700623
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1694700623
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1694700623
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1694700623
transform 1 0 6664 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_123
timestamp 1694700623
transform 1 0 7560 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1694700623
transform 1 0 1120 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1694700623
transform 1 0 1344 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1694700623
transform 1 0 3136 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_60
timestamp 1694700623
transform 1 0 4032 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1694700623
transform 1 0 4480 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_72
timestamp 1694700623
transform 1 0 4704 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_104
timestamp 1694700623
transform 1 0 6496 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_112
timestamp 1694700623
transform 1 0 6944 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1694700623
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1694700623
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1694700623
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1694700623
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_107
timestamp 1694700623
transform 1 0 6664 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_111
timestamp 1694700623
transform 1 0 6888 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_113
timestamp 1694700623
transform 1 0 7000 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1694700623
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1694700623
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1694700623
transform 1 0 4704 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_104
timestamp 1694700623
transform 1 0 6496 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1694700623
transform 1 0 1120 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1694700623
transform 1 0 1344 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1694700623
transform 1 0 2240 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1694700623
transform 1 0 2464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1694700623
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1694700623
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1694700623
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1694700623
transform 1 0 6664 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_115
timestamp 1694700623
transform 1 0 7112 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_117
timestamp 1694700623
transform 1 0 7224 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1694700623
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1694700623
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_72
timestamp 1694700623
transform 1 0 4704 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_104
timestamp 1694700623
transform 1 0 6496 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_112
timestamp 1694700623
transform 1 0 6944 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_148
timestamp 1694700623
transform 1 0 8960 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1694700623
transform 1 0 1120 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1694700623
transform 1 0 1344 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1694700623
transform 1 0 2240 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1694700623
transform 1 0 2464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1694700623
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1694700623
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1694700623
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_107
timestamp 1694700623
transform 1 0 6664 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_123
timestamp 1694700623
transform 1 0 7560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_125
timestamp 1694700623
transform 1 0 7672 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1694700623
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1694700623
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1694700623
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1694700623
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1694700623
transform 1 0 8848 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1694700623
transform 1 0 9072 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1694700623
transform 1 0 1120 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1694700623
transform 1 0 1344 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1694700623
transform 1 0 2240 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1694700623
transform 1 0 2464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1694700623
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1694700623
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1694700623
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1694700623
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1694700623
transform 1 0 7560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_125
timestamp 1694700623
transform 1 0 7672 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1694700623
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1694700623
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1694700623
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_104
timestamp 1694700623
transform 1 0 6496 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_112
timestamp 1694700623
transform 1 0 6944 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_8
timestamp 1694700623
transform 1 0 1120 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_12
timestamp 1694700623
transform 1 0 1344 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_28
timestamp 1694700623
transform 1 0 2240 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1694700623
transform 1 0 2464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1694700623
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1694700623
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1694700623
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1694700623
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1694700623
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1694700623
transform 1 0 7336 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1694700623
transform 1 0 7448 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1694700623
transform 1 0 784 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_8
timestamp 1694700623
transform 1 0 1120 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_40
timestamp 1694700623
transform 1 0 2912 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_56
timestamp 1694700623
transform 1 0 3808 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_64
timestamp 1694700623
transform 1 0 4256 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1694700623
transform 1 0 4480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1694700623
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_14
timestamp 1694700623
transform 1 0 1456 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_18
timestamp 1694700623
transform 1 0 1680 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_36
timestamp 1694700623
transform 1 0 2688 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_70
timestamp 1694700623
transform 1 0 4592 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_74
timestamp 1694700623
transform 1 0 4816 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_104
timestamp 1694700623
transform 1 0 6496 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_108
timestamp 1694700623
transform 1 0 6720 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_150
timestamp 1694700623
transform 1 0 9072 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1694700623
transform 1 0 784 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1694700623
transform 1 0 784 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1694700623
transform 1 0 784 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1694700623
transform 1 0 784 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1694700623
transform 1 0 784 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1694700623
transform 1 0 784 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1694700623
transform 1 0 784 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1694700623
transform 1 0 784 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1694700623
transform 1 0 1120 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1694700623
transform 1 0 784 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 7056 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1694700623
transform -1 0 9184 0 1 3920
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1694700623
transform 1 0 7056 0 -1 4704
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1694700623
transform -1 0 9184 0 1 3136
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1694700623
transform -1 0 8512 0 -1 3920
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1694700623
transform -1 0 9184 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1694700623
transform -1 0 8512 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1694700623
transform -1 0 8288 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1694700623
transform 1 0 7056 0 -1 3136
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1694700623
transform -1 0 6384 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1694700623
transform -1 0 8288 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1694700623
transform 1 0 7056 0 -1 5488
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1694700623
transform -1 0 9184 0 1 4704
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1694700623
transform 1 0 7728 0 1 5488
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1694700623
transform -1 0 9184 0 1 6272
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1694700623
transform -1 0 9184 0 1 7056
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1694700623
transform -1 0 8512 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1694700623
transform -1 0 8512 0 -1 7056
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1694700623
transform -1 0 7056 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1694700623
transform -1 0 6384 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 9296 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1694700623
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1694700623
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 9296 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1694700623
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 9296 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1694700623
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 9296 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1694700623
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 9296 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1694700623
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 9296 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1694700623
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 9296 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1694700623
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 9296 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1694700623
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 9296 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1694700623
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 9296 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1694700623
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 9296 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1694700623
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1694700623
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1694700623
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 9296 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1694700623
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1694700623
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 9296 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1694700623
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1694700623
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1694700623
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_38
timestamp 1694700623
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1694700623
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_40
timestamp 1694700623
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1694700623
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_42
timestamp 1694700623
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_43
timestamp 1694700623
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_44
timestamp 1694700623
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_45
timestamp 1694700623
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_46
timestamp 1694700623
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_47
timestamp 1694700623
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_48
timestamp 1694700623
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_49
timestamp 1694700623
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_50
timestamp 1694700623
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_51
timestamp 1694700623
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_52
timestamp 1694700623
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_53
timestamp 1694700623
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_54
timestamp 1694700623
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_55
timestamp 1694700623
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_56
timestamp 1694700623
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_57
timestamp 1694700623
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_58
timestamp 1694700623
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_59
timestamp 1694700623
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_60
timestamp 1694700623
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_61
timestamp 1694700623
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_62
timestamp 1694700623
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_63
timestamp 1694700623
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_64
timestamp 1694700623
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_65
timestamp 1694700623
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_66
timestamp 1694700623
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_67
timestamp 1694700623
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_68
timestamp 1694700623
transform 1 0 2576 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_69
timestamp 1694700623
transform 1 0 4480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_70
timestamp 1694700623
transform 1 0 6384 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_71
timestamp 1694700623
transform 1 0 8288 0 1 7840
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 896 400 952 0 FreeSans 224 0 0 0 input_signal[0]
port 0 nsew signal input
flabel metal3 s 0 1792 400 1848 0 FreeSans 224 0 0 0 input_signal[1]
port 1 nsew signal input
flabel metal3 s 0 2688 400 2744 0 FreeSans 224 0 0 0 input_signal[2]
port 2 nsew signal input
flabel metal3 s 0 3584 400 3640 0 FreeSans 224 0 0 0 input_signal[3]
port 3 nsew signal input
flabel metal3 s 0 4480 400 4536 0 FreeSans 224 0 0 0 input_signal[4]
port 4 nsew signal input
flabel metal3 s 0 5376 400 5432 0 FreeSans 224 0 0 0 input_signal[5]
port 5 nsew signal input
flabel metal3 s 0 6272 400 6328 0 FreeSans 224 0 0 0 input_signal[6]
port 6 nsew signal input
flabel metal3 s 0 7168 400 7224 0 FreeSans 224 0 0 0 input_signal[7]
port 7 nsew signal input
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 input_signal[8]
port 8 nsew signal input
flabel metal3 s 0 8960 400 9016 0 FreeSans 224 0 0 0 input_signal[9]
port 9 nsew signal input
flabel metal3 s 9600 672 10000 728 0 FreeSans 224 0 0 0 output_signal_minus[0]
port 10 nsew signal tristate
flabel metal3 s 9600 4704 10000 4760 0 FreeSans 224 0 0 0 output_signal_minus[1]
port 11 nsew signal tristate
flabel metal3 s 9600 4256 10000 4312 0 FreeSans 224 0 0 0 output_signal_minus[2]
port 12 nsew signal tristate
flabel metal3 s 9600 3808 10000 3864 0 FreeSans 224 0 0 0 output_signal_minus[3]
port 13 nsew signal tristate
flabel metal3 s 9600 3360 10000 3416 0 FreeSans 224 0 0 0 output_signal_minus[4]
port 14 nsew signal tristate
flabel metal3 s 9600 2912 10000 2968 0 FreeSans 224 0 0 0 output_signal_minus[5]
port 15 nsew signal tristate
flabel metal3 s 9600 2464 10000 2520 0 FreeSans 224 0 0 0 output_signal_minus[6]
port 16 nsew signal tristate
flabel metal3 s 9600 2016 10000 2072 0 FreeSans 224 0 0 0 output_signal_minus[7]
port 17 nsew signal tristate
flabel metal3 s 9600 1568 10000 1624 0 FreeSans 224 0 0 0 output_signal_minus[8]
port 18 nsew signal tristate
flabel metal3 s 9600 1120 10000 1176 0 FreeSans 224 0 0 0 output_signal_minus[9]
port 19 nsew signal tristate
flabel metal3 s 9600 9184 10000 9240 0 FreeSans 224 0 0 0 output_signal_plus[0]
port 20 nsew signal tristate
flabel metal3 s 9600 5152 10000 5208 0 FreeSans 224 0 0 0 output_signal_plus[1]
port 21 nsew signal tristate
flabel metal3 s 9600 5600 10000 5656 0 FreeSans 224 0 0 0 output_signal_plus[2]
port 22 nsew signal tristate
flabel metal3 s 9600 6048 10000 6104 0 FreeSans 224 0 0 0 output_signal_plus[3]
port 23 nsew signal tristate
flabel metal3 s 9600 6496 10000 6552 0 FreeSans 224 0 0 0 output_signal_plus[4]
port 24 nsew signal tristate
flabel metal3 s 9600 6944 10000 7000 0 FreeSans 224 0 0 0 output_signal_plus[5]
port 25 nsew signal tristate
flabel metal3 s 9600 7392 10000 7448 0 FreeSans 224 0 0 0 output_signal_plus[6]
port 26 nsew signal tristate
flabel metal3 s 9600 7840 10000 7896 0 FreeSans 224 0 0 0 output_signal_plus[7]
port 27 nsew signal tristate
flabel metal3 s 9600 8288 10000 8344 0 FreeSans 224 0 0 0 output_signal_plus[8]
port 28 nsew signal tristate
flabel metal3 s 9600 8736 10000 8792 0 FreeSans 224 0 0 0 output_signal_plus[9]
port 29 nsew signal tristate
flabel metal4 s 1670 1538 1830 8262 0 FreeSans 640 90 0 0 vdd
port 30 nsew power bidirectional
flabel metal4 s 3826 1538 3986 8262 0 FreeSans 640 90 0 0 vdd
port 30 nsew power bidirectional
flabel metal4 s 5982 1538 6142 8262 0 FreeSans 640 90 0 0 vdd
port 30 nsew power bidirectional
flabel metal4 s 8138 1538 8298 8262 0 FreeSans 640 90 0 0 vdd
port 30 nsew power bidirectional
flabel metal4 s 2748 1538 2908 8262 0 FreeSans 640 90 0 0 vss
port 31 nsew ground bidirectional
flabel metal4 s 4904 1538 5064 8262 0 FreeSans 640 90 0 0 vss
port 31 nsew ground bidirectional
flabel metal4 s 7060 1538 7220 8262 0 FreeSans 640 90 0 0 vss
port 31 nsew ground bidirectional
flabel metal4 s 9216 1538 9376 8262 0 FreeSans 640 90 0 0 vss
port 31 nsew ground bidirectional
rlabel metal1 4984 8232 4984 8232 0 vdd
rlabel via1 5024 7840 5024 7840 0 vss
rlabel metal2 868 1316 868 1316 0 input_signal[0]
rlabel metal2 868 1988 868 1988 0 input_signal[1]
rlabel metal2 868 2828 868 2828 0 input_signal[2]
rlabel metal2 868 3668 868 3668 0 input_signal[3]
rlabel metal2 868 4676 868 4676 0 input_signal[4]
rlabel metal2 868 5516 868 5516 0 input_signal[5]
rlabel metal2 868 6356 868 6356 0 input_signal[6]
rlabel metal3 623 7196 623 7196 0 input_signal[7]
rlabel metal2 1204 8064 1204 8064 0 input_signal[8]
rlabel metal2 868 8512 868 8512 0 input_signal[9]
rlabel metal2 1036 1764 1036 1764 0 net1
rlabel metal3 2618 7924 2618 7924 0 net10
rlabel metal2 8484 2016 8484 2016 0 net11
rlabel metal2 9044 3976 9044 3976 0 net12
rlabel metal2 7252 4368 7252 4368 0 net13
rlabel metal2 8988 3192 8988 3192 0 net14
rlabel metal3 8540 3052 8540 3052 0 net15
rlabel metal2 9016 3500 9016 3500 0 net16
rlabel metal2 8148 2156 8148 2156 0 net17
rlabel metal2 8204 1820 8204 1820 0 net18
rlabel metal2 7364 3570 7364 3570 0 net19
rlabel metal2 1064 2268 1064 2268 0 net2
rlabel metal3 7728 1764 7728 1764 0 net20
rlabel metal3 8344 2268 8344 2268 0 net21
rlabel metal2 7476 5068 7476 5068 0 net22
rlabel metal2 8708 4018 8708 4018 0 net23
rlabel metal2 7672 4060 7672 4060 0 net24
rlabel metal2 8708 4900 8708 4900 0 net25
rlabel metal2 8904 5404 8904 5404 0 net26
rlabel metal2 8680 6972 8680 6972 0 net27
rlabel metal2 8372 7280 8372 7280 0 net28
rlabel metal2 6972 7784 6972 7784 0 net29
rlabel metal2 1036 3276 1036 3276 0 net3
rlabel metal2 8820 8008 8820 8008 0 net30
rlabel metal2 7084 4004 7084 4004 0 net4
rlabel metal2 8764 3248 8764 3248 0 net5
rlabel metal2 1036 5656 1036 5656 0 net6
rlabel metal2 8764 6272 8764 6272 0 net7
rlabel metal2 1036 7224 1036 7224 0 net8
rlabel metal2 1372 7840 1372 7840 0 net9
rlabel metal2 6468 1456 6468 1456 0 output_signal_minus[0]
rlabel metal2 8596 4424 8596 4424 0 output_signal_minus[1]
rlabel metal2 8344 4396 8344 4396 0 output_signal_minus[2]
rlabel metal3 9121 3836 9121 3836 0 output_signal_minus[3]
rlabel metal2 7924 3500 7924 3500 0 output_signal_minus[4]
rlabel metal3 9009 2940 9009 2940 0 output_signal_minus[5]
rlabel metal2 7924 2380 7924 2380 0 output_signal_minus[6]
rlabel metal3 8589 2044 8589 2044 0 output_signal_minus[7]
rlabel metal2 7644 2688 7644 2688 0 output_signal_minus[8]
rlabel metal3 7721 1148 7721 1148 0 output_signal_minus[9]
rlabel metal3 8561 9212 8561 9212 0 output_signal_plus[0]
rlabel metal3 8981 5180 8981 5180 0 output_signal_plus[1]
rlabel metal3 9121 5628 9121 5628 0 output_signal_plus[2]
rlabel metal2 8988 5936 8988 5936 0 output_signal_plus[3]
rlabel metal3 9121 6524 9121 6524 0 output_signal_plus[4]
rlabel metal3 9121 6972 9121 6972 0 output_signal_plus[5]
rlabel metal3 7924 7560 7924 7560 0 output_signal_plus[6]
rlabel metal2 7812 7336 7812 7336 0 output_signal_plus[7]
rlabel metal2 6468 8036 6468 8036 0 output_signal_plus[8]
rlabel metal3 7721 8764 7721 8764 0 output_signal_plus[9]
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
