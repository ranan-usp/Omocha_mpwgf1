* NGSPICE file created from dac_in.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1 VDD VSS VPW VNW a_1380_472# a_36_472#
+ a_932_472# a_572_375# a_124_375# a_1468_375# a_1020_375# a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_1020_375# VNW 0.181468f
C1 a_932_472# a_484_472# 0.013276f
C2 a_36_472# a_484_472# 0.013276f
C3 a_124_375# VNW 0.180172f
C4 VSS VNW 0.017643f
C5 VSS a_1020_375# 0.134699f
C6 a_1468_375# VNW 0.18122f
C7 a_1020_375# a_1468_375# 0.012552f
C8 a_572_375# VNW 0.181468f
C9 VSS a_124_375# 0.134699f
C10 a_1380_472# VNW 0.024396f
C11 VNW VDD 0.217349f
C12 a_572_375# a_1020_375# 0.012552f
C13 a_1380_472# a_1020_375# 0.086905f
C14 a_1020_375# VDD 0.129962f
C15 VSS a_1468_375# 0.082091f
C16 a_484_472# VNW 0.024018f
C17 a_124_375# a_572_375# 0.012552f
C18 VSS a_572_375# 0.134699f
C19 a_124_375# VDD 0.12673f
C20 VSS a_1380_472# 0.144845f
C21 VSS VDD 0.026369f
C22 a_932_472# VNW 0.024018f
C23 a_932_472# a_1020_375# 0.285629f
C24 a_1380_472# a_1468_375# 0.285629f
C25 a_1468_375# VDD 0.129266f
C26 a_124_375# a_484_472# 0.086905f
C27 a_36_472# VNW 0.025611f
C28 VSS a_484_472# 0.148077f
C29 a_572_375# VDD 0.129962f
C30 a_1380_472# VDD 0.179463f
C31 VSS a_932_472# 0.148077f
C32 a_572_375# a_484_472# 0.285629f
C33 a_36_472# a_124_375# 0.285629f
C34 VSS a_36_472# 0.147381f
C35 a_484_472# VDD 0.179463f
C36 a_932_472# a_572_375# 0.086905f
C37 a_932_472# a_1380_472# 0.013276f
C38 a_932_472# VDD 0.179463f
C39 a_36_472# VDD 0.093681f
C40 VSS VSUBS 0.642184f
C41 VDD VSUBS 0.493288f
C42 VNW VSUBS 3.05206f
C43 a_1380_472# VSUBS 0.345058f
C44 a_932_472# VSUBS 0.33241f
C45 a_484_472# VSUBS 0.33241f
C46 a_36_472# VSUBS 0.404746f
C47 a_1468_375# VSUBS 0.233029f
C48 a_1020_375# VSUBS 0.171606f
C49 a_572_375# VSUBS 0.171606f
C50 a_124_375# VSUBS 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8$1 Z I VDD VSS VPW VNW a_224_472# VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 Z I 0.001907f
C1 VDD I 0.1311f
C2 I a_224_472# 0.796069f
C3 Z VSS 0.70427f
C4 Z VNW 0.038011f
C5 VDD VSS 0.031131f
C6 VDD VNW 0.305516f
C7 VSS a_224_472# 0.659695f
C8 a_224_472# VNW 1.14633f
C9 VSS I 0.158668f
C10 I VNW 0.55539f
C11 VSS VNW 0.01282f
C12 VDD Z 0.819024f
C13 Z a_224_472# 2.29481f
C14 VDD a_224_472# 0.74621f
C15 VSS VSUBS 0.910368f
C16 Z VSUBS 0.18914f
C17 VDD VSUBS 0.724491f
C18 I VSUBS 1.16773f
C19 VNW VSUBS 4.79254f
C20 a_224_472# VSUBS 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS VPW VNW a_1916_375# a_4516_472#
+ a_1380_472# a_3260_375# a_5860_472# a_36_472# a_932_472# a_2812_375# a_5412_472#
+ a_2276_472# a_4156_375# a_6756_472# a_1828_472# a_3708_375# a_3172_472# a_572_375#
+ a_6308_472# a_5052_375# a_2724_472# a_6396_375# a_4604_375# a_124_375# a_1468_375#
+ a_4068_472# a_5948_375# a_3620_472# a_1020_375# a_5500_375# a_4964_472# a_484_472#
+ a_2364_375# a_6844_375# VSUBS
X0 a_4604_375# a_4516_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3 a_4156_375# a_4068_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 a_5500_375# a_5412_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 VDD a_5052_375# a_4964_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 VDD a_6844_375# a_6756_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 a_5052_375# a_4964_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X11 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_4604_375# a_4516_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X14 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X15 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X16 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X17 a_5948_375# a_5860_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X18 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X19 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X20 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X21 VDD a_5500_375# a_5412_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X22 a_6844_375# a_6756_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X23 a_6396_375# a_6308_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X24 VDD a_6396_375# a_6308_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X25 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X26 VDD a_4156_375# a_4068_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X27 VDD a_5948_375# a_5860_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X28 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X29 a_3708_375# a_3620_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X30 VDD a_3708_375# a_3620_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X31 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_2276_472# VSS 0.144729f
C1 VDD a_572_375# 0.129962f
C2 a_3620_472# VSS 0.144729f
C3 VSS a_6308_472# 0.144729f
C4 a_4964_472# VDD 0.179463f
C5 a_5860_472# VSS 0.144729f
C6 VNW a_124_375# 0.180172f
C7 a_4068_472# a_3620_472# 0.013276f
C8 a_1916_375# VNW 0.181468f
C9 a_1828_472# VSS 0.144729f
C10 a_3620_472# a_3172_472# 0.013276f
C11 VSS a_484_472# 0.144729f
C12 a_3620_472# a_3260_375# 0.087066f
C13 a_4516_472# a_4964_472# 0.013276f
C14 a_2276_472# VNW 0.024018f
C15 a_3620_472# VNW 0.024018f
C16 a_572_375# VSS 0.132921f
C17 a_1468_375# a_1020_375# 0.012882f
C18 a_6756_472# a_6844_375# 0.285629f
C19 VNW a_6308_472# 0.024018f
C20 VNW a_5860_472# 0.024018f
C21 a_4964_472# VSS 0.144729f
C22 VDD a_1020_375# 0.129962f
C23 a_4964_472# a_4604_375# 0.087066f
C24 a_2812_375# a_2724_472# 0.285629f
C25 a_1380_472# a_1468_375# 0.285629f
C26 a_1828_472# VNW 0.024018f
C27 a_1380_472# VDD 0.179463f
C28 a_5412_472# a_5052_375# 0.087066f
C29 a_2276_472# a_1916_375# 0.087066f
C30 VNW a_484_472# 0.024018f
C31 VDD a_3708_375# 0.129962f
C32 VNW a_572_375# 0.181468f
C33 a_2812_375# VDD 0.129962f
C34 a_4964_472# VNW 0.024018f
C35 a_932_472# VDD 0.179463f
C36 VSS a_1020_375# 0.132921f
C37 VDD a_5052_375# 0.129962f
C38 a_1828_472# a_1916_375# 0.285629f
C39 a_124_375# a_484_472# 0.087066f
C40 a_2812_375# a_2364_375# 0.012882f
C41 a_5500_375# a_5052_375# 0.012882f
C42 a_6756_472# VDD 0.179463f
C43 a_1380_472# VSS 0.144729f
C44 a_124_375# a_572_375# 0.012882f
C45 a_5860_472# a_6308_472# 0.013276f
C46 a_6756_472# a_6396_375# 0.087066f
C47 a_1828_472# a_2276_472# 0.013276f
C48 a_3708_375# VSS 0.132921f
C49 VDD a_6844_375# 0.129266f
C50 a_6396_375# a_6844_375# 0.012882f
C51 a_4068_472# a_3708_375# 0.087066f
C52 a_2812_375# VSS 0.132921f
C53 VNW a_1020_375# 0.181468f
C54 a_932_472# VSS 0.144729f
C55 VSS a_5052_375# 0.132921f
C56 a_4604_375# a_5052_375# 0.012882f
C57 a_3708_375# a_4156_375# 0.012882f
C58 a_2812_375# a_3172_472# 0.087066f
C59 a_1380_472# VNW 0.024018f
C60 a_3260_375# a_3708_375# 0.012882f
C61 a_6756_472# VSS 0.141496f
C62 VDD a_2724_472# 0.179463f
C63 VDD a_5412_472# 0.179463f
C64 VNW a_3708_375# 0.181468f
C65 a_2812_375# a_3260_375# 0.012882f
C66 VSS a_6844_375# 0.081619f
C67 a_5500_375# a_5412_472# 0.285629f
C68 a_2812_375# VNW 0.181468f
C69 a_2724_472# a_2364_375# 0.087066f
C70 a_5948_375# VDD 0.129962f
C71 a_572_375# a_484_472# 0.285629f
C72 a_932_472# VNW 0.024018f
C73 a_5948_375# a_6396_375# 0.012882f
C74 VNW a_5052_375# 0.181468f
C75 VDD a_1468_375# 0.129962f
C76 a_5500_375# a_5948_375# 0.012882f
C77 VDD a_36_472# 0.093681f
C78 VDD a_6396_375# 0.129962f
C79 a_6756_472# VNW 0.024396f
C80 VSS a_2724_472# 0.144729f
C81 a_5500_375# VDD 0.129962f
C82 a_5412_472# VSS 0.144729f
C83 VDD a_2364_375# 0.129962f
C84 VNW a_6844_375# 0.18122f
C85 a_3620_472# a_3708_375# 0.285629f
C86 a_4516_472# VDD 0.179463f
C87 a_5948_375# VSS 0.132921f
C88 a_3172_472# a_2724_472# 0.013276f
C89 a_1468_375# VSS 0.132921f
C90 a_1828_472# a_1380_472# 0.013276f
C91 VSS a_36_472# 0.144033f
C92 VDD VSS 0.105475f
C93 VDD a_4604_375# 0.129962f
C94 a_6396_375# VSS 0.132921f
C95 a_572_375# a_1020_375# 0.012882f
C96 VNW a_2724_472# 0.024018f
C97 VNW a_5412_472# 0.024018f
C98 a_5500_375# VSS 0.132921f
C99 a_4068_472# VDD 0.179463f
C100 VSS a_2364_375# 0.132921f
C101 VDD a_3172_472# 0.179463f
C102 a_6756_472# a_6308_472# 0.013276f
C103 a_5948_375# VNW 0.181468f
C104 a_4516_472# VSS 0.144729f
C105 a_4516_472# a_4604_375# 0.285629f
C106 VDD a_4156_375# 0.129962f
C107 VDD a_3260_375# 0.129962f
C108 VNW a_1468_375# 0.181468f
C109 a_932_472# a_484_472# 0.013276f
C110 VNW a_36_472# 0.025611f
C111 VNW VDD 0.842606f
C112 a_4068_472# a_4516_472# 0.013276f
C113 VSS a_4604_375# 0.132921f
C114 VNW a_6396_375# 0.181468f
C115 a_932_472# a_572_375# 0.087066f
C116 a_5500_375# VNW 0.181468f
C117 a_4068_472# VSS 0.144729f
C118 VNW a_2364_375# 0.181468f
C119 a_4964_472# a_5052_375# 0.285629f
C120 a_4516_472# a_4156_375# 0.087066f
C121 a_2276_472# a_2724_472# 0.013276f
C122 VSS a_3172_472# 0.144729f
C123 a_124_375# a_36_472# 0.285629f
C124 VDD a_124_375# 0.12673f
C125 a_1916_375# a_1468_375# 0.012882f
C126 a_4516_472# VNW 0.024018f
C127 a_1380_472# a_1020_375# 0.087066f
C128 VSS a_4156_375# 0.132921f
C129 a_4156_375# a_4604_375# 0.012882f
C130 a_1916_375# VDD 0.129962f
C131 a_5412_472# a_5860_472# 0.013276f
C132 a_3260_375# VSS 0.132921f
C133 VNW VSS 0.070573f
C134 VNW a_4604_375# 0.181468f
C135 a_4068_472# a_4156_375# 0.285629f
C136 a_5948_375# a_6308_472# 0.087066f
C137 a_1916_375# a_2364_375# 0.012882f
C138 a_5948_375# a_5860_472# 0.285629f
C139 a_2276_472# VDD 0.179463f
C140 a_4068_472# VNW 0.024018f
C141 a_932_472# a_1020_375# 0.285629f
C142 a_3260_375# a_3172_472# 0.285629f
C143 a_3620_472# VDD 0.179463f
C144 VDD a_6308_472# 0.179463f
C145 VNW a_3172_472# 0.024018f
C146 VDD a_5860_472# 0.179463f
C147 a_6396_375# a_6308_472# 0.285629f
C148 a_2276_472# a_2364_375# 0.285629f
C149 a_932_472# a_1380_472# 0.013276f
C150 a_124_375# VSS 0.132921f
C151 a_1828_472# a_1468_375# 0.087066f
C152 VNW a_4156_375# 0.181468f
C153 a_4964_472# a_5412_472# 0.013276f
C154 VNW a_3260_375# 0.181468f
C155 a_1828_472# VDD 0.179463f
C156 a_1916_375# VSS 0.132921f
C157 a_5500_375# a_5860_472# 0.087066f
C158 a_36_472# a_484_472# 0.013276f
C159 VDD a_484_472# 0.179463f
C160 VSS VSUBS 2.33708f
C161 VDD VSUBS 1.73533f
C162 VNW VSUBS 11.406401f
C163 a_6756_472# VSUBS 0.345058f
C164 a_6308_472# VSUBS 0.33241f
C165 a_5860_472# VSUBS 0.33241f
C166 a_5412_472# VSUBS 0.33241f
C167 a_4964_472# VSUBS 0.33241f
C168 a_4516_472# VSUBS 0.33241f
C169 a_4068_472# VSUBS 0.33241f
C170 a_3620_472# VSUBS 0.33241f
C171 a_3172_472# VSUBS 0.33241f
C172 a_2724_472# VSUBS 0.33241f
C173 a_2276_472# VSUBS 0.33241f
C174 a_1828_472# VSUBS 0.33241f
C175 a_1380_472# VSUBS 0.33241f
C176 a_932_472# VSUBS 0.33241f
C177 a_484_472# VSUBS 0.33241f
C178 a_36_472# VSUBS 0.404746f
C179 a_6844_375# VSUBS 0.233068f
C180 a_6396_375# VSUBS 0.171644f
C181 a_5948_375# VSUBS 0.171644f
C182 a_5500_375# VSUBS 0.171644f
C183 a_5052_375# VSUBS 0.171644f
C184 a_4604_375# VSUBS 0.171644f
C185 a_4156_375# VSUBS 0.171644f
C186 a_3708_375# VSUBS 0.171644f
C187 a_3260_375# VSUBS 0.171644f
C188 a_2812_375# VSUBS 0.171644f
C189 a_2364_375# VSUBS 0.171644f
C190 a_1916_375# VSUBS 0.171644f
C191 a_1468_375# VSUBS 0.171644f
C192 a_1020_375# VSUBS 0.171644f
C193 a_572_375# VSUBS 0.171644f
C194 a_124_375# VSUBS 0.185708f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1 VDD VSS VPW VNW a_1916_375# a_1380_472#
+ a_3260_375# a_36_472# a_932_472# a_2812_375# a_2276_472# a_1828_472# a_3172_472#
+ a_572_375# a_2724_472# a_124_375# a_1468_375# a_1020_375# a_484_472# a_2364_375#
+ VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_124_375# a_484_472# 0.087174f
C1 a_2364_375# a_2724_472# 0.087174f
C2 a_2364_375# a_1916_375# 0.013103f
C3 a_3172_472# VNW 0.024396f
C4 a_1828_472# a_2276_472# 0.013276f
C5 a_2276_472# VNW 0.024018f
C6 a_124_375# a_36_472# 0.285629f
C7 a_1828_472# VSS 0.142721f
C8 VSS VNW 0.035286f
C9 a_2812_375# VDD 0.129962f
C10 a_1020_375# VNW 0.181468f
C11 a_36_472# a_484_472# 0.013276f
C12 a_3172_472# a_2724_472# 0.013276f
C13 VDD a_3260_375# 0.129266f
C14 a_2276_472# a_2724_472# 0.013276f
C15 VSS a_2724_472# 0.142721f
C16 a_1828_472# a_1380_472# 0.013276f
C17 VNW a_1380_472# 0.024018f
C18 a_2276_472# a_1916_375# 0.087174f
C19 VSS a_1916_375# 0.131736f
C20 a_124_375# VNW 0.180172f
C21 a_572_375# a_932_472# 0.087174f
C22 VNW a_484_472# 0.024018f
C23 a_2364_375# VDD 0.129962f
C24 a_572_375# VDD 0.129962f
C25 VSS a_1468_375# 0.131736f
C26 a_1020_375# a_1468_375# 0.013103f
C27 a_2812_375# a_3260_375# 0.013103f
C28 VNW a_36_472# 0.025611f
C29 VSS a_932_472# 0.142721f
C30 a_3172_472# VDD 0.179463f
C31 a_1468_375# a_1380_472# 0.285629f
C32 a_1020_375# a_932_472# 0.285629f
C33 a_2276_472# VDD 0.179463f
C34 VSS VDD 0.052737f
C35 a_1020_375# VDD 0.129962f
C36 a_2812_375# a_2364_375# 0.013103f
C37 a_932_472# a_1380_472# 0.013276f
C38 VDD a_1380_472# 0.179463f
C39 a_1828_472# VNW 0.024018f
C40 a_124_375# VDD 0.12673f
C41 a_484_472# a_932_472# 0.013276f
C42 a_3172_472# a_2812_375# 0.087174f
C43 VDD a_484_472# 0.179463f
C44 a_2812_375# VSS 0.131736f
C45 VNW a_2724_472# 0.024018f
C46 a_3172_472# a_3260_375# 0.285629f
C47 a_1828_472# a_1916_375# 0.285629f
C48 VNW a_1916_375# 0.181468f
C49 VSS a_3260_375# 0.081304f
C50 VDD a_36_472# 0.093681f
C51 a_1828_472# a_1468_375# 0.087174f
C52 VNW a_1468_375# 0.181468f
C53 a_2276_472# a_2364_375# 0.285629f
C54 VSS a_2364_375# 0.131736f
C55 a_572_375# VSS 0.131736f
C56 a_572_375# a_1020_375# 0.013103f
C57 VNW a_932_472# 0.024018f
C58 a_1468_375# a_1916_375# 0.013103f
C59 a_1828_472# VDD 0.179463f
C60 VNW VDD 0.425768f
C61 a_3172_472# VSS 0.139489f
C62 a_2276_472# VSS 0.142721f
C63 a_1020_375# VSS 0.131736f
C64 a_124_375# a_572_375# 0.013103f
C65 VDD a_2724_472# 0.179463f
C66 a_572_375# a_484_472# 0.285629f
C67 VDD a_1916_375# 0.129962f
C68 VSS a_1380_472# 0.142721f
C69 a_1020_375# a_1380_472# 0.087174f
C70 a_2812_375# VNW 0.181468f
C71 a_124_375# VSS 0.131736f
C72 VDD a_1468_375# 0.129962f
C73 VNW a_3260_375# 0.18122f
C74 VSS a_484_472# 0.142721f
C75 a_2812_375# a_2724_472# 0.285629f
C76 VDD a_932_472# 0.179463f
C77 VSS a_36_472# 0.142026f
C78 VNW a_2364_375# 0.181468f
C79 a_572_375# VNW 0.181468f
C80 VSS VSUBS 1.20585f
C81 VDD VSUBS 0.907304f
C82 VNW VSUBS 5.83682f
C83 a_3172_472# VSUBS 0.345058f
C84 a_2724_472# VSUBS 0.33241f
C85 a_2276_472# VSUBS 0.33241f
C86 a_1828_472# VSUBS 0.33241f
C87 a_1380_472# VSUBS 0.33241f
C88 a_932_472# VSUBS 0.33241f
C89 a_484_472# VSUBS 0.33241f
C90 a_36_472# VSUBS 0.404746f
C91 a_3260_375# VSUBS 0.233093f
C92 a_2812_375# VSUBS 0.17167f
C93 a_2364_375# VSUBS 0.17167f
C94 a_1916_375# VSUBS 0.17167f
C95 a_1468_375# VSUBS 0.17167f
C96 a_1020_375# VSUBS 0.17167f
C97 a_572_375# VSUBS 0.17167f
C98 a_124_375# VSUBS 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna$1 VSS I VDD VPW VNW VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 VSS VDD 0.009725f
C1 VDD VNW 0.048519f
C2 VDD I 0.017439f
C3 VSS VNW 0.007461f
C4 VSS I 0.031625f
C5 VNW I 0.027206f
C6 VSS VSUBS 0.12617f
C7 VDD VSUBS 0.087026f
C8 I VSUBS 0.139667f
C9 VNW VSUBS 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1 VDD VSS VPW VNW a_36_472# a_124_375#
+ VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VDD VNW 0.061035f
C1 VNW a_124_375# 0.179924f
C2 VSS VNW 0.004411f
C3 VNW a_36_472# 0.025989f
C4 VDD a_124_375# 0.126034f
C5 VDD VSS 0.006592f
C6 VSS a_124_375# 0.082879f
C7 VDD a_36_472# 0.093681f
C8 a_124_375# a_36_472# 0.285629f
C9 VSS a_36_472# 0.150876f
C10 VSS VSUBS 0.218985f
C11 VDD VSUBS 0.182777f
C12 VNW VSUBS 0.96348f
C13 a_36_472# VSUBS 0.417394f
C14 a_124_375# VSUBS 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1 VDD VSS VPW VNW a_36_472# a_572_375#
+ a_124_375# a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 a_484_472# a_36_472# 0.013276f
C1 VSS VDD 0.013184f
C2 a_36_472# a_124_375# 0.285629f
C3 VDD a_572_375# 0.129266f
C4 VNW a_36_472# 0.025611f
C5 VSS a_36_472# 0.151218f
C6 a_484_472# a_124_375# 0.086742f
C7 a_484_472# VNW 0.024396f
C8 VNW a_124_375# 0.180172f
C9 a_36_472# VDD 0.093681f
C10 VSS a_484_472# 0.148682f
C11 a_484_472# a_572_375# 0.285629f
C12 VSS a_124_375# 0.136476f
C13 VSS VNW 0.008822f
C14 a_124_375# a_572_375# 0.012222f
C15 VNW a_572_375# 0.18122f
C16 a_484_472# VDD 0.179463f
C17 VDD a_124_375# 0.12673f
C18 VSS a_572_375# 0.082563f
C19 VNW VDD 0.11314f
C20 VSS VSUBS 0.360066f
C21 VDD VSUBS 0.286281f
C22 VNW VSUBS 1.65967f
C23 a_484_472# VSUBS 0.345058f
C24 a_36_472# VSUBS 0.404746f
C25 a_572_375# VSUBS 0.232991f
C26 a_124_375# VSUBS 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1$1 VSS ZN I VDD VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD VNW 0.076257f
C1 VSS VNW 0.011339f
C2 VDD ZN 0.137375f
C3 I VDD 0.041847f
C4 VSS ZN 0.115297f
C5 I VSS 0.0533f
C6 VDD VSS 0.025626f
C7 ZN VNW 0.022202f
C8 I VNW 0.137757f
C9 I ZN 0.262199f
C10 VSS VSUBS 0.2316f
C11 ZN VSUBS 0.113404f
C12 VDD VSUBS 0.181139f
C13 I VSUBS 0.341982f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD VNW 0.076212f
C1 VSS VNW 0.011085f
C2 VDD ZN 0.098026f
C3 I VDD 0.157124f
C4 VSS ZN 0.077008f
C5 I VSS 0.058937f
C6 VDD VSS 0.025441f
C7 ZN VNW 0.031181f
C8 I VNW 0.135368f
C9 I ZN 0.47009f
C10 VSS VSUBS 0.242183f
C11 ZN VSUBS 0.095505f
C12 VDD VSUBS 0.182097f
C13 I VSUBS 0.355642f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1 VSS Z I VDD VPW VNW a_36_113# VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 I a_36_113# 0.476912f
C1 Z a_36_113# 0.191876f
C2 VSS a_36_113# 0.11114f
C3 I VDD 0.028968f
C4 VNW I 0.152645f
C5 Z VDD 0.085355f
C6 VNW Z 0.030118f
C7 VSS VDD 0.009561f
C8 VNW VSS 0.009307f
C9 I Z 0.031362f
C10 I VSS 0.070302f
C11 Z VSS 0.136942f
C12 VDD a_36_113# 0.278283f
C13 VNW a_36_113# 0.160792f
C14 VNW VDD 0.088196f
C15 VSS VSUBS 0.283681f
C16 Z VSUBS 0.117185f
C17 VDD VSUBS 0.180237f
C18 I VSUBS 0.336876f
C19 VNW VSUBS 1.31158f
C20 a_36_113# VSUBS 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1$1 VSS Z I VDD VPW VNW a_36_160# VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 I VSS 0.12329f
C1 I a_36_160# 0.545454f
C2 I VDD 0.02612f
C3 I VNW 0.2276f
C4 Z VSS 0.146199f
C5 a_36_160# Z 0.281838f
C6 VDD Z 0.128274f
C7 VNW Z 0.030347f
C8 a_36_160# VSS 0.074156f
C9 VDD VSS 0.009574f
C10 VNW VSS 0.009324f
C11 a_36_160# VDD 0.2736f
C12 I Z 0.041707f
C13 a_36_160# VNW 0.170864f
C14 VNW VDD 0.087464f
C15 VSS VSUBS 0.28275f
C16 Z VSUBS 0.10469f
C17 VDD VSUBS 0.178615f
C18 I VSUBS 0.323491f
C19 VNW VSUBS 1.31158f
C20 a_36_160# VSUBS 0.386641f
.ends

.subckt phase_inverter input_signal[0] input_signal[1] input_signal[2] input_signal[3]
+ input_signal[4] input_signal[5] input_signal[9] output_signal_minus[1] output_signal_minus[2]
+ output_signal_minus[3] output_signal_minus[4] output_signal_minus[5] output_signal_minus[6]
+ output_signal_minus[7] output_signal_minus[8] output_signal_minus[9] output_signal_plus[1]
+ output_signal_plus[2] output_signal_plus[3] output_signal_plus[4] output_signal_plus[5]
+ output_signal_plus[6] output_signal_plus[7] _10_/Z input_signal[7] _19_/Z FILLER_0_0_12/a_484_472#
+ FILLER_0_0_36/a_2276_472# _08_/ZN FILLER_0_16_36/a_2364_375# input_signal[8] output18/a_224_472#
+ _19_/I _00_/ZN output_signal_plus[0] _10_/I output_signal_plus[9] FILLER_0_16_36/a_124_375#
+ output20/a_224_472# output30/a_224_472# input_signal[6] FILLER_0_0_36/a_36_472#
+ output21/a_224_472# FILLER_0_16_18/a_124_375# output_signal_minus[0] output_signal_plus[8]
+ vdd vss
XFILLER_0_1_72 vdd vss FILLER_0_1_72/VPW vdd FILLER_0_1_72/a_1380_472# FILLER_0_1_72/a_36_472#
+ FILLER_0_1_72/a_932_472# FILLER_0_1_72/a_572_375# FILLER_0_1_72/a_124_375# FILLER_0_1_72/a_1468_375#
+ FILLER_0_1_72/a_1020_375# FILLER_0_1_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput20 output_signal_minus[9] _00_/ZN vdd vss output20/VPW vdd output20/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput21 output_signal_plus[0] _10_/Z vdd vss output21/VPW vdd output21/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_9_2 vdd vss FILLER_0_9_2/VPW vdd FILLER_0_9_2/a_1916_375# FILLER_0_9_2/a_4516_472#
+ FILLER_0_9_2/a_1380_472# FILLER_0_9_2/a_3260_375# FILLER_0_9_2/a_5860_472# FILLER_0_9_2/a_36_472#
+ FILLER_0_9_2/a_932_472# FILLER_0_9_2/a_2812_375# FILLER_0_9_2/a_5412_472# FILLER_0_9_2/a_2276_472#
+ FILLER_0_9_2/a_4156_375# FILLER_0_9_2/a_6756_472# FILLER_0_9_2/a_1828_472# FILLER_0_9_2/a_3708_375#
+ FILLER_0_9_2/a_3172_472# FILLER_0_9_2/a_572_375# FILLER_0_9_2/a_6308_472# FILLER_0_9_2/a_5052_375#
+ FILLER_0_9_2/a_2724_472# FILLER_0_9_2/a_6396_375# FILLER_0_9_2/a_4604_375# FILLER_0_9_2/a_124_375#
+ FILLER_0_9_2/a_1468_375# FILLER_0_9_2/a_4068_472# FILLER_0_9_2/a_5948_375# FILLER_0_9_2/a_3620_472#
+ FILLER_0_9_2/a_1020_375# FILLER_0_9_2/a_5500_375# FILLER_0_9_2/a_4964_472# FILLER_0_9_2/a_484_472#
+ FILLER_0_9_2/a_2364_375# FILLER_0_9_2/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_72 vdd vss FILLER_0_7_72/VPW vdd FILLER_0_7_72/a_1916_375# FILLER_0_7_72/a_1380_472#
+ FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472# FILLER_0_7_72/a_932_472# FILLER_0_7_72/a_2812_375#
+ FILLER_0_7_72/a_2276_472# FILLER_0_7_72/a_1828_472# FILLER_0_7_72/a_3172_472# FILLER_0_7_72/a_572_375#
+ FILLER_0_7_72/a_2724_472# FILLER_0_7_72/a_124_375# FILLER_0_7_72/a_1468_375# FILLER_0_7_72/a_1020_375#
+ FILLER_0_7_72/a_484_472# FILLER_0_7_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XANTENNA_input3_I vss input_signal[2] vdd ANTENNA_input3_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
Xoutput22 output_signal_plus[1] _11_/Z vdd vss output22/VPW vdd output22/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput11 output_signal_minus[0] _01_/ZN vdd vss output11/VPW vdd output11/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_12_101 vdd vss FILLER_0_12_101/VPW vdd FILLER_0_12_101/a_36_472# FILLER_0_12_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xoutput23 output_signal_plus[2] _12_/Z vdd vss output23/VPW vdd output23/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput12 output_signal_minus[1] _02_/ZN vdd vss output12/VPW vdd output12/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_13_66 vdd vss FILLER_0_13_66/VPW vdd FILLER_0_13_66/a_36_472# FILLER_0_13_66/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_10_12 vdd vss FILLER_0_10_12/VPW vdd FILLER_0_10_12/a_1380_472# FILLER_0_10_12/a_36_472#
+ FILLER_0_10_12/a_932_472# FILLER_0_10_12/a_572_375# FILLER_0_10_12/a_124_375# FILLER_0_10_12/a_1468_375#
+ FILLER_0_10_12/a_1020_375# FILLER_0_10_12/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput24 output_signal_plus[3] _13_/Z vdd vss output24/VPW vdd output24/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_8_107 vdd vss FILLER_0_8_107/VPW vdd FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_572_375#
+ FILLER_0_8_107/a_124_375# FILLER_0_8_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
Xoutput13 output_signal_minus[2] _03_/ZN vdd vss output13/VPW vdd output13/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_7_2 vdd vss FILLER_0_7_2/VPW vdd FILLER_0_7_2/a_1916_375# FILLER_0_7_2/a_4516_472#
+ FILLER_0_7_2/a_1380_472# FILLER_0_7_2/a_3260_375# FILLER_0_7_2/a_5860_472# FILLER_0_7_2/a_36_472#
+ FILLER_0_7_2/a_932_472# FILLER_0_7_2/a_2812_375# FILLER_0_7_2/a_5412_472# FILLER_0_7_2/a_2276_472#
+ FILLER_0_7_2/a_4156_375# FILLER_0_7_2/a_6756_472# FILLER_0_7_2/a_1828_472# FILLER_0_7_2/a_3708_375#
+ FILLER_0_7_2/a_3172_472# FILLER_0_7_2/a_572_375# FILLER_0_7_2/a_6308_472# FILLER_0_7_2/a_5052_375#
+ FILLER_0_7_2/a_2724_472# FILLER_0_7_2/a_6396_375# FILLER_0_7_2/a_4604_375# FILLER_0_7_2/a_124_375#
+ FILLER_0_7_2/a_1468_375# FILLER_0_7_2/a_4068_472# FILLER_0_7_2/a_5948_375# FILLER_0_7_2/a_3620_472#
+ FILLER_0_7_2/a_1020_375# FILLER_0_7_2/a_5500_375# FILLER_0_7_2/a_4964_472# FILLER_0_7_2/a_484_472#
+ FILLER_0_7_2/a_2364_375# FILLER_0_7_2/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I vss input_signal[0] vdd ANTENNA_input1_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_1_44 vdd vss FILLER_0_1_44/VPW vdd FILLER_0_1_44/a_1380_472# FILLER_0_1_44/a_36_472#
+ FILLER_0_1_44/a_932_472# FILLER_0_1_44/a_572_375# FILLER_0_1_44/a_124_375# FILLER_0_1_44/a_1468_375#
+ FILLER_0_1_44/a_1020_375# FILLER_0_1_44/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput25 output_signal_plus[4] _14_/Z vdd vss output25/VPW vdd output25/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput14 output_signal_minus[3] _04_/ZN vdd vss output14/VPW vdd output14/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_1_12 vdd vss FILLER_0_1_12/VPW vdd FILLER_0_1_12/a_1916_375# FILLER_0_1_12/a_1380_472#
+ FILLER_0_1_12/a_3260_375# FILLER_0_1_12/a_36_472# FILLER_0_1_12/a_932_472# FILLER_0_1_12/a_2812_375#
+ FILLER_0_1_12/a_2276_472# FILLER_0_1_12/a_1828_472# FILLER_0_1_12/a_3172_472# FILLER_0_1_12/a_572_375#
+ FILLER_0_1_12/a_2724_472# FILLER_0_1_12/a_124_375# FILLER_0_1_12/a_1468_375# FILLER_0_1_12/a_1020_375#
+ FILLER_0_1_12/a_484_472# FILLER_0_1_12/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xoutput26 output_signal_plus[5] _15_/Z vdd vss output26/VPW vdd output26/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_09_ vss _09_/ZN _18_/I vdd _09_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xoutput15 output_signal_minus[4] net15 vdd vss output15/VPW vdd output15/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_4_101 vdd vss FILLER_0_4_101/VPW vdd FILLER_0_4_101/a_36_472# FILLER_0_4_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_7_66 vdd vss FILLER_0_7_66/VPW vdd FILLER_0_7_66/a_36_472# FILLER_0_7_66/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_10_37 vdd vss FILLER_0_10_37/VPW vdd FILLER_0_10_37/a_1916_375# FILLER_0_10_37/a_4516_472#
+ FILLER_0_10_37/a_1380_472# FILLER_0_10_37/a_3260_375# FILLER_0_10_37/a_5860_472#
+ FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_932_472# FILLER_0_10_37/a_2812_375# FILLER_0_10_37/a_5412_472#
+ FILLER_0_10_37/a_2276_472# FILLER_0_10_37/a_4156_375# FILLER_0_10_37/a_6756_472#
+ FILLER_0_10_37/a_1828_472# FILLER_0_10_37/a_3708_375# FILLER_0_10_37/a_3172_472#
+ FILLER_0_10_37/a_572_375# FILLER_0_10_37/a_6308_472# FILLER_0_10_37/a_5052_375#
+ FILLER_0_10_37/a_2724_472# FILLER_0_10_37/a_6396_375# FILLER_0_10_37/a_4604_375#
+ FILLER_0_10_37/a_124_375# FILLER_0_10_37/a_1468_375# FILLER_0_10_37/a_4068_472#
+ FILLER_0_10_37/a_5948_375# FILLER_0_10_37/a_3620_472# FILLER_0_10_37/a_1020_375#
+ FILLER_0_10_37/a_5500_375# FILLER_0_10_37/a_4964_472# FILLER_0_10_37/a_484_472#
+ FILLER_0_10_37/a_2364_375# FILLER_0_10_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_36 vdd vss FILLER_0_16_36/VPW vdd FILLER_0_16_36/a_1916_375# FILLER_0_16_36/a_1380_472#
+ FILLER_0_16_36/a_3260_375# FILLER_0_16_36/a_36_472# FILLER_0_16_36/a_932_472# FILLER_0_16_36/a_2812_375#
+ FILLER_0_16_36/a_2276_472# FILLER_0_16_36/a_1828_472# FILLER_0_16_36/a_3172_472#
+ FILLER_0_16_36/a_572_375# FILLER_0_16_36/a_2724_472# FILLER_0_16_36/a_124_375# FILLER_0_16_36/a_1468_375#
+ FILLER_0_16_36/a_1020_375# FILLER_0_16_36/a_484_472# FILLER_0_16_36/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_08_ vss _08_/ZN _17_/I vdd _08_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xoutput27 output_signal_plus[6] _16_/Z vdd vss output27/VPW vdd output27/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput16 output_signal_minus[5] _06_/ZN vdd vss output16/VPW vdd output16/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput28 output_signal_plus[7] _17_/Z vdd vss output28/VPW vdd output28/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_07_ vss _07_/ZN _16_/I vdd _07_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xoutput17 output_signal_minus[6] _07_/ZN vdd vss output17/VPW vdd output17/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_10_28 vdd vss FILLER_0_10_28/VPW vdd FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_12_107 vdd vss FILLER_0_12_107/VPW vdd FILLER_0_12_107/a_1380_472# FILLER_0_12_107/a_36_472#
+ FILLER_0_12_107/a_932_472# FILLER_0_12_107/a_572_375# FILLER_0_12_107/a_124_375#
+ FILLER_0_12_107/a_1468_375# FILLER_0_12_107/a_1020_375# FILLER_0_12_107/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput29 output_signal_plus[8] _18_/Z vdd vss output29/VPW vdd output29/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_06_ vdd vss _15_/I _06_/ZN _06_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
Xoutput18 output_signal_minus[7] _08_/ZN vdd vss output18/VPW vdd output18/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_4_37 vdd vss FILLER_0_4_37/VPW vdd FILLER_0_4_37/a_1916_375# FILLER_0_4_37/a_4516_472#
+ FILLER_0_4_37/a_1380_472# FILLER_0_4_37/a_3260_375# FILLER_0_4_37/a_5860_472# FILLER_0_4_37/a_36_472#
+ FILLER_0_4_37/a_932_472# FILLER_0_4_37/a_2812_375# FILLER_0_4_37/a_5412_472# FILLER_0_4_37/a_2276_472#
+ FILLER_0_4_37/a_4156_375# FILLER_0_4_37/a_6756_472# FILLER_0_4_37/a_1828_472# FILLER_0_4_37/a_3708_375#
+ FILLER_0_4_37/a_3172_472# FILLER_0_4_37/a_572_375# FILLER_0_4_37/a_6308_472# FILLER_0_4_37/a_5052_375#
+ FILLER_0_4_37/a_2724_472# FILLER_0_4_37/a_6396_375# FILLER_0_4_37/a_4604_375# FILLER_0_4_37/a_124_375#
+ FILLER_0_4_37/a_1468_375# FILLER_0_4_37/a_4068_472# FILLER_0_4_37/a_5948_375# FILLER_0_4_37/a_3620_472#
+ FILLER_0_4_37/a_1020_375# FILLER_0_4_37/a_5500_375# FILLER_0_4_37/a_4964_472# FILLER_0_4_37/a_484_472#
+ FILLER_0_4_37/a_2364_375# FILLER_0_4_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_72 vdd vss FILLER_0_11_72/VPW vdd FILLER_0_11_72/a_1916_375# FILLER_0_11_72/a_4516_472#
+ FILLER_0_11_72/a_1380_472# FILLER_0_11_72/a_3260_375# FILLER_0_11_72/a_5860_472#
+ FILLER_0_11_72/a_36_472# FILLER_0_11_72/a_932_472# FILLER_0_11_72/a_2812_375# FILLER_0_11_72/a_5412_472#
+ FILLER_0_11_72/a_2276_472# FILLER_0_11_72/a_4156_375# FILLER_0_11_72/a_6756_472#
+ FILLER_0_11_72/a_1828_472# FILLER_0_11_72/a_3708_375# FILLER_0_11_72/a_3172_472#
+ FILLER_0_11_72/a_572_375# FILLER_0_11_72/a_6308_472# FILLER_0_11_72/a_5052_375#
+ FILLER_0_11_72/a_2724_472# FILLER_0_11_72/a_6396_375# FILLER_0_11_72/a_4604_375#
+ FILLER_0_11_72/a_124_375# FILLER_0_11_72/a_1468_375# FILLER_0_11_72/a_4068_472#
+ FILLER_0_11_72/a_5948_375# FILLER_0_11_72/a_3620_472# FILLER_0_11_72/a_1020_375#
+ FILLER_0_11_72/a_5500_375# FILLER_0_11_72/a_4964_472# FILLER_0_11_72/a_484_472#
+ FILLER_0_11_72/a_2364_375# FILLER_0_11_72/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__04__I vss _13_/I vdd ANTENNA__04__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
Xoutput19 output_signal_minus[8] _09_/ZN vdd vss output19/VPW vdd output19/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_05_ vdd vss _14_/I net15 _05_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
XFILLER_0_16_18 vdd vss FILLER_0_16_18/VPW vdd FILLER_0_16_18/a_1380_472# FILLER_0_16_18/a_36_472#
+ FILLER_0_16_18/a_932_472# FILLER_0_16_18/a_572_375# FILLER_0_16_18/a_124_375# FILLER_0_16_18/a_1468_375#
+ FILLER_0_16_18/a_1020_375# FILLER_0_16_18/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XANTENNA_input8_I vss input_signal[7] vdd ANTENNA_input8_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XANTENNA__15__I vss _15_/I vdd ANTENNA__15__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
X_04_ vdd vss _13_/I _04_/ZN _04_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
XFILLER_0_0_142 vdd vss FILLER_0_0_142/VPW vdd FILLER_0_0_142/a_36_472# FILLER_0_0_142/a_572_375#
+ FILLER_0_0_142/a_124_375# FILLER_0_0_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_5_60 vdd vss FILLER_0_5_60/VPW vdd FILLER_0_5_60/a_36_472# FILLER_0_5_60/a_572_375#
+ FILLER_0_5_60/a_124_375# FILLER_0_5_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_7_104 vdd vss FILLER_0_7_104/VPW vdd FILLER_0_7_104/a_36_472# FILLER_0_7_104/a_572_375#
+ FILLER_0_7_104/a_124_375# FILLER_0_7_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_03_ vdd vss _12_/I _03_/ZN _03_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
Xinput1 vss _10_/I input_signal[0] vdd input1/VPW vdd input1/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_4_107 vdd vss FILLER_0_4_107/VPW vdd FILLER_0_4_107/a_1380_472# FILLER_0_4_107/a_36_472#
+ FILLER_0_4_107/a_932_472# FILLER_0_4_107/a_572_375# FILLER_0_4_107/a_124_375# FILLER_0_4_107/a_1468_375#
+ FILLER_0_4_107/a_1020_375# FILLER_0_4_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_5_72 vdd vss FILLER_0_5_72/VPW vdd FILLER_0_5_72/a_1916_375# FILLER_0_5_72/a_1380_472#
+ FILLER_0_5_72/a_3260_375# FILLER_0_5_72/a_36_472# FILLER_0_5_72/a_932_472# FILLER_0_5_72/a_2812_375#
+ FILLER_0_5_72/a_2276_472# FILLER_0_5_72/a_1828_472# FILLER_0_5_72/a_3172_472# FILLER_0_5_72/a_572_375#
+ FILLER_0_5_72/a_2724_472# FILLER_0_5_72/a_124_375# FILLER_0_5_72/a_1468_375# FILLER_0_5_72/a_1020_375#
+ FILLER_0_5_72/a_484_472# FILLER_0_5_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xinput2 vss _11_/I input_signal[1] vdd input2/VPW vdd input2/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
X_02_ vdd vss _11_/I _02_/ZN _02_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
X_01_ vdd vss _10_/I _01_/ZN _01_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
Xinput3 vss _12_/I input_signal[2] vdd input3/VPW vdd input3/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA_input6_I vss input_signal[5] vdd ANTENNA_input6_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_11_66 vdd vss FILLER_0_11_66/VPW vdd FILLER_0_11_66/a_36_472# FILLER_0_11_66/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xinput4 vss _13_/I input_signal[3] vdd input4/VPW vdd input4/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
X_00_ vss _00_/ZN _19_/I vdd _00_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xinput5 vss _14_/I input_signal[4] vdd input5/VPW vdd input5/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_11_136 vdd vss FILLER_0_11_136/VPW vdd FILLER_0_11_136/a_36_472# FILLER_0_11_136/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_14_12 vdd vss FILLER_0_14_12/VPW vdd FILLER_0_14_12/a_1380_472# FILLER_0_14_12/a_36_472#
+ FILLER_0_14_12/a_932_472# FILLER_0_14_12/a_572_375# FILLER_0_14_12/a_124_375# FILLER_0_14_12/a_1468_375#
+ FILLER_0_14_12/a_1020_375# FILLER_0_14_12/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_14_101 vdd vss FILLER_0_14_101/VPW vdd FILLER_0_14_101/a_36_472# FILLER_0_14_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xinput6 vss _15_/I input_signal[5] vdd input6/VPW vdd input6/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_0_104 vdd vss FILLER_0_0_104/VPW vdd FILLER_0_0_104/a_36_472# FILLER_0_0_104/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA_input4_I vss input_signal[3] vdd ANTENNA_input4_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
Xinput7 vss _16_/I input_signal[6] vdd input7/VPW vdd input7/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_5_44 vdd vss FILLER_0_5_44/VPW vdd FILLER_0_5_44/a_1380_472# FILLER_0_5_44/a_36_472#
+ FILLER_0_5_44/a_932_472# FILLER_0_5_44/a_572_375# FILLER_0_5_44/a_124_375# FILLER_0_5_44/a_1468_375#
+ FILLER_0_5_44/a_1020_375# FILLER_0_5_44/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xinput10 vss _19_/I input_signal[9] vdd input10/VPW vdd input10/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_5_12 vdd vss FILLER_0_5_12/VPW vdd FILLER_0_5_12/a_1916_375# FILLER_0_5_12/a_1380_472#
+ FILLER_0_5_12/a_3260_375# FILLER_0_5_12/a_36_472# FILLER_0_5_12/a_932_472# FILLER_0_5_12/a_2812_375#
+ FILLER_0_5_12/a_2276_472# FILLER_0_5_12/a_1828_472# FILLER_0_5_12/a_3172_472# FILLER_0_5_12/a_572_375#
+ FILLER_0_5_12/a_2724_472# FILLER_0_5_12/a_124_375# FILLER_0_5_12/a_1468_375# FILLER_0_5_12/a_1020_375#
+ FILLER_0_5_12/a_484_472# FILLER_0_5_12/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xinput8 vss _17_/I input_signal[7] vdd input8/VPW vdd input8/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_14_37 vdd vss FILLER_0_14_37/VPW vdd FILLER_0_14_37/a_1916_375# FILLER_0_14_37/a_4516_472#
+ FILLER_0_14_37/a_1380_472# FILLER_0_14_37/a_3260_375# FILLER_0_14_37/a_5860_472#
+ FILLER_0_14_37/a_36_472# FILLER_0_14_37/a_932_472# FILLER_0_14_37/a_2812_375# FILLER_0_14_37/a_5412_472#
+ FILLER_0_14_37/a_2276_472# FILLER_0_14_37/a_4156_375# FILLER_0_14_37/a_6756_472#
+ FILLER_0_14_37/a_1828_472# FILLER_0_14_37/a_3708_375# FILLER_0_14_37/a_3172_472#
+ FILLER_0_14_37/a_572_375# FILLER_0_14_37/a_6308_472# FILLER_0_14_37/a_5052_375#
+ FILLER_0_14_37/a_2724_472# FILLER_0_14_37/a_6396_375# FILLER_0_14_37/a_4604_375#
+ FILLER_0_14_37/a_124_375# FILLER_0_14_37/a_1468_375# FILLER_0_14_37/a_4068_472#
+ FILLER_0_14_37/a_5948_375# FILLER_0_14_37/a_3620_472# FILLER_0_14_37/a_1020_375#
+ FILLER_0_14_37/a_5500_375# FILLER_0_14_37/a_4964_472# FILLER_0_14_37/a_484_472#
+ FILLER_0_14_37/a_2364_375# FILLER_0_14_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_12 vdd vss FILLER_0_8_12/VPW vdd FILLER_0_8_12/a_1380_472# FILLER_0_8_12/a_36_472#
+ FILLER_0_8_12/a_932_472# FILLER_0_8_12/a_572_375# FILLER_0_8_12/a_124_375# FILLER_0_8_12/a_1468_375#
+ FILLER_0_8_12/a_1020_375# FILLER_0_8_12/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xinput9 vss _18_/I input_signal[8] vdd input9/VPW vdd input9/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_14_115 vdd vss FILLER_0_14_115/VPW vdd FILLER_0_14_115/a_36_472# FILLER_0_14_115/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_6_101 vdd vss FILLER_0_6_101/VPW vdd FILLER_0_6_101/a_36_472# FILLER_0_6_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_3_104 vdd vss FILLER_0_3_104/VPW vdd FILLER_0_3_104/a_36_472# FILLER_0_3_104/a_572_375#
+ FILLER_0_3_104/a_124_375# FILLER_0_3_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XANTENNA_input10_I vss input_signal[9] vdd ANTENNA_input10_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XANTENNA_input2_I vss input_signal[1] vdd ANTENNA_input2_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_2_37 vdd vss FILLER_0_2_37/VPW vdd FILLER_0_2_37/a_1916_375# FILLER_0_2_37/a_4516_472#
+ FILLER_0_2_37/a_1380_472# FILLER_0_2_37/a_3260_375# FILLER_0_2_37/a_5860_472# FILLER_0_2_37/a_36_472#
+ FILLER_0_2_37/a_932_472# FILLER_0_2_37/a_2812_375# FILLER_0_2_37/a_5412_472# FILLER_0_2_37/a_2276_472#
+ FILLER_0_2_37/a_4156_375# FILLER_0_2_37/a_6756_472# FILLER_0_2_37/a_1828_472# FILLER_0_2_37/a_3708_375#
+ FILLER_0_2_37/a_3172_472# FILLER_0_2_37/a_572_375# FILLER_0_2_37/a_6308_472# FILLER_0_2_37/a_5052_375#
+ FILLER_0_2_37/a_2724_472# FILLER_0_2_37/a_6396_375# FILLER_0_2_37/a_4604_375# FILLER_0_2_37/a_124_375#
+ FILLER_0_2_37/a_1468_375# FILLER_0_2_37/a_4068_472# FILLER_0_2_37/a_5948_375# FILLER_0_2_37/a_3620_472#
+ FILLER_0_2_37/a_1020_375# FILLER_0_2_37/a_5500_375# FILLER_0_2_37/a_4964_472# FILLER_0_2_37/a_484_472#
+ FILLER_0_2_37/a_2364_375# FILLER_0_2_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_28 vdd vss FILLER_0_14_28/VPW vdd FILLER_0_14_28/a_36_472# FILLER_0_14_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_0_70 vdd vss FILLER_0_0_70/VPW vdd FILLER_0_0_70/a_36_472# FILLER_0_0_70/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA__02__I vss _11_/I vdd ANTENNA__02__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
X_19_ vss _19_/Z _19_/I vdd _19_/VPW vdd _19_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_8_37 vdd vss FILLER_0_8_37/VPW vdd FILLER_0_8_37/a_1916_375# FILLER_0_8_37/a_4516_472#
+ FILLER_0_8_37/a_1380_472# FILLER_0_8_37/a_3260_375# FILLER_0_8_37/a_5860_472# FILLER_0_8_37/a_36_472#
+ FILLER_0_8_37/a_932_472# FILLER_0_8_37/a_2812_375# FILLER_0_8_37/a_5412_472# FILLER_0_8_37/a_2276_472#
+ FILLER_0_8_37/a_4156_375# FILLER_0_8_37/a_6756_472# FILLER_0_8_37/a_1828_472# FILLER_0_8_37/a_3708_375#
+ FILLER_0_8_37/a_3172_472# FILLER_0_8_37/a_572_375# FILLER_0_8_37/a_6308_472# FILLER_0_8_37/a_5052_375#
+ FILLER_0_8_37/a_2724_472# FILLER_0_8_37/a_6396_375# FILLER_0_8_37/a_4604_375# FILLER_0_8_37/a_124_375#
+ FILLER_0_8_37/a_1468_375# FILLER_0_8_37/a_4068_472# FILLER_0_8_37/a_5948_375# FILLER_0_8_37/a_3620_472#
+ FILLER_0_8_37/a_1020_375# FILLER_0_8_37/a_5500_375# FILLER_0_8_37/a_4964_472# FILLER_0_8_37/a_484_472#
+ FILLER_0_8_37/a_2364_375# FILLER_0_8_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05__I vss _14_/I vdd ANTENNA__05__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_15_72 vdd vss FILLER_0_15_72/VPW vdd FILLER_0_15_72/a_1380_472# FILLER_0_15_72/a_36_472#
+ FILLER_0_15_72/a_932_472# FILLER_0_15_72/a_572_375# FILLER_0_15_72/a_124_375# FILLER_0_15_72/a_1468_375#
+ FILLER_0_15_72/a_1020_375# FILLER_0_15_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XANTENNA__13__I vss _13_/I vdd ANTENNA__13__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_14_107 vdd vss FILLER_0_14_107/VPW vdd FILLER_0_14_107/a_36_472# FILLER_0_14_107/a_572_375#
+ FILLER_0_14_107/a_124_375# FILLER_0_14_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_3_60 vdd vss FILLER_0_3_60/VPW vdd FILLER_0_3_60/a_36_472# FILLER_0_3_60/a_572_375#
+ FILLER_0_3_60/a_124_375# FILLER_0_3_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_18_ vss _18_/Z _18_/I vdd _18_/VPW vdd _18_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_40 vdd vss FILLER_0_15_40/VPW vdd FILLER_0_15_40/a_1380_472# FILLER_0_15_40/a_36_472#
+ FILLER_0_15_40/a_932_472# FILLER_0_15_40/a_572_375# FILLER_0_15_40/a_124_375# FILLER_0_15_40/a_1468_375#
+ FILLER_0_15_40/a_1020_375# FILLER_0_15_40/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_6_2 vdd vss FILLER_0_6_2/VPW vdd FILLER_0_6_2/a_1916_375# FILLER_0_6_2/a_1380_472#
+ FILLER_0_6_2/a_3260_375# FILLER_0_6_2/a_36_472# FILLER_0_6_2/a_932_472# FILLER_0_6_2/a_2812_375#
+ FILLER_0_6_2/a_2276_472# FILLER_0_6_2/a_1828_472# FILLER_0_6_2/a_3172_472# FILLER_0_6_2/a_572_375#
+ FILLER_0_6_2/a_2724_472# FILLER_0_6_2/a_124_375# FILLER_0_6_2/a_1468_375# FILLER_0_6_2/a_1020_375#
+ FILLER_0_6_2/a_484_472# FILLER_0_6_2/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_17_ vss _17_/Z _17_/I vdd _17_/VPW vdd _17_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_8_28 vdd vss FILLER_0_8_28/VPW vdd FILLER_0_8_28/a_36_472# FILLER_0_8_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_3_72 vdd vss FILLER_0_3_72/VPW vdd FILLER_0_3_72/a_1916_375# FILLER_0_3_72/a_1380_472#
+ FILLER_0_3_72/a_3260_375# FILLER_0_3_72/a_36_472# FILLER_0_3_72/a_932_472# FILLER_0_3_72/a_2812_375#
+ FILLER_0_3_72/a_2276_472# FILLER_0_3_72/a_1828_472# FILLER_0_3_72/a_3172_472# FILLER_0_3_72/a_572_375#
+ FILLER_0_3_72/a_2724_472# FILLER_0_3_72/a_124_375# FILLER_0_3_72/a_1468_375# FILLER_0_3_72/a_1020_375#
+ FILLER_0_3_72/a_484_472# FILLER_0_3_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_10_101 vdd vss FILLER_0_10_101/VPW vdd FILLER_0_10_101/a_36_472# FILLER_0_10_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_16_ vss _16_/Z _16_/I vdd _16_/VPW vdd _16_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_64 vdd vss FILLER_0_15_64/VPW vdd FILLER_0_15_64/a_36_472# FILLER_0_15_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_9_72 vdd vss FILLER_0_9_72/VPW vdd FILLER_0_9_72/a_1916_375# FILLER_0_9_72/a_1380_472#
+ FILLER_0_9_72/a_3260_375# FILLER_0_9_72/a_36_472# FILLER_0_9_72/a_932_472# FILLER_0_9_72/a_2812_375#
+ FILLER_0_9_72/a_2276_472# FILLER_0_9_72/a_1828_472# FILLER_0_9_72/a_3172_472# FILLER_0_9_72/a_572_375#
+ FILLER_0_9_72/a_2724_472# FILLER_0_9_72/a_124_375# FILLER_0_9_72/a_1468_375# FILLER_0_9_72/a_1020_375#
+ FILLER_0_9_72/a_484_472# FILLER_0_9_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_9_104 vdd vss FILLER_0_9_104/VPW vdd FILLER_0_9_104/a_36_472# FILLER_0_9_104/a_572_375#
+ FILLER_0_9_104/a_124_375# FILLER_0_9_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_6_107 vdd vss FILLER_0_6_107/VPW vdd FILLER_0_6_107/a_36_472# FILLER_0_6_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_15_ vss _15_/Z _15_/I vdd _15_/VPW vdd _15_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_2 vdd vss FILLER_0_15_2/VPW vdd FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_4_2 vdd vss FILLER_0_4_2/VPW vdd FILLER_0_4_2/a_1916_375# FILLER_0_4_2/a_1380_472#
+ FILLER_0_4_2/a_3260_375# FILLER_0_4_2/a_36_472# FILLER_0_4_2/a_932_472# FILLER_0_4_2/a_2812_375#
+ FILLER_0_4_2/a_2276_472# FILLER_0_4_2/a_1828_472# FILLER_0_4_2/a_3172_472# FILLER_0_4_2/a_572_375#
+ FILLER_0_4_2/a_2724_472# FILLER_0_4_2/a_124_375# FILLER_0_4_2/a_1468_375# FILLER_0_4_2/a_1020_375#
+ FILLER_0_4_2/a_484_472# FILLER_0_4_2/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_14_ vss _14_/Z _14_/I vdd _14_/VPW vdd _14_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA_input9_I vss input_signal[8] vdd ANTENNA_input9_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_12_12 vdd vss FILLER_0_12_12/VPW vdd FILLER_0_12_12/a_1380_472# FILLER_0_12_12/a_36_472#
+ FILLER_0_12_12/a_932_472# FILLER_0_12_12/a_572_375# FILLER_0_12_12/a_124_375# FILLER_0_12_12/a_1468_375#
+ FILLER_0_12_12/a_1020_375# FILLER_0_12_12/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_2_101 vdd vss FILLER_0_2_101/VPW vdd FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_13_ vss _13_/Z _13_/I vdd _13_/VPW vdd _13_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_56 vdd vss FILLER_0_15_56/VPW vdd FILLER_0_15_56/a_36_472# FILLER_0_15_56/a_572_375#
+ FILLER_0_15_56/a_124_375# FILLER_0_15_56/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_12_ vss _12_/Z _12_/I vdd _12_/VPW vdd _12_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_3_44 vdd vss FILLER_0_3_44/VPW vdd FILLER_0_3_44/a_1380_472# FILLER_0_3_44/a_36_472#
+ FILLER_0_3_44/a_932_472# FILLER_0_3_44/a_572_375# FILLER_0_3_44/a_124_375# FILLER_0_3_44/a_1468_375#
+ FILLER_0_3_44/a_1020_375# FILLER_0_3_44/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_0_12 vdd vss FILLER_0_0_12/VPW vdd FILLER_0_0_12/a_1380_472# FILLER_0_0_12/a_36_472#
+ FILLER_0_0_12/a_932_472# FILLER_0_0_12/a_572_375# FILLER_0_0_12/a_124_375# FILLER_0_0_12/a_1468_375#
+ FILLER_0_0_12/a_1020_375# FILLER_0_0_12/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_13_2 vdd vss FILLER_0_13_2/VPW vdd FILLER_0_13_2/a_1916_375# FILLER_0_13_2/a_4516_472#
+ FILLER_0_13_2/a_1380_472# FILLER_0_13_2/a_3260_375# FILLER_0_13_2/a_5860_472# FILLER_0_13_2/a_36_472#
+ FILLER_0_13_2/a_932_472# FILLER_0_13_2/a_2812_375# FILLER_0_13_2/a_5412_472# FILLER_0_13_2/a_2276_472#
+ FILLER_0_13_2/a_4156_375# FILLER_0_13_2/a_6756_472# FILLER_0_13_2/a_1828_472# FILLER_0_13_2/a_3708_375#
+ FILLER_0_13_2/a_3172_472# FILLER_0_13_2/a_572_375# FILLER_0_13_2/a_6308_472# FILLER_0_13_2/a_5052_375#
+ FILLER_0_13_2/a_2724_472# FILLER_0_13_2/a_6396_375# FILLER_0_13_2/a_4604_375# FILLER_0_13_2/a_124_375#
+ FILLER_0_13_2/a_1468_375# FILLER_0_13_2/a_4068_472# FILLER_0_13_2/a_5948_375# FILLER_0_13_2/a_3620_472#
+ FILLER_0_13_2/a_1020_375# FILLER_0_13_2/a_5500_375# FILLER_0_13_2/a_4964_472# FILLER_0_13_2/a_484_472#
+ FILLER_0_13_2/a_2364_375# FILLER_0_13_2/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_2 vdd vss FILLER_0_2_2/VPW vdd FILLER_0_2_2/a_1916_375# FILLER_0_2_2/a_1380_472#
+ FILLER_0_2_2/a_3260_375# FILLER_0_2_2/a_36_472# FILLER_0_2_2/a_932_472# FILLER_0_2_2/a_2812_375#
+ FILLER_0_2_2/a_2276_472# FILLER_0_2_2/a_1828_472# FILLER_0_2_2/a_3172_472# FILLER_0_2_2/a_572_375#
+ FILLER_0_2_2/a_2724_472# FILLER_0_2_2/a_124_375# FILLER_0_2_2/a_1468_375# FILLER_0_2_2/a_1020_375#
+ FILLER_0_2_2/a_484_472# FILLER_0_2_2/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_3_12 vdd vss FILLER_0_3_12/VPW vdd FILLER_0_3_12/a_1916_375# FILLER_0_3_12/a_1380_472#
+ FILLER_0_3_12/a_3260_375# FILLER_0_3_12/a_36_472# FILLER_0_3_12/a_932_472# FILLER_0_3_12/a_2812_375#
+ FILLER_0_3_12/a_2276_472# FILLER_0_3_12/a_1828_472# FILLER_0_3_12/a_3172_472# FILLER_0_3_12/a_572_375#
+ FILLER_0_3_12/a_2724_472# FILLER_0_3_12/a_124_375# FILLER_0_3_12/a_1468_375# FILLER_0_3_12/a_1020_375#
+ FILLER_0_3_12/a_484_472# FILLER_0_3_12/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_9_66 vdd vss FILLER_0_9_66/VPW vdd FILLER_0_9_66/a_36_472# FILLER_0_9_66/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_11_ vss _11_/Z _11_/I vdd _11_/VPW vdd _11_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA_input7_I vss input_signal[6] vdd ANTENNA_input7_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_13_104 vdd vss FILLER_0_13_104/VPW vdd FILLER_0_13_104/a_36_472# FILLER_0_13_104/a_572_375#
+ FILLER_0_13_104/a_124_375# FILLER_0_13_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_12_37 vdd vss FILLER_0_12_37/VPW vdd FILLER_0_12_37/a_1916_375# FILLER_0_12_37/a_4516_472#
+ FILLER_0_12_37/a_1380_472# FILLER_0_12_37/a_3260_375# FILLER_0_12_37/a_5860_472#
+ FILLER_0_12_37/a_36_472# FILLER_0_12_37/a_932_472# FILLER_0_12_37/a_2812_375# FILLER_0_12_37/a_5412_472#
+ FILLER_0_12_37/a_2276_472# FILLER_0_12_37/a_4156_375# FILLER_0_12_37/a_6756_472#
+ FILLER_0_12_37/a_1828_472# FILLER_0_12_37/a_3708_375# FILLER_0_12_37/a_3172_472#
+ FILLER_0_12_37/a_572_375# FILLER_0_12_37/a_6308_472# FILLER_0_12_37/a_5052_375#
+ FILLER_0_12_37/a_2724_472# FILLER_0_12_37/a_6396_375# FILLER_0_12_37/a_4604_375#
+ FILLER_0_12_37/a_124_375# FILLER_0_12_37/a_1468_375# FILLER_0_12_37/a_4068_472#
+ FILLER_0_12_37/a_5948_375# FILLER_0_12_37/a_3620_472# FILLER_0_12_37/a_1020_375#
+ FILLER_0_12_37/a_5500_375# FILLER_0_12_37/a_4964_472# FILLER_0_12_37/a_484_472#
+ FILLER_0_12_37/a_2364_375# FILLER_0_12_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_107 vdd vss FILLER_0_10_107/VPW vdd FILLER_0_10_107/a_1380_472# FILLER_0_10_107/a_36_472#
+ FILLER_0_10_107/a_932_472# FILLER_0_10_107/a_572_375# FILLER_0_10_107/a_124_375#
+ FILLER_0_10_107/a_1468_375# FILLER_0_10_107/a_1020_375# FILLER_0_10_107/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
X_10_ vss _10_/Z _10_/I vdd _10_/VPW vdd _10_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1$1
XFILLER_0_0_36 vdd vss FILLER_0_0_36/VPW vdd FILLER_0_0_36/a_1916_375# FILLER_0_0_36/a_1380_472#
+ FILLER_0_0_36/a_3260_375# FILLER_0_0_36/a_36_472# FILLER_0_0_36/a_932_472# FILLER_0_0_36/a_2812_375#
+ FILLER_0_0_36/a_2276_472# FILLER_0_0_36/a_1828_472# FILLER_0_0_36/a_3172_472# FILLER_0_0_36/a_572_375#
+ FILLER_0_0_36/a_2724_472# FILLER_0_0_36/a_124_375# FILLER_0_0_36/a_1468_375# FILLER_0_0_36/a_1020_375#
+ FILLER_0_0_36/a_484_472# FILLER_0_0_36/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_15_8 vdd vss FILLER_0_15_8/VPW vdd FILLER_0_15_8/a_1916_375# FILLER_0_15_8/a_1380_472#
+ FILLER_0_15_8/a_3260_375# FILLER_0_15_8/a_36_472# FILLER_0_15_8/a_932_472# FILLER_0_15_8/a_2812_375#
+ FILLER_0_15_8/a_2276_472# FILLER_0_15_8/a_1828_472# FILLER_0_15_8/a_3172_472# FILLER_0_15_8/a_572_375#
+ FILLER_0_15_8/a_2724_472# FILLER_0_15_8/a_124_375# FILLER_0_15_8/a_1468_375# FILLER_0_15_8/a_1020_375#
+ FILLER_0_15_8/a_484_472# FILLER_0_15_8/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_16_70 vdd vss FILLER_0_16_70/VPW vdd FILLER_0_16_70/a_36_472# FILLER_0_16_70/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_11_2 vdd vss FILLER_0_11_2/VPW vdd FILLER_0_11_2/a_1916_375# FILLER_0_11_2/a_4516_472#
+ FILLER_0_11_2/a_1380_472# FILLER_0_11_2/a_3260_375# FILLER_0_11_2/a_5860_472# FILLER_0_11_2/a_36_472#
+ FILLER_0_11_2/a_932_472# FILLER_0_11_2/a_2812_375# FILLER_0_11_2/a_5412_472# FILLER_0_11_2/a_2276_472#
+ FILLER_0_11_2/a_4156_375# FILLER_0_11_2/a_6756_472# FILLER_0_11_2/a_1828_472# FILLER_0_11_2/a_3708_375#
+ FILLER_0_11_2/a_3172_472# FILLER_0_11_2/a_572_375# FILLER_0_11_2/a_6308_472# FILLER_0_11_2/a_5052_375#
+ FILLER_0_11_2/a_2724_472# FILLER_0_11_2/a_6396_375# FILLER_0_11_2/a_4604_375# FILLER_0_11_2/a_124_375#
+ FILLER_0_11_2/a_1468_375# FILLER_0_11_2/a_4068_472# FILLER_0_11_2/a_5948_375# FILLER_0_11_2/a_3620_472#
+ FILLER_0_11_2/a_1020_375# FILLER_0_11_2/a_5500_375# FILLER_0_11_2/a_4964_472# FILLER_0_11_2/a_484_472#
+ FILLER_0_11_2/a_2364_375# FILLER_0_11_2/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_28 vdd vss FILLER_0_12_28/VPW vdd FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_16_104 vdd vss FILLER_0_16_104/VPW vdd FILLER_0_16_104/a_36_472# FILLER_0_16_104/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_8_101 vdd vss FILLER_0_8_101/VPW vdd FILLER_0_8_101/a_36_472# FILLER_0_8_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA_input5_I vss input_signal[4] vdd ANTENNA_input5_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_6_37 vdd vss FILLER_0_6_37/VPW vdd FILLER_0_6_37/a_1916_375# FILLER_0_6_37/a_4516_472#
+ FILLER_0_6_37/a_1380_472# FILLER_0_6_37/a_3260_375# FILLER_0_6_37/a_5860_472# FILLER_0_6_37/a_36_472#
+ FILLER_0_6_37/a_932_472# FILLER_0_6_37/a_2812_375# FILLER_0_6_37/a_5412_472# FILLER_0_6_37/a_2276_472#
+ FILLER_0_6_37/a_4156_375# FILLER_0_6_37/a_6756_472# FILLER_0_6_37/a_1828_472# FILLER_0_6_37/a_3708_375#
+ FILLER_0_6_37/a_3172_472# FILLER_0_6_37/a_572_375# FILLER_0_6_37/a_6308_472# FILLER_0_6_37/a_5052_375#
+ FILLER_0_6_37/a_2724_472# FILLER_0_6_37/a_6396_375# FILLER_0_6_37/a_4604_375# FILLER_0_6_37/a_124_375#
+ FILLER_0_6_37/a_1468_375# FILLER_0_6_37/a_4068_472# FILLER_0_6_37/a_5948_375# FILLER_0_6_37/a_3620_472#
+ FILLER_0_6_37/a_1020_375# FILLER_0_6_37/a_5500_375# FILLER_0_6_37/a_4964_472# FILLER_0_6_37/a_484_472#
+ FILLER_0_6_37/a_2364_375# FILLER_0_6_37/a_6844_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_104 vdd vss FILLER_0_5_104/VPW vdd FILLER_0_5_104/a_36_472# FILLER_0_5_104/a_572_375#
+ FILLER_0_5_104/a_124_375# FILLER_0_5_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_2_107 vdd vss FILLER_0_2_107/VPW vdd FILLER_0_2_107/a_1380_472# FILLER_0_2_107/a_36_472#
+ FILLER_0_2_107/a_932_472# FILLER_0_2_107/a_572_375# FILLER_0_2_107/a_124_375# FILLER_0_2_107/a_1468_375#
+ FILLER_0_2_107/a_1020_375# FILLER_0_2_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_13_72 vdd vss FILLER_0_13_72/VPW vdd FILLER_0_13_72/a_1916_375# FILLER_0_13_72/a_1380_472#
+ FILLER_0_13_72/a_3260_375# FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_932_472# FILLER_0_13_72/a_2812_375#
+ FILLER_0_13_72/a_2276_472# FILLER_0_13_72/a_1828_472# FILLER_0_13_72/a_3172_472#
+ FILLER_0_13_72/a_572_375# FILLER_0_13_72/a_2724_472# FILLER_0_13_72/a_124_375# FILLER_0_13_72/a_1468_375#
+ FILLER_0_13_72/a_1020_375# FILLER_0_13_72/a_484_472# FILLER_0_13_72/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XANTENNA__06__I vss _15_/I vdd ANTENNA__06__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XANTENNA__11__I vss _11_/I vdd ANTENNA__11__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_0_28 vdd vss FILLER_0_0_28/VPW vdd FILLER_0_0_28/a_36_472# FILLER_0_0_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_1_60 vdd vss FILLER_0_1_60/VPW vdd FILLER_0_1_60/a_36_472# FILLER_0_1_60/a_572_375#
+ FILLER_0_1_60/a_124_375# FILLER_0_1_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
Xoutput30 output_signal_plus[9] _19_/Z vdd vss output30/VPW vdd output30/a_224_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XANTENNA__14__I vss _14_/I vdd ANTENNA__14__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
C0 FILLER_0_4_37/a_4068_472# FILLER_0_5_72/a_124_375# 0.001723f
C1 FILLER_0_14_37/a_5412_472# vdd 0.006901f
C2 FILLER_0_4_37/a_4964_472# vdd 0.005164f
C3 FILLER_0_8_101/a_124_375# FILLER_0_9_72/a_3260_375# 0.026339f
C4 FILLER_0_3_12/a_3260_375# FILLER_0_4_37/a_484_472# 0.001597f
C5 FILLER_0_0_104/a_124_375# _01_/ZN 0.029999f
C6 _19_/I FILLER_0_15_8/a_2276_472# 0.00191f
C7 _17_/I FILLER_0_14_37/a_6844_375# 0.018729f
C8 _16_/I FILLER_0_13_72/a_1020_375# 0.006182f
C9 FILLER_0_14_37/a_5860_472# _17_/I 0.015502f
C10 FILLER_0_8_37/a_2724_472# vdd 0.009155f
C11 FILLER_0_9_2/a_4604_375# vdd 0.007327f
C12 FILLER_0_7_104/a_572_375# _03_/ZN 0.008517f
C13 _13_/I _14_/I 0.724249f
C14 output_signal_plus[8] output_signal_plus[0] 0.073184f
C15 FILLER_0_8_107/a_484_472# _14_/I 0.022901f
C16 FILLER_0_12_37/a_2724_472# FILLER_0_11_2/a_6756_472# 0.026657f
C17 _17_/Z _10_/Z 0.129159f
C18 _14_/I input5/a_36_113# 0.003003f
C19 _18_/I FILLER_0_16_18/a_932_472# 0.00191f
C20 FILLER_0_8_37/a_3708_375# vdd 0.021784f
C21 _15_/I FILLER_0_11_66/a_124_375# 0.007111f
C22 _12_/I FILLER_0_5_12/a_2276_472# 0.003915f
C23 FILLER_0_7_2/a_6844_375# FILLER_0_7_66/a_36_472# 0.086635f
C24 _17_/I FILLER_0_15_56/a_484_472# 0.004125f
C25 FILLER_0_7_2/a_1468_375# vdd -0.004303f
C26 FILLER_0_7_72/a_1020_375# FILLER_0_6_37/a_5052_375# 0.026339f
C27 _15_/I FILLER_0_10_37/a_5500_375# 0.018729f
C28 _07_/ZN output22/a_224_472# 0.058524f
C29 FILLER_0_12_37/a_5500_375# _16_/I 0.016091f
C30 FILLER_0_12_37/a_2812_375# FILLER_0_14_37/a_2724_472# 0.001512f
C31 FILLER_0_5_12/a_1916_375# _12_/I 0.001706f
C32 FILLER_0_3_60/a_572_375# FILLER_0_2_37/a_3172_472# 0.001723f
C33 _00_/ZN output_signal_plus[2] 0.044354f
C34 FILLER_0_6_37/a_5412_472# FILLER_0_5_72/a_1468_375# 0.001597f
C35 _18_/I output27/a_224_472# 0.176269f
C36 vdd FILLER_0_12_107/a_124_375# 0.01489f
C37 _18_/I FILLER_0_15_8/a_2276_472# 0.014431f
C38 _13_/Z FILLER_0_10_107/a_1468_375# 0.013159f
C39 output22/a_224_472# _11_/a_36_113# 0.002583f
C40 input1/a_36_113# vdd 0.102561f
C41 FILLER_0_16_70/a_36_472# FILLER_0_16_36/a_3260_375# 0.016748f
C42 FILLER_0_0_36/a_1468_375# vdd -0.00915f
C43 vdd FILLER_0_16_36/a_932_472# 0.00284f
C44 output21/a_224_472# _19_/I 0.051029f
C45 FILLER_0_6_2/a_1380_472# _13_/I 0.003872f
C46 _11_/I _12_/I 0.285453f
C47 FILLER_0_7_72/a_2276_472# _12_/I 0.004669f
C48 FILLER_0_7_66/a_124_375# _14_/I 0.008393f
C49 FILLER_0_1_12/a_124_375# vdd 0.001706f
C50 input_signal[2] vdd 0.32843f
C51 _11_/I output15/a_224_472# 0.08176f
C52 output_signal_plus[5] _18_/I 0.008007f
C53 _11_/I FILLER_0_4_37/a_572_375# 0.01418f
C54 FILLER_0_11_66/a_36_472# FILLER_0_12_37/a_3260_375# 0.001597f
C55 vdd FILLER_0_0_12/a_1020_375# -0.006653f
C56 vdd FILLER_0_5_72/a_1468_375# 0.007048f
C57 FILLER_0_14_37/a_1468_375# _17_/I 0.018729f
C58 _14_/Z output_signal_plus[2] 0.169713f
C59 input_signal[6] FILLER_0_11_2/a_572_375# 0.009765f
C60 _15_/a_36_113# vdd 0.118116f
C61 FILLER_0_10_107/a_36_472# FILLER_0_10_101/a_36_472# 0.003468f
C62 _07_/ZN _10_/I 0.002779f
C63 _13_/I FILLER_0_5_12/a_36_472# 0.027222f
C64 FILLER_0_8_28/a_36_472# FILLER_0_7_2/a_2812_375# 0.001543f
C65 FILLER_0_6_37/a_6756_472# _13_/I 0.004135f
C66 _18_/I FILLER_0_14_37/a_2364_375# 0.002015f
C67 input_signal[6] FILLER_0_12_12/a_124_375# 0.00628f
C68 FILLER_0_5_72/a_2812_375# FILLER_0_4_37/a_6844_375# 0.026339f
C69 FILLER_0_15_72/a_1020_375# FILLER_0_13_72/a_932_472# 0.001512f
C70 _13_/I FILLER_0_6_2/a_2724_472# 0.003872f
C71 _14_/I FILLER_0_9_2/a_3172_472# 0.004017f
C72 _18_/I FILLER_0_14_12/a_572_375# 0.001895f
C73 FILLER_0_12_12/a_1468_375# FILLER_0_14_12/a_1380_472# 0.0027f
C74 _18_/I FILLER_0_14_37/a_1380_472# 0.001526f
C75 FILLER_0_13_72/a_2364_375# _17_/I 0.006125f
C76 FILLER_0_5_12/a_1828_472# _12_/I 0.003872f
C77 _15_/I FILLER_0_12_37/a_932_472# 0.001368f
C78 output_signal_plus[7] vdd 0.303346f
C79 _16_/I FILLER_0_11_72/a_3620_472# 0.00769f
C80 FILLER_0_11_2/a_3172_472# FILLER_0_13_2/a_3260_375# 0.0027f
C81 _11_/I FILLER_0_3_104/a_124_375# 0.008393f
C82 _16_/I FILLER_0_10_37/a_2812_375# 0.002327f
C83 output22/a_224_472# FILLER_0_10_107/a_1380_472# 0.001007f
C84 _18_/I output21/a_224_472# 0.010936f
C85 FILLER_0_8_37/a_3172_472# FILLER_0_7_66/a_36_472# 0.026657f
C86 FILLER_0_16_70/a_36_472# vdd 0.115025f
C87 FILLER_0_7_2/a_3172_472# FILLER_0_9_2/a_3260_375# 0.0027f
C88 FILLER_0_10_37/a_1380_472# vdd 0.007845f
C89 FILLER_0_0_142/a_124_375# _01_/ZN 0.003537f
C90 FILLER_0_2_37/a_2364_375# FILLER_0_4_37/a_2276_472# 0.001512f
C91 FILLER_0_7_2/a_5860_472# _12_/I 0.004108f
C92 _13_/I FILLER_0_6_37/a_2812_375# 0.001706f
C93 FILLER_0_7_2/a_1380_472# _14_/I 0.008733f
C94 FILLER_0_13_2/a_932_472# vdd 0.011054f
C95 FILLER_0_11_136/a_36_472# _08_/ZN 0.020589f
C96 FILLER_0_2_2/a_2812_375# vdd 0.022556f
C97 FILLER_0_5_12/a_1916_375# FILLER_0_4_2/a_3172_472# 0.001684f
C98 FILLER_0_12_107/a_484_472# _16_/I 0.017477f
C99 FILLER_0_0_36/a_1020_375# vdd -0.011044f
C100 vdd FILLER_0_11_2/a_6396_375# 0.014009f
C101 _13_/I FILLER_0_6_107/a_124_375# 0.030385f
C102 FILLER_0_0_70/a_36_472# FILLER_0_0_36/a_3172_472# 0.003468f
C103 FILLER_0_1_60/a_124_375# vdd -0.002461f
C104 FILLER_0_10_37/a_2364_375# FILLER_0_12_37/a_2276_472# 0.001512f
C105 _16_/I FILLER_0_11_2/a_4964_472# 0.007542f
C106 FILLER_0_0_28/a_124_375# vdd 0.014408f
C107 FILLER_0_15_72/a_1380_472# vdd 0.004859f
C108 FILLER_0_13_104/a_124_375# _16_/I 0.006313f
C109 FILLER_0_12_37/a_124_375# _16_/I 0.016401f
C110 vdd FILLER_0_8_37/a_4604_375# 0.004103f
C111 FILLER_0_13_2/a_4964_472# FILLER_0_12_37/a_1020_375# 0.001723f
C112 _10_/Z FILLER_0_11_72/a_6756_472# 0.01497f
C113 _11_/I FILLER_0_4_2/a_3172_472# 0.014431f
C114 input8/a_36_113# vdd 0.120837f
C115 output12/a_224_472# _13_/Z 0.03322f
C116 FILLER_0_14_12/a_932_472# _17_/I 0.015529f
C117 FILLER_0_10_107/a_1020_375# FILLER_0_12_107/a_932_472# 0.001512f
C118 output_signal_plus[3] output_signal_plus[2] 0.22563f
C119 FILLER_0_10_37/a_572_375# FILLER_0_11_2/a_4516_472# 0.001723f
C120 _02_/ZN _12_/a_36_113# 0.146173f
C121 FILLER_0_11_2/a_5412_472# FILLER_0_12_37/a_1380_472# 0.026657f
C122 _08_/ZN output14/a_224_472# 0.061002f
C123 FILLER_0_2_2/a_3172_472# vdd 0.014746f
C124 FILLER_0_14_37/a_4964_472# FILLER_0_15_72/a_1020_375# 0.001723f
C125 FILLER_0_13_2/a_1380_472# _17_/I 0.00656f
C126 FILLER_0_9_2/a_1916_375# FILLER_0_8_12/a_932_472# 0.001684f
C127 _11_/I FILLER_0_5_12/a_1380_472# 0.001913f
C128 _19_/Z output_signal_plus[0] 0.056517f
C129 _15_/I FILLER_0_11_2/a_4516_472# 0.005458f
C130 _19_/I output_signal_plus[6] 0.00787f
C131 FILLER_0_6_37/a_1468_375# vdd 0.008961f
C132 _02_/ZN _12_/Z 0.031232f
C133 FILLER_0_12_28/a_124_375# FILLER_0_13_2/a_3172_472# 0.001684f
C134 FILLER_0_4_2/a_572_375# _12_/I 0.027023f
C135 _11_/I FILLER_0_4_37/a_124_375# 0.01418f
C136 _19_/I FILLER_0_15_40/a_484_472# 0.001782f
C137 input2/a_36_113# input1/a_36_113# 0.029417f
C138 _16_/I FILLER_0_11_72/a_5860_472# 0.00769f
C139 _15_/I FILLER_0_10_37/a_4068_472# 0.015502f
C140 _11_/I output19/a_224_472# 0.042992f
C141 _13_/Z _16_/I 0.003263f
C142 FILLER_0_9_2/a_1020_375# FILLER_0_8_12/a_36_472# 0.001684f
C143 _12_/I FILLER_0_6_37/a_1916_375# 0.016091f
C144 FILLER_0_6_37/a_4604_375# _12_/I 0.016091f
C145 output12/a_224_472# _14_/I 0.061774f
C146 output_signal_plus[5] _16_/a_36_113# 0.012925f
C147 _16_/I FILLER_0_11_72/a_2812_375# 0.007169f
C148 FILLER_0_4_2/a_1020_375# _12_/I 0.007331f
C149 _14_/I FILLER_0_8_12/a_36_472# 0.024093f
C150 input2/a_36_113# input_signal[2] 0.003542f
C151 input2/a_36_113# FILLER_0_1_12/a_124_375# 0.002124f
C152 _13_/I output16/a_224_472# 0.090122f
C153 vdd FILLER_0_1_12/a_932_472# 0.019027f
C154 output_signal_plus[8] _19_/Z 0.603273f
C155 _17_/I input_signal[8] 0.002921f
C156 _09_/ZN FILLER_0_12_107/a_124_375# 0.002085f
C157 FILLER_0_3_44/a_484_472# vdd 0.007487f
C158 FILLER_0_15_8/a_124_375# input_signal[8] 0.010194f
C159 FILLER_0_16_36/a_36_472# _19_/I 0.014431f
C160 FILLER_0_16_70/a_124_375# output30/a_224_472# 0.011959f
C161 _18_/I output_signal_plus[6] 0.334772f
C162 vdd FILLER_0_4_107/a_36_472# 0.110317f
C163 _18_/I FILLER_0_14_37/a_6396_375# 0.001895f
C164 _18_/I FILLER_0_14_37/a_4604_375# 0.003988f
C165 output20/a_224_472# FILLER_0_2_37/a_5412_472# 0.001058f
C166 FILLER_0_2_107/a_1380_472# _01_/ZN 0.005185f
C167 _18_/I FILLER_0_15_40/a_124_375# 0.01418f
C168 vdd FILLER_0_10_37/a_2724_472# 0.009656f
C169 _18_/I FILLER_0_15_40/a_484_472# 0.014431f
C170 FILLER_0_8_37/a_1916_375# FILLER_0_9_2/a_5948_375# 0.026339f
C171 FILLER_0_9_2/a_6756_472# FILLER_0_10_37/a_2724_472# 0.026657f
C172 FILLER_0_6_107/a_36_472# FILLER_0_6_101/a_124_375# 0.016748f
C173 _16_/I FILLER_0_10_12/a_124_375# 0.002327f
C174 FILLER_0_11_72/a_572_375# FILLER_0_10_37/a_4516_472# 0.001723f
C175 FILLER_0_2_37/a_932_472# FILLER_0_3_44/a_124_375# 0.001723f
C176 FILLER_0_6_37/a_484_472# vdd 0.004058f
C177 _00_/ZN _11_/I 0.456826f
C178 FILLER_0_16_36/a_2364_375# vdd 0.039333f
C179 vdd FILLER_0_7_2/a_1916_375# 0.017563f
C180 FILLER_0_3_72/a_3172_472# FILLER_0_3_104/a_36_472# 0.013276f
C181 input_signal[3] FILLER_0_5_12/a_572_375# 0.00242f
C182 FILLER_0_13_72/a_1468_375# _17_/I 0.006125f
C183 FILLER_0_10_37/a_1916_375# FILLER_0_12_37/a_1828_472# 0.001512f
C184 FILLER_0_3_44/a_1380_472# FILLER_0_3_60/a_36_472# 0.013276f
C185 FILLER_0_8_101/a_36_472# FILLER_0_6_101/a_124_375# 0.001512f
C186 _16_/I FILLER_0_11_72/a_4964_472# 0.006098f
C187 FILLER_0_2_2/a_2724_472# vdd 0.011159f
C188 FILLER_0_12_12/a_36_472# FILLER_0_11_2/a_1020_375# 0.001543f
C189 _15_/I output23/a_224_472# 0.035533f
C190 FILLER_0_4_37/a_5860_472# vdd 0.008331f
C191 FILLER_0_11_136/a_36_472# vdd 0.099264f
C192 FILLER_0_0_142/a_36_472# _01_/ZN 0.001973f
C193 FILLER_0_12_107/a_1380_472# output_signal_plus[4] 0.001294f
C194 _15_/I FILLER_0_9_104/a_124_375# 0.006125f
C195 _09_/ZN output_signal_plus[7] 0.210079f
C196 FILLER_0_11_72/a_1916_375# FILLER_0_12_37/a_5860_472# 0.001597f
C197 _17_/Z output_signal_plus[4] 0.002877f
C198 vdd FILLER_0_2_2/a_124_375# 0.012786f
C199 FILLER_0_11_136/a_124_375# _10_/Z 0.002831f
C200 FILLER_0_0_28/a_124_375# FILLER_0_1_12/a_1916_375# 0.05841f
C201 output_signal_minus[7] _06_/ZN 0.005232f
C202 output_signal_minus[9] output_signal_minus[0] 0.65109f
C203 _16_/I FILLER_0_13_2/a_3620_472# 0.004669f
C204 input6/a_36_113# vdd 0.120999f
C205 FILLER_0_2_101/a_36_472# vdd 0.096264f
C206 _10_/a_36_160# output_signal_minus[7] 0.024955f
C207 FILLER_0_9_72/a_572_375# FILLER_0_8_37/a_4604_375# 0.026339f
C208 input1/a_36_113# input_signal[1] 0.045824f
C209 FILLER_0_8_37/a_4068_472# FILLER_0_7_72/a_124_375# 0.001597f
C210 vdd FILLER_0_3_72/a_1828_472# 0.008296f
C211 output_signal_minus[6] _10_/Z 0.491295f
C212 FILLER_0_0_28/a_124_375# FILLER_0_0_36/a_36_472# 0.009654f
C213 _13_/I FILLER_0_5_44/a_124_375# 0.016091f
C214 vdd output14/a_224_472# 0.059712f
C215 FILLER_0_1_12/a_1380_472# vdd 0.01093f
C216 FILLER_0_3_60/a_572_375# FILLER_0_4_37/a_3172_472# 0.001597f
C217 FILLER_0_4_37/a_6756_472# FILLER_0_2_37/a_6844_375# 0.001512f
C218 vdd FILLER_0_5_72/a_1020_375# 0.005487f
C219 FILLER_0_2_2/a_3172_472# FILLER_0_1_12/a_1916_375# 0.001543f
C220 _11_/I FILLER_0_2_37/a_6756_472# 0.002136f
C221 FILLER_0_11_66/a_124_375# FILLER_0_10_37/a_3260_375# 0.026339f
C222 input_signal[2] input_signal[1] 0.055021f
C223 _11_/I FILLER_0_4_107/a_124_375# 0.01418f
C224 FILLER_0_1_12/a_124_375# input_signal[1] 0.009861f
C225 output26/a_224_472# _10_/Z 0.083702f
C226 FILLER_0_12_37/a_5412_472# vdd 0.00624f
C227 FILLER_0_11_2/a_5412_472# FILLER_0_13_2/a_5500_375# 0.001512f
C228 _13_/I FILLER_0_6_2/a_1828_472# 0.003872f
C229 FILLER_0_14_12/a_484_472# FILLER_0_13_2/a_1468_375# 0.001543f
C230 _16_/I FILLER_0_12_28/a_36_472# 0.018008f
C231 _15_/I FILLER_0_11_72/a_4068_472# 0.005458f
C232 FILLER_0_8_107/a_124_375# FILLER_0_9_104/a_484_472# 0.001723f
C233 FILLER_0_1_60/a_484_472# vdd 0.013043f
C234 FILLER_0_9_66/a_36_472# _15_/I 0.006506f
C235 _12_/a_36_113# _12_/I 0.010925f
C236 FILLER_0_3_72/a_3260_375# FILLER_0_2_101/a_36_472# 0.001723f
C237 FILLER_0_16_36/a_2812_375# _19_/I 0.017849f
C238 FILLER_0_12_37/a_4604_375# _16_/I 0.016091f
C239 FILLER_0_11_2/a_5948_375# _16_/I 0.007169f
C240 _16_/I FILLER_0_13_2/a_2276_472# 0.004669f
C241 FILLER_0_3_60/a_124_375# FILLER_0_1_60/a_36_472# 0.001512f
C242 FILLER_0_10_37/a_4964_472# FILLER_0_11_72/a_1020_375# 0.001723f
C243 FILLER_0_2_2/a_1020_375# FILLER_0_3_12/a_36_472# 0.001684f
C244 FILLER_0_2_2/a_1468_375# _10_/I 0.001886f
C245 _11_/I FILLER_0_3_44/a_572_375# 0.008393f
C246 _13_/I FILLER_0_6_37/a_2364_375# 0.001706f
C247 FILLER_0_4_37/a_124_375# FILLER_0_4_2/a_3260_375# 0.004426f
C248 FILLER_0_12_107/a_1468_375# _16_/I 0.01484f
C249 _12_/Z _12_/I 0.166374f
C250 FILLER_0_13_66/a_36_472# _17_/I 0.006506f
C251 input_signal[2] input_signal[3] 0.006057f
C252 output15/a_224_472# _12_/Z 0.004357f
C253 FILLER_0_5_104/a_572_375# output_signal_minus[4] 0.011852f
C254 FILLER_0_11_2/a_4068_472# _15_/I 0.005458f
C255 FILLER_0_9_72/a_3172_472# vdd 0.009151f
C256 _17_/a_36_113# output_signal_plus[7] 0.009958f
C257 FILLER_0_16_104/a_36_472# vdd 0.114072f
C258 FILLER_0_10_12/a_1380_472# vdd 0.010304f
C259 FILLER_0_5_12/a_3260_375# FILLER_0_3_12/a_3172_472# 0.001512f
C260 FILLER_0_9_2/a_4516_472# _14_/I 0.004017f
C261 FILLER_0_4_37/a_484_472# _13_/I 0.003497f
C262 FILLER_0_14_28/a_36_472# FILLER_0_14_37/a_36_472# 0.001963f
C263 FILLER_0_11_2/a_2364_375# FILLER_0_9_2/a_2276_472# 0.0027f
C264 FILLER_0_10_12/a_1468_375# _15_/I 0.018729f
C265 FILLER_0_1_72/a_484_472# vdd 0.002467f
C266 FILLER_0_12_28/a_124_375# vdd 0.046667f
C267 _19_/I FILLER_0_16_36/a_1380_472# 0.015152f
C268 _15_/I FILLER_0_8_37/a_2364_375# 0.001237f
C269 _18_/I FILLER_0_16_36/a_2812_375# 0.00153f
C270 FILLER_0_16_70/a_124_375# FILLER_0_15_72/a_36_472# 0.001543f
C271 _14_/I FILLER_0_9_72/a_1020_375# 0.005381f
C272 _08_/ZN _01_/ZN 0.319133f
C273 _09_/ZN FILLER_0_4_107/a_36_472# 0.002542f
C274 FILLER_0_16_70/a_36_472# output30/a_224_472# 0.003196f
C275 _17_/I FILLER_0_14_37/a_2724_472# 0.015502f
C276 _07_/ZN _13_/Z 0.041654f
C277 FILLER_0_15_8/a_2724_472# FILLER_0_16_18/a_1468_375# 0.001543f
C278 _17_/Z _17_/I 0.074565f
C279 FILLER_0_14_107/a_124_375# vdd 0.01514f
C280 output_signal_plus[4] FILLER_0_11_72/a_6756_472# 0.001108f
C281 FILLER_0_14_101/a_124_375# FILLER_0_14_37/a_6844_375# 0.012001f
C282 FILLER_0_15_72/a_572_375# FILLER_0_14_37/a_4516_472# 0.001723f
C283 _16_/I FILLER_0_11_66/a_124_375# 0.007169f
C284 _16_/I FILLER_0_10_37/a_5500_375# 0.002327f
C285 FILLER_0_10_37/a_3708_375# FILLER_0_12_37/a_3620_472# 0.0027f
C286 vdd FILLER_0_11_2/a_932_472# 0.009688f
C287 FILLER_0_10_37/a_2276_472# FILLER_0_9_2/a_6308_472# 0.026657f
C288 FILLER_0_1_12/a_3172_472# _10_/I 0.006408f
C289 FILLER_0_14_12/a_1468_375# FILLER_0_13_2/a_2724_472# 0.001543f
C290 input_signal[0] FILLER_0_0_12/a_36_472# 0.076453f
C291 FILLER_0_6_37/a_1468_375# FILLER_0_7_2/a_5500_375# 0.026339f
C292 vdd FILLER_0_6_37/a_572_375# 0.005339f
C293 FILLER_0_7_2/a_6844_375# _12_/I 0.006193f
C294 FILLER_0_15_72/a_1380_472# output30/a_224_472# 0.038484f
C295 _19_/I FILLER_0_16_18/a_1380_472# 0.014431f
C296 FILLER_0_8_37/a_1828_472# vdd 0.009805f
C297 FILLER_0_6_37/a_1020_375# FILLER_0_7_2/a_5052_375# 0.026339f
C298 FILLER_0_15_2/a_36_472# input_signal[8] 0.011959f
C299 FILLER_0_10_37/a_6844_375# FILLER_0_12_37/a_6756_472# 0.001512f
C300 _13_/Z _11_/a_36_113# 0.018722f
C301 _15_/I FILLER_0_10_37/a_572_375# 0.018729f
C302 FILLER_0_8_28/a_36_472# FILLER_0_9_2/a_2812_375# 0.001684f
C303 FILLER_0_12_37/a_5948_375# vdd 0.011644f
C304 _18_/I FILLER_0_16_36/a_1380_472# 0.001782f
C305 FILLER_0_4_2/a_2276_472# vdd 0.011739f
C306 _16_/I FILLER_0_13_104/a_572_375# 0.006193f
C307 FILLER_0_13_66/a_36_472# FILLER_0_12_37/a_3260_375# 0.001723f
C308 vdd FILLER_0_3_44/a_1020_375# 0.011772f
C309 _07_/ZN _14_/I 0.084253f
C310 FILLER_0_2_37/a_3708_375# _10_/I 0.001886f
C311 FILLER_0_2_37/a_484_472# vdd 0.005213f
C312 FILLER_0_4_37/a_2812_375# vdd 0.010742f
C313 FILLER_0_15_8/a_1916_375# _18_/I 0.014209f
C314 FILLER_0_1_12/a_2724_472# FILLER_0_3_12/a_2812_375# 0.001512f
C315 FILLER_0_7_2/a_3172_472# FILLER_0_8_28/a_124_375# 0.001543f
C316 _08_/ZN _16_/Z 0.013653f
C317 FILLER_0_11_72/a_2724_472# vdd 0.034098f
C318 FILLER_0_2_37/a_1380_472# _10_/I 0.002525f
C319 FILLER_0_12_37/a_572_375# FILLER_0_11_2/a_4516_472# 0.001597f
C320 _11_/I FILLER_0_4_37/a_6844_375# 0.01418f
C321 FILLER_0_14_37/a_5500_375# vdd 0.008584f
C322 FILLER_0_7_2/a_572_375# _14_/I 0.008393f
C323 vdd FILLER_0_5_72/a_3260_375# 0.009973f
C324 FILLER_0_8_37/a_4516_472# FILLER_0_6_37/a_4604_375# 0.001512f
C325 vdd FILLER_0_3_72/a_36_472# 0.109729f
C326 FILLER_0_6_2/a_2276_472# vdd 0.011126f
C327 _14_/I _11_/a_36_113# 0.004347f
C328 FILLER_0_0_28/a_124_375# FILLER_0_0_36/a_124_375# 0.003732f
C329 FILLER_0_7_2/a_1020_375# _12_/I 0.006134f
C330 _11_/I _13_/a_36_113# 0.050389f
C331 _18_/I FILLER_0_16_18/a_1380_472# 0.00191f
C332 FILLER_0_9_72/a_2812_375# FILLER_0_7_72/a_2724_472# 0.001512f
C333 FILLER_0_4_37/a_1380_472# FILLER_0_3_44/a_484_472# 0.026657f
C334 vdd FILLER_0_13_72/a_2724_472# 0.034847f
C335 FILLER_0_7_72/a_36_472# FILLER_0_7_66/a_124_375# 0.016748f
C336 FILLER_0_10_107/a_1380_472# _13_/Z 0.003128f
C337 vdd FILLER_0_9_2/a_5860_472# 0.017113f
C338 _11_/I output_signal_minus[5] 0.078891f
C339 FILLER_0_11_2/a_6308_472# FILLER_0_12_37/a_2364_375# 0.001597f
C340 FILLER_0_2_37/a_2724_472# FILLER_0_1_60/a_36_472# 0.026657f
C341 _13_/I FILLER_0_6_101/a_36_472# 0.005434f
C342 FILLER_0_15_8/a_1916_375# FILLER_0_14_12/a_1468_375# 0.05841f
C343 _13_/I FILLER_0_6_37/a_5860_472# 0.003818f
C344 FILLER_0_8_37/a_5948_375# vdd 0.011562f
C345 _18_/I FILLER_0_15_40/a_572_375# 0.01418f
C346 _16_/I FILLER_0_12_37/a_932_472# 0.017477f
C347 FILLER_0_9_2/a_1916_375# _14_/I 0.002004f
C348 output20/a_224_472# output_signal_minus[0] 0.013919f
C349 FILLER_0_15_8/a_3172_472# FILLER_0_16_36/a_36_472# 0.058411f
C350 FILLER_0_1_12/a_1020_375# FILLER_0_0_12/a_1020_375# 0.05841f
C351 FILLER_0_1_12/a_3260_375# _10_/I 0.008103f
C352 FILLER_0_14_37/a_6756_472# vdd 0.015534f
C353 _19_/I _18_/Z 1.423466f
C354 FILLER_0_7_2/a_4516_472# _12_/I 0.004669f
C355 _14_/I FILLER_0_8_37/a_932_472# 0.014431f
C356 FILLER_0_8_37/a_4068_472# _14_/I 0.014431f
C357 FILLER_0_10_28/a_124_375# FILLER_0_12_28/a_36_472# 0.0027f
C358 vdd FILLER_0_12_37/a_1020_375# 0.006813f
C359 FILLER_0_3_60/a_572_375# FILLER_0_3_72/a_124_375# 0.003732f
C360 FILLER_0_7_104/a_484_472# FILLER_0_8_107/a_36_472# 0.026657f
C361 _11_/I FILLER_0_2_37/a_3172_472# 0.002415f
C362 _14_/I FILLER_0_8_12/a_572_375# 0.014268f
C363 FILLER_0_2_37/a_4964_472# _10_/I 0.002486f
C364 input_signal[1] FILLER_0_2_2/a_124_375# 0.005045f
C365 FILLER_0_6_37/a_1020_375# _12_/I 0.016091f
C366 FILLER_0_6_37/a_4516_472# FILLER_0_5_72/a_572_375# 0.001597f
C367 _00_/ZN _12_/Z 0.006032f
C368 vdd _01_/ZN 0.423997f
C369 _15_/I FILLER_0_11_2/a_5500_375# 0.007111f
C370 FILLER_0_6_37/a_932_472# _12_/I 0.017477f
C371 FILLER_0_0_36/a_2812_375# vdd -0.007824f
C372 _11_/I FILLER_0_5_12/a_484_472# 0.001838f
C373 FILLER_0_16_70/a_124_375# _19_/I 0.018946f
C374 vdd FILLER_0_10_37/a_3172_472# 0.007139f
C375 output25/a_224_472# output24/a_224_472# 0.007f
C376 FILLER_0_10_37/a_6308_472# FILLER_0_9_72/a_2364_375# 0.001597f
C377 _11_/I FILLER_0_3_12/a_932_472# 0.00942f
C378 _13_/I FILLER_0_5_72/a_572_375# 0.016091f
C379 vdd FILLER_0_7_72/a_1380_472# 0.006325f
C380 FILLER_0_12_12/a_484_472# vdd 0.021419f
C381 FILLER_0_2_2/a_1380_472# FILLER_0_1_12/a_124_375# 0.001543f
C382 _18_/I _18_/Z 0.382716f
C383 FILLER_0_3_72/a_932_472# vdd 0.004803f
C384 FILLER_0_4_107/a_36_472# FILLER_0_4_101/a_124_375# 0.016748f
C385 FILLER_0_4_37/a_3172_472# FILLER_0_5_60/a_572_375# 0.001723f
C386 output_signal_minus[1] _13_/Z 0.029294f
C387 input_signal[5] input6/a_36_113# 0.026766f
C388 _11_/I FILLER_0_2_37/a_5860_472# 0.002415f
C389 _16_/I FILLER_0_11_2/a_4516_472# 0.007542f
C390 _15_/I FILLER_0_10_37/a_1468_375# 0.018729f
C391 _14_/Z _12_/Z 0.187331f
C392 FILLER_0_13_2/a_1020_375# _16_/I 0.006277f
C393 vdd FILLER_0_14_12/a_36_472# 0.015471f
C394 output29/a_224_472# FILLER_0_14_37/a_5948_375# 0.029497f
C395 FILLER_0_3_72/a_572_375# FILLER_0_2_37/a_4604_375# 0.026339f
C396 output19/a_224_472# FILLER_0_4_107/a_1380_472# 0.001007f
C397 vdd FILLER_0_1_72/a_36_472# 0.109729f
C398 _11_/I FILLER_0_4_37/a_3708_375# 0.01418f
C399 FILLER_0_6_37/a_1380_472# _13_/I 0.003818f
C400 FILLER_0_16_70/a_124_375# _18_/I 0.001989f
C401 FILLER_0_14_115/a_124_375# output27/a_224_472# 0.029497f
C402 FILLER_0_15_56/a_572_375# _17_/I 0.006589f
C403 FILLER_0_13_2/a_1828_472# vdd 0.048546f
C404 FILLER_0_7_72/a_1020_375# FILLER_0_8_37/a_4964_472# 0.001597f
C405 FILLER_0_15_40/a_1020_375# FILLER_0_14_37/a_1380_472# 0.001723f
C406 _16_/Z vdd 0.351819f
C407 FILLER_0_7_66/a_36_472# FILLER_0_9_66/a_124_375# 0.001512f
C408 output19/a_224_472# output_signal_minus[6] 0.007827f
C409 FILLER_0_6_107/a_36_472# vdd 0.112159f
C410 FILLER_0_16_36/a_3172_472# vdd 0.010244f
C411 FILLER_0_1_12/a_484_472# _11_/I 0.001094f
C412 net15 output_signal_minus[4] 0.045791f
C413 FILLER_0_11_72/a_5500_375# _10_/Z 0.001594f
C414 FILLER_0_3_60/a_484_472# FILLER_0_5_60/a_572_375# 0.001512f
C415 _11_/I FILLER_0_4_107/a_1468_375# 0.118948f
C416 _11_/I _03_/ZN 0.0092f
C417 FILLER_0_7_2/a_3620_472# _14_/I 0.008761f
C418 output_signal_minus[1] _14_/I 0.332908f
C419 FILLER_0_9_72/a_1468_375# FILLER_0_7_72/a_1380_472# 0.001512f
C420 FILLER_0_7_2/a_4156_375# FILLER_0_6_37/a_124_375# 0.026339f
C421 _18_/I FILLER_0_15_72/a_1020_375# 0.01418f
C422 FILLER_0_13_104/a_124_375# FILLER_0_13_72/a_3260_375# 0.012222f
C423 _13_/I FILLER_0_5_60/a_124_375# 0.016091f
C424 FILLER_0_15_8/a_3260_375# _18_/I 0.01418f
C425 vdd FILLER_0_8_101/a_36_472# 0.098287f
C426 output12/a_224_472# output23/a_224_472# 0.005712f
C427 FILLER_0_9_66/a_36_472# FILLER_0_10_37/a_3260_375# 0.001597f
C428 _11_/I FILLER_0_5_12/a_3260_375# 0.004712f
C429 output17/a_224_472# _01_/ZN 0.128071f
C430 vdd FILLER_0_5_44/a_484_472# 0.007356f
C431 _12_/I FILLER_0_7_72/a_1828_472# 0.004669f
C432 _14_/I FILLER_0_9_2/a_6844_375# 0.005381f
C433 FILLER_0_13_2/a_932_472# input_signal[7] 0.00143f
C434 FILLER_0_14_37/a_1468_375# FILLER_0_13_2/a_5412_472# 0.001597f
C435 _15_/I FILLER_0_9_2/a_484_472# 0.003226f
C436 FILLER_0_8_107/a_36_472# vdd 0.110317f
C437 _11_/Z vdd 0.193304f
C438 FILLER_0_14_37/a_5412_472# _18_/I 0.001526f
C439 FILLER_0_16_104/a_36_472# output30/a_224_472# 0.003176f
C440 _07_/ZN output16/a_224_472# 0.212108f
C441 vdd FILLER_0_6_37/a_3620_472# 0.007765f
C442 vdd FILLER_0_12_12/a_1380_472# 0.009391f
C443 FILLER_0_8_37/a_1916_375# vdd 0.015167f
C444 FILLER_0_7_2/a_5948_375# _12_/I 0.003867f
C445 FILLER_0_5_44/a_1468_375# vdd 0.043784f
C446 FILLER_0_11_2/a_5500_375# FILLER_0_10_37/a_1468_375# 0.026339f
C447 _11_/I FILLER_0_3_12/a_2364_375# 0.008393f
C448 _00_/ZN output_signal_minus[6] 0.0465f
C449 input8/a_36_113# input_signal[7] 0.02969f
C450 _19_/I FILLER_0_16_36/a_932_472# 0.014431f
C451 FILLER_0_8_37/a_6844_375# vdd 0.013417f
C452 FILLER_0_5_44/a_932_472# _11_/I 0.001913f
C453 _18_/a_36_113# _18_/Z 0.002435f
C454 FILLER_0_7_72/a_572_375# _12_/I 0.006182f
C455 _00_/ZN output26/a_224_472# 0.015084f
C456 FILLER_0_11_2/a_124_375# vdd 0.012902f
C457 _14_/I FILLER_0_9_72/a_2364_375# 0.004454f
C458 _11_/I FILLER_0_5_72/a_1916_375# 0.004712f
C459 _11_/I FILLER_0_4_2/a_1916_375# 0.01433f
C460 FILLER_0_3_72/a_2812_375# vdd 0.019956f
C461 FILLER_0_16_36/a_1468_375# vdd 0.005783f
C462 FILLER_0_12_37/a_36_472# FILLER_0_12_28/a_36_472# 0.001963f
C463 _10_/Z FILLER_0_11_72/a_6308_472# 0.036527f
C464 FILLER_0_2_37/a_6308_472# vdd 0.019321f
C465 _11_/I _06_/ZN 0.391549f
C466 _14_/I FILLER_0_8_12/a_1380_472# 0.014431f
C467 FILLER_0_3_60/a_36_472# FILLER_0_5_60/a_124_375# 0.001512f
C468 FILLER_0_13_72/a_1828_472# _16_/I 0.004669f
C469 FILLER_0_13_2/a_1916_375# vdd 0.051099f
C470 _15_/I FILLER_0_9_2/a_3172_472# 0.006606f
C471 _09_/ZN _01_/ZN 0.003503f
C472 _15_/I FILLER_0_10_107/a_1468_375# 0.017398f
C473 output_signal_plus[7] _19_/I 0.455107f
C474 FILLER_0_10_37/a_6756_472# vdd 0.015534f
C475 FILLER_0_0_142/a_572_375# output_signal_minus[7] 0.006638f
C476 FILLER_0_13_72/a_572_375# FILLER_0_11_72/a_484_472# 0.001512f
C477 _11_/Z output13/a_224_472# 0.00187f
C478 _11_/I FILLER_0_2_37/a_572_375# 0.00346f
C479 _11_/I FILLER_0_2_37/a_4068_472# 0.002301f
C480 _18_/I FILLER_0_16_36/a_932_472# 0.001782f
C481 FILLER_0_8_37/a_1380_472# vdd 0.007309f
C482 FILLER_0_16_70/a_36_472# _19_/I 0.020196f
C483 _17_/I output26/a_224_472# 0.176642f
C484 _16_/I FILLER_0_11_72/a_4068_472# 0.007542f
C485 output24/a_224_472# _15_/Z 0.052418f
C486 FILLER_0_5_60/a_36_472# _13_/I 0.017477f
C487 _11_/I FILLER_0_3_72/a_484_472# 0.002089f
C488 vdd FILLER_0_1_72/a_1020_375# 0.004358f
C489 FILLER_0_5_104/a_572_375# _12_/I 0.001706f
C490 _11_/I output_signal_minus[3] 0.086977f
C491 _11_/I FILLER_0_4_107/a_572_375# 0.01418f
C492 input_signal[2] FILLER_0_2_2/a_36_472# 0.011205f
C493 FILLER_0_5_104/a_572_375# output15/a_224_472# 0.011959f
C494 input10/a_36_113# input8/a_36_113# 0.001442f
C495 _15_/I FILLER_0_10_37/a_3260_375# 0.018729f
C496 output_signal_minus[7] FILLER_0_0_104/a_124_375# 0.011852f
C497 FILLER_0_6_2/a_3172_472# vdd 0.012828f
C498 FILLER_0_14_37/a_5500_375# output30/a_224_472# 0.001234f
C499 FILLER_0_15_72/a_1380_472# _19_/I 0.001641f
C500 output22/a_224_472# _15_/a_36_113# 0.006255f
C501 output_signal_plus[3] FILLER_0_11_136/a_124_375# 0.001077f
C502 FILLER_0_10_37/a_2364_375# vdd 0.025298f
C503 FILLER_0_4_2/a_36_472# vdd 0.105578f
C504 FILLER_0_11_2/a_4068_472# _16_/I 0.003315f
C505 output_signal_plus[7] _18_/I 0.679572f
C506 FILLER_0_13_2/a_2364_375# FILLER_0_12_12/a_1380_472# 0.001684f
C507 FILLER_0_0_36/a_1916_375# FILLER_0_1_44/a_1020_375# 0.05841f
C508 _13_/I FILLER_0_6_37/a_4516_472# 0.003481f
C509 _12_/I FILLER_0_6_2/a_3260_375# 0.017617f
C510 FILLER_0_1_44/a_1380_472# FILLER_0_1_60/a_36_472# 0.013276f
C511 FILLER_0_2_37/a_1916_375# FILLER_0_3_44/a_1020_375# 0.026339f
C512 FILLER_0_14_115/a_124_375# output_signal_plus[6] 0.001313f
C513 FILLER_0_8_12/a_124_375# _14_/I 0.014501f
C514 FILLER_0_16_70/a_36_472# _18_/I 0.004265f
C515 FILLER_0_13_66/a_36_472# FILLER_0_13_2/a_6756_472# 0.013277f
C516 output11/a_224_472# FILLER_0_2_101/a_36_472# 0.031813f
C517 FILLER_0_5_44/a_124_375# FILLER_0_3_44/a_36_472# 0.001512f
C518 FILLER_0_10_12/a_1468_375# _16_/I 0.002327f
C519 FILLER_0_12_12/a_1468_375# FILLER_0_11_2/a_2724_472# 0.001543f
C520 vdd FILLER_0_7_104/a_124_375# 0.027844f
C521 input1/a_36_113# _10_/I 0.018904f
C522 vdd FILLER_0_9_72/a_1916_375# 0.009597f
C523 FILLER_0_2_2/a_1916_375# FILLER_0_3_12/a_932_472# 0.001684f
C524 FILLER_0_0_36/a_1468_375# _10_/I 0.015932f
C525 input4/a_36_113# FILLER_0_5_12/a_124_375# 0.002124f
C526 _11_/I FILLER_0_3_60/a_124_375# 0.008393f
C527 _17_/I FILLER_0_14_37/a_4516_472# 0.015502f
C528 _11_/I FILLER_0_4_37/a_3172_472# 0.014431f
C529 vdd input4/a_36_113# 0.121449f
C530 vdd FILLER_0_5_104/a_36_472# 0.093124f
C531 FILLER_0_14_37/a_932_472# FILLER_0_13_2/a_4964_472# 0.026657f
C532 input_signal[6] vdd 0.096151f
C533 FILLER_0_1_12/a_124_375# _10_/I 0.008103f
C534 FILLER_0_15_72/a_1380_472# _18_/I 0.014431f
C535 _10_/I FILLER_0_0_12/a_1020_375# 0.015932f
C536 input1/a_36_113# FILLER_0_0_12/a_124_375# 0.002124f
C537 FILLER_0_4_37/a_4516_472# FILLER_0_5_72/a_572_375# 0.001723f
C538 FILLER_0_15_8/a_1020_375# vdd 0.019054f
C539 _14_/I _04_/ZN 0.059451f
C540 _14_/I FILLER_0_7_2/a_2364_375# 0.008393f
C541 FILLER_0_8_107/a_572_375# _14_/I 0.011425f
C542 FILLER_0_11_72/a_124_375# FILLER_0_11_66/a_124_375# 0.005439f
C543 output14/a_224_472# output_signal_minus[8] 0.005065f
C544 FILLER_0_4_101/a_124_375# FILLER_0_5_72/a_3260_375# 0.026339f
C545 _10_/Z net15 0.00699f
C546 _11_/Z _09_/ZN 0.466752f
C547 FILLER_0_1_12/a_3260_375# FILLER_0_1_44/a_124_375# 0.012552f
C548 FILLER_0_6_37/a_4068_472# vdd 0.002856f
C549 output25/a_224_472# _08_/ZN 0.097677f
C550 FILLER_0_1_12/a_124_375# FILLER_0_0_12/a_124_375# 0.05841f
C551 _11_/I FILLER_0_3_12/a_1468_375# 0.008393f
C552 FILLER_0_6_2/a_1020_375# _12_/I 0.017312f
C553 FILLER_0_6_2/a_2812_375# _14_/I 0.003099f
C554 FILLER_0_13_2/a_6756_472# FILLER_0_14_37/a_2724_472# 0.026657f
C555 _16_/I FILLER_0_10_37/a_572_375# 0.002327f
C556 output24/a_224_472# output_signal_plus[1] 0.004499f
C557 _11_/I FILLER_0_3_60/a_484_472# 0.008683f
C558 FILLER_0_6_2/a_1916_375# _12_/I 0.016383f
C559 _08_/ZN output28/a_224_472# 0.005132f
C560 FILLER_0_1_72/a_484_472# FILLER_0_2_37/a_4516_472# 0.026657f
C561 _11_/I FILLER_0_2_107/a_124_375# 0.00346f
C562 FILLER_0_6_37/a_3172_472# _14_/I 0.001219f
C563 _11_/I FILLER_0_3_44/a_124_375# 0.008393f
C564 FILLER_0_7_72/a_2364_375# FILLER_0_5_72/a_2276_472# 0.001512f
C565 FILLER_0_13_2/a_1380_472# FILLER_0_12_12/a_124_375# 0.001684f
C566 vdd FILLER_0_11_72/a_5412_472# 0.005202f
C567 _11_/I FILLER_0_3_72/a_3172_472# 0.008683f
C568 _15_/I _16_/I 0.580399f
C569 output27/a_224_472# output_signal_plus[0] 0.00179f
C570 FILLER_0_14_37/a_1020_375# FILLER_0_13_2/a_4964_472# 0.001597f
C571 FILLER_0_2_2/a_2812_375# _10_/I 0.001886f
C572 FILLER_0_16_36/a_2364_375# _19_/I 0.015268f
C573 FILLER_0_13_2/a_6308_472# vdd 0.028986f
C574 FILLER_0_0_36/a_1020_375# _10_/I 0.015932f
C575 _17_/a_36_113# _16_/Z 0.018643f
C576 _11_/I FILLER_0_2_107/a_36_472# 0.002415f
C577 FILLER_0_1_60/a_124_375# _10_/I 0.008103f
C578 FILLER_0_6_2/a_2364_375# vdd -0.007525f
C579 output_signal_plus[7] _18_/a_36_113# 0.008247f
C580 FILLER_0_11_2/a_124_375# FILLER_0_9_2/a_36_472# 0.00108f
C581 FILLER_0_0_28/a_124_375# _10_/I 0.015932f
C582 output18/a_224_472# output_signal_minus[0] 0.007272f
C583 _07_/ZN output23/a_224_472# 0.065632f
C584 FILLER_0_0_142/a_124_375# output_signal_minus[7] 0.004157f
C585 FILLER_0_12_37/a_5500_375# FILLER_0_14_37/a_5412_472# 0.001512f
C586 FILLER_0_3_12/a_3260_375# FILLER_0_3_44/a_36_472# 0.086905f
C587 FILLER_0_6_37/a_4068_472# FILLER_0_4_37/a_4156_375# 0.001512f
C588 FILLER_0_5_104/a_484_472# output_signal_minus[4] 0.002187f
C589 vdd FILLER_0_3_44/a_932_472# 0.009767f
C590 _17_/I output29/a_224_472# 0.036533f
C591 _14_/I FILLER_0_9_72/a_2812_375# 0.004386f
C592 FILLER_0_2_2/a_3172_472# _10_/I 0.002566f
C593 FILLER_0_7_72/a_3172_472# _12_/I 0.004669f
C594 output23/a_224_472# _11_/a_36_113# 0.021122f
C595 output_signal_minus[5] output_signal_minus[6] 0.357719f
C596 FILLER_0_3_72/a_124_375# FILLER_0_2_37/a_4156_375# 0.026339f
C597 FILLER_0_2_2/a_1020_375# FILLER_0_4_2/a_932_472# 0.0027f
C598 FILLER_0_2_101/a_36_472# FILLER_0_2_37/a_6844_375# 0.086635f
C599 _15_/I FILLER_0_10_12/a_572_375# 0.018846f
C600 FILLER_0_13_72/a_36_472# _16_/I 0.004669f
C601 output21/a_224_472# output_signal_plus[0] 0.027735f
C602 FILLER_0_13_2/a_4068_472# vdd 0.003435f
C603 vdd FILLER_0_11_2/a_6844_375# 0.011466f
C604 _11_/I FILLER_0_4_107/a_1020_375# 0.014156f
C605 vdd FILLER_0_6_37/a_3260_375# 0.007161f
C606 FILLER_0_12_101/a_36_472# _15_/I 0.001368f
C607 FILLER_0_1_12/a_3260_375# FILLER_0_0_36/a_572_375# 0.05841f
C608 FILLER_0_9_2/a_6756_472# FILLER_0_11_2/a_6844_375# 0.001512f
C609 FILLER_0_15_8/a_2724_472# vdd 0.007608f
C610 FILLER_0_13_72/a_2276_472# vdd 0.012304f
C611 _16_/I FILLER_0_11_2/a_5500_375# 0.007169f
C612 FILLER_0_11_2/a_4604_375# vdd 0.007327f
C613 FILLER_0_8_37/a_4068_472# FILLER_0_7_72/a_36_472# 0.026657f
C614 FILLER_0_10_37/a_1916_375# FILLER_0_11_2/a_5860_472# 0.001723f
C615 _10_/I FILLER_0_1_12/a_932_472# 0.0057f
C616 FILLER_0_6_37/a_6396_375# _14_/I 0.001418f
C617 _11_/I FILLER_0_2_37/a_2724_472# 0.002415f
C618 FILLER_0_6_2/a_572_375# _12_/I 0.024441f
C619 FILLER_0_6_37/a_6308_472# FILLER_0_5_72/a_2364_375# 0.001597f
C620 FILLER_0_7_72/a_572_375# FILLER_0_8_37/a_4516_472# 0.001597f
C621 FILLER_0_10_107/a_36_472# _15_/I 0.016097f
C622 _02_/ZN output_signal_minus[4] 0.004102f
C623 input_signal[5] FILLER_0_11_2/a_124_375# 0.034101f
C624 _10_/Z output_signal_minus[4] 0.300374f
C625 FILLER_0_13_72/a_1916_375# _16_/I 0.006182f
C626 output_signal_plus[4] FILLER_0_11_72/a_6308_472# 0.001069f
C627 FILLER_0_6_37/a_4068_472# FILLER_0_5_72/a_36_472# 0.026657f
C628 FILLER_0_13_72/a_1468_375# FILLER_0_11_72/a_1380_472# 0.001512f
C629 _12_/a_36_113# _06_/ZN 0.012603f
C630 output_signal_plus[8] output21/a_224_472# 0.036402f
C631 FILLER_0_11_2/a_3260_375# vdd 0.020842f
C632 FILLER_0_9_2/a_4516_472# FILLER_0_10_37/a_572_375# 0.001597f
C633 _12_/I FILLER_0_7_72/a_932_472# 0.004669f
C634 output25/a_224_472# vdd 0.081784f
C635 FILLER_0_14_28/a_124_375# FILLER_0_14_37/a_124_375# 0.003228f
C636 FILLER_0_10_12/a_1468_375# FILLER_0_10_28/a_124_375# 0.012001f
C637 FILLER_0_7_2/a_4156_375# _14_/I 0.00647f
C638 FILLER_0_16_104/a_36_472# _19_/I 0.016117f
C639 FILLER_0_7_2/a_6308_472# FILLER_0_9_2/a_6396_375# 0.001512f
C640 _16_/I FILLER_0_10_37/a_1468_375# 0.002327f
C641 FILLER_0_9_2/a_1916_375# FILLER_0_7_2/a_1828_472# 0.0027f
C642 _11_/I FILLER_0_3_72/a_1468_375# 0.008393f
C643 _12_/Z _06_/ZN 0.003398f
C644 FILLER_0_11_72/a_1916_375# FILLER_0_10_37/a_5860_472# 0.001723f
C645 vdd output_signal_plus[9] 0.181616f
C646 FILLER_0_9_2/a_4516_472# _15_/I 0.006506f
C647 output12/a_224_472# _13_/I 0.038811f
C648 vdd output28/a_224_472# 0.110606f
C649 FILLER_0_11_72/a_124_375# FILLER_0_10_37/a_4068_472# 0.001723f
C650 FILLER_0_10_12/a_484_472# FILLER_0_11_2/a_1468_375# 0.001684f
C651 FILLER_0_5_104/a_572_375# FILLER_0_4_107/a_124_375# 0.026339f
C652 FILLER_0_15_40/a_932_472# _17_/I 0.004125f
C653 FILLER_0_14_12/a_1380_472# vdd 0.010304f
C654 _15_/I FILLER_0_12_37/a_4516_472# 0.001245f
C655 output15/a_224_472# net15 0.036927f
C656 FILLER_0_8_12/a_36_472# input5/a_36_113# 0.001663f
C657 FILLER_0_12_37/a_1380_472# vdd 0.006949f
C658 _00_/ZN FILLER_0_0_142/a_484_472# 0.015062f
C659 FILLER_0_2_2/a_2724_472# _10_/I 0.002545f
C660 _13_/I FILLER_0_4_37/a_2364_375# 0.003204f
C661 _08_/ZN _15_/Z 0.077979f
C662 FILLER_0_13_104/a_36_472# vdd 0.094649f
C663 FILLER_0_7_2/a_1828_472# FILLER_0_8_12/a_572_375# 0.001543f
C664 output21/a_224_472# FILLER_0_14_107/a_572_375# 0.001234f
C665 _11_/I FILLER_0_2_37/a_5052_375# 0.00346f
C666 FILLER_0_3_72/a_1020_375# FILLER_0_2_37/a_5052_375# 0.026339f
C667 _15_/I FILLER_0_9_72/a_1020_375# 0.006125f
C668 _12_/a_36_113# output_signal_minus[3] 0.024933f
C669 FILLER_0_2_107/a_572_375# vdd 0.015888f
C670 _11_/I FILLER_0_3_72/a_124_375# 0.008393f
C671 FILLER_0_8_12/a_932_472# FILLER_0_7_2/a_1916_375# 0.001543f
C672 output11/a_224_472# _01_/ZN 0.003295f
C673 _09_/ZN FILLER_0_11_72/a_5412_472# 0.037136f
C674 _18_/I FILLER_0_16_104/a_36_472# 0.004186f
C675 _12_/Z output_signal_minus[3] 0.061138f
C676 FILLER_0_0_142/a_36_472# output_signal_minus[7] 0.002068f
C677 FILLER_0_5_12/a_1020_375# vdd 0.026014f
C678 FILLER_0_14_12/a_1020_375# vdd -0.007174f
C679 FILLER_0_2_101/a_36_472# _10_/I 0.002486f
C680 FILLER_0_3_72/a_36_472# FILLER_0_5_72/a_124_375# 0.001512f
C681 FILLER_0_7_2/a_4068_472# _12_/I 0.004669f
C682 output_signal_plus[0] output_signal_plus[6] 0.001007f
C683 _13_/I FILLER_0_4_37/a_4516_472# 0.003497f
C684 FILLER_0_5_44/a_1468_375# FILLER_0_6_37/a_2276_472# 0.001597f
C685 output_signal_minus[1] output23/a_224_472# 0.023062f
C686 FILLER_0_13_2/a_2812_375# FILLER_0_12_28/a_36_472# 0.001684f
C687 FILLER_0_2_37/a_1468_375# vdd 0.010794f
C688 FILLER_0_1_12/a_1380_472# _10_/I 0.006408f
C689 _15_/I FILLER_0_10_28/a_124_375# 0.021137f
C690 _01_/ZN output_signal_minus[8] 0.068703f
C691 FILLER_0_1_60/a_572_375# FILLER_0_1_72/a_36_472# 0.009654f
C692 FILLER_0_4_2/a_36_472# input_signal[3] 0.007536f
C693 _12_/I FILLER_0_6_2/a_1468_375# 0.016629f
C694 FILLER_0_9_72/a_1828_472# FILLER_0_10_37/a_5860_472# 0.026657f
C695 output_signal_minus[7] FILLER_0_0_104/a_36_472# 0.002187f
C696 input3/a_36_113# FILLER_0_3_12/a_124_375# 0.002124f
C697 _11_/I FILLER_0_5_72/a_2364_375# 0.00439f
C698 _14_/I FILLER_0_7_72/a_3260_375# 0.00911f
C699 _07_/ZN output18/a_224_472# 0.002857f
C700 FILLER_0_11_2/a_1828_472# _16_/I 0.007596f
C701 FILLER_0_10_37/a_124_375# FILLER_0_11_2/a_4156_375# 0.026339f
C702 FILLER_0_9_72/a_36_472# FILLER_0_9_66/a_124_375# 0.016748f
C703 FILLER_0_13_104/a_484_472# vdd 0.008043f
C704 FILLER_0_1_60/a_484_472# _10_/I 0.006408f
C705 FILLER_0_13_2/a_6308_472# FILLER_0_14_37/a_2276_472# 0.026657f
C706 _07_/ZN _15_/I 0.172972f
C707 _11_/Z FILLER_0_11_72/a_5052_375# 0.001366f
C708 output24/a_224_472# output_signal_plus[2] 0.046354f
C709 FILLER_0_13_66/a_124_375# _17_/I 0.006125f
C710 FILLER_0_13_72/a_572_375# FILLER_0_14_37/a_4516_472# 0.001597f
C711 vdd FILLER_0_7_72/a_484_472# 0.002467f
C712 output_signal_plus[8] FILLER_0_14_37/a_6396_375# 0.001633f
C713 input_signal[6] input_signal[5] 0.00646f
C714 FILLER_0_3_72/a_572_375# vdd 0.002455f
C715 FILLER_0_14_107/a_124_375# _18_/I 0.003997f
C716 FILLER_0_14_28/a_36_472# _17_/I 0.015502f
C717 input_signal[0] vdd 0.033193f
C718 FILLER_0_5_12/a_3172_472# FILLER_0_5_44/a_36_472# 0.013276f
C719 FILLER_0_14_37/a_3172_472# _16_/I 0.001667f
C720 FILLER_0_2_37/a_932_472# vdd 0.007211f
C721 input_signal[3] input4/a_36_113# 0.059344f
C722 input8/a_36_113# FILLER_0_14_12/a_124_375# 0.002124f
C723 _12_/I FILLER_0_7_66/a_36_472# 0.004669f
C724 vdd FILLER_0_7_104/a_572_375# 0.011639f
C725 _15_/I _11_/a_36_113# 0.001741f
C726 FILLER_0_14_12/a_1380_472# FILLER_0_13_2/a_2364_375# 0.001543f
C727 _11_/I FILLER_0_3_12/a_1916_375# 0.008393f
C728 FILLER_0_11_2/a_3708_375# FILLER_0_9_2/a_3620_472# 0.0027f
C729 vdd FILLER_0_7_72/a_2364_375# 0.022764f
C730 _11_/I FILLER_0_1_12/a_36_472# 0.011335f
C731 vdd FILLER_0_3_104/a_36_472# 0.093924f
C732 input_signal[7] FILLER_0_14_12/a_36_472# 0.073591f
C733 output_signal_minus[6] _06_/ZN 0.060667f
C734 FILLER_0_14_101/a_36_472# FILLER_0_14_107/a_36_472# 0.003468f
C735 _14_/I FILLER_0_8_37/a_2724_472# 0.014431f
C736 FILLER_0_4_2/a_2364_375# _13_/I 0.00577f
C737 _14_/I FILLER_0_9_2/a_4604_375# 0.005381f
C738 _16_/I FILLER_0_10_107/a_1468_375# 0.002311f
C739 _10_/a_36_160# output_signal_minus[6] 0.006519f
C740 _15_/I FILLER_0_11_2/a_2276_472# 0.005458f
C741 _08_/ZN output_signal_plus[1] 0.070201f
C742 FILLER_0_2_107/a_1468_375# _01_/ZN 0.005666f
C743 _15_/I FILLER_0_9_2/a_1916_375# 0.006125f
C744 FILLER_0_8_37/a_3708_375# _14_/I 0.01418f
C745 output19/a_224_472# net15 0.024146f
C746 FILLER_0_11_2/a_4068_472# FILLER_0_12_37/a_36_472# 0.026657f
C747 FILLER_0_1_72/a_484_472# _10_/I 0.006408f
C748 FILLER_0_11_72/a_572_375# FILLER_0_9_72/a_484_472# 0.001512f
C749 FILLER_0_9_72/a_124_375# FILLER_0_9_66/a_124_375# 0.005439f
C750 FILLER_0_11_2/a_1828_472# FILLER_0_10_12/a_572_375# 0.001684f
C751 FILLER_0_7_2/a_1468_375# _14_/I 0.008393f
C752 FILLER_0_9_66/a_36_472# FILLER_0_9_2/a_6844_375# 0.086635f
C753 _12_/I output_signal_minus[4] 0.003502f
C754 output21/a_224_472# _19_/Z 0.099292f
C755 FILLER_0_14_107/a_484_472# FILLER_0_14_115/a_36_472# 0.013276f
C756 FILLER_0_2_37/a_4964_472# output20/a_224_472# 0.001058f
C757 FILLER_0_7_2/a_4068_472# FILLER_0_8_37/a_124_375# 0.001597f
C758 FILLER_0_14_37/a_5500_375# _18_/I 0.003988f
C759 _17_/I FILLER_0_12_37/a_2364_375# 0.001237f
C760 output15/a_224_472# output_signal_minus[4] 0.025424f
C761 output25/a_224_472# _09_/ZN 0.008059f
C762 _11_/I FILLER_0_2_2/a_932_472# 0.01353f
C763 FILLER_0_3_72/a_3260_375# FILLER_0_3_104/a_36_472# 0.086742f
C764 FILLER_0_11_72/a_2276_472# FILLER_0_13_72/a_2364_375# 0.001512f
C765 _16_/I FILLER_0_12_37/a_572_375# 0.016091f
C766 _15_/I FILLER_0_8_12/a_572_375# 0.001106f
C767 vdd _15_/Z 0.260202f
C768 _16_/I FILLER_0_10_37/a_3260_375# 0.002327f
C769 _15_/I FILLER_0_10_107/a_1380_472# 0.015502f
C770 output_signal_minus[7] _08_/ZN 0.055873f
C771 _11_/I FILLER_0_3_12/a_1020_375# 0.008561f
C772 _11_/I FILLER_0_3_12/a_1380_472# 0.008733f
C773 _09_/ZN output28/a_224_472# 0.076073f
C774 vdd FILLER_0_13_2/a_5500_375# 0.011603f
C775 vdd FILLER_0_16_36/a_1020_375# 0.003818f
C776 FILLER_0_6_2/a_932_472# vdd 0.00868f
C777 FILLER_0_3_72/a_2812_375# output11/a_224_472# 0.001216f
C778 vdd FILLER_0_12_107/a_1020_375# 0.001984f
C779 output18/a_224_472# FILLER_0_2_107/a_484_472# 0.001058f
C780 FILLER_0_13_66/a_124_375# FILLER_0_12_37/a_3260_375# 0.026339f
C781 FILLER_0_2_37/a_6308_472# output11/a_224_472# 0.031813f
C782 FILLER_0_14_37/a_6756_472# _18_/I 0.001153f
C783 _15_/I FILLER_0_10_37/a_36_472# 0.01654f
C784 FILLER_0_0_36/a_1020_375# FILLER_0_1_44/a_124_375# 0.05841f
C785 FILLER_0_6_37/a_5500_375# vdd 0.009137f
C786 FILLER_0_14_37/a_932_472# vdd 0.006024f
C787 FILLER_0_5_12/a_2724_472# FILLER_0_6_37/a_36_472# 0.026657f
C788 FILLER_0_2_37/a_484_472# _10_/I 0.002525f
C789 vdd FILLER_0_9_72/a_3260_375# 0.010174f
C790 FILLER_0_11_2/a_6756_472# vdd 0.008994f
C791 FILLER_0_3_12/a_3260_375# FILLER_0_1_12/a_3172_472# 0.001512f
C792 vdd FILLER_0_6_37/a_4156_375# 0.004039f
C793 FILLER_0_7_72/a_1468_375# _12_/I 0.006182f
C794 _17_/I FILLER_0_15_8/a_1468_375# 0.006523f
C795 FILLER_0_10_37/a_4156_375# vdd 0.004039f
C796 FILLER_0_10_28/a_36_472# FILLER_0_8_28/a_124_375# 0.0027f
C797 FILLER_0_3_60/a_572_375# vdd 0.028687f
C798 FILLER_0_10_101/a_36_472# FILLER_0_9_72/a_3172_472# 0.026657f
C799 _11_/I FILLER_0_2_37/a_4604_375# 0.003196f
C800 FILLER_0_9_2/a_6396_375# vdd 0.014009f
C801 _19_/I _16_/Z 0.002019f
C802 input_signal[0] input2/a_36_113# 0.001293f
C803 FILLER_0_16_36/a_3172_472# _19_/I 0.020111f
C804 FILLER_0_6_37/a_2812_375# FILLER_0_8_37/a_2724_472# 0.001512f
C805 FILLER_0_13_2/a_5052_375# vdd 0.009047f
C806 _13_/I FILLER_0_4_2/a_932_472# 0.00186f
C807 _17_/I FILLER_0_13_2/a_484_472# 0.001747f
C808 _11_/I FILLER_0_5_72/a_1380_472# 0.001913f
C809 FILLER_0_11_72/a_1916_375# FILLER_0_9_72/a_1828_472# 0.001512f
C810 output_signal_minus[1] _15_/I 0.0418f
C811 FILLER_0_9_72/a_572_375# FILLER_0_7_72/a_484_472# 0.001512f
C812 _09_/ZN FILLER_0_13_104/a_484_472# 0.001886f
C813 vdd FILLER_0_9_2/a_1380_472# 0.012473f
C814 FILLER_0_14_37/a_1020_375# vdd 0.008411f
C815 _07_/ZN _13_/I 0.033539f
C816 FILLER_0_6_37/a_5052_375# vdd 0.007396f
C817 FILLER_0_0_12/a_572_375# FILLER_0_1_12/a_572_375# 0.05841f
C818 FILLER_0_16_36/a_2724_472# FILLER_0_15_56/a_484_472# 0.05841f
C819 _14_/I FILLER_0_8_37/a_4604_375# 0.01418f
C820 vdd FILLER_0_1_60/a_36_472# 0.094979f
C821 input_signal[6] FILLER_0_11_2/a_484_472# 0.009925f
C822 FILLER_0_11_72/a_124_375# _15_/I 0.007126f
C823 _15_/I FILLER_0_9_2/a_6844_375# 0.006125f
C824 _18_/I FILLER_0_14_12/a_36_472# 0.001469f
C825 output19/a_224_472# output_signal_minus[4] 0.002161f
C826 vdd output_signal_plus[1] 0.249902f
C827 FILLER_0_5_44/a_572_375# _11_/I 0.004712f
C828 FILLER_0_7_2/a_3172_472# vdd 0.007993f
C829 FILLER_0_8_107/a_484_472# _11_/a_36_113# 0.001212f
C830 FILLER_0_5_104/a_484_472# _12_/I 0.003818f
C831 _17_/I FILLER_0_14_37/a_36_472# 0.01654f
C832 output15/a_224_472# FILLER_0_5_104/a_484_472# 0.003196f
C833 output30/a_224_472# output_signal_plus[9] 0.027875f
C834 _18_/I _16_/Z 0.056478f
C835 FILLER_0_16_36/a_3172_472# _18_/I 0.004109f
C836 _09_/ZN FILLER_0_3_104/a_36_472# 0.001203f
C837 vdd FILLER_0_10_37/a_5948_375# 0.010867f
C838 _01_/ZN _10_/I 0.198927f
C839 FILLER_0_11_2/a_2364_375# _15_/I 0.007165f
C840 FILLER_0_0_36/a_2812_375# _10_/I 0.015932f
C841 _11_/I FILLER_0_5_44/a_36_472# 0.001913f
C842 FILLER_0_10_37/a_1916_375# vdd 0.01389f
C843 FILLER_0_9_2/a_1828_472# vdd 0.046365f
C844 FILLER_0_6_37/a_1468_375# _14_/I 0.003099f
C845 FILLER_0_5_72/a_484_472# FILLER_0_6_37/a_4516_472# 0.026657f
C846 _15_/I FILLER_0_9_72/a_2364_375# 0.006125f
C847 FILLER_0_16_36/a_1468_375# _19_/I 0.014393f
C848 output_signal_minus[7] vdd 0.53571f
C849 FILLER_0_3_72/a_2812_375# FILLER_0_2_37/a_6844_375# 0.026339f
C850 FILLER_0_13_2/a_4604_375# vdd 0.007327f
C851 FILLER_0_10_28/a_36_472# FILLER_0_11_2/a_2812_375# 0.001684f
C852 FILLER_0_10_28/a_124_375# FILLER_0_9_2/a_3172_472# 0.001543f
C853 FILLER_0_4_37/a_6756_472# FILLER_0_3_72/a_2724_472# 0.026657f
C854 _00_/ZN output_signal_minus[4] 0.040929f
C855 FILLER_0_14_101/a_124_375# output29/a_224_472# 0.029497f
C856 FILLER_0_4_37/a_1380_472# FILLER_0_2_37/a_1468_375# 0.001512f
C857 _13_/I FILLER_0_4_37/a_4068_472# 0.003497f
C858 _13_/I FILLER_0_5_72/a_484_472# 0.017477f
C859 input_signal[6] input_signal[7] 0.005521f
C860 FILLER_0_12_107/a_1468_375# output_signal_plus[7] 0.001633f
C861 FILLER_0_10_12/a_572_375# _16_/I 0.001124f
C862 FILLER_0_5_12/a_1020_375# input_signal[3] 0.001277f
C863 _17_/I FILLER_0_15_8/a_36_472# 0.005458f
C864 output22/a_224_472# _11_/Z 0.08038f
C865 FILLER_0_2_2/a_2812_375# FILLER_0_3_12/a_1828_472# 0.001684f
C866 FILLER_0_3_44/a_1020_375# FILLER_0_1_44/a_932_472# 0.001512f
C867 FILLER_0_4_2/a_484_472# vdd 0.006484f
C868 FILLER_0_5_72/a_2812_375# vdd 0.019423f
C869 FILLER_0_15_8/a_1380_472# vdd 0.018348f
C870 FILLER_0_5_72/a_3172_472# _12_/I 0.003805f
C871 _16_/I FILLER_0_13_72/a_2812_375# 0.005045f
C872 FILLER_0_1_72/a_36_472# _10_/I 0.006408f
C873 FILLER_0_7_2/a_6396_375# _12_/I 0.006193f
C874 FILLER_0_11_66/a_36_472# FILLER_0_12_37/a_3172_472# 0.026657f
C875 _15_/I FILLER_0_11_2/a_1916_375# 0.002702f
C876 output13/a_224_472# output_signal_plus[1] 0.001201f
C877 FILLER_0_8_37/a_5052_375# vdd 0.007304f
C878 input_signal[0] input_signal[1] 0.099155f
C879 _02_/ZN _12_/I 0.032964f
C880 _10_/Z _12_/I 0.032848f
C881 FILLER_0_6_37/a_2724_472# vdd 0.00885f
C882 _09_/ZN FILLER_0_12_107/a_1020_375# 0.009573f
C883 FILLER_0_12_101/a_36_472# _16_/I 0.017723f
C884 FILLER_0_7_2/a_5860_472# FILLER_0_9_2/a_5948_375# 0.001512f
C885 output15/a_224_472# _10_/Z 0.079849f
C886 FILLER_0_11_2/a_3172_472# vdd 0.007993f
C887 vdd FILLER_0_5_72/a_1828_472# 0.00716f
C888 vdd FILLER_0_7_2/a_3708_375# 0.019534f
C889 FILLER_0_6_37/a_6308_472# FILLER_0_5_72/a_2276_472# 0.026657f
C890 _08_/ZN output_signal_plus[2] 0.319854f
C891 _14_/I FILLER_0_6_37/a_484_472# 0.001219f
C892 _15_/I FILLER_0_11_2/a_1020_375# 0.007214f
C893 _14_/I FILLER_0_7_2/a_1916_375# 0.008393f
C894 FILLER_0_11_66/a_36_472# FILLER_0_11_72/a_36_472# 0.003468f
C895 FILLER_0_4_37/a_4604_375# vdd 0.004103f
C896 FILLER_0_13_104/a_572_375# FILLER_0_12_107/a_124_375# 0.026339f
C897 _13_/I FILLER_0_4_2/a_2724_472# 0.003497f
C898 FILLER_0_8_12/a_484_472# vdd 0.024606f
C899 output_signal_plus[0] _18_/Z 0.043315f
C900 _18_/a_36_113# _16_/Z 0.0047f
C901 FILLER_0_12_37/a_6396_375# vdd 0.038787f
C902 FILLER_0_6_37/a_4068_472# FILLER_0_5_72/a_124_375# 0.001597f
C903 FILLER_0_11_66/a_36_472# vdd 0.097097f
C904 FILLER_0_8_12/a_1468_375# FILLER_0_10_12/a_1380_472# 0.0027f
C905 FILLER_0_4_2/a_2812_375# vdd 0.022312f
C906 FILLER_0_5_12/a_572_375# FILLER_0_6_2/a_1828_472# 0.001543f
C907 FILLER_0_6_37/a_36_472# FILLER_0_6_2/a_3260_375# 0.012267f
C908 output17/a_224_472# output_signal_minus[7] 0.055621f
C909 _16_/I FILLER_0_12_37/a_4516_472# 0.017477f
C910 FILLER_0_12_37/a_124_375# FILLER_0_12_28/a_124_375# 0.003228f
C911 FILLER_0_8_12/a_124_375# _15_/I 0.002388f
C912 _11_/I FILLER_0_2_107/a_1380_472# 0.002075f
C913 FILLER_0_11_72/a_3708_375# vdd 0.023316f
C914 vdd FILLER_0_14_37/a_6844_375# 0.010412f
C915 _13_/I FILLER_0_5_72/a_932_472# 0.017477f
C916 output_signal_minus[1] _13_/I 0.036295f
C917 _16_/Z _16_/a_36_113# 0.004105f
C918 input6/a_36_113# FILLER_0_10_12/a_124_375# 0.002124f
C919 FILLER_0_14_37/a_5860_472# vdd 0.008907f
C920 input3/a_36_113# _12_/I 0.005228f
C921 _12_/I FILLER_0_7_2/a_5052_375# 0.006193f
C922 _17_/a_36_113# _15_/Z 0.021431f
C923 _14_/I output14/a_224_472# 0.120448f
C924 FILLER_0_1_12/a_1828_472# FILLER_0_3_12/a_1916_375# 0.0027f
C925 vdd FILLER_0_7_2/a_2812_375# -0.009557f
C926 output_signal_plus[7] FILLER_0_13_104/a_572_375# 0.011852f
C927 FILLER_0_10_107/a_124_375# FILLER_0_9_104/a_484_472# 0.001597f
C928 FILLER_0_8_37/a_3620_472# vdd 0.007892f
C929 output_signal_minus[5] net15 0.023926f
C930 output_signal_plus[8] _18_/Z 0.030779f
C931 _17_/I FILLER_0_12_37/a_6844_375# 0.002388f
C932 FILLER_0_15_56/a_484_472# vdd 0.007111f
C933 _17_/I FILLER_0_14_107/a_36_472# 0.016097f
C934 FILLER_0_2_37/a_6308_472# _10_/I 0.001464f
C935 FILLER_0_8_107/a_572_375# _15_/I 0.002302f
C936 FILLER_0_13_72/a_2276_472# FILLER_0_14_37/a_6308_472# 0.026657f
C937 _09_/ZN output_signal_plus[1] 0.020081f
C938 FILLER_0_2_2/a_2276_472# FILLER_0_3_12/a_1020_375# 0.001684f
C939 _07_/ZN output12/a_224_472# 0.062608f
C940 FILLER_0_16_18/a_124_375# input_signal[9] 0.007441f
C941 output_signal_plus[4] _10_/Z 0.095553f
C942 FILLER_0_6_37/a_3708_375# FILLER_0_8_37/a_3620_472# 0.0027f
C943 input_signal[6] FILLER_0_12_12/a_36_472# 0.073761f
C944 _11_/Z FILLER_0_9_104/a_572_375# 0.018997f
C945 vdd FILLER_0_3_12/a_3172_472# 0.002817f
C946 FILLER_0_11_72/a_1468_375# vdd 0.007205f
C947 _16_/I FILLER_0_10_28/a_124_375# 0.002327f
C948 FILLER_0_14_107/a_484_472# _17_/I 0.015502f
C949 _11_/I FILLER_0_5_72/a_2276_472# 0.001913f
C950 FILLER_0_7_2/a_124_375# input_signal[4] 0.028776f
C951 vdd FILLER_0_8_37/a_4156_375# 0.004039f
C952 FILLER_0_12_107/a_36_472# FILLER_0_10_107/a_124_375# 0.001512f
C953 FILLER_0_4_37/a_1828_472# FILLER_0_3_44/a_1020_375# 0.001597f
C954 FILLER_0_14_107/a_572_375# _18_/Z 0.0276f
C955 FILLER_0_11_72/a_1828_472# vdd 0.008296f
C956 output19/a_224_472# _10_/Z 0.041987f
C957 _15_/I FILLER_0_11_72/a_3172_472# 0.005458f
C958 _12_/Z _14_/a_36_113# 0.057599f
C959 FILLER_0_9_72/a_3172_472# _14_/I 0.004017f
C960 FILLER_0_15_72/a_1468_375# output29/a_224_472# 0.023259f
C961 _07_/ZN _16_/I 0.11878f
C962 FILLER_0_1_72/a_1020_375# _10_/I 0.008103f
C963 FILLER_0_2_2/a_1828_472# vdd 0.048778f
C964 vdd FILLER_0_5_60/a_572_375# 0.028544f
C965 vdd FILLER_0_2_37/a_3620_472# 0.008985f
C966 _18_/I FILLER_0_15_8/a_1020_375# 0.014659f
C967 FILLER_0_14_37/a_1468_375# vdd 0.010281f
C968 vdd FILLER_0_4_2/a_1828_472# 0.044032f
C969 _17_/I FILLER_0_14_37/a_572_375# 0.018729f
C970 output_signal_plus[2] vdd 0.272722f
C971 FILLER_0_16_104/a_124_375# vdd 0.026929f
C972 FILLER_0_13_72/a_2364_375# vdd 0.022764f
C973 FILLER_0_13_104/a_36_472# FILLER_0_13_72/a_3172_472# 0.013277f
C974 FILLER_0_9_2/a_932_472# vdd 0.009688f
C975 FILLER_0_5_12/a_3172_472# vdd 0.003484f
C976 input_signal[5] FILLER_0_9_2/a_1380_472# 0.002679f
C977 output15/a_224_472# _12_/I 0.0161f
C978 _15_/I FILLER_0_9_72/a_2812_375# 0.006125f
C979 FILLER_0_11_2/a_2276_472# _16_/I 0.007596f
C980 FILLER_0_5_104/a_484_472# FILLER_0_4_107/a_124_375# 0.001723f
C981 _00_/ZN _02_/ZN 0.166903f
C982 _00_/ZN _10_/Z 0.002152f
C983 vdd FILLER_0_16_18/a_1020_375# 0.004841f
C984 FILLER_0_10_12/a_1020_375# vdd 0.024939f
C985 FILLER_0_2_107/a_572_375# output_signal_minus[8] 0.003512f
C986 vdd FILLER_0_16_36/a_1828_472# 0.006448f
C987 output_signal_plus[5] _16_/I 0.022659f
C988 FILLER_0_11_2/a_4964_472# FILLER_0_12_37/a_1020_375# 0.001597f
C989 FILLER_0_7_2/a_4604_375# _12_/I 0.006193f
C990 FILLER_0_5_12/a_484_472# FILLER_0_6_2/a_1468_375# 0.001543f
C991 FILLER_0_11_72/a_4604_375# FILLER_0_10_107/a_572_375# 0.026339f
C992 _14_/I FILLER_0_6_37/a_572_375# 0.003099f
C993 FILLER_0_8_37/a_1828_472# _14_/I 0.014431f
C994 FILLER_0_15_8/a_36_472# FILLER_0_15_2/a_36_472# 0.003468f
C995 _15_/I FILLER_0_12_37/a_3620_472# 0.001368f
C996 FILLER_0_3_72/a_572_375# FILLER_0_2_37/a_4516_472# 0.001723f
C997 FILLER_0_6_101/a_36_472# FILLER_0_7_72/a_3260_375# 0.001723f
C998 FILLER_0_15_8/a_2364_375# _17_/I 0.006523f
C999 _19_/I FILLER_0_15_8/a_2724_472# 0.001938f
C1000 _16_/I FILLER_0_14_37/a_1380_472# 0.001667f
C1001 output_signal_minus[5] output_signal_minus[4] 0.115171f
C1002 _11_/I _08_/ZN 0.033163f
C1003 input_signal[5] FILLER_0_9_2/a_1828_472# 0.001351f
C1004 FILLER_0_14_12/a_932_472# vdd 0.017846f
C1005 FILLER_0_11_72/a_6844_375# FILLER_0_11_136/a_124_375# 0.012001f
C1006 FILLER_0_15_8/a_3260_375# FILLER_0_15_40/a_36_472# 0.086904f
C1007 FILLER_0_3_44/a_572_375# FILLER_0_1_44/a_484_472# 0.001512f
C1008 output_signal_plus[2] output13/a_224_472# 0.005065f
C1009 FILLER_0_10_101/a_36_472# FILLER_0_10_37/a_6756_472# 0.013277f
C1010 FILLER_0_5_44/a_1020_375# FILLER_0_3_44/a_932_472# 0.001512f
C1011 FILLER_0_8_12/a_124_375# input5/a_36_113# 0.002124f
C1012 _17_/I _10_/Z 0.043791f
C1013 FILLER_0_13_2/a_1380_472# vdd 0.013839f
C1014 output24/a_224_472# _12_/Z 0.005705f
C1015 _13_/I FILLER_0_5_60/a_484_472# 0.017924f
C1016 FILLER_0_12_12/a_932_472# _15_/I 0.001368f
C1017 _13_/I FILLER_0_4_37/a_6756_472# 0.002988f
C1018 FILLER_0_6_2/a_2276_472# _14_/I 0.001219f
C1019 _19_/Z _18_/Z 0.013331f
C1020 _15_/I FILLER_0_10_37/a_6396_375# 0.018729f
C1021 FILLER_0_0_70/a_124_375# vdd 0.042733f
C1022 input9/a_36_113# input_signal[8] 0.070332f
C1023 _13_/I FILLER_0_4_37/a_36_472# 0.003497f
C1024 _11_/I FILLER_0_4_37/a_5500_375# 0.01418f
C1025 _19_/I output_signal_plus[9] 0.130261f
C1026 _15_/I FILLER_0_11_72/a_1020_375# 0.007126f
C1027 _14_/I FILLER_0_9_2/a_5860_472# 0.003526f
C1028 FILLER_0_6_37/a_6308_472# vdd 0.019175f
C1029 output_signal_minus[1] output12/a_224_472# 0.015047f
C1030 FILLER_0_3_44/a_124_375# FILLER_0_1_44/a_36_472# 0.001512f
C1031 vdd FILLER_0_2_37/a_4156_375# 0.004039f
C1032 _13_/I _04_/ZN 0.364663f
C1033 FILLER_0_10_37/a_5052_375# FILLER_0_12_37/a_4964_472# 0.001512f
C1034 FILLER_0_8_37/a_5948_375# _14_/I 0.01418f
C1035 _18_/I FILLER_0_15_8/a_2724_472# 0.014431f
C1036 _17_/I FILLER_0_15_72/a_572_375# 0.006589f
C1037 _11_/I FILLER_0_5_12/a_1468_375# 0.004745f
C1038 _17_/I FILLER_0_12_37/a_2812_375# 0.002388f
C1039 FILLER_0_12_37/a_5412_472# FILLER_0_10_37/a_5500_375# 0.001512f
C1040 FILLER_0_10_101/a_124_375# FILLER_0_11_72/a_3260_375# 0.026339f
C1041 output_signal_minus[2] output_signal_plus[1] 0.002823f
C1042 FILLER_0_5_72/a_36_472# FILLER_0_5_60/a_572_375# 0.009654f
C1043 output23/a_224_472# _15_/a_36_113# 0.002892f
C1044 output14/a_224_472# output16/a_224_472# 0.005712f
C1045 _12_/I FILLER_0_5_12/a_1380_472# 0.003872f
C1046 FILLER_0_12_37/a_36_472# _16_/I 0.019816f
C1047 FILLER_0_1_44/a_1020_375# FILLER_0_2_37/a_1828_472# 0.001597f
C1048 FILLER_0_4_2/a_484_472# input_signal[3] 0.003397f
C1049 vdd FILLER_0_8_37/a_6396_375# 0.038694f
C1050 FILLER_0_6_2/a_2812_375# _13_/I 0.001706f
C1051 output_signal_plus[7] output_signal_plus[8] 0.171782f
C1052 vdd input_signal[8] 0.141473f
C1053 FILLER_0_3_72/a_1916_375# FILLER_0_2_37/a_5948_375# 0.026339f
C1054 FILLER_0_6_37/a_3172_472# _13_/I 0.003818f
C1055 FILLER_0_15_64/a_36_472# FILLER_0_16_36/a_3172_472# 0.05841f
C1056 vdd FILLER_0_4_37/a_1020_375# 0.008282f
C1057 FILLER_0_11_72/a_4068_472# FILLER_0_12_107/a_124_375# 0.001597f
C1058 FILLER_0_4_37/a_3620_472# _11_/I 0.014431f
C1059 output15/a_224_472# output19/a_224_472# 0.005204f
C1060 _14_/I _01_/ZN 0.003111f
C1061 input_signal[2] FILLER_0_2_2/a_1020_375# 0.001016f
C1062 _13_/I FILLER_0_4_37/a_5412_472# 0.003497f
C1063 _18_/I output_signal_plus[9] 0.016401f
C1064 _18_/I output28/a_224_472# 0.037282f
C1065 FILLER_0_11_72/a_124_375# _16_/I 0.007169f
C1066 _18_/I FILLER_0_14_12/a_1380_472# 0.001526f
C1067 _17_/I FILLER_0_14_115/a_36_472# 0.015502f
C1068 FILLER_0_15_8/a_3260_375# FILLER_0_14_37/a_124_375# 0.026339f
C1069 vdd FILLER_0_5_12/a_2276_472# 0.008296f
C1070 FILLER_0_13_72/a_1468_375# vdd 0.007205f
C1071 FILLER_0_3_72/a_1380_472# vdd 0.006325f
C1072 FILLER_0_14_101/a_36_472# _17_/I 0.015502f
C1073 FILLER_0_15_72/a_1380_472# output_signal_plus[8] 0.002792f
C1074 _17_/I FILLER_0_15_72/a_124_375# 0.006589f
C1075 output_signal_minus[3] net15 0.110724f
C1076 _14_/I FILLER_0_7_72/a_1380_472# 0.008683f
C1077 FILLER_0_11_72/a_3260_375# vdd 0.00923f
C1078 FILLER_0_4_107/a_1468_375# output_signal_minus[4] 0.002255f
C1079 FILLER_0_5_12/a_1916_375# vdd 0.021506f
C1080 _03_/ZN output_signal_minus[4] 0.001191f
C1081 _17_/Z _08_/ZN 0.007125f
C1082 output24/a_224_472# FILLER_0_11_136/a_124_375# 0.032639f
C1083 FILLER_0_9_72/a_484_472# FILLER_0_10_37/a_4516_472# 0.026657f
C1084 FILLER_0_8_12/a_124_375# FILLER_0_7_2/a_1380_472# 0.001543f
C1085 vdd FILLER_0_11_2/a_2724_472# 0.009793f
C1086 _17_/I FILLER_0_14_37/a_5948_375# 0.018729f
C1087 FILLER_0_11_2/a_2364_375# _16_/I 0.007169f
C1088 FILLER_0_7_72/a_1916_375# _12_/I 0.006182f
C1089 _13_/I FILLER_0_5_104/a_124_375# 0.017198f
C1090 _11_/I FILLER_0_5_12/a_124_375# 0.004745f
C1091 FILLER_0_14_12/a_1020_375# _18_/I 0.003935f
C1092 FILLER_0_13_2/a_6844_375# _16_/I 0.006193f
C1093 FILLER_0_11_2/a_5948_375# FILLER_0_9_2/a_5860_472# 0.001512f
C1094 FILLER_0_6_37/a_1020_375# FILLER_0_7_2/a_4964_472# 0.001723f
C1095 _11_/I vdd 2.106998f
C1096 FILLER_0_3_72/a_1020_375# vdd 0.00558f
C1097 vdd FILLER_0_7_72/a_2276_472# 0.011667f
C1098 FILLER_0_12_37/a_4964_472# FILLER_0_11_72/a_932_472# 0.026657f
C1099 FILLER_0_6_37/a_4068_472# FILLER_0_7_72/a_124_375# 0.001723f
C1100 FILLER_0_6_107/a_36_472# _14_/I 0.001219f
C1101 FILLER_0_8_37/a_1468_375# FILLER_0_9_2/a_5500_375# 0.026339f
C1102 _15_/I FILLER_0_9_2/a_4604_375# 0.006125f
C1103 _14_/I FILLER_0_8_101/a_36_472# 0.015237f
C1104 _16_/I FILLER_0_11_2/a_1916_375# 0.007169f
C1105 _13_/I FILLER_0_6_37/a_6396_375# 0.001706f
C1106 FILLER_0_8_37/a_3708_375# _15_/I 0.002388f
C1107 FILLER_0_13_72/a_3260_375# _16_/I 0.006182f
C1108 FILLER_0_5_12/a_1828_472# vdd 0.009457f
C1109 _11_/I FILLER_0_3_12/a_2276_472# 0.008787f
C1110 FILLER_0_9_2/a_572_375# input_signal[4] 0.005834f
C1111 _11_/I FILLER_0_3_72/a_3260_375# 0.008393f
C1112 _14_/I FILLER_0_8_107/a_36_472# 0.017114f
C1113 FILLER_0_3_60/a_572_375# FILLER_0_2_37/a_3260_375# 0.026339f
C1114 _17_/I FILLER_0_13_72/a_1380_472# 0.00652f
C1115 FILLER_0_4_37/a_6844_375# FILLER_0_4_101/a_36_472# 0.086635f
C1116 _11_/Z _14_/I 0.002864f
C1117 _06_/ZN output_signal_minus[4] 0.037168f
C1118 _16_/I FILLER_0_11_2/a_1020_375# 0.007169f
C1119 FILLER_0_6_37/a_932_472# FILLER_0_5_44/a_36_472# 0.026657f
C1120 FILLER_0_7_2/a_3260_375# FILLER_0_6_2/a_3260_375# 0.05841f
C1121 FILLER_0_13_66/a_36_472# vdd 0.097796f
C1122 FILLER_0_12_12/a_1020_375# FILLER_0_14_12/a_932_472# 0.0027f
C1123 FILLER_0_7_2/a_5860_472# vdd 0.017109f
C1124 _19_/I _15_/Z 0.029195f
C1125 _14_/I FILLER_0_6_37/a_3620_472# 0.001219f
C1126 FILLER_0_8_37/a_1916_375# _14_/I 0.01418f
C1127 output_signal_minus[5] _10_/Z 0.075569f
C1128 FILLER_0_12_37/a_6756_472# vdd 0.014295f
C1129 _11_/I FILLER_0_4_37/a_4156_375# 0.01418f
C1130 FILLER_0_8_37/a_1468_375# FILLER_0_7_2/a_5412_472# 0.001597f
C1131 FILLER_0_10_28/a_124_375# FILLER_0_10_37/a_36_472# 0.007947f
C1132 vdd FILLER_0_9_2/a_2812_375# 0.022556f
C1133 FILLER_0_7_2/a_6756_472# FILLER_0_7_66/a_36_472# 0.013276f
C1134 _19_/I FILLER_0_16_36/a_1020_375# 0.01418f
C1135 _11_/I FILLER_0_2_37/a_5500_375# 0.00346f
C1136 _11_/I output13/a_224_472# 0.083231f
C1137 FILLER_0_11_72/a_2364_375# vdd 0.02275f
C1138 FILLER_0_8_37/a_6844_375# _14_/I 0.014366f
C1139 FILLER_0_2_107/a_1020_375# _01_/ZN 0.004676f
C1140 FILLER_0_10_12/a_932_472# FILLER_0_8_12/a_1020_375# 0.0027f
C1141 FILLER_0_2_37/a_1468_375# _10_/I 0.001886f
C1142 input_signal[5] FILLER_0_9_2/a_932_472# 0.011077f
C1143 output_signal_plus[7] _19_/Z 0.01101f
C1144 FILLER_0_10_37/a_6756_472# FILLER_0_11_72/a_2812_375# 0.001723f
C1145 FILLER_0_16_104/a_124_375# output30/a_224_472# 0.001073f
C1146 _00_/ZN output_signal_plus[4] 0.046436f
C1147 FILLER_0_11_72/a_2276_472# FILLER_0_12_37/a_6308_472# 0.026657f
C1148 _15_/I _15_/a_36_113# 0.022654f
C1149 FILLER_0_8_37/a_5052_375# FILLER_0_10_37/a_4964_472# 0.001512f
C1150 FILLER_0_5_44/a_1468_375# FILLER_0_4_37/a_2276_472# 0.001723f
C1151 output_signal_minus[3] output_signal_minus[4] 0.324744f
C1152 output_signal_minus[7] output_signal_minus[8] 0.515416f
C1153 FILLER_0_12_107/a_1380_472# vdd 0.007259f
C1154 FILLER_0_2_107/a_1380_472# output_signal_minus[6] 0.002051f
C1155 vdd FILLER_0_14_37/a_2724_472# 0.009656f
C1156 _08_/ZN FILLER_0_11_72/a_6756_472# 0.00637f
C1157 FILLER_0_12_101/a_36_472# FILLER_0_13_72/a_3260_375# 0.001723f
C1158 output27/a_224_472# output21/a_224_472# 0.219442f
C1159 FILLER_0_4_2/a_572_375# vdd 0.019843f
C1160 input_signal[0] _10_/I 0.207716f
C1161 _17_/Z vdd 0.377565f
C1162 vdd FILLER_0_8_37/a_4964_472# 0.005164f
C1163 input_signal[2] FILLER_0_3_12/a_36_472# 0.075115f
C1164 FILLER_0_8_37/a_5412_472# FILLER_0_7_72/a_1380_472# 0.026657f
C1165 FILLER_0_2_37/a_932_472# _10_/I 0.002525f
C1166 FILLER_0_8_37/a_1380_472# _14_/I 0.014431f
C1167 FILLER_0_15_40/a_1380_472# _17_/I 0.004125f
C1168 _12_/a_36_113# _08_/ZN 0.001302f
C1169 _14_/Z output_signal_plus[4] 0.056171f
C1170 FILLER_0_11_72/a_5948_375# _10_/Z 0.013107f
C1171 vdd FILLER_0_6_37/a_1916_375# 0.014924f
C1172 vdd FILLER_0_6_37/a_4604_375# 0.004123f
C1173 vdd FILLER_0_0_36/a_2724_472# 0.007577f
C1174 _15_/I FILLER_0_10_37/a_1380_472# 0.015502f
C1175 _11_/I input2/a_36_113# 0.004615f
C1176 _11_/I FILLER_0_5_72/a_36_472# 0.001913f
C1177 FILLER_0_16_104/a_36_472# output_signal_plus[0] 0.002187f
C1178 vdd FILLER_0_11_72/a_484_472# 0.002467f
C1179 input_signal[0] FILLER_0_0_12/a_124_375# 0.006465f
C1180 FILLER_0_4_2/a_1020_375# vdd 0.021954f
C1181 output_signal_minus[2] output_signal_plus[2] 0.002124f
C1182 FILLER_0_12_37/a_1468_375# _17_/I 0.002388f
C1183 _01_/ZN output16/a_224_472# 0.006402f
C1184 _17_/I output_signal_plus[4] 0.008117f
C1185 FILLER_0_2_107/a_572_375# FILLER_0_4_107/a_484_472# 0.0027f
C1186 FILLER_0_4_2/a_124_375# _12_/I 0.029788f
C1187 FILLER_0_11_72/a_1468_375# FILLER_0_9_72/a_1380_472# 0.001512f
C1188 FILLER_0_7_2/a_36_472# input_signal[4] 0.061272f
C1189 FILLER_0_14_101/a_124_375# FILLER_0_14_107/a_36_472# 0.016748f
C1190 _12_/Z _08_/ZN 0.069554f
C1191 _07_/ZN output_signal_minus[1] 0.097037f
C1192 FILLER_0_14_37/a_932_472# _18_/I 0.001526f
C1193 FILLER_0_12_12/a_1380_472# FILLER_0_12_28/a_36_472# 0.013276f
C1194 _16_/I FILLER_0_13_2/a_2724_472# 0.004669f
C1195 _15_/I FILLER_0_11_2/a_6396_375# 0.007111f
C1196 _13_/I FILLER_0_5_12/a_572_375# 0.016091f
C1197 FILLER_0_8_37/a_3260_375# FILLER_0_9_66/a_124_375# 0.026339f
C1198 FILLER_0_6_2/a_3172_472# _14_/I 0.001219f
C1199 _13_/I FILLER_0_4_2/a_1380_472# 0.003497f
C1200 FILLER_0_11_72/a_3172_472# _16_/I 0.00753f
C1201 _15_/I FILLER_0_8_37/a_4604_375# 0.002181f
C1202 input_signal[9] FILLER_0_15_2/a_36_472# 0.021082f
C1203 vdd FILLER_0_4_2/a_3260_375# 0.043008f
C1204 FILLER_0_12_37/a_6396_375# FILLER_0_14_37/a_6308_472# 0.001512f
C1205 FILLER_0_13_2/a_1020_375# FILLER_0_11_2/a_932_472# 0.0027f
C1206 FILLER_0_8_37/a_5860_472# FILLER_0_9_72/a_1916_375# 0.001723f
C1207 _11_/I FILLER_0_4_37/a_932_472# 0.014431f
C1208 FILLER_0_7_2/a_5412_472# _12_/I 0.004669f
C1209 FILLER_0_6_107/a_124_375# FILLER_0_8_107/a_36_472# 0.001512f
C1210 _11_/I _09_/ZN 0.963184f
C1211 _11_/I FILLER_0_5_12/a_2812_375# 0.004712f
C1212 FILLER_0_12_37/a_4156_375# _17_/I 0.002049f
C1213 FILLER_0_4_37/a_5052_375# FILLER_0_6_37/a_4964_472# 0.001512f
C1214 _13_/I FILLER_0_4_37/a_4964_472# 0.003497f
C1215 _16_/I FILLER_0_13_2/a_1468_375# 0.006236f
C1216 output_signal_plus[8] FILLER_0_16_104/a_36_472# 0.03558f
C1217 _14_/I FILLER_0_7_104/a_124_375# 0.010093f
C1218 _14_/I FILLER_0_9_72/a_1916_375# 0.005381f
C1219 FILLER_0_4_37/a_1828_472# FILLER_0_3_44/a_932_472# 0.026657f
C1220 _18_/I FILLER_0_14_37/a_1020_375# 0.003988f
C1221 FILLER_0_14_37/a_572_375# FILLER_0_13_2/a_4516_472# 0.001597f
C1222 FILLER_0_3_12/a_2276_472# FILLER_0_4_2/a_3260_375# 0.001543f
C1223 output_signal_plus[3] output_signal_plus[4] 0.138344f
C1224 FILLER_0_10_37/a_2812_375# FILLER_0_11_2/a_6844_375# 0.026339f
C1225 _00_/ZN _14_/Z 0.037483f
C1226 _11_/I FILLER_0_3_44/a_1468_375# 0.008393f
C1227 FILLER_0_7_72/a_1020_375# _12_/I 0.006182f
C1228 _12_/I _13_/a_36_113# 0.082448f
C1229 FILLER_0_6_37/a_4068_472# _14_/I 0.001209f
C1230 _00_/ZN _17_/I 0.406419f
C1231 output15/a_224_472# _13_/a_36_113# 0.013428f
C1232 output27/a_224_472# output_signal_plus[6] 0.05886f
C1233 FILLER_0_7_66/a_36_472# FILLER_0_8_37/a_3260_375# 0.001597f
C1234 FILLER_0_7_72/a_3172_472# FILLER_0_7_104/a_36_472# 0.013276f
C1235 FILLER_0_2_2/a_1916_375# vdd 0.051352f
C1236 _17_/I FILLER_0_12_12/a_572_375# 0.001106f
C1237 output22/a_224_472# output_signal_plus[1] 0.02182f
C1238 FILLER_0_3_44/a_1380_472# FILLER_0_5_44/a_1468_375# 0.001512f
C1239 FILLER_0_15_8/a_1380_472# _19_/I 0.00191f
C1240 _16_/I FILLER_0_12_37/a_3620_472# 0.017477f
C1241 FILLER_0_12_37/a_124_375# FILLER_0_13_2/a_4068_472# 0.001723f
C1242 _15_/Z _16_/a_36_113# 0.070659f
C1243 FILLER_0_8_107/a_124_375# FILLER_0_8_101/a_124_375# 0.005439f
C1244 FILLER_0_12_101/a_36_472# FILLER_0_11_72/a_3172_472# 0.026657f
C1245 _11_/I input_signal[1] 0.077808f
C1246 _08_/ZN FILLER_0_11_136/a_124_375# 0.047331f
C1247 output_signal_plus[5] output_signal_plus[6] 0.13932f
C1248 vdd FILLER_0_11_72/a_6756_472# 0.022349f
C1249 _15_/I FILLER_0_10_37/a_2724_472# 0.015502f
C1250 FILLER_0_3_104/a_572_375# _01_/ZN 0.001549f
C1251 _02_/ZN _06_/ZN 0.405943f
C1252 FILLER_0_9_104/a_484_472# vdd 0.00781f
C1253 _13_/I FILLER_0_5_72/a_1468_375# 0.016091f
C1254 _17_/I _14_/Z 0.026798f
C1255 FILLER_0_3_12/a_3260_375# FILLER_0_2_37/a_484_472# 0.001723f
C1256 _10_/a_36_160# _10_/Z 0.003981f
C1257 _08_/ZN output_signal_minus[6] 0.047598f
C1258 _16_/I FILLER_0_13_2/a_2812_375# 0.006236f
C1259 FILLER_0_4_37/a_1380_472# _11_/I 0.014431f
C1260 _12_/a_36_113# vdd 0.015445f
C1261 FILLER_0_12_12/a_932_472# _16_/I 0.017483f
C1262 _11_/I FILLER_0_4_107/a_932_472# 0.014431f
C1263 FILLER_0_2_2/a_2276_472# vdd 0.013919f
C1264 FILLER_0_6_2/a_2364_375# _14_/I 0.003099f
C1265 _09_/ZN FILLER_0_12_107/a_1380_472# 0.020589f
C1266 _17_/I FILLER_0_15_8/a_124_375# 0.007193f
C1267 FILLER_0_5_12/a_36_472# input4/a_36_113# 0.001663f
C1268 _08_/ZN output26/a_224_472# 0.003213f
C1269 _16_/I FILLER_0_10_37/a_6396_375# 0.001124f
C1270 FILLER_0_1_60/a_36_472# _10_/I 0.006408f
C1271 _16_/I FILLER_0_13_2/a_3708_375# 0.006313f
C1272 _11_/I FILLER_0_5_12/a_932_472# 0.001494f
C1273 FILLER_0_5_12/a_484_472# _12_/I 0.006214f
C1274 FILLER_0_1_12/a_1468_375# FILLER_0_0_12/a_1468_375# 0.05841f
C1275 _11_/I input_signal[3] 0.035429f
C1276 FILLER_0_15_8/a_1380_472# _18_/I 0.015237f
C1277 FILLER_0_13_72/a_2364_375# FILLER_0_14_37/a_6308_472# 0.001597f
C1278 FILLER_0_9_2/a_4068_472# FILLER_0_11_2/a_4156_375# 0.001512f
C1279 _12_/Z vdd 0.273556f
C1280 _00_/ZN output_signal_plus[3] 0.062658f
C1281 output21/a_224_472# output_signal_plus[6] 0.002816f
C1282 _16_/I FILLER_0_11_72/a_1020_375# 0.007169f
C1283 FILLER_0_4_107/a_1020_375# output_signal_minus[4] 0.001688f
C1284 FILLER_0_4_37/a_36_472# FILLER_0_3_12/a_2812_375# 0.001597f
C1285 FILLER_0_15_56/a_572_375# vdd 0.011129f
C1286 FILLER_0_12_107/a_36_472# vdd 0.110178f
C1287 FILLER_0_7_2/a_932_472# input_signal[4] 0.004151f
C1288 _02_/ZN output_signal_minus[3] 0.045286f
C1289 FILLER_0_15_56/a_36_472# FILLER_0_16_36/a_2276_472# 0.05841f
C1290 output_signal_minus[3] _10_/Z 0.06108f
C1291 FILLER_0_10_28/a_36_472# vdd 0.097913f
C1292 FILLER_0_2_2/a_1468_375# FILLER_0_3_12/a_484_472# 0.001684f
C1293 FILLER_0_1_12/a_1828_472# vdd 0.008796f
C1294 _15_/I input6/a_36_113# 0.008411f
C1295 FILLER_0_0_36/a_1828_472# vdd 0.006872f
C1296 vdd FILLER_0_16_36/a_2276_472# 0.038168f
C1297 vdd FILLER_0_0_36/a_1916_375# -0.006107f
C1298 _11_/I FILLER_0_2_37/a_1916_375# 0.003339f
C1299 output25/a_224_472# _13_/Z 0.003776f
C1300 FILLER_0_13_2/a_6756_472# FILLER_0_12_37/a_2812_375# 0.001723f
C1301 FILLER_0_5_60/a_572_375# FILLER_0_5_72/a_124_375# 0.003732f
C1302 output_signal_plus[3] _14_/Z 0.096524f
C1303 FILLER_0_8_37/a_6756_472# FILLER_0_7_72/a_2812_375# 0.001597f
C1304 FILLER_0_15_56/a_484_472# _19_/I 0.001782f
C1305 FILLER_0_13_2/a_1020_375# FILLER_0_14_12/a_36_472# 0.001543f
C1306 output_signal_minus[7] _10_/I 0.480451f
C1307 _15_/I FILLER_0_12_37/a_5412_472# 0.001368f
C1308 FILLER_0_9_72/a_932_472# vdd 0.004803f
C1309 _14_/I FILLER_0_6_37/a_3260_375# 0.003099f
C1310 FILLER_0_11_72/a_5860_472# output28/a_224_472# 0.002432f
C1311 FILLER_0_16_104/a_36_472# _19_/Z 0.019249f
C1312 _11_/I FILLER_0_4_101/a_124_375# 0.014212f
C1313 FILLER_0_10_101/a_36_472# FILLER_0_9_72/a_3260_375# 0.001597f
C1314 _11_/I output_signal_minus[2] 0.034821f
C1315 _11_/I FILLER_0_2_37/a_1020_375# 0.00346f
C1316 _03_/ZN _12_/I 0.032657f
C1317 FILLER_0_12_101/a_124_375# _16_/I 0.017203f
C1318 output15/a_224_472# FILLER_0_4_107/a_1468_375# 0.029497f
C1319 output15/a_224_472# _03_/ZN 0.005522f
C1320 _18_/I FILLER_0_14_37/a_6844_375# 0.003935f
C1321 output_signal_minus[5] output19/a_224_472# 0.052257f
C1322 FILLER_0_6_37/a_1468_375# _13_/I 0.001706f
C1323 FILLER_0_6_101/a_36_472# FILLER_0_5_72/a_3260_375# 0.001597f
C1324 FILLER_0_7_2/a_6844_375# vdd 0.011885f
C1325 FILLER_0_14_37/a_5860_472# _18_/I 0.001526f
C1326 FILLER_0_12_107/a_1468_375# FILLER_0_11_72/a_5412_472# 0.001597f
C1327 FILLER_0_1_72/a_1020_375# output20/a_224_472# 0.03228f
C1328 FILLER_0_8_107/a_572_375# _11_/a_36_113# 0.002037f
C1329 _12_/I FILLER_0_5_12/a_3260_375# 0.001706f
C1330 _17_/I FILLER_0_12_37/a_3260_375# 0.002388f
C1331 FILLER_0_7_2/a_4068_472# FILLER_0_9_2/a_4156_375# 0.001512f
C1332 FILLER_0_8_12/a_484_472# FILLER_0_9_2/a_1468_375# 0.001684f
C1333 FILLER_0_4_37/a_572_375# FILLER_0_5_12/a_3260_375# 0.026339f
C1334 _17_/a_36_113# _17_/Z 0.004248f
C1335 _15_/I FILLER_0_9_72/a_3172_472# 0.00652f
C1336 _15_/I FILLER_0_10_12/a_1380_472# 0.015502f
C1337 _18_/I FILLER_0_15_56/a_484_472# 0.014431f
C1338 FILLER_0_15_72/a_124_375# FILLER_0_14_37/a_4068_472# 0.001723f
C1339 FILLER_0_7_72/a_124_375# FILLER_0_6_37/a_4156_375# 0.026339f
C1340 FILLER_0_12_37/a_5860_472# vdd 0.007851f
C1341 FILLER_0_4_37/a_6396_375# FILLER_0_6_37/a_6308_472# 0.001512f
C1342 FILLER_0_6_2/a_484_472# FILLER_0_4_2/a_572_375# 0.0027f
C1343 FILLER_0_11_136/a_124_375# vdd 0.042415f
C1344 FILLER_0_10_107/a_124_375# FILLER_0_11_72/a_4156_375# 0.026339f
C1345 vdd FILLER_0_4_107/a_1380_472# 0.002196f
C1346 FILLER_0_10_37/a_5412_472# FILLER_0_8_37/a_5500_375# 0.001512f
C1347 FILLER_0_14_37/a_5412_472# _16_/I 0.001667f
C1348 input_signal[3] FILLER_0_4_2/a_572_375# 0.008479f
C1349 output28/a_224_472# FILLER_0_11_72/a_4964_472# 0.001463f
C1350 FILLER_0_16_104/a_124_375# _19_/I 0.009128f
C1351 output_signal_minus[6] vdd 0.31108f
C1352 FILLER_0_5_44/a_932_472# _12_/I 0.003805f
C1353 _13_/I FILLER_0_4_107/a_36_472# 0.003497f
C1354 vdd FILLER_0_7_2/a_1020_375# -0.008191f
C1355 _00_/ZN output_signal_minus[5] 0.043945f
C1356 _12_/I FILLER_0_5_72/a_1916_375# 0.001706f
C1357 FILLER_0_4_2/a_1916_375# _12_/I 0.001625f
C1358 FILLER_0_11_2/a_6308_472# FILLER_0_12_37/a_2276_472# 0.026657f
C1359 FILLER_0_6_37/a_36_472# _12_/I 0.019129f
C1360 vdd output26/a_224_472# 0.059563f
C1361 FILLER_0_15_8/a_1916_375# FILLER_0_16_18/a_932_472# 0.001543f
C1362 _09_/ZN FILLER_0_9_104/a_484_472# 0.001414f
C1363 _06_/ZN _12_/I 0.001685f
C1364 _19_/I FILLER_0_16_18/a_1020_375# 0.01418f
C1365 _13_/I FILLER_0_6_37/a_484_472# 0.003818f
C1366 input_signal[2] FILLER_0_3_12/a_572_375# 0.003342f
C1367 _19_/I FILLER_0_16_36/a_1828_472# 0.01568f
C1368 FILLER_0_2_37/a_932_472# FILLER_0_1_44/a_124_375# 0.001597f
C1369 FILLER_0_3_72/a_3172_472# FILLER_0_4_101/a_36_472# 0.026657f
C1370 FILLER_0_14_37/a_1468_375# _18_/I 0.003988f
C1371 _15_/I FILLER_0_11_2/a_932_472# 0.005458f
C1372 FILLER_0_9_66/a_36_472# FILLER_0_10_37/a_3172_472# 0.026657f
C1373 FILLER_0_1_12/a_2364_375# vdd 0.018969f
C1374 FILLER_0_13_2/a_3260_375# _17_/I 0.006125f
C1375 _11_/I FILLER_0_4_37/a_1468_375# 0.01418f
C1376 FILLER_0_3_72/a_2364_375# vdd 0.022764f
C1377 FILLER_0_16_70/a_36_472# FILLER_0_14_37/a_3708_375# 0.001436f
C1378 FILLER_0_7_2/a_4516_472# vdd 0.005419f
C1379 vdd FILLER_0_1_12/a_1468_375# -0.00845f
C1380 FILLER_0_12_37/a_6308_472# vdd 0.019363f
C1381 FILLER_0_8_37/a_1468_375# FILLER_0_9_2/a_5412_472# 0.001723f
C1382 _13_/I FILLER_0_4_37/a_5860_472# 0.003497f
C1383 FILLER_0_16_104/a_124_375# _18_/I 0.001989f
C1384 _11_/I FILLER_0_2_37/a_4516_472# 0.001106f
C1385 vdd FILLER_0_8_37/a_3172_472# 0.006745f
C1386 FILLER_0_1_12/a_1380_472# FILLER_0_2_2/a_2364_375# 0.001543f
C1387 _16_/I FILLER_0_12_107/a_124_375# 0.016256f
C1388 output22/a_224_472# output_signal_plus[2] 0.007987f
C1389 _11_/I FILLER_0_4_2/a_1468_375# 0.014453f
C1390 FILLER_0_6_37/a_1020_375# vdd 0.006813f
C1391 FILLER_0_12_107/a_36_472# _09_/ZN 0.001273f
C1392 FILLER_0_11_2/a_6756_472# FILLER_0_10_37/a_2812_375# 0.001723f
C1393 FILLER_0_6_37/a_932_472# vdd 0.005743f
C1394 FILLER_0_11_72/a_4604_375# vdd 0.00451f
C1395 vdd FILLER_0_3_12/a_2724_472# 0.002467f
C1396 FILLER_0_4_37/a_2812_375# FILLER_0_5_60/a_124_375# 0.026339f
C1397 _15_/I FILLER_0_11_72/a_2724_472# 0.00215f
C1398 output_signal_minus[3] _12_/I 0.048486f
C1399 _14_/I FILLER_0_7_72/a_484_472# 0.002089f
C1400 FILLER_0_12_107/a_1468_375# output25/a_224_472# 0.009488f
C1401 FILLER_0_7_2/a_6756_472# _12_/I 0.004669f
C1402 output15/a_224_472# output_signal_minus[3] 0.006135f
C1403 input6/a_36_113# input5/a_36_113# 0.001442f
C1404 _18_/I FILLER_0_16_36/a_1828_472# 0.001782f
C1405 FILLER_0_7_2/a_5412_472# FILLER_0_9_2/a_5500_375# 0.001512f
C1406 vdd FILLER_0_10_37/a_484_472# 0.004128f
C1407 FILLER_0_1_12/a_36_472# FILLER_0_3_12/a_124_375# 0.0027f
C1408 FILLER_0_9_72/a_2724_472# vdd 0.034112f
C1409 FILLER_0_2_2/a_1380_472# _11_/I 0.00653f
C1410 _13_/I output14/a_224_472# 0.057064f
C1411 vdd FILLER_0_14_37/a_4516_472# 0.002735f
C1412 FILLER_0_13_2/a_572_375# vdd 0.02016f
C1413 vdd FILLER_0_9_2/a_6308_472# 0.028286f
C1414 _11_/I FILLER_0_4_37/a_6396_375# 0.01418f
C1415 _13_/I FILLER_0_5_72/a_1020_375# 0.016091f
C1416 FILLER_0_6_107/a_36_472# FILLER_0_6_101/a_36_472# 0.003468f
C1417 _14_/I FILLER_0_7_104/a_572_375# 0.207187f
C1418 FILLER_0_14_115/a_124_375# output28/a_224_472# 0.001597f
C1419 FILLER_0_12_107/a_1468_375# output28/a_224_472# 0.029497f
C1420 FILLER_0_8_37/a_36_472# FILLER_0_7_2/a_4068_472# 0.026657f
C1421 input_signal[6] FILLER_0_11_2/a_36_472# 0.027333f
C1422 FILLER_0_4_37/a_1916_375# FILLER_0_6_37/a_1828_472# 0.001512f
C1423 output17/a_224_472# output_signal_minus[6] 0.022663f
C1424 FILLER_0_5_12/a_2724_472# vdd 0.003283f
C1425 _14_/I FILLER_0_7_72/a_2364_375# 0.008393f
C1426 _11_/I output_signal_minus[8] 0.0259f
C1427 FILLER_0_2_37/a_3620_472# _10_/I 0.002517f
C1428 FILLER_0_1_72/a_932_472# vdd 0.004803f
C1429 _11_/I FILLER_0_4_37/a_6308_472# 0.014431f
C1430 input10/a_36_113# input_signal[8] 0.042822f
C1431 _15_/I FILLER_0_9_2/a_5860_472# 0.006506f
C1432 _15_/I FILLER_0_8_37/a_5948_375# 0.002388f
C1433 FILLER_0_11_66/a_124_375# FILLER_0_11_2/a_6844_375# 0.012001f
C1434 FILLER_0_14_12/a_932_472# _18_/I 0.001153f
C1435 output_signal_plus[7] _16_/I 0.023741f
C1436 FILLER_0_13_2/a_5052_375# FILLER_0_11_2/a_4964_472# 0.001512f
C1437 _19_/I input_signal[8] 0.137832f
C1438 FILLER_0_11_72/a_572_375# vdd 0.002455f
C1439 _11_/I FILLER_0_2_37/a_3260_375# 0.00346f
C1440 FILLER_0_14_12/a_1020_375# FILLER_0_13_2/a_2276_472# 0.001543f
C1441 FILLER_0_13_2/a_932_472# _16_/I 0.004669f
C1442 FILLER_0_4_37/a_124_375# FILLER_0_6_37/a_36_472# 0.001512f
C1443 output18/a_224_472# _01_/ZN 0.044051f
C1444 FILLER_0_5_44/a_1380_472# _12_/I 0.003805f
C1445 _16_/I FILLER_0_11_2/a_6396_375# 0.007169f
C1446 _11_/I FILLER_0_5_72/a_124_375# 0.004712f
C1447 _17_/I FILLER_0_13_72/a_572_375# 0.003577f
C1448 FILLER_0_12_37/a_5948_375# FILLER_0_13_72/a_1916_375# 0.026339f
C1449 vdd FILLER_0_7_72/a_1828_472# 0.008296f
C1450 _15_/I FILLER_0_10_37/a_3172_472# 0.015502f
C1451 FILLER_0_6_2/a_932_472# _14_/I 0.001219f
C1452 output27/a_224_472# _18_/Z 0.04012f
C1453 _09_/ZN FILLER_0_4_107/a_1380_472# 0.082253f
C1454 FILLER_0_8_37/a_572_375# vdd 0.00526f
C1455 _11_/I FILLER_0_2_107/a_1468_375# 0.003258f
C1456 _18_/I input_signal[8] 0.041737f
C1457 FILLER_0_7_2/a_2364_375# FILLER_0_8_12/a_1380_472# 0.001543f
C1458 _19_/Z _16_/Z 0.001069f
C1459 FILLER_0_12_107/a_1020_375# FILLER_0_11_72/a_4964_472# 0.001597f
C1460 FILLER_0_6_37/a_5500_375# _14_/I 0.003099f
C1461 vdd output29/a_224_472# 0.100233f
C1462 FILLER_0_3_104/a_484_472# FILLER_0_4_107/a_36_472# 0.026657f
C1463 FILLER_0_13_104/a_572_375# output28/a_224_472# 0.011959f
C1464 FILLER_0_7_2/a_5948_375# vdd 0.032854f
C1465 FILLER_0_12_37/a_4156_375# FILLER_0_14_37/a_4068_472# 0.001512f
C1466 _14_/I FILLER_0_9_72/a_3260_375# 0.005381f
C1467 FILLER_0_4_2/a_2276_472# FILLER_0_2_2/a_2364_375# 0.0027f
C1468 FILLER_0_10_12/a_1468_375# FILLER_0_12_12/a_1380_472# 0.0027f
C1469 _14_/I FILLER_0_6_37/a_4156_375# 0.002629f
C1470 output19/a_224_472# output_signal_minus[3] 0.005065f
C1471 FILLER_0_7_72/a_572_375# vdd 0.002455f
C1472 FILLER_0_7_72/a_2812_375# _12_/I 0.005045f
C1473 vdd FILLER_0_0_12/a_932_472# 0.012458f
C1474 FILLER_0_2_2/a_572_375# input_signal[2] 0.010396f
C1475 _11_/I FILLER_0_4_37/a_2724_472# 0.014431f
C1476 FILLER_0_6_37/a_4964_472# _12_/I 0.017477f
C1477 _00_/ZN _06_/ZN 0.473117f
C1478 _17_/I FILLER_0_15_72/a_484_472# 0.004125f
C1479 _13_/Z output_signal_plus[1] 0.098465f
C1480 _11_/I FILLER_0_2_37/a_6844_375# 0.00346f
C1481 _13_/I FILLER_0_6_37/a_572_375# 0.001706f
C1482 _14_/I FILLER_0_9_2/a_6396_375# 0.005381f
C1483 FILLER_0_0_70/a_124_375# _10_/I 0.015932f
C1484 FILLER_0_15_72/a_1468_375# FILLER_0_13_72/a_1380_472# 0.001512f
C1485 FILLER_0_6_37/a_1380_472# FILLER_0_5_44/a_484_472# 0.026657f
C1486 _00_/ZN _10_/a_36_160# 0.006235f
C1487 FILLER_0_4_37/a_5860_472# FILLER_0_2_37/a_5948_375# 0.001512f
C1488 FILLER_0_14_107/a_484_472# FILLER_0_12_107/a_572_375# 0.0027f
C1489 FILLER_0_6_107/a_124_375# FILLER_0_7_104/a_572_375# 0.026339f
C1490 vdd FILLER_0_11_2/a_4156_375# 0.004039f
C1491 FILLER_0_10_12/a_1020_375# FILLER_0_9_2/a_2276_472# 0.001543f
C1492 FILLER_0_4_2/a_2276_472# _13_/I 0.003497f
C1493 output21/a_224_472# _18_/Z 0.102793f
C1494 vdd FILLER_0_13_2/a_124_375# 0.012902f
C1495 _14_/I FILLER_0_9_2/a_1380_472# 0.004017f
C1496 _12_/Z output_signal_minus[2] 0.047494f
C1497 FILLER_0_10_12/a_124_375# FILLER_0_9_2/a_1380_472# 0.001543f
C1498 FILLER_0_13_72/a_3260_375# FILLER_0_11_72/a_3172_472# 0.001512f
C1499 _14_/I FILLER_0_6_37/a_5052_375# 0.003099f
C1500 _13_/I FILLER_0_4_37/a_2812_375# 0.005726f
C1501 FILLER_0_15_8/a_572_375# _17_/I 0.006523f
C1502 FILLER_0_11_72/a_4604_375# _09_/ZN 0.004803f
C1503 FILLER_0_5_12/a_2812_375# FILLER_0_3_12/a_2724_472# 0.001512f
C1504 _13_/I FILLER_0_5_72/a_3260_375# 0.01659f
C1505 _14_/I output_signal_plus[1] 0.037728f
C1506 _13_/I FILLER_0_6_2/a_2276_472# 0.003872f
C1507 _15_/I _11_/Z 0.015538f
C1508 FILLER_0_7_2/a_3172_472# _14_/I 0.008787f
C1509 _00_/ZN output_signal_minus[3] 0.044218f
C1510 FILLER_0_5_12/a_572_375# FILLER_0_3_12/a_484_472# 0.0027f
C1511 FILLER_0_7_72/a_1468_375# FILLER_0_5_72/a_1380_472# 0.001512f
C1512 FILLER_0_5_104/a_572_375# vdd 0.020942f
C1513 _15_/I FILLER_0_12_12/a_1380_472# 0.001368f
C1514 _11_/I FILLER_0_2_2/a_36_472# 0.010829f
C1515 _15_/I FILLER_0_8_37/a_1916_375# 0.002367f
C1516 _11_/I output22/a_224_472# 0.016465f
C1517 _11_/I FILLER_0_5_44/a_1020_375# 0.004712f
C1518 output15/a_224_472# FILLER_0_4_107/a_1020_375# 0.029497f
C1519 FILLER_0_11_72/a_572_375# FILLER_0_10_37/a_4604_375# 0.026339f
C1520 FILLER_0_5_44/a_1468_375# FILLER_0_5_60/a_124_375# 0.012222f
C1521 FILLER_0_1_72/a_124_375# FILLER_0_2_37/a_4068_472# 0.001597f
C1522 FILLER_0_11_136/a_36_472# _16_/I 0.009708f
C1523 output12/a_224_472# output14/a_224_472# 0.005408f
C1524 FILLER_0_15_40/a_932_472# vdd 0.004364f
C1525 FILLER_0_8_37/a_6844_375# _15_/I 0.002388f
C1526 _17_/I FILLER_0_13_2/a_4516_472# 0.006506f
C1527 FILLER_0_13_2/a_6756_472# _17_/I 0.006506f
C1528 FILLER_0_14_101/a_124_375# _17_/I 0.019472f
C1529 _17_/I FILLER_0_14_37/a_4068_472# 0.015502f
C1530 FILLER_0_12_37/a_1468_375# FILLER_0_13_2/a_5412_472# 0.001723f
C1531 vdd FILLER_0_6_2/a_3260_375# 0.010972f
C1532 FILLER_0_11_2/a_5412_472# FILLER_0_12_37/a_1468_375# 0.001597f
C1533 FILLER_0_1_12/a_1020_375# FILLER_0_2_2/a_2276_472# 0.001543f
C1534 FILLER_0_10_107/a_1020_375# vdd 0.002455f
C1535 FILLER_0_16_36/a_36_472# FILLER_0_16_18/a_1380_472# 0.003468f
C1536 FILLER_0_6_37/a_3172_472# FILLER_0_5_60/a_484_472# 0.026657f
C1537 FILLER_0_7_2/a_484_472# input_signal[4] 0.008159f
C1538 FILLER_0_11_72/a_5500_375# vdd 0.007282f
C1539 output_signal_minus[9] output_signal_minus[7] 0.005128f
C1540 FILLER_0_1_72/a_1380_472# FILLER_0_3_72/a_1468_375# 0.001512f
C1541 FILLER_0_4_37/a_3260_375# vdd 0.008639f
C1542 _11_/I FILLER_0_4_37/a_5948_375# 0.01418f
C1543 _17_/Z _19_/I 0.006359f
C1544 _15_/I FILLER_0_10_37/a_6756_472# 0.015502f
C1545 FILLER_0_8_37/a_5052_375# _14_/I 0.01418f
C1546 FILLER_0_8_37/a_124_375# FILLER_0_8_28/a_124_375# 0.003228f
C1547 FILLER_0_11_72/a_6844_375# _10_/Z 0.008557f
C1548 _11_/I _10_/I 0.007761f
C1549 FILLER_0_6_37/a_2724_472# _14_/I 0.001219f
C1550 FILLER_0_12_37/a_5412_472# _16_/I 0.017477f
C1551 _11_/I FILLER_0_5_12/a_2364_375# 0.004781f
C1552 _02_/ZN _14_/a_36_113# 0.020254f
C1553 vdd FILLER_0_1_44/a_36_472# 0.089951f
C1554 output_signal_plus[6] _18_/Z 0.011292f
C1555 _14_/I FILLER_0_7_2/a_3708_375# 0.006303f
C1556 FILLER_0_6_37/a_5500_375# FILLER_0_8_37/a_5412_472# 0.001512f
C1557 FILLER_0_15_64/a_36_472# FILLER_0_15_56/a_484_472# 0.013277f
C1558 FILLER_0_12_12/a_932_472# FILLER_0_11_2/a_1916_375# 0.001543f
C1559 vdd FILLER_0_0_142/a_484_472# 0.007827f
C1560 FILLER_0_2_101/a_36_472# output_signal_minus[0] 0.002109f
C1561 output_signal_plus[0] output_signal_plus[9] 0.433936f
C1562 FILLER_0_9_2/a_124_375# input_signal[4] 0.035733f
C1563 FILLER_0_6_2/a_1020_375# vdd -0.008425f
C1564 FILLER_0_8_12/a_484_472# _14_/I 0.014741f
C1565 input_signal[2] FILLER_0_3_12/a_484_472# 0.001534f
C1566 _03_/ZN _13_/a_36_113# 0.002627f
C1567 output_signal_plus[7] output27/a_224_472# 0.065176f
C1568 _18_/I FILLER_0_14_37/a_2724_472# 0.001526f
C1569 FILLER_0_9_72/a_2276_472# vdd 0.011667f
C1570 FILLER_0_13_66/a_124_375# vdd 0.042248f
C1571 FILLER_0_6_2/a_1916_375# vdd 0.017057f
C1572 vdd FILLER_0_10_37/a_5412_472# 0.006901f
C1573 _15_/I FILLER_0_10_37/a_2364_375# 0.018729f
C1574 _08_/ZN net15 0.722542f
C1575 _17_/Z _18_/I 0.24858f
C1576 _17_/I FILLER_0_12_37/a_1916_375# 0.002367f
C1577 FILLER_0_14_28/a_36_472# vdd 0.097913f
C1578 FILLER_0_12_12/a_1468_375# _17_/I 0.002388f
C1579 FILLER_0_5_60/a_36_472# FILLER_0_5_44/a_1468_375# 0.086742f
C1580 vdd FILLER_0_9_2/a_2364_375# 0.024816f
C1581 FILLER_0_11_2/a_5948_375# FILLER_0_10_37/a_1916_375# 0.026339f
C1582 FILLER_0_7_2/a_3260_375# _12_/I 0.006134f
C1583 output_signal_plus[5] output_signal_plus[7] 0.01783f
C1584 vdd FILLER_0_11_72/a_6308_472# 0.005474f
C1585 FILLER_0_6_107/a_36_472# _13_/I 0.011739f
C1586 output_signal_plus[8] output_signal_plus[9] 0.551989f
C1587 _12_/I FILLER_0_5_72/a_2364_375# 0.001706f
C1588 _17_/I FILLER_0_15_8/a_2812_375# 0.006723f
C1589 _17_/I FILLER_0_15_40/a_1468_375# 0.006589f
C1590 _16_/I FILLER_0_12_28/a_124_375# 0.018215f
C1591 FILLER_0_13_2/a_1380_472# FILLER_0_14_12/a_124_375# 0.001543f
C1592 FILLER_0_9_72/a_932_472# FILLER_0_10_37/a_4964_472# 0.026657f
C1593 _15_/I FILLER_0_9_72/a_1916_375# 0.006125f
C1594 vdd input_signal[4] 0.128179f
C1595 FILLER_0_6_37/a_6756_472# FILLER_0_5_72/a_2812_375# 0.001597f
C1596 vdd FILLER_0_0_36/a_1380_472# 0.004747f
C1597 _14_/I FILLER_0_7_2/a_2812_375# 0.008393f
C1598 FILLER_0_15_8/a_3260_375# FILLER_0_15_40/a_124_375# 0.012552f
C1599 _13_/I FILLER_0_5_44/a_484_472# 0.017477f
C1600 FILLER_0_8_37/a_3620_472# _14_/I 0.014431f
C1601 _11_/I FILLER_0_3_72/a_2276_472# 0.008683f
C1602 FILLER_0_10_101/a_36_472# FILLER_0_11_72/a_3260_375# 0.001723f
C1603 input_signal[6] _15_/I 0.030463f
C1604 FILLER_0_12_107/a_932_472# vdd 0.002467f
C1605 vdd FILLER_0_12_37/a_2364_375# 0.027535f
C1606 _11_/I FILLER_0_4_107/a_484_472# 0.014431f
C1607 FILLER_0_9_72/a_1468_375# FILLER_0_10_37/a_5412_472# 0.001597f
C1608 FILLER_0_7_104/a_36_472# _12_/I 0.004669f
C1609 FILLER_0_12_101/a_124_375# FILLER_0_13_72/a_3260_375# 0.026339f
C1610 FILLER_0_8_107/a_484_472# _11_/Z 0.001795f
C1611 output_signal_plus[7] output21/a_224_472# 0.00756f
C1612 FILLER_0_6_37/a_1828_472# _12_/I 0.017477f
C1613 FILLER_0_7_72/a_3172_472# vdd 0.009151f
C1614 _17_/I FILLER_0_13_2/a_5412_472# 0.006506f
C1615 _16_/I FILLER_0_11_2/a_932_472# 0.005931f
C1616 _13_/I FILLER_0_6_37/a_3620_472# 0.003965f
C1617 FILLER_0_5_104/a_572_375# _09_/ZN 0.003262f
C1618 FILLER_0_12_12/a_124_375# input7/a_36_113# 0.002124f
C1619 FILLER_0_5_44/a_1468_375# _13_/I 0.016091f
C1620 FILLER_0_0_142/a_124_375# _10_/Z 0.003267f
C1621 _13_/Z output_signal_plus[2] 0.021201f
C1622 output24/a_224_472# _10_/Z 0.053005f
C1623 FILLER_0_15_72/a_1468_375# _17_/I 0.006589f
C1624 FILLER_0_13_72/a_1468_375# FILLER_0_12_37/a_5500_375# 0.026339f
C1625 _14_/I FILLER_0_8_37/a_4156_375# 0.01418f
C1626 output_signal_minus[5] _06_/ZN 0.051053f
C1627 FILLER_0_12_37/a_5948_375# _16_/I 0.016091f
C1628 FILLER_0_8_37/a_484_472# vdd 0.003786f
C1629 FILLER_0_2_2/a_1468_375# FILLER_0_4_2/a_1380_472# 0.0027f
C1630 _15_/I FILLER_0_11_72/a_5412_472# 0.004676f
C1631 FILLER_0_10_12/a_484_472# vdd 0.023895f
C1632 FILLER_0_0_36/a_2724_472# _10_/I 0.016187f
C1633 FILLER_0_4_2/a_2812_375# FILLER_0_6_2/a_2724_472# 0.0027f
C1634 output30/a_224_472# output29/a_224_472# 0.072646f
C1635 FILLER_0_10_107/a_1020_375# _09_/ZN 0.009573f
C1636 FILLER_0_11_72/a_2724_472# _16_/I 0.00753f
C1637 FILLER_0_4_2/a_2812_375# FILLER_0_3_12/a_1828_472# 0.001543f
C1638 FILLER_0_2_2/a_2812_375# FILLER_0_4_2/a_2724_472# 0.0027f
C1639 FILLER_0_6_2/a_572_375# vdd -0.010507f
C1640 _09_/ZN FILLER_0_11_72/a_5500_375# 0.048757f
C1641 _17_/Z _18_/a_36_113# 0.001822f
C1642 _14_/I output_signal_plus[2] 0.028537f
C1643 output11/a_224_472# output_signal_minus[6] 0.010207f
C1644 FILLER_0_10_37/a_6308_472# FILLER_0_8_37/a_6396_375# 0.001512f
C1645 output_signal_minus[7] output16/a_224_472# 0.003702f
C1646 _07_/ZN FILLER_0_11_136/a_36_472# 0.013793f
C1647 vdd FILLER_0_7_72/a_932_472# 0.004803f
C1648 vdd FILLER_0_15_8/a_1468_375# -0.006196f
C1649 _16_/I FILLER_0_13_72/a_2724_472# 0.00187f
C1650 FILLER_0_9_2/a_932_472# _14_/I 0.002651f
C1651 _17_/Z _16_/a_36_113# 0.007498f
C1652 FILLER_0_15_40/a_484_472# FILLER_0_16_36/a_932_472# 0.05841f
C1653 FILLER_0_4_2/a_1916_375# FILLER_0_3_12/a_932_472# 0.001543f
C1654 _08_/ZN output_signal_minus[4] 0.036684f
C1655 _11_/Z FILLER_0_10_107/a_1468_375# 0.003499f
C1656 output_signal_minus[6] output_signal_minus[8] 0.165904f
C1657 FILLER_0_13_2/a_4068_472# FILLER_0_14_37/a_124_375# 0.001597f
C1658 FILLER_0_7_2/a_2276_472# FILLER_0_9_2/a_2364_375# 0.0027f
C1659 FILLER_0_1_72/a_1468_375# vdd 0.014833f
C1660 vdd net15 0.264485f
C1661 FILLER_0_11_2/a_1828_472# FILLER_0_13_2/a_1916_375# 0.0027f
C1662 FILLER_0_3_12/a_1916_375# FILLER_0_4_2/a_3172_472# 0.001543f
C1663 _19_/I FILLER_0_16_36/a_2276_472# 0.016804f
C1664 FILLER_0_13_2/a_484_472# vdd 0.009126f
C1665 FILLER_0_14_37/a_6756_472# _16_/I 0.001653f
C1666 output11/a_224_472# FILLER_0_3_72/a_2364_375# 0.001216f
C1667 output22/a_224_472# FILLER_0_9_104/a_484_472# 0.002002f
C1668 FILLER_0_8_37/a_124_375# FILLER_0_9_2/a_4156_375# 0.026339f
C1669 FILLER_0_7_2/a_2724_472# FILLER_0_9_2/a_2812_375# 0.0027f
C1670 FILLER_0_2_37/a_2276_472# FILLER_0_1_44/a_1468_375# 0.001597f
C1671 FILLER_0_7_2/a_932_472# _12_/I 0.004669f
C1672 _13_/I FILLER_0_6_2/a_3172_472# 0.003872f
C1673 FILLER_0_13_2/a_572_375# FILLER_0_11_2/a_484_472# 0.0027f
C1674 _07_/ZN output14/a_224_472# 0.05996f
C1675 FILLER_0_11_2/a_4604_375# FILLER_0_10_37/a_572_375# 0.026339f
C1676 FILLER_0_14_37/a_1468_375# FILLER_0_15_40/a_1020_375# 0.026339f
C1677 _16_/I FILLER_0_12_37/a_1020_375# 0.016091f
C1678 FILLER_0_11_72/a_4156_375# vdd 0.007088f
C1679 FILLER_0_8_12/a_1020_375# vdd 0.02589f
C1680 output_signal_plus[7] output_signal_plus[6] 0.27768f
C1681 _15_/I FILLER_0_11_2/a_6844_375# 0.007111f
C1682 _17_/I FILLER_0_14_37/a_1916_375# 0.018729f
C1683 FILLER_0_11_72/a_2724_472# FILLER_0_13_72/a_2812_375# 0.001512f
C1684 vdd FILLER_0_9_66/a_124_375# 0.042248f
C1685 _15_/I FILLER_0_11_2/a_4604_375# 0.007111f
C1686 FILLER_0_4_37/a_6308_472# FILLER_0_3_72/a_2364_375# 0.001597f
C1687 _19_/Z output_signal_plus[9] 0.025942f
C1688 FILLER_0_15_56/a_572_375# _18_/I 0.01418f
C1689 FILLER_0_12_12/a_124_375# _17_/I 0.002388f
C1690 FILLER_0_15_64/a_124_375# FILLER_0_15_56/a_572_375# 0.012001f
C1691 _09_/ZN FILLER_0_11_72/a_6308_472# 0.004262f
C1692 FILLER_0_7_2/a_6756_472# FILLER_0_8_37/a_2812_375# 0.001597f
C1693 vdd FILLER_0_14_37/a_36_472# 0.108844f
C1694 FILLER_0_11_72/a_6396_375# _10_/Z 0.048359f
C1695 FILLER_0_2_2/a_1916_375# _10_/I 0.001061f
C1696 _12_/I FILLER_0_5_72/a_1380_472# 0.003805f
C1697 FILLER_0_7_2/a_4068_472# vdd 0.002735f
C1698 FILLER_0_7_2/a_4964_472# _12_/I 0.004669f
C1699 _18_/I FILLER_0_16_36/a_2276_472# 0.001782f
C1700 FILLER_0_4_2/a_2364_375# FILLER_0_6_2/a_2276_472# 0.0027f
C1701 _16_/I FILLER_0_12_12/a_484_472# 0.01779f
C1702 _15_/I FILLER_0_11_2/a_3260_375# 0.007211f
C1703 output25/a_224_472# _15_/I 0.002599f
C1704 _13_/I input4/a_36_113# 0.004042f
C1705 vdd FILLER_0_6_2/a_1468_375# -0.00495f
C1706 input_signal[2] FILLER_0_2_2/a_484_472# 0.009373f
C1707 _01_/ZN output_signal_minus[0] 0.005845f
C1708 FILLER_0_2_107/a_1468_375# output_signal_minus[6] 0.001064f
C1709 _13_/I FILLER_0_5_104/a_36_472# 0.020094f
C1710 _09_/ZN FILLER_0_12_107/a_932_472# 0.006746f
C1711 FILLER_0_6_37/a_6308_472# _14_/I 0.001167f
C1712 FILLER_0_5_44/a_572_375# _12_/I 0.001706f
C1713 FILLER_0_4_37/a_5052_375# vdd 0.007304f
C1714 FILLER_0_14_37/a_6756_472# FILLER_0_13_72/a_2812_375# 0.001597f
C1715 output_signal_minus[9] FILLER_0_0_70/a_124_375# 0.011852f
C1716 _16_/I FILLER_0_14_12/a_36_472# 0.001667f
C1717 _11_/I FILLER_0_4_37/a_1828_472# 0.014431f
C1718 _13_/I FILLER_0_6_37/a_4068_472# 0.003481f
C1719 FILLER_0_9_2/a_36_472# input_signal[4] 0.001957f
C1720 FILLER_0_13_2/a_572_375# input_signal[7] 0.007169f
C1721 _12_/I FILLER_0_5_72/a_2724_472# 0.003805f
C1722 FILLER_0_2_2/a_2276_472# _10_/I 0.002545f
C1723 _15_/I FILLER_0_12_37/a_1380_472# 0.001368f
C1724 _14_/I FILLER_0_8_37/a_6396_375# 0.01418f
C1725 FILLER_0_5_44/a_36_472# _12_/I 0.003805f
C1726 FILLER_0_15_8/a_36_472# vdd 0.022495f
C1727 _16_/I _16_/Z 0.018114f
C1728 vdd FILLER_0_7_66/a_36_472# 0.097097f
C1729 FILLER_0_7_72/a_1020_375# FILLER_0_6_37/a_4964_472# 0.001723f
C1730 FILLER_0_11_72/a_1468_375# FILLER_0_10_37/a_5500_375# 0.026339f
C1731 FILLER_0_9_104/a_124_375# FILLER_0_9_72/a_3260_375# 0.012222f
C1732 FILLER_0_14_37/a_2276_472# FILLER_0_12_37/a_2364_375# 0.001512f
C1733 vdd FILLER_0_9_2/a_3620_472# 0.005895f
C1734 _11_/I FILLER_0_2_37/a_6396_375# 0.001418f
C1735 FILLER_0_13_2/a_4604_375# FILLER_0_11_2/a_4516_472# 0.001512f
C1736 FILLER_0_0_142/a_572_375# _00_/ZN 0.028887f
C1737 FILLER_0_11_2/a_6308_472# vdd 0.028286f
C1738 FILLER_0_10_12/a_572_375# FILLER_0_12_12/a_484_472# 0.0027f
C1739 FILLER_0_1_12/a_1828_472# _10_/I 0.006408f
C1740 FILLER_0_0_36/a_1828_472# _10_/I 0.016187f
C1741 FILLER_0_11_72/a_2364_375# FILLER_0_10_37/a_6308_472# 0.001723f
C1742 FILLER_0_0_36/a_1916_375# _10_/I 0.015932f
C1743 FILLER_0_6_2/a_1916_375# FILLER_0_5_12/a_932_472# 0.001543f
C1744 FILLER_0_5_44/a_1468_375# FILLER_0_4_37/a_2364_375# 0.026339f
C1745 _11_/I _13_/Z 0.287692f
C1746 _13_/I FILLER_0_6_2/a_2364_375# 0.001706f
C1747 vdd output_signal_minus[4] 0.437957f
C1748 _10_/a_36_160# _06_/ZN 0.022884f
C1749 _12_/I FILLER_0_6_101/a_124_375# 0.017235f
C1750 _16_/I FILLER_0_12_12/a_1380_472# 0.017477f
C1751 _00_/ZN FILLER_0_0_104/a_124_375# 0.01937f
C1752 FILLER_0_7_2/a_2276_472# FILLER_0_8_12/a_1020_375# 0.001543f
C1753 input_signal[5] input_signal[4] 0.060075f
C1754 FILLER_0_10_37/a_4516_472# vdd 0.002735f
C1755 output23/a_224_472# output_signal_plus[1] 0.045278f
C1756 _18_/I output26/a_224_472# 0.026338f
C1757 vdd FILLER_0_10_37/a_5860_472# 0.008907f
C1758 vdd FILLER_0_3_12/a_124_375# 0.03382f
C1759 FILLER_0_13_72/a_3172_472# output29/a_224_472# 0.001243f
C1760 output21/a_224_472# FILLER_0_16_104/a_36_472# 0.003196f
C1761 input_signal[3] input_signal[4] 0.002245f
C1762 _00_/ZN _14_/a_36_113# 0.001745f
C1763 _11_/I _14_/I 0.380222f
C1764 FILLER_0_4_37/a_1916_375# vdd 0.016751f
C1765 output_signal_minus[3] _06_/ZN 0.034329f
C1766 FILLER_0_6_37/a_5412_472# FILLER_0_7_72/a_1468_375# 0.001723f
C1767 _14_/I FILLER_0_7_72/a_2276_472# 0.008683f
C1768 FILLER_0_2_107/a_932_472# _01_/ZN 0.002848f
C1769 FILLER_0_4_37/a_5412_472# FILLER_0_5_72/a_1468_375# 0.001723f
C1770 _09_/ZN FILLER_0_11_72/a_4156_375# 0.002408f
C1771 vdd FILLER_0_12_37/a_6844_375# 0.013514f
C1772 _16_/I FILLER_0_13_2/a_1916_375# 0.00233f
C1773 _13_/I FILLER_0_6_37/a_3260_375# 0.001706f
C1774 FILLER_0_14_107/a_36_472# vdd 0.110617f
C1775 output24/a_224_472# output_signal_plus[4] 0.001204f
C1776 _08_/ZN _10_/Z 0.121907f
C1777 FILLER_0_3_72/a_1916_375# FILLER_0_4_37/a_5860_472# 0.001597f
C1778 FILLER_0_10_107/a_1468_375# FILLER_0_11_72/a_5412_472# 0.001723f
C1779 FILLER_0_11_72/a_2812_375# FILLER_0_12_37/a_6756_472# 0.001597f
C1780 FILLER_0_10_107/a_1020_375# FILLER_0_11_72/a_5052_375# 0.026339f
C1781 FILLER_0_12_37/a_1380_472# FILLER_0_10_37/a_1468_375# 0.001512f
C1782 FILLER_0_7_72/a_1468_375# vdd 0.007205f
C1783 _14_/Z _14_/a_36_113# 0.005715f
C1784 _11_/I FILLER_0_4_37/a_2276_472# 0.014431f
C1785 FILLER_0_2_37/a_6308_472# output_signal_minus[0] 0.001292f
C1786 FILLER_0_13_2/a_124_375# input_signal[7] 0.007233f
C1787 input_signal[5] FILLER_0_10_12/a_484_472# 0.001984f
C1788 FILLER_0_14_107/a_484_472# vdd 0.004716f
C1789 output_signal_minus[6] _10_/I 0.015552f
C1790 FILLER_0_12_107/a_572_375# _17_/I 0.002302f
C1791 FILLER_0_7_2/a_4964_472# FILLER_0_8_37/a_1020_375# 0.001597f
C1792 FILLER_0_7_2/a_5860_472# _14_/I 0.008683f
C1793 _18_/I FILLER_0_14_37/a_4516_472# 0.001526f
C1794 FILLER_0_12_37/a_36_472# FILLER_0_12_28/a_124_375# 0.007947f
C1795 input_signal[0] FILLER_0_0_12/a_484_472# 0.002568f
C1796 FILLER_0_13_72/a_484_472# FILLER_0_14_37/a_4516_472# 0.026657f
C1797 vdd FILLER_0_8_37/a_6756_472# 0.015684f
C1798 vdd FILLER_0_2_37/a_1828_472# 0.011772f
C1799 _15_/I _15_/Z 0.269871f
C1800 FILLER_0_9_2/a_6396_375# FILLER_0_8_37/a_2364_375# 0.026339f
C1801 _14_/I FILLER_0_9_2/a_2812_375# 0.005414f
C1802 FILLER_0_5_12/a_1916_375# FILLER_0_3_12/a_1828_472# 0.0027f
C1803 _07_/ZN _01_/ZN 0.077572f
C1804 FILLER_0_9_72/a_1380_472# FILLER_0_10_37/a_5412_472# 0.026657f
C1805 FILLER_0_1_12/a_2364_375# _10_/I 0.008299f
C1806 _16_/I FILLER_0_10_37/a_2364_375# 0.001157f
C1807 FILLER_0_7_66/a_124_375# FILLER_0_6_37/a_3260_375# 0.026339f
C1808 _11_/I FILLER_0_5_12/a_36_472# 0.001913f
C1809 FILLER_0_14_37/a_572_375# vdd 0.007106f
C1810 FILLER_0_4_37/a_4068_472# FILLER_0_3_72/a_36_472# 0.026657f
C1811 _10_/I FILLER_0_1_12/a_1468_375# 0.008103f
C1812 _12_/I FILLER_0_5_72/a_2276_472# 0.003805f
C1813 FILLER_0_8_37/a_124_375# FILLER_0_9_2/a_4068_472# 0.001723f
C1814 _11_/I FILLER_0_3_12/a_1828_472# 0.008733f
C1815 _18_/a_36_113# output26/a_224_472# 0.001339f
C1816 FILLER_0_12_37/a_4964_472# vdd 0.005073f
C1817 FILLER_0_5_104/a_484_472# vdd 0.007483f
C1818 FILLER_0_4_37/a_484_472# FILLER_0_3_12/a_3172_472# 0.026657f
C1819 FILLER_0_7_2/a_6308_472# _12_/I 0.002625f
C1820 _19_/I output29/a_224_472# 0.010052f
C1821 FILLER_0_11_2/a_2364_375# FILLER_0_10_12/a_1380_472# 0.001684f
C1822 _00_/ZN FILLER_0_0_142/a_124_375# 0.012159f
C1823 _00_/ZN output24/a_224_472# 0.008306f
C1824 FILLER_0_10_37/a_4068_472# FILLER_0_8_37/a_4156_375# 0.001512f
C1825 output_signal_plus[8] FILLER_0_14_37/a_6844_375# 0.001633f
C1826 _15_/I FILLER_0_9_72/a_3260_375# 0.006125f
C1827 vdd FILLER_0_1_44/a_484_472# 0.007487f
C1828 _15_/I FILLER_0_11_2/a_6756_472# 0.005458f
C1829 FILLER_0_0_70/a_124_375# output20/a_224_472# 0.011959f
C1830 _13_/I FILLER_0_5_12/a_1020_375# 0.016091f
C1831 _14_/I FILLER_0_8_37/a_4964_472# 0.014431f
C1832 input_signal[6] _16_/I 0.233494f
C1833 _15_/I FILLER_0_10_37/a_4156_375# 0.018729f
C1834 _11_/I FILLER_0_2_2/a_3260_375# 0.00346f
C1835 _09_/ZN output_signal_minus[4] 0.091457f
C1836 _15_/I FILLER_0_9_2/a_6396_375# 0.006125f
C1837 _14_/I FILLER_0_6_37/a_4604_375# 0.002835f
C1838 _11_/I FILLER_0_2_107/a_1020_375# 0.002387f
C1839 FILLER_0_6_37/a_5860_472# FILLER_0_5_72/a_1828_472# 0.026657f
C1840 _14_/I FILLER_0_6_37/a_1916_375# 0.003066f
C1841 FILLER_0_6_37/a_6844_375# FILLER_0_8_37/a_6756_472# 0.001512f
C1842 FILLER_0_11_2/a_3260_375# FILLER_0_9_2/a_3172_472# 0.0027f
C1843 FILLER_0_9_72/a_572_375# FILLER_0_10_37/a_4516_472# 0.001597f
C1844 FILLER_0_3_72/a_2724_472# FILLER_0_5_72/a_2812_375# 0.001512f
C1845 output24/a_224_472# _14_/Z 0.061535f
C1846 FILLER_0_0_36/a_3260_375# vdd 0.019402f
C1847 FILLER_0_1_72/a_932_472# _10_/I 0.006408f
C1848 FILLER_0_15_8/a_2364_375# vdd -0.010699f
C1849 _15_/I FILLER_0_9_2/a_1380_472# 0.00656f
C1850 _18_/I output29/a_224_472# 0.111864f
C1851 output_signal_minus[8] FILLER_0_0_142/a_484_472# 0.012073f
C1852 FILLER_0_5_72/a_3172_472# vdd 0.007853f
C1853 FILLER_0_7_2/a_6396_375# vdd 0.014428f
C1854 _02_/ZN vdd 0.034615f
C1855 FILLER_0_12_101/a_124_375# FILLER_0_12_107/a_124_375# 0.005439f
C1856 FILLER_0_11_72/a_1916_375# vdd 0.009594f
C1857 vdd _10_/Z 1.197471f
C1858 FILLER_0_14_37/a_5860_472# FILLER_0_13_72/a_1828_472# 0.026657f
C1859 _16_/I FILLER_0_11_72/a_5412_472# 0.006073f
C1860 output_signal_minus[2] net15 0.003648f
C1861 FILLER_0_16_104/a_124_375# output_signal_plus[0] 0.011852f
C1862 _15_/I output_signal_plus[1] 0.266874f
C1863 _11_/I FILLER_0_3_44/a_1380_472# 0.008683f
C1864 FILLER_0_8_37/a_36_472# FILLER_0_8_28/a_36_472# 0.001963f
C1865 FILLER_0_13_2/a_6308_472# _16_/I 0.002625f
C1866 FILLER_0_8_37/a_1020_375# FILLER_0_10_37/a_932_472# 0.001512f
C1867 FILLER_0_2_107/a_484_472# _01_/ZN 0.030904f
C1868 vdd FILLER_0_1_44/a_1468_375# 0.02682f
C1869 vdd FILLER_0_4_101/a_36_472# 0.098288f
C1870 _17_/I FILLER_0_14_37/a_1828_472# 0.015502f
C1871 FILLER_0_10_12/a_36_472# vdd 0.015471f
C1872 output_signal_plus[7] _18_/Z 0.66687f
C1873 vdd FILLER_0_1_12/a_572_375# 0.020697f
C1874 _15_/I FILLER_0_10_37/a_5948_375# 0.018729f
C1875 _08_/ZN _12_/I 0.046319f
C1876 output_signal_plus[5] _16_/Z 0.157485f
C1877 output14/a_224_472# _04_/ZN 0.019697f
C1878 FILLER_0_15_40/a_932_472# _19_/I 0.001782f
C1879 _17_/I FILLER_0_13_2/a_4964_472# 0.006506f
C1880 _15_/I FILLER_0_10_37/a_1916_375# 0.018729f
C1881 FILLER_0_9_2/a_1828_472# _15_/I 0.00656f
C1882 output15/a_224_472# _08_/ZN 0.016157f
C1883 FILLER_0_15_72/a_572_375# vdd 0.002455f
C1884 FILLER_0_10_37/a_2276_472# vdd 0.037602f
C1885 vdd FILLER_0_12_37/a_2812_375# 0.009304f
C1886 _11_/Z _11_/a_36_113# 0.027105f
C1887 output18/a_224_472# output_signal_minus[7] 0.031258f
C1888 FILLER_0_16_104/a_124_375# output_signal_plus[8] 0.023881f
C1889 _17_/I FILLER_0_12_37/a_5052_375# 0.002388f
C1890 FILLER_0_13_2/a_1828_472# FILLER_0_14_12/a_572_375# 0.001543f
C1891 FILLER_0_3_60/a_484_472# FILLER_0_4_37/a_3172_472# 0.026657f
C1892 FILLER_0_4_37/a_4604_375# FILLER_0_5_72/a_572_375# 0.026339f
C1893 FILLER_0_4_2/a_1020_375# FILLER_0_5_12/a_36_472# 0.001684f
C1894 input_signal[9] input9/a_36_113# 0.01895f
C1895 FILLER_0_14_107/a_484_472# _09_/ZN 0.001293f
C1896 FILLER_0_10_107/a_484_472# vdd 0.005094f
C1897 output23/a_224_472# output_signal_plus[2] 0.014303f
C1898 FILLER_0_3_72/a_3260_375# FILLER_0_4_101/a_36_472# 0.001597f
C1899 FILLER_0_15_64/a_36_472# FILLER_0_15_56/a_572_375# 0.086635f
C1900 FILLER_0_15_8/a_1020_375# FILLER_0_16_18/a_36_472# 0.001543f
C1901 output24/a_224_472# output_signal_plus[3] 0.008471f
C1902 FILLER_0_7_104/a_484_472# _12_/I 0.004669f
C1903 FILLER_0_0_12/a_572_375# vdd 0.016551f
C1904 FILLER_0_8_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001597f
C1905 FILLER_0_5_44/a_124_375# FILLER_0_4_37/a_1020_375# 0.026339f
C1906 FILLER_0_8_37/a_1468_375# vdd 0.008806f
C1907 vdd FILLER_0_9_72/a_1828_472# 0.008296f
C1908 input3/a_36_113# vdd 0.121003f
C1909 vdd FILLER_0_7_2/a_5052_375# 0.009467f
C1910 output13/a_224_472# _10_/Z 0.029067f
C1911 FILLER_0_12_37/a_4068_472# FILLER_0_11_72/a_36_472# 0.026657f
C1912 FILLER_0_8_37/a_6308_472# vdd 0.020611f
C1913 FILLER_0_5_12/a_1468_375# _12_/I 0.001706f
C1914 vdd input_signal[9] 0.217952f
C1915 vdd FILLER_0_16_18/a_572_375# 0.006965f
C1916 FILLER_0_8_37/a_5052_375# _15_/I 0.002388f
C1917 FILLER_0_0_12/a_932_472# _10_/I 0.016279f
C1918 _16_/I FILLER_0_13_2/a_4068_472# 0.004669f
C1919 FILLER_0_7_2/a_484_472# _12_/I 0.002259f
C1920 _13_/I FILLER_0_6_2/a_932_472# 0.003922f
C1921 FILLER_0_15_40/a_932_472# _18_/I 0.014431f
C1922 _16_/I FILLER_0_11_2/a_6844_375# 0.007169f
C1923 FILLER_0_14_115/a_36_472# vdd 0.086171f
C1924 FILLER_0_6_37/a_2724_472# FILLER_0_5_60/a_124_375# 0.001597f
C1925 FILLER_0_0_142/a_36_472# _00_/ZN 0.009873f
C1926 _15_/I FILLER_0_11_2/a_3172_472# 0.005458f
C1927 output17/a_224_472# _10_/Z 0.040736f
C1928 FILLER_0_14_101/a_36_472# vdd 0.098751f
C1929 FILLER_0_13_72/a_2276_472# _16_/I 0.004669f
C1930 FILLER_0_11_2/a_4604_375# _16_/I 0.007169f
C1931 FILLER_0_9_104/a_484_472# _14_/I 0.004017f
C1932 vdd FILLER_0_15_72/a_124_375# 0.013594f
C1933 _11_/Z FILLER_0_10_107/a_1380_472# 0.038912f
C1934 FILLER_0_12_37/a_4068_472# vdd 0.002856f
C1935 _13_/I FILLER_0_6_37/a_5500_375# 0.001706f
C1936 _12_/a_36_113# _14_/I 0.044553f
C1937 _17_/I FILLER_0_15_8/a_932_472# 0.00338f
C1938 vdd FILLER_0_14_37/a_5948_375# 0.008812f
C1939 _00_/ZN FILLER_0_0_104/a_36_472# 0.02331f
C1940 _16_/I FILLER_0_11_2/a_3260_375# 0.007169f
C1941 _19_/a_36_113# _17_/I 0.00777f
C1942 output25/a_224_472# _16_/I 0.171365f
C1943 _12_/Z _14_/I 0.476815f
C1944 _08_/ZN output_signal_plus[4] 0.266951f
C1945 _15_/I FILLER_0_11_66/a_36_472# 0.005458f
C1946 FILLER_0_13_2/a_6396_375# FILLER_0_12_37/a_2364_375# 0.026339f
C1947 _11_/I FILLER_0_5_44/a_124_375# 0.004712f
C1948 _16_/I output28/a_224_472# 0.035719f
C1949 FILLER_0_1_72/a_1468_375# output11/a_224_472# 0.023259f
C1950 FILLER_0_14_12/a_1380_472# _16_/I 0.001667f
C1951 FILLER_0_6_37/a_5412_472# _12_/I 0.017477f
C1952 FILLER_0_3_72/a_124_375# FILLER_0_2_37/a_4068_472# 0.001723f
C1953 FILLER_0_12_37/a_1380_472# _16_/I 0.017477f
C1954 _15_/I FILLER_0_11_72/a_3708_375# 0.007218f
C1955 _11_/I FILLER_0_3_104/a_572_375# 0.008393f
C1956 _17_/I FILLER_0_14_37/a_5052_375# 0.018729f
C1957 FILLER_0_3_60/a_124_375# FILLER_0_2_37/a_2724_472# 0.001723f
C1958 FILLER_0_13_104/a_36_472# _16_/I 0.004669f
C1959 output19/a_224_472# _08_/ZN 0.016961f
C1960 _13_/I FILLER_0_6_37/a_5052_375# 0.001706f
C1961 FILLER_0_1_12/a_3172_472# FILLER_0_2_37/a_484_472# 0.026657f
C1962 output_signal_minus[8] net15 0.00927f
C1963 _12_/I FILLER_0_5_12/a_124_375# 0.005257f
C1964 FILLER_0_16_18/a_124_375# input9/a_36_113# 0.002124f
C1965 FILLER_0_9_72/a_932_472# _14_/I 0.004017f
C1966 _09_/ZN _10_/Z 0.128015f
C1967 FILLER_0_13_2/a_484_472# input_signal[7] 0.007674f
C1968 vdd _12_/I 1.548303f
C1969 FILLER_0_11_2/a_3708_375# vdd 0.018728f
C1970 FILLER_0_14_28/a_36_472# _18_/I 0.001526f
C1971 FILLER_0_13_72/a_1380_472# vdd 0.006325f
C1972 FILLER_0_1_72/a_1380_472# vdd 0.007849f
C1973 FILLER_0_5_44/a_932_472# FILLER_0_6_37/a_1828_472# 0.026657f
C1974 output15/a_224_472# vdd 0.106428f
C1975 FILLER_0_8_107/a_124_375# vdd 0.014813f
C1976 vdd FILLER_0_4_37/a_572_375# 0.006843f
C1977 _16_/Z output_signal_plus[6] 0.087721f
C1978 FILLER_0_6_37/a_124_375# FILLER_0_6_2/a_3260_375# 0.004426f
C1979 FILLER_0_5_60/a_36_472# FILLER_0_6_37/a_2724_472# 0.026657f
C1980 FILLER_0_6_37/a_3708_375# _12_/I 0.016091f
C1981 FILLER_0_11_72/a_1468_375# _15_/I 0.007126f
C1982 FILLER_0_7_2/a_4604_375# vdd 0.007747f
C1983 vdd FILLER_0_16_18/a_124_375# 0.039949f
C1984 FILLER_0_4_37/a_484_472# _11_/I 0.014431f
C1985 _14_/I FILLER_0_7_2/a_6844_375# 0.008393f
C1986 _15_/I FILLER_0_8_37/a_4156_375# 0.002049f
C1987 FILLER_0_10_37/a_124_375# FILLER_0_9_2/a_4068_472# 0.001597f
C1988 _17_/I FILLER_0_13_2/a_3172_472# 0.006606f
C1989 FILLER_0_16_104/a_124_375# _19_/Z 0.022181f
C1990 input2/a_36_113# input3/a_36_113# 0.001442f
C1991 FILLER_0_14_37/a_1916_375# FILLER_0_15_40/a_1468_375# 0.026339f
C1992 FILLER_0_11_72/a_1828_472# _15_/I 0.005458f
C1993 FILLER_0_1_44/a_36_472# _10_/I 0.006408f
C1994 FILLER_0_14_28/a_36_472# FILLER_0_14_12/a_1468_375# 0.086635f
C1995 _16_/I FILLER_0_13_104/a_484_472# 0.004669f
C1996 _00_/ZN _08_/ZN 0.104462f
C1997 FILLER_0_9_72/a_36_472# vdd 0.108637f
C1998 vdd FILLER_0_3_104/a_124_375# 0.028196f
C1999 FILLER_0_3_72/a_2364_375# FILLER_0_2_37/a_6396_375# 0.026339f
C2000 FILLER_0_0_142/a_572_375# _06_/ZN 0.002444f
C2001 _10_/I FILLER_0_0_142/a_484_472# 0.010562f
C2002 _13_/I output_signal_minus[7] 0.009819f
C2003 FILLER_0_9_2/a_4516_472# FILLER_0_11_2/a_4604_375# 0.001512f
C2004 _09_/ZN FILLER_0_10_107/a_484_472# 0.003007f
C2005 FILLER_0_0_142/a_572_375# _10_/a_36_160# 0.001925f
C2006 vdd FILLER_0_11_2/a_1468_375# 0.027811f
C2007 FILLER_0_11_2/a_2364_375# FILLER_0_12_12/a_1380_472# 0.001543f
C2008 FILLER_0_3_12/a_3260_375# _11_/I 0.008393f
C2009 _15_/I output_signal_plus[2] 0.39846f
C2010 FILLER_0_1_12/a_3260_375# FILLER_0_2_37/a_484_472# 0.001597f
C2011 _13_/I FILLER_0_5_72/a_2812_375# 0.016337f
C2012 output13/a_224_472# _12_/I 0.019965f
C2013 FILLER_0_3_72/a_572_375# FILLER_0_4_37/a_4516_472# 0.001597f
C2014 _14_/I output_signal_minus[6] 0.048085f
C2015 output15/a_224_472# output13/a_224_472# 0.004177f
C2016 FILLER_0_15_40/a_1380_472# FILLER_0_15_56/a_36_472# 0.013277f
C2017 FILLER_0_13_66/a_124_375# FILLER_0_13_72/a_124_375# 0.005439f
C2018 FILLER_0_4_37/a_4604_375# FILLER_0_6_37/a_4516_472# 0.001512f
C2019 _14_/I FILLER_0_7_2/a_1020_375# 0.008393f
C2020 _14_/Z _08_/ZN 0.135194f
C2021 _13_/I FILLER_0_6_37/a_2724_472# 0.003818f
C2022 FILLER_0_6_37/a_6844_375# _12_/I 0.016091f
C2023 FILLER_0_14_37/a_5860_472# FILLER_0_13_72/a_1916_375# 0.001597f
C2024 FILLER_0_3_72/a_3260_375# FILLER_0_3_104/a_124_375# 0.012221f
C2025 _09_/ZN FILLER_0_14_115/a_36_472# 0.006052f
C2026 FILLER_0_15_8/a_1020_375# FILLER_0_14_12/a_572_375# 0.05841f
C2027 FILLER_0_11_2/a_3620_472# vdd 0.005895f
C2028 FILLER_0_9_2/a_932_472# _15_/I 0.005193f
C2029 vdd FILLER_0_4_2/a_3172_472# 0.012967f
C2030 FILLER_0_15_40/a_1380_472# vdd 0.00607f
C2031 _11_/I output23/a_224_472# 0.010749f
C2032 _13_/I FILLER_0_5_72/a_1828_472# 0.017477f
C2033 FILLER_0_15_8/a_1468_375# FILLER_0_16_18/a_484_472# 0.001543f
C2034 _17_/I _08_/ZN 0.032158f
C2035 FILLER_0_8_37/a_124_375# vdd 0.013676f
C2036 FILLER_0_12_37/a_1468_375# vdd 0.008961f
C2037 FILLER_0_10_12/a_1020_375# _15_/I 0.018729f
C2038 input_signal[1] FILLER_0_1_12/a_572_375# 0.00186f
C2039 _14_/a_36_113# _06_/ZN 0.137199f
C2040 vdd FILLER_0_13_2/a_36_472# 0.105578f
C2041 output_signal_plus[4] vdd 0.184117f
C2042 _13_/I FILLER_0_4_37/a_4604_375# 0.005726f
C2043 FILLER_0_9_72/a_124_375# vdd 0.011994f
C2044 vdd FILLER_0_5_12/a_1380_472# 0.011134f
C2045 FILLER_0_16_104/a_36_472# _18_/Z 0.037282f
C2046 FILLER_0_9_104/a_36_472# vdd 0.093924f
C2047 FILLER_0_0_36/a_1380_472# _10_/I 0.016187f
C2048 FILLER_0_7_2/a_4516_472# _14_/I 0.008683f
C2049 FILLER_0_5_104/a_124_375# FILLER_0_5_72/a_3260_375# 0.012222f
C2050 input7/a_36_113# vdd 0.12101f
C2051 FILLER_0_10_12/a_36_472# input_signal[5] 0.074078f
C2052 FILLER_0_4_37/a_124_375# vdd 0.014132f
C2053 FILLER_0_9_72/a_2724_472# FILLER_0_11_72/a_2812_375# 0.001512f
C2054 vdd FILLER_0_12_37/a_484_472# 0.00379f
C2055 _14_/I FILLER_0_8_37/a_3172_472# 0.014431f
C2056 _16_/I _15_/Z 0.161007f
C2057 _18_/I FILLER_0_15_8/a_1468_375# 0.014412f
C2058 output19/a_224_472# vdd 0.155541f
C2059 FILLER_0_13_2/a_6308_472# FILLER_0_14_37/a_2364_375# 0.001597f
C2060 _13_/I FILLER_0_4_2/a_2812_375# 0.00577f
C2061 FILLER_0_6_37/a_1020_375# _14_/I 0.003099f
C2062 FILLER_0_12_37/a_4156_375# vdd 0.004039f
C2063 _11_/I FILLER_0_2_2/a_1020_375# 0.012735f
C2064 _16_/I FILLER_0_13_2/a_5500_375# 0.006193f
C2065 FILLER_0_10_12/a_484_472# FILLER_0_9_2/a_1468_375# 0.001543f
C2066 FILLER_0_7_2/a_2276_472# _12_/I 0.004669f
C2067 FILLER_0_5_72/a_36_472# _12_/I 0.003805f
C2068 FILLER_0_11_72/a_1828_472# FILLER_0_13_72/a_1916_375# 0.001512f
C2069 FILLER_0_4_37/a_4964_472# FILLER_0_5_72/a_1020_375# 0.001723f
C2070 FILLER_0_6_37/a_932_472# _14_/I 0.001219f
C2071 _16_/I FILLER_0_12_107/a_1020_375# 0.016091f
C2072 FILLER_0_5_44/a_36_472# FILLER_0_5_12/a_3260_375# 0.086905f
C2073 FILLER_0_6_37/a_2812_375# FILLER_0_7_2/a_6844_375# 0.026339f
C2074 FILLER_0_2_2/a_1380_472# FILLER_0_3_12/a_124_375# 0.001684f
C2075 FILLER_0_9_72/a_2724_472# _14_/I 0.001634f
C2076 output_signal_plus[3] _08_/ZN 0.107889f
C2077 _14_/I FILLER_0_9_2/a_6308_472# 0.002295f
C2078 FILLER_0_14_107/a_124_375# _18_/Z 0.029638f
C2079 _07_/ZN output25/a_224_472# 0.00885f
C2080 FILLER_0_14_37/a_932_472# _16_/I 0.001667f
C2081 FILLER_0_12_12/a_484_472# FILLER_0_13_2/a_1468_375# 0.001684f
C2082 FILLER_0_13_2/a_4604_375# FILLER_0_12_37/a_572_375# 0.026339f
C2083 _09_/ZN _12_/I 0.10888f
C2084 _02_/ZN output_signal_minus[2] 0.027053f
C2085 FILLER_0_11_2/a_6756_472# _16_/I 0.007542f
C2086 FILLER_0_11_2/a_6308_472# FILLER_0_13_2/a_6396_375# 0.001512f
C2087 _11_/I FILLER_0_3_72/a_2724_472# 0.008683f
C2088 output15/a_224_472# _09_/ZN 0.083396f
C2089 output_signal_minus[2] _10_/Z 0.100524f
C2090 vdd FILLER_0_7_72/a_1916_375# 0.009597f
C2091 FILLER_0_10_12/a_1468_375# FILLER_0_11_2/a_2724_472# 0.001684f
C2092 vdd FILLER_0_8_37/a_1020_375# 0.006698f
C2093 _00_/ZN vdd 1.606974f
C2094 _16_/I FILLER_0_10_37/a_4156_375# 0.002086f
C2095 _18_/I FILLER_0_14_37/a_36_472# 0.001526f
C2096 input3/a_36_113# input_signal[3] 0.003334f
C2097 FILLER_0_15_8/a_36_472# _19_/I 0.008641f
C2098 FILLER_0_12_12/a_572_375# vdd 0.052349f
C2099 _15_/I FILLER_0_8_37/a_6396_375# 0.001106f
C2100 input_signal[2] FILLER_0_2_2/a_124_375# 0.045794f
C2101 FILLER_0_8_107/a_572_375# _11_/Z 0.005144f
C2102 FILLER_0_13_2/a_5052_375# _16_/I 0.006193f
C2103 FILLER_0_8_37/a_5860_472# FILLER_0_7_72/a_1828_472# 0.026657f
C2104 output27/a_224_472# output28/a_224_472# 0.010315f
C2105 FILLER_0_0_142/a_124_375# _10_/a_36_160# 0.02985f
C2106 FILLER_0_3_72/a_2812_375# FILLER_0_4_37/a_6756_472# 0.001597f
C2107 _13_/I FILLER_0_5_60/a_572_375# 0.017949f
C2108 _11_/I FILLER_0_5_72/a_572_375# 0.004712f
C2109 output17/a_224_472# output19/a_224_472# 0.005241f
C2110 FILLER_0_1_72/a_1468_375# _10_/I 0.008103f
C2111 FILLER_0_1_72/a_124_375# vdd 0.028611f
C2112 _14_/Z vdd 0.422708f
C2113 _14_/I FILLER_0_7_72/a_1828_472# 0.008683f
C2114 output_signal_plus[5] output28/a_224_472# 0.002451f
C2115 _17_/I vdd 2.044431f
C2116 FILLER_0_8_37/a_572_375# _14_/I 0.01418f
C2117 vdd FILLER_0_15_8/a_124_375# 0.029156f
C2118 _18_/I FILLER_0_15_8/a_36_472# 0.004473f
C2119 FILLER_0_10_101/a_124_375# FILLER_0_10_37/a_6844_375# 0.012001f
C2120 FILLER_0_2_37/a_6756_472# vdd 0.013974f
C2121 _15_/I FILLER_0_11_72/a_3260_375# 0.007126f
C2122 vdd FILLER_0_4_107/a_124_375# 0.014813f
C2123 _16_/I FILLER_0_10_37/a_5948_375# 0.002327f
C2124 FILLER_0_11_66/a_36_472# FILLER_0_10_37/a_3260_375# 0.001723f
C2125 FILLER_0_7_2/a_5500_375# _12_/I 0.006193f
C2126 _15_/I FILLER_0_11_2/a_2724_472# 0.005458f
C2127 _13_/I FILLER_0_5_12/a_3172_472# 0.017477f
C2128 FILLER_0_7_2/a_5948_375# _14_/I 0.008393f
C2129 FILLER_0_12_37/a_4604_375# FILLER_0_14_37/a_4516_472# 0.001512f
C2130 FILLER_0_10_37/a_1916_375# _16_/I 0.002323f
C2131 FILLER_0_0_36/a_3260_375# FILLER_0_1_60/a_572_375# 0.05841f
C2132 FILLER_0_12_37/a_1828_472# FILLER_0_11_2/a_5860_472# 0.026657f
C2133 _09_/ZN output_signal_plus[4] 0.003516f
C2134 output_signal_minus[6] output16/a_224_472# 0.105215f
C2135 FILLER_0_7_72/a_572_375# _14_/I 0.005f
C2136 FILLER_0_8_37/a_4516_472# vdd 0.002735f
C2137 FILLER_0_6_2/a_484_472# _12_/I 0.027722f
C2138 FILLER_0_7_2/a_4068_472# FILLER_0_6_37/a_124_375# 0.001723f
C2139 FILLER_0_13_2/a_4604_375# _16_/I 0.006193f
C2140 _11_/I FILLER_0_5_60/a_124_375# 0.004712f
C2141 _11_/I _15_/I 0.002206f
C2142 output_signal_minus[5] _08_/ZN 0.420191f
C2143 FILLER_0_3_44/a_572_375# vdd 0.008603f
C2144 _12_/I FILLER_0_5_12/a_932_472# 0.004687f
C2145 FILLER_0_12_12/a_124_375# FILLER_0_11_2/a_1380_472# 0.001543f
C2146 input_signal[3] _12_/I 0.120616f
C2147 FILLER_0_5_12/a_2812_375# FILLER_0_4_37/a_124_375# 0.026339f
C2148 _14_/Z output13/a_224_472# 0.00595f
C2149 _09_/ZN output19/a_224_472# 0.052368f
C2150 output_signal_plus[3] vdd 0.152275f
C2151 FILLER_0_15_2/a_124_375# input_signal[8] 0.080164f
C2152 FILLER_0_8_37/a_6844_375# FILLER_0_9_72/a_2812_375# 0.026339f
C2153 FILLER_0_10_37/a_6844_375# vdd 0.012466f
C2154 FILLER_0_8_28/a_36_472# vdd 0.098927f
C2155 FILLER_0_8_12/a_1020_375# FILLER_0_9_2/a_2276_472# 0.001684f
C2156 output_signal_minus[7] output_signal_minus[0] 0.0035f
C2157 _11_/I FILLER_0_3_12/a_36_472# 0.013673f
C2158 FILLER_0_9_72/a_2276_472# FILLER_0_10_37/a_6308_472# 0.026657f
C2159 FILLER_0_11_2/a_3172_472# _16_/I 0.007639f
C2160 FILLER_0_9_2/a_5500_375# vdd 0.011603f
C2161 _11_/I FILLER_0_2_101/a_124_375# 0.00346f
C2162 FILLER_0_13_66/a_36_472# FILLER_0_14_37/a_3260_375# 0.001597f
C2163 FILLER_0_9_2/a_1828_472# FILLER_0_10_12/a_572_375# 0.001543f
C2164 _17_/I FILLER_0_13_2/a_5860_472# 0.006506f
C2165 vdd FILLER_0_12_37/a_3260_375# 0.007161f
C2166 FILLER_0_10_37/a_5052_375# vdd 0.00705f
C2167 _10_/Z output_signal_minus[8] 0.116523f
C2168 FILLER_0_4_2/a_124_375# vdd 0.012902f
C2169 _15_/I FILLER_0_12_37/a_6756_472# 0.001368f
C2170 _13_/I FILLER_0_6_37/a_6308_472# 0.003818f
C2171 FILLER_0_4_37/a_1916_375# FILLER_0_5_44/a_1020_375# 0.026339f
C2172 _15_/I FILLER_0_9_2/a_2812_375# 0.006125f
C2173 _18_/I FILLER_0_14_107/a_36_472# 0.001526f
C2174 _17_/I FILLER_0_13_2/a_2364_375# 0.006125f
C2175 output_signal_minus[2] _12_/I 0.152514f
C2176 _16_/Z _18_/Z 0.008221f
C2177 FILLER_0_12_37/a_1916_375# FILLER_0_14_37/a_1828_472# 0.001512f
C2178 FILLER_0_11_72/a_2364_375# _15_/I 0.005833f
C2179 FILLER_0_10_37/a_6756_472# FILLER_0_9_72/a_2812_375# 0.001597f
C2180 output15/a_224_472# output_signal_minus[2] 0.001224f
C2181 FILLER_0_12_37/a_6396_375# _16_/I 0.016091f
C2182 FILLER_0_0_36/a_2364_375# FILLER_0_1_44/a_1468_375# 0.05841f
C2183 FILLER_0_11_66/a_36_472# _16_/I 0.007542f
C2184 FILLER_0_8_37/a_36_472# FILLER_0_8_28/a_124_375# 0.007947f
C2185 FILLER_0_7_2/a_5412_472# vdd 0.008843f
C2186 _17_/I FILLER_0_13_72/a_932_472# 0.00652f
C2187 vdd FILLER_0_10_37/a_124_375# 0.013676f
C2188 _14_/I FILLER_0_6_2/a_3260_375# 0.003099f
C2189 FILLER_0_14_107/a_484_472# _18_/I 0.002069f
C2190 FILLER_0_14_37/a_1828_472# FILLER_0_15_40/a_1468_375# 0.001723f
C2191 FILLER_0_9_2/a_5052_375# FILLER_0_8_37/a_1020_375# 0.026339f
C2192 FILLER_0_2_37/a_4964_472# FILLER_0_1_72/a_1020_375# 0.001597f
C2193 FILLER_0_7_72/a_2812_375# FILLER_0_5_72/a_2724_472# 0.001512f
C2194 _16_/I FILLER_0_11_72/a_3708_375# 0.007169f
C2195 vdd FILLER_0_10_37/a_3620_472# 0.00818f
C2196 output23/a_224_472# _12_/Z 0.065277f
C2197 _11_/I FILLER_0_2_37/a_2812_375# 0.00346f
C2198 _13_/I FILLER_0_4_37/a_1020_375# 0.005726f
C2199 FILLER_0_6_37/a_2276_472# _12_/I 0.017477f
C2200 FILLER_0_14_37/a_5860_472# _16_/I 0.001667f
C2201 vdd FILLER_0_1_44/a_1020_375# -0.005325f
C2202 FILLER_0_5_60/a_36_472# _11_/I 0.001913f
C2203 FILLER_0_10_37/a_1828_472# vdd 0.010403f
C2204 _15_/I FILLER_0_12_107/a_1380_472# 0.001368f
C2205 FILLER_0_10_107/a_1020_375# FILLER_0_11_72/a_4964_472# 0.001723f
C2206 FILLER_0_2_2/a_1828_472# FILLER_0_3_12/a_572_375# 0.001684f
C2207 output_signal_plus[5] _15_/Z 0.05851f
C2208 FILLER_0_12_12/a_932_472# FILLER_0_13_2/a_1916_375# 0.001684f
C2209 FILLER_0_4_37/a_4964_472# FILLER_0_3_72/a_932_472# 0.026657f
C2210 FILLER_0_13_66/a_36_472# FILLER_0_13_72/a_36_472# 0.003468f
C2211 FILLER_0_12_37/a_1916_375# FILLER_0_11_2/a_5860_472# 0.001597f
C2212 _13_/I FILLER_0_5_12/a_2276_472# 0.017477f
C2213 FILLER_0_4_37/a_6844_375# vdd 0.013417f
C2214 FILLER_0_13_2/a_3260_375# vdd 0.020842f
C2215 FILLER_0_1_72/a_932_472# output20/a_224_472# 0.001699f
C2216 FILLER_0_3_12/a_572_375# FILLER_0_4_2/a_1828_472# 0.001543f
C2217 _18_/I FILLER_0_14_37/a_572_375# 0.003988f
C2218 _09_/ZN _17_/I 0.024311f
C2219 _17_/I FILLER_0_12_37/a_3708_375# 0.002388f
C2220 FILLER_0_10_107/a_572_375# FILLER_0_11_72/a_4516_472# 0.001723f
C2221 FILLER_0_8_37/a_6756_472# FILLER_0_7_72/a_2724_472# 0.026657f
C2222 _11_/I FILLER_0_2_2/a_2364_375# 0.00346f
C2223 FILLER_0_4_37/a_5860_472# FILLER_0_3_72/a_1828_472# 0.026657f
C2224 _15_/I FILLER_0_11_72/a_484_472# 0.005458f
C2225 FILLER_0_7_72/a_1020_375# vdd 0.00558f
C2226 FILLER_0_7_72/a_3260_375# FILLER_0_8_101/a_36_472# 0.001597f
C2227 vdd _13_/a_36_113# 0.089652f
C2228 input_signal[7] input_signal[9] 0.003454f
C2229 _13_/I FILLER_0_5_12/a_1916_375# 0.016091f
C2230 FILLER_0_14_101/a_36_472# FILLER_0_13_72/a_3172_472# 0.026657f
C2231 FILLER_0_11_72/a_1468_375# _16_/I 0.007169f
C2232 _09_/ZN FILLER_0_4_107/a_124_375# 0.003315f
C2233 _14_/I FILLER_0_6_2/a_1020_375# 0.003099f
C2234 FILLER_0_6_2/a_2364_375# FILLER_0_7_2/a_2364_375# 0.05841f
C2235 FILLER_0_9_72/a_572_375# FILLER_0_8_37/a_4516_472# 0.001723f
C2236 FILLER_0_2_2/a_572_375# FILLER_0_4_2/a_484_472# 0.0027f
C2237 output_signal_minus[5] vdd 0.328106f
C2238 vdd FILLER_0_8_101/a_124_375# 0.043777f
C2239 output_signal_minus[9] FILLER_0_0_142/a_484_472# 0.001011f
C2240 FILLER_0_7_104/a_484_472# _03_/ZN 0.004342f
C2241 FILLER_0_9_72/a_2276_472# _14_/I 0.004017f
C2242 FILLER_0_12_12/a_1020_375# _17_/I 0.002388f
C2243 FILLER_0_11_72/a_1828_472# _16_/I 0.00753f
C2244 FILLER_0_6_37/a_932_472# FILLER_0_5_44/a_124_375# 0.001597f
C2245 _19_/I _10_/Z 0.04379f
C2246 _11_/I FILLER_0_2_37/a_5412_472# 0.002415f
C2247 FILLER_0_14_37/a_2276_472# _17_/I 0.015502f
C2248 _00_/ZN _17_/a_36_113# 0.139977f
C2249 FILLER_0_14_37/a_4964_472# _17_/I 0.015502f
C2250 _11_/I _13_/I 0.839309f
C2251 vdd FILLER_0_11_72/a_932_472# 0.004803f
C2252 _14_/I FILLER_0_9_2/a_2364_375# 0.005414f
C2253 FILLER_0_12_37/a_2724_472# vdd 0.008581f
C2254 _11_/I FILLER_0_8_107/a_484_472# 0.004233f
C2255 FILLER_0_12_107/a_36_472# FILLER_0_11_72/a_4068_472# 0.026657f
C2256 _07_/ZN output_signal_plus[1] 0.114015f
C2257 FILLER_0_4_2/a_1020_375# FILLER_0_3_12/a_36_472# 0.001543f
C2258 vdd FILLER_0_15_2/a_36_472# 0.10601f
C2259 FILLER_0_8_37/a_4068_472# FILLER_0_6_37/a_4156_375# 0.001512f
C2260 FILLER_0_13_104/a_36_472# FILLER_0_13_72/a_3260_375# 0.086742f
C2261 FILLER_0_2_37/a_1828_472# _10_/I 0.002525f
C2262 FILLER_0_8_37/a_5052_375# FILLER_0_9_72/a_1020_375# 0.026339f
C2263 FILLER_0_2_37/a_3172_472# vdd 0.008405f
C2264 FILLER_0_4_2/a_1468_375# _12_/I 0.003251f
C2265 _14_/I input_signal[4] 0.32954f
C2266 FILLER_0_15_8/a_2364_375# _18_/I 0.01418f
C2267 _16_/I output_signal_plus[2] 0.009099f
C2268 FILLER_0_13_72/a_2364_375# _16_/I 0.005093f
C2269 FILLER_0_5_12/a_484_472# vdd 0.0232f
C2270 _08_/ZN _06_/ZN 0.008635f
C2271 _13_/I FILLER_0_5_12/a_1828_472# 0.017477f
C2272 vdd FILLER_0_8_37/a_2812_375# 0.009158f
C2273 FILLER_0_9_2/a_6756_472# FILLER_0_8_37/a_2812_375# 0.001723f
C2274 output11/a_224_472# FILLER_0_1_72/a_1380_472# 0.005437f
C2275 FILLER_0_9_2/a_3260_375# vdd 0.020842f
C2276 _10_/a_36_160# _08_/ZN 0.001823f
C2277 output13/a_224_472# _13_/a_36_113# 0.020123f
C2278 _18_/I _10_/Z 0.06196f
C2279 _07_/ZN output_signal_minus[7] 0.020942f
C2280 FILLER_0_3_12/a_932_472# vdd 0.018883f
C2281 _17_/a_36_113# _17_/I 0.041373f
C2282 input10/a_36_113# input_signal[9] 0.052126f
C2283 FILLER_0_10_12/a_1020_375# _16_/I 0.002327f
C2284 FILLER_0_11_72/a_5948_375# vdd 0.022968f
C2285 FILLER_0_7_72/a_3172_472# _14_/I 0.010748f
C2286 FILLER_0_5_12/a_36_472# FILLER_0_6_2/a_1020_375# 0.001543f
C2287 output22/a_224_472# _10_/Z 0.029269f
C2288 FILLER_0_12_107/a_932_472# FILLER_0_11_72/a_4964_472# 0.026657f
C2289 vdd FILLER_0_2_37/a_5860_472# 0.006386f
C2290 FILLER_0_11_2/a_3172_472# FILLER_0_10_28/a_124_375# 0.001684f
C2291 FILLER_0_1_44/a_484_472# _10_/I 0.006408f
C2292 FILLER_0_10_12/a_1468_375# FILLER_0_10_28/a_36_472# 0.086635f
C2293 _19_/I input_signal[9] 0.339232f
C2294 FILLER_0_13_72/a_572_375# vdd 0.002455f
C2295 output17/a_224_472# output_signal_minus[5] 0.001272f
C2296 _19_/I FILLER_0_16_18/a_572_375# 0.01418f
C2297 _11_/I FILLER_0_3_60/a_36_472# 0.008683f
C2298 FILLER_0_1_60/a_124_375# FILLER_0_0_36/a_2812_375# 0.05841f
C2299 _11_/I FILLER_0_2_37/a_2364_375# 0.001984f
C2300 _18_/I FILLER_0_15_72/a_572_375# 0.01418f
C2301 FILLER_0_9_72/a_484_472# vdd 0.002467f
C2302 FILLER_0_8_37/a_484_472# _14_/I 0.014431f
C2303 FILLER_0_13_72/a_484_472# FILLER_0_15_72/a_572_375# 0.001512f
C2304 FILLER_0_12_107/a_572_375# FILLER_0_11_72/a_4516_472# 0.001597f
C2305 _08_/ZN output_signal_minus[3] 0.162335f
C2306 FILLER_0_12_37/a_124_375# FILLER_0_14_37/a_36_472# 0.001512f
C2307 _00_/ZN output_signal_minus[2] 0.043339f
C2308 FILLER_0_4_37/a_3708_375# vdd 0.021784f
C2309 FILLER_0_14_12/a_932_472# _16_/I 0.001653f
C2310 _15_/I FILLER_0_9_104/a_484_472# 0.006506f
C2311 FILLER_0_0_36/a_3260_375# _10_/I 0.015932f
C2312 FILLER_0_1_12/a_484_472# vdd 0.024695f
C2313 vdd FILLER_0_4_107/a_1468_375# 0.014222f
C2314 _14_/I FILLER_0_6_2/a_572_375# 0.003099f
C2315 vdd _03_/ZN 0.186524f
C2316 FILLER_0_13_2/a_1380_472# _16_/I 0.004669f
C2317 FILLER_0_9_2/a_1828_472# FILLER_0_8_12/a_572_375# 0.001684f
C2318 output_signal_plus[7] _16_/Z 0.006948f
C2319 _15_/Z output_signal_plus[6] 0.016592f
C2320 vdd FILLER_0_1_72/a_572_375# 0.00206f
C2321 FILLER_0_4_37/a_1380_472# FILLER_0_3_44/a_572_375# 0.001597f
C2322 _12_/I FILLER_0_5_72/a_124_375# 0.001706f
C2323 _10_/Z _10_/I 0.014664f
C2324 vdd FILLER_0_5_12/a_3260_375# 0.005051f
C2325 _14_/I FILLER_0_7_72/a_932_472# 0.008683f
C2326 FILLER_0_16_36/a_3172_472# FILLER_0_16_70/a_36_472# 0.003468f
C2327 FILLER_0_13_66/a_36_472# FILLER_0_14_37/a_3172_472# 0.026657f
C2328 _15_/I _12_/Z 0.15773f
C2329 _18_/I input_signal[9] 0.065423f
C2330 _18_/I FILLER_0_16_18/a_572_375# 0.001052f
C2331 _14_/Z output_signal_minus[2] 0.010158f
C2332 _18_/I FILLER_0_14_115/a_36_472# 0.004893f
C2333 vdd FILLER_0_15_72/a_484_472# 0.002143f
C2334 FILLER_0_12_107/a_36_472# _15_/I 0.001368f
C2335 FILLER_0_7_104/a_124_375# FILLER_0_7_72/a_3260_375# 0.012222f
C2336 FILLER_0_1_44/a_1468_375# _10_/I 0.001498f
C2337 _13_/I FILLER_0_6_37/a_4604_375# 0.001706f
C2338 FILLER_0_11_72/a_124_375# FILLER_0_10_37/a_4156_375# 0.026339f
C2339 _13_/I FILLER_0_6_37/a_1916_375# 0.001706f
C2340 FILLER_0_7_2/a_124_375# vdd -0.003842f
C2341 FILLER_0_14_101/a_36_472# _18_/I 0.001526f
C2342 _18_/I FILLER_0_15_72/a_124_375# 0.01418f
C2343 input8/a_36_113# FILLER_0_14_12/a_36_472# 0.001663f
C2344 FILLER_0_4_2/a_1020_375# _13_/I 0.005811f
C2345 FILLER_0_15_64/a_124_375# FILLER_0_15_72/a_124_375# 0.003732f
C2346 _14_/I net15 0.406952f
C2347 _15_/I FILLER_0_10_28/a_36_472# 0.015502f
C2348 _10_/I FILLER_0_1_12/a_572_375# 0.003137f
C2349 _09_/ZN _13_/a_36_113# 0.067564f
C2350 FILLER_0_11_2/a_36_472# FILLER_0_13_2/a_124_375# 0.00108f
C2351 FILLER_0_4_107/a_124_375# FILLER_0_4_101/a_124_375# 0.005439f
C2352 FILLER_0_1_44/a_932_472# FILLER_0_2_37/a_1828_472# 0.026657f
C2353 FILLER_0_3_12/a_2364_375# vdd 0.019634f
C2354 _18_/a_36_113# _10_/Z 0.007031f
C2355 _18_/I FILLER_0_14_37/a_5948_375# 0.003935f
C2356 _14_/I FILLER_0_8_12/a_1020_375# 0.01418f
C2357 FILLER_0_1_72/a_1468_375# output_signal_minus[9] 0.001027f
C2358 FILLER_0_5_44/a_932_472# vdd 0.009085f
C2359 FILLER_0_15_8/a_572_375# vdd -0.007105f
C2360 FILLER_0_12_37/a_1828_472# vdd 0.008978f
C2361 output_signal_minus[1] output_signal_plus[1] 0.176107f
C2362 _13_/I FILLER_0_4_2/a_3260_375# 0.00577f
C2363 FILLER_0_13_2/a_36_472# input_signal[7] 0.024466f
C2364 FILLER_0_13_2/a_6844_375# FILLER_0_11_2/a_6756_472# 0.001512f
C2365 _15_/I FILLER_0_9_72/a_932_472# 0.00652f
C2366 _11_/I FILLER_0_2_37/a_5948_375# 0.00346f
C2367 vdd FILLER_0_5_72/a_1916_375# 0.009315f
C2368 _14_/I FILLER_0_9_66/a_124_375# 0.005381f
C2369 FILLER_0_4_2/a_1916_375# vdd 0.050516f
C2370 vdd FILLER_0_6_37/a_36_472# 0.10831f
C2371 output13/a_224_472# _03_/ZN 0.038831f
C2372 FILLER_0_12_37/a_4964_472# FILLER_0_13_72/a_1020_375# 0.001723f
C2373 FILLER_0_0_12/a_572_375# _10_/I 0.016605f
C2374 _11_/I FILLER_0_3_12/a_572_375# 0.009462f
C2375 FILLER_0_4_2/a_124_375# input_signal[3] 0.040128f
C2376 _11_/I FILLER_0_3_104/a_484_472# 0.008683f
C2377 vdd _06_/ZN 0.305391f
C2378 _17_/I FILLER_0_14_37/a_484_472# 0.015502f
C2379 input7/a_36_113# input_signal[7] 0.002947f
C2380 _10_/a_36_160# vdd 0.03433f
C2381 FILLER_0_7_2/a_4068_472# _14_/I 0.003726f
C2382 _19_/I FILLER_0_16_18/a_124_375# 0.01418f
C2383 FILLER_0_13_72/a_1468_375# _16_/I 0.006182f
C2384 output19/a_224_472# output_signal_minus[8] 0.021278f
C2385 _11_/I output12/a_224_472# 0.003296f
C2386 FILLER_0_12_107/a_1380_472# FILLER_0_10_107/a_1468_375# 0.001512f
C2387 _14_/I FILLER_0_6_2/a_1468_375# 0.003099f
C2388 _16_/I FILLER_0_11_72/a_3260_375# 0.007169f
C2389 _16_/I FILLER_0_11_2/a_2724_472# 0.007596f
C2390 FILLER_0_2_37/a_572_375# vdd 0.007011f
C2391 FILLER_0_3_44/a_36_472# FILLER_0_3_12/a_3172_472# 0.013276f
C2392 vdd FILLER_0_13_2/a_4516_472# 0.006118f
C2393 vdd FILLER_0_2_37/a_4068_472# 0.00356f
C2394 _11_/I FILLER_0_4_37/a_2364_375# 0.01418f
C2395 FILLER_0_14_101/a_124_375# vdd 0.041136f
C2396 FILLER_0_13_2/a_6756_472# vdd 0.009694f
C2397 output_signal_plus[8] output29/a_224_472# 0.027343f
C2398 vdd FILLER_0_14_37/a_4068_472# 0.002855f
C2399 FILLER_0_2_37/a_124_375# vdd 0.014132f
C2400 _15_/I FILLER_0_12_37/a_5860_472# 0.001368f
C2401 _00_/ZN output11/a_224_472# 0.125198f
C2402 FILLER_0_3_72/a_484_472# vdd 0.002467f
C2403 FILLER_0_12_37/a_4068_472# FILLER_0_13_72/a_124_375# 0.001723f
C2404 _09_/ZN FILLER_0_11_72/a_5948_375# 0.012909f
C2405 FILLER_0_4_2/a_36_472# input_signal[2] 0.020769f
C2406 _15_/I FILLER_0_11_136/a_124_375# 0.001503f
C2407 FILLER_0_1_60/a_572_375# FILLER_0_1_72/a_124_375# 0.003732f
C2408 output_signal_minus[3] vdd 0.273026f
C2409 vdd FILLER_0_4_107/a_572_375# 0.016637f
C2410 FILLER_0_7_2/a_6756_472# vdd 0.008994f
C2411 FILLER_0_9_2/a_4964_472# FILLER_0_8_37/a_1020_375# 0.001723f
C2412 output18/a_224_472# output_signal_minus[6] 0.002784f
C2413 FILLER_0_5_44/a_1020_375# _12_/I 0.001706f
C2414 _13_/Z output_signal_minus[4] 0.005716f
C2415 _07_/ZN output_signal_plus[2] 0.098743f
C2416 _18_/I FILLER_0_16_18/a_124_375# 0.00145f
C2417 _17_/I FILLER_0_14_37/a_3620_472# 0.015502f
C2418 _00_/ZN output_signal_minus[8] 0.915677f
C2419 FILLER_0_7_72/a_2724_472# _12_/I 0.00187f
C2420 _14_/I FILLER_0_7_66/a_36_472# 0.008683f
C2421 _11_/I FILLER_0_4_37/a_4516_472# 0.014431f
C2422 _17_/I FILLER_0_15_72/a_36_472# 0.004125f
C2423 _14_/I FILLER_0_9_2/a_3620_472# 0.004017f
C2424 FILLER_0_15_40/a_1380_472# _19_/I 0.001782f
C2425 output19/a_224_472# FILLER_0_2_107/a_1468_375# 0.00135f
C2426 output_signal_plus[2] _11_/a_36_113# 0.023343f
C2427 FILLER_0_8_37/a_2364_375# FILLER_0_9_2/a_6308_472# 0.001723f
C2428 _13_/I _12_/a_36_113# 0.050349f
C2429 _09_/ZN _03_/ZN 0.109721f
C2430 _09_/ZN FILLER_0_4_107/a_1468_375# 0.023526f
C2431 FILLER_0_3_72/a_932_472# FILLER_0_5_72/a_1020_375# 0.001512f
C2432 _14_/I output_signal_minus[4] 0.049921f
C2433 _17_/I FILLER_0_14_37/a_6308_472# 0.015502f
C2434 FILLER_0_15_56/a_572_375# FILLER_0_14_37/a_2812_375# 0.026339f
C2435 FILLER_0_12_101/a_36_472# FILLER_0_11_72/a_3260_375# 0.001597f
C2436 FILLER_0_2_37/a_6756_472# output11/a_224_472# 0.031813f
C2437 FILLER_0_3_60/a_124_375# vdd 0.014636f
C2438 FILLER_0_10_37/a_2364_375# FILLER_0_11_2/a_6396_375# 0.026339f
C2439 FILLER_0_13_66/a_36_472# _16_/I 0.004669f
C2440 FILLER_0_9_2/a_1828_472# FILLER_0_11_2/a_1916_375# 0.0027f
C2441 vdd FILLER_0_4_37/a_3172_472# 0.007014f
C2442 _13_/I _12_/Z 0.031103f
C2443 FILLER_0_5_12/a_2364_375# _12_/I 0.001706f
C2444 FILLER_0_13_72/a_3172_472# _17_/I 0.00652f
C2445 _16_/I FILLER_0_12_37/a_6756_472# 0.017477f
C2446 FILLER_0_1_72/a_1380_472# _10_/I 0.006408f
C2447 FILLER_0_5_44/a_1380_472# vdd 0.040664f
C2448 FILLER_0_12_37/a_1916_375# vdd 0.015021f
C2449 FILLER_0_12_12/a_1468_375# vdd 0.024432f
C2450 FILLER_0_6_37/a_1468_375# FILLER_0_8_37/a_1380_472# 0.001512f
C2451 FILLER_0_4_37/a_6844_375# FILLER_0_4_101/a_124_375# 0.012001f
C2452 FILLER_0_6_37/a_124_375# _12_/I 0.016315f
C2453 FILLER_0_16_18/a_1020_375# FILLER_0_15_8/a_2276_472# 0.001543f
C2454 FILLER_0_5_104/a_124_375# FILLER_0_3_104/a_36_472# 0.0027f
C2455 FILLER_0_15_40/a_1380_472# _18_/I 0.014431f
C2456 FILLER_0_13_104/a_36_472# _18_/Z 0.001538f
C2457 FILLER_0_8_12/a_124_375# FILLER_0_9_2/a_1380_472# 0.001684f
C2458 _17_/I input_signal[7] 0.353802f
C2459 FILLER_0_12_12/a_36_472# input7/a_36_113# 0.001663f
C2460 input_signal[7] FILLER_0_15_8/a_124_375# 0.002912f
C2461 FILLER_0_11_72/a_2364_375# _16_/I 0.007169f
C2462 FILLER_0_15_56/a_36_472# FILLER_0_15_40/a_1468_375# 0.086743f
C2463 vdd FILLER_0_9_2/a_5412_472# 0.008843f
C2464 FILLER_0_11_72/a_4604_375# _15_/I 0.007111f
C2465 FILLER_0_16_70/a_124_375# output_signal_plus[9] 0.011852f
C2466 vdd FILLER_0_15_8/a_2812_375# 0.018843f
C2467 FILLER_0_10_12/a_1020_375# FILLER_0_11_2/a_2276_472# 0.001684f
C2468 FILLER_0_14_12/a_484_472# FILLER_0_12_12/a_572_375# 0.0027f
C2469 vdd FILLER_0_3_12/a_1468_375# 0.023663f
C2470 FILLER_0_4_2/a_2364_375# _11_/I 0.01418f
C2471 vdd FILLER_0_15_40/a_1468_375# 0.012652f
C2472 FILLER_0_1_60/a_484_472# FILLER_0_1_72/a_36_472# 0.002296f
C2473 FILLER_0_13_72/a_1916_375# FILLER_0_12_37/a_5860_472# 0.001723f
C2474 FILLER_0_5_12/a_484_472# input_signal[3] 0.001168f
C2475 _15_/I FILLER_0_10_37/a_484_472# 0.015502f
C2476 vdd FILLER_0_2_37/a_36_472# 0.109127f
C2477 _15_/I FILLER_0_9_72/a_2724_472# 0.00652f
C2478 _15_/I FILLER_0_9_2/a_6308_472# 0.006506f
C2479 FILLER_0_10_12/a_932_472# vdd 0.017846f
C2480 FILLER_0_3_60/a_484_472# vdd 0.013043f
C2481 vdd FILLER_0_2_107/a_124_375# 0.01497f
C2482 FILLER_0_7_2/a_484_472# FILLER_0_9_2/a_572_375# 0.0027f
C2483 FILLER_0_12_107/a_1380_472# _16_/I 0.017919f
C2484 FILLER_0_6_37/a_6396_375# FILLER_0_7_72/a_2364_375# 0.026339f
C2485 _16_/I FILLER_0_14_37/a_2724_472# 0.001667f
C2486 FILLER_0_3_44/a_124_375# vdd 0.011034f
C2487 FILLER_0_16_104/a_124_375# output21/a_224_472# 0.01196f
C2488 vdd FILLER_0_3_72/a_3172_472# 0.009151f
C2489 FILLER_0_5_12/a_2812_375# FILLER_0_6_37/a_36_472# 0.001597f
C2490 FILLER_0_8_107/a_124_375# FILLER_0_9_104/a_572_375# 0.026339f
C2491 _00_/ZN _19_/I 0.049372f
C2492 vdd FILLER_0_13_2/a_5412_472# 0.009543f
C2493 _17_/Z _16_/I 0.02009f
C2494 FILLER_0_7_72/a_1468_375# _14_/I 0.008393f
C2495 FILLER_0_11_2/a_5412_472# vdd 0.008843f
C2496 FILLER_0_2_2/a_572_375# _11_/I 0.04168f
C2497 FILLER_0_13_104/a_484_472# _18_/Z 0.001466f
C2498 FILLER_0_14_12/a_484_472# _17_/I 0.015594f
C2499 vdd FILLER_0_7_72/a_2812_375# 0.019859f
C2500 vdd FILLER_0_2_107/a_36_472# 0.108263f
C2501 _17_/I FILLER_0_13_2/a_6396_375# 0.006125f
C2502 _15_/I FILLER_0_11_72/a_572_375# 0.007126f
C2503 FILLER_0_6_37/a_4964_472# vdd 0.005073f
C2504 FILLER_0_15_72/a_1468_375# vdd 0.015779f
C2505 FILLER_0_12_37/a_6756_472# FILLER_0_13_72/a_2812_375# 0.001723f
C2506 FILLER_0_1_44/a_1380_472# FILLER_0_2_37/a_2276_472# 0.026657f
C2507 _16_/I FILLER_0_11_72/a_484_472# 0.001852f
C2508 FILLER_0_1_72/a_1468_375# output20/a_224_472# 0.03228f
C2509 FILLER_0_12_101/a_36_472# FILLER_0_12_37/a_6756_472# 0.013277f
C2510 _14_/I FILLER_0_8_37/a_6756_472# 0.014868f
C2511 _19_/Z output29/a_224_472# 0.148069f
C2512 FILLER_0_13_2/a_5860_472# FILLER_0_12_37/a_1916_375# 0.001723f
C2513 FILLER_0_8_28/a_124_375# vdd 0.046575f
C2514 vdd FILLER_0_8_37/a_3260_375# 0.007055f
C2515 FILLER_0_14_37/a_6756_472# FILLER_0_13_72/a_2724_472# 0.026657f
C2516 _13_/I FILLER_0_4_107/a_1380_472# 0.001318f
C2517 output_signal_minus[1] output_signal_plus[2] 0.006826f
C2518 _17_/I _19_/I 0.054381f
C2519 _09_/ZN FILLER_0_4_107/a_572_375# 0.007439f
C2520 _19_/I FILLER_0_15_8/a_124_375# 0.008393f
C2521 FILLER_0_0_36/a_3260_375# FILLER_0_0_70/a_36_472# 0.016748f
C2522 _15_/I FILLER_0_8_37/a_572_375# 0.002388f
C2523 _13_/I output_signal_minus[6] 0.060548f
C2524 FILLER_0_4_37/a_6756_472# FILLER_0_5_72/a_2812_375# 0.001723f
C2525 FILLER_0_14_37/a_932_472# FILLER_0_15_40/a_572_375# 0.001723f
C2526 output30/a_224_472# FILLER_0_15_72/a_484_472# 0.035046f
C2527 FILLER_0_4_37/a_4068_472# FILLER_0_2_37/a_4156_375# 0.001512f
C2528 vdd FILLER_0_9_2/a_572_375# 0.019913f
C2529 FILLER_0_7_2/a_124_375# input_signal[3] 0.001163f
C2530 vdd FILLER_0_4_107/a_1020_375# 0.001984f
C2531 FILLER_0_7_2/a_2724_472# _12_/I 0.004669f
C2532 FILLER_0_7_66/a_124_375# FILLER_0_7_2/a_6844_375# 0.012001f
C2533 FILLER_0_13_2/a_4156_375# _17_/I 0.004676f
C2534 FILLER_0_12_37/a_4156_375# FILLER_0_13_72/a_124_375# 0.026339f
C2535 _17_/I FILLER_0_15_8/a_484_472# 0.004125f
C2536 _11_/I FILLER_0_4_2/a_932_472# 0.016612f
C2537 _10_/Z FILLER_0_11_72/a_5860_472# 0.008573f
C2538 FILLER_0_2_37/a_2724_472# vdd 0.01103f
C2539 FILLER_0_4_2/a_36_472# FILLER_0_2_2/a_124_375# 0.00108f
C2540 FILLER_0_6_37/a_6844_375# FILLER_0_7_72/a_2812_375# 0.026339f
C2541 _13_/Z _10_/Z 0.521439f
C2542 FILLER_0_7_72/a_124_375# _12_/I 0.006182f
C2543 output_signal_plus[4] _16_/a_36_113# 0.001039f
C2544 _07_/ZN _11_/I 0.037277f
C2545 FILLER_0_4_2/a_1916_375# FILLER_0_5_12/a_932_472# 0.001684f
C2546 _17_/I _18_/I 0.867795f
C2547 _18_/I FILLER_0_15_8/a_124_375# 0.0037f
C2548 _17_/I FILLER_0_13_72/a_484_472# 0.001644f
C2549 FILLER_0_15_64/a_124_375# _17_/I 0.006589f
C2550 _15_/I FILLER_0_11_2/a_4156_375# 0.007111f
C2551 FILLER_0_14_37/a_1916_375# vdd 0.01595f
C2552 vdd FILLER_0_11_2/a_572_375# 0.02016f
C2553 FILLER_0_14_37/a_1020_375# FILLER_0_15_40/a_572_375# 0.026339f
C2554 vdd FILLER_0_3_72/a_1468_375# 0.007205f
C2555 _13_/I FILLER_0_6_37/a_1020_375# 0.001706f
C2556 _11_/I FILLER_0_3_44/a_36_472# 0.008683f
C2557 _11_/I _11_/a_36_113# 0.016972f
C2558 FILLER_0_2_37/a_3172_472# FILLER_0_1_60/a_572_375# 0.001597f
C2559 FILLER_0_12_12/a_124_375# vdd 0.033413f
C2560 _00_/ZN _10_/I 2.433093f
C2561 _13_/I FILLER_0_6_37/a_932_472# 0.003818f
C2562 FILLER_0_7_2/a_36_472# FILLER_0_9_2/a_124_375# 0.00108f
C2563 _14_/I FILLER_0_7_2/a_6396_375# 0.008393f
C2564 vdd FILLER_0_11_2/a_2812_375# 0.022556f
C2565 output12/a_224_472# _12_/Z 0.11967f
C2566 _02_/ZN _14_/I 0.076469f
C2567 output_signal_plus[7] output28/a_224_472# 0.053836f
C2568 _16_/I FILLER_0_11_72/a_6756_472# 0.006872f
C2569 _14_/I _10_/Z 0.155363f
C2570 vdd FILLER_0_1_44/a_572_375# -0.008493f
C2571 _17_/I FILLER_0_14_12/a_1468_375# 0.018729f
C2572 output_signal_minus[5] output_signal_minus[8] 0.021693f
C2573 FILLER_0_16_70/a_36_472# output_signal_plus[9] 0.002187f
C2574 vdd FILLER_0_11_72/a_1380_472# 0.006325f
C2575 FILLER_0_10_12/a_36_472# FILLER_0_9_2/a_1020_375# 0.001543f
C2576 input_signal[6] input6/a_36_113# 0.004439f
C2577 vdd FILLER_0_2_37/a_5052_375# 0.007501f
C2578 FILLER_0_5_12/a_484_472# FILLER_0_4_2/a_1468_375# 0.001684f
C2579 FILLER_0_3_60/a_124_375# FILLER_0_3_44/a_1468_375# 0.012222f
C2580 FILLER_0_3_72/a_124_375# vdd 0.013594f
C2581 _13_/I FILLER_0_5_12/a_2724_472# 0.017477f
C2582 FILLER_0_6_37/a_5948_375# _12_/I 0.016091f
C2583 FILLER_0_13_104/a_484_472# FILLER_0_12_107/a_124_375# 0.001723f
C2584 FILLER_0_12_37/a_4516_472# FILLER_0_11_72/a_484_472# 0.026657f
C2585 FILLER_0_8_37/a_4964_472# FILLER_0_9_72/a_1020_375# 0.001723f
C2586 FILLER_0_3_44/a_124_375# FILLER_0_4_37/a_932_472# 0.001597f
C2587 FILLER_0_1_72/a_124_375# _10_/I 0.008292f
C2588 FILLER_0_7_72/a_1468_375# FILLER_0_8_37/a_5412_472# 0.001597f
C2589 FILLER_0_11_72/a_6844_375# _08_/ZN 0.009573f
C2590 _11_/I FILLER_0_3_12/a_484_472# 0.010838f
C2591 input_signal[7] FILLER_0_15_2/a_36_472# 0.004572f
C2592 _11_/I FILLER_0_4_37/a_4068_472# 0.014431f
C2593 _11_/I FILLER_0_5_72/a_484_472# 0.001913f
C2594 FILLER_0_7_2/a_36_472# vdd 0.105401f
C2595 output_signal_minus[2] _06_/ZN 0.047281f
C2596 input_signal[0] input1/a_36_113# 0.023145f
C2597 FILLER_0_12_107/a_36_472# _16_/I 0.018669f
C2598 _17_/I FILLER_0_13_72/a_124_375# 0.006125f
C2599 FILLER_0_9_2/a_932_472# FILLER_0_11_2/a_1020_375# 0.0027f
C2600 FILLER_0_0_12/a_36_472# vdd 0.010651f
C2601 FILLER_0_6_2/a_2812_375# FILLER_0_7_2/a_2812_375# 0.05841f
C2602 FILLER_0_2_37/a_6756_472# _10_/I 0.002386f
C2603 vdd FILLER_0_7_2/a_3260_375# -0.011271f
C2604 FILLER_0_10_107/a_1020_375# _15_/I 0.018729f
C2605 FILLER_0_2_37/a_5500_375# FILLER_0_3_72/a_1468_375# 0.026339f
C2606 FILLER_0_10_107/a_572_375# vdd 0.002455f
C2607 FILLER_0_6_107/a_124_375# FILLER_0_5_104/a_484_472# 0.001597f
C2608 output11/a_224_472# FILLER_0_2_37/a_5860_472# 0.031509f
C2609 vdd FILLER_0_5_72/a_2364_375# 0.021274f
C2610 FILLER_0_8_37/a_1916_375# FILLER_0_9_2/a_5860_472# 0.001723f
C2611 FILLER_0_5_12/a_1468_375# FILLER_0_3_12/a_1380_472# 0.0027f
C2612 _15_/I FILLER_0_11_72/a_5500_375# 0.005506f
C2613 FILLER_0_8_37/a_1468_375# _14_/I 0.01418f
C2614 vdd FILLER_0_11_2/a_1380_472# 0.012473f
C2615 _11_/I FILLER_0_2_107/a_484_472# 0.002415f
C2616 _14_/I FILLER_0_9_72/a_1828_472# 0.004017f
C2617 FILLER_0_13_2/a_5860_472# FILLER_0_14_37/a_1916_375# 0.001597f
C2618 _14_/I FILLER_0_7_2/a_5052_375# 0.008393f
C2619 FILLER_0_8_37/a_6308_472# _14_/I 0.014431f
C2620 output_signal_plus[7] FILLER_0_13_104/a_484_472# 0.002187f
C2621 vdd FILLER_0_12_37/a_2276_472# 0.035321f
C2622 FILLER_0_2_37/a_4516_472# FILLER_0_1_72/a_572_375# 0.001597f
C2623 _14_/Z _16_/a_36_113# 0.020822f
C2624 _11_/I FILLER_0_4_2/a_2724_472# 0.014431f
C2625 output_signal_minus[2] output_signal_minus[3] 0.140198f
C2626 FILLER_0_10_107/a_124_375# FILLER_0_10_101/a_124_375# 0.005439f
C2627 FILLER_0_7_104/a_36_472# vdd 0.093924f
C2628 _17_/I _16_/a_36_113# 0.001886f
C2629 FILLER_0_9_72/a_2364_375# FILLER_0_8_37/a_6396_375# 0.026339f
C2630 FILLER_0_7_72/a_572_375# FILLER_0_6_37/a_4516_472# 0.001723f
C2631 FILLER_0_10_107/a_36_472# FILLER_0_9_104/a_484_472# 0.026657f
C2632 FILLER_0_6_37/a_1828_472# vdd 0.009247f
C2633 FILLER_0_3_12/a_1916_375# vdd 0.021609f
C2634 FILLER_0_10_107/a_932_472# _09_/ZN 0.006746f
C2635 FILLER_0_9_2/a_4156_375# vdd 0.004039f
C2636 FILLER_0_1_12/a_36_472# vdd 0.015685f
C2637 _09_/ZN FILLER_0_4_107/a_1020_375# 0.030288f
C2638 _17_/I FILLER_0_13_2/a_5948_375# 0.006125f
C2639 _17_/Z output27/a_224_472# 0.051576f
C2640 _15_/I FILLER_0_9_72/a_2276_472# 0.00652f
C2641 FILLER_0_13_2/a_4516_472# FILLER_0_14_37/a_484_472# 0.026657f
C2642 FILLER_0_0_142/a_572_375# vdd 0.039381f
C2643 _11_/I FILLER_0_5_72/a_932_472# 0.001913f
C2644 output_signal_minus[1] _11_/I 0.00156f
C2645 vdd FILLER_0_11_72/a_4516_472# 0.003435f
C2646 _15_/I FILLER_0_10_37/a_5412_472# 0.015502f
C2647 FILLER_0_12_107/a_36_472# FILLER_0_12_101/a_36_472# 0.003468f
C2648 _13_/Z _12_/I 0.055269f
C2649 FILLER_0_6_37/a_3172_472# FILLER_0_5_60/a_572_375# 0.001597f
C2650 FILLER_0_7_2/a_1020_375# FILLER_0_8_12/a_36_472# 0.001543f
C2651 _15_/I FILLER_0_9_2/a_2364_375# 0.006125f
C2652 output15/a_224_472# _13_/Z 0.00998f
C2653 _16_/I FILLER_0_12_37/a_5860_472# 0.017477f
C2654 _17_/Z output_signal_plus[5] 0.145667f
C2655 input_signal[6] FILLER_0_11_2/a_932_472# 0.002507f
C2656 _15_/I FILLER_0_11_72/a_6308_472# 0.004676f
C2657 _15_/a_36_113# _15_/Z 0.002665f
C2658 _16_/I FILLER_0_11_136/a_124_375# 0.007308f
C2659 output24/a_224_472# _08_/ZN 0.083176f
C2660 vdd FILLER_0_2_2/a_932_472# 0.010864f
C2661 output25/a_224_472# FILLER_0_11_136/a_36_472# 0.038484f
C2662 FILLER_0_6_2/a_36_472# input_signal[4] 0.00404f
C2663 vdd FILLER_0_0_104/a_124_375# 0.028958f
C2664 FILLER_0_3_12/a_1020_375# vdd 0.026369f
C2665 vdd FILLER_0_3_12/a_1380_472# 0.01093f
C2666 FILLER_0_10_107/a_124_375# vdd 0.014533f
C2667 _17_/I FILLER_0_13_72/a_1020_375# 0.006125f
C2668 FILLER_0_11_72/a_6844_375# vdd 0.043757f
C2669 _14_/I _12_/I 1.049906f
C2670 _16_/I output26/a_224_472# 0.006813f
C2671 FILLER_0_8_107/a_36_472# FILLER_0_8_101/a_36_472# 0.003468f
C2672 FILLER_0_8_107/a_124_375# _14_/I 0.015759f
C2673 vdd _14_/a_36_113# 0.016371f
C2674 output_signal_plus[7] FILLER_0_12_107/a_1020_375# 0.001313f
C2675 FILLER_0_12_107/a_572_375# vdd 0.015888f
C2676 vdd FILLER_0_16_18/a_1468_375# 0.032537f
C2677 FILLER_0_3_72/a_1916_375# _11_/I 0.008393f
C2678 FILLER_0_5_104/a_36_472# FILLER_0_5_72/a_3260_375# 0.086742f
C2679 FILLER_0_7_72/a_36_472# FILLER_0_7_66/a_36_472# 0.003468f
C2680 FILLER_0_13_66/a_124_375# FILLER_0_13_72/a_36_472# 0.016748f
C2681 FILLER_0_9_72/a_2364_375# FILLER_0_7_72/a_2276_472# 0.001512f
C2682 FILLER_0_1_44/a_1020_375# _10_/I 0.008103f
C2683 FILLER_0_5_44/a_1380_472# FILLER_0_6_37/a_2276_472# 0.026657f
C2684 _13_/I FILLER_0_5_104/a_572_375# 0.02241f
C2685 FILLER_0_7_2/a_4604_375# _14_/I 0.008393f
C2686 _10_/Z output16/a_224_472# 0.068033f
C2687 FILLER_0_15_8/a_3172_472# _17_/I 0.004125f
C2688 FILLER_0_8_37/a_5948_375# FILLER_0_9_72/a_1916_375# 0.026339f
C2689 FILLER_0_6_37/a_5948_375# FILLER_0_7_72/a_1916_375# 0.026339f
C2690 FILLER_0_12_37/a_5500_375# _17_/I 0.002388f
C2691 _16_/I FILLER_0_12_37/a_6308_472# 0.017477f
C2692 FILLER_0_7_2/a_932_472# vdd 0.009688f
C2693 FILLER_0_6_37/a_5412_472# FILLER_0_5_72/a_1380_472# 0.026657f
C2694 FILLER_0_8_37/a_6844_375# FILLER_0_8_101/a_36_472# 0.086635f
C2695 FILLER_0_3_44/a_124_375# FILLER_0_2_37/a_1020_375# 0.026339f
C2696 FILLER_0_9_72/a_36_472# _14_/I 0.004017f
C2697 input_signal[5] FILLER_0_9_2/a_572_375# 0.017676f
C2698 _07_/ZN FILLER_0_11_72/a_6756_472# 0.023101f
C2699 FILLER_0_2_37/a_4604_375# vdd 0.004128f
C2700 _15_/I FILLER_0_10_12/a_484_472# 0.016023f
C2701 _13_/I FILLER_0_6_2/a_3260_375# 0.001706f
C2702 _11_/I FILLER_0_2_2/a_1468_375# 0.007381f
C2703 FILLER_0_11_72/a_4604_375# _16_/I 0.002848f
C2704 FILLER_0_10_101/a_36_472# FILLER_0_10_37/a_6844_375# 0.086635f
C2705 FILLER_0_6_2/a_1380_472# _12_/I 0.019649f
C2706 _09_/ZN FILLER_0_10_107/a_572_375# 0.003962f
C2707 FILLER_0_1_44/a_1380_472# vdd 0.043943f
C2708 vdd FILLER_0_5_72/a_1380_472# 0.005631f
C2709 FILLER_0_8_37/a_36_472# vdd 0.108844f
C2710 FILLER_0_7_2/a_4964_472# vdd 0.006804f
C2711 _13_/I FILLER_0_4_37/a_3260_375# 0.005726f
C2712 _17_/I FILLER_0_14_12/a_124_375# 0.019386f
C2713 _16_/I FILLER_0_14_37/a_4516_472# 0.001424f
C2714 FILLER_0_13_66/a_36_472# FILLER_0_13_2/a_6844_375# 0.086635f
C2715 FILLER_0_13_2/a_572_375# _16_/I 0.006828f
C2716 output22/a_224_472# FILLER_0_11_72/a_5948_375# 0.002409f
C2717 input2/a_36_113# FILLER_0_1_12/a_36_472# 0.001663f
C2718 _15_/a_36_113# output_signal_plus[1] 0.021353f
C2719 _11_/I FILLER_0_2_2/a_484_472# 0.05086f
C2720 FILLER_0_5_12/a_36_472# _12_/I 0.009334f
C2721 output13/a_224_472# _14_/a_36_113# 0.004186f
C2722 FILLER_0_6_37/a_6756_472# _12_/I 0.017477f
C2723 FILLER_0_11_72/a_6396_375# _08_/ZN 0.001164f
C2724 FILLER_0_6_2/a_2724_472# _12_/I 0.017477f
C2725 _13_/I FILLER_0_0_142/a_484_472# 0.001188f
C2726 FILLER_0_8_37/a_124_375# _14_/I 0.01418f
C2727 FILLER_0_5_44/a_572_375# vdd 0.008383f
C2728 FILLER_0_11_2/a_2812_375# FILLER_0_9_2/a_2724_472# 0.0027f
C2729 FILLER_0_2_37/a_3172_472# _10_/I 0.002525f
C2730 vdd FILLER_0_5_72/a_2724_472# 0.030585f
C2731 input_signal[6] FILLER_0_12_12/a_484_472# 0.001912f
C2732 FILLER_0_9_72/a_124_375# _14_/I 0.005381f
C2733 _13_/I FILLER_0_6_2/a_1020_375# 0.001706f
C2734 _16_/I FILLER_0_11_72/a_572_375# 0.004231f
C2735 FILLER_0_9_104/a_36_472# _14_/I 0.004017f
C2736 vdd FILLER_0_16_36/a_572_375# 0.00158f
C2737 FILLER_0_5_44/a_36_472# vdd 0.090189f
C2738 FILLER_0_12_12/a_932_472# FILLER_0_10_12/a_1020_375# 0.0027f
C2739 FILLER_0_9_2/a_5948_375# vdd 0.032271f
C2740 FILLER_0_0_142/a_124_375# vdd 0.009175f
C2741 FILLER_0_6_37/a_2812_375# _12_/I 0.016091f
C2742 output24/a_224_472# vdd 0.165069f
C2743 _15_/I FILLER_0_11_72/a_4156_375# 0.007111f
C2744 _15_/I FILLER_0_8_12/a_1020_375# 0.002388f
C2745 _13_/I FILLER_0_6_2/a_1916_375# 0.001706f
C2746 _17_/Z output_signal_plus[6] 0.16562f
C2747 _09_/ZN FILLER_0_11_72/a_4516_472# 0.003603f
C2748 _11_/I FILLER_0_5_60/a_484_472# 0.001913f
C2749 FILLER_0_8_37/a_6844_375# FILLER_0_10_37/a_6756_472# 0.001512f
C2750 FILLER_0_7_2/a_1468_375# FILLER_0_8_12/a_484_472# 0.001543f
C2751 _15_/I FILLER_0_9_66/a_124_375# 0.006125f
C2752 output19/a_224_472# _14_/I 0.128014f
C2753 FILLER_0_6_107/a_124_375# _12_/I 0.019881f
C2754 _11_/I FILLER_0_4_37/a_6756_472# 0.014431f
C2755 FILLER_0_4_2/a_484_472# input_signal[2] 0.001108f
C2756 _18_/I FILLER_0_15_72/a_484_472# 0.014431f
C2757 FILLER_0_16_104/a_124_375# _18_/Z 0.001719f
C2758 FILLER_0_2_37/a_5860_472# _10_/I 0.002486f
C2759 FILLER_0_13_104/a_124_375# _17_/I 0.006125f
C2760 vdd FILLER_0_14_37/a_1828_472# 0.010403f
C2761 FILLER_0_2_107/a_932_472# output_signal_minus[6] 0.001473f
C2762 _11_/I FILLER_0_4_37/a_36_472# 0.014431f
C2763 _11_/I _04_/ZN 0.120439f
C2764 FILLER_0_10_107/a_1468_375# FILLER_0_11_72/a_5500_375# 0.026339f
C2765 FILLER_0_8_107/a_572_375# _11_/I 0.02657f
C2766 FILLER_0_3_72/a_1380_472# FILLER_0_4_37/a_5412_472# 0.026657f
C2767 FILLER_0_8_37/a_5860_472# FILLER_0_7_72/a_1916_375# 0.001597f
C2768 input_signal[4] input5/a_36_113# 0.028434f
C2769 FILLER_0_13_2/a_4964_472# vdd 0.007504f
C2770 FILLER_0_15_64/a_36_472# _17_/I 0.004125f
C2771 FILLER_0_10_107/a_124_375# _09_/ZN 0.002085f
C2772 vdd FILLER_0_8_37/a_5500_375# 0.009007f
C2773 _11_/I FILLER_0_2_37/a_3708_375# 0.00346f
C2774 FILLER_0_2_37/a_3260_375# FILLER_0_4_37/a_3172_472# 0.001512f
C2775 FILLER_0_6_37/a_2364_375# FILLER_0_7_2/a_6396_375# 0.026339f
C2776 vdd FILLER_0_6_101/a_124_375# 0.043907f
C2777 _11_/I FILLER_0_2_37/a_1380_472# 0.002415f
C2778 FILLER_0_9_2/a_484_472# input_signal[4] 0.003497f
C2779 FILLER_0_15_8/a_572_375# _18_/I 0.015448f
C2780 vdd FILLER_0_12_37/a_5052_375# 0.007396f
C2781 FILLER_0_10_101/a_36_472# FILLER_0_8_101/a_124_375# 0.001512f
C2782 FILLER_0_11_72/a_2276_472# vdd 0.011667f
C2783 FILLER_0_1_12/a_484_472# _10_/I 0.004764f
C2784 FILLER_0_12_107/a_572_375# _09_/ZN 0.003962f
C2785 FILLER_0_1_12/a_36_472# input_signal[1] 0.071895f
C2786 _14_/I FILLER_0_7_72/a_1916_375# 0.008393f
C2787 _07_/ZN FILLER_0_11_136/a_124_375# 0.030177f
C2788 _14_/I FILLER_0_8_37/a_1020_375# 0.01418f
C2789 _00_/ZN _14_/I 0.022453f
C2790 vdd FILLER_0_2_37/a_2276_472# 0.04006f
C2791 FILLER_0_5_12/a_572_375# FILLER_0_4_2/a_1828_472# 0.001684f
C2792 FILLER_0_1_72/a_572_375# _10_/I 0.008197f
C2793 vdd FILLER_0_10_37/a_932_472# 0.006024f
C2794 vdd FILLER_0_11_2/a_5860_472# 0.017111f
C2795 vdd FILLER_0_9_2/a_4068_472# 0.002735f
C2796 FILLER_0_9_2/a_4516_472# FILLER_0_10_37/a_484_472# 0.026657f
C2797 _11_/I FILLER_0_4_37/a_5412_472# 0.014431f
C2798 FILLER_0_5_104/a_572_375# FILLER_0_3_104/a_484_472# 0.001512f
C2799 output_signal_plus[0] _10_/Z 0.00741f
C2800 FILLER_0_1_72/a_484_472# FILLER_0_3_72/a_572_375# 0.001512f
C2801 _16_/I FILLER_0_11_2/a_4156_375# 0.005501f
C2802 output_signal_minus[9] _00_/ZN 0.136507f
C2803 _07_/ZN output_signal_minus[6] 0.049342f
C2804 FILLER_0_6_2/a_2812_375# FILLER_0_5_12/a_1828_472# 0.001543f
C2805 FILLER_0_10_28/a_36_472# FILLER_0_10_37/a_36_472# 0.001963f
C2806 FILLER_0_15_56/a_124_375# FILLER_0_15_40/a_1468_375# 0.012222f
C2807 FILLER_0_11_72/a_932_472# FILLER_0_13_72/a_1020_375# 0.001512f
C2808 _15_/I FILLER_0_9_2/a_3620_472# 0.006613f
C2809 FILLER_0_2_107/a_36_472# output_signal_minus[8] 0.001447f
C2810 FILLER_0_9_72/a_1468_375# FILLER_0_8_37/a_5500_375# 0.026339f
C2811 FILLER_0_12_107/a_1468_375# output_signal_plus[4] 0.010183f
C2812 FILLER_0_2_2/a_3260_375# FILLER_0_4_2/a_3172_472# 0.0027f
C2813 FILLER_0_4_2/a_2276_472# FILLER_0_5_12/a_1020_375# 0.001684f
C2814 FILLER_0_14_101/a_124_375# _18_/I 0.003935f
C2815 FILLER_0_14_107/a_124_375# FILLER_0_13_104/a_484_472# 0.001597f
C2816 input_signal[6] FILLER_0_11_2/a_124_375# 0.010061f
C2817 _15_/I FILLER_0_11_2/a_6308_472# 0.003016f
C2818 _18_/I FILLER_0_14_37/a_4068_472# 0.001526f
C2819 _14_/Z _14_/I 0.017631f
C2820 FILLER_0_8_12/a_1468_375# FILLER_0_8_28/a_36_472# 0.086635f
C2821 FILLER_0_2_107/a_1380_472# vdd 0.003184f
C2822 _13_/I FILLER_0_6_2/a_572_375# 0.001839f
C2823 FILLER_0_11_72/a_6396_375# vdd 0.008108f
C2824 vdd FILLER_0_15_8/a_932_472# 0.022599f
C2825 FILLER_0_13_2/a_5860_472# FILLER_0_14_37/a_1828_472# 0.026657f
C2826 FILLER_0_1_72/a_1380_472# output20/a_224_472# 0.001699f
C2827 _11_/I FILLER_0_2_37/a_4964_472# 0.002415f
C2828 FILLER_0_3_72/a_1020_375# FILLER_0_2_37/a_4964_472# 0.001723f
C2829 FILLER_0_4_37/a_5948_375# FILLER_0_5_72/a_1916_375# 0.026339f
C2830 output_signal_minus[1] _12_/Z 0.156466f
C2831 output_signal_plus[8] _10_/Z 0.008894f
C2832 FILLER_0_3_60/a_124_375# FILLER_0_4_37/a_2724_472# 0.001597f
C2833 _19_/a_36_113# vdd 0.060195f
C2834 FILLER_0_11_72/a_572_375# FILLER_0_12_37/a_4516_472# 0.001597f
C2835 _11_/I FILLER_0_5_104/a_124_375# 0.004764f
C2836 FILLER_0_6_37/a_6844_375# FILLER_0_6_101/a_124_375# 0.012001f
C2837 FILLER_0_6_2/a_2276_472# FILLER_0_5_12/a_1020_375# 0.001543f
C2838 output27/a_224_472# output26/a_224_472# 0.061459f
C2839 output23/a_224_472# _10_/Z 0.061631f
C2840 FILLER_0_9_2/a_5052_375# FILLER_0_7_2/a_4964_472# 0.001512f
C2841 _06_/ZN _10_/I 0.011118f
C2842 _15_/I FILLER_0_10_37/a_4516_472# 0.015502f
C2843 FILLER_0_1_72/a_1468_375# FILLER_0_2_37/a_5412_472# 0.001597f
C2844 _15_/I FILLER_0_10_37/a_5860_472# 0.015502f
C2845 FILLER_0_0_142/a_36_472# vdd 0.090744f
C2846 FILLER_0_2_107/a_1020_375# output19/a_224_472# 0.001274f
C2847 FILLER_0_16_36/a_124_375# FILLER_0_16_18/a_1468_375# 0.005439f
C2848 FILLER_0_13_2/a_2812_375# FILLER_0_11_2/a_2724_472# 0.0027f
C2849 FILLER_0_7_2/a_1380_472# input_signal[4] 0.001545f
C2850 _10_/a_36_160# _10_/I 0.04652f
C2851 _13_/I net15 0.02696f
C2852 output_signal_plus[5] output26/a_224_472# 0.03317f
C2853 FILLER_0_10_37/a_6844_375# FILLER_0_11_72/a_2812_375# 0.026339f
C2854 FILLER_0_1_44/a_1380_472# FILLER_0_3_44/a_1468_375# 0.001512f
C2855 FILLER_0_14_37/a_5052_375# vdd 0.00705f
C2856 FILLER_0_8_37/a_4516_472# _14_/I 0.014431f
C2857 FILLER_0_9_2/a_4516_472# FILLER_0_8_37/a_572_375# 0.001723f
C2858 FILLER_0_3_60/a_572_375# FILLER_0_1_60/a_484_472# 0.001512f
C2859 FILLER_0_10_107/a_1020_375# _16_/I 0.001478f
C2860 vdd FILLER_0_5_72/a_2276_472# 0.009744f
C2861 output24/a_224_472# _09_/ZN 0.002668f
C2862 FILLER_0_2_37/a_572_375# _10_/I 0.001886f
C2863 FILLER_0_2_37/a_4068_472# _10_/I 0.002354f
C2864 FILLER_0_0_104/a_36_472# vdd 0.112334f
C2865 _17_/I FILLER_0_13_2/a_3620_472# 0.006613f
C2866 FILLER_0_2_107/a_572_375# _01_/ZN 0.004526f
C2867 _16_/I FILLER_0_11_72/a_5500_375# 0.005899f
C2868 FILLER_0_7_2/a_6308_472# vdd 0.028286f
C2869 _17_/I FILLER_0_15_40/a_1020_375# 0.006589f
C2870 FILLER_0_5_44/a_124_375# _12_/I 0.001706f
C2871 FILLER_0_13_72/a_124_375# FILLER_0_14_37/a_4068_472# 0.001597f
C2872 FILLER_0_7_2/a_6308_472# FILLER_0_8_37/a_2276_472# 0.026657f
C2873 _15_/a_36_113# output_signal_plus[2] 0.039665f
C2874 FILLER_0_4_37/a_36_472# FILLER_0_4_2/a_3260_375# 0.012267f
C2875 FILLER_0_6_101/a_36_472# FILLER_0_5_72/a_3172_472# 0.026657f
C2876 _14_/I FILLER_0_8_28/a_36_472# 0.014431f
C2877 output25/a_224_472# _16_/Z 0.003213f
C2878 output17/a_224_472# FILLER_0_2_107/a_1380_472# 0.031813f
C2879 _18_/I FILLER_0_15_8/a_2812_375# 0.01418f
C2880 _14_/I FILLER_0_9_2/a_5500_375# 0.005381f
C2881 _12_/I FILLER_0_6_2/a_1828_472# 0.018605f
C2882 FILLER_0_6_37/a_1020_375# FILLER_0_8_37/a_932_472# 0.001512f
C2883 FILLER_0_12_37/a_2724_472# FILLER_0_10_37/a_2812_375# 0.001512f
C2884 _18_/I FILLER_0_15_40/a_1468_375# 0.01418f
C2885 FILLER_0_7_104/a_124_375# FILLER_0_5_104/a_36_472# 0.0027f
C2886 output19/a_224_472# output16/a_224_472# 0.031309f
C2887 _16_/Z output28/a_224_472# 0.004477f
C2888 FILLER_0_13_2/a_3172_472# vdd 0.00936f
C2889 _13_/I FILLER_0_6_2/a_1468_375# 0.001706f
C2890 FILLER_0_12_37/a_4604_375# _17_/I 0.002181f
C2891 _17_/I FILLER_0_13_2/a_2276_472# 0.00656f
C2892 FILLER_0_6_37/a_2364_375# _12_/I 0.016091f
C2893 _13_/I FILLER_0_4_37/a_5052_375# 0.005726f
C2894 FILLER_0_15_8/a_1828_472# FILLER_0_16_18/a_572_375# 0.001543f
C2895 FILLER_0_8_12/a_36_472# input_signal[4] 0.073974f
C2896 FILLER_0_12_107/a_1468_375# _17_/I 0.002307f
C2897 FILLER_0_14_115/a_124_375# _17_/I 0.021021f
C2898 output_signal_plus[8] FILLER_0_14_37/a_5948_375# 0.001313f
C2899 FILLER_0_13_66/a_124_375# _16_/I 0.006193f
C2900 output_signal_minus[2] _14_/a_36_113# 0.011258f
C2901 FILLER_0_14_28/a_36_472# _16_/I 0.001667f
C2902 FILLER_0_16_36/a_2724_472# vdd 0.00736f
C2903 FILLER_0_16_36/a_1916_375# vdd 0.00889f
C2904 FILLER_0_4_37/a_1380_472# FILLER_0_5_44/a_572_375# 0.001723f
C2905 FILLER_0_7_2/a_5412_472# _14_/I 0.008683f
C2906 vdd FILLER_0_0_12/a_1468_375# -0.008218f
C2907 FILLER_0_14_115/a_36_472# FILLER_0_14_107/a_572_375# 0.086635f
C2908 _16_/I FILLER_0_11_72/a_6308_472# 0.006064f
C2909 FILLER_0_15_72/a_1468_375# _18_/I 0.014337f
C2910 _15_/I FILLER_0_12_37/a_4964_472# 0.001368f
C2911 _13_/Z _13_/a_36_113# 0.008917f
C2912 FILLER_0_11_72/a_2364_375# FILLER_0_10_37/a_6396_375# 0.026339f
C2913 FILLER_0_14_37/a_4964_472# FILLER_0_12_37/a_5052_375# 0.001512f
C2914 FILLER_0_13_72/a_1468_375# FILLER_0_14_37/a_5412_472# 0.001597f
C2915 _00_/ZN output16/a_224_472# 0.007567f
C2916 FILLER_0_4_37/a_6396_375# FILLER_0_5_72/a_2364_375# 0.026339f
C2917 _08_/ZN vdd 1.437655f
C2918 FILLER_0_9_72/a_36_472# FILLER_0_10_37/a_4068_472# 0.026657f
C2919 FILLER_0_6_37/a_5412_472# FILLER_0_4_37/a_5500_375# 0.001512f
C2920 _09_/ZN FILLER_0_2_107/a_1380_472# 0.003056f
C2921 FILLER_0_12_107/a_932_472# _16_/I 0.017477f
C2922 _09_/ZN FILLER_0_11_72/a_6396_375# 0.002937f
C2923 FILLER_0_4_37/a_6308_472# FILLER_0_5_72/a_2364_375# 0.001723f
C2924 _16_/I FILLER_0_12_37/a_2364_375# 0.016091f
C2925 FILLER_0_3_44/a_1468_375# FILLER_0_2_37/a_2276_472# 0.001723f
C2926 _11_/I FILLER_0_5_12/a_572_375# 0.002201f
C2927 _19_/Z _10_/Z 0.063499f
C2928 _13_/I output_signal_minus[4] 0.141656f
C2929 _11_/I FILLER_0_4_2/a_1380_472# 0.015395f
C2930 FILLER_0_2_107/a_124_375# _10_/I 0.001886f
C2931 output27/a_224_472# output29/a_224_472# 0.001691f
C2932 FILLER_0_10_37/a_2276_472# FILLER_0_8_37/a_2364_375# 0.001512f
C2933 _00_/ZN output20/a_224_472# 0.003458f
C2934 FILLER_0_7_72/a_1020_375# _14_/I 0.008393f
C2935 _12_/a_36_113# _04_/ZN 0.020254f
C2936 FILLER_0_7_104/a_484_472# vdd 0.005198f
C2937 _14_/I _13_/a_36_113# 0.004071f
C2938 FILLER_0_3_60/a_572_375# FILLER_0_3_72/a_36_472# 0.009654f
C2939 FILLER_0_7_72/a_36_472# _12_/I 0.004669f
C2940 FILLER_0_4_37/a_5500_375# vdd 0.009007f
C2941 _11_/I FILLER_0_4_37/a_4964_472# 0.014431f
C2942 output26/a_224_472# output_signal_plus[6] 0.029342f
C2943 FILLER_0_3_72/a_1020_375# FILLER_0_4_37/a_4964_472# 0.001597f
C2944 output_signal_minus[5] _14_/I 0.440158f
C2945 _14_/I FILLER_0_8_101/a_124_375# 0.014572f
C2946 vdd FILLER_0_5_12/a_1468_375# 0.023488f
C2947 FILLER_0_2_107/a_36_472# _10_/I 0.002486f
C2948 output19/a_224_472# FILLER_0_3_104/a_572_375# 0.011584f
C2949 _15_/I _02_/ZN 0.031709f
C2950 FILLER_0_15_8/a_572_375# FILLER_0_14_12/a_124_375# 0.05841f
C2951 FILLER_0_11_72/a_1916_375# _15_/I 0.007126f
C2952 FILLER_0_12_37/a_1916_375# FILLER_0_13_2/a_5948_375# 0.026339f
C2953 _15_/I _10_/Z 0.041954f
C2954 FILLER_0_7_2/a_484_472# vdd 0.007876f
C2955 _17_/I FILLER_0_13_104/a_572_375# 0.006125f
C2956 FILLER_0_14_37/a_932_472# FILLER_0_12_37/a_1020_375# 0.001512f
C2957 FILLER_0_4_37/a_1916_375# _13_/I 0.005593f
C2958 _13_/Z FILLER_0_11_72/a_5948_375# 0.001136f
C2959 FILLER_0_12_37/a_484_472# FILLER_0_11_2/a_4516_472# 0.026657f
C2960 FILLER_0_9_72/a_124_375# FILLER_0_10_37/a_4068_472# 0.001597f
C2961 FILLER_0_10_12/a_36_472# _15_/I 0.02621f
C2962 FILLER_0_0_142/a_572_375# output_signal_minus[8] 0.006083f
C2963 output12/a_224_472# net15 0.145749f
C2964 _08_/ZN output13/a_224_472# 0.02808f
C2965 FILLER_0_11_2/a_3172_472# FILLER_0_12_28/a_124_375# 0.001543f
C2966 FILLER_0_10_101/a_124_375# vdd 0.04319f
C2967 FILLER_0_3_72/a_1380_472# FILLER_0_5_72/a_1468_375# 0.001512f
C2968 _18_/I FILLER_0_14_37/a_1916_375# 0.003979f
C2969 FILLER_0_4_37/a_3620_472# vdd 0.007892f
C2970 vdd FILLER_0_16_36/a_3260_375# 0.03453f
C2971 _15_/I FILLER_0_10_37/a_2276_472# 0.015502f
C2972 output17/a_224_472# _08_/ZN 0.104017f
C2973 FILLER_0_7_72/a_572_375# FILLER_0_5_72/a_484_472# 0.001512f
C2974 FILLER_0_6_37/a_6756_472# FILLER_0_4_37/a_6844_375# 0.001512f
C2975 _14_/I FILLER_0_8_37/a_2812_375# 0.01418f
C2976 vdd FILLER_0_12_37/a_3172_472# 0.006466f
C2977 vdd FILLER_0_9_2/a_124_375# 0.012743f
C2978 FILLER_0_13_2/a_5052_375# FILLER_0_12_37/a_1020_375# 0.026339f
C2979 FILLER_0_6_101/a_36_472# _12_/I 0.017723f
C2980 FILLER_0_9_2/a_3260_375# _14_/I 0.005451f
C2981 _12_/I FILLER_0_6_37/a_5860_472# 0.017477f
C2982 _16_/Z _15_/Z 0.065695f
C2983 FILLER_0_5_12/a_3172_472# FILLER_0_6_37/a_484_472# 0.026657f
C2984 _15_/I FILLER_0_10_107/a_484_472# 0.015502f
C2985 FILLER_0_14_37/a_4156_375# FILLER_0_15_72/a_124_375# 0.026339f
C2986 FILLER_0_2_101/a_124_375# FILLER_0_4_101/a_36_472# 0.001512f
C2987 FILLER_0_6_37/a_5412_472# vdd 0.00624f
C2988 FILLER_0_11_72/a_1468_375# FILLER_0_12_37/a_5412_472# 0.001597f
C2989 _16_/I FILLER_0_13_2/a_484_472# 0.004373f
C2990 vdd input9/a_36_113# 0.017835f
C2991 _11_/I input_signal[2] 0.204298f
C2992 FILLER_0_11_72/a_36_472# vdd 0.108637f
C2993 FILLER_0_8_37/a_1468_375# _15_/I 0.002388f
C2994 _11_/I FILLER_0_5_72/a_1468_375# 0.004712f
C2995 FILLER_0_10_37/a_1916_375# FILLER_0_9_2/a_5860_472# 0.001597f
C2996 _15_/I FILLER_0_9_72/a_1828_472# 0.00652f
C2997 FILLER_0_2_37/a_2724_472# _10_/I 0.002525f
C2998 _16_/I FILLER_0_11_72/a_4156_375# 0.007169f
C2999 FILLER_0_9_72/a_484_472# _14_/I 0.004017f
C3000 FILLER_0_15_56/a_36_472# vdd 0.122339f
C3001 vdd FILLER_0_5_12/a_124_375# 0.033446f
C3002 FILLER_0_7_72/a_36_472# FILLER_0_9_72/a_124_375# 0.001512f
C3003 FILLER_0_1_72/a_1468_375# output_signal_minus[0] 0.017765f
C3004 FILLER_0_6_37/a_2724_472# FILLER_0_4_37/a_2812_375# 0.001512f
C3005 FILLER_0_9_66/a_36_472# FILLER_0_9_72/a_36_472# 0.003468f
C3006 FILLER_0_5_44/a_572_375# FILLER_0_4_37/a_1468_375# 0.026339f
C3007 FILLER_0_9_2/a_6756_472# vdd 0.008994f
C3008 FILLER_0_12_37/a_4068_472# _15_/I 0.001245f
C3009 _13_/I FILLER_0_5_104/a_484_472# 0.023864f
C3010 _14_/I _03_/ZN 0.087081f
C3011 FILLER_0_8_37/a_2276_472# vdd 0.037216f
C3012 input3/a_36_113# FILLER_0_3_12/a_36_472# 0.001663f
C3013 _12_/I FILLER_0_5_72/a_572_375# 0.001706f
C3014 FILLER_0_6_37/a_3708_375# vdd 0.021857f
C3015 FILLER_0_9_72/a_3260_375# FILLER_0_8_101/a_36_472# 0.001723f
C3016 output_signal_minus[6] _04_/ZN 0.002008f
C3017 FILLER_0_14_37/a_5052_375# output30/a_224_472# 0.001234f
C3018 _11_/I FILLER_0_2_2/a_2812_375# 0.00346f
C3019 FILLER_0_1_44/a_572_375# _10_/I 0.008103f
C3020 FILLER_0_3_12/a_2276_472# vdd 0.007367f
C3021 FILLER_0_3_72/a_3260_375# vdd 0.010174f
C3022 FILLER_0_2_37/a_5052_375# _10_/I 0.001886f
C3023 FILLER_0_11_72/a_5412_472# output28/a_224_472# 0.001463f
C3024 output_signal_minus[7] _01_/ZN 0.562775f
C3025 FILLER_0_13_2/a_1020_375# _17_/I 0.006125f
C3026 FILLER_0_14_37/a_5860_472# FILLER_0_12_37/a_5948_375# 0.001512f
C3027 FILLER_0_9_72/a_1468_375# vdd 0.007205f
C3028 FILLER_0_6_37/a_1380_472# _12_/I 0.017477f
C3029 output_signal_plus[6] output29/a_224_472# 0.010207f
C3030 FILLER_0_14_37/a_6396_375# output29/a_224_472# 0.029497f
C3031 FILLER_0_4_37/a_4156_375# vdd 0.004039f
C3032 output12/a_224_472# output_signal_minus[4] 0.001853f
C3033 FILLER_0_13_72/a_36_472# FILLER_0_15_72/a_124_375# 0.001512f
C3034 FILLER_0_2_37/a_5500_375# vdd 0.009317f
C3035 _11_/I FILLER_0_2_2/a_3172_472# 0.002415f
C3036 output13/a_224_472# vdd 0.141765f
C3037 _13_/I FILLER_0_5_72/a_3172_472# 0.018781f
C3038 FILLER_0_5_44/a_1020_375# FILLER_0_6_37/a_1828_472# 0.001597f
C3039 _13_/I _02_/ZN 0.018952f
C3040 _00_/ZN output23/a_224_472# 0.001144f
C3041 _13_/I _10_/Z 0.039074f
C3042 FILLER_0_6_37/a_6844_375# vdd 0.013514f
C3043 FILLER_0_6_2/a_36_472# _12_/I 0.008006f
C3044 FILLER_0_7_2/a_572_375# input_signal[4] 0.003261f
C3045 FILLER_0_0_12/a_36_472# _10_/I 0.025518f
C3046 _12_/I FILLER_0_5_60/a_124_375# 0.001706f
C3047 FILLER_0_12_37/a_4604_375# FILLER_0_13_72/a_572_375# 0.026339f
C3048 _15_/I FILLER_0_11_2/a_3708_375# 0.007218f
C3049 FILLER_0_11_2/a_6308_472# _16_/I 0.007542f
C3050 _19_/I FILLER_0_16_18/a_1468_375# 0.014212f
C3051 FILLER_0_8_107/a_124_375# _15_/I 0.002388f
C3052 FILLER_0_0_142/a_124_375# output_signal_minus[8] 0.005664f
C3053 FILLER_0_4_37/a_36_472# FILLER_0_3_12/a_2724_472# 0.026657f
C3054 output17/a_224_472# vdd 0.03125f
C3055 FILLER_0_13_2/a_5860_472# vdd 0.017991f
C3056 _13_/I FILLER_0_4_101/a_36_472# 0.003497f
C3057 _14_/I _06_/ZN 0.17731f
C3058 output_signal_minus[5] output16/a_224_472# 0.032268f
C3059 FILLER_0_15_2/a_124_375# input_signal[9] 0.005994f
C3060 FILLER_0_7_72/a_932_472# FILLER_0_9_72/a_1020_375# 0.001512f
C3061 FILLER_0_13_2/a_2364_375# vdd 0.024816f
C3062 _17_/I output_signal_plus[8] 0.019638f
C3063 FILLER_0_9_72/a_932_472# FILLER_0_11_72/a_1020_375# 0.001512f
C3064 output23/a_224_472# _14_/Z 0.093853f
C3065 _12_/I FILLER_0_3_12/a_36_472# 0.009048f
C3066 _15_/I FILLER_0_9_72/a_36_472# 0.00652f
C3067 _11_/I FILLER_0_3_44/a_484_472# 0.008683f
C3068 _17_/Z output_signal_plus[7] 0.035866f
C3069 vdd FILLER_0_13_72/a_932_472# 0.004803f
C3070 _11_/I FILLER_0_4_107/a_36_472# 0.014431f
C3071 _15_/I FILLER_0_11_2/a_1468_375# 0.007165f
C3072 FILLER_0_1_12/a_36_472# _10_/I 0.006408f
C3073 input2/a_36_113# vdd 0.104921f
C3074 vdd FILLER_0_5_72/a_36_472# 0.109579f
C3075 FILLER_0_7_2/a_2276_472# vdd 0.012553f
C3076 FILLER_0_7_72/a_1916_375# FILLER_0_6_37/a_5860_472# 0.001723f
C3077 FILLER_0_12_101/a_124_375# FILLER_0_12_107/a_36_472# 0.016748f
C3078 FILLER_0_6_107/a_124_375# _03_/ZN 0.002229f
C3079 _17_/I FILLER_0_15_8/a_1828_472# 0.004125f
C3080 _14_/I output_signal_minus[3] 0.101323f
C3081 FILLER_0_7_2/a_6756_472# _14_/I 0.008683f
C3082 FILLER_0_1_12/a_1916_375# vdd -0.010505f
C3083 vdd FILLER_0_10_37/a_4604_375# 0.004123f
C3084 FILLER_0_14_28/a_124_375# FILLER_0_14_37/a_36_472# 0.007947f
C3085 FILLER_0_9_2/a_4964_472# FILLER_0_10_37/a_932_472# 0.026657f
C3086 FILLER_0_9_72/a_572_375# vdd 0.002455f
C3087 FILLER_0_0_142/a_572_375# _10_/I 0.008906f
C3088 _17_/I FILLER_0_14_107/a_572_375# 0.018729f
C3089 output25/a_224_472# output28/a_224_472# 0.061459f
C3090 FILLER_0_7_2/a_572_375# FILLER_0_6_2/a_572_375# 0.05841f
C3091 _16_/I FILLER_0_12_37/a_6844_375# 0.016091f
C3092 _16_/I FILLER_0_14_107/a_36_472# 0.001667f
C3093 FILLER_0_13_72/a_1828_472# _17_/I 0.00652f
C3094 _15_/I FILLER_0_11_2/a_3620_472# 0.005458f
C3095 vdd FILLER_0_0_36/a_36_472# 0.106034f
C3096 FILLER_0_4_37/a_932_472# vdd 0.005895f
C3097 FILLER_0_2_2/a_2724_472# _11_/I 0.002415f
C3098 _09_/ZN vdd 0.830474f
C3099 FILLER_0_12_37/a_3708_375# vdd 0.021857f
C3100 _11_/I FILLER_0_4_37/a_5860_472# 0.014431f
C3101 FILLER_0_5_12/a_2812_375# vdd 0.002455f
C3102 FILLER_0_3_72/a_2276_472# FILLER_0_5_72/a_2364_375# 0.001512f
C3103 FILLER_0_2_2/a_932_472# _10_/I 0.002192f
C3104 _07_/ZN net15 0.159456f
C3105 FILLER_0_13_72/a_1468_375# FILLER_0_12_37/a_5412_472# 0.001723f
C3106 _15_/I output_signal_plus[4] 0.002234f
C3107 FILLER_0_1_12/a_2812_375# FILLER_0_2_37/a_36_472# 0.001597f
C3108 _15_/I FILLER_0_9_72/a_124_375# 0.006125f
C3109 FILLER_0_0_104/a_124_375# _10_/I 0.010439f
C3110 FILLER_0_5_60/a_36_472# _12_/I 0.003805f
C3111 _19_/I FILLER_0_16_36/a_572_375# 0.01418f
C3112 FILLER_0_10_37/a_572_375# FILLER_0_12_37/a_484_472# 0.001512f
C3113 _15_/I FILLER_0_9_104/a_36_472# 0.006613f
C3114 FILLER_0_9_2/a_5052_375# vdd 0.009047f
C3115 _11_/I FILLER_0_2_2/a_124_375# 0.018139f
C3116 FILLER_0_14_107/a_484_472# _16_/I 0.001667f
C3117 vdd FILLER_0_10_37/a_1020_375# 0.006351f
C3118 FILLER_0_15_40/a_36_472# _17_/I 0.004125f
C3119 FILLER_0_12_12/a_1020_375# vdd 0.025987f
C3120 FILLER_0_2_107/a_1380_472# output_signal_minus[8] 0.031957f
C3121 vdd FILLER_0_9_2/a_36_472# 0.105264f
C3122 _11_/I FILLER_0_2_101/a_36_472# 0.002415f
C3123 _08_/ZN output_signal_minus[2] 0.118532f
C3124 FILLER_0_10_12/a_484_472# FILLER_0_8_12/a_572_375# 0.0027f
C3125 _15_/I FILLER_0_12_37/a_484_472# 0.001368f
C3126 FILLER_0_14_37/a_2276_472# vdd 0.037602f
C3127 _11_/I FILLER_0_3_72/a_1828_472# 0.008683f
C3128 FILLER_0_14_37/a_4964_472# vdd 0.005482f
C3129 FILLER_0_2_37/a_4964_472# FILLER_0_1_72/a_932_472# 0.026657f
C3130 _11_/I output14/a_224_472# 0.097904f
C3131 _11_/I FILLER_0_5_72/a_1020_375# 0.004712f
C3132 FILLER_0_8_12/a_1468_375# FILLER_0_8_28/a_124_375# 0.012001f
C3133 FILLER_0_3_44/a_1468_375# vdd 0.044773f
C3134 _14_/I FILLER_0_9_2/a_5412_472# 0.004017f
C3135 FILLER_0_12_37/a_6308_472# FILLER_0_10_37/a_6396_375# 0.001512f
C3136 FILLER_0_6_37/a_4516_472# _12_/I 0.017477f
C3137 input_signal[5] FILLER_0_9_2/a_124_375# 0.018827f
C3138 FILLER_0_13_72/a_2812_375# FILLER_0_12_37/a_6844_375# 0.026339f
C3139 FILLER_0_9_72/a_3172_472# FILLER_0_11_72/a_3260_375# 0.001512f
C3140 FILLER_0_0_142/a_36_472# output_signal_minus[8] 0.011481f
C3141 FILLER_0_12_37/a_4964_472# _16_/I 0.017477f
C3142 output11/a_224_472# FILLER_0_0_104/a_36_472# 0.001684f
C3143 FILLER_0_12_101/a_36_472# FILLER_0_12_37/a_6844_375# 0.086635f
C3144 _09_/ZN output13/a_224_472# 0.072849f
C3145 FILLER_0_2_37/a_4604_375# _10_/I 0.001788f
C3146 vdd input_signal[1] 0.289969f
C3147 FILLER_0_1_72/a_1380_472# FILLER_0_2_37/a_5412_472# 0.026657f
C3148 FILLER_0_1_72/a_572_375# output20/a_224_472# 0.030009f
C3149 FILLER_0_7_2/a_5500_375# vdd 0.012022f
C3150 _13_/I _12_/I 3.156494f
C3151 FILLER_0_13_104/a_484_472# output28/a_224_472# 0.003196f
C3152 vdd FILLER_0_16_36/a_124_375# 0.009145f
C3153 _00_/ZN output18/a_224_472# 0.089168f
C3154 _13_/I output15/a_224_472# 0.068599f
C3155 FILLER_0_13_66/a_124_375# FILLER_0_13_2/a_6844_375# 0.012001f
C3156 output22/a_224_472# output24/a_224_472# 0.072646f
C3157 FILLER_0_2_2/a_3260_375# FILLER_0_2_37/a_124_375# 0.004426f
C3158 _13_/I FILLER_0_4_37/a_572_375# 0.005726f
C3159 FILLER_0_7_2/a_6756_472# FILLER_0_6_37/a_2812_375# 0.001723f
C3160 _17_/a_36_113# vdd 0.0171f
C3161 output17/a_224_472# _09_/ZN 0.003258f
C3162 _15_/I FILLER_0_8_37/a_1020_375# 0.002388f
C3163 _00_/ZN _15_/I 1.070977f
C3164 vdd FILLER_0_9_2/a_2724_472# 0.009793f
C3165 FILLER_0_4_37/a_1380_472# vdd 0.007577f
C3166 output12/a_224_472# _02_/ZN 0.018348f
C3167 _18_/I FILLER_0_14_37/a_1828_472# 0.001526f
C3168 FILLER_0_8_37/a_36_472# FILLER_0_6_37/a_124_375# 0.001512f
C3169 _14_/I FILLER_0_7_72/a_2812_375# 0.008773f
C3170 output12/a_224_472# _10_/Z 0.061442f
C3171 _15_/a_36_113# _12_/Z 0.016436f
C3172 FILLER_0_6_2/a_484_472# vdd 0.00694f
C3173 _14_/I FILLER_0_6_37/a_4964_472# 0.001219f
C3174 input_signal[5] vdd 0.10807f
C3175 _17_/I _19_/Z 0.004704f
C3176 FILLER_0_14_37/a_4156_375# _17_/I 0.018729f
C3177 input_signal[3] FILLER_0_5_12/a_124_375# 0.010583f
C3178 FILLER_0_9_2/a_2364_375# FILLER_0_8_12/a_1380_472# 0.001684f
C3179 vdd FILLER_0_5_12/a_932_472# 0.01798f
C3180 FILLER_0_1_12/a_2724_472# FILLER_0_2_37/a_36_472# 0.026657f
C3181 input_signal[3] vdd 0.191982f
C3182 output30/a_224_472# vdd 0.098146f
C3183 FILLER_0_6_2/a_124_375# input_signal[4] 0.004381f
C3184 _17_/I FILLER_0_14_37/a_124_375# 0.01911f
C3185 _06_/ZN output16/a_224_472# 0.038768f
C3186 FILLER_0_15_2/a_124_375# FILLER_0_13_2/a_36_472# 0.00108f
C3187 FILLER_0_12_12/a_1468_375# FILLER_0_12_28/a_36_472# 0.086635f
C3188 _14_/I FILLER_0_8_28/a_124_375# 0.014501f
C3189 _14_/I FILLER_0_8_37/a_3260_375# 0.01418f
C3190 _17_/I FILLER_0_14_37/a_3260_375# 0.018729f
C3191 _15_/I _14_/Z 0.321844f
C3192 FILLER_0_11_2/a_5052_375# vdd 0.009047f
C3193 _19_/I FILLER_0_15_8/a_932_472# 0.001964f
C3194 FILLER_0_11_72/a_1916_375# _16_/I 0.007169f
C3195 FILLER_0_7_66/a_124_375# _12_/I 0.006193f
C3196 _16_/I _10_/Z 0.052605f
C3197 FILLER_0_0_142/a_124_375# _10_/I 0.037069f
C3198 _07_/ZN output_signal_minus[4] 0.03949f
C3199 _19_/a_36_113# _19_/I 0.05363f
C3200 output25/a_224_472# _15_/Z 0.059652f
C3201 vdd FILLER_0_2_37/a_1916_375# 0.017898f
C3202 FILLER_0_5_44/a_124_375# FILLER_0_5_12/a_3260_375# 0.012552f
C3203 vdd FILLER_0_0_36/a_124_375# -0.003896f
C3204 _13_/I FILLER_0_4_2/a_3172_472# 0.003497f
C3205 FILLER_0_14_37/a_4964_472# FILLER_0_13_72/a_932_472# 0.026657f
C3206 FILLER_0_12_107/a_484_472# FILLER_0_10_107/a_572_375# 0.001512f
C3207 FILLER_0_1_12/a_1828_472# FILLER_0_2_2/a_2812_375# 0.001543f
C3208 FILLER_0_1_12/a_3172_472# FILLER_0_1_44/a_36_472# 0.013276f
C3209 vdd FILLER_0_4_101/a_124_375# 0.043777f
C3210 output_signal_minus[1] net15 0.002666f
C3211 FILLER_0_2_2/a_1916_375# FILLER_0_1_12/a_932_472# 0.001543f
C3212 _16_/I FILLER_0_12_37/a_2812_375# 0.016091f
C3213 output_signal_minus[2] vdd 0.319435f
C3214 FILLER_0_4_2/a_2276_472# _11_/I 0.014431f
C3215 FILLER_0_2_37/a_1020_375# vdd 0.008544f
C3216 FILLER_0_6_37/a_6756_472# FILLER_0_7_72/a_2812_375# 0.001723f
C3217 FILLER_0_12_107/a_1020_375# output28/a_224_472# 0.029497f
C3218 _11_/I FILLER_0_3_44/a_1020_375# 0.008393f
C3219 _13_/I FILLER_0_5_12/a_1380_472# 0.017477f
C3220 FILLER_0_11_2/a_4068_472# FILLER_0_10_37/a_124_375# 0.001723f
C3221 _18_/I FILLER_0_15_8/a_932_472# 0.016191f
C3222 FILLER_0_7_2/a_4516_472# FILLER_0_9_2/a_4604_375# 0.001512f
C3223 _11_/I FILLER_0_2_37/a_484_472# 0.002415f
C3224 _08_/ZN output_signal_minus[8] 0.043157f
C3225 FILLER_0_2_2/a_3260_375# FILLER_0_2_37/a_36_472# 0.012267f
C3226 _11_/I FILLER_0_4_37/a_2812_375# 0.01418f
C3227 FILLER_0_7_2/a_1380_472# _12_/I 0.004669f
C3228 _19_/a_36_113# _18_/I 0.014821f
C3229 _13_/I FILLER_0_4_37/a_124_375# 0.005726f
C3230 FILLER_0_15_40/a_932_472# FILLER_0_16_36/a_1380_472# 0.05841f
C3231 FILLER_0_9_2/a_3708_375# vdd 0.018728f
C3232 FILLER_0_6_37/a_3172_472# FILLER_0_4_37/a_3260_375# 0.001512f
C3233 _11_/I FILLER_0_5_72/a_3260_375# 0.004712f
C3234 FILLER_0_6_37/a_2276_472# vdd 0.034863f
C3235 FILLER_0_0_70/a_124_375# FILLER_0_1_72/a_36_472# 0.001684f
C3236 _11_/I FILLER_0_3_72/a_36_472# 0.008683f
C3237 FILLER_0_13_72/a_36_472# _17_/I 0.00652f
C3238 _15_/I output_signal_plus[3] 0.398979f
C3239 input2/a_36_113# input_signal[1] 0.059503f
C3240 FILLER_0_8_12/a_124_375# input_signal[4] 0.005753f
C3241 FILLER_0_9_2/a_6844_375# FILLER_0_9_66/a_124_375# 0.012001f
C3242 FILLER_0_2_37/a_2276_472# _10_/I 0.001022f
C3243 _15_/I FILLER_0_10_37/a_6844_375# 0.018729f
C3244 FILLER_0_4_37/a_484_472# FILLER_0_5_12/a_3260_375# 0.001723f
C3245 FILLER_0_8_37/a_1828_472# FILLER_0_7_2/a_5860_472# 0.026657f
C3246 output29/a_224_472# _18_/Z 0.019031f
C3247 vdd FILLER_0_14_37/a_484_472# 0.004128f
C3248 FILLER_0_14_101/a_36_472# _16_/I 0.001667f
C3249 _15_/I FILLER_0_9_2/a_5500_375# 0.006125f
C3250 FILLER_0_9_72/a_1380_472# vdd 0.006325f
C3251 FILLER_0_4_2/a_1916_375# FILLER_0_6_2/a_1828_472# 0.0027f
C3252 _18_/I FILLER_0_14_37/a_5052_375# 0.003988f
C3253 FILLER_0_12_107/a_484_472# FILLER_0_11_72/a_4516_472# 0.026657f
C3254 FILLER_0_12_37/a_4068_472# _16_/I 0.017477f
C3255 FILLER_0_4_2/a_124_375# FILLER_0_6_2/a_36_472# 0.00108f
C3256 FILLER_0_10_37/a_5052_375# _15_/I 0.018729f
C3257 _17_/I FILLER_0_13_72/a_1916_375# 0.006125f
C3258 FILLER_0_1_12/a_3260_375# FILLER_0_1_44/a_36_472# 0.086905f
C3259 output_signal_minus[2] output13/a_224_472# 0.028204f
C3260 FILLER_0_11_72/a_5052_375# vdd 0.004637f
C3261 FILLER_0_11_136/a_36_472# FILLER_0_11_72/a_6756_472# 0.013276f
C3262 FILLER_0_11_72/a_2724_472# FILLER_0_12_37/a_6756_472# 0.026657f
C3263 FILLER_0_1_12/a_1020_375# vdd -0.005745f
C3264 FILLER_0_14_28/a_124_375# FILLER_0_15_8/a_2364_375# 0.05841f
C3265 FILLER_0_15_2/a_124_375# FILLER_0_15_8/a_124_375# 0.003598f
C3266 output_signal_plus[7] output26/a_224_472# 0.030595f
C3267 _00_/ZN _13_/I 0.18426f
C3268 FILLER_0_16_36/a_2724_472# _19_/I 0.019067f
C3269 FILLER_0_16_36/a_1916_375# _19_/I 0.014588f
C3270 vdd FILLER_0_4_37/a_1468_375# 0.01039f
C3271 vdd FILLER_0_11_2/a_484_472# 0.007876f
C3272 _09_/ZN FILLER_0_4_107/a_932_472# 0.047259f
C3273 output12/a_224_472# _12_/I 0.09633f
C3274 _15_/I FILLER_0_10_37/a_124_375# 0.01911f
C3275 output12/a_224_472# output15/a_224_472# 0.072646f
C3276 _14_/I FILLER_0_7_2/a_3260_375# 0.008393f
C3277 vdd FILLER_0_14_37/a_3620_472# 0.00818f
C3278 FILLER_0_1_60/a_572_375# vdd 0.011591f
C3279 _15_/I FILLER_0_10_37/a_3620_472# 0.015502f
C3280 FILLER_0_15_72/a_36_472# vdd 0.112218f
C3281 FILLER_0_2_37/a_4516_472# vdd 0.003374f
C3282 FILLER_0_14_12/a_932_472# FILLER_0_13_2/a_1916_375# 0.001543f
C3283 _15_/I FILLER_0_10_37/a_1828_472# 0.015502f
C3284 FILLER_0_13_2/a_5948_375# FILLER_0_11_2/a_5860_472# 0.001512f
C3285 FILLER_0_0_142/a_36_472# _10_/I 0.072794f
C3286 FILLER_0_4_2/a_1468_375# vdd 0.027303f
C3287 FILLER_0_14_37/a_2812_375# _17_/I 0.018729f
C3288 FILLER_0_10_37/a_4964_472# vdd 0.005482f
C3289 FILLER_0_10_12/a_124_375# FILLER_0_11_2/a_1380_472# 0.001684f
C3290 FILLER_0_8_37/a_1828_472# FILLER_0_6_37/a_1916_375# 0.001512f
C3291 _11_/I FILLER_0_3_72/a_932_472# 0.008683f
C3292 input_signal[5] FILLER_0_9_2/a_36_472# 0.039749f
C3293 FILLER_0_11_2/a_1828_472# FILLER_0_12_12/a_572_375# 0.001543f
C3294 _19_/a_36_113# _18_/a_36_113# 0.001578f
C3295 output_signal_minus[1] output_signal_minus[4] 0.001687f
C3296 FILLER_0_16_18/a_36_472# input_signal[9] 0.070705f
C3297 output11/a_224_472# vdd 0.07857f
C3298 FILLER_0_4_37/a_484_472# FILLER_0_2_37/a_572_375# 0.001512f
C3299 FILLER_0_11_2/a_2812_375# FILLER_0_12_28/a_36_472# 0.001543f
C3300 FILLER_0_11_2/a_3708_375# _16_/I 0.005447f
C3301 FILLER_0_8_37/a_572_375# FILLER_0_9_2/a_4604_375# 0.026339f
C3302 _16_/I FILLER_0_13_72/a_1380_472# 0.004669f
C3303 FILLER_0_0_12/a_1380_472# vdd 0.005476f
C3304 FILLER_0_16_36/a_2724_472# _18_/I 0.001782f
C3305 vdd FILLER_0_14_37/a_6308_472# 0.021839f
C3306 FILLER_0_0_104/a_36_472# _10_/I 0.007714f
C3307 FILLER_0_2_2/a_1380_472# vdd 0.013839f
C3308 FILLER_0_7_104/a_36_472# _14_/I 0.013033f
C3309 FILLER_0_4_37/a_6396_375# vdd 0.038622f
C3310 FILLER_0_9_2/a_4964_472# vdd 0.006804f
C3311 FILLER_0_6_37/a_1828_472# _14_/I 0.001219f
C3312 FILLER_0_12_37/a_5052_375# FILLER_0_13_72/a_1020_375# 0.026339f
C3313 _13_/I FILLER_0_4_107/a_124_375# 0.005716f
C3314 FILLER_0_13_72/a_3172_472# vdd 0.009788f
C3315 FILLER_0_11_2/a_5052_375# FILLER_0_10_37/a_1020_375# 0.026339f
C3316 _14_/I FILLER_0_9_2/a_4156_375# 0.005381f
C3317 vdd output_signal_minus[8] 0.451417f
C3318 FILLER_0_4_37/a_6308_472# vdd 0.020611f
C3319 FILLER_0_0_36/a_2364_375# vdd 0.020934f
C3320 _15_/I FILLER_0_8_101/a_124_375# 0.002388f
C3321 vdd input_signal[7] 0.09759f
C3322 output23/a_224_472# _06_/ZN 0.001429f
C3323 FILLER_0_11_66/a_36_472# FILLER_0_11_2/a_6844_375# 0.086635f
C3324 _09_/ZN output_signal_minus[2] 0.002008f
C3325 FILLER_0_1_72/a_1380_472# output_signal_minus[0] 0.002792f
C3326 FILLER_0_2_37/a_1020_375# FILLER_0_4_37/a_932_472# 0.001512f
C3327 FILLER_0_3_72/a_3260_375# output11/a_224_472# 0.001216f
C3328 FILLER_0_11_72/a_6844_375# _13_/Z 0.029766f
C3329 _07_/ZN _10_/Z 1.66841f
C3330 FILLER_0_3_12/a_3260_375# FILLER_0_2_37/a_572_375# 0.026339f
C3331 _15_/I FILLER_0_11_72/a_932_472# 0.005458f
C3332 FILLER_0_12_37/a_2724_472# _15_/I 0.001368f
C3333 FILLER_0_9_2/a_6308_472# FILLER_0_11_2/a_6396_375# 0.001512f
C3334 output22/a_224_472# _08_/ZN 0.030901f
C3335 FILLER_0_2_37/a_3260_375# vdd 0.008869f
C3336 _16_/I FILLER_0_11_2/a_1468_375# 0.007169f
C3337 _11_/I FILLER_0_5_44/a_484_472# 0.001913f
C3338 FILLER_0_14_101/a_124_375# output_signal_plus[8] 0.002612f
C3339 FILLER_0_14_28/a_36_472# FILLER_0_13_2/a_2812_375# 0.001543f
C3340 FILLER_0_15_56/a_124_375# vdd 0.048221f
C3341 FILLER_0_14_37/a_3172_472# _17_/I 0.015502f
C3342 _11_/I _11_/Z 0.208356f
C3343 _19_/I FILLER_0_16_36/a_3260_375# 0.018198f
C3344 FILLER_0_3_104/a_572_375# FILLER_0_2_107/a_124_375# 0.026339f
C3345 vdd FILLER_0_5_72/a_124_375# 0.013594f
C3346 output19/a_224_472# FILLER_0_3_104/a_484_472# 0.002002f
C3347 output27/a_224_472# _10_/Z 0.166209f
C3348 FILLER_0_11_2/a_3620_472# _16_/I 0.00769f
C3349 _15_/I FILLER_0_8_37/a_2812_375# 0.002388f
C3350 input10/a_36_113# input9/a_36_113# 0.001578f
C3351 FILLER_0_14_12/a_484_472# vdd 0.023895f
C3352 _10_/I FILLER_0_0_12/a_1468_375# 0.015932f
C3353 FILLER_0_6_37/a_5860_472# FILLER_0_5_72/a_1916_375# 0.001597f
C3354 vdd FILLER_0_13_2/a_6396_375# 0.014009f
C3355 _15_/I FILLER_0_9_2/a_3260_375# 0.006125f
C3356 output17/a_224_472# output11/a_224_472# 0.001691f
C3357 FILLER_0_2_107/a_1468_375# vdd 0.016357f
C3358 _14_/I _14_/a_36_113# 0.046735f
C3359 _15_/I FILLER_0_11_72/a_5948_375# 0.00726f
C3360 FILLER_0_10_28/a_36_472# FILLER_0_10_12/a_1380_472# 0.013277f
C3361 output_signal_plus[5] _10_/Z 0.093318f
C3362 FILLER_0_12_37/a_1468_375# _16_/I 0.016091f
C3363 _19_/I input9/a_36_113# 0.18911f
C3364 _16_/I output_signal_plus[4] 0.256241f
C3365 FILLER_0_10_107/a_36_472# FILLER_0_8_107/a_124_375# 0.001512f
C3366 _11_/I FILLER_0_3_72/a_2812_375# 0.008393f
C3367 _08_/ZN _10_/I 0.099908f
C3368 FILLER_0_9_2/a_1020_375# FILLER_0_7_2/a_932_472# 0.0027f
C3369 input10/a_36_113# vdd 0.107237f
C3370 _09_/ZN FILLER_0_11_72/a_5052_375# 0.013107f
C3371 _11_/I FILLER_0_2_37/a_6308_472# 0.001793f
C3372 output17/a_224_472# output_signal_minus[8] 0.084186f
C3373 _14_/I FILLER_0_7_2/a_932_472# 0.008787f
C3374 input7/a_36_113# _16_/I 0.003764f
C3375 FILLER_0_15_56/a_36_472# _19_/I 0.001782f
C3376 FILLER_0_10_37/a_3708_375# vdd 0.021519f
C3377 _18_/I FILLER_0_16_36/a_3260_375# 0.001989f
C3378 _16_/I FILLER_0_12_37/a_484_472# 0.017477f
C3379 FILLER_0_1_12/a_2276_472# FILLER_0_3_12/a_2364_375# 0.0027f
C3380 _15_/I FILLER_0_9_72/a_484_472# 0.001644f
C3381 _17_/I FILLER_0_12_37/a_572_375# 0.002388f
C3382 _15_/Z output_signal_plus[1] 0.012051f
C3383 _19_/I vdd 1.003458f
C3384 output14/a_224_472# FILLER_0_4_107/a_1380_472# 0.002338f
C3385 vdd FILLER_0_4_37/a_2724_472# 0.009424f
C3386 FILLER_0_12_37/a_4156_375# _16_/I 0.016091f
C3387 FILLER_0_2_37/a_6844_375# vdd 0.013868f
C3388 FILLER_0_7_2/a_5860_472# FILLER_0_8_37/a_1916_375# 0.001597f
C3389 FILLER_0_4_37/a_4156_375# FILLER_0_5_72/a_124_375# 0.026339f
C3390 FILLER_0_2_2/a_2724_472# FILLER_0_1_12/a_1468_375# 0.001543f
C3391 output21/a_224_472# _10_/Z 0.055413f
C3392 FILLER_0_12_37/a_3708_375# FILLER_0_14_37/a_3620_472# 0.0027f
C3393 vdd FILLER_0_16_18/a_484_472# 0.013106f
C3394 FILLER_0_5_12/a_1916_375# FILLER_0_6_2/a_3172_472# 0.001543f
C3395 FILLER_0_8_37/a_36_472# _14_/I 0.014431f
C3396 _00_/ZN output12/a_224_472# 0.004121f
C3397 _17_/Z _16_/Z 0.301563f
C3398 FILLER_0_12_12/a_36_472# vdd 0.014415f
C3399 _14_/I FILLER_0_7_2/a_4964_472# 0.008683f
C3400 _18_/I input9/a_36_113# 0.004981f
C3401 _17_/I FILLER_0_14_37/a_3708_375# 0.018729f
C3402 FILLER_0_15_72/a_1380_472# output29/a_224_472# 0.005437f
C3403 FILLER_0_13_2/a_4156_375# vdd 0.004039f
C3404 output24/a_224_472# _13_/Z 0.010438f
C3405 vdd FILLER_0_15_8/a_484_472# 0.010346f
C3406 FILLER_0_14_37/a_3172_472# FILLER_0_12_37/a_3260_375# 0.001512f
C3407 _08_/ZN _16_/a_36_113# 0.152085f
C3408 _13_/I FILLER_0_4_37/a_6844_375# 0.005726f
C3409 _18_/I FILLER_0_15_56/a_36_472# 0.014431f
C3410 FILLER_0_3_12/a_3260_375# FILLER_0_3_44/a_124_375# 0.012552f
C3411 FILLER_0_14_37/a_572_375# FILLER_0_15_40/a_124_375# 0.026339f
C3412 _18_/I vdd 1.307286f
C3413 FILLER_0_15_64/a_124_375# vdd 0.033433f
C3414 FILLER_0_13_72/a_484_472# vdd 0.002467f
C3415 output17/a_224_472# FILLER_0_2_107/a_1468_375# 0.001597f
C3416 FILLER_0_4_2/a_36_472# _11_/I 0.001145f
C3417 _13_/I _13_/a_36_113# 0.011803f
C3418 FILLER_0_4_2/a_2364_375# FILLER_0_5_12/a_1380_472# 0.001684f
C3419 FILLER_0_2_2/a_36_472# vdd 0.106171f
C3420 _16_/I FILLER_0_12_12/a_572_375# 0.016141f
C3421 FILLER_0_9_104/a_572_375# FILLER_0_7_104/a_484_472# 0.001512f
C3422 _04_/ZN output_signal_minus[4] 0.033175f
C3423 output22/a_224_472# vdd 0.157202f
C3424 _09_/ZN output_signal_minus[8] 0.012193f
C3425 FILLER_0_5_44/a_1020_375# vdd 0.011235f
C3426 output_signal_minus[5] _13_/I 0.054563f
C3427 FILLER_0_3_104/a_484_472# FILLER_0_4_107/a_124_375# 0.001597f
C3428 _14_/I FILLER_0_9_2/a_5948_375# 0.003376f
C3429 _12_/I FILLER_0_4_2/a_932_472# 0.005926f
C3430 output_signal_minus[1] _02_/ZN 0.002436f
C3431 output_signal_minus[1] _10_/Z 0.070547f
C3432 FILLER_0_3_72/a_484_472# FILLER_0_5_72/a_572_375# 0.001512f
C3433 FILLER_0_15_72/a_1468_375# output_signal_plus[8] 0.017765f
C3434 FILLER_0_9_2/a_4964_472# FILLER_0_10_37/a_1020_375# 0.001597f
C3435 _15_/I FILLER_0_12_37/a_1828_472# 0.001368f
C3436 vdd FILLER_0_7_72/a_2724_472# 0.034108f
C3437 _07_/ZN _12_/I 0.033218f
C3438 vdd FILLER_0_14_12/a_1468_375# -0.008399f
C3439 _00_/ZN output_signal_minus[0] 0.074904f
C3440 _07_/ZN output15/a_224_472# 0.083164f
C3441 _16_/I _14_/Z 0.44239f
C3442 _15_/I _06_/ZN 0.015378f
C3443 FILLER_0_9_2/a_1468_375# vdd 0.027811f
C3444 _11_/I FILLER_0_5_104/a_36_472# 0.001913f
C3445 FILLER_0_7_2/a_572_375# _12_/I 0.006109f
C3446 _17_/I _16_/I 0.016418f
C3447 FILLER_0_11_72/a_36_472# FILLER_0_13_72/a_124_375# 0.001512f
C3448 FILLER_0_4_37/a_5948_375# vdd 0.011562f
C3449 _14_/I FILLER_0_8_37/a_5500_375# 0.01418f
C3450 FILLER_0_5_12/a_484_472# _13_/I 0.017477f
C3451 _14_/I FILLER_0_6_101/a_124_375# 0.003099f
C3452 vdd _10_/I 1.971103f
C3453 output_signal_plus[6] _10_/Z 0.112218f
C3454 FILLER_0_5_12/a_2364_375# vdd 0.019634f
C3455 FILLER_0_13_72/a_124_375# vdd 0.011994f
C3456 _09_/ZN FILLER_0_2_107/a_1468_375# 0.028929f
C3457 FILLER_0_6_37/a_124_375# vdd 0.012548f
C3458 output22/a_224_472# output13/a_224_472# 0.004655f
C3459 FILLER_0_6_37/a_6756_472# FILLER_0_5_72/a_2724_472# 0.026657f
C3460 FILLER_0_14_37/a_2276_472# FILLER_0_15_56/a_124_375# 0.001723f
C3461 _13_/Z FILLER_0_11_72/a_6396_375# 0.032765f
C3462 _14_/I FILLER_0_9_2/a_4068_472# 0.004017f
C3463 FILLER_0_2_37/a_6756_472# output_signal_minus[0] 0.001292f
C3464 FILLER_0_8_12/a_932_472# vdd 0.019362f
C3465 _18_/a_36_113# vdd 0.018573f
C3466 FILLER_0_14_37/a_4604_375# FILLER_0_15_72/a_572_375# 0.026339f
C3467 FILLER_0_5_12/a_2364_375# FILLER_0_3_12/a_2276_472# 0.0027f
C3468 FILLER_0_5_72/a_484_472# _12_/I 0.001371f
C3469 FILLER_0_11_2/a_6756_472# FILLER_0_11_66/a_36_472# 0.013276f
C3470 _16_/I output_signal_plus[3] 0.005193f
C3471 _13_/I FILLER_0_4_37/a_3708_375# 0.005846f
C3472 output20/a_224_472# FILLER_0_0_104/a_124_375# 0.001073f
C3473 FILLER_0_7_2/a_4516_472# FILLER_0_6_37/a_572_375# 0.001723f
C3474 FILLER_0_13_2/a_6844_375# FILLER_0_12_37/a_2812_375# 0.026339f
C3475 _17_/I FILLER_0_13_72/a_2812_375# 0.006125f
C3476 FILLER_0_9_104/a_572_375# vdd 0.018731f
C3477 vdd _16_/a_36_113# 0.013616f
C3478 _16_/I FILLER_0_10_37/a_6844_375# 0.002327f
C3479 _11_/I FILLER_0_3_44/a_932_472# 0.008683f
C3480 FILLER_0_9_66/a_36_472# FILLER_0_8_37/a_3260_375# 0.001723f
C3481 FILLER_0_2_107/a_1380_472# _14_/I 0.004574f
C3482 _13_/I FILLER_0_4_107/a_1468_375# 0.003168f
C3483 _13_/I _03_/ZN 0.152144f
C3484 _07_/ZN output_signal_plus[4] 0.005998f
C3485 FILLER_0_11_72/a_124_375# FILLER_0_12_37/a_4068_472# 0.001597f
C3486 FILLER_0_9_2/a_4964_472# FILLER_0_11_2/a_5052_375# 0.001512f
C3487 FILLER_0_2_37/a_5500_375# _10_/I 0.001886f
C3488 FILLER_0_13_2/a_5948_375# vdd 0.032268f
C3489 FILLER_0_13_72/a_36_472# FILLER_0_14_37/a_4068_472# 0.026657f
C3490 _11_/Z FILLER_0_9_104/a_484_472# 0.004443f
C3491 vdd FILLER_0_9_2/a_2276_472# 0.012553f
C3492 _16_/I FILLER_0_12_37/a_3260_375# 0.016091f
C3493 _13_/I FILLER_0_5_12/a_3260_375# 0.016091f
C3494 FILLER_0_3_72/a_2276_472# vdd 0.011667f
C3495 FILLER_0_10_37/a_5052_375# _16_/I 0.002327f
C3496 FILLER_0_10_12/a_36_472# FILLER_0_11_2/a_1020_375# 0.001684f
C3497 FILLER_0_8_37/a_6308_472# FILLER_0_9_72/a_2364_375# 0.001723f
C3498 FILLER_0_6_2/a_3172_472# FILLER_0_4_2/a_3260_375# 0.0027f
C3499 output17/a_224_472# _10_/I 0.012887f
C3500 _07_/ZN output19/a_224_472# 0.05503f
C3501 vdd FILLER_0_4_107/a_484_472# 0.005163f
C3502 FILLER_0_15_8/a_3260_375# FILLER_0_14_37/a_36_472# 0.001723f
C3503 _09_/ZN _18_/I 0.028145f
C3504 _15_/I FILLER_0_9_2/a_5412_472# 0.006506f
C3505 output_signal_plus[2] _15_/Z 0.042147f
C3506 output22/a_224_472# _09_/ZN 0.076985f
C3507 FILLER_0_2_37/a_1380_472# FILLER_0_1_44/a_484_472# 0.026657f
C3508 FILLER_0_10_101/a_36_472# vdd 0.098751f
C3509 output_signal_minus[9] FILLER_0_0_142/a_36_472# 0.001011f
C3510 output_signal_plus[5] output_signal_plus[4] 0.147694f
C3511 _15_/I FILLER_0_10_12/a_932_472# 0.015565f
C3512 output_signal_minus[6] _01_/ZN 0.094353f
C3513 FILLER_0_5_44/a_932_472# _13_/I 0.017477f
C3514 FILLER_0_5_72/a_932_472# _12_/I 0.003805f
C3515 FILLER_0_16_104/a_36_472# output29/a_224_472# 0.001178f
C3516 FILLER_0_9_72/a_2812_375# FILLER_0_8_37/a_6756_472# 0.001723f
C3517 FILLER_0_7_2/a_3620_472# _12_/I 0.004669f
C3518 output_signal_minus[1] _12_/I 0.079399f
C3519 output12/a_224_472# _13_/a_36_113# 0.008132f
C3520 FILLER_0_14_28/a_124_375# _17_/I 0.021137f
C3521 FILLER_0_7_2/a_6308_472# _14_/I 0.008683f
C3522 FILLER_0_6_107/a_124_375# FILLER_0_6_101/a_124_375# 0.005439f
C3523 FILLER_0_12_107/a_1380_472# FILLER_0_11_72/a_5412_472# 0.026657f
C3524 FILLER_0_8_37/a_4068_472# FILLER_0_9_72/a_124_375# 0.001723f
C3525 FILLER_0_10_12/a_36_472# FILLER_0_8_12/a_124_375# 0.0027f
C3526 _13_/I FILLER_0_5_72/a_1916_375# 0.016091f
C3527 _19_/I FILLER_0_16_36/a_124_375# 0.01418f
C3528 vdd FILLER_0_13_72/a_1020_375# 0.00558f
C3529 _13_/I FILLER_0_4_2/a_1916_375# 0.001863f
C3530 FILLER_0_7_2/a_2724_472# vdd 0.009793f
C3531 _17_/a_36_113# _19_/I 0.006856f
C3532 FILLER_0_14_37/a_4964_472# _18_/I 0.001526f
C3533 vdd FILLER_0_1_44/a_932_472# 0.009767f
C3534 _13_/I _06_/ZN 0.88854f
C3535 FILLER_0_14_101/a_36_472# FILLER_0_13_72/a_3260_375# 0.001597f
C3536 output_signal_minus[9] FILLER_0_0_104/a_36_472# 0.002951f
C3537 FILLER_0_12_37/a_1468_375# FILLER_0_14_37/a_1380_472# 0.001512f
C3538 FILLER_0_4_37/a_6756_472# FILLER_0_4_101/a_36_472# 0.013277f
C3539 _02_/ZN _04_/ZN 0.005252f
C3540 FILLER_0_1_12/a_1916_375# _10_/I 0.008103f
C3541 FILLER_0_13_2/a_3260_375# _16_/I 0.006272f
C3542 _13_/I _10_/a_36_160# 0.058633f
C3543 FILLER_0_11_2/a_5412_472# _15_/I 0.005458f
C3544 FILLER_0_7_72/a_124_375# vdd 0.011994f
C3545 FILLER_0_14_37/a_2812_375# FILLER_0_13_2/a_6756_472# 0.001597f
C3546 _17_/I FILLER_0_15_72/a_932_472# 0.004125f
C3547 FILLER_0_12_37/a_5500_375# vdd 0.009137f
C3548 FILLER_0_8_37/a_124_375# FILLER_0_10_37/a_36_472# 0.001512f
C3549 _19_/I output30/a_224_472# 0.121547f
C3550 FILLER_0_6_37/a_6308_472# FILLER_0_7_72/a_2364_375# 0.001723f
C3551 FILLER_0_2_101/a_124_375# FILLER_0_2_107/a_124_375# 0.005439f
C3552 FILLER_0_0_36/a_36_472# _10_/I 0.0157f
C3553 _13_/Z _08_/ZN 0.004526f
C3554 FILLER_0_2_37/a_2812_375# FILLER_0_3_60/a_124_375# 0.026339f
C3555 FILLER_0_7_2/a_1468_375# FILLER_0_6_2/a_1468_375# 0.05841f
C3556 _15_/I FILLER_0_8_28/a_124_375# 0.002388f
C3557 _15_/I FILLER_0_8_37/a_3260_375# 0.002388f
C3558 FILLER_0_11_72/a_124_375# FILLER_0_9_72/a_36_472# 0.001512f
C3559 _11_/I FILLER_0_2_107/a_572_375# 0.003106f
C3560 _07_/ZN _14_/Z 0.032414f
C3561 FILLER_0_11_2/a_5500_375# FILLER_0_9_2/a_5412_472# 0.001512f
C3562 FILLER_0_2_2/a_36_472# input_signal[1] 0.021174f
C3563 _17_/a_36_113# _18_/I 0.002684f
C3564 FILLER_0_6_2/a_124_375# _12_/I 0.005373f
C3565 FILLER_0_5_60/a_36_472# FILLER_0_5_44/a_1380_472# 0.013276f
C3566 _13_/I output_signal_minus[3] 0.171411f
C3567 _16_/I FILLER_0_11_72/a_932_472# 0.00753f
C3568 FILLER_0_7_104/a_36_472# FILLER_0_9_104/a_124_375# 0.0027f
C3569 FILLER_0_2_101/a_124_375# FILLER_0_2_107/a_36_472# 0.016748f
C3570 _13_/I FILLER_0_4_107/a_572_375# 0.005848f
C3571 FILLER_0_6_2/a_1916_375# FILLER_0_7_2/a_1916_375# 0.05841f
C3572 FILLER_0_12_37/a_2724_472# _16_/I 0.017477f
C3573 _11_/I FILLER_0_5_12/a_1020_375# 0.004745f
C3574 FILLER_0_8_107/a_572_375# FILLER_0_10_107/a_484_472# 0.0027f
C3575 _16_/Z output26/a_224_472# 0.227699f
C3576 _00_/ZN output_signal_plus[5] 0.041491f
C3577 FILLER_0_10_107/a_932_472# _15_/I 0.015502f
C3578 _11_/I FILLER_0_2_37/a_1468_375# 0.00346f
C3579 FILLER_0_6_37/a_5948_375# vdd 0.011644f
C3580 _18_/I output30/a_224_472# 0.023746f
C3581 output_signal_plus[2] output_signal_plus[1] 0.186309f
C3582 FILLER_0_14_107/a_484_472# _18_/Z 0.001168f
C3583 FILLER_0_9_2/a_5412_472# FILLER_0_10_37/a_1468_375# 0.001597f
C3584 _08_/ZN _14_/I 0.130623f
C3585 FILLER_0_12_101/a_124_375# FILLER_0_12_37/a_6844_375# 0.012001f
C3586 _17_/I output27/a_224_472# 0.024557f
C3587 vdd FILLER_0_11_72/a_3620_472# 0.009735f
C3588 FILLER_0_4_2/a_1380_472# FILLER_0_3_12/a_124_375# 0.001543f
C3589 _17_/I FILLER_0_15_8/a_2276_472# 0.004125f
C3590 FILLER_0_1_12/a_484_472# FILLER_0_3_12/a_572_375# 0.0027f
C3591 FILLER_0_15_8/a_2364_375# FILLER_0_16_18/a_1380_472# 0.001543f
C3592 vdd FILLER_0_10_37/a_2812_375# 0.008466f
C3593 FILLER_0_2_2/a_1020_375# FILLER_0_1_12/a_36_472# 0.001543f
C3594 output_signal_minus[9] _08_/ZN 0.002843f
C3595 output_signal_plus[5] _14_/Z 0.001613f
C3596 FILLER_0_12_37/a_4964_472# FILLER_0_11_72/a_1020_375# 0.001597f
C3597 FILLER_0_9_2/a_6756_472# FILLER_0_10_37/a_2812_375# 0.001597f
C3598 output25/a_224_472# FILLER_0_12_107/a_1380_472# 0.002618f
C3599 _16_/I FILLER_0_11_72/a_5948_375# 0.007169f
C3600 vdd FILLER_0_10_37/a_6308_472# 0.021839f
C3601 input_signal[1] _10_/I 0.089061f
C3602 _13_/I FILLER_0_4_37/a_3172_472# 0.003497f
C3603 output29/a_224_472# FILLER_0_13_72/a_2724_472# 0.001243f
C3604 FILLER_0_3_72/a_572_375# _11_/I 0.005f
C3605 FILLER_0_7_104/a_484_472# _14_/I 0.026299f
C3606 output_signal_plus[5] _17_/I 0.253985f
C3607 FILLER_0_12_107/a_484_472# vdd 0.003157f
C3608 output11/a_224_472# output_signal_minus[8] 0.002981f
C3609 _13_/I FILLER_0_5_44/a_1380_472# 0.017477f
C3610 output25/a_224_472# _17_/Z 0.12295f
C3611 _15_/I FILLER_0_11_2/a_572_375# 0.007774f
C3612 FILLER_0_2_107/a_1380_472# output16/a_224_472# 0.002338f
C3613 FILLER_0_2_37/a_932_472# _11_/I 0.002415f
C3614 _16_/I FILLER_0_13_72/a_572_375# 0.006182f
C3615 _07_/ZN output_signal_plus[3] 0.023981f
C3616 _09_/ZN FILLER_0_4_107/a_484_472# 0.005391f
C3617 FILLER_0_0_12/a_124_375# input_signal[1] 0.001377f
C3618 vdd FILLER_0_11_2/a_4964_472# 0.006804f
C3619 _11_/I FILLER_0_3_104/a_36_472# 0.008761f
C3620 FILLER_0_4_37/a_1828_472# vdd 0.010074f
C3621 FILLER_0_13_104/a_124_375# vdd 0.027844f
C3622 _17_/I FILLER_0_14_37/a_2364_375# 0.018729f
C3623 FILLER_0_12_37/a_124_375# vdd 0.013676f
C3624 FILLER_0_11_2/a_5412_472# FILLER_0_10_37/a_1468_375# 0.001723f
C3625 _17_/Z output28/a_224_472# 0.032609f
C3626 _15_/I FILLER_0_11_2/a_2812_375# 0.007165f
C3627 FILLER_0_7_2/a_484_472# _14_/I 0.009189f
C3628 _17_/I FILLER_0_14_12/a_572_375# 0.018801f
C3629 _17_/I FILLER_0_14_37/a_1380_472# 0.015502f
C3630 FILLER_0_8_12/a_1468_375# vdd 0.024301f
C3631 _15_/I FILLER_0_11_72/a_1380_472# 0.005458f
C3632 FILLER_0_7_72/a_124_375# FILLER_0_5_72/a_36_472# 0.001512f
C3633 FILLER_0_2_37/a_5860_472# output_signal_minus[0] 0.001069f
C3634 FILLER_0_15_64/a_36_472# vdd 0.094137f
C3635 FILLER_0_12_37/a_572_375# FILLER_0_13_2/a_4516_472# 0.001723f
C3636 _12_/I FILLER_0_5_60/a_484_472# 0.003805f
C3637 vdd FILLER_0_2_37/a_6396_375# 0.040336f
C3638 FILLER_0_10_37/a_124_375# FILLER_0_10_28/a_124_375# 0.003228f
C3639 vdd FILLER_0_0_70/a_36_472# 0.109853f
C3640 _00_/ZN output_signal_minus[1] 0.041447f
C3641 FILLER_0_2_37/a_6308_472# FILLER_0_3_72/a_2364_375# 0.001723f
C3642 FILLER_0_10_107/a_124_375# FILLER_0_11_72/a_4068_472# 0.001723f
C3643 vdd FILLER_0_1_44/a_124_375# -0.006062f
C3644 FILLER_0_1_12/a_2812_375# vdd -0.014642f
C3645 vdd FILLER_0_11_72/a_5860_472# 0.009498f
C3646 FILLER_0_10_12/a_1380_472# FILLER_0_9_2/a_2364_375# 0.001543f
C3647 _12_/I _04_/ZN 0.024687f
C3648 _12_/I FILLER_0_7_2/a_2364_375# 0.006134f
C3649 _13_/I FILLER_0_6_37/a_4964_472# 0.003818f
C3650 _18_/I FILLER_0_14_37/a_484_472# 0.001526f
C3651 _13_/Z vdd 0.376215f
C3652 FILLER_0_2_37/a_1916_375# _10_/I 0.001695f
C3653 input_signal[2] FILLER_0_3_12/a_124_375# 0.013212f
C3654 FILLER_0_11_72/a_2812_375# vdd 0.01985f
C3655 output12/a_224_472# _06_/ZN 0.062433f
C3656 FILLER_0_15_72/a_36_472# _19_/I 0.001811f
C3657 FILLER_0_14_28/a_36_472# FILLER_0_12_28/a_124_375# 0.0027f
C3658 _15_/I FILLER_0_10_107/a_572_375# 0.018729f
C3659 FILLER_0_6_37/a_5412_472# _14_/I 0.001219f
C3660 FILLER_0_0_36/a_124_375# _10_/I 0.015932f
C3661 FILLER_0_14_107/a_36_472# FILLER_0_12_107/a_124_375# 0.001512f
C3662 FILLER_0_14_37/a_4964_472# FILLER_0_13_72/a_1020_375# 0.001597f
C3663 FILLER_0_6_2/a_2812_375# _12_/I 0.016091f
C3664 _10_/Z _18_/Z 0.054871f
C3665 FILLER_0_8_37/a_5860_472# vdd 0.008331f
C3666 output_signal_minus[1] _14_/Z 0.080696f
C3667 FILLER_0_14_12/a_484_472# input_signal[7] 0.001645f
C3668 FILLER_0_12_37/a_6396_375# FILLER_0_13_72/a_2364_375# 0.026339f
C3669 _15_/I FILLER_0_11_2/a_1380_472# 0.005458f
C3670 FILLER_0_2_107/a_1468_375# output_signal_minus[8] 0.06111f
C3671 FILLER_0_2_37/a_1020_375# _10_/I 0.001886f
C3672 FILLER_0_0_104/a_36_472# output20/a_224_472# 0.003176f
C3673 FILLER_0_6_2/a_2724_472# FILLER_0_5_12/a_1468_375# 0.001543f
C3674 FILLER_0_6_37/a_3172_472# _12_/I 0.017477f
C3675 FILLER_0_8_37/a_6308_472# FILLER_0_6_37/a_6396_375# 0.001512f
C3676 _00_/ZN output_signal_plus[6] 0.058952f
C3677 FILLER_0_12_37/a_1828_472# _16_/I 0.017477f
C3678 FILLER_0_9_2/a_1020_375# vdd 0.022339f
C3679 output11/a_224_472# FILLER_0_2_37/a_6844_375# 0.001597f
C3680 FILLER_0_10_12/a_124_375# vdd 0.032635f
C3681 _14_/I vdd 2.279909f
C3682 FILLER_0_9_2/a_6756_472# _14_/I 0.004017f
C3683 input10/a_36_113# input_signal[7] 0.001014f
C3684 output24/a_224_472# output23/a_224_472# 0.005335f
C3685 FILLER_0_9_72/a_2724_472# FILLER_0_10_37/a_6756_472# 0.026657f
C3686 _11_/I FILLER_0_3_60/a_572_375# 0.008393f
C3687 FILLER_0_6_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001723f
C3688 _18_/I FILLER_0_14_37/a_3620_472# 0.001526f
C3689 _14_/I FILLER_0_8_37/a_2276_472# 0.014431f
C3690 _15_/I FILLER_0_9_2/a_4156_375# 0.004676f
C3691 _13_/I FILLER_0_4_107/a_1020_375# 0.002197f
C3692 output_signal_minus[9] vdd 0.03452f
C3693 output12/a_224_472# output_signal_minus[3] 0.005251f
C3694 FILLER_0_5_72/a_3172_472# FILLER_0_7_72/a_3260_375# 0.001512f
C3695 _18_/I FILLER_0_15_72/a_36_472# 0.014431f
C3696 vdd FILLER_0_11_72/a_4964_472# 0.002804f
C3697 FILLER_0_6_37/a_3708_375# _14_/I 0.003099f
C3698 _07_/ZN output_signal_minus[5] 0.149064f
C3699 FILLER_0_15_64/a_124_375# FILLER_0_15_72/a_36_472# 0.009654f
C3700 output25/a_224_472# FILLER_0_11_72/a_6756_472# 0.038484f
C3701 _13_/Z output13/a_224_472# 0.077824f
C3702 FILLER_0_10_37/a_4516_472# FILLER_0_8_37/a_4604_375# 0.001512f
C3703 FILLER_0_4_37/a_36_472# FILLER_0_4_2/a_3172_472# 0.002765f
C3704 output14/a_224_472# net15 0.16627f
C3705 FILLER_0_13_72/a_572_375# FILLER_0_12_37/a_4516_472# 0.001723f
C3706 _16_/I FILLER_0_13_2/a_4516_472# 0.004669f
C3707 _15_/I FILLER_0_11_72/a_4516_472# 0.005458f
C3708 FILLER_0_4_37/a_2276_472# vdd 0.036902f
C3709 FILLER_0_13_2/a_6756_472# _16_/I 0.004669f
C3710 _17_/I output_signal_plus[6] 0.419279f
C3711 _16_/I FILLER_0_14_37/a_4068_472# 0.001522f
C3712 _17_/I FILLER_0_14_37/a_6396_375# 0.018729f
C3713 _17_/I FILLER_0_14_37/a_4604_375# 0.018729f
C3714 FILLER_0_1_12/a_2724_472# vdd 0.002467f
C3715 FILLER_0_6_2/a_1380_472# FILLER_0_5_12/a_124_375# 0.001543f
C3716 _12_/I FILLER_0_5_104/a_124_375# 0.001706f
C3717 _18_/I FILLER_0_14_37/a_6308_472# 0.001526f
C3718 _17_/I FILLER_0_15_40/a_124_375# 0.006589f
C3719 _17_/I FILLER_0_15_40/a_484_472# 0.004125f
C3720 _08_/ZN output16/a_224_472# 0.087095f
C3721 FILLER_0_6_2/a_1380_472# vdd 0.010848f
C3722 FILLER_0_13_2/a_6844_375# _17_/I 0.006125f
C3723 vdd FILLER_0_13_2/a_3620_472# 0.007261f
C3724 FILLER_0_9_72/a_1468_375# _14_/I 0.005381f
C3725 output18/a_224_472# FILLER_0_0_104/a_124_375# 0.01196f
C3726 FILLER_0_2_37/a_5412_472# FILLER_0_3_72/a_1468_375# 0.001723f
C3727 FILLER_0_12_107/a_484_472# _09_/ZN 0.003007f
C3728 FILLER_0_10_37/a_2364_375# FILLER_0_9_2/a_6308_472# 0.001597f
C3729 FILLER_0_15_40/a_1020_375# vdd 0.008714f
C3730 FILLER_0_0_36/a_572_375# vdd -0.013067f
C3731 FILLER_0_3_72/a_484_472# FILLER_0_4_37/a_4516_472# 0.026657f
C3732 FILLER_0_1_12/a_1020_375# _10_/I 0.008103f
C3733 _17_/Z _15_/Z 0.007036f
C3734 _15_/I FILLER_0_10_107/a_124_375# 0.01888f
C3735 FILLER_0_8_28/a_124_375# FILLER_0_9_2/a_3172_472# 0.001684f
C3736 _14_/I output13/a_224_472# 0.130298f
C3737 FILLER_0_9_2/a_484_472# FILLER_0_11_2/a_572_375# 0.0027f
C3738 FILLER_0_5_12/a_36_472# vdd 0.015781f
C3739 FILLER_0_6_37/a_6844_375# _14_/I 0.003099f
C3740 FILLER_0_6_37/a_6756_472# vdd 0.014295f
C3741 vdd FILLER_0_6_2/a_2724_472# 0.008883f
C3742 FILLER_0_1_60/a_572_375# _10_/I 0.008103f
C3743 FILLER_0_6_37/a_6396_375# _12_/I 0.016091f
C3744 vdd FILLER_0_12_28/a_36_472# 0.097355f
C3745 _15_/I _14_/a_36_113# 0.004083f
C3746 output17/a_224_472# _14_/I 0.002386f
C3747 FILLER_0_2_37/a_4516_472# _10_/I 0.001843f
C3748 FILLER_0_13_72/a_3260_375# _17_/I 0.006125f
C3749 vdd FILLER_0_3_12/a_1828_472# 0.008796f
C3750 FILLER_0_11_2/a_4964_472# FILLER_0_10_37/a_1020_375# 0.001723f
C3751 FILLER_0_8_37/a_484_472# FILLER_0_6_37/a_572_375# 0.001512f
C3752 FILLER_0_12_101/a_124_375# FILLER_0_14_101/a_36_472# 0.001512f
C3753 FILLER_0_12_37/a_4604_375# vdd 0.004123f
C3754 FILLER_0_7_2/a_6308_472# FILLER_0_6_37/a_2364_375# 0.001723f
C3755 input10/a_36_113# _19_/I 0.003449f
C3756 vdd FILLER_0_13_2/a_2276_472# 0.013919f
C3757 FILLER_0_11_2/a_5948_375# vdd 0.032266f
C3758 FILLER_0_4_2/a_1020_375# FILLER_0_6_2/a_932_472# 0.0027f
C3759 FILLER_0_12_37/a_36_472# FILLER_0_10_37/a_124_375# 0.001512f
C3760 FILLER_0_3_104/a_484_472# FILLER_0_2_107/a_124_375# 0.001723f
C3761 _18_/I FILLER_0_15_56/a_124_375# 0.01418f
C3762 FILLER_0_14_115/a_124_375# vdd 0.020723f
C3763 FILLER_0_12_107/a_1468_375# vdd 0.020319f
C3764 FILLER_0_4_37/a_5052_375# FILLER_0_5_72/a_1020_375# 0.026339f
C3765 FILLER_0_6_37/a_2812_375# vdd 0.009304f
C3766 output11/a_224_472# _10_/I 0.050446f
C3767 FILLER_0_7_2/a_4156_375# _12_/I 0.006193f
C3768 FILLER_0_0_12/a_1380_472# _10_/I 0.016187f
C3769 _19_/a_36_113# output_signal_plus[8] 0.01001f
C3770 _16_/I FILLER_0_12_37/a_1916_375# 0.016091f
C3771 FILLER_0_12_12/a_1468_375# _16_/I 0.016091f
C3772 _09_/ZN FILLER_0_11_72/a_5860_472# 0.017841f
C3773 FILLER_0_2_2/a_3260_375# vdd 0.043165f
C3774 _09_/ZN _13_/Z 0.13814f
C3775 FILLER_0_2_2/a_1380_472# _10_/I 0.002545f
C3776 FILLER_0_4_2/a_484_472# _11_/I 0.017918f
C3777 _11_/I FILLER_0_5_72/a_2812_375# 0.003717f
C3778 FILLER_0_6_107/a_124_375# vdd 0.030073f
C3779 FILLER_0_14_12/a_484_472# _18_/I 0.001526f
C3780 FILLER_0_2_107/a_1020_375# vdd 0.002032f
C3781 _00_/ZN _04_/ZN 0.011799f
C3782 FILLER_0_7_2/a_2276_472# _14_/I 0.008733f
C3783 _19_/I FILLER_0_16_18/a_484_472# 0.014431f
C3784 _13_/I FILLER_0_5_72/a_2364_375# 0.016091f
C3785 output_signal_minus[8] _10_/I 0.038812f
C3786 FILLER_0_0_36/a_2364_375# _10_/I 0.015932f
C3787 FILLER_0_8_28/a_36_472# FILLER_0_8_12/a_1380_472# 0.013277f
C3788 _11_/I FILLER_0_5_72/a_1828_472# 0.001913f
C3789 FILLER_0_6_37/a_1380_472# FILLER_0_5_44/a_572_375# 0.001597f
C3790 _19_/I FILLER_0_15_8/a_484_472# 0.002002f
C3791 FILLER_0_9_72/a_572_375# _14_/I 0.005381f
C3792 FILLER_0_11_72/a_36_472# FILLER_0_11_66/a_124_375# 0.016748f
C3793 FILLER_0_9_72/a_1916_375# FILLER_0_7_72/a_1828_472# 0.001512f
C3794 FILLER_0_0_70/a_124_375# FILLER_0_2_37/a_3620_472# 0.001188f
C3795 FILLER_0_8_37/a_5412_472# vdd 0.006451f
C3796 _11_/I FILLER_0_4_37/a_4604_375# 0.01418f
C3797 FILLER_0_6_37/a_5052_375# FILLER_0_8_37/a_4964_472# 0.001512f
C3798 FILLER_0_2_37/a_3260_375# _10_/I 0.001886f
C3799 FILLER_0_2_2/a_3260_375# FILLER_0_3_12/a_2276_472# 0.001684f
C3800 _03_/ZN _11_/a_36_113# 0.010162f
C3801 _11_/Z FILLER_0_11_72/a_5500_375# 0.001101f
C3802 FILLER_0_7_72/a_1020_375# FILLER_0_5_72/a_932_472# 0.001512f
C3803 _09_/ZN _14_/I 0.074384f
C3804 _18_/I _19_/I 1.858695f
C3805 output14/a_224_472# output_signal_minus[4] 0.076067f
C3806 FILLER_0_3_44/a_1380_472# vdd 0.043709f
C3807 output_signal_plus[7] _10_/Z 0.368064f
C3808 _16_/I FILLER_0_13_2/a_5412_472# 0.004669f
C3809 FILLER_0_11_66/a_124_375# vdd 0.042248f
C3810 _13_/I FILLER_0_6_37/a_1828_472# 0.003818f
C3811 FILLER_0_11_2/a_5412_472# _16_/I 0.007542f
C3812 vdd FILLER_0_10_37/a_5500_375# 0.008584f
C3813 FILLER_0_8_12/a_1468_375# FILLER_0_9_2/a_2724_472# 0.001684f
C3814 _11_/I FILLER_0_4_2/a_2812_375# 0.01418f
C3815 FILLER_0_9_2/a_5052_375# _14_/I 0.005381f
C3816 _18_/I FILLER_0_16_18/a_484_472# 0.002853f
C3817 _09_/ZN FILLER_0_11_72/a_4964_472# 0.008573f
C3818 FILLER_0_11_2/a_3620_472# FILLER_0_13_2/a_3708_375# 0.0027f
C3819 output25/a_224_472# output26/a_224_472# 0.005408f
C3820 _15_/I output24/a_224_472# 0.17689f
C3821 _15_/I FILLER_0_9_2/a_5948_375# 0.006125f
C3822 FILLER_0_7_72/a_3260_375# _12_/I 0.006182f
C3823 vdd output16/a_224_472# 0.14761f
C3824 FILLER_0_8_37/a_3172_472# FILLER_0_6_37/a_3260_375# 0.001512f
C3825 FILLER_0_0_142/a_572_375# _13_/I 0.003279f
C3826 _18_/I FILLER_0_15_8/a_484_472# 0.020978f
C3827 FILLER_0_2_2/a_2364_375# FILLER_0_3_12/a_1380_472# 0.001684f
C3828 FILLER_0_13_104/a_572_375# vdd 0.021013f
C3829 FILLER_0_5_12/a_572_375# _12_/I 0.003304f
C3830 _17_/I FILLER_0_13_2/a_2724_472# 0.00656f
C3831 input_signal[2] input3/a_36_113# 0.060061f
C3832 FILLER_0_4_2/a_1380_472# _12_/I 0.002217f
C3833 output26/a_224_472# output28/a_224_472# 0.072646f
C3834 FILLER_0_9_72/a_1468_375# FILLER_0_8_37/a_5412_472# 0.001723f
C3835 FILLER_0_2_37/a_124_375# FILLER_0_3_12/a_2812_375# 0.026339f
C3836 FILLER_0_5_12/a_1828_472# FILLER_0_4_2/a_2812_375# 0.001684f
C3837 FILLER_0_1_60/a_124_375# FILLER_0_1_44/a_1468_375# 0.012222f
C3838 output17/a_224_472# FILLER_0_2_107/a_1020_375# 0.001597f
C3839 FILLER_0_4_37/a_6308_472# FILLER_0_3_72/a_2276_472# 0.026657f
C3840 FILLER_0_15_64/a_124_375# _18_/I 0.014423f
C3841 _07_/ZN _10_/a_36_160# 0.007113f
C3842 vdd output20/a_224_472# 0.077827f
C3843 FILLER_0_4_37/a_1828_472# FILLER_0_2_37/a_1916_375# 0.001512f
C3844 FILLER_0_14_37/a_5412_472# FILLER_0_13_72/a_1380_472# 0.026657f
C3845 _17_/I FILLER_0_13_2/a_1468_375# 0.006125f
C3846 input_signal[6] FILLER_0_13_2/a_124_375# 0.035039f
C3847 _12_/Z _15_/Z 0.007766f
C3848 _11_/I FILLER_0_3_12/a_3172_472# 0.008683f
C3849 _15_/I FILLER_0_8_37/a_5500_375# 0.002388f
C3850 FILLER_0_2_37/a_6844_375# _10_/I 0.001886f
C3851 FILLER_0_7_2/a_5500_375# _14_/I 0.008393f
C3852 FILLER_0_4_37/a_2276_472# FILLER_0_3_44/a_1468_375# 0.001597f
C3853 FILLER_0_3_44/a_572_375# FILLER_0_2_37/a_1380_472# 0.001723f
C3854 FILLER_0_8_37/a_2812_375# FILLER_0_9_2/a_6844_375# 0.026339f
C3855 FILLER_0_8_37/a_1468_375# FILLER_0_10_37/a_1380_472# 0.001512f
C3856 _18_/I FILLER_0_14_12/a_1468_375# 0.003935f
C3857 output_signal_plus[7] FILLER_0_14_115/a_36_472# 0.001892f
C3858 FILLER_0_11_72/a_2276_472# _15_/I 0.005458f
C3859 vdd FILLER_0_12_37/a_932_472# 0.005474f
C3860 FILLER_0_7_72/a_3172_472# FILLER_0_8_101/a_36_472# 0.026657f
C3861 FILLER_0_7_2/a_1468_375# _12_/I 0.006134f
C3862 input_signal[5] FILLER_0_9_2/a_1020_375# 0.001965f
C3863 _07_/ZN output_signal_minus[3] 0.094076f
C3864 _14_/I FILLER_0_9_2/a_2724_472# 0.004017f
C3865 _15_/I FILLER_0_10_37/a_932_472# 0.015502f
C3866 FILLER_0_2_2/a_1828_472# _11_/I 0.002292f
C3867 _11_/I FILLER_0_5_60/a_572_375# 0.004712f
C3868 FILLER_0_6_2/a_484_472# _14_/I 0.001099f
C3869 _11_/I FILLER_0_2_37/a_3620_472# 0.002415f
C3870 FILLER_0_15_8/a_1916_375# _17_/I 0.006523f
C3871 _15_/I FILLER_0_11_2/a_5860_472# 0.004815f
C3872 _15_/I FILLER_0_9_2/a_4068_472# 0.0029f
C3873 input_signal[5] FILLER_0_10_12/a_124_375# 0.006359f
C3874 input_signal[5] _14_/I 0.002261f
C3875 _18_/a_36_113# _19_/I 0.009548f
C3876 FILLER_0_14_115/a_124_375# _09_/ZN 0.029414f
C3877 FILLER_0_12_107/a_1468_375# _09_/ZN 0.047331f
C3878 output23/a_224_472# _08_/ZN 0.079965f
C3879 FILLER_0_1_12/a_2812_375# FILLER_0_0_36/a_124_375# 0.058411f
C3880 _11_/I FILLER_0_4_2/a_1828_472# 0.014933f
C3881 _19_/a_36_113# _19_/Z 0.007578f
C3882 output17/a_224_472# output16/a_224_472# 0.072646f
C3883 FILLER_0_11_2/a_36_472# vdd 0.105578f
C3884 _11_/I output_signal_plus[2] 0.001778f
C3885 FILLER_0_5_44/a_124_375# vdd 0.010906f
C3886 FILLER_0_6_107/a_124_375# _09_/ZN 0.001551f
C3887 FILLER_0_12_12/a_124_375# _16_/I 0.016409f
C3888 input8/a_36_113# input_signal[9] 0.001325f
C3889 FILLER_0_12_12/a_1020_375# FILLER_0_13_2/a_2276_472# 0.001684f
C3890 _13_/Z output_signal_minus[2] 0.102232f
C3891 _09_/ZN FILLER_0_2_107/a_1020_375# 0.029277f
C3892 _16_/I FILLER_0_11_2/a_2812_375# 0.007169f
C3893 _15_/I FILLER_0_11_72/a_6396_375# 0.005476f
C3894 input_signal[2] _12_/I 0.065697f
C3895 _11_/I FILLER_0_5_12/a_3172_472# 0.001913f
C3896 FILLER_0_4_101/a_36_472# FILLER_0_4_107/a_36_472# 0.003468f
C3897 FILLER_0_3_104/a_572_375# vdd 0.018731f
C3898 FILLER_0_7_2/a_6308_472# FILLER_0_8_37/a_2364_375# 0.001597f
C3899 _13_/I FILLER_0_5_72/a_1380_472# 0.017477f
C3900 _17_/I FILLER_0_15_40/a_572_375# 0.006589f
C3901 FILLER_0_5_72/a_1468_375# _12_/I 0.001706f
C3902 _16_/I FILLER_0_11_72/a_1380_472# 0.00753f
C3903 vdd FILLER_0_6_2/a_1828_472# 0.0419f
C3904 FILLER_0_2_37/a_36_472# FILLER_0_3_12/a_2812_375# 0.001723f
C3905 FILLER_0_3_72/a_1916_375# FILLER_0_2_37/a_5860_472# 0.001723f
C3906 _17_/I FILLER_0_13_2/a_2812_375# 0.006125f
C3907 _18_/I _18_/a_36_113# 0.017913f
C3908 FILLER_0_13_72/a_2276_472# output29/a_224_472# 0.001243f
C3909 vdd FILLER_0_11_2/a_4516_472# 0.005419f
C3910 FILLER_0_11_136/a_36_472# _10_/Z 0.004421f
C3911 FILLER_0_6_37/a_2364_375# vdd 0.027535f
C3912 FILLER_0_13_2/a_1020_375# vdd 0.022339f
C3913 _17_/I FILLER_0_13_2/a_3708_375# 0.00471f
C3914 FILLER_0_5_44/a_572_375# _13_/I 0.016091f
C3915 FILLER_0_14_12/a_124_375# input_signal[7] 0.005639f
C3916 _14_/I output_signal_minus[2] 0.249844f
C3917 _12_/Z output_signal_plus[1] 0.023126f
C3918 _13_/I FILLER_0_5_72/a_2724_472# 0.017477f
C3919 FILLER_0_10_37/a_4068_472# vdd 0.002855f
C3920 FILLER_0_6_37/a_2364_375# FILLER_0_8_37/a_2276_472# 0.001512f
C3921 output18/a_224_472# FILLER_0_0_104/a_36_472# 0.003196f
C3922 FILLER_0_4_37/a_484_472# vdd 0.004055f
C3923 _13_/I FILLER_0_5_44/a_36_472# 0.017477f
C3924 output22/a_224_472# FILLER_0_9_104/a_572_375# 0.011584f
C3925 FILLER_0_5_12/a_36_472# input_signal[3] 0.073201f
C3926 _16_/I FILLER_0_10_107/a_572_375# 0.00231f
C3927 vdd output_signal_plus[0] 0.123495f
C3928 _15_/Z output26/a_224_472# 0.034465f
C3929 FILLER_0_9_2/a_3708_375# _14_/I 0.005433f
C3930 _10_/Z output14/a_224_472# 0.056447f
C3931 _09_/ZN FILLER_0_13_104/a_572_375# 0.002462f
C3932 output_signal_minus[5] _04_/ZN 0.020416f
C3933 FILLER_0_15_64/a_36_472# FILLER_0_15_72/a_36_472# 0.002296f
C3934 _17_/I _18_/Z 0.015713f
C3935 _16_/I FILLER_0_11_2/a_1380_472# 0.007596f
C3936 output_signal_minus[1] _06_/ZN 0.0113f
C3937 FILLER_0_10_12/a_36_472# input6/a_36_113# 0.001663f
C3938 FILLER_0_0_12/a_124_375# _10_/I 0.017538f
C3939 FILLER_0_8_37/a_5948_375# FILLER_0_10_37/a_5860_472# 0.001512f
C3940 _16_/I FILLER_0_12_37/a_2276_472# 0.017477f
C3941 _11_/I FILLER_0_2_37/a_4156_375# 0.002629f
C3942 FILLER_0_9_72/a_1380_472# _14_/I 0.004017f
C3943 FILLER_0_1_12/a_484_472# FILLER_0_2_2/a_1468_375# 0.001543f
C3944 FILLER_0_7_2/a_124_375# FILLER_0_6_2/a_124_375# 0.05841f
C3945 FILLER_0_3_12/a_3260_375# vdd 0.005129f
C3946 output_signal_plus[8] vdd 0.659222f
C3947 FILLER_0_12_101/a_124_375# _17_/I 0.002388f
C3948 FILLER_0_9_2/a_1916_375# FILLER_0_10_12/a_932_472# 0.001543f
C3949 output11/a_224_472# FILLER_0_2_37/a_6396_375# 0.001597f
C3950 _13_/I FILLER_0_6_101/a_124_375# 0.002413f
C3951 FILLER_0_3_44/a_1020_375# FILLER_0_2_37/a_1828_472# 0.001723f
C3952 FILLER_0_6_37/a_1468_375# _12_/I 0.016091f
C3953 FILLER_0_7_72/a_36_472# vdd 0.108637f
C3954 output23/a_224_472# vdd 0.147266f
C3955 FILLER_0_14_37/a_6756_472# FILLER_0_12_37/a_6844_375# 0.001512f
C3956 output_signal_minus[1] output_signal_minus[3] 0.004865f
C3957 _16_/I FILLER_0_11_72/a_4516_472# 0.005646f
C3958 vdd FILLER_0_9_104/a_124_375# 0.027844f
C3959 _11_/I FILLER_0_4_37/a_1020_375# 0.01418f
C3960 vdd FILLER_0_15_8/a_1828_472# 0.010564f
C3961 _17_/I FILLER_0_15_72/a_1020_375# 0.006589f
C3962 FILLER_0_15_8/a_3260_375# _17_/I 0.006589f
C3963 FILLER_0_4_37/a_6308_472# FILLER_0_2_37/a_6396_375# 0.001512f
C3964 FILLER_0_7_2/a_6756_472# FILLER_0_9_2/a_6844_375# 0.001512f
C3965 FILLER_0_15_8/a_3172_472# _18_/I 0.014431f
C3966 output24/a_224_472# FILLER_0_10_107/a_1468_375# 0.009867f
C3967 vdd FILLER_0_14_107/a_572_375# 0.004919f
C3968 FILLER_0_10_37/a_5052_375# FILLER_0_11_72/a_1020_375# 0.026339f
C3969 FILLER_0_10_37/a_1020_375# FILLER_0_12_37/a_932_472# 0.001512f
C3970 _11_/I FILLER_0_5_12/a_2276_472# 0.001913f
C3971 output18/a_224_472# _08_/ZN 0.020259f
C3972 _11_/I FILLER_0_3_72/a_1380_472# 0.008683f
C3973 FILLER_0_13_72/a_1828_472# vdd 0.00902f
C3974 _17_/I FILLER_0_14_37/a_5412_472# 0.015502f
C3975 FILLER_0_12_37/a_5860_472# FILLER_0_10_37/a_5948_375# 0.001512f
C3976 FILLER_0_5_44/a_124_375# FILLER_0_4_37/a_932_472# 0.001723f
C3977 FILLER_0_10_107/a_124_375# _16_/I 0.002327f
C3978 FILLER_0_2_2/a_1020_375# vdd 0.022339f
C3979 _15_/I _08_/ZN 0.094861f
C3980 FILLER_0_13_2/a_5412_472# FILLER_0_14_37/a_1380_472# 0.026657f
C3981 _11_/I FILLER_0_5_12/a_1916_375# 0.004745f
C3982 FILLER_0_7_2/a_1828_472# vdd 0.046351f
C3983 FILLER_0_11_72/a_6844_375# _16_/I 0.005677f
C3984 FILLER_0_4_2/a_2724_472# FILLER_0_3_12/a_1468_375# 0.001543f
C3985 _09_/ZN FILLER_0_3_104/a_572_375# 0.018071f
C3986 vdd FILLER_0_6_37/a_5860_472# 0.007851f
C3987 FILLER_0_6_101/a_36_472# vdd 0.097837f
C3988 vdd FILLER_0_11_72/a_4068_472# 0.005722f
C3989 FILLER_0_6_37/a_484_472# _12_/I 0.017477f
C3990 FILLER_0_12_107/a_572_375# _16_/I 0.016091f
C3991 FILLER_0_13_2/a_6308_472# FILLER_0_12_37/a_2364_375# 0.001723f
C3992 FILLER_0_9_66/a_36_472# vdd 0.097097f
C3993 _12_/I FILLER_0_7_2/a_1916_375# 0.002227f
C3994 FILLER_0_15_40/a_36_472# vdd 0.084762f
C3995 _18_/I FILLER_0_14_12/a_124_375# 0.003935f
C3996 FILLER_0_9_2/a_4964_472# _14_/I 0.004017f
C3997 FILLER_0_9_66/a_36_472# FILLER_0_9_2/a_6756_472# 0.013276f
C3998 FILLER_0_6_37/a_484_472# FILLER_0_4_37/a_572_375# 0.001512f
C3999 output23/a_224_472# output13/a_224_472# 0.09755f
C4000 input_signal[0] FILLER_0_0_12/a_932_472# 0.001215f
C4001 FILLER_0_0_104/a_124_375# output_signal_minus[0] 0.017182f
C4002 FILLER_0_1_44/a_932_472# _10_/I 0.006408f
C4003 _11_/I FILLER_0_3_72/a_1020_375# 0.008393f
C4004 _14_/I output_signal_minus[8] 0.370182f
C4005 FILLER_0_3_72/a_2724_472# vdd 0.034108f
C4006 output_signal_minus[7] output_signal_minus[6] 0.214325f
C4007 FILLER_0_2_2/a_1916_375# FILLER_0_4_2/a_1828_472# 0.0027f
C4008 input8/a_36_113# input7/a_36_113# 0.001442f
C4009 FILLER_0_11_2/a_4068_472# vdd 0.002735f
C4010 FILLER_0_6_2/a_1380_472# FILLER_0_4_2/a_1468_375# 0.0027f
C4011 output_signal_minus[9] output_signal_minus[8] 0.328708f
C4012 _17_/I FILLER_0_12_107/a_124_375# 0.002388f
C4013 _00_/ZN output_signal_plus[7] 0.006625f
C4014 FILLER_0_15_64/a_36_472# _19_/I 0.001641f
C4015 _13_/I FILLER_0_5_72/a_2276_472# 0.017477f
C4016 FILLER_0_1_12/a_2276_472# vdd 0.007367f
C4017 _11_/I FILLER_0_5_12/a_1828_472# 0.001913f
C4018 FILLER_0_10_12/a_1468_375# vdd 0.023715f
C4019 FILLER_0_2_37/a_4604_375# FILLER_0_4_37/a_4516_472# 0.001512f
C4020 FILLER_0_12_37/a_124_375# FILLER_0_13_2/a_4156_375# 0.026339f
C4021 _14_/Z _15_/a_36_113# 0.074239f
C4022 _15_/I FILLER_0_10_101/a_124_375# 0.019472f
C4023 vdd FILLER_0_8_37/a_2364_375# 0.027463f
C4024 FILLER_0_4_2/a_2364_375# FILLER_0_3_12/a_1380_472# 0.001543f
C4025 vdd FILLER_0_5_72/a_572_375# 0.002455f
C4026 _12_/I FILLER_0_5_72/a_1020_375# 0.001706f
C4027 output15/a_224_472# output14/a_224_472# 0.061459f
C4028 FILLER_0_4_101/a_36_472# FILLER_0_5_72/a_3260_375# 0.001723f
C4029 output25/a_224_472# FILLER_0_11_72/a_6308_472# 0.038484f
C4030 FILLER_0_6_37/a_4964_472# FILLER_0_5_72/a_932_472# 0.026657f
C4031 _15_/I FILLER_0_12_37/a_3172_472# 0.001368f
C4032 FILLER_0_6_37/a_6844_375# FILLER_0_6_101/a_36_472# 0.086635f
C4033 input_signal[5] FILLER_0_11_2/a_36_472# 0.002659f
C4034 FILLER_0_14_28/a_36_472# FILLER_0_14_12/a_1380_472# 0.013276f
C4035 _19_/Z vdd 0.461606f
C4036 FILLER_0_2_107/a_1468_375# _14_/I 0.042058f
C4037 _06_/ZN _04_/ZN 0.383359f
C4038 FILLER_0_14_37/a_4156_375# vdd 0.004458f
C4039 output_signal_plus[7] _17_/I 0.077237f
C4040 FILLER_0_0_12/a_1468_375# FILLER_0_0_28/a_36_472# 0.086635f
C4041 FILLER_0_5_44/a_1020_375# FILLER_0_4_37/a_1828_472# 0.001723f
C4042 FILLER_0_15_64/a_36_472# _18_/I 0.014431f
C4043 vdd FILLER_0_14_37/a_124_375# 0.015736f
C4044 FILLER_0_8_37/a_6756_472# FILLER_0_8_101/a_36_472# 0.013277f
C4045 FILLER_0_6_37/a_1380_472# vdd 0.007218f
C4046 _15_/I FILLER_0_11_72/a_36_472# 0.005458f
C4047 output24/a_224_472# _16_/I 0.010638f
C4048 FILLER_0_10_37/a_572_375# vdd 0.005046f
C4049 FILLER_0_14_37/a_3260_375# vdd 0.008684f
C4050 FILLER_0_13_2/a_932_472# _17_/I 0.005193f
C4051 output18/a_224_472# vdd 0.009481f
C4052 FILLER_0_11_2/a_6308_472# FILLER_0_10_37/a_2364_375# 0.001723f
C4053 FILLER_0_2_37/a_124_375# FILLER_0_4_37/a_36_472# 0.001512f
C4054 FILLER_0_6_107/a_36_472# FILLER_0_5_104/a_484_472# 0.026657f
C4055 _10_/Z _01_/ZN 0.293785f
C4056 FILLER_0_11_136/a_36_472# output_signal_plus[4] 0.001108f
C4057 vdd FILLER_0_6_2/a_36_472# 0.105578f
C4058 vdd FILLER_0_5_60/a_124_375# 0.014393f
C4059 _15_/I vdd 2.230738f
C4060 _11_/I FILLER_0_4_2/a_572_375# 0.017531f
C4061 FILLER_0_9_2/a_6756_472# _15_/I 0.006506f
C4062 FILLER_0_3_72/a_124_375# FILLER_0_4_37/a_4068_472# 0.001597f
C4063 FILLER_0_15_72/a_1380_472# _17_/I 0.004125f
C4064 FILLER_0_4_2/a_3260_375# FILLER_0_5_12/a_2276_472# 0.001684f
C4065 _16_/I FILLER_0_14_37/a_1828_472# 0.001667f
C4066 FILLER_0_11_2/a_1916_375# FILLER_0_10_12/a_932_472# 0.001684f
C4067 output_signal_minus[3] _04_/ZN 0.004026f
C4068 output22/a_224_472# _13_/Z 0.220782f
C4069 input8/a_36_113# _17_/I 0.008318f
C4070 FILLER_0_12_12/a_36_472# FILLER_0_10_12/a_124_375# 0.0027f
C4071 FILLER_0_8_37/a_3708_375# FILLER_0_10_37/a_3620_472# 0.0027f
C4072 FILLER_0_2_37/a_932_472# FILLER_0_1_44/a_36_472# 0.026657f
C4073 _16_/I FILLER_0_13_2/a_4964_472# 0.004669f
C4074 _13_/I _08_/ZN 0.098939f
C4075 FILLER_0_4_2/a_1020_375# _11_/I 0.014773f
C4076 FILLER_0_2_107/a_1020_375# output_signal_minus[8] 0.00945f
C4077 FILLER_0_3_12/a_36_472# FILLER_0_5_12/a_124_375# 0.0027f
C4078 input_signal[2] FILLER_0_4_2/a_124_375# 0.003817f
C4079 FILLER_0_11_72/a_1828_472# FILLER_0_12_37/a_5860_472# 0.026657f
C4080 _16_/I FILLER_0_12_37/a_5052_375# 0.016091f
C4081 vdd FILLER_0_3_12/a_36_472# 0.015685f
C4082 vdd FILLER_0_2_101/a_124_375# 0.044083f
C4083 input6/a_36_113# input7/a_36_113# 0.001442f
C4084 FILLER_0_11_72/a_2276_472# _16_/I 0.00753f
C4085 _09_/ZN FILLER_0_11_72/a_4068_472# 0.001875f
C4086 FILLER_0_9_72/a_1468_375# _15_/I 0.006125f
C4087 _11_/I FILLER_0_4_2/a_3260_375# 0.014327f
C4088 FILLER_0_14_37/a_6756_472# FILLER_0_14_101/a_36_472# 0.013277f
C4089 FILLER_0_0_12/a_484_472# vdd 0.016427f
C4090 _12_/I FILLER_0_6_37/a_572_375# 0.016091f
C4091 _13_/I FILLER_0_4_37/a_5500_375# 0.005726f
C4092 _16_/I FILLER_0_11_2/a_5860_472# 0.007542f
C4093 output22/a_224_472# _14_/I 0.007248f
C4094 FILLER_0_0_70/a_36_472# _10_/I 0.016219f
C4095 _16_/Z _10_/Z 0.099778f
C4096 FILLER_0_1_44/a_124_375# _10_/I 0.008103f
C4097 output19/a_224_472# output14/a_224_472# 0.09755f
C4098 FILLER_0_13_72/a_36_472# vdd 0.108638f
C4099 FILLER_0_9_72/a_1916_375# FILLER_0_10_37/a_5860_472# 0.001597f
C4100 FILLER_0_1_12/a_2812_375# _10_/I 0.008103f
C4101 _19_/I FILLER_0_16_36/a_484_472# 0.014431f
C4102 _13_/I FILLER_0_5_12/a_1468_375# 0.016091f
C4103 FILLER_0_2_37/a_4516_472# output20/a_224_472# 0.001058f
C4104 FILLER_0_7_2/a_5860_472# FILLER_0_6_37/a_1916_375# 0.001723f
C4105 _14_/I FILLER_0_7_72/a_2724_472# 0.009305f
C4106 output17/a_224_472# output18/a_224_472# 0.185233f
C4107 _07_/ZN FILLER_0_11_72/a_6844_375# 0.018746f
C4108 FILLER_0_3_72/a_3260_375# FILLER_0_2_101/a_124_375# 0.026339f
C4109 FILLER_0_7_2/a_4604_375# FILLER_0_6_37/a_572_375# 0.026339f
C4110 FILLER_0_13_2/a_4068_472# FILLER_0_14_37/a_36_472# 0.026657f
C4111 FILLER_0_0_36/a_2276_472# vdd 0.035285f
C4112 output_signal_plus[8] output30/a_224_472# 0.013948f
C4113 FILLER_0_11_2/a_5500_375# vdd 0.011603f
C4114 output_signal_minus[8] output16/a_224_472# 0.011966f
C4115 _14_/I FILLER_0_9_2/a_1468_375# 0.005414f
C4116 FILLER_0_9_104/a_36_472# FILLER_0_9_72/a_3172_472# 0.013276f
C4117 _16_/I FILLER_0_11_72/a_6396_375# 0.005912f
C4118 output11/a_224_472# output20/a_224_472# 0.061459f
C4119 FILLER_0_12_12/a_1468_375# FILLER_0_13_2/a_2724_472# 0.001684f
C4120 _12_/I FILLER_0_5_72/a_3260_375# 0.001706f
C4121 FILLER_0_13_72/a_1916_375# vdd 0.009597f
C4122 FILLER_0_2_37/a_2812_375# vdd 0.011102f
C4123 FILLER_0_5_60/a_36_472# vdd 0.094274f
C4124 FILLER_0_6_2/a_2276_472# _12_/I 0.017477f
C4125 FILLER_0_4_37/a_3620_472# _13_/I 0.003497f
C4126 _18_/I FILLER_0_15_40/a_1020_375# 0.01418f
C4127 FILLER_0_15_2/a_124_375# vdd 0.020228f
C4128 _11_/I FILLER_0_2_2/a_1916_375# 0.003213f
C4129 _00_/ZN output14/a_224_472# 0.001232f
C4130 _18_/I FILLER_0_16_36/a_484_472# 0.001782f
C4131 FILLER_0_14_12/a_1020_375# FILLER_0_15_8/a_1468_375# 0.05841f
C4132 vdd FILLER_0_10_37/a_1468_375# 0.008221f
C4133 vdd FILLER_0_0_28/a_36_472# 0.093232f
C4134 vdd FILLER_0_2_2/a_2364_375# 0.024816f
C4135 FILLER_0_6_37/a_5412_472# _13_/I 0.003818f
C4136 FILLER_0_13_72/a_2364_375# FILLER_0_12_37/a_6308_472# 0.001723f
C4137 output_signal_minus[9] _10_/I 0.15211f
C4138 vdd FILLER_0_6_37/a_4516_472# 0.002735f
C4139 _15_/I FILLER_0_10_37/a_4604_375# 0.018729f
C4140 FILLER_0_14_37/a_2812_375# vdd 0.010526f
C4141 FILLER_0_6_37/a_3260_375# FILLER_0_7_66/a_36_472# 0.001723f
C4142 _14_/I FILLER_0_8_12/a_932_472# 0.014431f
C4143 FILLER_0_9_72/a_572_375# _15_/I 0.003577f
C4144 FILLER_0_0_36/a_484_472# _10_/I 0.016187f
C4145 output23/a_224_472# output_signal_minus[2] 0.007286f
C4146 FILLER_0_2_107/a_1468_375# output16/a_224_472# 0.002622f
C4147 _11_/I _12_/a_36_113# 0.001358f
C4148 FILLER_0_14_115/a_124_375# _18_/I 0.011194f
C4149 vdd FILLER_0_2_37/a_5412_472# 0.007665f
C4150 _13_/I FILLER_0_5_12/a_124_375# 0.01631f
C4151 _11_/I FILLER_0_2_2/a_2276_472# 0.002415f
C4152 FILLER_0_1_12/a_2724_472# _10_/I 0.006408f
C4153 FILLER_0_8_12/a_1468_375# FILLER_0_7_2/a_2724_472# 0.001543f
C4154 _13_/I vdd 1.572923f
C4155 _15_/I _09_/ZN 0.047804f
C4156 FILLER_0_6_37/a_1468_375# FILLER_0_7_2/a_5412_472# 0.001723f
C4157 FILLER_0_8_107/a_484_472# vdd 0.008393f
C4158 FILLER_0_2_37/a_6756_472# FILLER_0_2_101/a_36_472# 0.013277f
C4159 FILLER_0_14_37/a_6844_375# output29/a_224_472# 0.029497f
C4160 FILLER_0_9_104/a_572_375# _14_/I 0.005381f
C4161 vdd input5/a_36_113# 0.121506f
C4162 FILLER_0_0_36/a_572_375# _10_/I 0.015932f
C4163 vdd FILLER_0_9_2/a_484_472# 0.0074f
C4164 _15_/I FILLER_0_9_2/a_5052_375# 0.006125f
C4165 _13_/I FILLER_0_6_37/a_3708_375# 0.001706f
C4166 _12_/I FILLER_0_7_72/a_1380_472# 0.004669f
C4167 FILLER_0_0_104/a_36_472# output_signal_minus[0] 0.032681f
C4168 _14_/I FILLER_0_9_2/a_2276_472# 0.004017f
C4169 _16_/I FILLER_0_13_2/a_3172_472# 0.004669f
C4170 _07_/ZN output24/a_224_472# 0.12199f
C4171 _15_/I FILLER_0_10_37/a_1020_375# 0.018729f
C4172 FILLER_0_10_12/a_1468_375# FILLER_0_9_2/a_2724_472# 0.001543f
C4173 FILLER_0_11_2/a_1828_472# vdd 0.046348f
C4174 FILLER_0_7_2/a_4964_472# FILLER_0_8_37/a_932_472# 0.026657f
C4175 FILLER_0_3_104/a_124_375# _01_/ZN 0.001664f
C4176 FILLER_0_6_101/a_36_472# FILLER_0_4_101/a_124_375# 0.001512f
C4177 output12/a_224_472# _08_/ZN 0.08546f
C4178 FILLER_0_7_72/a_3172_472# FILLER_0_9_72/a_3260_375# 0.001512f
C4179 FILLER_0_7_66/a_124_375# vdd 0.042668f
C4180 FILLER_0_14_37/a_3172_472# vdd 0.007139f
C4181 _13_/I FILLER_0_4_37/a_4156_375# 0.005726f
C4182 output_signal_minus[7] FILLER_0_0_142/a_484_472# 0.002964f
C4183 FILLER_0_6_107/a_36_472# _12_/I 0.020616f
C4184 vdd FILLER_0_3_60/a_36_472# 0.094979f
C4185 FILLER_0_12_12/a_484_472# FILLER_0_11_2/a_1468_375# 0.001543f
C4186 FILLER_0_2_37/a_2364_375# vdd 0.029138f
C4187 _17_/I FILLER_0_12_28/a_124_375# 0.002388f
C4188 FILLER_0_10_37/a_3260_375# FILLER_0_12_37/a_3172_472# 0.001512f
C4189 FILLER_0_2_2/a_3260_375# _10_/I 0.001886f
C4190 FILLER_0_6_37/a_6844_375# _13_/I 0.001944f
C4191 _19_/Z output30/a_224_472# 0.003458f
C4192 output_signal_minus[1] _14_/a_36_113# 0.023164f
C4193 FILLER_0_5_72/a_3172_472# FILLER_0_5_104/a_36_472# 0.013276f
C4194 FILLER_0_7_2/a_2724_472# _14_/I 0.008733f
C4195 _16_/I _08_/ZN 0.226887f
C4196 FILLER_0_13_104/a_124_375# FILLER_0_11_72/a_3620_472# 0.0027f
C4197 FILLER_0_10_107/a_1468_375# vdd 0.018648f
C4198 vdd FILLER_0_9_2/a_3172_472# 0.007993f
C4199 FILLER_0_5_44/a_484_472# _12_/I 0.003805f
C4200 FILLER_0_10_28/a_36_472# FILLER_0_9_2/a_2812_375# 0.001543f
C4201 vdd FILLER_0_0_36/a_932_472# 0.00312f
C4202 _15_/I FILLER_0_9_2/a_2724_472# 0.00656f
C4203 FILLER_0_7_72/a_124_375# _14_/I 0.008393f
C4204 input_signal[5] _15_/I 0.154964f
C4205 output24/a_224_472# FILLER_0_10_107/a_1380_472# 0.001826f
C4206 FILLER_0_8_107/a_124_375# _11_/Z 0.002001f
C4207 FILLER_0_14_107/a_124_375# _17_/I 0.01888f
C4208 _12_/I FILLER_0_6_37/a_3620_472# 0.017477f
C4209 FILLER_0_7_2/a_1380_472# vdd 0.012473f
C4210 input_signal[3] FILLER_0_6_2/a_36_472# 0.021747f
C4211 FILLER_0_2_37/a_1380_472# FILLER_0_1_44/a_572_375# 0.001597f
C4212 _11_/I FILLER_0_4_107/a_1380_472# 0.028098f
C4213 FILLER_0_5_44/a_1468_375# _12_/I 0.001706f
C4214 FILLER_0_12_37/a_572_375# vdd 0.005339f
C4215 FILLER_0_15_56/a_572_375# FILLER_0_14_37/a_2724_472# 0.001723f
C4216 output19/a_224_472# _01_/ZN 0.005567f
C4217 vdd FILLER_0_10_37/a_3260_375# 0.006624f
C4218 FILLER_0_6_37/a_932_472# FILLER_0_4_37/a_1020_375# 0.001512f
C4219 FILLER_0_4_37/a_5412_472# FILLER_0_3_72/a_1468_375# 0.001597f
C4220 FILLER_0_0_36/a_36_472# FILLER_0_0_28/a_36_472# 0.002296f
C4221 _13_/I FILLER_0_5_72/a_36_472# 0.019507f
C4222 _17_/I FILLER_0_12_37/a_5948_375# 0.002388f
C4223 _15_/I FILLER_0_11_2/a_5052_375# 0.007111f
C4224 FILLER_0_7_2/a_6756_472# FILLER_0_8_37/a_2724_472# 0.026657f
C4225 FILLER_0_8_37/a_5860_472# FILLER_0_6_37/a_5948_375# 0.001512f
C4226 _07_/ZN FILLER_0_11_72/a_6396_375# 0.001195f
C4227 vdd FILLER_0_14_37/a_3708_375# 0.021939f
C4228 output16/a_224_472# _10_/I 0.00369f
C4229 input3/a_36_113# input4/a_36_113# 0.001442f
C4230 FILLER_0_14_37/a_5500_375# _17_/I 0.018729f
C4231 FILLER_0_6_37/a_5948_375# _14_/I 0.003099f
C4232 _16_/I FILLER_0_10_101/a_124_375# 0.002327f
C4233 vdd FILLER_0_2_37/a_5948_375# 0.012018f
C4234 _11_/I FILLER_0_3_72/a_2364_375# 0.008393f
C4235 _13_/I FILLER_0_4_37/a_932_472# 0.003497f
C4236 _13_/I _09_/ZN 0.151561f
C4237 _13_/I FILLER_0_5_12/a_2812_375# 0.016091f
C4238 FILLER_0_14_28/a_124_375# FILLER_0_13_2/a_3172_472# 0.001543f
C4239 FILLER_0_13_66/a_124_375# FILLER_0_11_66/a_36_472# 0.001512f
C4240 FILLER_0_10_37/a_2724_472# FILLER_0_8_37/a_2812_375# 0.001512f
C4241 FILLER_0_3_12/a_572_375# vdd 0.053784f
C4242 _15_/I output_signal_minus[2] 0.00664f
C4243 vdd FILLER_0_3_104/a_484_472# 0.00781f
C4244 output20/a_224_472# _10_/I 0.114068f
C4245 FILLER_0_16_36/a_36_472# FILLER_0_16_18/a_1468_375# 0.016748f
C4246 _16_/I FILLER_0_12_37/a_3172_472# 0.017477f
C4247 _00_/ZN _01_/ZN 0.009066f
C4248 _17_/I FILLER_0_13_72/a_2724_472# 0.00652f
C4249 vdd FILLER_0_0_36/a_3172_472# 0.010866f
C4250 FILLER_0_8_12/a_484_472# input_signal[4] 0.001762f
C4251 FILLER_0_12_12/a_36_472# FILLER_0_13_2/a_1020_375# 0.001684f
C4252 output12/a_224_472# vdd 0.137446f
C4253 output_signal_minus[5] output14/a_224_472# 0.001472f
C4254 vdd FILLER_0_8_12/a_36_472# 0.016261f
C4255 _11_/I FILLER_0_3_12/a_2724_472# 0.003282f
C4256 _19_/I output_signal_plus[0] 0.052365f
C4257 FILLER_0_13_104/a_484_472# FILLER_0_14_107/a_36_472# 0.026657f
C4258 FILLER_0_14_37/a_6756_472# _17_/I 0.015502f
C4259 _16_/I FILLER_0_11_72/a_36_472# 0.00753f
C4260 _15_/I FILLER_0_9_2/a_3708_375# 0.00471f
C4261 FILLER_0_6_2/a_3172_472# _12_/I 0.01783f
C4262 FILLER_0_4_37/a_2364_375# vdd 0.028423f
C4263 FILLER_0_9_2/a_4068_472# FILLER_0_10_37/a_36_472# 0.026657f
C4264 FILLER_0_4_37/a_3260_375# FILLER_0_5_60/a_572_375# 0.026339f
C4265 _17_/I FILLER_0_12_37/a_1020_375# 0.002388f
C4266 FILLER_0_13_2/a_1468_375# FILLER_0_11_2/a_1380_472# 0.0027f
C4267 FILLER_0_4_2/a_36_472# _12_/I 0.014911f
C4268 _11_/I FILLER_0_5_12/a_2724_472# 0.001913f
C4269 FILLER_0_3_72/a_1020_375# FILLER_0_1_72/a_932_472# 0.001512f
C4270 _16_/I vdd 1.882731f
C4271 FILLER_0_9_72/a_1380_472# _15_/I 0.00652f
C4272 FILLER_0_8_12/a_1468_375# _14_/I 0.01418f
C4273 output_signal_plus[8] _19_/I 0.068849f
C4274 FILLER_0_11_72/a_1468_375# FILLER_0_10_37/a_5412_472# 0.001723f
C4275 FILLER_0_7_104/a_124_375# _12_/I 0.006313f
C4276 FILLER_0_11_72/a_2364_375# FILLER_0_12_37/a_6308_472# 0.001597f
C4277 FILLER_0_12_101/a_36_472# FILLER_0_10_101/a_124_375# 0.001512f
C4278 FILLER_0_6_37/a_1380_472# FILLER_0_4_37/a_1468_375# 0.001512f
C4279 FILLER_0_4_37/a_4516_472# vdd 0.002735f
C4280 FILLER_0_13_2/a_1828_472# FILLER_0_12_12/a_572_375# 0.001684f
C4281 _18_/I output_signal_plus[0] 0.004162f
C4282 _15_/I FILLER_0_11_72/a_5052_375# 0.007111f
C4283 FILLER_0_2_37/a_3172_472# FILLER_0_1_60/a_484_472# 0.026657f
C4284 FILLER_0_15_72/a_1468_375# FILLER_0_14_37/a_5412_472# 0.001723f
C4285 output25/a_224_472# _10_/Z 0.086381f
C4286 _09_/ZN FILLER_0_10_107/a_1468_375# 0.047331f
C4287 _12_/I input4/a_36_113# 0.019215f
C4288 FILLER_0_10_107/a_36_472# FILLER_0_10_101/a_124_375# 0.016748f
C4289 _12_/I FILLER_0_5_104/a_36_472# 0.003965f
C4290 _17_/Z output26/a_224_472# 0.219393f
C4291 vdd output_signal_minus[0] 0.291987f
C4292 output12/a_224_472# output13/a_224_472# 0.031309f
C4293 _19_/I FILLER_0_15_8/a_1828_472# 0.00191f
C4294 FILLER_0_6_37/a_484_472# FILLER_0_5_12/a_3260_375# 0.001597f
C4295 FILLER_0_4_37/a_1380_472# _13_/I 0.003497f
C4296 _10_/Z output28/a_224_472# 0.099085f
C4297 _13_/I FILLER_0_6_2/a_484_472# 0.005378f
C4298 _13_/Z _14_/I 0.047735f
C4299 _15_/I FILLER_0_11_2/a_484_472# 0.005205f
C4300 _12_/a_36_113# _12_/Z 0.007219f
C4301 output_signal_minus[9] FILLER_0_0_70/a_36_472# 0.002187f
C4302 input_signal[5] input5/a_36_113# 0.005377f
C4303 FILLER_0_6_37/a_4068_472# _12_/I 0.017477f
C4304 _13_/I FILLER_0_5_12/a_932_472# 0.017477f
C4305 _17_/I FILLER_0_14_12/a_36_472# 0.025249f
C4306 _13_/I input_signal[3] 0.176165f
C4307 _18_/I output_signal_plus[8] 0.117587f
C4308 FILLER_0_3_44/a_1468_375# FILLER_0_3_60/a_36_472# 0.086742f
C4309 FILLER_0_2_37/a_2364_375# FILLER_0_3_44/a_1468_375# 0.026339f
C4310 FILLER_0_8_37/a_5860_472# _14_/I 0.014431f
C4311 input_signal[5] FILLER_0_9_2/a_484_472# 0.020188f
C4312 FILLER_0_13_2/a_1828_472# _17_/I 0.00656f
C4313 FILLER_0_10_12/a_572_375# vdd 0.050148f
C4314 FILLER_0_16_18/a_36_472# input9/a_36_113# 0.001663f
C4315 _15_/I FILLER_0_10_37/a_4964_472# 0.015502f
C4316 _17_/I _16_/Z 0.16387f
C4317 _07_/ZN _08_/ZN 0.540896f
C4318 vdd FILLER_0_13_72/a_2812_375# 0.019859f
C4319 FILLER_0_9_2/a_1020_375# _14_/I 0.005451f
C4320 output14/a_224_472# FILLER_0_4_107/a_1468_375# 0.002622f
C4321 FILLER_0_5_104/a_484_472# FILLER_0_7_104/a_572_375# 0.001512f
C4322 FILLER_0_12_101/a_36_472# vdd 0.097837f
C4323 FILLER_0_4_2/a_2364_375# vdd 0.024437f
C4324 FILLER_0_6_107/a_36_472# FILLER_0_4_107/a_124_375# 0.001512f
C4325 output22/a_224_472# output23/a_224_472# 0.031309f
C4326 _18_/I FILLER_0_15_8/a_1828_472# 0.014868f
C4327 FILLER_0_15_40/a_36_472# _19_/I 0.001782f
C4328 vdd FILLER_0_16_18/a_36_472# 0.050638f
C4329 _16_/I FILLER_0_13_2/a_5860_472# 0.004108f
C4330 output18/a_224_472# output_signal_minus[8] 0.115179f
C4331 FILLER_0_9_2/a_4964_472# _15_/I 0.006506f
C4332 FILLER_0_10_107/a_36_472# vdd 0.110617f
C4333 FILLER_0_10_37/a_1380_472# FILLER_0_9_2/a_5412_472# 0.026657f
C4334 FILLER_0_9_2/a_932_472# input_signal[4] 0.001342f
C4335 FILLER_0_6_2/a_2364_375# _12_/I 0.016091f
C4336 _18_/I FILLER_0_14_107/a_572_375# 0.006259f
C4337 FILLER_0_10_37/a_1828_472# FILLER_0_9_2/a_5860_472# 0.026657f
C4338 _16_/I FILLER_0_13_2/a_2364_375# 0.006236f
C4339 FILLER_0_4_37/a_5860_472# FILLER_0_5_72/a_1916_375# 0.001723f
C4340 FILLER_0_6_37/a_5500_375# FILLER_0_7_72/a_1468_375# 0.026339f
C4341 _13_/I FILLER_0_4_101/a_124_375# 0.005726f
C4342 _13_/I output_signal_minus[2] 0.026885f
C4343 _09_/ZN FILLER_0_3_104/a_484_472# 0.006246f
C4344 output11/a_224_472# FILLER_0_2_101/a_124_375# 0.001597f
C4345 FILLER_0_14_115/a_36_472# output28/a_224_472# 0.031509f
C4346 FILLER_0_2_2/a_572_375# vdd 0.019216f
C4347 output_signal_plus[5] _08_/ZN 0.150908f
C4348 FILLER_0_9_2/a_4516_472# vdd 0.005419f
C4349 _16_/I FILLER_0_13_72/a_932_472# 0.004669f
C4350 input_signal[6] FILLER_0_13_2/a_36_472# 0.003542f
C4351 vdd FILLER_0_12_37/a_4516_472# 0.002735f
C4352 FILLER_0_6_2/a_1380_472# _14_/I 0.001219f
C4353 FILLER_0_15_40/a_36_472# _18_/I 0.014431f
C4354 FILLER_0_14_28/a_124_375# vdd 0.014104f
C4355 FILLER_0_11_2/a_4068_472# FILLER_0_13_2/a_4156_375# 0.001512f
C4356 _13_/I FILLER_0_6_37/a_2276_472# 0.003818f
C4357 FILLER_0_3_72/a_1828_472# FILLER_0_5_72/a_1916_375# 0.001512f
C4358 FILLER_0_6_2/a_3260_375# FILLER_0_5_12/a_2276_472# 0.001543f
C4359 _16_/I FILLER_0_10_37/a_4604_375# 0.002119f
C4360 input_signal[6] input7/a_36_113# 0.030631f
C4361 vdd FILLER_0_9_72/a_1020_375# 0.00558f
C4362 FILLER_0_3_72/a_2812_375# FILLER_0_2_37/a_6756_472# 0.001723f
C4363 FILLER_0_4_37/a_4964_472# FILLER_0_2_37/a_5052_375# 0.001512f
C4364 _11_/I FILLER_0_5_104/a_572_375# 0.004712f
C4365 _06_/ZN output14/a_224_472# 0.050195f
C4366 _12_/I FILLER_0_6_37/a_3260_375# 0.016091f
C4367 FILLER_0_2_2/a_3172_472# FILLER_0_2_37/a_36_472# 0.002765f
C4368 _17_/I FILLER_0_13_2/a_1916_375# 0.006125f
C4369 output_signal_plus[8] _18_/a_36_113# 0.008442f
C4370 _09_/ZN _16_/I 0.049108f
C4371 _16_/I FILLER_0_12_37/a_3708_375# 0.016091f
C4372 _14_/I FILLER_0_6_2/a_2724_472# 0.001219f
C4373 _19_/I _19_/Z 2.434557f
C4374 vdd FILLER_0_3_12/a_2812_375# 0.002455f
C4375 vdd FILLER_0_15_72/a_932_472# 0.001979f
C4376 FILLER_0_2_2/a_1020_375# _10_/I 0.001886f
C4377 vdd FILLER_0_10_28/a_124_375# 0.046217f
C4378 _16_/I FILLER_0_10_37/a_1020_375# 0.002327f
C4379 output_signal_minus[5] _01_/ZN 0.001785f
C4380 FILLER_0_12_12/a_1020_375# _16_/I 0.016091f
C4381 vdd FILLER_0_4_2/a_932_472# 0.009004f
C4382 FILLER_0_4_37/a_5948_375# FILLER_0_6_37/a_5860_472# 0.001512f
C4383 FILLER_0_6_37/a_2812_375# _14_/I 0.003099f
C4384 _15_/I FILLER_0_10_37/a_3708_375# 0.018729f
C4385 FILLER_0_6_2/a_2364_375# FILLER_0_5_12/a_1380_472# 0.001543f
C4386 FILLER_0_7_104/a_36_472# FILLER_0_7_72/a_3260_375# 0.086742f
C4387 FILLER_0_14_37/a_4964_472# _16_/I 0.001667f
C4388 _13_/I FILLER_0_4_37/a_1468_375# 0.005726f
C4389 output_signal_minus[3] output14/a_224_472# 0.018548f
C4390 _11_/I FILLER_0_4_37/a_3260_375# 0.01418f
C4391 vdd FILLER_0_16_18/a_932_472# 0.010558f
C4392 FILLER_0_4_37/a_2724_472# FILLER_0_5_60/a_124_375# 0.001723f
C4393 FILLER_0_7_2/a_5948_375# FILLER_0_6_37/a_1916_375# 0.026339f
C4394 FILLER_0_6_107/a_124_375# _14_/I 0.003099f
C4395 _07_/ZN vdd 1.363583f
C4396 FILLER_0_0_12/a_1380_472# FILLER_0_0_28/a_36_472# 0.013276f
C4397 FILLER_0_0_36/a_1468_375# FILLER_0_1_44/a_572_375# 0.05841f
C4398 _18_/I _19_/Z 0.07203f
C4399 FILLER_0_14_37/a_4156_375# _18_/I 0.003988f
C4400 FILLER_0_15_2/a_124_375# input_signal[7] 0.036284f
C4401 FILLER_0_7_72/a_572_375# FILLER_0_6_37/a_4604_375# 0.026339f
C4402 FILLER_0_8_37/a_6308_472# FILLER_0_7_72/a_2364_375# 0.001597f
C4403 FILLER_0_12_12/a_36_472# _15_/I 0.001368f
C4404 FILLER_0_2_107/a_124_375# FILLER_0_4_107/a_36_472# 0.001512f
C4405 FILLER_0_7_2/a_572_375# vdd -0.01037f
C4406 output_signal_minus[1] _08_/ZN 0.303139f
C4407 _18_/I FILLER_0_14_37/a_124_375# 0.003988f
C4408 _13_/I FILLER_0_4_2/a_1468_375# 0.00577f
C4409 vdd FILLER_0_3_44/a_36_472# 0.089951f
C4410 vdd _11_/a_36_113# 0.063638f
C4411 output17/a_224_472# FILLER_0_2_107/a_932_472# 0.031509f
C4412 FILLER_0_4_2/a_2724_472# FILLER_0_5_12/a_1468_375# 0.001684f
C4413 _14_/I FILLER_0_8_37/a_5412_472# 0.014431f
C4414 output27/a_224_472# vdd 0.078796f
C4415 FILLER_0_11_2/a_4964_472# FILLER_0_12_37/a_932_472# 0.026657f
C4416 FILLER_0_1_60/a_124_375# FILLER_0_2_37/a_2724_472# 0.001597f
C4417 _18_/I FILLER_0_14_37/a_3260_375# 0.003988f
C4418 vdd FILLER_0_15_8/a_2276_472# 0.008643f
C4419 FILLER_0_15_64/a_124_375# FILLER_0_14_37/a_3260_375# 0.026339f
C4420 FILLER_0_2_2/a_2724_472# FILLER_0_3_12/a_1468_375# 0.001684f
C4421 FILLER_0_0_70/a_36_472# output20/a_224_472# 0.003196f
C4422 FILLER_0_5_12/a_1020_375# _12_/I 0.002038f
C4423 FILLER_0_11_2/a_2276_472# vdd 0.012553f
C4424 FILLER_0_1_12/a_2276_472# _10_/I 0.006408f
C4425 FILLER_0_2_37/a_6844_375# FILLER_0_2_101/a_124_375# 0.012001f
C4426 FILLER_0_9_2/a_1916_375# vdd 0.051114f
C4427 FILLER_0_0_12/a_36_472# input1/a_36_113# 0.001663f
C4428 _13_/I FILLER_0_4_37/a_6396_375# 0.002482f
C4429 FILLER_0_10_107/a_36_472# _09_/ZN 0.001273f
C4430 FILLER_0_10_37/a_1828_472# FILLER_0_8_37/a_1916_375# 0.001512f
C4431 output_signal_plus[5] vdd 0.127396f
C4432 _17_/I FILLER_0_15_8/a_1020_375# 0.002766f
C4433 vdd FILLER_0_8_37/a_932_472# 0.005627f
C4434 output22/a_224_472# _15_/I 0.047946f
C4435 FILLER_0_8_37/a_4068_472# vdd 0.00286f
C4436 FILLER_0_4_37/a_6308_472# _13_/I 0.002855f
C4437 vdd FILLER_0_3_12/a_484_472# 0.024462f
C4438 _14_/I output16/a_224_472# 0.039773f
C4439 FILLER_0_12_37/a_4516_472# FILLER_0_10_37/a_4604_375# 0.001512f
C4440 _07_/ZN output13/a_224_472# 0.05796f
C4441 FILLER_0_12_37/a_572_375# FILLER_0_14_37/a_484_472# 0.001512f
C4442 vdd FILLER_0_14_37/a_2364_375# 0.026924f
C4443 FILLER_0_11_2/a_6756_472# FILLER_0_12_37/a_2812_375# 0.001597f
C4444 FILLER_0_4_37/a_4068_472# vdd 0.00286f
C4445 vdd FILLER_0_8_12/a_572_375# 0.052255f
C4446 FILLER_0_5_72/a_484_472# vdd 0.002467f
C4447 FILLER_0_14_12/a_572_375# vdd 0.01694f
C4448 vdd FILLER_0_14_37/a_1380_472# 0.007845f
C4449 output25/a_224_472# output_signal_plus[4] 0.059516f
C4450 FILLER_0_10_107/a_1380_472# vdd 0.005026f
C4451 FILLER_0_8_107/a_36_472# FILLER_0_8_101/a_124_375# 0.016748f
C4452 FILLER_0_3_44/a_1380_472# FILLER_0_4_37/a_2276_472# 0.026657f
C4453 FILLER_0_1_12/a_1380_472# FILLER_0_3_12/a_1468_375# 0.0027f
C4454 _07_/ZN output17/a_224_472# 0.097325f
C4455 FILLER_0_14_107/a_124_375# FILLER_0_14_101/a_124_375# 0.005439f
C4456 FILLER_0_7_72/a_484_472# _12_/I 0.004669f
C4457 _16_/I FILLER_0_11_2/a_5052_375# 0.007169f
C4458 _15_/I FILLER_0_9_2/a_1468_375# 0.006125f
C4459 output12/a_224_472# output_signal_minus[2] 0.044725f
C4460 output13/a_224_472# _11_/a_36_113# 0.002131f
C4461 output21/a_224_472# vdd 0.049021f
C4462 _10_/Z output_signal_plus[1] 0.100575f
C4463 FILLER_0_7_2/a_5412_472# FILLER_0_8_37/a_1380_472# 0.026657f
C4464 FILLER_0_1_60/a_36_472# FILLER_0_1_44/a_1468_375# 0.086742f
C4465 FILLER_0_2_37/a_2812_375# FILLER_0_4_37/a_2724_472# 0.001512f
C4466 vdd FILLER_0_10_37/a_36_472# 0.108844f
C4467 FILLER_0_2_107/a_484_472# vdd 0.004107f
C4468 FILLER_0_7_104/a_572_375# _12_/I 0.006193f
C4469 output18/a_224_472# _10_/I 0.053716f
C4470 FILLER_0_2_107/a_932_472# _09_/ZN 0.001711f
C4471 _13_/I FILLER_0_5_72/a_124_375# 0.016362f
C4472 FILLER_0_13_2/a_6308_472# _17_/I 0.006506f
C4473 FILLER_0_11_72/a_1916_375# FILLER_0_10_37/a_5948_375# 0.026339f
C4474 FILLER_0_8_37/a_6844_375# FILLER_0_8_101/a_124_375# 0.012001f
C4475 _12_/I FILLER_0_7_72/a_2364_375# 0.005093f
C4476 FILLER_0_2_101/a_36_472# FILLER_0_2_107/a_36_472# 0.003468f
C4477 _18_/a_36_113# _19_/Z 0.201005f
C4478 FILLER_0_11_72/a_2364_375# FILLER_0_9_72/a_2276_472# 0.001512f
C4479 output_signal_minus[9] output20/a_224_472# 0.03334f
C4480 FILLER_0_4_2/a_2724_472# vdd 0.009191f
C4481 FILLER_0_6_37/a_4964_472# FILLER_0_5_72/a_1020_375# 0.001597f
C4482 FILLER_0_12_12/a_1468_375# FILLER_0_12_28/a_124_375# 0.012001f
C4483 output_signal_minus[7] _10_/Z 0.079577f
C4484 FILLER_0_12_37/a_36_472# vdd 0.108844f
C4485 FILLER_0_6_37/a_2276_472# FILLER_0_4_37/a_2364_375# 0.001512f
C4486 FILLER_0_12_37/a_4068_472# FILLER_0_10_37/a_4156_375# 0.001512f
C4487 FILLER_0_11_2/a_2276_472# FILLER_0_13_2/a_2364_375# 0.0027f
C4488 input_signal[2] FILLER_0_2_2/a_932_472# 0.008791f
C4489 FILLER_0_15_8/a_3172_472# FILLER_0_15_40/a_36_472# 0.013277f
C4490 FILLER_0_2_2/a_572_375# input_signal[1] 0.004159f
C4491 FILLER_0_5_72/a_932_472# vdd 0.004382f
C4492 FILLER_0_7_2/a_3620_472# vdd 0.005895f
C4493 output_signal_minus[1] vdd 0.25191f
C4494 FILLER_0_2_101/a_124_375# _10_/I 0.001886f
C4495 _00_/ZN output25/a_224_472# 0.014879f
C4496 _13_/I FILLER_0_4_37/a_2724_472# 0.003497f
C4497 input_signal[2] FILLER_0_3_12/a_1020_375# 0.001668f
C4498 _15_/I FILLER_0_9_104/a_572_375# 0.006125f
C4499 FILLER_0_6_2/a_932_472# _12_/I 0.022465f
C4500 _17_/I FILLER_0_13_2/a_4068_472# 0.0029f
C4501 FILLER_0_11_72/a_124_375# vdd 0.011994f
C4502 vdd FILLER_0_9_2/a_6844_375# 0.011466f
C4503 FILLER_0_0_12/a_484_472# _10_/I 0.016407f
C4504 _16_/I FILLER_0_14_37/a_484_472# 0.001667f
C4505 _10_/a_36_160# _01_/ZN 0.004846f
C4506 FILLER_0_13_72/a_2276_472# _17_/I 0.00652f
C4507 _17_/I FILLER_0_15_8/a_2724_472# 0.004125f
C4508 FILLER_0_4_37/a_932_472# FILLER_0_3_44/a_36_472# 0.026657f
C4509 _15_/I FILLER_0_9_2/a_2276_472# 0.00656f
C4510 FILLER_0_14_37/a_2812_375# _18_/I 0.003988f
C4511 _09_/ZN _11_/a_36_113# 0.057411f
C4512 FILLER_0_6_37/a_5500_375# _12_/I 0.016091f
C4513 _11_/I net15 0.172728f
C4514 FILLER_0_0_36/a_2276_472# _10_/I 0.016187f
C4515 FILLER_0_4_37/a_3708_375# FILLER_0_6_37/a_3620_472# 0.0027f
C4516 _09_/ZN output27/a_224_472# 0.002783f
C4517 output25/a_224_472# _14_/Z 0.049204f
C4518 output11/a_224_472# FILLER_0_2_37/a_5948_375# 0.001597f
C4519 _11_/Z _03_/ZN 0.012887f
C4520 FILLER_0_11_2/a_2364_375# vdd 0.024816f
C4521 FILLER_0_15_8/a_36_472# input_signal[8] 0.197185f
C4522 _16_/I FILLER_0_11_72/a_5052_375# 0.007169f
C4523 vdd output_signal_plus[6] 0.512148f
C4524 FILLER_0_2_2/a_3172_472# FILLER_0_3_12/a_1916_375# 0.001684f
C4525 _08_/ZN _04_/ZN 0.00174f
C4526 FILLER_0_6_37/a_2364_375# _14_/I 0.001623f
C4527 vdd FILLER_0_14_37/a_6396_375# 0.034034f
C4528 FILLER_0_6_37/a_4156_375# _12_/I 0.016091f
C4529 FILLER_0_14_37/a_4604_375# vdd 0.004123f
C4530 output25/a_224_472# _17_/I 0.005345f
C4531 vdd FILLER_0_15_40/a_124_375# 0.009039f
C4532 vdd FILLER_0_9_72/a_2364_375# 0.022764f
C4533 FILLER_0_2_37/a_2812_375# _10_/I 0.001886f
C4534 FILLER_0_3_72/a_1916_375# vdd 0.009949f
C4535 FILLER_0_15_40/a_484_472# vdd 0.00284f
C4536 FILLER_0_13_2/a_6844_375# vdd 0.011466f
C4537 vdd FILLER_0_6_2/a_124_375# -0.003794f
C4538 output_signal_plus[5] _09_/ZN 0.004194f
C4539 _16_/I FILLER_0_11_2/a_484_472# 0.001841f
C4540 _13_/I FILLER_0_5_44/a_1020_375# 0.016091f
C4541 output_signal_minus[1] output13/a_224_472# 0.009261f
C4542 _17_/I output28/a_224_472# 0.038566f
C4543 _15_/I FILLER_0_10_101/a_36_472# 0.015502f
C4544 FILLER_0_7_72/a_3260_375# FILLER_0_6_101/a_124_375# 0.026339f
C4545 _17_/I FILLER_0_14_12/a_1380_472# 0.015502f
C4546 _16_/I FILLER_0_14_37/a_3620_472# 0.001667f
C4547 vdd FILLER_0_8_12/a_1380_472# 0.011207f
C4548 FILLER_0_4_37/a_2724_472# FILLER_0_3_60/a_36_472# 0.026657f
C4549 FILLER_0_11_2/a_2276_472# FILLER_0_12_12/a_1020_375# 0.001543f
C4550 output30/a_224_472# FILLER_0_15_72/a_932_472# 0.038484f
C4551 FILLER_0_13_104/a_36_472# _17_/I 0.006613f
C4552 FILLER_0_10_107/a_1380_472# _09_/ZN 0.020589f
C4553 output23/a_224_472# _13_/Z 0.030239f
C4554 _10_/I FILLER_0_0_28/a_36_472# 0.016494f
C4555 FILLER_0_6_37/a_5052_375# _12_/I 0.016091f
C4556 FILLER_0_2_2/a_2364_375# _10_/I 0.001886f
C4557 FILLER_0_16_36/a_36_472# vdd 0.104943f
C4558 output_signal_plus[4] _15_/Z 0.04198f
C4559 FILLER_0_11_2/a_1916_375# vdd 0.051101f
C4560 FILLER_0_2_2/a_1468_375# vdd 0.027835f
C4561 FILLER_0_13_72/a_3260_375# vdd 0.010174f
C4562 FILLER_0_1_72/a_36_472# FILLER_0_2_37/a_4068_472# 0.026657f
C4563 FILLER_0_3_60/a_484_472# FILLER_0_3_72/a_36_472# 0.002296f
C4564 FILLER_0_12_37/a_1468_375# FILLER_0_13_2/a_5500_375# 0.026339f
C4565 FILLER_0_12_37/a_5412_472# FILLER_0_11_72/a_1380_472# 0.026657f
C4566 _11_/I FILLER_0_4_37/a_5052_375# 0.01418f
C4567 input_signal[3] FILLER_0_4_2/a_932_472# 0.003222f
C4568 FILLER_0_3_72/a_3172_472# FILLER_0_5_72/a_3260_375# 0.001512f
C4569 FILLER_0_7_2/a_3172_472# _12_/I 0.004669f
C4570 FILLER_0_14_37/a_3172_472# _18_/I 0.001526f
C4571 FILLER_0_14_12/a_1020_375# _17_/I 0.018729f
C4572 _13_/I FILLER_0_4_37/a_5948_375# 0.005726f
C4573 output25/a_224_472# output_signal_plus[3] 0.002485f
C4574 FILLER_0_2_37/a_5412_472# _10_/I 0.002486f
C4575 FILLER_0_15_64/a_124_375# FILLER_0_14_37/a_3172_472# 0.001723f
C4576 vdd FILLER_0_11_2/a_1020_375# 0.022339f
C4577 FILLER_0_2_2/a_484_472# vdd 0.008472f
C4578 FILLER_0_14_37/a_5500_375# FILLER_0_15_72/a_1468_375# 0.026339f
C4579 FILLER_0_13_72/a_3172_472# _16_/I 0.004669f
C4580 _13_/I _10_/I 0.007137f
C4581 _13_/I FILLER_0_5_12/a_2364_375# 0.016091f
C4582 FILLER_0_8_37/a_4964_472# FILLER_0_7_72/a_932_472# 0.026657f
C4583 FILLER_0_7_72/a_36_472# _14_/I 0.008683f
C4584 FILLER_0_7_2/a_4516_472# FILLER_0_8_37/a_572_375# 0.001597f
C4585 output23/a_224_472# _14_/I 0.031637f
C4586 _16_/I input_signal[7] 0.024419f
C4587 FILLER_0_12_37/a_124_375# FILLER_0_11_2/a_4068_472# 0.001597f
C4588 FILLER_0_11_2/a_1468_375# FILLER_0_9_2/a_1380_472# 0.0027f
C4589 _13_/I FILLER_0_6_37/a_124_375# 0.001706f
C4590 output11/a_224_472# output_signal_minus[0] 0.024072f
C4591 _14_/I FILLER_0_9_104/a_124_375# 0.005433f
C4592 FILLER_0_3_12/a_1020_375# FILLER_0_1_12/a_932_472# 0.0027f
C4593 _17_/I FILLER_0_13_104/a_484_472# 0.006506f
C4594 output24/a_224_472# _15_/a_36_113# 0.012996f
C4595 FILLER_0_4_37/a_3620_472# FILLER_0_2_37/a_3708_375# 0.0027f
C4596 FILLER_0_9_104/a_36_472# FILLER_0_9_72/a_3260_375# 0.086742f
C4597 FILLER_0_8_12/a_124_375# vdd 0.033331f
C4598 FILLER_0_14_101/a_36_472# FILLER_0_14_37/a_6844_375# 0.086635f
C4599 _01_/ZN FILLER_0_2_107/a_124_375# 0.001597f
C4600 output_signal_plus[2] _10_/Z 0.070884f
C4601 vdd FILLER_0_5_60/a_484_472# 0.012891f
C4602 FILLER_0_2_2/a_1828_472# FILLER_0_1_12/a_572_375# 0.001543f
C4603 _11_/I output_signal_minus[4] 0.664575f
C4604 FILLER_0_8_37/a_572_375# FILLER_0_10_37/a_484_472# 0.001512f
C4605 FILLER_0_2_37/a_1468_375# FILLER_0_3_44/a_572_375# 0.026339f
C4606 FILLER_0_4_2/a_484_472# _12_/I 0.049518f
C4607 FILLER_0_5_72/a_2812_375# _12_/I 0.001706f
C4608 FILLER_0_1_12/a_3172_472# vdd 0.002817f
C4609 FILLER_0_4_37/a_6756_472# vdd 0.015684f
C4610 FILLER_0_7_104/a_124_375# _03_/ZN 0.002258f
C4611 _00_/ZN _15_/Z 0.184979f
C4612 _07_/ZN output_signal_minus[2] 0.123667f
C4613 FILLER_0_14_37/a_5052_375# FILLER_0_15_72/a_1020_375# 0.026339f
C4614 FILLER_0_6_37/a_2724_472# _12_/I 0.017477f
C4615 FILLER_0_7_2/a_1828_472# _14_/I 0.008733f
C4616 _15_/I FILLER_0_11_72/a_3620_472# 0.005458f
C4617 vdd FILLER_0_4_37/a_36_472# 0.10831f
C4618 _16_/I FILLER_0_13_2/a_6396_375# 0.006193f
C4619 vdd _04_/ZN 0.082622f
C4620 FILLER_0_7_2/a_3708_375# _12_/I 0.006313f
C4621 _01_/ZN FILLER_0_2_107/a_36_472# 0.031889f
C4622 _12_/I FILLER_0_5_72/a_1828_472# 0.003805f
C4623 vdd FILLER_0_7_2/a_2364_375# -0.007297f
C4624 _15_/I FILLER_0_10_37/a_2812_375# 0.018729f
C4625 FILLER_0_8_107/a_572_375# vdd 0.030961f
C4626 FILLER_0_6_101/a_36_472# _14_/I 0.001219f
C4627 _14_/I FILLER_0_6_37/a_5860_472# 0.001219f
C4628 FILLER_0_15_8/a_1380_472# FILLER_0_16_18/a_124_375# 0.001543f
C4629 _11_/I FILLER_0_3_12/a_124_375# 0.010835f
C4630 FILLER_0_9_66/a_36_472# _14_/I 0.004017f
C4631 _18_/I FILLER_0_14_37/a_3708_375# 0.00404f
C4632 FILLER_0_2_37/a_2364_375# _10_/I 0.001352f
C4633 FILLER_0_8_37/a_4516_472# FILLER_0_7_72/a_484_472# 0.026657f
C4634 _15_/I FILLER_0_10_37/a_6308_472# 0.015502f
C4635 FILLER_0_2_37/a_3708_375# vdd 0.021933f
C4636 FILLER_0_12_107/a_484_472# _15_/I 0.001368f
C4637 FILLER_0_2_37/a_1380_472# vdd 0.009105f
C4638 FILLER_0_4_37/a_1916_375# _11_/I 0.01418f
C4639 FILLER_0_6_2/a_2812_375# vdd -0.009691f
C4640 FILLER_0_16_36/a_2812_375# vdd 0.007113f
C4641 FILLER_0_7_2/a_1380_472# FILLER_0_9_2/a_1468_375# 0.0027f
C4642 vdd FILLER_0_13_2/a_2724_472# 0.011159f
C4643 FILLER_0_6_2/a_3172_472# FILLER_0_6_37/a_36_472# 0.002765f
C4644 _09_/ZN output_signal_plus[6] 0.001179f
C4645 _13_/I FILLER_0_4_107/a_484_472# 0.003777f
C4646 _14_/Z _15_/Z 0.611858f
C4647 FILLER_0_11_136/a_36_472# FILLER_0_11_72/a_6844_375# 0.086635f
C4648 _16_/I FILLER_0_10_37/a_3708_375# 0.002327f
C4649 _15_/I FILLER_0_11_2/a_4964_472# 0.005458f
C4650 FILLER_0_0_36/a_932_472# _10_/I 0.016187f
C4651 FILLER_0_11_72/a_3172_472# vdd 0.009528f
C4652 FILLER_0_6_37/a_3172_472# vdd 0.006735f
C4653 _17_/I _15_/Z 0.317682f
C4654 FILLER_0_10_37/a_3172_472# FILLER_0_8_37/a_3260_375# 0.001512f
C4655 FILLER_0_0_70/a_124_375# FILLER_0_0_36/a_3260_375# 0.005439f
C4656 FILLER_0_8_12/a_1468_375# _15_/I 0.002388f
C4657 FILLER_0_4_37/a_5412_472# vdd 0.006451f
C4658 _17_/I FILLER_0_13_2/a_5500_375# 0.006125f
C4659 vdd FILLER_0_13_2/a_1468_375# 0.027811f
C4660 FILLER_0_10_37/a_4964_472# FILLER_0_9_72/a_1020_375# 0.001597f
C4661 _17_/I FILLER_0_12_107/a_1020_375# 0.001551f
C4662 FILLER_0_12_12/a_36_472# _16_/I 0.027902f
C4663 FILLER_0_1_12/a_3260_375# vdd -0.011968f
C4664 FILLER_0_13_2/a_4156_375# _16_/I 0.006193f
C4665 _14_/I FILLER_0_8_37/a_2364_375# 0.01418f
C4666 _12_/I FILLER_0_7_2/a_2812_375# 0.006134f
C4667 vdd FILLER_0_16_36/a_1380_472# 0.004364f
C4668 FILLER_0_5_44/a_572_375# FILLER_0_3_44/a_484_472# 0.001512f
C4669 FILLER_0_14_37/a_932_472# _17_/I 0.015502f
C4670 _15_/I FILLER_0_11_72/a_5860_472# 0.005458f
C4671 _11_/I FILLER_0_2_37/a_1828_472# 0.002415f
C4672 FILLER_0_14_115/a_124_375# FILLER_0_14_107/a_572_375# 0.012001f
C4673 FILLER_0_6_37/a_6756_472# FILLER_0_6_101/a_36_472# 0.013277f
C4674 FILLER_0_15_40/a_36_472# FILLER_0_16_36/a_484_472# 0.05841f
C4675 _15_/I _13_/Z 0.076848f
C4676 FILLER_0_9_72/a_2812_375# vdd 0.019868f
C4677 FILLER_0_2_37/a_4964_472# vdd 0.006196f
C4678 FILLER_0_15_8/a_1916_375# vdd -0.008756f
C4679 FILLER_0_2_107/a_932_472# output_signal_minus[8] 0.007707f
C4680 _16_/I FILLER_0_13_72/a_484_472# 0.004669f
C4681 FILLER_0_6_2/a_1020_375# FILLER_0_7_2/a_1020_375# 0.05841f
C4682 _15_/I FILLER_0_11_72/a_2812_375# 0.00583f
C4683 vdd FILLER_0_5_104/a_124_375# 0.027728f
C4684 _00_/ZN output_signal_plus[1] 0.041288f
C4685 FILLER_0_2_37/a_5948_375# _10_/I 0.001886f
C4686 _19_/a_36_113# output_signal_plus[7] 0.014264f
C4687 output_signal_plus[3] _15_/Z 0.350581f
C4688 FILLER_0_6_37/a_1380_472# _14_/I 0.001219f
C4689 _12_/a_36_113# net15 0.006186f
C4690 vdd FILLER_0_12_37/a_3620_472# 0.007765f
C4691 FILLER_0_5_72/a_36_472# FILLER_0_5_60/a_484_472# 0.002296f
C4692 _17_/a_36_113# output_signal_plus[6] 0.015529f
C4693 vdd FILLER_0_16_18/a_1380_472# 0.014764f
C4694 _11_/I FILLER_0_5_104/a_484_472# 0.001913f
C4695 FILLER_0_13_2/a_5052_375# _17_/I 0.006125f
C4696 FILLER_0_9_104/a_484_472# FILLER_0_11_72/a_4156_375# 0.001512f
C4697 FILLER_0_4_37/a_5412_472# FILLER_0_2_37/a_5500_375# 0.001512f
C4698 FILLER_0_0_36/a_3172_472# _10_/I 0.01623f
C4699 _15_/I FILLER_0_9_2/a_1020_375# 0.006125f
C4700 _17_/I FILLER_0_14_37/a_1020_375# 0.018729f
C4701 _12_/I FILLER_0_5_60/a_572_375# 0.001706f
C4702 _12_/Z net15 0.009957f
C4703 vdd FILLER_0_15_40/a_572_375# 0.006749f
C4704 _15_/I FILLER_0_10_12/a_124_375# 0.01948f
C4705 _15_/I _14_/I 0.025535f
C4706 _19_/I FILLER_0_16_18/a_36_472# 0.014431f
C4707 FILLER_0_6_37/a_6396_375# vdd 0.038787f
C4708 output_signal_minus[9] output18/a_224_472# 0.008677f
C4709 FILLER_0_4_2/a_1828_472# _12_/I 0.001124f
C4710 _14_/Z output_signal_plus[1] 0.057785f
C4711 _00_/ZN output_signal_minus[7] 0.174901f
C4712 FILLER_0_7_2/a_1020_375# input_signal[4] 0.001353f
C4713 FILLER_0_13_2/a_2812_375# vdd 0.022556f
C4714 FILLER_0_7_66/a_124_375# FILLER_0_7_72/a_124_375# 0.005439f
C4715 _13_/I FILLER_0_6_37/a_5948_375# 0.001706f
C4716 FILLER_0_14_37/a_4604_375# output30/a_224_472# 0.001234f
C4717 FILLER_0_12_12/a_932_472# vdd 0.016607f
C4718 _15_/I FILLER_0_11_72/a_4964_472# 0.005458f
C4719 _07_/ZN output_signal_minus[8] 0.113708f
C4720 output_signal_minus[1] output_signal_minus[2] 0.253585f
C4721 FILLER_0_10_37/a_6396_375# vdd 0.036586f
C4722 input_signal[3] FILLER_0_6_2/a_124_375# 0.004728f
C4723 FILLER_0_13_2/a_3708_375# vdd 0.018728f
C4724 FILLER_0_9_104/a_36_472# FILLER_0_11_72/a_3708_375# 0.0027f
C4725 FILLER_0_5_12/a_3172_472# _12_/I 0.003805f
C4726 FILLER_0_7_2/a_4156_375# vdd 0.004458f
C4727 FILLER_0_12_12/a_124_375# FILLER_0_14_12/a_36_472# 0.0027f
C4728 FILLER_0_10_107/a_932_472# _11_/Z 0.032348f
C4729 vdd FILLER_0_11_72/a_1020_375# 0.00558f
C4730 FILLER_0_5_12/a_2812_375# FILLER_0_4_37/a_36_472# 0.001723f
C4731 FILLER_0_16_70/a_124_375# FILLER_0_16_36/a_3260_375# 0.005439f
C4732 _16_/I FILLER_0_13_72/a_124_375# 0.006182f
C4733 _11_/I FILLER_0_5_72/a_3172_472# 0.001913f
C4734 input_signal[9] input_signal[8] 0.472617f
C4735 FILLER_0_2_2/a_484_472# input_signal[1] 0.004572f
C4736 FILLER_0_4_2/a_1468_375# FILLER_0_3_12/a_484_472# 0.001543f
C4737 _11_/I _02_/ZN 0.032042f
C4738 FILLER_0_7_72/a_1916_375# FILLER_0_5_72/a_1828_472# 0.001512f
C4739 FILLER_0_7_2/a_3620_472# FILLER_0_9_2/a_3708_375# 0.0027f
C4740 FILLER_0_2_2/a_3260_375# FILLER_0_1_12/a_2276_472# 0.001543f
C4741 FILLER_0_5_12/a_1020_375# FILLER_0_3_12/a_932_472# 0.0027f
C4742 _18_/I FILLER_0_16_18/a_36_472# 0.012849f
C4743 _11_/I _10_/Z 0.111253f
C4744 FILLER_0_9_66/a_36_472# FILLER_0_11_66/a_124_375# 0.001512f
C4745 FILLER_0_4_2/a_2276_472# FILLER_0_3_12/a_1020_375# 0.001543f
C4746 FILLER_0_13_2/a_4604_375# _17_/I 0.006125f
C4747 vdd _18_/Z 0.203096f
C4748 output_signal_minus[0] _10_/I 0.062197f
C4749 _11_/I FILLER_0_4_101/a_36_472# 0.014431f
C4750 FILLER_0_3_72/a_124_375# FILLER_0_1_72/a_36_472# 0.001512f
C4751 _13_/I FILLER_0_4_37/a_1828_472# 0.003497f
C4752 FILLER_0_13_104/a_572_375# FILLER_0_11_72/a_4068_472# 0.001512f
C4753 FILLER_0_9_72/a_124_375# FILLER_0_8_37/a_4156_375# 0.026339f
C4754 _19_/I FILLER_0_15_72/a_932_472# 0.001678f
C4755 output_signal_plus[3] output_signal_plus[1] 0.005056f
C4756 FILLER_0_15_8/a_1380_472# _17_/I 0.003525f
C4757 _15_/I FILLER_0_12_28/a_36_472# 0.001368f
C4758 _16_/I _16_/a_36_113# 0.049132f
C4759 FILLER_0_16_70/a_124_375# vdd 0.025757f
C4760 FILLER_0_12_101/a_124_375# vdd 0.043908f
C4761 _15_/a_36_113# _08_/ZN 0.001057f
C4762 FILLER_0_8_37/a_484_472# FILLER_0_7_2/a_4516_472# 0.026657f
C4763 _15_/I FILLER_0_11_2/a_5948_375# 0.004401f
C4764 FILLER_0_14_28/a_124_375# _18_/I 0.003935f
C4765 _16_/I FILLER_0_13_2/a_5948_375# 0.003867f
C4766 vdd FILLER_0_7_72/a_3260_375# 0.010174f
C4767 _12_/a_36_113# output_signal_minus[4] 0.007124f
C4768 FILLER_0_6_37/a_6308_472# _12_/I 0.017477f
C4769 vdd FILLER_0_15_72/a_1020_375# 0.005404f
C4770 output_signal_minus[6] net15 0.002062f
C4771 _19_/I FILLER_0_16_18/a_932_472# 0.014431f
C4772 FILLER_0_15_8/a_3260_375# vdd 0.003875f
C4773 FILLER_0_4_2/a_1380_472# FILLER_0_5_12/a_124_375# 0.001684f
C4774 _13_/I _13_/Z 0.01597f
C4775 _11_/I input3/a_36_113# 0.016795f
C4776 FILLER_0_4_37/a_5500_375# FILLER_0_5_72/a_1468_375# 0.026339f
C4777 vdd FILLER_0_5_12/a_572_375# 0.052283f
C4778 FILLER_0_14_37/a_484_472# FILLER_0_15_40/a_124_375# 0.001723f
C4779 FILLER_0_2_107/a_484_472# output_signal_minus[8] 0.003305f
C4780 FILLER_0_4_2/a_1380_472# vdd 0.011604f
C4781 FILLER_0_8_37/a_6308_472# FILLER_0_7_72/a_2276_472# 0.026657f
C4782 FILLER_0_15_56/a_124_375# FILLER_0_14_37/a_2364_375# 0.026339f
C4783 FILLER_0_15_40/a_1380_472# FILLER_0_16_36/a_1828_472# 0.05841f
C4784 _12_/Z output_signal_minus[4] 0.004744f
C4785 _09_/ZN FILLER_0_5_104/a_124_375# 0.001685f
C4786 _18_/I FILLER_0_15_72/a_932_472# 0.014431f
C4787 FILLER_0_0_28/a_124_375# FILLER_0_0_12/a_1468_375# 0.012001f
C4788 FILLER_0_12_37/a_6396_375# _17_/I 0.001106f
C4789 FILLER_0_14_28/a_124_375# FILLER_0_14_12/a_1468_375# 0.012001f
C4790 output_signal_plus[9] vss 0.405805f
C4791 _19_/Z vss 1.30414f
C4792 output30/a_224_472# vss 2.434601f
C4793 FILLER_0_1_60/a_484_472# vss 0.351448f
C4794 FILLER_0_1_60/a_36_472# vss 0.407263f
C4795 FILLER_0_1_60/a_572_375# vss 0.254574f
C4796 FILLER_0_1_60/a_124_375# vss 0.187795f
C4797 FILLER_0_0_28/a_36_472# vss 0.424906f
C4798 FILLER_0_0_28/a_124_375# vss 0.268784f
C4799 FILLER_0_13_72/a_3172_472# vss 0.351491f
C4800 FILLER_0_13_72/a_2724_472# vss 0.332816f
C4801 FILLER_0_13_72/a_2276_472# vss 0.333278f
C4802 FILLER_0_13_72/a_1828_472# vss 0.336102f
C4803 FILLER_0_13_72/a_1380_472# vss 0.337801f
C4804 FILLER_0_13_72/a_932_472# vss 0.340498f
C4805 FILLER_0_13_72/a_484_472# vss 0.371346f
C4806 FILLER_0_13_72/a_36_472# vss 0.415873f
C4807 FILLER_0_13_72/a_3260_375# vss 0.290708f
C4808 FILLER_0_13_72/a_2812_375# vss 0.171987f
C4809 FILLER_0_13_72/a_2364_375# vss 0.171987f
C4810 FILLER_0_13_72/a_1916_375# vss 0.175274f
C4811 FILLER_0_13_72/a_1468_375# vss 0.176943f
C4812 FILLER_0_13_72/a_1020_375# vss 0.179193f
C4813 FILLER_0_13_72/a_572_375# vss 0.198742f
C4814 FILLER_0_13_72/a_124_375# vss 0.200509f
C4815 FILLER_0_2_107/a_1380_472# vss 0.352409f
C4816 FILLER_0_2_107/a_932_472# vss 0.363161f
C4817 FILLER_0_2_107/a_484_472# vss 0.341341f
C4818 FILLER_0_2_107/a_36_472# vss 0.413257f
C4819 FILLER_0_2_107/a_1468_375# vss 0.24369f
C4820 FILLER_0_2_107/a_1020_375# vss 0.191476f
C4821 FILLER_0_2_107/a_572_375# vss 0.191665f
C4822 FILLER_0_2_107/a_124_375# vss 0.195323f
C4823 FILLER_0_5_104/a_484_472# vss 0.352309f
C4824 FILLER_0_5_104/a_36_472# vss 0.410889f
C4825 FILLER_0_5_104/a_572_375# vss 0.249887f
C4826 FILLER_0_5_104/a_124_375# vss 0.190626f
C4827 FILLER_0_6_37/a_6756_472# vss 0.347527f
C4828 FILLER_0_6_37/a_6308_472# vss 0.331577f
C4829 FILLER_0_6_37/a_5860_472# vss 0.33401f
C4830 FILLER_0_6_37/a_5412_472# vss 0.335276f
C4831 FILLER_0_6_37/a_4964_472# vss 0.337162f
C4832 FILLER_0_6_37/a_4516_472# vss 0.353881f
C4833 FILLER_0_6_37/a_4068_472# vss 0.341294f
C4834 FILLER_0_6_37/a_3620_472# vss 0.339239f
C4835 FILLER_0_6_37/a_3172_472# vss 0.334823f
C4836 FILLER_0_6_37/a_2724_472# vss 0.333748f
C4837 FILLER_0_6_37/a_2276_472# vss 0.331577f
C4838 FILLER_0_6_37/a_1828_472# vss 0.332467f
C4839 FILLER_0_6_37/a_1380_472# vss 0.334418f
C4840 FILLER_0_6_37/a_932_472# vss 0.335895f
C4841 FILLER_0_6_37/a_484_472# vss 0.338195f
C4842 FILLER_0_6_37/a_36_472# vss 0.446096f
C4843 FILLER_0_6_37/a_6844_375# vss 0.288762f
C4844 FILLER_0_6_37/a_6396_375# vss 0.171802f
C4845 FILLER_0_6_37/a_5948_375# vss 0.174707f
C4846 FILLER_0_6_37/a_5500_375# vss 0.17616f
C4847 FILLER_0_6_37/a_5052_375# vss 0.178237f
C4848 FILLER_0_6_37/a_4604_375# vss 0.183967f
C4849 FILLER_0_6_37/a_4156_375# vss 0.198537f
C4850 FILLER_0_6_37/a_3708_375# vss 0.179261f
C4851 FILLER_0_6_37/a_3260_375# vss 0.176687f
C4852 FILLER_0_6_37/a_2812_375# vss 0.175071f
C4853 FILLER_0_6_37/a_2364_375# vss 0.171961f
C4854 FILLER_0_6_37/a_1916_375# vss 0.172079f
C4855 FILLER_0_6_37/a_1468_375# vss 0.175335f
C4856 FILLER_0_6_37/a_1020_375# vss 0.177038f
C4857 FILLER_0_6_37/a_572_375# vss 0.179211f
C4858 FILLER_0_6_37/a_124_375# vss 0.222087f
C4859 input_signal[4] vss 1.247059f
C4860 FILLER_0_8_101/a_36_472# vss 0.423424f
C4861 FILLER_0_8_101/a_124_375# vss 0.298762f
C4862 FILLER_0_16_104/a_36_472# vss 0.425296f
C4863 FILLER_0_16_104/a_124_375# vss 0.259163f
C4864 FILLER_0_12_28/a_36_472# vss 0.425395f
C4865 FILLER_0_12_28/a_124_375# vss 0.265471f
C4866 FILLER_0_11_2/a_6756_472# vss 0.350352f
C4867 FILLER_0_11_2/a_6308_472# vss 0.331577f
C4868 FILLER_0_11_2/a_5860_472# vss 0.331577f
C4869 FILLER_0_11_2/a_5412_472# vss 0.334643f
C4870 FILLER_0_11_2/a_4964_472# vss 0.336301f
C4871 FILLER_0_11_2/a_4516_472# vss 0.338848f
C4872 FILLER_0_11_2/a_4068_472# vss 0.363177f
C4873 FILLER_0_11_2/a_3620_472# vss 0.342921f
C4874 FILLER_0_11_2/a_3172_472# vss 0.338101f
C4875 FILLER_0_11_2/a_2724_472# vss 0.33745f
C4876 FILLER_0_11_2/a_2276_472# vss 0.335621f
C4877 FILLER_0_11_2/a_1828_472# vss 0.333666f
C4878 FILLER_0_11_2/a_1380_472# vss 0.333666f
C4879 FILLER_0_11_2/a_932_472# vss 0.333666f
C4880 FILLER_0_11_2/a_484_472# vss 0.33241f
C4881 FILLER_0_11_2/a_36_472# vss 0.408581f
C4882 FILLER_0_11_2/a_6844_375# vss 0.291562f
C4883 FILLER_0_11_2/a_6396_375# vss 0.172168f
C4884 FILLER_0_11_2/a_5948_375# vss 0.171802f
C4885 FILLER_0_11_2/a_5500_375# vss 0.174928f
C4886 FILLER_0_11_2/a_5052_375# vss 0.17651f
C4887 FILLER_0_11_2/a_4604_375# vss 0.178722f
C4888 FILLER_0_11_2/a_4156_375# vss 0.191165f
C4889 FILLER_0_11_2/a_3708_375# vss 0.191898f
C4890 FILLER_0_11_2/a_3260_375# vss 0.178853f
C4891 FILLER_0_11_2/a_2812_375# vss 0.176722f
C4892 FILLER_0_11_2/a_2364_375# vss 0.175137f
C4893 FILLER_0_11_2/a_1916_375# vss 0.17209f
C4894 FILLER_0_11_2/a_1468_375# vss 0.17209f
C4895 FILLER_0_11_2/a_1020_375# vss 0.17209f
C4896 FILLER_0_11_2/a_572_375# vss 0.171927f
C4897 FILLER_0_11_2/a_124_375# vss 0.188994f
C4898 FILLER_0_16_70/a_36_472# vss 0.429713f
C4899 FILLER_0_16_70/a_124_375# vss 0.265239f
C4900 FILLER_0_15_8/a_3172_472# vss 0.37487f
C4901 FILLER_0_15_8/a_2724_472# vss 0.339039f
C4902 FILLER_0_15_8/a_2276_472# vss 0.337695f
C4903 FILLER_0_15_8/a_1828_472# vss 0.336291f
C4904 FILLER_0_15_8/a_1380_472# vss 0.333736f
C4905 FILLER_0_15_8/a_932_472# vss 0.333666f
C4906 FILLER_0_15_8/a_484_472# vss 0.33241f
C4907 FILLER_0_15_8/a_36_472# vss 0.40747f
C4908 FILLER_0_15_8/a_3260_375# vss 0.331787f
C4909 FILLER_0_15_8/a_2812_375# vss 0.180266f
C4910 FILLER_0_15_8/a_2364_375# vss 0.177037f
C4911 FILLER_0_15_8/a_1916_375# vss 0.175199f
C4912 FILLER_0_15_8/a_1468_375# vss 0.172355f
C4913 FILLER_0_15_8/a_1020_375# vss 0.17167f
C4914 FILLER_0_15_8/a_572_375# vss 0.17167f
C4915 FILLER_0_15_8/a_124_375# vss 0.186386f
C4916 vdd vss 0.39933p
C4917 FILLER_0_0_36/a_3172_472# vss 0.351976f
C4918 FILLER_0_0_36/a_2724_472# vss 0.333825f
C4919 FILLER_0_0_36/a_2276_472# vss 0.33241f
C4920 FILLER_0_0_36/a_1828_472# vss 0.334216f
C4921 FILLER_0_0_36/a_1380_472# vss 0.33597f
C4922 FILLER_0_0_36/a_932_472# vss 0.337858f
C4923 FILLER_0_0_36/a_484_472# vss 0.340851f
C4924 FILLER_0_0_36/a_36_472# vss 0.437752f
C4925 FILLER_0_0_36/a_3260_375# vss 0.28576f
C4926 FILLER_0_0_36/a_2812_375# vss 0.174073f
C4927 FILLER_0_0_36/a_2364_375# vss 0.17167f
C4928 FILLER_0_0_36/a_1916_375# vss 0.172727f
C4929 FILLER_0_0_36/a_1468_375# vss 0.175034f
C4930 FILLER_0_0_36/a_1020_375# vss 0.176762f
C4931 FILLER_0_0_36/a_572_375# vss 0.179053f
C4932 FILLER_0_0_36/a_124_375# vss 0.232475f
C4933 _10_/a_36_160# vss 0.395723f
C4934 FILLER_0_10_107/a_1380_472# vss 0.353246f
C4935 FILLER_0_10_107/a_932_472# vss 0.361941f
C4936 FILLER_0_10_107/a_484_472# vss 0.340589f
C4937 FILLER_0_10_107/a_36_472# vss 0.413139f
C4938 FILLER_0_10_107/a_1468_375# vss 0.243852f
C4939 FILLER_0_10_107/a_1020_375# vss 0.189352f
C4940 FILLER_0_10_107/a_572_375# vss 0.189181f
C4941 FILLER_0_10_107/a_124_375# vss 0.194299f
C4942 FILLER_0_12_37/a_6756_472# vss 0.347527f
C4943 FILLER_0_12_37/a_6308_472# vss 0.331577f
C4944 FILLER_0_12_37/a_5860_472# vss 0.33401f
C4945 FILLER_0_12_37/a_5412_472# vss 0.335276f
C4946 FILLER_0_12_37/a_4964_472# vss 0.337162f
C4947 FILLER_0_12_37/a_4516_472# vss 0.353881f
C4948 FILLER_0_12_37/a_4068_472# vss 0.341338f
C4949 FILLER_0_12_37/a_3620_472# vss 0.339239f
C4950 FILLER_0_12_37/a_3172_472# vss 0.336106f
C4951 FILLER_0_12_37/a_2724_472# vss 0.334988f
C4952 FILLER_0_12_37/a_2276_472# vss 0.332816f
C4953 FILLER_0_12_37/a_1828_472# vss 0.333707f
C4954 FILLER_0_12_37/a_1380_472# vss 0.335658f
C4955 FILLER_0_12_37/a_932_472# vss 0.337134f
C4956 FILLER_0_12_37/a_484_472# vss 0.339435f
C4957 FILLER_0_12_37/a_36_472# vss 0.447577f
C4958 FILLER_0_12_37/a_6844_375# vss 0.288762f
C4959 FILLER_0_12_37/a_6396_375# vss 0.171802f
C4960 FILLER_0_12_37/a_5948_375# vss 0.174707f
C4961 FILLER_0_12_37/a_5500_375# vss 0.17616f
C4962 FILLER_0_12_37/a_5052_375# vss 0.178237f
C4963 FILLER_0_12_37/a_4604_375# vss 0.183967f
C4964 FILLER_0_12_37/a_4156_375# vss 0.198537f
C4965 FILLER_0_12_37/a_3708_375# vss 0.179261f
C4966 FILLER_0_12_37/a_3260_375# vss 0.176687f
C4967 FILLER_0_12_37/a_2812_375# vss 0.175071f
C4968 FILLER_0_12_37/a_2364_375# vss 0.171961f
C4969 FILLER_0_12_37/a_1916_375# vss 0.172079f
C4970 FILLER_0_12_37/a_1468_375# vss 0.175335f
C4971 FILLER_0_12_37/a_1020_375# vss 0.177038f
C4972 FILLER_0_12_37/a_572_375# vss 0.179212f
C4973 FILLER_0_12_37/a_124_375# vss 0.222087f
C4974 FILLER_0_13_104/a_484_472# vss 0.353546f
C4975 FILLER_0_13_104/a_36_472# vss 0.411703f
C4976 FILLER_0_13_104/a_572_375# vss 0.25017f
C4977 FILLER_0_13_104/a_124_375# vss 0.190801f
C4978 input_signal[6] vss 1.179258f
C4979 _11_/Z vss 1.237957f
C4980 _11_/a_36_113# vss 0.437095f
C4981 FILLER_0_9_66/a_36_472# vss 0.425205f
C4982 FILLER_0_9_66/a_124_375# vss 0.300651f
C4983 FILLER_0_3_12/a_3172_472# vss 0.358005f
C4984 FILLER_0_3_12/a_2724_472# vss 0.365013f
C4985 FILLER_0_3_12/a_2276_472# vss 0.339207f
C4986 FILLER_0_3_12/a_1828_472# vss 0.338282f
C4987 FILLER_0_3_12/a_1380_472# vss 0.336686f
C4988 FILLER_0_3_12/a_932_472# vss 0.333727f
C4989 FILLER_0_3_12/a_484_472# vss 0.333639f
C4990 FILLER_0_3_12/a_36_472# vss 0.407776f
C4991 FILLER_0_3_12/a_3260_375# vss 0.294263f
C4992 FILLER_0_3_12/a_2812_375# vss 0.219231f
C4993 FILLER_0_3_12/a_2364_375# vss 0.180554f
C4994 FILLER_0_3_12/a_1916_375# vss 0.177813f
C4995 FILLER_0_3_12/a_1468_375# vss 0.175853f
C4996 FILLER_0_3_12/a_1020_375# vss 0.172934f
C4997 FILLER_0_3_12/a_572_375# vss 0.172109f
C4998 FILLER_0_3_12/a_124_375# vss 0.186354f
C4999 FILLER_0_2_2/a_3172_472# vss 0.354973f
C5000 FILLER_0_2_2/a_2724_472# vss 0.337495f
C5001 FILLER_0_2_2/a_2276_472# vss 0.335691f
C5002 FILLER_0_2_2/a_1828_472# vss 0.333736f
C5003 FILLER_0_2_2/a_1380_472# vss 0.333736f
C5004 FILLER_0_2_2/a_932_472# vss 0.333736f
C5005 FILLER_0_2_2/a_484_472# vss 0.332471f
C5006 FILLER_0_2_2/a_36_472# vss 0.408737f
C5007 FILLER_0_2_2/a_3260_375# vss 0.266669f
C5008 FILLER_0_2_2/a_2812_375# vss 0.176735f
C5009 FILLER_0_2_2/a_2364_375# vss 0.175157f
C5010 FILLER_0_2_2/a_1916_375# vss 0.172109f
C5011 FILLER_0_2_2/a_1468_375# vss 0.172109f
C5012 FILLER_0_2_2/a_1020_375# vss 0.172109f
C5013 FILLER_0_2_2/a_572_375# vss 0.171953f
C5014 FILLER_0_2_2/a_124_375# vss 0.189405f
C5015 FILLER_0_13_2/a_6756_472# vss 0.350424f
C5016 FILLER_0_13_2/a_6308_472# vss 0.331648f
C5017 FILLER_0_13_2/a_5860_472# vss 0.331648f
C5018 FILLER_0_13_2/a_5412_472# vss 0.334714f
C5019 FILLER_0_13_2/a_4964_472# vss 0.336371f
C5020 FILLER_0_13_2/a_4516_472# vss 0.338919f
C5021 FILLER_0_13_2/a_4068_472# vss 0.363279f
C5022 FILLER_0_13_2/a_3620_472# vss 0.343017f
C5023 FILLER_0_13_2/a_3172_472# vss 0.338197f
C5024 FILLER_0_13_2/a_2724_472# vss 0.337546f
C5025 FILLER_0_13_2/a_2276_472# vss 0.335717f
C5026 FILLER_0_13_2/a_1828_472# vss 0.333762f
C5027 FILLER_0_13_2/a_1380_472# vss 0.333762f
C5028 FILLER_0_13_2/a_932_472# vss 0.333762f
C5029 FILLER_0_13_2/a_484_472# vss 0.332506f
C5030 FILLER_0_13_2/a_36_472# vss 0.408581f
C5031 FILLER_0_13_2/a_6844_375# vss 0.291562f
C5032 FILLER_0_13_2/a_6396_375# vss 0.172168f
C5033 FILLER_0_13_2/a_5948_375# vss 0.171802f
C5034 FILLER_0_13_2/a_5500_375# vss 0.174928f
C5035 FILLER_0_13_2/a_5052_375# vss 0.17651f
C5036 FILLER_0_13_2/a_4604_375# vss 0.178722f
C5037 FILLER_0_13_2/a_4156_375# vss 0.191163f
C5038 FILLER_0_13_2/a_3708_375# vss 0.191898f
C5039 FILLER_0_13_2/a_3260_375# vss 0.178853f
C5040 FILLER_0_13_2/a_2812_375# vss 0.176722f
C5041 FILLER_0_13_2/a_2364_375# vss 0.175137f
C5042 FILLER_0_13_2/a_1916_375# vss 0.17209f
C5043 FILLER_0_13_2/a_1468_375# vss 0.17209f
C5044 FILLER_0_13_2/a_1020_375# vss 0.17209f
C5045 FILLER_0_13_2/a_572_375# vss 0.171927f
C5046 FILLER_0_13_2/a_124_375# vss 0.188994f
C5047 FILLER_0_0_12/a_1380_472# vss 0.351176f
C5048 FILLER_0_0_12/a_932_472# vss 0.332499f
C5049 FILLER_0_0_12/a_484_472# vss 0.33241f
C5050 FILLER_0_0_12/a_36_472# vss 0.406548f
C5051 FILLER_0_0_12/a_1468_375# vss 0.291133f
C5052 FILLER_0_0_12/a_1020_375# vss 0.172412f
C5053 FILLER_0_0_12/a_572_375# vss 0.171606f
C5054 FILLER_0_0_12/a_124_375# vss 0.185399f
C5055 FILLER_0_3_44/a_1380_472# vss 0.348697f
C5056 FILLER_0_3_44/a_932_472# vss 0.334777f
C5057 FILLER_0_3_44/a_484_472# vss 0.336616f
C5058 FILLER_0_3_44/a_36_472# vss 0.41167f
C5059 FILLER_0_3_44/a_1468_375# vss 0.287259f
C5060 FILLER_0_3_44/a_1020_375# vss 0.173184f
C5061 FILLER_0_3_44/a_572_375# vss 0.175752f
C5062 FILLER_0_3_44/a_124_375# vss 0.191478f
C5063 _12_/Z vss 1.360286f
C5064 _12_/a_36_113# vss 0.424895f
C5065 FILLER_0_15_56/a_484_472# vss 0.347509f
C5066 FILLER_0_15_56/a_36_472# vss 0.403547f
C5067 FILLER_0_15_56/a_572_375# vss 0.290693f
C5068 FILLER_0_15_56/a_124_375# vss 0.185465f
C5069 _13_/Z vss 1.333857f
C5070 _13_/a_36_113# vss 0.469366f
C5071 FILLER_0_2_101/a_36_472# vss 0.423771f
C5072 FILLER_0_2_101/a_124_375# vss 0.298976f
C5073 FILLER_0_12_12/a_1380_472# vss 0.352048f
C5074 FILLER_0_12_12/a_932_472# vss 0.33372f
C5075 FILLER_0_12_12/a_484_472# vss 0.33365f
C5076 FILLER_0_12_12/a_36_472# vss 0.407787f
C5077 FILLER_0_12_12/a_1468_375# vss 0.291881f
C5078 FILLER_0_12_12/a_1020_375# vss 0.172801f
C5079 FILLER_0_12_12/a_572_375# vss 0.172048f
C5080 FILLER_0_12_12/a_124_375# vss 0.185841f
C5081 input_signal[8] vss 1.234047f
C5082 _14_/Z vss 1.447568f
C5083 _14_/a_36_113# vss 0.426025f
C5084 FILLER_0_4_2/a_3172_472# vss 0.354187f
C5085 FILLER_0_4_2/a_2724_472# vss 0.336885f
C5086 FILLER_0_4_2/a_2276_472# vss 0.335244f
C5087 FILLER_0_4_2/a_1828_472# vss 0.333639f
C5088 FILLER_0_4_2/a_1380_472# vss 0.333639f
C5089 FILLER_0_4_2/a_932_472# vss 0.333639f
C5090 FILLER_0_4_2/a_484_472# vss 0.33241f
C5091 FILLER_0_4_2/a_36_472# vss 0.408673f
C5092 FILLER_0_4_2/a_3260_375# vss 0.266256f
C5093 FILLER_0_4_2/a_2812_375# vss 0.176466f
C5094 FILLER_0_4_2/a_2364_375# vss 0.174985f
C5095 FILLER_0_4_2/a_1916_375# vss 0.172109f
C5096 FILLER_0_4_2/a_1468_375# vss 0.172109f
C5097 FILLER_0_4_2/a_1020_375# vss 0.172109f
C5098 FILLER_0_4_2/a_572_375# vss 0.171953f
C5099 FILLER_0_4_2/a_124_375# vss 0.189405f
C5100 FILLER_0_15_2/a_36_472# vss 0.4231f
C5101 FILLER_0_15_2/a_124_375# vss 0.252646f
C5102 _15_/Z vss 1.428789f
C5103 _15_/a_36_113# vss 0.46837f
C5104 FILLER_0_6_107/a_36_472# vss 0.427063f
C5105 FILLER_0_6_107/a_124_375# vss 0.257842f
C5106 FILLER_0_9_104/a_484_472# vss 0.353529f
C5107 FILLER_0_9_104/a_36_472# vss 0.41165f
C5108 FILLER_0_9_104/a_572_375# vss 0.25109f
C5109 FILLER_0_9_104/a_124_375# vss 0.190801f
C5110 FILLER_0_9_72/a_3172_472# vss 0.351491f
C5111 FILLER_0_9_72/a_2724_472# vss 0.332816f
C5112 FILLER_0_9_72/a_2276_472# vss 0.333278f
C5113 FILLER_0_9_72/a_1828_472# vss 0.336049f
C5114 FILLER_0_9_72/a_1380_472# vss 0.337801f
C5115 FILLER_0_9_72/a_932_472# vss 0.340498f
C5116 FILLER_0_9_72/a_484_472# vss 0.371346f
C5117 FILLER_0_9_72/a_36_472# vss 0.415873f
C5118 FILLER_0_9_72/a_3260_375# vss 0.290708f
C5119 FILLER_0_9_72/a_2812_375# vss 0.171987f
C5120 FILLER_0_9_72/a_2364_375# vss 0.171987f
C5121 FILLER_0_9_72/a_1916_375# vss 0.175274f
C5122 FILLER_0_9_72/a_1468_375# vss 0.176943f
C5123 FILLER_0_9_72/a_1020_375# vss 0.179193f
C5124 FILLER_0_9_72/a_572_375# vss 0.198734f
C5125 FILLER_0_9_72/a_124_375# vss 0.200509f
C5126 FILLER_0_15_64/a_36_472# vss 0.421692f
C5127 FILLER_0_15_64/a_124_375# vss 0.268011f
C5128 _16_/Z vss 1.33333f
C5129 _16_/a_36_113# vss 0.423308f
C5130 FILLER_0_10_101/a_36_472# vss 0.423764f
C5131 FILLER_0_10_101/a_124_375# vss 0.298484f
C5132 FILLER_0_3_72/a_3172_472# vss 0.351491f
C5133 FILLER_0_3_72/a_2724_472# vss 0.332816f
C5134 FILLER_0_3_72/a_2276_472# vss 0.333278f
C5135 FILLER_0_3_72/a_1828_472# vss 0.336049f
C5136 FILLER_0_3_72/a_1380_472# vss 0.337801f
C5137 FILLER_0_3_72/a_932_472# vss 0.340498f
C5138 FILLER_0_3_72/a_484_472# vss 0.371425f
C5139 FILLER_0_3_72/a_36_472# vss 0.416116f
C5140 FILLER_0_3_72/a_3260_375# vss 0.290823f
C5141 FILLER_0_3_72/a_2812_375# vss 0.172103f
C5142 FILLER_0_3_72/a_2364_375# vss 0.172103f
C5143 FILLER_0_3_72/a_1916_375# vss 0.175389f
C5144 FILLER_0_3_72/a_1468_375# vss 0.176943f
C5145 FILLER_0_3_72/a_1020_375# vss 0.179193f
C5146 FILLER_0_3_72/a_572_375# vss 0.198976f
C5147 FILLER_0_3_72/a_124_375# vss 0.200509f
C5148 FILLER_0_8_28/a_36_472# vss 0.425794f
C5149 FILLER_0_8_28/a_124_375# vss 0.265502f
C5150 _17_/a_36_113# vss 0.426785f
C5151 FILLER_0_6_2/a_3172_472# vss 0.353745f
C5152 FILLER_0_6_2/a_2724_472# vss 0.336724f
C5153 FILLER_0_6_2/a_2276_472# vss 0.335214f
C5154 FILLER_0_6_2/a_1828_472# vss 0.333639f
C5155 FILLER_0_6_2/a_1380_472# vss 0.333639f
C5156 FILLER_0_6_2/a_932_472# vss 0.333639f
C5157 FILLER_0_6_2/a_484_472# vss 0.33241f
C5158 FILLER_0_6_2/a_36_472# vss 0.408673f
C5159 FILLER_0_6_2/a_3260_375# vss 0.265756f
C5160 FILLER_0_6_2/a_2812_375# vss 0.176144f
C5161 FILLER_0_6_2/a_2364_375# vss 0.174627f
C5162 FILLER_0_6_2/a_1916_375# vss 0.17167f
C5163 FILLER_0_6_2/a_1468_375# vss 0.17167f
C5164 FILLER_0_6_2/a_1020_375# vss 0.17167f
C5165 FILLER_0_6_2/a_572_375# vss 0.17167f
C5166 FILLER_0_6_2/a_124_375# vss 0.189122f
C5167 FILLER_0_15_40/a_1380_472# vss 0.348153f
C5168 FILLER_0_15_40/a_932_472# vss 0.333851f
C5169 FILLER_0_15_40/a_484_472# vss 0.335669f
C5170 FILLER_0_15_40/a_36_472# vss 0.411995f
C5171 FILLER_0_15_40/a_1468_375# vss 0.288579f
C5172 FILLER_0_15_40/a_1020_375# vss 0.175632f
C5173 FILLER_0_15_40/a_572_375# vss 0.177463f
C5174 FILLER_0_15_40/a_124_375# vss 0.193585f
C5175 _18_/a_36_113# vss 0.42374f
C5176 FILLER_0_3_60/a_484_472# vss 0.351448f
C5177 FILLER_0_3_60/a_36_472# vss 0.407263f
C5178 FILLER_0_3_60/a_572_375# vss 0.254892f
C5179 FILLER_0_3_60/a_124_375# vss 0.188112f
C5180 FILLER_0_14_107/a_484_472# vss 0.356469f
C5181 FILLER_0_14_107/a_36_472# vss 0.412998f
C5182 FILLER_0_14_107/a_572_375# vss 0.30533f
C5183 FILLER_0_14_107/a_124_375# vss 0.193359f
C5184 FILLER_0_15_72/a_1380_472# vss 0.3523f
C5185 FILLER_0_15_72/a_932_472# vss 0.339324f
C5186 FILLER_0_15_72/a_484_472# vss 0.368354f
C5187 FILLER_0_15_72/a_36_472# vss 0.4146f
C5188 FILLER_0_15_72/a_1468_375# vss 0.252733f
C5189 FILLER_0_15_72/a_1020_375# vss 0.178759f
C5190 FILLER_0_15_72/a_572_375# vss 0.197724f
C5191 FILLER_0_15_72/a_124_375# vss 0.198786f
C5192 _14_/I vss 3.171133f
C5193 FILLER_0_8_37/a_6756_472# vss 0.347527f
C5194 FILLER_0_8_37/a_6308_472# vss 0.331577f
C5195 FILLER_0_8_37/a_5860_472# vss 0.33412f
C5196 FILLER_0_8_37/a_5412_472# vss 0.335515f
C5197 FILLER_0_8_37/a_4964_472# vss 0.337674f
C5198 FILLER_0_8_37/a_4516_472# vss 0.355495f
C5199 FILLER_0_8_37/a_4068_472# vss 0.342266f
C5200 FILLER_0_8_37/a_3620_472# vss 0.339657f
C5201 FILLER_0_8_37/a_3172_472# vss 0.336286f
C5202 FILLER_0_8_37/a_2724_472# vss 0.335067f
C5203 FILLER_0_8_37/a_2276_472# vss 0.332816f
C5204 FILLER_0_8_37/a_1828_472# vss 0.333794f
C5205 FILLER_0_8_37/a_1380_472# vss 0.335804f
C5206 FILLER_0_8_37/a_932_472# vss 0.337458f
C5207 FILLER_0_8_37/a_484_472# vss 0.340073f
C5208 FILLER_0_8_37/a_36_472# vss 0.449284f
C5209 FILLER_0_8_37/a_6844_375# vss 0.288694f
C5210 FILLER_0_8_37/a_6396_375# vss 0.171802f
C5211 FILLER_0_8_37/a_5948_375# vss 0.174639f
C5212 FILLER_0_8_37/a_5500_375# vss 0.176062f
C5213 FILLER_0_8_37/a_5052_375# vss 0.178099f
C5214 FILLER_0_8_37/a_4604_375# vss 0.183886f
C5215 FILLER_0_8_37/a_4156_375# vss 0.198485f
C5216 FILLER_0_8_37/a_3708_375# vss 0.179135f
C5217 FILLER_0_8_37/a_3260_375# vss 0.176565f
C5218 FILLER_0_8_37/a_2812_375# vss 0.174986f
C5219 FILLER_0_8_37/a_2364_375# vss 0.171961f
C5220 FILLER_0_8_37/a_1916_375# vss 0.172079f
C5221 FILLER_0_8_37/a_1468_375# vss 0.175257f
C5222 FILLER_0_8_37/a_1020_375# vss 0.176926f
C5223 FILLER_0_8_37/a_572_375# vss 0.179058f
C5224 FILLER_0_8_37/a_124_375# vss 0.222024f
C5225 _19_/a_36_113# vss 0.443847f
C5226 FILLER_0_0_70/a_36_472# vss 0.428778f
C5227 FILLER_0_0_70/a_124_375# vss 0.266077f
C5228 FILLER_0_14_28/a_36_472# vss 0.426175f
C5229 FILLER_0_14_28/a_124_375# vss 0.264513f
C5230 FILLER_0_2_37/a_6756_472# vss 0.34747f
C5231 FILLER_0_2_37/a_6308_472# vss 0.331501f
C5232 FILLER_0_2_37/a_5860_472# vss 0.334411f
C5233 FILLER_0_2_37/a_5412_472# vss 0.336051f
C5234 FILLER_0_2_37/a_4964_472# vss 0.338426f
C5235 FILLER_0_2_37/a_4516_472# vss 0.357104f
C5236 FILLER_0_2_37/a_4068_472# vss 0.343998f
C5237 FILLER_0_2_37/a_3620_472# vss 0.340481f
C5238 FILLER_0_2_37/a_3172_472# vss 0.335573f
C5239 FILLER_0_2_37/a_2724_472# vss 0.334228f
C5240 FILLER_0_2_37/a_2276_472# vss 0.331611f
C5241 FILLER_0_2_37/a_1828_472# vss 0.332607f
C5242 FILLER_0_2_37/a_1380_472# vss 0.335021f
C5243 FILLER_0_2_37/a_932_472# vss 0.336867f
C5244 FILLER_0_2_37/a_484_472# vss 0.339691f
C5245 FILLER_0_2_37/a_36_472# vss 0.451256f
C5246 FILLER_0_2_37/a_6844_375# vss 0.288834f
C5247 FILLER_0_2_37/a_6396_375# vss 0.171802f
C5248 FILLER_0_2_37/a_5948_375# vss 0.174777f
C5249 FILLER_0_2_37/a_5500_375# vss 0.176273f
C5250 FILLER_0_2_37/a_5052_375# vss 0.178431f
C5251 FILLER_0_2_37/a_4604_375# vss 0.184694f
C5252 FILLER_0_2_37/a_4156_375# vss 0.200289f
C5253 FILLER_0_2_37/a_3708_375# vss 0.179566f
C5254 FILLER_0_2_37/a_3260_375# vss 0.17668f
C5255 FILLER_0_2_37/a_2812_375# vss 0.175008f
C5256 FILLER_0_2_37/a_2364_375# vss 0.171802f
C5257 FILLER_0_2_37/a_1916_375# vss 0.17192f
C5258 FILLER_0_2_37/a_1468_375# vss 0.175259f
C5259 FILLER_0_2_37/a_1020_375# vss 0.177017f
C5260 FILLER_0_2_37/a_572_375# vss 0.179288f
C5261 FILLER_0_2_37/a_124_375# vss 0.222892f
C5262 input_signal[9] vss 1.750877f
C5263 FILLER_0_3_104/a_484_472# vss 0.353529f
C5264 FILLER_0_3_104/a_36_472# vss 0.41165f
C5265 FILLER_0_3_104/a_572_375# vss 0.25109f
C5266 FILLER_0_3_104/a_124_375# vss 0.190916f
C5267 FILLER_0_6_101/a_36_472# vss 0.423318f
C5268 FILLER_0_6_101/a_124_375# vss 0.29886f
C5269 FILLER_0_14_115/a_36_472# vss 0.449039f
C5270 FILLER_0_14_115/a_124_375# vss 0.263041f
C5271 input9/a_36_113# vss 0.418606f
C5272 FILLER_0_8_12/a_1380_472# vss 0.352251f
C5273 FILLER_0_8_12/a_932_472# vss 0.333816f
C5274 FILLER_0_8_12/a_484_472# vss 0.333746f
C5275 FILLER_0_8_12/a_36_472# vss 0.407883f
C5276 FILLER_0_8_12/a_1468_375# vss 0.291783f
C5277 FILLER_0_8_12/a_1020_375# vss 0.172733f
C5278 FILLER_0_8_12/a_572_375# vss 0.172048f
C5279 FILLER_0_8_12/a_124_375# vss 0.185841f
C5280 FILLER_0_14_37/a_6756_472# vss 0.347546f
C5281 FILLER_0_14_37/a_6308_472# vss 0.331577f
C5282 FILLER_0_14_37/a_5860_472# vss 0.334391f
C5283 FILLER_0_14_37/a_5412_472# vss 0.335888f
C5284 FILLER_0_14_37/a_4964_472# vss 0.338157f
C5285 FILLER_0_14_37/a_4516_472# vss 0.355623f
C5286 FILLER_0_14_37/a_4068_472# vss 0.343211f
C5287 FILLER_0_14_37/a_3620_472# vss 0.340215f
C5288 FILLER_0_14_37/a_3172_472# vss 0.336709f
C5289 FILLER_0_14_37/a_2724_472# vss 0.335364f
C5290 FILLER_0_14_37/a_2276_472# vss 0.332816f
C5291 FILLER_0_14_37/a_1828_472# vss 0.333741f
C5292 FILLER_0_14_37/a_1380_472# vss 0.33611f
C5293 FILLER_0_14_37/a_932_472# vss 0.337873f
C5294 FILLER_0_14_37/a_484_472# vss 0.340592f
C5295 FILLER_0_14_37/a_36_472# vss 0.450529f
C5296 FILLER_0_14_37/a_6844_375# vss 0.288568f
C5297 FILLER_0_14_37/a_6396_375# vss 0.171644f
C5298 FILLER_0_14_37/a_5948_375# vss 0.174238f
C5299 FILLER_0_14_37/a_5500_375# vss 0.175724f
C5300 FILLER_0_14_37/a_5052_375# vss 0.177514f
C5301 FILLER_0_14_37/a_4604_375# vss 0.182367f
C5302 FILLER_0_14_37/a_4156_375# vss 0.197225f
C5303 FILLER_0_14_37/a_3708_375# vss 0.178641f
C5304 FILLER_0_14_37/a_3260_375# vss 0.176071f
C5305 FILLER_0_14_37/a_2812_375# vss 0.174653f
C5306 FILLER_0_14_37/a_2364_375# vss 0.171861f
C5307 FILLER_0_14_37/a_1916_375# vss 0.171963f
C5308 FILLER_0_14_37/a_1468_375# vss 0.174868f
C5309 FILLER_0_14_37/a_1020_375# vss 0.176352f
C5310 FILLER_0_14_37/a_572_375# vss 0.178212f
C5311 FILLER_0_14_37/a_124_375# vss 0.219478f
C5312 input8/a_36_113# vss 0.46218f
C5313 FILLER_0_5_12/a_3172_472# vss 0.356303f
C5314 FILLER_0_5_12/a_2724_472# vss 0.361652f
C5315 FILLER_0_5_12/a_2276_472# vss 0.337933f
C5316 FILLER_0_5_12/a_1828_472# vss 0.337516f
C5317 FILLER_0_5_12/a_1380_472# vss 0.336254f
C5318 FILLER_0_5_12/a_932_472# vss 0.333805f
C5319 FILLER_0_5_12/a_484_472# vss 0.333735f
C5320 FILLER_0_5_12/a_36_472# vss 0.407873f
C5321 FILLER_0_5_12/a_3260_375# vss 0.293977f
C5322 FILLER_0_5_12/a_2812_375# vss 0.217378f
C5323 FILLER_0_5_12/a_2364_375# vss 0.180111f
C5324 FILLER_0_5_12/a_1916_375# vss 0.177613f
C5325 FILLER_0_5_12/a_1468_375# vss 0.175736f
C5326 FILLER_0_5_12/a_1020_375# vss 0.172862f
C5327 FILLER_0_5_12/a_572_375# vss 0.172109f
C5328 FILLER_0_5_12/a_124_375# vss 0.186354f
C5329 input10/a_36_113# vss 0.462031f
C5330 FILLER_0_5_44/a_1380_472# vss 0.348731f
C5331 FILLER_0_5_44/a_932_472# vss 0.334518f
C5332 FILLER_0_5_44/a_484_472# vss 0.336007f
C5333 FILLER_0_5_44/a_36_472# vss 0.410642f
C5334 FILLER_0_5_44/a_1468_375# vss 0.287259f
C5335 FILLER_0_5_44/a_1020_375# vss 0.173184f
C5336 FILLER_0_5_44/a_572_375# vss 0.175659f
C5337 FILLER_0_5_44/a_124_375# vss 0.19132f
C5338 input7/a_36_113# vss 0.462188f
C5339 FILLER_0_0_104/a_36_472# vss 0.425761f
C5340 FILLER_0_0_104/a_124_375# vss 0.259262f
C5341 input_signal[5] vss 1.32071f
C5342 input6/a_36_113# vss 0.462188f
C5343 FILLER_0_14_101/a_36_472# vss 0.423764f
C5344 FILLER_0_14_101/a_124_375# vss 0.298325f
C5345 FILLER_0_14_12/a_1380_472# vss 0.352495f
C5346 FILLER_0_14_12/a_932_472# vss 0.333738f
C5347 FILLER_0_14_12/a_484_472# vss 0.33365f
C5348 FILLER_0_14_12/a_36_472# vss 0.407787f
C5349 FILLER_0_14_12/a_1468_375# vss 0.291063f
C5350 FILLER_0_14_12/a_1020_375# vss 0.172323f
C5351 FILLER_0_14_12/a_572_375# vss 0.171606f
C5352 FILLER_0_14_12/a_124_375# vss 0.185399f
C5353 FILLER_0_11_136/a_36_472# vss 0.421095f
C5354 FILLER_0_11_136/a_124_375# vss 0.295936f
C5355 input5/a_36_113# vss 0.462205f
C5356 _19_/I vss 2.157633f
C5357 input_signal[3] vss 1.010588f
C5358 input4/a_36_113# vss 0.462201f
C5359 FILLER_0_11_66/a_36_472# vss 0.425205f
C5360 FILLER_0_11_66/a_124_375# vss 0.300651f
C5361 _12_/I vss 2.384244f
C5362 input3/a_36_113# vss 0.462184f
C5363 _11_/I vss 3.38813f
C5364 input_signal[1] vss 1.077806f
C5365 input2/a_36_113# vss 0.461966f
C5366 FILLER_0_5_72/a_3172_472# vss 0.35102f
C5367 FILLER_0_5_72/a_2724_472# vss 0.332816f
C5368 FILLER_0_5_72/a_2276_472# vss 0.333243f
C5369 FILLER_0_5_72/a_1828_472# vss 0.335514f
C5370 FILLER_0_5_72/a_1380_472# vss 0.33692f
C5371 FILLER_0_5_72/a_932_472# vss 0.339102f
C5372 FILLER_0_5_72/a_484_472# vss 0.36718f
C5373 FILLER_0_5_72/a_36_472# vss 0.414431f
C5374 FILLER_0_5_72/a_3260_375# vss 0.290606f
C5375 FILLER_0_5_72/a_2812_375# vss 0.171987f
C5376 FILLER_0_5_72/a_2364_375# vss 0.171987f
C5377 FILLER_0_5_72/a_1916_375# vss 0.175196f
C5378 FILLER_0_5_72/a_1468_375# vss 0.176814f
C5379 FILLER_0_5_72/a_1020_375# vss 0.178972f
C5380 FILLER_0_5_72/a_572_375# vss 0.197898f
C5381 FILLER_0_5_72/a_124_375# vss 0.199772f
C5382 FILLER_0_4_107/a_1380_472# vss 0.350765f
C5383 FILLER_0_4_107/a_932_472# vss 0.361484f
C5384 FILLER_0_4_107/a_484_472# vss 0.340004f
C5385 FILLER_0_4_107/a_36_472# vss 0.412595f
C5386 FILLER_0_4_107/a_1468_375# vss 0.241948f
C5387 FILLER_0_4_107/a_1020_375# vss 0.190237f
C5388 FILLER_0_4_107/a_572_375# vss 0.189988f
C5389 FILLER_0_4_107/a_124_375# vss 0.19491f
C5390 _10_/I vss 1.83604f
C5391 input_signal[0] vss 1.802519f
C5392 input1/a_36_113# vss 0.46182f
C5393 _03_/ZN vss 1.204896f
C5394 FILLER_0_7_104/a_484_472# vss 0.352854f
C5395 FILLER_0_7_104/a_36_472# vss 0.41165f
C5396 FILLER_0_7_104/a_572_375# vss 0.244875f
C5397 FILLER_0_7_104/a_124_375# vss 0.190801f
C5398 FILLER_0_5_60/a_484_472# vss 0.35085f
C5399 FILLER_0_5_60/a_36_472# vss 0.407006f
C5400 FILLER_0_5_60/a_572_375# vss 0.254749f
C5401 FILLER_0_5_60/a_124_375# vss 0.188027f
C5402 FILLER_0_0_142/a_484_472# vss 0.353124f
C5403 FILLER_0_0_142/a_36_472# vss 0.409555f
C5404 FILLER_0_0_142/a_572_375# vss 0.258541f
C5405 FILLER_0_0_142/a_124_375# vss 0.188874f
C5406 _04_/ZN vss 1.185082f
C5407 input_signal[7] vss 1.044541f
C5408 FILLER_0_16_18/a_1380_472# vss 0.354861f
C5409 FILLER_0_16_18/a_932_472# vss 0.336984f
C5410 FILLER_0_16_18/a_484_472# vss 0.335341f
C5411 FILLER_0_16_18/a_36_472# vss 0.407893f
C5412 FILLER_0_16_18/a_1468_375# vss 0.28854f
C5413 FILLER_0_16_18/a_1020_375# vss 0.175963f
C5414 FILLER_0_16_18/a_572_375# vss 0.174482f
C5415 FILLER_0_16_18/a_124_375# vss 0.185399f
C5416 net15 vss 1.184586f
C5417 output_signal_minus[8] vss 1.122171f
C5418 _09_/ZN vss 2.178702f
C5419 output19/a_224_472# vss 2.431075f
C5420 _13_/I vss 2.759121f
C5421 FILLER_0_11_72/a_6756_472# vss 0.347154f
C5422 FILLER_0_11_72/a_6308_472# vss 0.333601f
C5423 FILLER_0_11_72/a_5860_472# vss 0.336647f
C5424 FILLER_0_11_72/a_5412_472# vss 0.337039f
C5425 FILLER_0_11_72/a_4964_472# vss 0.349809f
C5426 FILLER_0_11_72/a_4516_472# vss 0.350891f
C5427 FILLER_0_11_72/a_4068_472# vss 0.337824f
C5428 FILLER_0_11_72/a_3620_472# vss 0.338619f
C5429 FILLER_0_11_72/a_3172_472# vss 0.335611f
C5430 FILLER_0_11_72/a_2724_472# vss 0.332816f
C5431 FILLER_0_11_72/a_2276_472# vss 0.333278f
C5432 FILLER_0_11_72/a_1828_472# vss 0.336049f
C5433 FILLER_0_11_72/a_1380_472# vss 0.337801f
C5434 FILLER_0_11_72/a_932_472# vss 0.340498f
C5435 FILLER_0_11_72/a_484_472# vss 0.371351f
C5436 FILLER_0_11_72/a_36_472# vss 0.415779f
C5437 FILLER_0_11_72/a_6844_375# vss 0.288201f
C5438 FILLER_0_11_72/a_6396_375# vss 0.173472f
C5439 FILLER_0_11_72/a_5948_375# vss 0.176409f
C5440 FILLER_0_11_72/a_5500_375# vss 0.176994f
C5441 FILLER_0_11_72/a_5052_375# vss 0.181061f
C5442 FILLER_0_11_72/a_4604_375# vss 0.207297f
C5443 FILLER_0_11_72/a_4156_375# vss 0.179575f
C5444 FILLER_0_11_72/a_3708_375# vss 0.177356f
C5445 FILLER_0_11_72/a_3260_375# vss 0.175346f
C5446 FILLER_0_11_72/a_2812_375# vss 0.171961f
C5447 FILLER_0_11_72/a_2364_375# vss 0.171961f
C5448 FILLER_0_11_72/a_1916_375# vss 0.175248f
C5449 FILLER_0_11_72/a_1468_375# vss 0.176917f
C5450 FILLER_0_11_72/a_1020_375# vss 0.179167f
C5451 FILLER_0_11_72/a_572_375# vss 0.198686f
C5452 FILLER_0_11_72/a_124_375# vss 0.200072f
C5453 FILLER_0_4_37/a_6756_472# vss 0.347527f
C5454 FILLER_0_4_37/a_6308_472# vss 0.331577f
C5455 FILLER_0_4_37/a_5860_472# vss 0.33412f
C5456 FILLER_0_4_37/a_5412_472# vss 0.335515f
C5457 FILLER_0_4_37/a_4964_472# vss 0.337674f
C5458 FILLER_0_4_37/a_4516_472# vss 0.355451f
C5459 FILLER_0_4_37/a_4068_472# vss 0.34222f
C5460 FILLER_0_4_37/a_3620_472# vss 0.339657f
C5461 FILLER_0_4_37/a_3172_472# vss 0.335003f
C5462 FILLER_0_4_37/a_2724_472# vss 0.333827f
C5463 FILLER_0_4_37/a_2276_472# vss 0.331577f
C5464 FILLER_0_4_37/a_1828_472# vss 0.332554f
C5465 FILLER_0_4_37/a_1380_472# vss 0.334564f
C5466 FILLER_0_4_37/a_932_472# vss 0.336218f
C5467 FILLER_0_4_37/a_484_472# vss 0.338833f
C5468 FILLER_0_4_37/a_36_472# vss 0.447838f
C5469 FILLER_0_4_37/a_6844_375# vss 0.288694f
C5470 FILLER_0_4_37/a_6396_375# vss 0.171802f
C5471 FILLER_0_4_37/a_5948_375# vss 0.174639f
C5472 FILLER_0_4_37/a_5500_375# vss 0.176062f
C5473 FILLER_0_4_37/a_5052_375# vss 0.178099f
C5474 FILLER_0_4_37/a_4604_375# vss 0.183708f
C5475 FILLER_0_4_37/a_4156_375# vss 0.19827f
C5476 FILLER_0_4_37/a_3708_375# vss 0.179135f
C5477 FILLER_0_4_37/a_3260_375# vss 0.176395f
C5478 FILLER_0_4_37/a_2812_375# vss 0.174827f
C5479 FILLER_0_4_37/a_2364_375# vss 0.171802f
C5480 FILLER_0_4_37/a_1916_375# vss 0.17192f
C5481 FILLER_0_4_37/a_1468_375# vss 0.175098f
C5482 FILLER_0_4_37/a_1020_375# vss 0.176767f
C5483 FILLER_0_4_37/a_572_375# vss 0.178899f
C5484 FILLER_0_4_37/a_124_375# vss 0.221614f
C5485 output_signal_minus[7] vss 0.274217f
C5486 _08_/ZN vss 1.925324f
C5487 output18/a_224_472# vss 2.463949f
C5488 _15_/I vss 2.585433f
C5489 output_signal_plus[8] vss 0.64573f
C5490 _18_/Z vss 1.637627f
C5491 output29/a_224_472# vss 2.403936f
C5492 FILLER_0_12_107/a_1380_472# vss 0.35344f
C5493 FILLER_0_12_107/a_932_472# vss 0.361419f
C5494 FILLER_0_12_107/a_484_472# vss 0.339537f
C5495 FILLER_0_12_107/a_36_472# vss 0.412184f
C5496 FILLER_0_12_107/a_1468_375# vss 0.243384f
C5497 FILLER_0_12_107/a_1020_375# vss 0.190312f
C5498 FILLER_0_12_107/a_572_375# vss 0.190062f
C5499 FILLER_0_12_107/a_124_375# vss 0.195063f
C5500 FILLER_0_10_28/a_36_472# vss 0.426175f
C5501 FILLER_0_10_28/a_124_375# vss 0.264954f
C5502 output_signal_minus[6] vss 0.610572f
C5503 _07_/ZN vss 1.557929f
C5504 output17/a_224_472# vss 2.439832f
C5505 _16_/I vss 2.274916f
C5506 output_signal_plus[7] vss 0.809631f
C5507 _17_/Z vss 1.264877f
C5508 output28/a_224_472# vss 2.451366f
C5509 output_signal_minus[5] vss 0.420391f
C5510 _06_/ZN vss 1.278708f
C5511 output16/a_224_472# vss 2.411456f
C5512 output_signal_plus[6] vss 0.462068f
C5513 output27/a_224_472# vss 2.441884f
C5514 _17_/I vss 2.050051f
C5515 FILLER_0_16_36/a_3172_472# vss 0.349639f
C5516 FILLER_0_16_36/a_2724_472# vss 0.331571f
C5517 FILLER_0_16_36/a_2276_472# vss 0.330516f
C5518 FILLER_0_16_36/a_1828_472# vss 0.332273f
C5519 FILLER_0_16_36/a_1380_472# vss 0.333851f
C5520 FILLER_0_16_36/a_932_472# vss 0.335669f
C5521 FILLER_0_16_36/a_484_472# vss 0.338963f
C5522 FILLER_0_16_36/a_36_472# vss 0.432767f
C5523 FILLER_0_16_36/a_3260_375# vss 0.286106f
C5524 FILLER_0_16_36/a_2812_375# vss 0.174164f
C5525 FILLER_0_16_36/a_2364_375# vss 0.17167f
C5526 FILLER_0_16_36/a_1916_375# vss 0.172931f
C5527 FILLER_0_16_36/a_1468_375# vss 0.17532f
C5528 FILLER_0_16_36/a_1020_375# vss 0.177151f
C5529 FILLER_0_16_36/a_572_375# vss 0.179489f
C5530 FILLER_0_16_36/a_124_375# vss 0.22997f
C5531 FILLER_0_10_37/a_6756_472# vss 0.347546f
C5532 FILLER_0_10_37/a_6308_472# vss 0.331577f
C5533 FILLER_0_10_37/a_5860_472# vss 0.334391f
C5534 FILLER_0_10_37/a_5412_472# vss 0.335888f
C5535 FILLER_0_10_37/a_4964_472# vss 0.338157f
C5536 FILLER_0_10_37/a_4516_472# vss 0.355623f
C5537 FILLER_0_10_37/a_4068_472# vss 0.343211f
C5538 FILLER_0_10_37/a_3620_472# vss 0.340215f
C5539 FILLER_0_10_37/a_3172_472# vss 0.336709f
C5540 FILLER_0_10_37/a_2724_472# vss 0.335364f
C5541 FILLER_0_10_37/a_2276_472# vss 0.332816f
C5542 FILLER_0_10_37/a_1828_472# vss 0.333741f
C5543 FILLER_0_10_37/a_1380_472# vss 0.33611f
C5544 FILLER_0_10_37/a_932_472# vss 0.337873f
C5545 FILLER_0_10_37/a_484_472# vss 0.340592f
C5546 FILLER_0_10_37/a_36_472# vss 0.450529f
C5547 FILLER_0_10_37/a_6844_375# vss 0.288726f
C5548 FILLER_0_10_37/a_6396_375# vss 0.171802f
C5549 FILLER_0_10_37/a_5948_375# vss 0.174396f
C5550 FILLER_0_10_37/a_5500_375# vss 0.175669f
C5551 FILLER_0_10_37/a_5052_375# vss 0.17746f
C5552 FILLER_0_10_37/a_4604_375# vss 0.182472f
C5553 FILLER_0_10_37/a_4156_375# vss 0.197111f
C5554 FILLER_0_10_37/a_3708_375# vss 0.178495f
C5555 FILLER_0_10_37/a_3260_375# vss 0.176182f
C5556 FILLER_0_10_37/a_2812_375# vss 0.174753f
C5557 FILLER_0_10_37/a_2364_375# vss 0.171961f
C5558 FILLER_0_10_37/a_1916_375# vss 0.172063f
C5559 FILLER_0_10_37/a_1468_375# vss 0.174968f
C5560 FILLER_0_10_37/a_1020_375# vss 0.176452f
C5561 FILLER_0_10_37/a_572_375# vss 0.178313f
C5562 FILLER_0_10_37/a_124_375# vss 0.219307f
C5563 FILLER_0_7_66/a_36_472# vss 0.425205f
C5564 FILLER_0_7_66/a_124_375# vss 0.300709f
C5565 FILLER_0_4_101/a_36_472# vss 0.423424f
C5566 FILLER_0_4_101/a_124_375# vss 0.298762f
C5567 output_signal_minus[4] vss 0.438303f
C5568 output15/a_224_472# vss 2.457798f
C5569 _18_/I vss 2.388747f
C5570 output_signal_plus[5] vss 0.628454f
C5571 output26/a_224_472# vss 2.407613f
C5572 FILLER_0_1_12/a_3172_472# vss 0.358005f
C5573 FILLER_0_1_12/a_2724_472# vss 0.36501f
C5574 FILLER_0_1_12/a_2276_472# vss 0.339207f
C5575 FILLER_0_1_12/a_1828_472# vss 0.338282f
C5576 FILLER_0_1_12/a_1380_472# vss 0.336686f
C5577 FILLER_0_1_12/a_932_472# vss 0.333727f
C5578 FILLER_0_1_12/a_484_472# vss 0.333639f
C5579 FILLER_0_1_12/a_36_472# vss 0.407776f
C5580 FILLER_0_1_12/a_3260_375# vss 0.293945f
C5581 FILLER_0_1_12/a_2812_375# vss 0.217772f
C5582 FILLER_0_1_12/a_2364_375# vss 0.180752f
C5583 FILLER_0_1_12/a_1916_375# vss 0.177374f
C5584 FILLER_0_1_12/a_1468_375# vss 0.175414f
C5585 FILLER_0_1_12/a_1020_375# vss 0.172495f
C5586 FILLER_0_1_12/a_572_375# vss 0.17167f
C5587 FILLER_0_1_12/a_124_375# vss 0.185915f
C5588 output_signal_minus[3] vss 0.543172f
C5589 output14/a_224_472# vss 2.413605f
C5590 output_signal_plus[4] vss 0.442006f
C5591 output25/a_224_472# vss 2.415915f
C5592 FILLER_0_1_44/a_1380_472# vss 0.348697f
C5593 FILLER_0_1_44/a_932_472# vss 0.334777f
C5594 FILLER_0_1_44/a_484_472# vss 0.336616f
C5595 FILLER_0_1_44/a_36_472# vss 0.41167f
C5596 FILLER_0_1_44/a_1468_375# vss 0.286942f
C5597 FILLER_0_1_44/a_1020_375# vss 0.172867f
C5598 FILLER_0_1_44/a_572_375# vss 0.175435f
C5599 FILLER_0_1_44/a_124_375# vss 0.191161f
C5600 FILLER_0_7_2/a_6756_472# vss 0.350352f
C5601 FILLER_0_7_2/a_6308_472# vss 0.331577f
C5602 FILLER_0_7_2/a_5860_472# vss 0.331577f
C5603 FILLER_0_7_2/a_5412_472# vss 0.334643f
C5604 FILLER_0_7_2/a_4964_472# vss 0.336301f
C5605 FILLER_0_7_2/a_4516_472# vss 0.338848f
C5606 FILLER_0_7_2/a_4068_472# vss 0.363177f
C5607 FILLER_0_7_2/a_3620_472# vss 0.342921f
C5608 FILLER_0_7_2/a_3172_472# vss 0.338101f
C5609 FILLER_0_7_2/a_2724_472# vss 0.33745f
C5610 FILLER_0_7_2/a_2276_472# vss 0.335621f
C5611 FILLER_0_7_2/a_1828_472# vss 0.333666f
C5612 FILLER_0_7_2/a_1380_472# vss 0.333666f
C5613 FILLER_0_7_2/a_932_472# vss 0.333666f
C5614 FILLER_0_7_2/a_484_472# vss 0.33241f
C5615 FILLER_0_7_2/a_36_472# vss 0.408581f
C5616 FILLER_0_7_2/a_6844_375# vss 0.291708f
C5617 FILLER_0_7_2/a_6396_375# vss 0.172313f
C5618 FILLER_0_7_2/a_5948_375# vss 0.171946f
C5619 FILLER_0_7_2/a_5500_375# vss 0.175072f
C5620 FILLER_0_7_2/a_5052_375# vss 0.176654f
C5621 FILLER_0_7_2/a_4604_375# vss 0.178866f
C5622 FILLER_0_7_2/a_4156_375# vss 0.191332f
C5623 FILLER_0_7_2/a_3708_375# vss 0.192086f
C5624 FILLER_0_7_2/a_3260_375# vss 0.17857f
C5625 FILLER_0_7_2/a_2812_375# vss 0.17627f
C5626 FILLER_0_7_2/a_2364_375# vss 0.174691f
C5627 FILLER_0_7_2/a_1916_375# vss 0.171644f
C5628 FILLER_0_7_2/a_1468_375# vss 0.171644f
C5629 FILLER_0_7_2/a_1020_375# vss 0.171644f
C5630 FILLER_0_7_2/a_572_375# vss 0.171644f
C5631 FILLER_0_7_2/a_124_375# vss 0.18871f
C5632 output_signal_minus[2] vss 0.566155f
C5633 output13/a_224_472# vss 2.428023f
C5634 FILLER_0_8_107/a_484_472# vss 0.355546f
C5635 FILLER_0_8_107/a_36_472# vss 0.412454f
C5636 FILLER_0_8_107/a_572_375# vss 0.255691f
C5637 FILLER_0_8_107/a_124_375# vss 0.194287f
C5638 output_signal_plus[3] vss 0.604963f
C5639 output24/a_224_472# vss 2.405173f
C5640 FILLER_0_10_12/a_1380_472# vss 0.352495f
C5641 FILLER_0_10_12/a_932_472# vss 0.333738f
C5642 FILLER_0_10_12/a_484_472# vss 0.33365f
C5643 FILLER_0_10_12/a_36_472# vss 0.407787f
C5644 FILLER_0_10_12/a_1468_375# vss 0.291504f
C5645 FILLER_0_10_12/a_1020_375# vss 0.172765f
C5646 FILLER_0_10_12/a_572_375# vss 0.172048f
C5647 FILLER_0_10_12/a_124_375# vss 0.185841f
C5648 FILLER_0_13_66/a_36_472# vss 0.425239f
C5649 FILLER_0_13_66/a_124_375# vss 0.300651f
C5650 output_signal_minus[1] vss 0.580262f
C5651 _02_/ZN vss 1.150216f
C5652 output12/a_224_472# vss 2.407854f
C5653 output_signal_plus[2] vss 0.613956f
C5654 output23/a_224_472# vss 2.420832f
C5655 FILLER_0_12_101/a_36_472# vss 0.423318f
C5656 FILLER_0_12_101/a_124_375# vss 0.29886f
C5657 output_signal_minus[0] vss 2.173901f
C5658 _01_/ZN vss 1.536046f
C5659 output11/a_224_472# vss 2.409127f
C5660 output_signal_plus[1] vss 0.63321f
C5661 output22/a_224_472# vss 2.423755f
C5662 input_signal[2] vss 1.040925f
C5663 FILLER_0_7_72/a_3172_472# vss 0.351491f
C5664 FILLER_0_7_72/a_2724_472# vss 0.332816f
C5665 FILLER_0_7_72/a_2276_472# vss 0.333278f
C5666 FILLER_0_7_72/a_1828_472# vss 0.336049f
C5667 FILLER_0_7_72/a_1380_472# vss 0.337801f
C5668 FILLER_0_7_72/a_932_472# vss 0.340498f
C5669 FILLER_0_7_72/a_484_472# vss 0.371338f
C5670 FILLER_0_7_72/a_36_472# vss 0.415873f
C5671 FILLER_0_7_72/a_3260_375# vss 0.290708f
C5672 FILLER_0_7_72/a_2812_375# vss 0.171987f
C5673 FILLER_0_7_72/a_2364_375# vss 0.171987f
C5674 FILLER_0_7_72/a_1916_375# vss 0.175274f
C5675 FILLER_0_7_72/a_1468_375# vss 0.176943f
C5676 FILLER_0_7_72/a_1020_375# vss 0.179193f
C5677 FILLER_0_7_72/a_572_375# vss 0.198742f
C5678 FILLER_0_7_72/a_124_375# vss 0.200509f
C5679 FILLER_0_9_2/a_6756_472# vss 0.350352f
C5680 FILLER_0_9_2/a_6308_472# vss 0.331577f
C5681 FILLER_0_9_2/a_5860_472# vss 0.331577f
C5682 FILLER_0_9_2/a_5412_472# vss 0.334643f
C5683 FILLER_0_9_2/a_4964_472# vss 0.336301f
C5684 FILLER_0_9_2/a_4516_472# vss 0.338848f
C5685 FILLER_0_9_2/a_4068_472# vss 0.36318f
C5686 FILLER_0_9_2/a_3620_472# vss 0.342921f
C5687 FILLER_0_9_2/a_3172_472# vss 0.338101f
C5688 FILLER_0_9_2/a_2724_472# vss 0.33745f
C5689 FILLER_0_9_2/a_2276_472# vss 0.335621f
C5690 FILLER_0_9_2/a_1828_472# vss 0.333666f
C5691 FILLER_0_9_2/a_1380_472# vss 0.333666f
C5692 FILLER_0_9_2/a_932_472# vss 0.333666f
C5693 FILLER_0_9_2/a_484_472# vss 0.33241f
C5694 FILLER_0_9_2/a_36_472# vss 0.408581f
C5695 FILLER_0_9_2/a_6844_375# vss 0.291562f
C5696 FILLER_0_9_2/a_6396_375# vss 0.172168f
C5697 FILLER_0_9_2/a_5948_375# vss 0.171802f
C5698 FILLER_0_9_2/a_5500_375# vss 0.174928f
C5699 FILLER_0_9_2/a_5052_375# vss 0.17651f
C5700 FILLER_0_9_2/a_4604_375# vss 0.178722f
C5701 FILLER_0_9_2/a_4156_375# vss 0.191163f
C5702 FILLER_0_9_2/a_3708_375# vss 0.191898f
C5703 FILLER_0_9_2/a_3260_375# vss 0.178853f
C5704 FILLER_0_9_2/a_2812_375# vss 0.176722f
C5705 FILLER_0_9_2/a_2364_375# vss 0.175137f
C5706 FILLER_0_9_2/a_1916_375# vss 0.17209f
C5707 FILLER_0_9_2/a_1468_375# vss 0.17209f
C5708 FILLER_0_9_2/a_1020_375# vss 0.17209f
C5709 FILLER_0_9_2/a_572_375# vss 0.171927f
C5710 FILLER_0_9_2/a_124_375# vss 0.188994f
C5711 output_signal_plus[0] vss 1.372481f
C5712 _10_/Z vss 1.956451f
C5713 output21/a_224_472# vss 2.447125f
C5714 output_signal_minus[9] vss 0.550324f
C5715 _00_/ZN vss 3.111761f
C5716 output20/a_224_472# vss 2.438489f
C5717 FILLER_0_1_72/a_1380_472# vss 0.353259f
C5718 FILLER_0_1_72/a_932_472# vss 0.340498f
C5719 FILLER_0_1_72/a_484_472# vss 0.37141f
C5720 FILLER_0_1_72/a_36_472# vss 0.415882f
C5721 FILLER_0_1_72/a_1468_375# vss 0.252653f
C5722 FILLER_0_1_72/a_1020_375# vss 0.178811f
C5723 FILLER_0_1_72/a_572_375# vss 0.198504f
C5724 FILLER_0_1_72/a_124_375# vss 0.19949f
.ends

.subckt dac_in inputp inputm vss vdd input_signal[0] input_signal[1] input_signal[2]
+ input_signal[3] input_signal[4] input_signal[5] input_signal[6] input_signal[7]
+ input_signal[8] input_signal[9]
Xphase_inverter_0 input_signal[0] input_signal[1] input_signal[2] input_signal[3]
+ input_signal[4] input_signal[5] input_signal[9] carray_in_1/n1 carray_in_1/n2 carray_in_1/n3
+ carray_in_1/n4 carray_in_1/n5 carray_in_1/n6 carray_in_1/n7 carray_in_1/n8 carray_in_1/n9
+ carray_in_0/n1 carray_in_0/n2 carray_in_0/n3 carray_in_0/n4 carray_in_0/n5 carray_in_0/n6
+ carray_in_0/n7 phase_inverter_0/_10_/Z input_signal[7] phase_inverter_0/_19_/Z phase_inverter_0/FILLER_0_0_12/a_484_472#
+ phase_inverter_0/FILLER_0_0_36/a_2276_472# phase_inverter_0/_08_/ZN phase_inverter_0/FILLER_0_16_36/a_2364_375#
+ input_signal[8] phase_inverter_0/output18/a_224_472# phase_inverter_0/_19_/I phase_inverter_0/_00_/ZN
+ carray_in_0/n0 phase_inverter_0/_10_/I carray_in_0/n9 phase_inverter_0/FILLER_0_16_36/a_124_375#
+ phase_inverter_0/output20/a_224_472# phase_inverter_0/output30/a_224_472# input_signal[6]
+ phase_inverter_0/FILLER_0_0_36/a_36_472# phase_inverter_0/output21/a_224_472# phase_inverter_0/FILLER_0_16_18/a_124_375#
+ carray_in_1/n0 carray_in_0/n8 vdd vss phase_inverter
C0 carray_in_1/n0 carray_in_1/n3 0.047411f
C1 carray_in_0/n7 inputp 0.209952p
C2 inputp carray_in_0/n1 3.280347f
C3 inputp carray_in_0/n4 26.242765f
C4 carray_in_0/n5 carray_in_0/n0 0.025424f
C5 carray_in_0/n7 carray_in_0/n1 0.243006f
C6 carray_in_0/n7 carray_in_0/n4 1.70684f
C7 phase_inverter_0/_00_/ZN vdd 0.006089f
C8 carray_in_0/n1 carray_in_0/n4 0.145617f
C9 carray_in_0/n5 carray_in_0/n6 29.200403f
C10 carray_in_1/n0 carray_in_1/n1 8.401715f
C11 carray_in_0/n8 vdd 0.117452f
C12 carray_in_1/n0 carray_in_1/n5 0.025424f
C13 inputm carray_in_1/n2 6.560692f
C14 vdd phase_inverter_0/FILLER_0_16_36/a_2364_375# 0.004729f
C15 carray_in_0/n8 carray_in_0/n3 1.46349f
C16 carray_in_0/n0 carray_in_0/n2 0.089469f
C17 carray_in_1/n0 carray_in_1/n9 0.82611f
C18 carray_in_1/n0 carray_in_1/n6 0.025424f
C19 carray_in_0/n0 carray_in_0/n9 0.82611f
C20 carray_in_1/n0 carray_in_1/n8 0.097254f
C21 inputm carray_in_1/n7 0.209952p
C22 carray_in_0/n2 carray_in_0/n6 0.210444f
C23 carray_in_0/n6 carray_in_0/n9 14.718489f
C24 inputm carray_in_1/n4 26.242765f
C25 carray_in_1/n3 inputm 13.12139f
C26 inputp carray_in_0/n0 1.640173f
C27 carray_in_1/n7 carray_in_1/n2 0.487626f
C28 vdd phase_inverter_0/_08_/ZN 0.009745f
C29 phase_inverter_0/FILLER_0_16_18/a_124_375# vdd 0.004162f
C30 inputp carray_in_0/n6 0.104976p
C31 carray_in_1/n4 carray_in_1/n2 0.215946f
C32 carray_in_0/n7 carray_in_0/n0 0.06073f
C33 carray_in_0/n0 carray_in_0/n1 8.401715f
C34 carray_in_0/n0 carray_in_0/n4 0.03814f
C35 vdd phase_inverter_0/FILLER_0_0_12/a_484_472# 0.002838f
C36 carray_in_1/n3 carray_in_1/n2 23.465405f
C37 carray_in_1/n0 vdd 0.193605f
C38 carray_in_0/n7 carray_in_0/n6 34.900005f
C39 carray_in_0/n1 carray_in_0/n6 0.145088f
C40 carray_in_0/n4 carray_in_0/n6 0.617028f
C41 carray_in_0/n8 carray_in_0/n5 5.6103f
C42 inputm carray_in_1/n1 3.280347f
C43 carray_in_1/n4 carray_in_1/n7 1.70684f
C44 inputm carray_in_1/n5 52.485596f
C45 input_signal[0] vdd 0.001009f
C46 carray_in_0/n1 carray_in_1/n1 5.901133f
C47 carray_in_0/n5 carray_in_0/n3 0.350346f
C48 carray_in_1/n3 carray_in_1/n7 0.894213f
C49 phase_inverter_0/_19_/I vdd 0.002267f
C50 carray_in_1/n9 inputm 0.846091p
C51 inputm carray_in_1/n6 0.104976p
C52 carray_in_1/n3 carray_in_1/n4 26.505903f
C53 inputm carray_in_1/n8 0.420079p
C54 carray_in_1/n1 carray_in_1/n2 15.574605f
C55 carray_in_0/n8 carray_in_0/n2 0.772498f
C56 carray_in_1/n2 carray_in_1/n5 0.210974f
C57 carray_in_0/n8 carray_in_0/n9 87.65757f
C58 vdd carray_in_0/n9 0.358842f
C59 carray_in_0/n3 carray_in_0/n2 23.465405f
C60 carray_in_1/n9 carray_in_1/n2 0.997758f
C61 carray_in_1/n2 carray_in_1/n6 0.210444f
C62 carray_in_0/n3 carray_in_0/n9 1.912414f
C63 carray_in_1/n1 carray_in_1/n7 0.243006f
C64 carray_in_1/n8 carray_in_1/n2 0.772498f
C65 carray_in_1/n7 carray_in_1/n5 3.37237f
C66 vdd input_signal[9] 0.00119f
C67 carray_in_1/n4 carray_in_1/n1 0.145617f
C68 vdd phase_inverter_0/FILLER_0_0_36/a_2276_472# 0.004729f
C69 carray_in_1/n9 carray_in_1/n7 29.520088f
C70 carray_in_1/n7 carray_in_1/n6 34.900005f
C71 carray_in_1/n4 carray_in_1/n5 28.094206f
C72 carray_in_0/n8 inputp 0.420079p
C73 carray_in_1/n3 carray_in_1/n1 0.148119f
C74 phase_inverter_0/_10_/I vdd 0.023473f
C75 carray_in_1/n8 carray_in_1/n7 50.742203f
C76 carray_in_1/n3 carray_in_1/n5 0.350346f
C77 carray_in_0/n0 carray_in_0/n6 0.025424f
C78 inputp carray_in_0/n3 13.12139f
C79 carray_in_1/n9 carray_in_1/n4 3.741774f
C80 carray_in_1/n4 carray_in_1/n6 0.617028f
C81 carray_in_0/n8 carray_in_0/n7 50.742203f
C82 carray_in_0/n8 carray_in_0/n1 0.333459f
C83 carray_in_0/n8 carray_in_0/n4 2.84594f
C84 carray_in_1/n9 carray_in_1/n3 1.912414f
C85 carray_in_1/n3 carray_in_1/n6 0.339322f
C86 carray_in_1/n8 carray_in_1/n4 2.84594f
C87 phase_inverter_0/_19_/Z vdd 0.005964f
C88 carray_in_0/n7 carray_in_0/n3 0.894213f
C89 carray_in_0/n3 carray_in_0/n1 0.148119f
C90 carray_in_0/n3 carray_in_0/n4 26.505903f
C91 carray_in_1/n3 carray_in_1/n8 1.46349f
C92 carray_in_1/n1 carray_in_1/n5 0.145556f
C93 carray_in_0/n5 carray_in_0/n2 0.210974f
C94 vdd phase_inverter_0/_10_/Z 0.003245f
C95 carray_in_0/n5 carray_in_0/n9 7.400846f
C96 carray_in_1/n9 carray_in_1/n1 0.39415f
C97 carray_in_1/n1 carray_in_1/n6 0.145088f
C98 carray_in_1/n9 carray_in_1/n5 7.400846f
C99 carray_in_1/n6 carray_in_1/n5 29.200403f
C100 carray_in_1/n8 carray_in_1/n1 0.333459f
C101 carray_in_1/n8 carray_in_1/n5 5.6103f
C102 carray_in_1/n9 carray_in_1/n6 14.718489f
C103 carray_in_1/n9 carray_in_1/n8 87.65758f
C104 carray_in_1/n8 carray_in_1/n6 11.2197f
C105 carray_in_0/n5 inputp 52.485596f
C106 carray_in_0/n2 carray_in_0/n9 0.997758f
C107 carray_in_1/n0 inputm 1.640173f
C108 carray_in_0/n8 carray_in_0/n0 0.097254f
C109 vdd carray_in_0/n0 0.177806f
C110 carray_in_0/n5 carray_in_0/n7 3.37237f
C111 carray_in_0/n5 carray_in_0/n1 0.145556f
C112 carray_in_0/n5 carray_in_0/n4 28.094206f
C113 carray_in_0/n3 carray_in_0/n0 0.047411f
C114 carray_in_0/n8 carray_in_0/n6 11.2197f
C115 inputp carray_in_0/n2 6.560692f
C116 carray_in_1/n0 carray_in_1/n2 0.089469f
C117 carray_in_0/n3 carray_in_0/n6 0.339322f
C118 inputp carray_in_0/n9 0.846091p
C119 carray_in_0/n7 carray_in_0/n2 0.487626f
C120 carray_in_0/n2 carray_in_0/n1 15.574605f
C121 carray_in_0/n2 carray_in_0/n4 0.215946f
C122 vdd carray_in_1/n9 0.348295f
C123 carray_in_1/n0 carray_in_1/n7 0.06073f
C124 carray_in_0/n7 carray_in_0/n9 29.520088f
C125 carray_in_0/n1 carray_in_0/n9 0.39415f
C126 carray_in_0/n4 carray_in_0/n9 3.741774f
C127 vdd carray_in_1/n8 0.021439f
C128 carray_in_1/n0 carray_in_1/n4 0.03814f
C129 phase_inverter_0/_19_/Z vss 1.174253f
C130 phase_inverter_0/output30/a_224_472# vss 2.386102f
C131 phase_inverter_0/FILLER_0_1_60/a_484_472# vss 0.345058f
C132 phase_inverter_0/FILLER_0_1_60/a_36_472# vss 0.404746f
C133 phase_inverter_0/FILLER_0_1_60/a_572_375# vss 0.232991f
C134 phase_inverter_0/FILLER_0_1_60/a_124_375# vss 0.185089f
C135 phase_inverter_0/FILLER_0_0_28/a_36_472# vss 0.417394f
C136 phase_inverter_0/FILLER_0_0_28/a_124_375# vss 0.246306f
C137 phase_inverter_0/FILLER_0_13_72/a_3172_472# vss 0.345058f
C138 phase_inverter_0/FILLER_0_13_72/a_2724_472# vss 0.33241f
C139 phase_inverter_0/FILLER_0_13_72/a_2276_472# vss 0.33241f
C140 phase_inverter_0/FILLER_0_13_72/a_1828_472# vss 0.33241f
C141 phase_inverter_0/FILLER_0_13_72/a_1380_472# vss 0.33241f
C142 phase_inverter_0/FILLER_0_13_72/a_932_472# vss 0.33241f
C143 phase_inverter_0/FILLER_0_13_72/a_484_472# vss 0.33241f
C144 phase_inverter_0/FILLER_0_13_72/a_36_472# vss 0.404746f
C145 phase_inverter_0/FILLER_0_13_72/a_3260_375# vss 0.233093f
C146 phase_inverter_0/FILLER_0_13_72/a_2812_375# vss 0.17167f
C147 phase_inverter_0/FILLER_0_13_72/a_2364_375# vss 0.17167f
C148 phase_inverter_0/FILLER_0_13_72/a_1916_375# vss 0.17167f
C149 phase_inverter_0/FILLER_0_13_72/a_1468_375# vss 0.17167f
C150 phase_inverter_0/FILLER_0_13_72/a_1020_375# vss 0.17167f
C151 phase_inverter_0/FILLER_0_13_72/a_572_375# vss 0.17167f
C152 phase_inverter_0/FILLER_0_13_72/a_124_375# vss 0.185915f
C153 phase_inverter_0/FILLER_0_2_107/a_1380_472# vss 0.345058f
C154 phase_inverter_0/FILLER_0_2_107/a_932_472# vss 0.33241f
C155 phase_inverter_0/FILLER_0_2_107/a_484_472# vss 0.33241f
C156 phase_inverter_0/FILLER_0_2_107/a_36_472# vss 0.404746f
C157 phase_inverter_0/FILLER_0_2_107/a_1468_375# vss 0.233029f
C158 phase_inverter_0/FILLER_0_2_107/a_1020_375# vss 0.171606f
C159 phase_inverter_0/FILLER_0_2_107/a_572_375# vss 0.171606f
C160 phase_inverter_0/FILLER_0_2_107/a_124_375# vss 0.185399f
C161 phase_inverter_0/FILLER_0_5_104/a_484_472# vss 0.345058f
C162 phase_inverter_0/FILLER_0_5_104/a_36_472# vss 0.404746f
C163 phase_inverter_0/FILLER_0_5_104/a_572_375# vss 0.232991f
C164 phase_inverter_0/FILLER_0_5_104/a_124_375# vss 0.185089f
C165 phase_inverter_0/FILLER_0_6_37/a_6756_472# vss 0.345058f
C166 phase_inverter_0/FILLER_0_6_37/a_6308_472# vss 0.33241f
C167 phase_inverter_0/FILLER_0_6_37/a_5860_472# vss 0.33241f
C168 phase_inverter_0/FILLER_0_6_37/a_5412_472# vss 0.33241f
C169 phase_inverter_0/FILLER_0_6_37/a_4964_472# vss 0.33241f
C170 phase_inverter_0/FILLER_0_6_37/a_4516_472# vss 0.33241f
C171 phase_inverter_0/FILLER_0_6_37/a_4068_472# vss 0.33241f
C172 phase_inverter_0/FILLER_0_6_37/a_3620_472# vss 0.33241f
C173 phase_inverter_0/FILLER_0_6_37/a_3172_472# vss 0.33241f
C174 phase_inverter_0/FILLER_0_6_37/a_2724_472# vss 0.33241f
C175 phase_inverter_0/FILLER_0_6_37/a_2276_472# vss 0.33241f
C176 phase_inverter_0/FILLER_0_6_37/a_1828_472# vss 0.33241f
C177 phase_inverter_0/FILLER_0_6_37/a_1380_472# vss 0.33241f
C178 phase_inverter_0/FILLER_0_6_37/a_932_472# vss 0.33241f
C179 phase_inverter_0/FILLER_0_6_37/a_484_472# vss 0.33241f
C180 phase_inverter_0/FILLER_0_6_37/a_36_472# vss 0.404746f
C181 phase_inverter_0/FILLER_0_6_37/a_6844_375# vss 0.233068f
C182 phase_inverter_0/FILLER_0_6_37/a_6396_375# vss 0.171644f
C183 phase_inverter_0/FILLER_0_6_37/a_5948_375# vss 0.171644f
C184 phase_inverter_0/FILLER_0_6_37/a_5500_375# vss 0.171644f
C185 phase_inverter_0/FILLER_0_6_37/a_5052_375# vss 0.171644f
C186 phase_inverter_0/FILLER_0_6_37/a_4604_375# vss 0.171644f
C187 phase_inverter_0/FILLER_0_6_37/a_4156_375# vss 0.171644f
C188 phase_inverter_0/FILLER_0_6_37/a_3708_375# vss 0.171644f
C189 phase_inverter_0/FILLER_0_6_37/a_3260_375# vss 0.171644f
C190 phase_inverter_0/FILLER_0_6_37/a_2812_375# vss 0.171644f
C191 phase_inverter_0/FILLER_0_6_37/a_2364_375# vss 0.171644f
C192 phase_inverter_0/FILLER_0_6_37/a_1916_375# vss 0.171644f
C193 phase_inverter_0/FILLER_0_6_37/a_1468_375# vss 0.171644f
C194 phase_inverter_0/FILLER_0_6_37/a_1020_375# vss 0.171644f
C195 phase_inverter_0/FILLER_0_6_37/a_572_375# vss 0.171644f
C196 phase_inverter_0/FILLER_0_6_37/a_124_375# vss 0.185708f
C197 input_signal[4] vss 1.095436f
C198 phase_inverter_0/FILLER_0_8_101/a_36_472# vss 0.417394f
C199 phase_inverter_0/FILLER_0_8_101/a_124_375# vss 0.246306f
C200 phase_inverter_0/FILLER_0_16_104/a_36_472# vss 0.417394f
C201 phase_inverter_0/FILLER_0_16_104/a_124_375# vss 0.246306f
C202 phase_inverter_0/FILLER_0_12_28/a_36_472# vss 0.417394f
C203 phase_inverter_0/FILLER_0_12_28/a_124_375# vss 0.246306f
C204 phase_inverter_0/FILLER_0_11_2/a_6756_472# vss 0.345058f
C205 phase_inverter_0/FILLER_0_11_2/a_6308_472# vss 0.33241f
C206 phase_inverter_0/FILLER_0_11_2/a_5860_472# vss 0.33241f
C207 phase_inverter_0/FILLER_0_11_2/a_5412_472# vss 0.33241f
C208 phase_inverter_0/FILLER_0_11_2/a_4964_472# vss 0.33241f
C209 phase_inverter_0/FILLER_0_11_2/a_4516_472# vss 0.33241f
C210 phase_inverter_0/FILLER_0_11_2/a_4068_472# vss 0.33241f
C211 phase_inverter_0/FILLER_0_11_2/a_3620_472# vss 0.33241f
C212 phase_inverter_0/FILLER_0_11_2/a_3172_472# vss 0.33241f
C213 phase_inverter_0/FILLER_0_11_2/a_2724_472# vss 0.33241f
C214 phase_inverter_0/FILLER_0_11_2/a_2276_472# vss 0.33241f
C215 phase_inverter_0/FILLER_0_11_2/a_1828_472# vss 0.33241f
C216 phase_inverter_0/FILLER_0_11_2/a_1380_472# vss 0.33241f
C217 phase_inverter_0/FILLER_0_11_2/a_932_472# vss 0.33241f
C218 phase_inverter_0/FILLER_0_11_2/a_484_472# vss 0.33241f
C219 phase_inverter_0/FILLER_0_11_2/a_36_472# vss 0.404746f
C220 phase_inverter_0/FILLER_0_11_2/a_6844_375# vss 0.233068f
C221 phase_inverter_0/FILLER_0_11_2/a_6396_375# vss 0.171644f
C222 phase_inverter_0/FILLER_0_11_2/a_5948_375# vss 0.171644f
C223 phase_inverter_0/FILLER_0_11_2/a_5500_375# vss 0.171644f
C224 phase_inverter_0/FILLER_0_11_2/a_5052_375# vss 0.171644f
C225 phase_inverter_0/FILLER_0_11_2/a_4604_375# vss 0.171644f
C226 phase_inverter_0/FILLER_0_11_2/a_4156_375# vss 0.171644f
C227 phase_inverter_0/FILLER_0_11_2/a_3708_375# vss 0.171644f
C228 phase_inverter_0/FILLER_0_11_2/a_3260_375# vss 0.171644f
C229 phase_inverter_0/FILLER_0_11_2/a_2812_375# vss 0.171644f
C230 phase_inverter_0/FILLER_0_11_2/a_2364_375# vss 0.171644f
C231 phase_inverter_0/FILLER_0_11_2/a_1916_375# vss 0.171644f
C232 phase_inverter_0/FILLER_0_11_2/a_1468_375# vss 0.171644f
C233 phase_inverter_0/FILLER_0_11_2/a_1020_375# vss 0.171644f
C234 phase_inverter_0/FILLER_0_11_2/a_572_375# vss 0.171644f
C235 phase_inverter_0/FILLER_0_11_2/a_124_375# vss 0.185708f
C236 phase_inverter_0/FILLER_0_16_70/a_36_472# vss 0.417394f
C237 phase_inverter_0/FILLER_0_16_70/a_124_375# vss 0.246306f
C238 phase_inverter_0/FILLER_0_15_8/a_3172_472# vss 0.345058f
C239 phase_inverter_0/FILLER_0_15_8/a_2724_472# vss 0.33241f
C240 phase_inverter_0/FILLER_0_15_8/a_2276_472# vss 0.33241f
C241 phase_inverter_0/FILLER_0_15_8/a_1828_472# vss 0.33241f
C242 phase_inverter_0/FILLER_0_15_8/a_1380_472# vss 0.33241f
C243 phase_inverter_0/FILLER_0_15_8/a_932_472# vss 0.33241f
C244 phase_inverter_0/FILLER_0_15_8/a_484_472# vss 0.33241f
C245 phase_inverter_0/FILLER_0_15_8/a_36_472# vss 0.404746f
C246 phase_inverter_0/FILLER_0_15_8/a_3260_375# vss 0.233093f
C247 phase_inverter_0/FILLER_0_15_8/a_2812_375# vss 0.17167f
C248 phase_inverter_0/FILLER_0_15_8/a_2364_375# vss 0.17167f
C249 phase_inverter_0/FILLER_0_15_8/a_1916_375# vss 0.17167f
C250 phase_inverter_0/FILLER_0_15_8/a_1468_375# vss 0.17167f
C251 phase_inverter_0/FILLER_0_15_8/a_1020_375# vss 0.17167f
C252 phase_inverter_0/FILLER_0_15_8/a_572_375# vss 0.17167f
C253 phase_inverter_0/FILLER_0_15_8/a_124_375# vss 0.185915f
C254 vdd vss 0.426348p
C255 phase_inverter_0/FILLER_0_0_36/a_3172_472# vss 0.345058f
C256 phase_inverter_0/FILLER_0_0_36/a_2724_472# vss 0.33241f
C257 phase_inverter_0/FILLER_0_0_36/a_2276_472# vss 0.33241f
C258 phase_inverter_0/FILLER_0_0_36/a_1828_472# vss 0.33241f
C259 phase_inverter_0/FILLER_0_0_36/a_1380_472# vss 0.33241f
C260 phase_inverter_0/FILLER_0_0_36/a_932_472# vss 0.33241f
C261 phase_inverter_0/FILLER_0_0_36/a_484_472# vss 0.33241f
C262 phase_inverter_0/FILLER_0_0_36/a_36_472# vss 0.409475f
C263 phase_inverter_0/FILLER_0_0_36/a_3260_375# vss 0.233093f
C264 phase_inverter_0/FILLER_0_0_36/a_2812_375# vss 0.17167f
C265 phase_inverter_0/FILLER_0_0_36/a_2364_375# vss 0.17167f
C266 phase_inverter_0/FILLER_0_0_36/a_1916_375# vss 0.17167f
C267 phase_inverter_0/FILLER_0_0_36/a_1468_375# vss 0.17167f
C268 phase_inverter_0/FILLER_0_0_36/a_1020_375# vss 0.17167f
C269 phase_inverter_0/FILLER_0_0_36/a_572_375# vss 0.17167f
C270 phase_inverter_0/FILLER_0_0_36/a_124_375# vss 0.185915f
C271 phase_inverter_0/_10_/a_36_160# vss 0.386641f
C272 phase_inverter_0/FILLER_0_10_107/a_1380_472# vss 0.345058f
C273 phase_inverter_0/FILLER_0_10_107/a_932_472# vss 0.33241f
C274 phase_inverter_0/FILLER_0_10_107/a_484_472# vss 0.33241f
C275 phase_inverter_0/FILLER_0_10_107/a_36_472# vss 0.404746f
C276 phase_inverter_0/FILLER_0_10_107/a_1468_375# vss 0.233029f
C277 phase_inverter_0/FILLER_0_10_107/a_1020_375# vss 0.171606f
C278 phase_inverter_0/FILLER_0_10_107/a_572_375# vss 0.171606f
C279 phase_inverter_0/FILLER_0_10_107/a_124_375# vss 0.185399f
C280 phase_inverter_0/FILLER_0_12_37/a_6756_472# vss 0.345058f
C281 phase_inverter_0/FILLER_0_12_37/a_6308_472# vss 0.33241f
C282 phase_inverter_0/FILLER_0_12_37/a_5860_472# vss 0.33241f
C283 phase_inverter_0/FILLER_0_12_37/a_5412_472# vss 0.33241f
C284 phase_inverter_0/FILLER_0_12_37/a_4964_472# vss 0.33241f
C285 phase_inverter_0/FILLER_0_12_37/a_4516_472# vss 0.33241f
C286 phase_inverter_0/FILLER_0_12_37/a_4068_472# vss 0.33241f
C287 phase_inverter_0/FILLER_0_12_37/a_3620_472# vss 0.33241f
C288 phase_inverter_0/FILLER_0_12_37/a_3172_472# vss 0.33241f
C289 phase_inverter_0/FILLER_0_12_37/a_2724_472# vss 0.33241f
C290 phase_inverter_0/FILLER_0_12_37/a_2276_472# vss 0.33241f
C291 phase_inverter_0/FILLER_0_12_37/a_1828_472# vss 0.33241f
C292 phase_inverter_0/FILLER_0_12_37/a_1380_472# vss 0.33241f
C293 phase_inverter_0/FILLER_0_12_37/a_932_472# vss 0.33241f
C294 phase_inverter_0/FILLER_0_12_37/a_484_472# vss 0.33241f
C295 phase_inverter_0/FILLER_0_12_37/a_36_472# vss 0.404746f
C296 phase_inverter_0/FILLER_0_12_37/a_6844_375# vss 0.233068f
C297 phase_inverter_0/FILLER_0_12_37/a_6396_375# vss 0.171644f
C298 phase_inverter_0/FILLER_0_12_37/a_5948_375# vss 0.171644f
C299 phase_inverter_0/FILLER_0_12_37/a_5500_375# vss 0.171644f
C300 phase_inverter_0/FILLER_0_12_37/a_5052_375# vss 0.171644f
C301 phase_inverter_0/FILLER_0_12_37/a_4604_375# vss 0.171644f
C302 phase_inverter_0/FILLER_0_12_37/a_4156_375# vss 0.171644f
C303 phase_inverter_0/FILLER_0_12_37/a_3708_375# vss 0.171644f
C304 phase_inverter_0/FILLER_0_12_37/a_3260_375# vss 0.171644f
C305 phase_inverter_0/FILLER_0_12_37/a_2812_375# vss 0.171644f
C306 phase_inverter_0/FILLER_0_12_37/a_2364_375# vss 0.171644f
C307 phase_inverter_0/FILLER_0_12_37/a_1916_375# vss 0.171644f
C308 phase_inverter_0/FILLER_0_12_37/a_1468_375# vss 0.171644f
C309 phase_inverter_0/FILLER_0_12_37/a_1020_375# vss 0.171644f
C310 phase_inverter_0/FILLER_0_12_37/a_572_375# vss 0.171644f
C311 phase_inverter_0/FILLER_0_12_37/a_124_375# vss 0.185708f
C312 phase_inverter_0/FILLER_0_13_104/a_484_472# vss 0.345058f
C313 phase_inverter_0/FILLER_0_13_104/a_36_472# vss 0.404746f
C314 phase_inverter_0/FILLER_0_13_104/a_572_375# vss 0.232991f
C315 phase_inverter_0/FILLER_0_13_104/a_124_375# vss 0.185089f
C316 input_signal[6] vss 1.014523f
C317 phase_inverter_0/_11_/Z vss 1.137333f
C318 phase_inverter_0/_11_/a_36_113# vss 0.418095f
C319 phase_inverter_0/FILLER_0_9_66/a_36_472# vss 0.417394f
C320 phase_inverter_0/FILLER_0_9_66/a_124_375# vss 0.246306f
C321 phase_inverter_0/FILLER_0_3_12/a_3172_472# vss 0.345058f
C322 phase_inverter_0/FILLER_0_3_12/a_2724_472# vss 0.33241f
C323 phase_inverter_0/FILLER_0_3_12/a_2276_472# vss 0.33241f
C324 phase_inverter_0/FILLER_0_3_12/a_1828_472# vss 0.33241f
C325 phase_inverter_0/FILLER_0_3_12/a_1380_472# vss 0.33241f
C326 phase_inverter_0/FILLER_0_3_12/a_932_472# vss 0.33241f
C327 phase_inverter_0/FILLER_0_3_12/a_484_472# vss 0.33241f
C328 phase_inverter_0/FILLER_0_3_12/a_36_472# vss 0.404746f
C329 phase_inverter_0/FILLER_0_3_12/a_3260_375# vss 0.233093f
C330 phase_inverter_0/FILLER_0_3_12/a_2812_375# vss 0.17167f
C331 phase_inverter_0/FILLER_0_3_12/a_2364_375# vss 0.17167f
C332 phase_inverter_0/FILLER_0_3_12/a_1916_375# vss 0.17167f
C333 phase_inverter_0/FILLER_0_3_12/a_1468_375# vss 0.17167f
C334 phase_inverter_0/FILLER_0_3_12/a_1020_375# vss 0.17167f
C335 phase_inverter_0/FILLER_0_3_12/a_572_375# vss 0.17167f
C336 phase_inverter_0/FILLER_0_3_12/a_124_375# vss 0.185915f
C337 phase_inverter_0/FILLER_0_2_2/a_3172_472# vss 0.345058f
C338 phase_inverter_0/FILLER_0_2_2/a_2724_472# vss 0.33241f
C339 phase_inverter_0/FILLER_0_2_2/a_2276_472# vss 0.33241f
C340 phase_inverter_0/FILLER_0_2_2/a_1828_472# vss 0.33241f
C341 phase_inverter_0/FILLER_0_2_2/a_1380_472# vss 0.33241f
C342 phase_inverter_0/FILLER_0_2_2/a_932_472# vss 0.33241f
C343 phase_inverter_0/FILLER_0_2_2/a_484_472# vss 0.33241f
C344 phase_inverter_0/FILLER_0_2_2/a_36_472# vss 0.404746f
C345 phase_inverter_0/FILLER_0_2_2/a_3260_375# vss 0.233093f
C346 phase_inverter_0/FILLER_0_2_2/a_2812_375# vss 0.17167f
C347 phase_inverter_0/FILLER_0_2_2/a_2364_375# vss 0.17167f
C348 phase_inverter_0/FILLER_0_2_2/a_1916_375# vss 0.17167f
C349 phase_inverter_0/FILLER_0_2_2/a_1468_375# vss 0.17167f
C350 phase_inverter_0/FILLER_0_2_2/a_1020_375# vss 0.17167f
C351 phase_inverter_0/FILLER_0_2_2/a_572_375# vss 0.17167f
C352 phase_inverter_0/FILLER_0_2_2/a_124_375# vss 0.185915f
C353 phase_inverter_0/FILLER_0_13_2/a_6756_472# vss 0.345058f
C354 phase_inverter_0/FILLER_0_13_2/a_6308_472# vss 0.33241f
C355 phase_inverter_0/FILLER_0_13_2/a_5860_472# vss 0.33241f
C356 phase_inverter_0/FILLER_0_13_2/a_5412_472# vss 0.33241f
C357 phase_inverter_0/FILLER_0_13_2/a_4964_472# vss 0.33241f
C358 phase_inverter_0/FILLER_0_13_2/a_4516_472# vss 0.33241f
C359 phase_inverter_0/FILLER_0_13_2/a_4068_472# vss 0.33241f
C360 phase_inverter_0/FILLER_0_13_2/a_3620_472# vss 0.33241f
C361 phase_inverter_0/FILLER_0_13_2/a_3172_472# vss 0.33241f
C362 phase_inverter_0/FILLER_0_13_2/a_2724_472# vss 0.33241f
C363 phase_inverter_0/FILLER_0_13_2/a_2276_472# vss 0.33241f
C364 phase_inverter_0/FILLER_0_13_2/a_1828_472# vss 0.33241f
C365 phase_inverter_0/FILLER_0_13_2/a_1380_472# vss 0.33241f
C366 phase_inverter_0/FILLER_0_13_2/a_932_472# vss 0.33241f
C367 phase_inverter_0/FILLER_0_13_2/a_484_472# vss 0.33241f
C368 phase_inverter_0/FILLER_0_13_2/a_36_472# vss 0.404746f
C369 phase_inverter_0/FILLER_0_13_2/a_6844_375# vss 0.233068f
C370 phase_inverter_0/FILLER_0_13_2/a_6396_375# vss 0.171644f
C371 phase_inverter_0/FILLER_0_13_2/a_5948_375# vss 0.171644f
C372 phase_inverter_0/FILLER_0_13_2/a_5500_375# vss 0.171644f
C373 phase_inverter_0/FILLER_0_13_2/a_5052_375# vss 0.171644f
C374 phase_inverter_0/FILLER_0_13_2/a_4604_375# vss 0.171644f
C375 phase_inverter_0/FILLER_0_13_2/a_4156_375# vss 0.171644f
C376 phase_inverter_0/FILLER_0_13_2/a_3708_375# vss 0.171644f
C377 phase_inverter_0/FILLER_0_13_2/a_3260_375# vss 0.171644f
C378 phase_inverter_0/FILLER_0_13_2/a_2812_375# vss 0.171644f
C379 phase_inverter_0/FILLER_0_13_2/a_2364_375# vss 0.171644f
C380 phase_inverter_0/FILLER_0_13_2/a_1916_375# vss 0.171644f
C381 phase_inverter_0/FILLER_0_13_2/a_1468_375# vss 0.171644f
C382 phase_inverter_0/FILLER_0_13_2/a_1020_375# vss 0.171644f
C383 phase_inverter_0/FILLER_0_13_2/a_572_375# vss 0.171644f
C384 phase_inverter_0/FILLER_0_13_2/a_124_375# vss 0.185708f
C385 phase_inverter_0/FILLER_0_0_12/a_1380_472# vss 0.345058f
C386 phase_inverter_0/FILLER_0_0_12/a_932_472# vss 0.33241f
C387 phase_inverter_0/FILLER_0_0_12/a_484_472# vss 0.33241f
C388 phase_inverter_0/FILLER_0_0_12/a_36_472# vss 0.404746f
C389 phase_inverter_0/FILLER_0_0_12/a_1468_375# vss 0.233029f
C390 phase_inverter_0/FILLER_0_0_12/a_1020_375# vss 0.171606f
C391 phase_inverter_0/FILLER_0_0_12/a_572_375# vss 0.171606f
C392 phase_inverter_0/FILLER_0_0_12/a_124_375# vss 0.185399f
C393 phase_inverter_0/FILLER_0_3_44/a_1380_472# vss 0.345058f
C394 phase_inverter_0/FILLER_0_3_44/a_932_472# vss 0.33241f
C395 phase_inverter_0/FILLER_0_3_44/a_484_472# vss 0.33241f
C396 phase_inverter_0/FILLER_0_3_44/a_36_472# vss 0.404746f
C397 phase_inverter_0/FILLER_0_3_44/a_1468_375# vss 0.233029f
C398 phase_inverter_0/FILLER_0_3_44/a_1020_375# vss 0.171606f
C399 phase_inverter_0/FILLER_0_3_44/a_572_375# vss 0.171606f
C400 phase_inverter_0/FILLER_0_3_44/a_124_375# vss 0.185399f
C401 phase_inverter_0/_12_/Z vss 1.135084f
C402 phase_inverter_0/_12_/a_36_113# vss 0.418095f
C403 phase_inverter_0/FILLER_0_15_56/a_484_472# vss 0.345058f
C404 phase_inverter_0/FILLER_0_15_56/a_36_472# vss 0.404746f
C405 phase_inverter_0/FILLER_0_15_56/a_572_375# vss 0.232991f
C406 phase_inverter_0/FILLER_0_15_56/a_124_375# vss 0.185089f
C407 phase_inverter_0/_13_/Z vss 1.131177f
C408 phase_inverter_0/_13_/a_36_113# vss 0.418095f
C409 phase_inverter_0/FILLER_0_2_101/a_36_472# vss 0.417394f
C410 phase_inverter_0/FILLER_0_2_101/a_124_375# vss 0.246306f
C411 phase_inverter_0/FILLER_0_12_12/a_1380_472# vss 0.345058f
C412 phase_inverter_0/FILLER_0_12_12/a_932_472# vss 0.33241f
C413 phase_inverter_0/FILLER_0_12_12/a_484_472# vss 0.33241f
C414 phase_inverter_0/FILLER_0_12_12/a_36_472# vss 0.404746f
C415 phase_inverter_0/FILLER_0_12_12/a_1468_375# vss 0.233029f
C416 phase_inverter_0/FILLER_0_12_12/a_1020_375# vss 0.171606f
C417 phase_inverter_0/FILLER_0_12_12/a_572_375# vss 0.171606f
C418 phase_inverter_0/FILLER_0_12_12/a_124_375# vss 0.185399f
C419 input_signal[8] vss 1.074195f
C420 phase_inverter_0/_14_/Z vss 1.171827f
C421 phase_inverter_0/_14_/a_36_113# vss 0.418095f
C422 phase_inverter_0/FILLER_0_4_2/a_3172_472# vss 0.345058f
C423 phase_inverter_0/FILLER_0_4_2/a_2724_472# vss 0.33241f
C424 phase_inverter_0/FILLER_0_4_2/a_2276_472# vss 0.33241f
C425 phase_inverter_0/FILLER_0_4_2/a_1828_472# vss 0.33241f
C426 phase_inverter_0/FILLER_0_4_2/a_1380_472# vss 0.33241f
C427 phase_inverter_0/FILLER_0_4_2/a_932_472# vss 0.33241f
C428 phase_inverter_0/FILLER_0_4_2/a_484_472# vss 0.33241f
C429 phase_inverter_0/FILLER_0_4_2/a_36_472# vss 0.404746f
C430 phase_inverter_0/FILLER_0_4_2/a_3260_375# vss 0.233093f
C431 phase_inverter_0/FILLER_0_4_2/a_2812_375# vss 0.17167f
C432 phase_inverter_0/FILLER_0_4_2/a_2364_375# vss 0.17167f
C433 phase_inverter_0/FILLER_0_4_2/a_1916_375# vss 0.17167f
C434 phase_inverter_0/FILLER_0_4_2/a_1468_375# vss 0.17167f
C435 phase_inverter_0/FILLER_0_4_2/a_1020_375# vss 0.17167f
C436 phase_inverter_0/FILLER_0_4_2/a_572_375# vss 0.17167f
C437 phase_inverter_0/FILLER_0_4_2/a_124_375# vss 0.185915f
C438 phase_inverter_0/FILLER_0_15_2/a_36_472# vss 0.417394f
C439 phase_inverter_0/FILLER_0_15_2/a_124_375# vss 0.246306f
C440 phase_inverter_0/_15_/Z vss 1.167741f
C441 phase_inverter_0/_15_/a_36_113# vss 0.418095f
C442 phase_inverter_0/FILLER_0_6_107/a_36_472# vss 0.417394f
C443 phase_inverter_0/FILLER_0_6_107/a_124_375# vss 0.246306f
C444 phase_inverter_0/FILLER_0_9_104/a_484_472# vss 0.345058f
C445 phase_inverter_0/FILLER_0_9_104/a_36_472# vss 0.404746f
C446 phase_inverter_0/FILLER_0_9_104/a_572_375# vss 0.232991f
C447 phase_inverter_0/FILLER_0_9_104/a_124_375# vss 0.185089f
C448 phase_inverter_0/FILLER_0_9_72/a_3172_472# vss 0.345058f
C449 phase_inverter_0/FILLER_0_9_72/a_2724_472# vss 0.33241f
C450 phase_inverter_0/FILLER_0_9_72/a_2276_472# vss 0.33241f
C451 phase_inverter_0/FILLER_0_9_72/a_1828_472# vss 0.33241f
C452 phase_inverter_0/FILLER_0_9_72/a_1380_472# vss 0.33241f
C453 phase_inverter_0/FILLER_0_9_72/a_932_472# vss 0.33241f
C454 phase_inverter_0/FILLER_0_9_72/a_484_472# vss 0.33241f
C455 phase_inverter_0/FILLER_0_9_72/a_36_472# vss 0.404746f
C456 phase_inverter_0/FILLER_0_9_72/a_3260_375# vss 0.233093f
C457 phase_inverter_0/FILLER_0_9_72/a_2812_375# vss 0.17167f
C458 phase_inverter_0/FILLER_0_9_72/a_2364_375# vss 0.17167f
C459 phase_inverter_0/FILLER_0_9_72/a_1916_375# vss 0.17167f
C460 phase_inverter_0/FILLER_0_9_72/a_1468_375# vss 0.17167f
C461 phase_inverter_0/FILLER_0_9_72/a_1020_375# vss 0.17167f
C462 phase_inverter_0/FILLER_0_9_72/a_572_375# vss 0.17167f
C463 phase_inverter_0/FILLER_0_9_72/a_124_375# vss 0.185915f
C464 phase_inverter_0/FILLER_0_15_64/a_36_472# vss 0.417394f
C465 phase_inverter_0/FILLER_0_15_64/a_124_375# vss 0.246306f
C466 phase_inverter_0/_16_/Z vss 1.160526f
C467 phase_inverter_0/_16_/a_36_113# vss 0.418095f
C468 phase_inverter_0/FILLER_0_10_101/a_36_472# vss 0.417394f
C469 phase_inverter_0/FILLER_0_10_101/a_124_375# vss 0.246306f
C470 phase_inverter_0/FILLER_0_3_72/a_3172_472# vss 0.345058f
C471 phase_inverter_0/FILLER_0_3_72/a_2724_472# vss 0.33241f
C472 phase_inverter_0/FILLER_0_3_72/a_2276_472# vss 0.33241f
C473 phase_inverter_0/FILLER_0_3_72/a_1828_472# vss 0.33241f
C474 phase_inverter_0/FILLER_0_3_72/a_1380_472# vss 0.33241f
C475 phase_inverter_0/FILLER_0_3_72/a_932_472# vss 0.33241f
C476 phase_inverter_0/FILLER_0_3_72/a_484_472# vss 0.33241f
C477 phase_inverter_0/FILLER_0_3_72/a_36_472# vss 0.404746f
C478 phase_inverter_0/FILLER_0_3_72/a_3260_375# vss 0.233093f
C479 phase_inverter_0/FILLER_0_3_72/a_2812_375# vss 0.17167f
C480 phase_inverter_0/FILLER_0_3_72/a_2364_375# vss 0.17167f
C481 phase_inverter_0/FILLER_0_3_72/a_1916_375# vss 0.17167f
C482 phase_inverter_0/FILLER_0_3_72/a_1468_375# vss 0.17167f
C483 phase_inverter_0/FILLER_0_3_72/a_1020_375# vss 0.17167f
C484 phase_inverter_0/FILLER_0_3_72/a_572_375# vss 0.17167f
C485 phase_inverter_0/FILLER_0_3_72/a_124_375# vss 0.185915f
C486 phase_inverter_0/FILLER_0_8_28/a_36_472# vss 0.417394f
C487 phase_inverter_0/FILLER_0_8_28/a_124_375# vss 0.246306f
C488 phase_inverter_0/_17_/a_36_113# vss 0.418095f
C489 phase_inverter_0/FILLER_0_6_2/a_3172_472# vss 0.345058f
C490 phase_inverter_0/FILLER_0_6_2/a_2724_472# vss 0.33241f
C491 phase_inverter_0/FILLER_0_6_2/a_2276_472# vss 0.33241f
C492 phase_inverter_0/FILLER_0_6_2/a_1828_472# vss 0.33241f
C493 phase_inverter_0/FILLER_0_6_2/a_1380_472# vss 0.33241f
C494 phase_inverter_0/FILLER_0_6_2/a_932_472# vss 0.33241f
C495 phase_inverter_0/FILLER_0_6_2/a_484_472# vss 0.33241f
C496 phase_inverter_0/FILLER_0_6_2/a_36_472# vss 0.404746f
C497 phase_inverter_0/FILLER_0_6_2/a_3260_375# vss 0.233093f
C498 phase_inverter_0/FILLER_0_6_2/a_2812_375# vss 0.17167f
C499 phase_inverter_0/FILLER_0_6_2/a_2364_375# vss 0.17167f
C500 phase_inverter_0/FILLER_0_6_2/a_1916_375# vss 0.17167f
C501 phase_inverter_0/FILLER_0_6_2/a_1468_375# vss 0.17167f
C502 phase_inverter_0/FILLER_0_6_2/a_1020_375# vss 0.17167f
C503 phase_inverter_0/FILLER_0_6_2/a_572_375# vss 0.17167f
C504 phase_inverter_0/FILLER_0_6_2/a_124_375# vss 0.185915f
C505 phase_inverter_0/FILLER_0_15_40/a_1380_472# vss 0.345058f
C506 phase_inverter_0/FILLER_0_15_40/a_932_472# vss 0.33241f
C507 phase_inverter_0/FILLER_0_15_40/a_484_472# vss 0.33241f
C508 phase_inverter_0/FILLER_0_15_40/a_36_472# vss 0.404746f
C509 phase_inverter_0/FILLER_0_15_40/a_1468_375# vss 0.233029f
C510 phase_inverter_0/FILLER_0_15_40/a_1020_375# vss 0.171606f
C511 phase_inverter_0/FILLER_0_15_40/a_572_375# vss 0.171606f
C512 phase_inverter_0/FILLER_0_15_40/a_124_375# vss 0.185399f
C513 phase_inverter_0/_18_/a_36_113# vss 0.418095f
C514 phase_inverter_0/FILLER_0_3_60/a_484_472# vss 0.345058f
C515 phase_inverter_0/FILLER_0_3_60/a_36_472# vss 0.404746f
C516 phase_inverter_0/FILLER_0_3_60/a_572_375# vss 0.232991f
C517 phase_inverter_0/FILLER_0_3_60/a_124_375# vss 0.185089f
C518 phase_inverter_0/FILLER_0_14_107/a_484_472# vss 0.345058f
C519 phase_inverter_0/FILLER_0_14_107/a_36_472# vss 0.404746f
C520 phase_inverter_0/FILLER_0_14_107/a_572_375# vss 0.232991f
C521 phase_inverter_0/FILLER_0_14_107/a_124_375# vss 0.185089f
C522 phase_inverter_0/FILLER_0_15_72/a_1380_472# vss 0.345058f
C523 phase_inverter_0/FILLER_0_15_72/a_932_472# vss 0.33241f
C524 phase_inverter_0/FILLER_0_15_72/a_484_472# vss 0.333066f
C525 phase_inverter_0/FILLER_0_15_72/a_36_472# vss 0.404746f
C526 phase_inverter_0/FILLER_0_15_72/a_1468_375# vss 0.233029f
C527 phase_inverter_0/FILLER_0_15_72/a_1020_375# vss 0.171606f
C528 phase_inverter_0/FILLER_0_15_72/a_572_375# vss 0.171606f
C529 phase_inverter_0/FILLER_0_15_72/a_124_375# vss 0.185399f
C530 phase_inverter_0/_14_/I vss 1.424187f
C531 phase_inverter_0/FILLER_0_8_37/a_6756_472# vss 0.345058f
C532 phase_inverter_0/FILLER_0_8_37/a_6308_472# vss 0.33241f
C533 phase_inverter_0/FILLER_0_8_37/a_5860_472# vss 0.33241f
C534 phase_inverter_0/FILLER_0_8_37/a_5412_472# vss 0.33241f
C535 phase_inverter_0/FILLER_0_8_37/a_4964_472# vss 0.33241f
C536 phase_inverter_0/FILLER_0_8_37/a_4516_472# vss 0.33241f
C537 phase_inverter_0/FILLER_0_8_37/a_4068_472# vss 0.33241f
C538 phase_inverter_0/FILLER_0_8_37/a_3620_472# vss 0.33241f
C539 phase_inverter_0/FILLER_0_8_37/a_3172_472# vss 0.33241f
C540 phase_inverter_0/FILLER_0_8_37/a_2724_472# vss 0.33241f
C541 phase_inverter_0/FILLER_0_8_37/a_2276_472# vss 0.33241f
C542 phase_inverter_0/FILLER_0_8_37/a_1828_472# vss 0.33241f
C543 phase_inverter_0/FILLER_0_8_37/a_1380_472# vss 0.33241f
C544 phase_inverter_0/FILLER_0_8_37/a_932_472# vss 0.33241f
C545 phase_inverter_0/FILLER_0_8_37/a_484_472# vss 0.33241f
C546 phase_inverter_0/FILLER_0_8_37/a_36_472# vss 0.404746f
C547 phase_inverter_0/FILLER_0_8_37/a_6844_375# vss 0.233068f
C548 phase_inverter_0/FILLER_0_8_37/a_6396_375# vss 0.171644f
C549 phase_inverter_0/FILLER_0_8_37/a_5948_375# vss 0.171644f
C550 phase_inverter_0/FILLER_0_8_37/a_5500_375# vss 0.171644f
C551 phase_inverter_0/FILLER_0_8_37/a_5052_375# vss 0.171644f
C552 phase_inverter_0/FILLER_0_8_37/a_4604_375# vss 0.171644f
C553 phase_inverter_0/FILLER_0_8_37/a_4156_375# vss 0.171644f
C554 phase_inverter_0/FILLER_0_8_37/a_3708_375# vss 0.171644f
C555 phase_inverter_0/FILLER_0_8_37/a_3260_375# vss 0.171644f
C556 phase_inverter_0/FILLER_0_8_37/a_2812_375# vss 0.171644f
C557 phase_inverter_0/FILLER_0_8_37/a_2364_375# vss 0.171644f
C558 phase_inverter_0/FILLER_0_8_37/a_1916_375# vss 0.171644f
C559 phase_inverter_0/FILLER_0_8_37/a_1468_375# vss 0.171644f
C560 phase_inverter_0/FILLER_0_8_37/a_1020_375# vss 0.171644f
C561 phase_inverter_0/FILLER_0_8_37/a_572_375# vss 0.171644f
C562 phase_inverter_0/FILLER_0_8_37/a_124_375# vss 0.185708f
C563 phase_inverter_0/_19_/a_36_113# vss 0.418095f
C564 phase_inverter_0/FILLER_0_0_70/a_36_472# vss 0.417394f
C565 phase_inverter_0/FILLER_0_0_70/a_124_375# vss 0.246306f
C566 phase_inverter_0/FILLER_0_14_28/a_36_472# vss 0.417394f
C567 phase_inverter_0/FILLER_0_14_28/a_124_375# vss 0.246306f
C568 phase_inverter_0/FILLER_0_2_37/a_6756_472# vss 0.345058f
C569 phase_inverter_0/FILLER_0_2_37/a_6308_472# vss 0.33241f
C570 phase_inverter_0/FILLER_0_2_37/a_5860_472# vss 0.33241f
C571 phase_inverter_0/FILLER_0_2_37/a_5412_472# vss 0.33241f
C572 phase_inverter_0/FILLER_0_2_37/a_4964_472# vss 0.33241f
C573 phase_inverter_0/FILLER_0_2_37/a_4516_472# vss 0.33241f
C574 phase_inverter_0/FILLER_0_2_37/a_4068_472# vss 0.33241f
C575 phase_inverter_0/FILLER_0_2_37/a_3620_472# vss 0.33241f
C576 phase_inverter_0/FILLER_0_2_37/a_3172_472# vss 0.33241f
C577 phase_inverter_0/FILLER_0_2_37/a_2724_472# vss 0.33241f
C578 phase_inverter_0/FILLER_0_2_37/a_2276_472# vss 0.33241f
C579 phase_inverter_0/FILLER_0_2_37/a_1828_472# vss 0.33241f
C580 phase_inverter_0/FILLER_0_2_37/a_1380_472# vss 0.33241f
C581 phase_inverter_0/FILLER_0_2_37/a_932_472# vss 0.33241f
C582 phase_inverter_0/FILLER_0_2_37/a_484_472# vss 0.33241f
C583 phase_inverter_0/FILLER_0_2_37/a_36_472# vss 0.404746f
C584 phase_inverter_0/FILLER_0_2_37/a_6844_375# vss 0.233068f
C585 phase_inverter_0/FILLER_0_2_37/a_6396_375# vss 0.171644f
C586 phase_inverter_0/FILLER_0_2_37/a_5948_375# vss 0.171644f
C587 phase_inverter_0/FILLER_0_2_37/a_5500_375# vss 0.171644f
C588 phase_inverter_0/FILLER_0_2_37/a_5052_375# vss 0.171644f
C589 phase_inverter_0/FILLER_0_2_37/a_4604_375# vss 0.171644f
C590 phase_inverter_0/FILLER_0_2_37/a_4156_375# vss 0.171644f
C591 phase_inverter_0/FILLER_0_2_37/a_3708_375# vss 0.171644f
C592 phase_inverter_0/FILLER_0_2_37/a_3260_375# vss 0.171644f
C593 phase_inverter_0/FILLER_0_2_37/a_2812_375# vss 0.171644f
C594 phase_inverter_0/FILLER_0_2_37/a_2364_375# vss 0.171644f
C595 phase_inverter_0/FILLER_0_2_37/a_1916_375# vss 0.171644f
C596 phase_inverter_0/FILLER_0_2_37/a_1468_375# vss 0.171644f
C597 phase_inverter_0/FILLER_0_2_37/a_1020_375# vss 0.171644f
C598 phase_inverter_0/FILLER_0_2_37/a_572_375# vss 0.171644f
C599 phase_inverter_0/FILLER_0_2_37/a_124_375# vss 0.185708f
C600 input_signal[9] vss 1.722228f
C601 phase_inverter_0/FILLER_0_3_104/a_484_472# vss 0.345058f
C602 phase_inverter_0/FILLER_0_3_104/a_36_472# vss 0.404746f
C603 phase_inverter_0/FILLER_0_3_104/a_572_375# vss 0.232991f
C604 phase_inverter_0/FILLER_0_3_104/a_124_375# vss 0.185089f
C605 phase_inverter_0/FILLER_0_6_101/a_36_472# vss 0.417394f
C606 phase_inverter_0/FILLER_0_6_101/a_124_375# vss 0.246306f
C607 phase_inverter_0/FILLER_0_14_115/a_36_472# vss 0.417394f
C608 phase_inverter_0/FILLER_0_14_115/a_124_375# vss 0.246306f
C609 phase_inverter_0/input9/a_36_113# vss 0.418095f
C610 phase_inverter_0/FILLER_0_8_12/a_1380_472# vss 0.345058f
C611 phase_inverter_0/FILLER_0_8_12/a_932_472# vss 0.33241f
C612 phase_inverter_0/FILLER_0_8_12/a_484_472# vss 0.33241f
C613 phase_inverter_0/FILLER_0_8_12/a_36_472# vss 0.404746f
C614 phase_inverter_0/FILLER_0_8_12/a_1468_375# vss 0.233029f
C615 phase_inverter_0/FILLER_0_8_12/a_1020_375# vss 0.171606f
C616 phase_inverter_0/FILLER_0_8_12/a_572_375# vss 0.171606f
C617 phase_inverter_0/FILLER_0_8_12/a_124_375# vss 0.185399f
C618 phase_inverter_0/FILLER_0_14_37/a_6756_472# vss 0.345058f
C619 phase_inverter_0/FILLER_0_14_37/a_6308_472# vss 0.33241f
C620 phase_inverter_0/FILLER_0_14_37/a_5860_472# vss 0.33241f
C621 phase_inverter_0/FILLER_0_14_37/a_5412_472# vss 0.33241f
C622 phase_inverter_0/FILLER_0_14_37/a_4964_472# vss 0.33241f
C623 phase_inverter_0/FILLER_0_14_37/a_4516_472# vss 0.33241f
C624 phase_inverter_0/FILLER_0_14_37/a_4068_472# vss 0.33241f
C625 phase_inverter_0/FILLER_0_14_37/a_3620_472# vss 0.33241f
C626 phase_inverter_0/FILLER_0_14_37/a_3172_472# vss 0.33241f
C627 phase_inverter_0/FILLER_0_14_37/a_2724_472# vss 0.33241f
C628 phase_inverter_0/FILLER_0_14_37/a_2276_472# vss 0.33241f
C629 phase_inverter_0/FILLER_0_14_37/a_1828_472# vss 0.33241f
C630 phase_inverter_0/FILLER_0_14_37/a_1380_472# vss 0.33241f
C631 phase_inverter_0/FILLER_0_14_37/a_932_472# vss 0.33241f
C632 phase_inverter_0/FILLER_0_14_37/a_484_472# vss 0.33241f
C633 phase_inverter_0/FILLER_0_14_37/a_36_472# vss 0.404746f
C634 phase_inverter_0/FILLER_0_14_37/a_6844_375# vss 0.233068f
C635 phase_inverter_0/FILLER_0_14_37/a_6396_375# vss 0.171644f
C636 phase_inverter_0/FILLER_0_14_37/a_5948_375# vss 0.171644f
C637 phase_inverter_0/FILLER_0_14_37/a_5500_375# vss 0.171644f
C638 phase_inverter_0/FILLER_0_14_37/a_5052_375# vss 0.171644f
C639 phase_inverter_0/FILLER_0_14_37/a_4604_375# vss 0.171644f
C640 phase_inverter_0/FILLER_0_14_37/a_4156_375# vss 0.171644f
C641 phase_inverter_0/FILLER_0_14_37/a_3708_375# vss 0.171644f
C642 phase_inverter_0/FILLER_0_14_37/a_3260_375# vss 0.171644f
C643 phase_inverter_0/FILLER_0_14_37/a_2812_375# vss 0.171644f
C644 phase_inverter_0/FILLER_0_14_37/a_2364_375# vss 0.171644f
C645 phase_inverter_0/FILLER_0_14_37/a_1916_375# vss 0.171644f
C646 phase_inverter_0/FILLER_0_14_37/a_1468_375# vss 0.171644f
C647 phase_inverter_0/FILLER_0_14_37/a_1020_375# vss 0.171644f
C648 phase_inverter_0/FILLER_0_14_37/a_572_375# vss 0.171644f
C649 phase_inverter_0/FILLER_0_14_37/a_124_375# vss 0.185708f
C650 phase_inverter_0/input8/a_36_113# vss 0.418095f
C651 phase_inverter_0/FILLER_0_5_12/a_3172_472# vss 0.345058f
C652 phase_inverter_0/FILLER_0_5_12/a_2724_472# vss 0.33241f
C653 phase_inverter_0/FILLER_0_5_12/a_2276_472# vss 0.33241f
C654 phase_inverter_0/FILLER_0_5_12/a_1828_472# vss 0.33241f
C655 phase_inverter_0/FILLER_0_5_12/a_1380_472# vss 0.33241f
C656 phase_inverter_0/FILLER_0_5_12/a_932_472# vss 0.33241f
C657 phase_inverter_0/FILLER_0_5_12/a_484_472# vss 0.33241f
C658 phase_inverter_0/FILLER_0_5_12/a_36_472# vss 0.404746f
C659 phase_inverter_0/FILLER_0_5_12/a_3260_375# vss 0.233093f
C660 phase_inverter_0/FILLER_0_5_12/a_2812_375# vss 0.17167f
C661 phase_inverter_0/FILLER_0_5_12/a_2364_375# vss 0.17167f
C662 phase_inverter_0/FILLER_0_5_12/a_1916_375# vss 0.17167f
C663 phase_inverter_0/FILLER_0_5_12/a_1468_375# vss 0.17167f
C664 phase_inverter_0/FILLER_0_5_12/a_1020_375# vss 0.17167f
C665 phase_inverter_0/FILLER_0_5_12/a_572_375# vss 0.17167f
C666 phase_inverter_0/FILLER_0_5_12/a_124_375# vss 0.185915f
C667 phase_inverter_0/input10/a_36_113# vss 0.418095f
C668 phase_inverter_0/FILLER_0_5_44/a_1380_472# vss 0.345058f
C669 phase_inverter_0/FILLER_0_5_44/a_932_472# vss 0.33241f
C670 phase_inverter_0/FILLER_0_5_44/a_484_472# vss 0.33241f
C671 phase_inverter_0/FILLER_0_5_44/a_36_472# vss 0.404746f
C672 phase_inverter_0/FILLER_0_5_44/a_1468_375# vss 0.233029f
C673 phase_inverter_0/FILLER_0_5_44/a_1020_375# vss 0.171606f
C674 phase_inverter_0/FILLER_0_5_44/a_572_375# vss 0.171606f
C675 phase_inverter_0/FILLER_0_5_44/a_124_375# vss 0.185399f
C676 phase_inverter_0/input7/a_36_113# vss 0.418095f
C677 phase_inverter_0/FILLER_0_0_104/a_36_472# vss 0.417394f
C678 phase_inverter_0/FILLER_0_0_104/a_124_375# vss 0.246306f
C679 input_signal[5] vss 1.048828f
C680 phase_inverter_0/input6/a_36_113# vss 0.418095f
C681 phase_inverter_0/FILLER_0_14_101/a_36_472# vss 0.417394f
C682 phase_inverter_0/FILLER_0_14_101/a_124_375# vss 0.246306f
C683 phase_inverter_0/FILLER_0_14_12/a_1380_472# vss 0.345058f
C684 phase_inverter_0/FILLER_0_14_12/a_932_472# vss 0.33241f
C685 phase_inverter_0/FILLER_0_14_12/a_484_472# vss 0.33241f
C686 phase_inverter_0/FILLER_0_14_12/a_36_472# vss 0.404746f
C687 phase_inverter_0/FILLER_0_14_12/a_1468_375# vss 0.233029f
C688 phase_inverter_0/FILLER_0_14_12/a_1020_375# vss 0.171606f
C689 phase_inverter_0/FILLER_0_14_12/a_572_375# vss 0.171606f
C690 phase_inverter_0/FILLER_0_14_12/a_124_375# vss 0.185399f
C691 phase_inverter_0/FILLER_0_11_136/a_36_472# vss 0.417394f
C692 phase_inverter_0/FILLER_0_11_136/a_124_375# vss 0.246306f
C693 phase_inverter_0/input5/a_36_113# vss 0.418095f
C694 phase_inverter_0/_19_/I vss 1.019585f
C695 input_signal[3] vss 0.969415f
C696 phase_inverter_0/input4/a_36_113# vss 0.418095f
C697 phase_inverter_0/FILLER_0_11_66/a_36_472# vss 0.417394f
C698 phase_inverter_0/FILLER_0_11_66/a_124_375# vss 0.246306f
C699 phase_inverter_0/_12_/I vss 1.059653f
C700 phase_inverter_0/input3/a_36_113# vss 0.418095f
C701 phase_inverter_0/_11_/I vss 1.493507f
C702 input_signal[1] vss 1.033314f
C703 phase_inverter_0/input2/a_36_113# vss 0.418095f
C704 phase_inverter_0/FILLER_0_5_72/a_3172_472# vss 0.345058f
C705 phase_inverter_0/FILLER_0_5_72/a_2724_472# vss 0.33241f
C706 phase_inverter_0/FILLER_0_5_72/a_2276_472# vss 0.33241f
C707 phase_inverter_0/FILLER_0_5_72/a_1828_472# vss 0.33241f
C708 phase_inverter_0/FILLER_0_5_72/a_1380_472# vss 0.33241f
C709 phase_inverter_0/FILLER_0_5_72/a_932_472# vss 0.33241f
C710 phase_inverter_0/FILLER_0_5_72/a_484_472# vss 0.33241f
C711 phase_inverter_0/FILLER_0_5_72/a_36_472# vss 0.404746f
C712 phase_inverter_0/FILLER_0_5_72/a_3260_375# vss 0.233093f
C713 phase_inverter_0/FILLER_0_5_72/a_2812_375# vss 0.17167f
C714 phase_inverter_0/FILLER_0_5_72/a_2364_375# vss 0.17167f
C715 phase_inverter_0/FILLER_0_5_72/a_1916_375# vss 0.17167f
C716 phase_inverter_0/FILLER_0_5_72/a_1468_375# vss 0.17167f
C717 phase_inverter_0/FILLER_0_5_72/a_1020_375# vss 0.17167f
C718 phase_inverter_0/FILLER_0_5_72/a_572_375# vss 0.17167f
C719 phase_inverter_0/FILLER_0_5_72/a_124_375# vss 0.185915f
C720 phase_inverter_0/FILLER_0_4_107/a_1380_472# vss 0.345058f
C721 phase_inverter_0/FILLER_0_4_107/a_932_472# vss 0.33241f
C722 phase_inverter_0/FILLER_0_4_107/a_484_472# vss 0.33241f
C723 phase_inverter_0/FILLER_0_4_107/a_36_472# vss 0.404746f
C724 phase_inverter_0/FILLER_0_4_107/a_1468_375# vss 0.233029f
C725 phase_inverter_0/FILLER_0_4_107/a_1020_375# vss 0.171606f
C726 phase_inverter_0/FILLER_0_4_107/a_572_375# vss 0.171606f
C727 phase_inverter_0/FILLER_0_4_107/a_124_375# vss 0.185399f
C728 phase_inverter_0/_10_/I vss 0.979826f
C729 input_signal[0] vss 1.665667f
C730 phase_inverter_0/input1/a_36_113# vss 0.418095f
C731 phase_inverter_0/_03_/ZN vss 1.105776f
C732 phase_inverter_0/FILLER_0_7_104/a_484_472# vss 0.345058f
C733 phase_inverter_0/FILLER_0_7_104/a_36_472# vss 0.404746f
C734 phase_inverter_0/FILLER_0_7_104/a_572_375# vss 0.232991f
C735 phase_inverter_0/FILLER_0_7_104/a_124_375# vss 0.185089f
C736 phase_inverter_0/FILLER_0_5_60/a_484_472# vss 0.345058f
C737 phase_inverter_0/FILLER_0_5_60/a_36_472# vss 0.404746f
C738 phase_inverter_0/FILLER_0_5_60/a_572_375# vss 0.232991f
C739 phase_inverter_0/FILLER_0_5_60/a_124_375# vss 0.185089f
C740 phase_inverter_0/FILLER_0_0_142/a_484_472# vss 0.345058f
C741 phase_inverter_0/FILLER_0_0_142/a_36_472# vss 0.404746f
C742 phase_inverter_0/FILLER_0_0_142/a_572_375# vss 0.232991f
C743 phase_inverter_0/FILLER_0_0_142/a_124_375# vss 0.185089f
C744 phase_inverter_0/_04_/ZN vss 1.111802f
C745 input_signal[7] vss 0.974241f
C746 phase_inverter_0/FILLER_0_16_18/a_1380_472# vss 0.345058f
C747 phase_inverter_0/FILLER_0_16_18/a_932_472# vss 0.33241f
C748 phase_inverter_0/FILLER_0_16_18/a_484_472# vss 0.33241f
C749 phase_inverter_0/FILLER_0_16_18/a_36_472# vss 0.404746f
C750 phase_inverter_0/FILLER_0_16_18/a_1468_375# vss 0.233029f
C751 phase_inverter_0/FILLER_0_16_18/a_1020_375# vss 0.171606f
C752 phase_inverter_0/FILLER_0_16_18/a_572_375# vss 0.171606f
C753 phase_inverter_0/FILLER_0_16_18/a_124_375# vss 0.185399f
C754 phase_inverter_0/net15 vss 1.058175f
C755 phase_inverter_0/_09_/ZN vss 1.363364f
C756 phase_inverter_0/output19/a_224_472# vss 2.38465f
C757 phase_inverter_0/_13_/I vss 1.115417f
C758 phase_inverter_0/FILLER_0_11_72/a_6756_472# vss 0.345058f
C759 phase_inverter_0/FILLER_0_11_72/a_6308_472# vss 0.33241f
C760 phase_inverter_0/FILLER_0_11_72/a_5860_472# vss 0.33241f
C761 phase_inverter_0/FILLER_0_11_72/a_5412_472# vss 0.33241f
C762 phase_inverter_0/FILLER_0_11_72/a_4964_472# vss 0.33241f
C763 phase_inverter_0/FILLER_0_11_72/a_4516_472# vss 0.33241f
C764 phase_inverter_0/FILLER_0_11_72/a_4068_472# vss 0.33241f
C765 phase_inverter_0/FILLER_0_11_72/a_3620_472# vss 0.33241f
C766 phase_inverter_0/FILLER_0_11_72/a_3172_472# vss 0.33241f
C767 phase_inverter_0/FILLER_0_11_72/a_2724_472# vss 0.33241f
C768 phase_inverter_0/FILLER_0_11_72/a_2276_472# vss 0.33241f
C769 phase_inverter_0/FILLER_0_11_72/a_1828_472# vss 0.33241f
C770 phase_inverter_0/FILLER_0_11_72/a_1380_472# vss 0.33241f
C771 phase_inverter_0/FILLER_0_11_72/a_932_472# vss 0.33241f
C772 phase_inverter_0/FILLER_0_11_72/a_484_472# vss 0.33241f
C773 phase_inverter_0/FILLER_0_11_72/a_36_472# vss 0.404746f
C774 phase_inverter_0/FILLER_0_11_72/a_6844_375# vss 0.233068f
C775 phase_inverter_0/FILLER_0_11_72/a_6396_375# vss 0.171644f
C776 phase_inverter_0/FILLER_0_11_72/a_5948_375# vss 0.171644f
C777 phase_inverter_0/FILLER_0_11_72/a_5500_375# vss 0.171644f
C778 phase_inverter_0/FILLER_0_11_72/a_5052_375# vss 0.171644f
C779 phase_inverter_0/FILLER_0_11_72/a_4604_375# vss 0.171644f
C780 phase_inverter_0/FILLER_0_11_72/a_4156_375# vss 0.171644f
C781 phase_inverter_0/FILLER_0_11_72/a_3708_375# vss 0.171644f
C782 phase_inverter_0/FILLER_0_11_72/a_3260_375# vss 0.171644f
C783 phase_inverter_0/FILLER_0_11_72/a_2812_375# vss 0.171644f
C784 phase_inverter_0/FILLER_0_11_72/a_2364_375# vss 0.171644f
C785 phase_inverter_0/FILLER_0_11_72/a_1916_375# vss 0.171644f
C786 phase_inverter_0/FILLER_0_11_72/a_1468_375# vss 0.171644f
C787 phase_inverter_0/FILLER_0_11_72/a_1020_375# vss 0.171644f
C788 phase_inverter_0/FILLER_0_11_72/a_572_375# vss 0.171644f
C789 phase_inverter_0/FILLER_0_11_72/a_124_375# vss 0.185708f
C790 phase_inverter_0/FILLER_0_4_37/a_6756_472# vss 0.345058f
C791 phase_inverter_0/FILLER_0_4_37/a_6308_472# vss 0.33241f
C792 phase_inverter_0/FILLER_0_4_37/a_5860_472# vss 0.33241f
C793 phase_inverter_0/FILLER_0_4_37/a_5412_472# vss 0.33241f
C794 phase_inverter_0/FILLER_0_4_37/a_4964_472# vss 0.33241f
C795 phase_inverter_0/FILLER_0_4_37/a_4516_472# vss 0.33241f
C796 phase_inverter_0/FILLER_0_4_37/a_4068_472# vss 0.33241f
C797 phase_inverter_0/FILLER_0_4_37/a_3620_472# vss 0.33241f
C798 phase_inverter_0/FILLER_0_4_37/a_3172_472# vss 0.33241f
C799 phase_inverter_0/FILLER_0_4_37/a_2724_472# vss 0.33241f
C800 phase_inverter_0/FILLER_0_4_37/a_2276_472# vss 0.33241f
C801 phase_inverter_0/FILLER_0_4_37/a_1828_472# vss 0.33241f
C802 phase_inverter_0/FILLER_0_4_37/a_1380_472# vss 0.33241f
C803 phase_inverter_0/FILLER_0_4_37/a_932_472# vss 0.33241f
C804 phase_inverter_0/FILLER_0_4_37/a_484_472# vss 0.33241f
C805 phase_inverter_0/FILLER_0_4_37/a_36_472# vss 0.404746f
C806 phase_inverter_0/FILLER_0_4_37/a_6844_375# vss 0.233068f
C807 phase_inverter_0/FILLER_0_4_37/a_6396_375# vss 0.171644f
C808 phase_inverter_0/FILLER_0_4_37/a_5948_375# vss 0.171644f
C809 phase_inverter_0/FILLER_0_4_37/a_5500_375# vss 0.171644f
C810 phase_inverter_0/FILLER_0_4_37/a_5052_375# vss 0.171644f
C811 phase_inverter_0/FILLER_0_4_37/a_4604_375# vss 0.171644f
C812 phase_inverter_0/FILLER_0_4_37/a_4156_375# vss 0.171644f
C813 phase_inverter_0/FILLER_0_4_37/a_3708_375# vss 0.171644f
C814 phase_inverter_0/FILLER_0_4_37/a_3260_375# vss 0.171644f
C815 phase_inverter_0/FILLER_0_4_37/a_2812_375# vss 0.171644f
C816 phase_inverter_0/FILLER_0_4_37/a_2364_375# vss 0.171644f
C817 phase_inverter_0/FILLER_0_4_37/a_1916_375# vss 0.171644f
C818 phase_inverter_0/FILLER_0_4_37/a_1468_375# vss 0.171644f
C819 phase_inverter_0/FILLER_0_4_37/a_1020_375# vss 0.171644f
C820 phase_inverter_0/FILLER_0_4_37/a_572_375# vss 0.171644f
C821 phase_inverter_0/FILLER_0_4_37/a_124_375# vss 0.185708f
C822 phase_inverter_0/_08_/ZN vss 1.295594f
C823 phase_inverter_0/output18/a_224_472# vss 2.39122f
C824 phase_inverter_0/_15_/I vss 1.113137f
C825 phase_inverter_0/_18_/Z vss 1.167483f
C826 phase_inverter_0/output29/a_224_472# vss 2.38465f
C827 phase_inverter_0/FILLER_0_12_107/a_1380_472# vss 0.345058f
C828 phase_inverter_0/FILLER_0_12_107/a_932_472# vss 0.33241f
C829 phase_inverter_0/FILLER_0_12_107/a_484_472# vss 0.33241f
C830 phase_inverter_0/FILLER_0_12_107/a_36_472# vss 0.404746f
C831 phase_inverter_0/FILLER_0_12_107/a_1468_375# vss 0.233029f
C832 phase_inverter_0/FILLER_0_12_107/a_1020_375# vss 0.171606f
C833 phase_inverter_0/FILLER_0_12_107/a_572_375# vss 0.171606f
C834 phase_inverter_0/FILLER_0_12_107/a_124_375# vss 0.185399f
C835 phase_inverter_0/FILLER_0_10_28/a_36_472# vss 0.417394f
C836 phase_inverter_0/FILLER_0_10_28/a_124_375# vss 0.246306f
C837 phase_inverter_0/_07_/ZN vss 1.113234f
C838 phase_inverter_0/output17/a_224_472# vss 2.38465f
C839 phase_inverter_0/_16_/I vss 0.912843f
C840 phase_inverter_0/_17_/Z vss 1.120758f
C841 phase_inverter_0/output28/a_224_472# vss 2.38465f
C842 phase_inverter_0/_06_/ZN vss 1.134591f
C843 phase_inverter_0/output16/a_224_472# vss 2.38465f
C844 phase_inverter_0/output27/a_224_472# vss 2.38465f
C845 phase_inverter_0/_17_/I vss 0.917813f
C846 phase_inverter_0/FILLER_0_16_36/a_3172_472# vss 0.345058f
C847 phase_inverter_0/FILLER_0_16_36/a_2724_472# vss 0.33241f
C848 phase_inverter_0/FILLER_0_16_36/a_2276_472# vss 0.33241f
C849 phase_inverter_0/FILLER_0_16_36/a_1828_472# vss 0.33241f
C850 phase_inverter_0/FILLER_0_16_36/a_1380_472# vss 0.33241f
C851 phase_inverter_0/FILLER_0_16_36/a_932_472# vss 0.33241f
C852 phase_inverter_0/FILLER_0_16_36/a_484_472# vss 0.33241f
C853 phase_inverter_0/FILLER_0_16_36/a_36_472# vss 0.404746f
C854 phase_inverter_0/FILLER_0_16_36/a_3260_375# vss 0.233093f
C855 phase_inverter_0/FILLER_0_16_36/a_2812_375# vss 0.17167f
C856 phase_inverter_0/FILLER_0_16_36/a_2364_375# vss 0.17167f
C857 phase_inverter_0/FILLER_0_16_36/a_1916_375# vss 0.17167f
C858 phase_inverter_0/FILLER_0_16_36/a_1468_375# vss 0.17167f
C859 phase_inverter_0/FILLER_0_16_36/a_1020_375# vss 0.17167f
C860 phase_inverter_0/FILLER_0_16_36/a_572_375# vss 0.17167f
C861 phase_inverter_0/FILLER_0_16_36/a_124_375# vss 0.190644f
C862 phase_inverter_0/FILLER_0_10_37/a_6756_472# vss 0.345058f
C863 phase_inverter_0/FILLER_0_10_37/a_6308_472# vss 0.33241f
C864 phase_inverter_0/FILLER_0_10_37/a_5860_472# vss 0.33241f
C865 phase_inverter_0/FILLER_0_10_37/a_5412_472# vss 0.33241f
C866 phase_inverter_0/FILLER_0_10_37/a_4964_472# vss 0.33241f
C867 phase_inverter_0/FILLER_0_10_37/a_4516_472# vss 0.33241f
C868 phase_inverter_0/FILLER_0_10_37/a_4068_472# vss 0.33241f
C869 phase_inverter_0/FILLER_0_10_37/a_3620_472# vss 0.33241f
C870 phase_inverter_0/FILLER_0_10_37/a_3172_472# vss 0.33241f
C871 phase_inverter_0/FILLER_0_10_37/a_2724_472# vss 0.33241f
C872 phase_inverter_0/FILLER_0_10_37/a_2276_472# vss 0.33241f
C873 phase_inverter_0/FILLER_0_10_37/a_1828_472# vss 0.33241f
C874 phase_inverter_0/FILLER_0_10_37/a_1380_472# vss 0.33241f
C875 phase_inverter_0/FILLER_0_10_37/a_932_472# vss 0.33241f
C876 phase_inverter_0/FILLER_0_10_37/a_484_472# vss 0.33241f
C877 phase_inverter_0/FILLER_0_10_37/a_36_472# vss 0.404746f
C878 phase_inverter_0/FILLER_0_10_37/a_6844_375# vss 0.233068f
C879 phase_inverter_0/FILLER_0_10_37/a_6396_375# vss 0.171644f
C880 phase_inverter_0/FILLER_0_10_37/a_5948_375# vss 0.171644f
C881 phase_inverter_0/FILLER_0_10_37/a_5500_375# vss 0.171644f
C882 phase_inverter_0/FILLER_0_10_37/a_5052_375# vss 0.171644f
C883 phase_inverter_0/FILLER_0_10_37/a_4604_375# vss 0.171644f
C884 phase_inverter_0/FILLER_0_10_37/a_4156_375# vss 0.171644f
C885 phase_inverter_0/FILLER_0_10_37/a_3708_375# vss 0.171644f
C886 phase_inverter_0/FILLER_0_10_37/a_3260_375# vss 0.171644f
C887 phase_inverter_0/FILLER_0_10_37/a_2812_375# vss 0.171644f
C888 phase_inverter_0/FILLER_0_10_37/a_2364_375# vss 0.171644f
C889 phase_inverter_0/FILLER_0_10_37/a_1916_375# vss 0.171644f
C890 phase_inverter_0/FILLER_0_10_37/a_1468_375# vss 0.171644f
C891 phase_inverter_0/FILLER_0_10_37/a_1020_375# vss 0.171644f
C892 phase_inverter_0/FILLER_0_10_37/a_572_375# vss 0.171644f
C893 phase_inverter_0/FILLER_0_10_37/a_124_375# vss 0.185708f
C894 phase_inverter_0/FILLER_0_7_66/a_36_472# vss 0.417394f
C895 phase_inverter_0/FILLER_0_7_66/a_124_375# vss 0.246306f
C896 phase_inverter_0/FILLER_0_4_101/a_36_472# vss 0.417394f
C897 phase_inverter_0/FILLER_0_4_101/a_124_375# vss 0.246306f
C898 phase_inverter_0/output15/a_224_472# vss 2.38465f
C899 phase_inverter_0/_18_/I vss 0.865773f
C900 phase_inverter_0/output26/a_224_472# vss 2.38465f
C901 phase_inverter_0/FILLER_0_1_12/a_3172_472# vss 0.345058f
C902 phase_inverter_0/FILLER_0_1_12/a_2724_472# vss 0.33241f
C903 phase_inverter_0/FILLER_0_1_12/a_2276_472# vss 0.33241f
C904 phase_inverter_0/FILLER_0_1_12/a_1828_472# vss 0.33241f
C905 phase_inverter_0/FILLER_0_1_12/a_1380_472# vss 0.33241f
C906 phase_inverter_0/FILLER_0_1_12/a_932_472# vss 0.33241f
C907 phase_inverter_0/FILLER_0_1_12/a_484_472# vss 0.33241f
C908 phase_inverter_0/FILLER_0_1_12/a_36_472# vss 0.404746f
C909 phase_inverter_0/FILLER_0_1_12/a_3260_375# vss 0.233093f
C910 phase_inverter_0/FILLER_0_1_12/a_2812_375# vss 0.17167f
C911 phase_inverter_0/FILLER_0_1_12/a_2364_375# vss 0.17167f
C912 phase_inverter_0/FILLER_0_1_12/a_1916_375# vss 0.17167f
C913 phase_inverter_0/FILLER_0_1_12/a_1468_375# vss 0.17167f
C914 phase_inverter_0/FILLER_0_1_12/a_1020_375# vss 0.17167f
C915 phase_inverter_0/FILLER_0_1_12/a_572_375# vss 0.17167f
C916 phase_inverter_0/FILLER_0_1_12/a_124_375# vss 0.185915f
C917 phase_inverter_0/output14/a_224_472# vss 2.38465f
C918 phase_inverter_0/output25/a_224_472# vss 2.38465f
C919 phase_inverter_0/FILLER_0_1_44/a_1380_472# vss 0.345058f
C920 phase_inverter_0/FILLER_0_1_44/a_932_472# vss 0.33241f
C921 phase_inverter_0/FILLER_0_1_44/a_484_472# vss 0.33241f
C922 phase_inverter_0/FILLER_0_1_44/a_36_472# vss 0.404746f
C923 phase_inverter_0/FILLER_0_1_44/a_1468_375# vss 0.233029f
C924 phase_inverter_0/FILLER_0_1_44/a_1020_375# vss 0.171606f
C925 phase_inverter_0/FILLER_0_1_44/a_572_375# vss 0.171606f
C926 phase_inverter_0/FILLER_0_1_44/a_124_375# vss 0.185399f
C927 phase_inverter_0/FILLER_0_7_2/a_6756_472# vss 0.345058f
C928 phase_inverter_0/FILLER_0_7_2/a_6308_472# vss 0.33241f
C929 phase_inverter_0/FILLER_0_7_2/a_5860_472# vss 0.33241f
C930 phase_inverter_0/FILLER_0_7_2/a_5412_472# vss 0.33241f
C931 phase_inverter_0/FILLER_0_7_2/a_4964_472# vss 0.33241f
C932 phase_inverter_0/FILLER_0_7_2/a_4516_472# vss 0.33241f
C933 phase_inverter_0/FILLER_0_7_2/a_4068_472# vss 0.33241f
C934 phase_inverter_0/FILLER_0_7_2/a_3620_472# vss 0.33241f
C935 phase_inverter_0/FILLER_0_7_2/a_3172_472# vss 0.33241f
C936 phase_inverter_0/FILLER_0_7_2/a_2724_472# vss 0.33241f
C937 phase_inverter_0/FILLER_0_7_2/a_2276_472# vss 0.33241f
C938 phase_inverter_0/FILLER_0_7_2/a_1828_472# vss 0.33241f
C939 phase_inverter_0/FILLER_0_7_2/a_1380_472# vss 0.33241f
C940 phase_inverter_0/FILLER_0_7_2/a_932_472# vss 0.33241f
C941 phase_inverter_0/FILLER_0_7_2/a_484_472# vss 0.33241f
C942 phase_inverter_0/FILLER_0_7_2/a_36_472# vss 0.404746f
C943 phase_inverter_0/FILLER_0_7_2/a_6844_375# vss 0.233068f
C944 phase_inverter_0/FILLER_0_7_2/a_6396_375# vss 0.171644f
C945 phase_inverter_0/FILLER_0_7_2/a_5948_375# vss 0.171644f
C946 phase_inverter_0/FILLER_0_7_2/a_5500_375# vss 0.171644f
C947 phase_inverter_0/FILLER_0_7_2/a_5052_375# vss 0.171644f
C948 phase_inverter_0/FILLER_0_7_2/a_4604_375# vss 0.171644f
C949 phase_inverter_0/FILLER_0_7_2/a_4156_375# vss 0.171644f
C950 phase_inverter_0/FILLER_0_7_2/a_3708_375# vss 0.171644f
C951 phase_inverter_0/FILLER_0_7_2/a_3260_375# vss 0.171644f
C952 phase_inverter_0/FILLER_0_7_2/a_2812_375# vss 0.171644f
C953 phase_inverter_0/FILLER_0_7_2/a_2364_375# vss 0.171644f
C954 phase_inverter_0/FILLER_0_7_2/a_1916_375# vss 0.171644f
C955 phase_inverter_0/FILLER_0_7_2/a_1468_375# vss 0.171644f
C956 phase_inverter_0/FILLER_0_7_2/a_1020_375# vss 0.171644f
C957 phase_inverter_0/FILLER_0_7_2/a_572_375# vss 0.171644f
C958 phase_inverter_0/FILLER_0_7_2/a_124_375# vss 0.185708f
C959 phase_inverter_0/output13/a_224_472# vss 2.38465f
C960 phase_inverter_0/FILLER_0_8_107/a_484_472# vss 0.345058f
C961 phase_inverter_0/FILLER_0_8_107/a_36_472# vss 0.404746f
C962 phase_inverter_0/FILLER_0_8_107/a_572_375# vss 0.232991f
C963 phase_inverter_0/FILLER_0_8_107/a_124_375# vss 0.185089f
C964 phase_inverter_0/output24/a_224_472# vss 2.38465f
C965 phase_inverter_0/FILLER_0_10_12/a_1380_472# vss 0.345058f
C966 phase_inverter_0/FILLER_0_10_12/a_932_472# vss 0.33241f
C967 phase_inverter_0/FILLER_0_10_12/a_484_472# vss 0.33241f
C968 phase_inverter_0/FILLER_0_10_12/a_36_472# vss 0.404746f
C969 phase_inverter_0/FILLER_0_10_12/a_1468_375# vss 0.233029f
C970 phase_inverter_0/FILLER_0_10_12/a_1020_375# vss 0.171606f
C971 phase_inverter_0/FILLER_0_10_12/a_572_375# vss 0.171606f
C972 phase_inverter_0/FILLER_0_10_12/a_124_375# vss 0.185399f
C973 phase_inverter_0/FILLER_0_13_66/a_36_472# vss 0.417394f
C974 phase_inverter_0/FILLER_0_13_66/a_124_375# vss 0.246306f
C975 phase_inverter_0/_02_/ZN vss 1.077381f
C976 phase_inverter_0/output12/a_224_472# vss 2.38465f
C977 phase_inverter_0/output23/a_224_472# vss 2.38465f
C978 phase_inverter_0/FILLER_0_12_101/a_36_472# vss 0.417394f
C979 phase_inverter_0/FILLER_0_12_101/a_124_375# vss 0.246306f
C980 carray_in_1/n0 vss 19.828964f
C981 phase_inverter_0/_01_/ZN vss 1.235885f
C982 phase_inverter_0/output11/a_224_472# vss 2.38465f
C983 phase_inverter_0/output22/a_224_472# vss 2.38465f
C984 input_signal[2] vss 0.99345f
C985 phase_inverter_0/FILLER_0_7_72/a_3172_472# vss 0.345058f
C986 phase_inverter_0/FILLER_0_7_72/a_2724_472# vss 0.33241f
C987 phase_inverter_0/FILLER_0_7_72/a_2276_472# vss 0.33241f
C988 phase_inverter_0/FILLER_0_7_72/a_1828_472# vss 0.33241f
C989 phase_inverter_0/FILLER_0_7_72/a_1380_472# vss 0.33241f
C990 phase_inverter_0/FILLER_0_7_72/a_932_472# vss 0.33241f
C991 phase_inverter_0/FILLER_0_7_72/a_484_472# vss 0.33241f
C992 phase_inverter_0/FILLER_0_7_72/a_36_472# vss 0.404746f
C993 phase_inverter_0/FILLER_0_7_72/a_3260_375# vss 0.233093f
C994 phase_inverter_0/FILLER_0_7_72/a_2812_375# vss 0.17167f
C995 phase_inverter_0/FILLER_0_7_72/a_2364_375# vss 0.17167f
C996 phase_inverter_0/FILLER_0_7_72/a_1916_375# vss 0.17167f
C997 phase_inverter_0/FILLER_0_7_72/a_1468_375# vss 0.17167f
C998 phase_inverter_0/FILLER_0_7_72/a_1020_375# vss 0.17167f
C999 phase_inverter_0/FILLER_0_7_72/a_572_375# vss 0.17167f
C1000 phase_inverter_0/FILLER_0_7_72/a_124_375# vss 0.185915f
C1001 phase_inverter_0/FILLER_0_9_2/a_6756_472# vss 0.345058f
C1002 phase_inverter_0/FILLER_0_9_2/a_6308_472# vss 0.33241f
C1003 phase_inverter_0/FILLER_0_9_2/a_5860_472# vss 0.33241f
C1004 phase_inverter_0/FILLER_0_9_2/a_5412_472# vss 0.33241f
C1005 phase_inverter_0/FILLER_0_9_2/a_4964_472# vss 0.33241f
C1006 phase_inverter_0/FILLER_0_9_2/a_4516_472# vss 0.33241f
C1007 phase_inverter_0/FILLER_0_9_2/a_4068_472# vss 0.33241f
C1008 phase_inverter_0/FILLER_0_9_2/a_3620_472# vss 0.33241f
C1009 phase_inverter_0/FILLER_0_9_2/a_3172_472# vss 0.33241f
C1010 phase_inverter_0/FILLER_0_9_2/a_2724_472# vss 0.33241f
C1011 phase_inverter_0/FILLER_0_9_2/a_2276_472# vss 0.33241f
C1012 phase_inverter_0/FILLER_0_9_2/a_1828_472# vss 0.33241f
C1013 phase_inverter_0/FILLER_0_9_2/a_1380_472# vss 0.33241f
C1014 phase_inverter_0/FILLER_0_9_2/a_932_472# vss 0.33241f
C1015 phase_inverter_0/FILLER_0_9_2/a_484_472# vss 0.33241f
C1016 phase_inverter_0/FILLER_0_9_2/a_36_472# vss 0.404746f
C1017 phase_inverter_0/FILLER_0_9_2/a_6844_375# vss 0.233068f
C1018 phase_inverter_0/FILLER_0_9_2/a_6396_375# vss 0.171644f
C1019 phase_inverter_0/FILLER_0_9_2/a_5948_375# vss 0.171644f
C1020 phase_inverter_0/FILLER_0_9_2/a_5500_375# vss 0.171644f
C1021 phase_inverter_0/FILLER_0_9_2/a_5052_375# vss 0.171644f
C1022 phase_inverter_0/FILLER_0_9_2/a_4604_375# vss 0.171644f
C1023 phase_inverter_0/FILLER_0_9_2/a_4156_375# vss 0.171644f
C1024 phase_inverter_0/FILLER_0_9_2/a_3708_375# vss 0.171644f
C1025 phase_inverter_0/FILLER_0_9_2/a_3260_375# vss 0.171644f
C1026 phase_inverter_0/FILLER_0_9_2/a_2812_375# vss 0.171644f
C1027 phase_inverter_0/FILLER_0_9_2/a_2364_375# vss 0.171644f
C1028 phase_inverter_0/FILLER_0_9_2/a_1916_375# vss 0.171644f
C1029 phase_inverter_0/FILLER_0_9_2/a_1468_375# vss 0.171644f
C1030 phase_inverter_0/FILLER_0_9_2/a_1020_375# vss 0.171644f
C1031 phase_inverter_0/FILLER_0_9_2/a_572_375# vss 0.171644f
C1032 phase_inverter_0/FILLER_0_9_2/a_124_375# vss 0.185708f
C1033 carray_in_0/n0 vss 18.960093f
C1034 phase_inverter_0/_10_/Z vss 1.18279f
C1035 phase_inverter_0/output21/a_224_472# vss 2.390638f
C1036 phase_inverter_0/_00_/ZN vss 1.56724f
C1037 phase_inverter_0/output20/a_224_472# vss 2.386258f
C1038 phase_inverter_0/FILLER_0_1_72/a_1380_472# vss 0.345058f
C1039 phase_inverter_0/FILLER_0_1_72/a_932_472# vss 0.33241f
C1040 phase_inverter_0/FILLER_0_1_72/a_484_472# vss 0.33241f
C1041 phase_inverter_0/FILLER_0_1_72/a_36_472# vss 0.404746f
C1042 phase_inverter_0/FILLER_0_1_72/a_1468_375# vss 0.233029f
C1043 phase_inverter_0/FILLER_0_1_72/a_1020_375# vss 0.171606f
C1044 phase_inverter_0/FILLER_0_1_72/a_572_375# vss 0.172262f
C1045 phase_inverter_0/FILLER_0_1_72/a_124_375# vss 0.185399f
C1046 carray_in_1/n1 vss 26.054531f
C1047 carray_in_1/n4 vss 40.26557f
C1048 carray_in_1/n5 vss 48.29981f
C1049 carray_in_1/n2 vss 31.908575f
C1050 carray_in_1/n3 vss 34.573807f
C1051 carray_in_1/n9 vss 15.677258f
C1052 inputm vss -0.686844p
C1053 carray_in_1/n8 vss 41.236954f
C1054 carray_in_1/n7 vss 56.976776f
C1055 carray_in_1/n6 vss 53.73989f
C1056 carray_in_0/n1 vss 26.210373f
C1057 carray_in_0/n4 vss 40.29222f
C1058 carray_in_0/n5 vss 48.35306f
C1059 carray_in_0/n2 vss 31.825562f
C1060 carray_in_0/n3 vss 34.694798f
C1061 carray_in_0/n9 vss 15.763344f
C1062 inputp vss -0.686844p
C1063 carray_in_0/n8 vss 41.365013f
C1064 carray_in_0/n7 vss 57.173172f
C1065 carray_in_0/n6 vss 53.727947f
.ends

