* NGSPICE file created from saradc.ext - technology: gf180mcuD

.subckt XM2_latch_x4 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 S G 0.143803f
C2 S D 0.09188f
C3 D VSUBS 0.04225f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.56551f
.ends

.subckt XM1_latch_x4 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.226575f
.ends

.subckt x4_latch vdd out in vss
XXM2_latch_x4_0 in out vdd vss XM2_latch_x4
XXM1_latch_x4_0 in out vss XM1_latch_x4
C0 vdd out 0.102755f
C1 out in 0.057341f
C2 vdd in 0.039699f
C3 out vss 0.49906f
C4 in vss 0.450066f
C5 vdd vss 1.7619f
.ends

.subckt XM2_latch_x3 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 S D 0.09188f
C2 S G 0.143803f
C3 D VSUBS 0.04225f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.56551f
.ends

.subckt XM1_latch_x3 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.226575f
.ends

.subckt x3_latch out in vdd vss
XXM2_latch_x3_0 in out vdd vss XM2_latch_x3
XXM1_latch_x3_0 in out vss XM1_latch_x3
C0 in out 0.057341f
C1 vdd out 0.102755f
C2 vdd in 0.039699f
C3 out vss 0.49906f
C4 in vss 0.450066f
C5 vdd vss 1.761853f
.ends

.subckt XM4_latch G D a_258_n1293# S
X0 S G D S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt XM2_latch_x2 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 S D 0.091354f
C2 S G 0.143685f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.5328f
.ends

.subckt XM1_latch_x2 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt x2_latch vdd out in vss
XXM2_latch_x2_0 in out vdd vss XM2_latch_x2
XXM1_latch_x2_0 in out vss XM1_latch_x2
C0 in out 0.057341f
C1 vdd out 0.088354f
C2 vdd in 0.039609f
C3 out vss 0.511014f
C4 in vss 0.449897f
C5 vdd vss 1.73873f
.ends

.subckt XM3_latch G D a_n349_n1268# S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt XM2_latch_x1 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 S D 0.091354f
C2 S G 0.143685f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.082818f
C5 S VSUBS 1.5328f
.ends

.subckt XM1_latch_x1 G D S a_n254_114#
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134096f
C2 G S 0.22648f
.ends

.subckt x1_latch out in XM1_latch_x1_0/a_n254_114# vdd vss
XXM2_latch_x1_0 in out vdd vss XM2_latch_x1
XXM1_latch_x1_0 in out vss XM1_latch_x1_0/a_n254_114# XM1_latch_x1
C0 in out 0.057341f
C1 vdd out 0.088354f
C2 vdd in 0.039609f
C3 out vss 0.511014f
C4 in vss 0.449897f
C5 vdd vss 1.738608f
.ends

.subckt latch tutyuu1 tutyuu2 Qn Q S R vdd vss
Xx4_latch_0 vdd tutyuu1 S vss x4_latch
Xx3_latch_0 tutyuu2 R vdd vss x3_latch
XXM4_latch_0 tutyuu2 Q vss vss XM4_latch
Xx2_latch_0 vdd Qn Q vss x2_latch
XXM3_latch_0 tutyuu1 Qn vss vss XM3_latch
Xx1_latch_0 Q Qn vss vdd vss x1_latch
C0 tutyuu1 vdd 0.101448f
C1 tutyuu1 S 0.115854f
C2 R Q 0.011346f
C3 Qn Q 1.472762f
C4 R tutyuu2 0.115854f
C5 Qn tutyuu2 0.060761f
C6 R vdd 0.053607f
C7 Q tutyuu2 0.109341f
C8 Qn vdd 0.059024f
C9 Qn S 0.011276f
C10 Q vdd 0.35434f
C11 Qn tutyuu1 0.109231f
C12 tutyuu1 Q 0.060871f
C13 vdd tutyuu2 0.101384f
C14 vdd S 0.053607f
C15 vdd vss 5.959083f
C16 Qn vss 0.913293f
C17 Q vss 0.942836f
C18 tutyuu2 vss 0.702253f
C19 R vss 0.476811f
C20 tutyuu1 vss 0.702189f
C21 S vss 0.476811f
.ends

.subckt XM2_buffer_inv2 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S G 0.138578f
C1 D G 0.001764f
C2 D S 0.090564f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.08816f
C5 S VSUBS 1.2321f
.ends

.subckt XM1_buffer_inv2 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt buffer_inv2 vdd out in vss
XXM2_buffer_inv2_0 in out vdd vss XM2_buffer_inv2
XXM1_buffer_inv2_0 in out vss XM1_buffer_inv2
C0 vdd in 0.034991f
C1 out in 0.057341f
C2 out vdd 0.086562f
C3 out vss 0.51823f
C4 in vss 0.460091f
C5 vdd vss 1.392287f
.ends

.subckt XM1_buffer_inv1 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt buffer_inv1 vdd out in XM2_buffer_inv1_0/w_n90_n162# vss
XXM1_buffer_inv1_0 in out vss XM1_buffer_inv1
C0 XM2_buffer_inv1_0/w_n90_n162# vdd 0.009724f
C1 XM2_buffer_inv1_0/w_n90_n162# in 0.049713f
C2 vdd out 0.142029f
C3 in out 0.058676f
C4 XM2_buffer_inv1_0/w_n90_n162# out 0.007628f
C5 in vdd 0.040357f
C6 out vss 0.548612f
C7 in vss 0.543919f
C8 vdd vss 0.438255f
C9 XM2_buffer_inv1_0/w_n90_n162# vss 0.176185f
.ends

.subckt buffer middle out in vdd vss buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162#
Xbuffer_inv2_0 vdd out middle vss buffer_inv2
Xbuffer_inv1_0 vdd middle in buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vss buffer_inv1
C0 middle buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# 0.003733f
C1 middle out 0.160929f
C2 vdd buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# 0.007171f
C3 in buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# 0.051621f
C4 out vdd 0.039935f
C5 middle vdd 0.190904f
C6 middle in 0.119536f
C7 vdd in 0.054064f
C8 middle vss 0.950535f
C9 in vss 0.600677f
C10 vdd vss 1.632177f
C11 buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vss 0.17473f
C12 out vss 0.56762f
.ends

.subckt inv_p VNW VPW VSS ZN I VDD VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 ZN VSS 0.180794f
C1 VDD VSS 0.029045f
C2 ZN VDD 0.271625f
C3 VNW VSS 0.006277f
C4 VNW ZN 0.023676f
C5 VNW VDD 0.082022f
C6 I VSS 0.091531f
C7 I ZN 0.58604f
C8 I VDD 0.074838f
C9 VNW I 0.285482f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu_p inv_p_7/I inv_p_9/ZN inv_p_6/ZN inv_p_3/ZN inv_p_0/ZN inv_p_0/I
+ inv_p_10/I inv_p_4/I inv_p_8/ZN inv_p_2/ZN inv_p_5/ZN inv_p_6/I inv_p_2/I inv_p_10/ZN
+ inv_p_8/I inv_p_1/I inv_p_9/I inv_p_7/ZN inv_p_4/ZN inv_p_1/ZN inv_p_3/I inv_p_5/I
+ vss vdd
Xinv_p_0 vdd inv_p_0/VPW vss inv_p_0/ZN inv_p_0/I vdd vss inv_p
Xinv_p_1 vdd inv_p_1/VPW vss inv_p_1/ZN inv_p_1/I vdd vss inv_p
Xinv_p_2 vdd inv_p_2/VPW vss inv_p_2/ZN inv_p_2/I vdd vss inv_p
Xinv_p_3 vdd inv_p_3/VPW vss inv_p_3/ZN inv_p_3/I vdd vss inv_p
Xinv_p_4 vdd inv_p_4/VPW vss inv_p_4/ZN inv_p_4/I vdd vss inv_p
Xinv_p_5 vdd inv_p_5/VPW vss inv_p_5/ZN inv_p_5/I vdd vss inv_p
Xinv_p_6 vdd inv_p_6/VPW vss inv_p_6/ZN inv_p_6/I vdd vss inv_p
Xinv_p_7 vdd inv_p_7/VPW vss inv_p_7/ZN inv_p_7/I vdd vss inv_p
Xinv_p_8 vdd inv_p_8/VPW vss inv_p_8/ZN inv_p_8/I vdd vss inv_p
Xinv_p_9 vdd inv_p_9/VPW vss inv_p_9/ZN inv_p_9/I vdd vss inv_p
Xinv_p_10 vdd inv_p_10/VPW vss inv_p_10/ZN inv_p_10/I vdd vss inv_p
C0 inv_p_9/I inv_p_10/I 0.084161f
C1 vss inv_p_10/ZN 0.003326f
C2 inv_p_4/ZN inv_p_4/I 0.029333f
C3 vdd inv_p_4/ZN 0.159176f
C4 inv_p_0/ZN inv_p_3/I 0.002086f
C5 inv_p_9/I inv_p_10/ZN 0.028928f
C6 inv_p_4/I inv_p_5/I 0.084161f
C7 vdd inv_p_5/I 0.019437f
C8 inv_p_6/ZN inv_p_6/I 0.029333f
C9 inv_p_9/ZN inv_p_10/I 0.002086f
C10 inv_p_3/I inv_p_1/I 0.084161f
C11 inv_p_6/ZN vss 0.003326f
C12 inv_p_1/ZN inv_p_3/I 0.028928f
C13 inv_p_9/ZN inv_p_10/ZN 0.080571f
C14 inv_p_1/I inv_p_4/ZN 0.028928f
C15 inv_p_4/I inv_p_5/ZN 0.028928f
C16 vdd inv_p_5/ZN 0.159176f
C17 inv_p_6/ZN inv_p_7/I 0.002086f
C18 inv_p_1/ZN inv_p_4/ZN 0.080571f
C19 inv_p_2/ZN inv_p_2/I 0.029333f
C20 vdd inv_p_4/I 0.019437f
C21 inv_p_6/ZN inv_p_7/ZN 0.080571f
C22 vss inv_p_3/ZN 0.003326f
C23 inv_p_0/ZN vdd 0.184001f
C24 inv_p_2/I vss 0.164788f
C25 inv_p_2/ZN vss 0.005014f
C26 inv_p_6/I vss 0.166388f
C27 inv_p_0/I inv_p_3/ZN 0.028928f
C28 inv_p_1/I inv_p_4/I 0.084161f
C29 vdd inv_p_1/I 0.019437f
C30 inv_p_6/I inv_p_7/I 0.084161f
C31 inv_p_1/ZN inv_p_4/I 0.002086f
C32 inv_p_1/ZN vdd 0.159176f
C33 vss inv_p_8/I 0.166388f
C34 inv_p_7/I vss 0.166388f
C35 vss inv_p_9/I 0.166388f
C36 inv_p_7/I inv_p_8/I 0.084161f
C37 inv_p_9/I inv_p_8/I 0.084161f
C38 inv_p_6/I inv_p_7/ZN 0.028928f
C39 inv_p_0/I vss 0.170492f
C40 inv_p_1/ZN inv_p_1/I 0.029333f
C41 vss inv_p_8/ZN 0.003326f
C42 inv_p_6/ZN inv_p_5/I 0.028928f
C43 inv_p_7/ZN vss 0.003326f
C44 vdd inv_p_10/I 0.019437f
C45 inv_p_8/I inv_p_8/ZN 0.029333f
C46 vss inv_p_9/ZN 0.003326f
C47 inv_p_7/ZN inv_p_8/I 0.002086f
C48 inv_p_7/I inv_p_8/ZN 0.028928f
C49 inv_p_9/ZN inv_p_8/I 0.028928f
C50 inv_p_9/I inv_p_8/ZN 0.002086f
C51 inv_p_7/I inv_p_7/ZN 0.029333f
C52 inv_p_9/I inv_p_9/ZN 0.029333f
C53 vdd inv_p_10/ZN 0.159176f
C54 inv_p_3/I inv_p_3/ZN 0.029333f
C55 inv_p_6/ZN inv_p_5/ZN 0.080571f
C56 inv_p_7/ZN inv_p_8/ZN 0.080571f
C57 inv_p_9/ZN inv_p_8/ZN 0.080571f
C58 inv_p_6/ZN vdd 0.159176f
C59 vss inv_p_3/I 0.166388f
C60 inv_p_6/I inv_p_5/I 0.084161f
C61 vss inv_p_4/ZN 0.003326f
C62 vss inv_p_5/I 0.166388f
C63 inv_p_0/I inv_p_3/I 0.08416f
C64 inv_p_6/I inv_p_5/ZN 0.002086f
C65 vdd inv_p_3/ZN 0.159176f
C66 inv_p_2/I vdd 0.035575f
C67 inv_p_10/I inv_p_10/ZN 0.029333f
C68 vss inv_p_5/ZN 0.003326f
C69 inv_p_2/ZN vdd 0.174722f
C70 inv_p_0/ZN inv_p_3/ZN 0.080571f
C71 inv_p_6/I vdd 0.019437f
C72 inv_p_1/I inv_p_3/ZN 0.002086f
C73 vss inv_p_4/I 0.166388f
C74 vdd vss 0.009518f
C75 vdd inv_p_8/I 0.019437f
C76 inv_p_1/ZN inv_p_3/ZN 0.080571f
C77 inv_p_7/I vdd 0.019437f
C78 vdd inv_p_9/I 0.019437f
C79 inv_p_0/ZN vss 0.005399f
C80 inv_p_0/I vdd 0.026972f
C81 vdd inv_p_8/ZN 0.159176f
C82 inv_p_0/I inv_p_0/ZN 0.029333f
C83 vss inv_p_1/I 0.166388f
C84 inv_p_7/ZN vdd 0.159176f
C85 vdd inv_p_9/ZN 0.159176f
C86 inv_p_1/ZN vss 0.003326f
C87 inv_p_4/ZN inv_p_5/I 0.002086f
C88 inv_p_2/I inv_p_10/I 0.084161f
C89 inv_p_2/ZN inv_p_10/I 0.028928f
C90 inv_p_2/I inv_p_10/ZN 0.002086f
C91 inv_p_2/ZN inv_p_10/ZN 0.080571f
C92 inv_p_4/ZN inv_p_5/ZN 0.080571f
C93 vss inv_p_10/I 0.166388f
C94 inv_p_5/I inv_p_5/ZN 0.029333f
C95 vdd inv_p_3/I 0.019437f
C96 inv_p_10/ZN 0 0.131999f
C97 inv_p_10/I 0 0.64919f
C98 inv_p_9/ZN 0 0.131999f
C99 inv_p_9/I 0 0.64919f
C100 inv_p_8/ZN 0 0.131999f
C101 inv_p_8/I 0 0.64919f
C102 inv_p_7/ZN 0 0.131999f
C103 inv_p_7/I 0 0.64919f
C104 inv_p_6/ZN 0 0.131999f
C105 inv_p_6/I 0 0.64919f
C106 inv_p_5/ZN 0 0.131999f
C107 inv_p_5/I 0 0.64919f
C108 inv_p_4/ZN 0 0.131999f
C109 inv_p_4/I 0 0.64919f
C110 inv_p_3/ZN 0 0.131999f
C111 inv_p_3/I 0 0.64919f
C112 vss 0 3.02573f
C113 inv_p_2/ZN 0 0.206166f
C114 vdd 0 16.013325f
C115 inv_p_2/I 0 0.750024f
C116 inv_p_1/ZN 0 0.131999f
C117 inv_p_1/I 0 0.64919f
C118 inv_p_0/ZN 0 0.209411f
C119 inv_p_0/I 0 0.731246f
.ends

.subckt XM1_bs G D a_811_3903# S a_1507_3903#
X0 D G S a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D S 0.103318f
C1 G S 0.002993f
C2 G D 0.002993f
C3 S a_811_3903# 0.109266f
C4 G a_811_3903# 0.288275f
C5 D a_811_3903# 0.109266f
.ends

.subckt XM4_bs G D S VSUBS
X0 D G S S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D G 0.002993f
C1 S G 0.180042f
C2 D S 0.127372f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.66703f
.ends

.subckt XMs1_bs G D S a_n2855_n800#
X0 D G S a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D S 0.103318f
C1 G S 0.002993f
C2 D G 0.002993f
C3 D a_n2855_n800# 0.109266f
C4 S a_n2855_n800# 0.177295f
C5 G a_n2855_n800# 0.288368f
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668# VSUBS
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0fF c_width=8u c_length=8u
C0 m4_n3800_n668# m4_n3440_n548# 0.646322f
C1 m4_n3440_n548# VSUBS 1.17298f
C2 m4_n3800_n668# VSUBS 1.64833f
.ends

.subckt sw_cap_unit in out VSUBS
Xcap_mim_2p0fF_8JNR63_0 out in VSUBS cap_mim_2p0fF_8JNR63
C0 out VSUBS 1.17298f
C1 in VSUBS 1.64833f
.ends

.subckt sw_cap out in VSUBS
Xsw_cap_unit_0 in out VSUBS sw_cap_unit
Xsw_cap_unit_1 in out VSUBS sw_cap_unit
Xsw_cap_unit_2 in out VSUBS sw_cap_unit
Xsw_cap_unit_3 in out VSUBS sw_cap_unit
Xsw_cap_unit_4 in out VSUBS sw_cap_unit
C0 in out 2.231591f
C1 out VSUBS 6.064711f
C2 in VSUBS 7.39096f
.ends

.subckt XM3_bs G D S VSUBS
X0 S G D S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D S 0.127372f
C1 D G 0.002993f
C2 S G 0.175929f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.68221f
.ends

.subckt XMs_bs G D S a_846_4542#
X0 S G D a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D S 0.103318f
C1 D G 0.002993f
C2 S G 0.002993f
C3 D a_846_4542# 0.387117f
C4 G a_846_4542# 0.288368f
C5 S a_846_4542# 0.109266f
.ends

.subckt XM1_bs_inv G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt XM2_bs_inv G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.090564f
C1 D G 0.001764f
C2 S G 0.138578f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.08816f
C5 S VSUBS 1.2321f
.ends

.subckt bs_inv out in vdd vss
XXM1_bs_inv_0 in out vss XM1_bs_inv
XXM2_bs_inv_0 in out vdd vss XM2_bs_inv
C0 out in 0.057341f
C1 in vdd 0.034991f
C2 out vdd 0.086562f
C3 in vss 0.019395f
C4 out vss 0.056311f
C5 vss vdd 0.050184f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt XM2_bs G D a_811_3460# a_1507_3460# S
X0 S G D a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 G D 0.002993f
C1 S D 0.103318f
C2 G S 0.002993f
C3 D a_811_3460# 0.109266f
C4 G a_811_3460# 0.288275f
C5 S a_811_3460# 0.109266f
.ends

.subckt XMs2_bs G D a_n3988_469# S a_n3988_1165#
X0 D G S a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S D 0.103318f
C1 G D 0.002993f
C2 S G 0.002993f
C3 D a_n3988_469# 0.109266f
C4 S a_n3988_469# 0.109266f
C5 G a_n3988_469# 0.288275f
.ends

.subckt bootstrapped_sw_p in vss en enb vs vg vdd out vbsh vbsl
XXM1_bs_0 vg vbsl vss in vss XM1_bs
XXM4_bs_0 enb vg vbsh vss XM4_bs
XXMs1_bs_0 vdd vs vg vss XMs1_bs
Xsw_cap_0 vbsh vbsl vss sw_cap
XXM3_bs_0 vg vdd vbsh vss XM3_bs
XXMs_bs_0 vg out in vss XMs_bs
Xbs_inv_0 enb en vdd vss bs_inv
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 enb vss vss vs vss XMs2_bs
C0 vbsh out 0.106418f
C1 enb vg 0.612108f
C2 vdd vg 0.447811f
C3 enb vs 0.00376f
C4 enb vbsl 0.017274f
C5 vbsl vdd 0.005409f
C6 vbsh vg 0.225467f
C7 vg in 0.075595f
C8 enb vdd 0.448382f
C9 out vg 0.04429f
C10 vbsh vbsl 0.035648f
C11 vbsl in 0.299565f
C12 out vbsl 0.058082f
C13 vbsh enb 0.079647f
C14 vbsh vdd 0.216342f
C15 vs vg 0.01049f
C16 out vdd 0.017908f
C17 vbsl vg 0.046114f
C18 enb en 0.025502f
C19 vbsl vs 0.001422f
C20 vbsh in 0.008752f
C21 en vdd 0.062309f
C22 vs vss 0.072259f
C23 enb vss 1.595622f
C24 en vss 0.636177f
C25 out vss 1.088543f
C26 vdd vss 3.10752f
C27 vg vss 1.218874f
C28 vbsh vss 9.044386f
C29 vbsl vss 8.368301f
C30 in vss 0.308876f
.ends

.subckt dacp dum ctl7 ctl8 ctl9 ctl10 in sample ctl2 ctl1 carray_p_0/n0 carray_p_0/ndum
+ ctl4 ctl6 bootstrapped_sw_p_0/enb out bootstrapped_sw_p_0/vbsl ctl3 bootstrapped_sw_p_0/vg
+ bootstrapped_sw_p_0/vbsh carray_p_0/n8 carray_p_0/n9 ctl5 vdd vss
Xinv_renketu_p_0 ctl6 carray_p_0/n8 carray_p_0/n5 carray_p_0/n1 carray_p_0/ndum dum
+ ctl9 ctl3 carray_p_0/n7 carray_p_0/n0 carray_p_0/n4 ctl5 ctl10 carray_p_0/n9 ctl7
+ ctl2 ctl8 carray_p_0/n6 carray_p_0/n3 carray_p_0/n2 ctl1 ctl4 vss vdd inv_renketu_p
Xbootstrapped_sw_p_0 in vss sample bootstrapped_sw_p_0/enb bootstrapped_sw_p_0/vs
+ bootstrapped_sw_p_0/vg vdd out bootstrapped_sw_p_0/vbsh bootstrapped_sw_p_0/vbsl
+ bootstrapped_sw_p
C0 out carray_p_0/n8 0.420152p
C1 carray_p_0/n5 vdd 0.002151f
C2 out carray_p_0/n9 0.846161p
C3 carray_p_0/n5 carray_p_0/n2 0.208112f
C4 carray_p_0/ndum carray_p_0/n7 0.06073f
C5 vdd carray_p_0/n2 0.002151f
C6 carray_p_0/ndum carray_p_0/n4 0.025424f
C7 carray_p_0/n8 carray_p_0/n7 50.514606f
C8 carray_p_0/n9 carray_p_0/n7 29.51607f
C9 ctl7 ctl6 0.104537f
C10 ctl3 ctl4 0.104537f
C11 carray_p_0/n6 out 0.105055p
C12 carray_p_0/n8 carray_p_0/n4 2.84323f
C13 out carray_p_0/n3 13.201303f
C14 carray_p_0/n9 carray_p_0/n4 3.740571f
C15 ctl5 ctl4 0.104537f
C16 ctl9 ctl8 0.104537f
C17 bootstrapped_sw_p_0/vbsh out 0.137967f
C18 carray_p_0/n0 out 1.750611f
C19 carray_p_0/n1 out 3.367623f
C20 ctl10 ctl9 0.104537f
C21 carray_p_0/n6 carray_p_0/n7 34.66261f
C22 carray_p_0/n8 carray_p_0/ndum 0.097254f
C23 carray_p_0/n9 carray_p_0/ndum 0.127951f
C24 carray_p_0/n7 carray_p_0/n3 0.891504f
C25 sample carray_p_0/ndum 0.045492f
C26 carray_p_0/n5 out 52.565495f
C27 carray_p_0/n6 carray_p_0/n4 0.614078f
C28 carray_p_0/n0 carray_p_0/n7 0.06073f
C29 carray_p_0/n1 carray_p_0/n7 0.212822f
C30 carray_p_0/n4 carray_p_0/n3 26.229404f
C31 ctl2 ctl1 0.104537f
C32 carray_p_0/n9 carray_p_0/n8 87.43916f
C33 carray_p_0/n0 carray_p_0/n4 0.040502f
C34 carray_p_0/n1 carray_p_0/n4 0.142475f
C35 out carray_p_0/n2 6.640605f
C36 carray_p_0/n5 carray_p_0/n7 3.36878f
C37 carray_p_0/n6 carray_p_0/ndum 0.025424f
C38 carray_p_0/ndum carray_p_0/n3 0.025424f
C39 carray_p_0/n5 carray_p_0/n4 27.828503f
C40 carray_p_0/n6 carray_p_0/n8 11.2161f
C41 carray_p_0/n6 carray_p_0/n9 14.716781f
C42 carray_p_0/n1 carray_p_0/ndum 8.4982f
C43 vdd carray_p_0/n7 0.002151f
C44 carray_p_0/n8 carray_p_0/n3 1.46111f
C45 carray_p_0/n9 carray_p_0/n3 1.911225f
C46 carray_p_0/n7 carray_p_0/n2 0.485355f
C47 carray_p_0/n0 carray_p_0/n8 0.097254f
C48 vdd carray_p_0/n4 0.002151f
C49 carray_p_0/n1 carray_p_0/n8 0.28587f
C50 carray_p_0/n0 carray_p_0/n9 0.521489f
C51 carray_p_0/n1 carray_p_0/n9 0.350042f
C52 carray_p_0/n4 carray_p_0/n2 0.213209f
C53 carray_p_0/n5 carray_p_0/ndum 0.025424f
C54 ctl2 ctl3 0.104537f
C55 carray_p_0/n5 carray_p_0/n8 5.60732f
C56 carray_p_0/n5 carray_p_0/n9 7.39935f
C57 ctl7 ctl8 0.104537f
C58 carray_p_0/n6 carray_p_0/n3 0.336612f
C59 vdd carray_p_0/ndum 0.004405f
C60 carray_p_0/n6 carray_p_0/n0 0.025424f
C61 carray_p_0/ndum carray_p_0/n2 0.041162f
C62 carray_p_0/n6 carray_p_0/n1 0.142211f
C63 carray_p_0/n8 vdd 0.002151f
C64 carray_p_0/n0 carray_p_0/n3 0.051666f
C65 carray_p_0/n9 vdd 0.002151f
C66 carray_p_0/n1 carray_p_0/n3 0.145048f
C67 carray_p_0/n8 carray_p_0/n2 0.770227f
C68 carray_p_0/n1 carray_p_0/n0 8.476913f
C69 carray_p_0/n9 carray_p_0/n2 0.996681f
C70 carray_p_0/n5 carray_p_0/n6 28.925903f
C71 out carray_p_0/n7 0.210032p
C72 carray_p_0/n5 carray_p_0/n3 0.346757f
C73 carray_p_0/n5 carray_p_0/n0 0.025424f
C74 out carray_p_0/n4 26.32268f
C75 carray_p_0/n5 carray_p_0/n1 0.142354f
C76 carray_p_0/n6 vdd 0.002151f
C77 vdd carray_p_0/n3 0.002151f
C78 dum ctl1 0.104537f
C79 carray_p_0/n6 carray_p_0/n2 0.20799f
C80 bootstrapped_sw_p_0/vbsl out 0.061234f
C81 carray_p_0/n0 vdd 0.002151f
C82 carray_p_0/n3 carray_p_0/n2 23.177216f
C83 carray_p_0/n1 vdd 0.002151f
C84 carray_p_0/n0 carray_p_0/n2 0.099314f
C85 carray_p_0/n1 carray_p_0/n2 16.941956f
C86 out carray_p_0/ndum 1.640173f
C87 carray_p_0/n7 carray_p_0/n4 1.70387f
C88 ctl6 ctl5 0.104537f
C89 carray_p_0/n2 vss 30.239845f
C90 carray_p_0/n3 vss 33.722244f
C91 carray_p_0/n4 vss 39.983227f
C92 carray_p_0/n5 vss 47.48966f
C93 carray_p_0/n9 vss 14.559587f
C94 out vss -0.683569p
C95 carray_p_0/n8 vss 40.389835f
C96 carray_p_0/n7 vss 57.16868f
C97 carray_p_0/n6 vss 53.444874f
C98 carray_p_0/n0 vss 17.398035f
C99 carray_p_0/n1 vss 16.427063f
C100 bootstrapped_sw_p_0/vs vss 0.065021f
C101 bootstrapped_sw_p_0/enb vss 1.52928f
C102 sample vss 20.507322f
C103 bootstrapped_sw_p_0/vg vss 1.162193f
C104 bootstrapped_sw_p_0/vbsh vss 9.037161f
C105 bootstrapped_sw_p_0/vbsl vss 8.446682f
C106 in vss 0.297821f
C107 ctl9 vss 0.916847f
C108 ctl8 vss 0.916847f
C109 ctl7 vss 0.916847f
C110 ctl6 vss 0.916847f
C111 ctl5 vss 0.916847f
C112 ctl4 vss 0.916847f
C113 ctl3 vss 0.916847f
C114 ctl1 vss 0.916847f
C115 vdd vss 19.487324f
C116 ctl10 vss 1.146163f
C117 ctl2 vss 0.916847f
C118 carray_p_0/ndum vss 14.881927f
C119 dum vss 1.125528f
.ends

.subckt XM0_trim_right G D a_n484_399# a_n484_895# S
X0 S G D a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.14243f
C1 G S 0.005902f
C2 G D 0.011845f
C3 S a_n484_399# 0.098801f
C4 D a_n484_399# 0.215099f
C5 G a_n484_399# 0.21851f
.ends

.subckt XM1_trim_right G D a_n484_399# a_n484_895# S
X0 D G S a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.075352f
C1 G D 0.011845f
C2 G S 0.001764f
C3 D a_n484_399# 0.24117f
C4 S a_n484_399# 0.057381f
C5 G a_n484_399# 0.21851f
.ends

.subckt XM2_trim_right G D a_n375_n620# a_n375_n1116# S
X0 D G S a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.263094f
C1 G D 0.011804f
C2 G S 0.011804f
C3 D a_n375_n1116# 0.365155f
C4 S a_n375_n1116# 0.043869f
C5 G a_n375_n1116# 0.382504f
.ends

.subckt XM3_trim_right G D a_n778_n975# S
X0 D G S a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 D G S a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 S G D a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 S G 0.023608f
C1 D G 0.023608f
C2 S D 0.526188f
C3 D a_n778_n975# 0.557521f
C4 S a_n778_n975# 0.087739f
C5 G a_n778_n975# 0.718155f
.ends

.subckt XM4_trim_right G D a_1072_n1100# S
X0 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 S G D a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 D G 0.047215f
C1 S G 0.047215f
C2 D S 1.052376f
C3 S a_1072_n1100# 0.425359f
C4 D a_1072_n1100# 0.448822f
C5 G a_1072_n1100# 1.37423f
.ends

.subckt trim_switch_right XM3_trim_right_0/D XM0_trim_right_0/G XM4_trim_right_0/G
+ XM0_trim_right_0/D XM4_trim_right_0/D XM1_trim_right_0/G XM1_trim_right_0/D XM2_trim_right_0/G
+ XM2_trim_right_0/D XM3_trim_right_0/G VSUBS
XXM0_trim_right_0 XM0_trim_right_0/G XM0_trim_right_0/D VSUBS VSUBS VSUBS XM0_trim_right
XXM1_trim_right_0 XM1_trim_right_0/G XM1_trim_right_0/D VSUBS VSUBS VSUBS XM1_trim_right
XXM2_trim_right_0 XM2_trim_right_0/G XM2_trim_right_0/D VSUBS VSUBS VSUBS XM2_trim_right
XXM3_trim_right_0 XM3_trim_right_0/G XM3_trim_right_0/D VSUBS VSUBS XM3_trim_right
XXM4_trim_right_0 XM4_trim_right_0/G XM4_trim_right_0/D VSUBS VSUBS XM4_trim_right
C0 XM0_trim_right_0/D XM2_trim_right_0/D 0.039382f
C1 XM1_trim_right_0/D XM1_trim_right_0/G 0.07096f
C2 XM0_trim_right_0/G XM2_trim_right_0/G 0.041018f
C3 XM4_trim_right_0/D XM4_trim_right_0/G 0.272119f
C4 XM3_trim_right_0/G XM3_trim_right_0/D 0.092062f
C5 XM0_trim_right_0/D XM1_trim_right_0/D 0.027386f
C6 XM3_trim_right_0/G XM2_trim_right_0/G 0.027949f
C7 XM0_trim_right_0/G XM1_trim_right_0/G 0.123582f
C8 XM0_trim_right_0/G XM0_trim_right_0/D 0.07096f
C9 XM4_trim_right_0/D XM1_trim_right_0/D 0.00859f
C10 XM2_trim_right_0/D XM3_trim_right_0/D 0.040124f
C11 XM2_trim_right_0/G XM2_trim_right_0/D 0.014034f
C12 XM1_trim_right_0/G XM4_trim_right_0/G 0.02663f
C13 XM4_trim_right_0/D VSUBS 1.278621f
C14 XM4_trim_right_0/G VSUBS 1.959711f
C15 XM3_trim_right_0/D VSUBS 1.12292f
C16 XM3_trim_right_0/G VSUBS 1.128649f
C17 XM2_trim_right_0/D VSUBS 0.604021f
C18 XM2_trim_right_0/G VSUBS 0.637566f
C19 XM1_trim_right_0/D VSUBS 0.42776f
C20 XM1_trim_right_0/G VSUBS 0.407201f
C21 XM0_trim_right_0/D VSUBS 0.314559f
C22 XM0_trim_right_0/G VSUBS 0.388025f
.ends

.subckt trim_right d_4 d_1 d_0 d_2 d_3 trim_switch_right_0/XM3_trim_right_0/D trim_switch_right_0/XM2_trim_right_0/D
+ trim_switch_right_0/XM4_trim_right_0/D VSUBS ip
Xtrim_switch_right_0 trim_switch_right_0/XM3_trim_right_0/D d_0 d_4 trim_switch_right_0/XM0_trim_right_0/D
+ trim_switch_right_0/XM4_trim_right_0/D d_1 trim_switch_right_0/XM1_trim_right_0/D
+ d_2 trim_switch_right_0/XM2_trim_right_0/D d_3 VSUBS trim_switch_right
C0 trim_switch_right_0/XM4_trim_right_0/D ip 12.877382f
C1 trim_switch_right_0/XM2_trim_right_0/D trim_switch_right_0/XM1_trim_right_0/D 0.081094f
C2 d_4 trim_switch_right_0/XM2_trim_right_0/D 0.00312f
C3 trim_switch_right_0/XM3_trim_right_0/D trim_switch_right_0/XM0_trim_right_0/D 0.087807f
C4 ip trim_switch_right_0/XM2_trim_right_0/D 3.213024f
C5 trim_switch_right_0/XM4_trim_right_0/D trim_switch_right_0/XM3_trim_right_0/D 1.600475f
C6 d_0 trim_switch_right_0/XM2_trim_right_0/D 0.002632f
C7 ip trim_switch_right_0/XM1_trim_right_0/D 1.60623f
C8 trim_switch_right_0/XM4_trim_right_0/D trim_switch_right_0/XM0_trim_right_0/D 0.166348f
C9 trim_switch_right_0/XM3_trim_right_0/D trim_switch_right_0/XM2_trim_right_0/D 0.58337f
C10 trim_switch_right_0/XM2_trim_right_0/D trim_switch_right_0/XM0_trim_right_0/D 0.103369f
C11 trim_switch_right_0/XM3_trim_right_0/D trim_switch_right_0/XM1_trim_right_0/D 0.087807f
C12 trim_switch_right_0/XM1_trim_right_0/D trim_switch_right_0/XM0_trim_right_0/D 0.520979f
C13 trim_switch_right_0/XM4_trim_right_0/D trim_switch_right_0/XM2_trim_right_0/D 0.596682f
C14 trim_switch_right_0/XM4_trim_right_0/D trim_switch_right_0/XM1_trim_right_0/D 0.169398f
C15 ip trim_switch_right_0/XM3_trim_right_0/D 6.427485f
C16 d_1 trim_switch_right_0/XM2_trim_right_0/D 0.003137f
C17 ip trim_switch_right_0/XM0_trim_right_0/D 1.60623f
C18 d_0 trim_switch_right_0/XM0_trim_right_0/D 0.004139f
C19 d_1 trim_switch_right_0/XM1_trim_right_0/D 0.003099f
C20 d_4 VSUBS 1.64786f
C21 d_3 VSUBS 0.927186f
C22 d_2 VSUBS 0.513348f
C23 d_1 VSUBS 0.345562f
C24 d_0 VSUBS 0.33412f
C25 trim_switch_right_0/XM0_trim_right_0/D VSUBS 0.689164f
C26 trim_switch_right_0/XM1_trim_right_0/D VSUBS 0.727243f
C27 trim_switch_right_0/XM4_trim_right_0/D VSUBS 4.36705f
C28 ip VSUBS -5.906306f
C29 trim_switch_right_0/XM3_trim_right_0/D VSUBS 3.463846f
C30 trim_switch_right_0/XM2_trim_right_0/D VSUBS 2.037146f
.ends

.subckt XMdiff_com G D a_439_n1281# S
X0 D G S a_439_n1281# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 S G D a_439_n1281# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
C0 S G 0.003527f
C1 S D 0.137081f
C2 G D 0.003527f
C3 S a_439_n1281# 0.230614f
C4 D a_439_n1281# 0.02923f
C5 G a_439_n1281# 0.382694f
.ends

.subckt XMinp_com a_251_n1284# G D a_251_n788# S
X0 D G S a_251_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.06854f
C1 S G 0.001764f
C2 G D 0.001764f
C3 D a_251_n1284# 0.057707f
C4 S a_251_n1284# 0.057707f
C5 G a_251_n1284# 0.21851f
.ends

.subckt XMl4_com G D S w_n198_790# VSUBS
X0 D G S w_n198_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.06854f
C1 S w_n198_790# 0.008358f
C2 w_n198_790# D 0.010275f
C3 S G 0.001764f
C4 G D 0.001764f
C5 w_n198_790# G 0.131025f
C6 D VSUBS 0.047486f
C7 S VSUBS 0.049403f
C8 G VSUBS 0.087507f
C9 w_n198_790# VSUBS 1.54752f
.ends

.subckt XM4_com G D w_1022_790# S VSUBS
X0 D G S w_1022_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.06854f
C1 S w_1022_790# 0.021497f
C2 w_1022_790# D 0.022441f
C3 S G 0.001764f
C4 G D 0.001764f
C5 w_1022_790# G 0.132558f
C6 D VSUBS 0.043675f
C7 S VSUBS 0.043675f
C8 G VSUBS 0.08816f
C9 w_1022_790# VSUBS 1.17557f
.ends

.subckt XMl3_com G D w_n634_790# S VSUBS
X0 S G D w_n634_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.06854f
C1 D w_n634_790# 0.024248f
C2 w_n634_790# S 0.021497f
C3 D G 0.001764f
C4 G S 0.001764f
C5 w_n634_790# G 0.139286f
C6 S VSUBS 0.043675f
C7 D VSUBS 0.041759f
C8 G VSUBS 0.081314f
C9 w_n634_790# VSUBS 1.68331f
.ends

.subckt XM3_com G D w_n509_n1092# S VSUBS
X0 S G D w_n509_n1092# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.06854f
C1 D w_n509_n1092# 0.010275f
C2 w_n509_n1092# S 0.008358f
C3 D G 0.001764f
C4 G S 0.001764f
C5 w_n509_n1092# G 0.131025f
C6 S VSUBS 0.049403f
C7 D VSUBS 0.047486f
C8 G VSUBS 0.087507f
C9 w_n509_n1092# VSUBS 1.54752f
.ends

.subckt XMinn_com G a_719_n1284# D S a_719_n788#
X0 S G D a_719_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.06854f
C1 D G 0.001764f
C2 G S 0.001764f
C3 S a_719_n1284# 0.057707f
C4 D a_719_n1284# 0.057707f
C5 G a_719_n1284# 0.21851f
.ends

.subckt XM4_trim_left G D a_1072_n1100# S
X0 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 S G D a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 S G D a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 D G S a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 S G 0.047215f
C1 S D 1.052376f
C2 G D 0.047215f
C3 S a_1072_n1100# 0.425359f
C4 D a_1072_n1100# 0.448822f
C5 G a_1072_n1100# 1.37423f
.ends

.subckt XM3_trim_left G D a_n778_n975# S
X0 D G S a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 D G S a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 S G D a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.023608f
C1 D S 0.526188f
C2 G S 0.023608f
C3 D a_n778_n975# 0.557521f
C4 S a_n778_n975# 0.087739f
C5 G a_n778_n975# 0.718155f
.ends

.subckt XM2_trim_left G D a_n375_n620# a_n375_n1116# S
X0 D G S a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 S G D a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.263094f
C1 S G 0.011804f
C2 G D 0.011804f
C3 D a_n375_n1116# 0.365155f
C4 S a_n375_n1116# 0.043869f
C5 G a_n375_n1116# 0.382504f
.ends

.subckt XM1_trim_left G D a_n484_399# a_n484_895# S
X0 D G S a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.075352f
C1 S G 0.001764f
C2 G D 0.011845f
C3 D a_n484_399# 0.24117f
C4 S a_n484_399# 0.057381f
C5 G a_n484_399# 0.21851f
.ends

.subckt XM0_trim_left G D a_n484_399# a_n484_895# S
X0 S G D a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.14243f
C1 D G 0.011845f
C2 G S 0.005902f
C3 S a_n484_399# 0.098801f
C4 D a_n484_399# 0.215099f
C5 G a_n484_399# 0.21851f
.ends

.subckt trim_switch_left n1 n0 n2 n3 XM0_trim_left_0/G XM3_trim_left_0/G XM1_trim_left_0/G
+ XM4_trim_left_0/G n4 XM2_trim_left_0/G VSUBS
XXM4_trim_left_0 XM4_trim_left_0/G n4 VSUBS VSUBS XM4_trim_left
XXM3_trim_left_0 XM3_trim_left_0/G n3 VSUBS VSUBS XM3_trim_left
XXM2_trim_left_0 XM2_trim_left_0/G n2 VSUBS VSUBS VSUBS XM2_trim_left
XXM1_trim_left_0 XM1_trim_left_0/G n1 VSUBS VSUBS VSUBS XM1_trim_left
XXM0_trim_left_0 XM0_trim_left_0/G n0 VSUBS VSUBS VSUBS XM0_trim_left
C0 n1 n0 0.037109f
C1 XM2_trim_left_0/G XM0_trim_left_0/G 0.041018f
C2 n3 XM3_trim_left_0/G 0.092062f
C3 n2 n0 0.043322f
C4 XM4_trim_left_0/G n4 0.272119f
C5 n1 n4 0.01164f
C6 XM2_trim_left_0/G XM3_trim_left_0/G 0.027949f
C7 n3 n2 0.040124f
C8 XM1_trim_left_0/G XM0_trim_left_0/G 0.123582f
C9 XM1_trim_left_0/G XM4_trim_left_0/G 0.02663f
C10 XM2_trim_left_0/G n2 0.014034f
C11 XM1_trim_left_0/G n1 0.07096f
C12 XM0_trim_left_0/G n0 0.07096f
C13 n0 VSUBS 0.245304f
C14 XM0_trim_left_0/G VSUBS 0.388025f
C15 n1 VSUBS 0.34349f
C16 XM1_trim_left_0/G VSUBS 0.4072f
C17 n2 VSUBS 0.600267f
C18 XM2_trim_left_0/G VSUBS 0.637566f
C19 n3 VSUBS 1.12292f
C20 XM3_trim_left_0/G VSUBS 1.128649f
C21 n4 VSUBS 1.275608f
C22 XM4_trim_left_0/G VSUBS 1.959711f
.ends

.subckt trim_left in d_4 d_1 d_0 d_2 d_3 trim_switch_left_0/n3 trim_switch_left_0/n4
+ trim_switch_left_0/n2 VSUBS
Xtrim_switch_left_0 trim_switch_left_0/n1 trim_switch_left_0/n0 trim_switch_left_0/n2
+ trim_switch_left_0/n3 d_0 d_3 d_1 d_4 trim_switch_left_0/n4 d_2 VSUBS trim_switch_left
C0 trim_switch_left_0/n1 trim_switch_left_0/n3 0.087807f
C1 trim_switch_left_0/n1 in 1.60623f
C2 trim_switch_left_0/n2 d_4 0.00312f
C3 trim_switch_left_0/n0 trim_switch_left_0/n4 0.166348f
C4 trim_switch_left_0/n2 trim_switch_left_0/n4 0.596682f
C5 d_0 trim_switch_left_0/n0 0.004139f
C6 trim_switch_left_0/n2 d_0 0.002632f
C7 trim_switch_left_0/n1 trim_switch_left_0/n4 0.166348f
C8 in trim_switch_left_0/n3 6.427485f
C9 trim_switch_left_0/n2 trim_switch_left_0/n0 0.09943f
C10 trim_switch_left_0/n1 trim_switch_left_0/n0 0.511256f
C11 trim_switch_left_0/n1 trim_switch_left_0/n2 0.081094f
C12 trim_switch_left_0/n4 trim_switch_left_0/n3 1.600475f
C13 in trim_switch_left_0/n4 12.877382f
C14 d_1 trim_switch_left_0/n2 0.003137f
C15 trim_switch_left_0/n0 trim_switch_left_0/n3 0.087807f
C16 in trim_switch_left_0/n0 1.60623f
C17 trim_switch_left_0/n2 trim_switch_left_0/n3 0.58337f
C18 d_1 trim_switch_left_0/n1 0.003099f
C19 trim_switch_left_0/n2 in 3.213024f
C20 trim_switch_left_0/n0 VSUBS 0.60229f
C21 trim_switch_left_0/n1 VSUBS 0.624612f
C22 trim_switch_left_0/n4 VSUBS 4.36705f
C23 in VSUBS -5.906306f
C24 trim_switch_left_0/n3 VSUBS 3.463846f
C25 trim_switch_left_0/n2 VSUBS 2.037146f
C26 d_0 VSUBS 0.33412f
C27 d_1 VSUBS 0.345561f
C28 d_2 VSUBS 0.513348f
C29 d_3 VSUBS 0.927186f
C30 d_4 VSUBS 1.64786f
.ends

.subckt XM2_com G D w_n237_n1121# S VSUBS
X0 D G S w_n237_n1121# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.06854f
C1 D G 0.001764f
C2 S G 0.001764f
C3 D w_n237_n1121# 0.010275f
C4 S w_n237_n1121# 0.008358f
C5 G w_n237_n1121# 0.131025f
C6 D VSUBS 0.047486f
C7 S VSUBS 0.049403f
C8 G VSUBS 0.087507f
C9 w_n237_n1121# VSUBS 1.54752f
.ends

.subckt XMl2_com G D S a_n249_n1284#
X0 D G S a_n249_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D S 0.06854f
C1 D G 0.001764f
C2 S G 0.001764f
C3 D a_n249_n1284# 0.066395f
C4 S a_n249_n1284# 0.057707f
C5 G a_n249_n1284# 0.218606f
.ends

.subckt XM1_com G D S w_n1578_790# VSUBS
X0 S G D w_n1578_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.06854f
C1 S G 0.001764f
C2 D G 0.001764f
C3 S w_n1578_790# 0.021497f
C4 D w_n1578_790# 0.022441f
C5 G w_n1578_790# 0.132558f
C6 S VSUBS 0.043675f
C7 D VSUBS 0.043675f
C8 G VSUBS 0.08816f
C9 w_n1578_790# VSUBS 1.17557f
.ends

.subckt XMl1_com G D a_1224_n1284# S
X0 S G D a_1224_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.06854f
C1 S G 0.001764f
C2 D G 0.001764f
C3 S a_1224_n1284# 0.057707f
C4 D a_1224_n1284# 0.066395f
C5 G a_1224_n1284# 0.218606f
.ends

.subckt comparator vdd vp vn trim4 trim1 trim0 trimb4 trimb1 trimb0 trimb2 trimb3
+ diff in trim_right_0/trim_switch_right_0/XM2_trim_right_0/D trim_right_0/trim_switch_right_0/XM3_trim_right_0/D
+ clkc trim_right_0/trim_switch_right_0/XM4_trim_right_0/D outp outn trim_left_0/trim_switch_left_0/n4
+ trim_left_0/trim_switch_left_0/n3 trim_left_0/trim_switch_left_0/n2 ip trim3 trim2
+ vss
Xtrim_right_0 trimb4 trimb1 trimb0 trimb2 trimb3 trim_right_0/trim_switch_right_0/XM3_trim_right_0/D
+ trim_right_0/trim_switch_right_0/XM2_trim_right_0/D trim_right_0/trim_switch_right_0/XM4_trim_right_0/D
+ vss ip trim_right
XXMdiff_com_0 clkc diff vss vss XMdiff_com
XXMinp_com_0 vss vp ip vss diff XMinp_com
XXMl4_com_0 outn outp vdd vdd vss XMl4_com
XXM4_com_0 clkc ip vdd vdd vss XM4_com
XXMl3_com_0 outp outn vdd vdd vss XMl3_com
XXM3_com_0 clkc outp vdd vdd vss XM3_com
XXMinn_com_0 vn vss in diff vss XMinn_com
Xtrim_left_0 in trim4 trim1 trim0 trim2 trim3 trim_left_0/trim_switch_left_0/n3 trim_left_0/trim_switch_left_0/n4
+ trim_left_0/trim_switch_left_0/n2 vss trim_left
XXM2_com_0 clkc outn vdd vdd vss XM2_com
XXMl2_com_0 outn outp ip vss XMl2_com
XXM1_com_0 clkc in vdd vdd vss XM1_com
XXMl1_com_0 outp outn vss in XMl1_com
C0 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D trimb4 0.002224f
C1 in outp 0.016739f
C2 vp vn 0.217155f
C3 clkc outn 0.223756f
C4 vn vdd 0.059928f
C5 vp diff 0.004194f
C6 trimb4 trimb0 0.001193f
C7 ip outp 0.120151f
C8 trim_left_0/trim_switch_left_0/n1 trim_left_0/trim_switch_left_0/n4 0.032158f
C9 trim_left_0/trim_switch_left_0/n1 trim_left_0/trim_switch_left_0/n0 0.032158f
C10 vp clkc 0.104887f
C11 clkc vdd 0.233505f
C12 vn outp 0.238674f
C13 ip trim_right_0/trim_switch_right_0/XM3_trim_right_0/D 6.427209f
C14 diff outp 0.006112f
C15 ip trim_right_0/trim_switch_right_0/XM0_trim_right_0/D 1.606993f
C16 vn in 0.542295f
C17 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D ip 12.853658f
C18 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D trim_right_0/trim_switch_right_0/XM3_trim_right_0/D 0.241184f
C19 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D trim_right_0/trim_switch_right_0/XM0_trim_right_0/D 0.032158f
C20 in diff 0.133902f
C21 clkc outp 0.22388f
C22 trim_left_0/trim_switch_left_0/n1 in 1.606993f
C23 vp outn 0.212506f
C24 outn vdd 0.464524f
C25 trimb1 trimb4 0.420884f
C26 ip diff 0.133902f
C27 in clkc 0.467511f
C28 trim_left_0/trim_switch_left_0/n2 trim_left_0/trim_switch_left_0/n4 0.128631f
C29 trimb2 trimb0 0.78245f
C30 ip clkc 0.46748f
C31 vn diff 0.004194f
C32 vp vdd 0.059928f
C33 outn outp 1.248977f
C34 trimb3 trimb2 0.919951f
C35 trim_left_0/trim_switch_left_0/n4 trim_left_0/trim_switch_left_0/n0 0.032158f
C36 vn clkc 0.104888f
C37 in outn 0.120156f
C38 diff clkc 0.071648f
C39 trim_left_0/trim_switch_left_0/n4 trim1 0.001374f
C40 in trim_left_0/trim_switch_left_0/n2 3.21681f
C41 trim_left_0/trim_switch_left_0/n3 trim_left_0/trim_switch_left_0/n4 0.241184f
C42 trim_left_0/trim_switch_left_0/n4 trim4 0.002224f
C43 vp outp 0.245635f
C44 ip outn 0.016739f
C45 vdd outp 0.441033f
C46 ip trim_right_0/trim_switch_right_0/XM2_trim_right_0/D 3.21681f
C47 trim_right_0/trim_switch_right_0/XM1_trim_right_0/D ip 1.606993f
C48 trim_right_0/trim_switch_right_0/XM1_trim_right_0/D trim_right_0/trim_switch_right_0/XM0_trim_right_0/D 0.032158f
C49 trim3 trim2 0.919951f
C50 trim0 trim2 0.78245f
C51 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D trimb1 0.001374f
C52 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D trim_right_0/trim_switch_right_0/XM2_trim_right_0/D 0.128631f
C53 trim4 trim1 0.420884f
C54 in vdd 0.088929f
C55 in trim_left_0/trim_switch_left_0/n4 12.853658f
C56 trim_right_0/trim_switch_right_0/XM1_trim_right_0/D trim_right_0/trim_switch_right_0/XM4_trim_right_0/D 0.032158f
C57 vn outn 0.198266f
C58 in trim_left_0/trim_switch_left_0/n0 1.606993f
C59 vp ip 0.542294f
C60 trimb1 trimb0 0.720503f
C61 diff outn 0.003297f
C62 trim0 trim1 0.720503f
C63 ip vdd 0.088929f
C64 trim0 trim4 0.001193f
C65 in trim_left_0/trim_switch_left_0/n3 6.427209f
C66 outn vss 2.441227f
C67 outp vss 2.475127f
C68 vdd vss 7.878819f
C69 trim_left_0/trim_switch_left_0/n0 vss 0.59175f
C70 trim_left_0/trim_switch_left_0/n1 vss 0.614476f
C71 trim_left_0/trim_switch_left_0/n4 vss 4.199547f
C72 in vss -4.381556f
C73 trim_left_0/trim_switch_left_0/n3 vss 3.310533f
C74 trim_left_0/trim_switch_left_0/n2 vss 1.980191f
C75 trim0 vss 0.985146f
C76 trim1 vss 0.998489f
C77 trim2 vss 1.41065f
C78 trim3 vss 2.983196f
C79 trim4 vss 2.263372f
C80 diff vss 0.21339f
C81 vn vss 1.131511f
C82 vp vss 1.115711f
C83 clkc vss 4.18047f
C84 trimb4 vss 2.263372f
C85 trimb3 vss 2.983196f
C86 trimb2 vss 1.41065f
C87 trimb1 vss 0.99849f
C88 trimb0 vss 0.985146f
C89 trim_right_0/trim_switch_right_0/XM0_trim_right_0/D vss 0.677622f
C90 trim_right_0/trim_switch_right_0/XM1_trim_right_0/D vss 0.716105f
C91 trim_right_0/trim_switch_right_0/XM4_trim_right_0/D vss 4.199547f
C92 ip vss -4.381578f
C93 trim_right_0/trim_switch_right_0/XM3_trim_right_0/D vss 3.310533f
C94 trim_right_0/trim_switch_right_0/XM2_trim_right_0/D vss 1.980191f
.ends

.subckt inv_n VNW VPW VSS ZN I VDD VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VDD I 0.074838f
C1 VNW I 0.285482f
C2 VSS I 0.091531f
C3 ZN I 0.58604f
C4 VNW VDD 0.082022f
C5 VSS VDD 0.029045f
C6 ZN VDD 0.271625f
C7 VSS VNW 0.006277f
C8 ZN VNW 0.023676f
C9 VSS ZN 0.180794f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu_n inv_n_8/I inv_n_1/I inv_n_4/ZN inv_n_1/ZN inv_n_3/I inv_n_5/I
+ inv_n_7/I inv_n_9/ZN inv_n_6/ZN inv_n_10/ZN inv_n_3/ZN inv_n_0/ZN inv_n_0/I inv_n_10/I
+ inv_n_2/I inv_n_9/I inv_n_4/I vdd inv_n_7/ZN inv_n_8/ZN inv_n_5/ZN inv_n_6/I inv_n_2/ZN
+ vss
Xinv_n_0 vdd inv_n_0/VPW vss inv_n_0/ZN inv_n_0/I vdd vss inv_n
Xinv_n_1 vdd inv_n_1/VPW vss inv_n_1/ZN inv_n_1/I vdd vss inv_n
Xinv_n_2 vdd inv_n_2/VPW vss inv_n_2/ZN inv_n_2/I vdd vss inv_n
Xinv_n_3 vdd inv_n_3/VPW vss inv_n_3/ZN inv_n_3/I vdd vss inv_n
Xinv_n_4 vdd inv_n_4/VPW vss inv_n_4/ZN inv_n_4/I vdd vss inv_n
Xinv_n_5 vdd inv_n_5/VPW vss inv_n_5/ZN inv_n_5/I vdd vss inv_n
Xinv_n_6 vdd inv_n_6/VPW vss inv_n_6/ZN inv_n_6/I vdd vss inv_n
Xinv_n_7 vdd inv_n_7/VPW vss inv_n_7/ZN inv_n_7/I vdd vss inv_n
Xinv_n_8 vdd inv_n_8/VPW vss inv_n_8/ZN inv_n_8/I vdd vss inv_n
Xinv_n_9 vdd inv_n_9/VPW vss inv_n_9/ZN inv_n_9/I vdd vss inv_n
Xinv_n_10 vdd inv_n_10/VPW vss inv_n_10/ZN inv_n_10/I vdd vss inv_n
C0 inv_n_6/ZN inv_n_5/I 0.028928f
C1 inv_n_9/ZN inv_n_9/I 0.029333f
C2 inv_n_10/ZN vss 0.003326f
C3 inv_n_0/ZN vdd 0.184001f
C4 inv_n_7/I inv_n_7/ZN 0.029333f
C5 inv_n_4/ZN inv_n_5/I 0.002086f
C6 inv_n_8/I vdd 0.019437f
C7 inv_n_10/I inv_n_9/I 0.084161f
C8 inv_n_4/I inv_n_1/I 0.084161f
C9 vdd inv_n_1/ZN 0.159176f
C10 inv_n_8/I inv_n_7/ZN 0.002086f
C11 inv_n_5/ZN inv_n_5/I 0.029333f
C12 vdd inv_n_7/ZN 0.159176f
C13 inv_n_6/I inv_n_5/I 0.084161f
C14 vdd inv_n_2/I 0.035575f
C15 vss inv_n_6/ZN 0.003326f
C16 vss inv_n_9/ZN 0.003326f
C17 inv_n_3/I inv_n_3/ZN 0.029333f
C18 inv_n_2/ZN inv_n_10/I 0.028928f
C19 inv_n_8/ZN inv_n_7/I 0.028928f
C20 inv_n_4/I inv_n_5/I 0.084161f
C21 inv_n_4/ZN vss 0.003326f
C22 inv_n_3/I vss 0.166388f
C23 inv_n_10/ZN inv_n_9/ZN 0.080571f
C24 inv_n_10/I vss 0.166388f
C25 inv_n_3/I inv_n_0/I 0.08416f
C26 vdd inv_n_1/I 0.019437f
C27 inv_n_10/ZN inv_n_10/I 0.029333f
C28 inv_n_8/I inv_n_8/ZN 0.029333f
C29 inv_n_1/ZN inv_n_1/I 0.029333f
C30 inv_n_8/ZN vdd 0.159176f
C31 vss inv_n_5/ZN 0.003326f
C32 vss inv_n_6/I 0.166388f
C33 inv_n_8/I inv_n_9/I 0.084161f
C34 vdd inv_n_9/I 0.019437f
C35 inv_n_8/ZN inv_n_7/ZN 0.080571f
C36 vdd inv_n_5/I 0.019437f
C37 inv_n_4/I vss 0.166388f
C38 vss inv_n_7/I 0.166388f
C39 inv_n_10/I inv_n_9/ZN 0.002086f
C40 inv_n_0/ZN inv_n_3/ZN 0.080571f
C41 vss inv_n_0/ZN 0.005399f
C42 inv_n_2/ZN vdd 0.174722f
C43 inv_n_6/ZN inv_n_5/ZN 0.080571f
C44 vdd inv_n_3/ZN 0.159176f
C45 inv_n_0/ZN inv_n_0/I 0.029333f
C46 inv_n_8/I vss 0.166388f
C47 inv_n_6/I inv_n_6/ZN 0.029333f
C48 inv_n_4/ZN inv_n_5/ZN 0.080571f
C49 vss vdd 0.009518f
C50 inv_n_3/ZN inv_n_1/ZN 0.080571f
C51 vdd inv_n_0/I 0.026972f
C52 vss inv_n_1/ZN 0.003326f
C53 inv_n_10/ZN vdd 0.159176f
C54 inv_n_8/ZN inv_n_9/I 0.002086f
C55 inv_n_4/ZN inv_n_4/I 0.029333f
C56 inv_n_2/ZN inv_n_2/I 0.029333f
C57 vss inv_n_7/ZN 0.003326f
C58 vss inv_n_2/I 0.164788f
C59 inv_n_7/I inv_n_6/ZN 0.002086f
C60 inv_n_6/I inv_n_5/ZN 0.002086f
C61 inv_n_10/ZN inv_n_2/I 0.002086f
C62 inv_n_4/I inv_n_5/ZN 0.028928f
C63 inv_n_3/ZN inv_n_1/I 0.002086f
C64 vss inv_n_1/I 0.166388f
C65 inv_n_3/I inv_n_0/ZN 0.002086f
C66 inv_n_8/I inv_n_9/ZN 0.028928f
C67 vdd inv_n_6/ZN 0.159176f
C68 vdd inv_n_9/ZN 0.159176f
C69 inv_n_4/ZN vdd 0.159176f
C70 vss inv_n_8/ZN 0.003326f
C71 inv_n_3/I vdd 0.019437f
C72 inv_n_7/I inv_n_6/I 0.084161f
C73 inv_n_10/I vdd 0.019437f
C74 inv_n_4/ZN inv_n_1/ZN 0.080571f
C75 inv_n_3/I inv_n_1/ZN 0.028928f
C76 inv_n_6/ZN inv_n_7/ZN 0.080571f
C77 vss inv_n_9/I 0.166388f
C78 vss inv_n_5/I 0.166388f
C79 vdd inv_n_5/ZN 0.159176f
C80 inv_n_10/ZN inv_n_9/I 0.028928f
C81 vdd inv_n_6/I 0.019437f
C82 inv_n_10/I inv_n_2/I 0.084161f
C83 inv_n_4/I vdd 0.019437f
C84 inv_n_6/I inv_n_7/ZN 0.028928f
C85 inv_n_4/ZN inv_n_1/I 0.028928f
C86 inv_n_4/I inv_n_1/ZN 0.002086f
C87 inv_n_2/ZN vss 0.005014f
C88 inv_n_3/I inv_n_1/I 0.084161f
C89 inv_n_8/ZN inv_n_9/ZN 0.080571f
C90 vss inv_n_3/ZN 0.003326f
C91 inv_n_8/I inv_n_7/I 0.084161f
C92 vdd inv_n_7/I 0.019437f
C93 inv_n_3/ZN inv_n_0/I 0.028928f
C94 inv_n_2/ZN inv_n_10/ZN 0.080571f
C95 vss inv_n_0/I 0.170492f
C96 inv_n_10/ZN 0 0.131999f
C97 inv_n_10/I 0 0.64919f
C98 inv_n_9/ZN 0 0.131999f
C99 inv_n_9/I 0 0.64919f
C100 inv_n_8/ZN 0 0.131999f
C101 inv_n_8/I 0 0.64919f
C102 inv_n_7/ZN 0 0.131999f
C103 inv_n_7/I 0 0.64919f
C104 inv_n_6/ZN 0 0.131999f
C105 inv_n_6/I 0 0.64919f
C106 inv_n_5/ZN 0 0.131999f
C107 inv_n_5/I 0 0.64919f
C108 inv_n_4/ZN 0 0.131999f
C109 inv_n_4/I 0 0.64919f
C110 inv_n_3/ZN 0 0.131999f
C111 inv_n_3/I 0 0.64919f
C112 vss 0 3.02573f
C113 inv_n_2/ZN 0 0.206166f
C114 vdd 0 16.013325f
C115 inv_n_2/I 0 0.750024f
C116 inv_n_1/ZN 0 0.131999f
C117 inv_n_1/I 0 0.64919f
C118 inv_n_0/ZN 0 0.209411f
C119 inv_n_0/I 0 0.731246f
.ends

.subckt XM1_bs$1 G D a_811_3903# S a_1507_3903#
X0 D G S a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D G 0.002993f
C1 G S 0.002993f
C2 D S 0.103318f
C3 S a_811_3903# 0.109266f
C4 G a_811_3903# 0.288275f
C5 D a_811_3903# 0.109266f
.ends

.subckt XMs1_bs$1 G D S a_n2855_n800#
X0 D G S a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 G D 0.002993f
C1 S D 0.103318f
C2 S G 0.002993f
C3 D a_n2855_n800# 0.109266f
C4 S a_n2855_n800# 0.177295f
C5 G a_n2855_n800# 0.288368f
.ends

.subckt XM2_bs$1 G D a_811_3460# a_1507_3460# S
X0 S G D a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S G 0.002993f
C1 G D 0.002993f
C2 S D 0.103318f
C3 D a_811_3460# 0.109266f
C4 G a_811_3460# 0.288275f
C5 S a_811_3460# 0.109266f
.ends

.subckt XMs2_bs$1 G D a_n3988_469# S a_n3988_1165#
X0 D G S a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 G S 0.002993f
C1 S D 0.103318f
C2 G D 0.002993f
C3 D a_n3988_469# 0.109266f
C4 S a_n3988_469# 0.109266f
C5 G a_n3988_469# 0.288275f
.ends

.subckt XM3_bs$1 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S D 0.127372f
C1 G D 0.002993f
C2 G S 0.175929f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.68221f
.ends

.subckt cap_mim_2p0fF_8JNR63$1 m4_n3440_n548# m4_n3800_n668# VSUBS
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0fF c_width=8u c_length=8u
C0 m4_n3440_n548# m4_n3800_n668# 0.646322f
C1 m4_n3440_n548# VSUBS 1.17298f
C2 m4_n3800_n668# VSUBS 1.64833f
.ends

.subckt sw_cap_unit$1 in out VSUBS
Xcap_mim_2p0fF_8JNR63_0 out in VSUBS cap_mim_2p0fF_8JNR63$1
C0 out VSUBS 1.17298f
C1 in VSUBS 1.64833f
.ends

.subckt sw_cap$1 out in VSUBS
Xsw_cap_unit$1_0 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_1 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_2 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_3 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_4 in out VSUBS sw_cap_unit$1
C0 out in 2.231591f
C1 out VSUBS 6.064711f
C2 in VSUBS 7.39096f
.ends

.subckt XM2_bs_inv$1 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G S 0.138578f
C1 D S 0.090564f
C2 G D 0.001764f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.08816f
C5 S VSUBS 1.2321f
.ends

.subckt XM1_bs_inv$1 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt bs_inv$1 out in vdd vss
XXM2_bs_inv$1_0 in out vdd vss XM2_bs_inv$1
XXM1_bs_inv$1_0 in out vss XM1_bs_inv$1
C0 in vss 0.019395f
C1 vss out 0.056311f
C2 in out 0.057341f
C3 vss vdd 0.050184f
C4 in vdd 0.034991f
C5 out vdd 0.086562f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt XM4_bs$1 G D S VSUBS
X0 D G S S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S G 0.180042f
C1 S D 0.127372f
C2 G D 0.002993f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.66703f
.ends

.subckt XMs_bs$1 G D S a_846_4542#
X0 S G D a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S G 0.002993f
C1 S D 0.103318f
C2 G D 0.002993f
C3 D a_846_4542# 0.387117f
C4 G a_846_4542# 0.288368f
C5 S a_846_4542# 0.109266f
.ends

.subckt bootstrapped_sw_n in en enb vs vg vss out vdd vbsl vbsh
XXM1_bs$1_0 vg vbsl vss in vss XM1_bs$1
XXMs1_bs$1_0 vdd vs vg vss XMs1_bs$1
XXM2_bs$1_0 enb vbsl vss vss vss XM2_bs$1
XXMs2_bs$1_0 enb vss vss vs vss XMs2_bs$1
XXM3_bs$1_0 vg vdd vbsh vss XM3_bs$1
Xsw_cap$1_0 vbsh vbsl vss sw_cap$1
Xbs_inv$1_0 enb en vdd vss bs_inv$1
XXM4_bs$1_0 enb vg vbsh vss XM4_bs$1
XXMs_bs$1_0 vg out in vss XMs_bs$1
C0 vdd en 0.062309f
C1 vbsh out 0.106418f
C2 in vg 0.075595f
C3 enb en 0.025502f
C4 out vg 0.04429f
C5 vdd vbsl 0.005409f
C6 vs vbsl 0.001422f
C7 vbsl enb 0.017274f
C8 vbsh vbsl 0.035648f
C9 vbsl in 0.299565f
C10 vbsl vg 0.046114f
C11 vdd enb 0.448382f
C12 vdd vbsh 0.216342f
C13 vs enb 0.00376f
C14 vbsh enb 0.079647f
C15 vbsl out 0.058082f
C16 vdd vg 0.447811f
C17 vs vg 0.01049f
C18 vbsh in 0.008752f
C19 enb vg 0.612108f
C20 vbsh vg 0.225467f
C21 vdd out 0.017908f
C22 out vss 1.088543f
C23 en vss 0.636177f
C24 vbsh vss 9.044386f
C25 vbsl vss 8.368301f
C26 vdd vss 3.10752f
C27 vg vss 1.218874f
C28 vs vss 0.072259f
C29 enb vss 1.595622f
C30 in vss 0.308876f
.ends

.subckt dacn ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10 in bootstrapped_sw_n_0/vg
+ bootstrapped_sw_n_0/enb carray_n_0/n9 sample carray_n_0/n0 out carray_n_0/n8 dum
+ vdd bootstrapped_sw_n_0/vbsh vss bootstrapped_sw_n_0/vbsl carray_n_0/ndum
Xinv_renketu_n_0 ctl7 ctl2 carray_n_0/n3 carray_n_0/n2 ctl1 ctl4 ctl6 carray_n_0/n8
+ carray_n_0/n5 carray_n_0/n9 carray_n_0/n1 carray_n_0/ndum dum ctl9 ctl10 ctl8 ctl3
+ vdd carray_n_0/n6 carray_n_0/n7 carray_n_0/n4 ctl5 carray_n_0/n0 vss inv_renketu_n
Xbootstrapped_sw_n_0 in sample bootstrapped_sw_n_0/enb bootstrapped_sw_n_0/vs bootstrapped_sw_n_0/vg
+ vss out vdd bootstrapped_sw_n_0/vbsl bootstrapped_sw_n_0/vbsh bootstrapped_sw_n
C0 carray_n_0/n4 carray_n_0/n7 1.70387f
C1 carray_n_0/n0 vdd 0.002151f
C2 carray_n_0/n2 carray_n_0/n5 0.208112f
C3 carray_n_0/n6 carray_n_0/n7 34.66261f
C4 carray_n_0/n4 vdd 0.002151f
C5 carray_n_0/ndum out 1.640173f
C6 carray_n_0/n2 carray_n_0/n8 0.770227f
C7 carray_n_0/n5 carray_n_0/n9 7.39935f
C8 vdd carray_n_0/n6 0.002151f
C9 carray_n_0/n1 carray_n_0/n7 0.212822f
C10 carray_n_0/n8 carray_n_0/n9 87.43916f
C11 carray_n_0/n5 carray_n_0/n0 0.025424f
C12 carray_n_0/n2 carray_n_0/n3 23.177216f
C13 vdd carray_n_0/n1 0.002151f
C14 carray_n_0/n4 carray_n_0/n5 27.828503f
C15 carray_n_0/n0 carray_n_0/n8 0.097254f
C16 ctl10 ctl9 0.104537f
C17 carray_n_0/n3 carray_n_0/n9 1.911225f
C18 carray_n_0/n4 carray_n_0/n8 2.84323f
C19 carray_n_0/n5 carray_n_0/n6 28.925903f
C20 bootstrapped_sw_n_0/vbsh out 0.137967f
C21 carray_n_0/n2 out 6.640605f
C22 carray_n_0/n3 carray_n_0/n0 0.051666f
C23 vdd carray_n_0/n7 0.002151f
C24 sample carray_n_0/ndum 0.045492f
C25 carray_n_0/n6 carray_n_0/n8 11.2161f
C26 carray_n_0/n5 carray_n_0/n1 0.142354f
C27 carray_n_0/n2 carray_n_0/ndum 0.041162f
C28 carray_n_0/n4 carray_n_0/n3 26.229404f
C29 out carray_n_0/n9 0.846161p
C30 carray_n_0/n1 carray_n_0/n8 0.28587f
C31 ctl7 ctl6 0.104537f
C32 carray_n_0/n3 carray_n_0/n6 0.336612f
C33 carray_n_0/ndum carray_n_0/n9 0.127951f
C34 ctl1 ctl2 0.104537f
C35 carray_n_0/n0 out 1.750611f
C36 carray_n_0/n4 out 26.32268f
C37 carray_n_0/n3 carray_n_0/n1 0.145048f
C38 carray_n_0/n5 carray_n_0/n7 3.36878f
C39 carray_n_0/ndum carray_n_0/n4 0.025424f
C40 carray_n_0/n7 carray_n_0/n8 50.514606f
C41 carray_n_0/n6 out 0.105055p
C42 carray_n_0/n5 vdd 0.002151f
C43 carray_n_0/ndum carray_n_0/n6 0.025424f
C44 vdd carray_n_0/n8 0.002151f
C45 carray_n_0/n1 out 3.367623f
C46 carray_n_0/n3 carray_n_0/n7 0.891504f
C47 ctl1 dum 0.104537f
C48 carray_n_0/n2 carray_n_0/n9 0.996681f
C49 carray_n_0/ndum carray_n_0/n1 8.4982f
C50 carray_n_0/n3 vdd 0.002151f
C51 ctl6 ctl5 0.104537f
C52 carray_n_0/n2 carray_n_0/n0 0.099314f
C53 carray_n_0/n2 carray_n_0/n4 0.213209f
C54 carray_n_0/n7 out 0.210032p
C55 carray_n_0/n5 carray_n_0/n8 5.60732f
C56 carray_n_0/n0 carray_n_0/n9 0.521489f
C57 carray_n_0/ndum carray_n_0/n7 0.06073f
C58 carray_n_0/n2 carray_n_0/n6 0.20799f
C59 carray_n_0/n4 carray_n_0/n9 3.740571f
C60 carray_n_0/n3 carray_n_0/n5 0.346757f
C61 bootstrapped_sw_n_0/vbsl out 0.061234f
C62 carray_n_0/ndum vdd 0.004405f
C63 carray_n_0/n2 carray_n_0/n1 16.941956f
C64 carray_n_0/n6 carray_n_0/n9 14.716781f
C65 carray_n_0/n4 carray_n_0/n0 0.040502f
C66 carray_n_0/n3 carray_n_0/n8 1.46111f
C67 carray_n_0/n0 carray_n_0/n6 0.025424f
C68 carray_n_0/n1 carray_n_0/n9 0.350042f
C69 ctl3 ctl4 0.104537f
C70 carray_n_0/n5 out 52.565495f
C71 carray_n_0/n4 carray_n_0/n6 0.614078f
C72 ctl4 ctl5 0.104537f
C73 ctl3 ctl2 0.104537f
C74 carray_n_0/n0 carray_n_0/n1 8.476913f
C75 carray_n_0/ndum carray_n_0/n5 0.025424f
C76 carray_n_0/n2 carray_n_0/n7 0.485355f
C77 carray_n_0/n8 out 0.420152p
C78 carray_n_0/n4 carray_n_0/n1 0.142475f
C79 ctl9 ctl8 0.104537f
C80 carray_n_0/ndum carray_n_0/n8 0.097254f
C81 carray_n_0/n2 vdd 0.002151f
C82 carray_n_0/n7 carray_n_0/n9 29.51607f
C83 carray_n_0/n3 out 13.201303f
C84 ctl7 ctl8 0.104537f
C85 carray_n_0/n1 carray_n_0/n6 0.142211f
C86 vdd carray_n_0/n9 0.002151f
C87 carray_n_0/n0 carray_n_0/n7 0.06073f
C88 carray_n_0/ndum carray_n_0/n3 0.025424f
C89 carray_n_0/n9 vss 14.559587f
C90 out vss -0.683569p
C91 carray_n_0/n8 vss 40.389835f
C92 carray_n_0/n7 vss 57.16868f
C93 carray_n_0/n6 vss 53.444874f
C94 carray_n_0/n0 vss 17.398035f
C95 carray_n_0/n1 vss 16.427063f
C96 carray_n_0/n2 vss 30.239845f
C97 carray_n_0/n3 vss 33.722244f
C98 carray_n_0/n4 vss 39.983227f
C99 carray_n_0/n5 vss 47.48966f
C100 sample vss 20.507322f
C101 bootstrapped_sw_n_0/vbsh vss 9.037161f
C102 bootstrapped_sw_n_0/vbsl vss 8.446682f
C103 bootstrapped_sw_n_0/vg vss 1.162193f
C104 bootstrapped_sw_n_0/vs vss 0.065021f
C105 bootstrapped_sw_n_0/enb vss 1.52928f
C106 in vss 0.297821f
C107 ctl9 vss 0.916847f
C108 ctl8 vss 0.916847f
C109 ctl7 vss 0.916847f
C110 ctl6 vss 0.916847f
C111 ctl5 vss 0.916847f
C112 ctl4 vss 0.916847f
C113 ctl3 vss 0.916847f
C114 ctl1 vss 0.916847f
C115 vdd vss 19.487324f
C116 ctl10 vss 1.146163f
C117 ctl2 vss 0.916847f
C118 carray_n_0/ndum vss 14.881927f
C119 dum vss 1.125528f
.ends

.subckt cap_mim_2p0fF_RCWXT2$1 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3240_n3120# m4_n3120_n3000# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30_flip cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$1
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_RCWXT2 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3240_n3120# m4_n3120_n3000# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap1 vss vdd VSUBS
Xmim_cap_30_30_flip_233 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_222 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_200 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_211 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_68 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_57 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_79 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_13 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_24 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_46 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_35 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_213 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_224 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_202 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_235 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_212 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_234 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_223 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_201 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_58 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_69 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_14 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_25 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_47 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_36 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_214 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_225 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_203 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_236 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_224 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_213 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_235 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_202 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_59 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_15 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_48 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_26 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_37 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_226 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_204 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_237 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_215 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_225 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_214 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_236 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_203 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_16 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_49 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_38 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_27 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_227 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_238 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_205 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_216 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_226 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_215 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_237 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_204 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_17 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_28 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_39 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_228 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_217 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_239 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_206 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_227 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_216 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_238 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_205 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_18 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_29 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_229 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_218 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_207 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_228 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_217 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_206 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_239 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_19 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_219 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_208 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_229 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_218 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_207 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_209 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_219 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_208 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_190 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_209 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_90 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_180 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_191 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_80 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_91 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_190 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_170 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_181 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_192 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_81 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_70 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_92 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_0 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_191 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_180 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_0 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_160 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_193 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_182 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_171 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_60 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_82 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_71 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_93 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_1 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_170 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_192 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_181 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_1 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_183 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_172 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_150 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_194 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_161 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_83 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_72 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_94 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_50 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_61 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_2 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_160 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_193 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_182 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_171 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_2 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_173 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_162 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_184 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_195 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_140 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_151 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_73 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_84 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_95 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_51 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_40 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_62 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_3 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_161 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_172 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_194 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_183 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_150 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_3 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_174 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_152 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_141 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_196 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_130 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_185 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_163 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_30 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_74 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_85 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_52 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_96 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_41 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_63 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_4 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_151 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_162 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_140 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_173 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_184 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_195 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_4 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_131 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_120 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_153 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_186 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_142 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_197 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_164 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_175 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_31 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_75 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_20 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_64 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_86 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_42 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_53 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_97 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_5 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_152 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_163 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_141 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_174 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_130 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_196 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_185 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_5 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_154 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_176 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_165 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_110 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_132 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_121 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_143 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_198 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_187 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_76 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_21 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_65 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_10 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_32 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_43 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_54 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_87 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_98 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_6 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_153 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_164 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_175 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_131 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_142 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_120 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_197 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_186 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_6 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_155 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_166 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_111 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_100 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_133 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_144 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_122 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_199 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_188 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_177 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_77 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_22 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_66 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_11 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_99 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_33 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_44 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_55 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_88 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_7 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_110 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_121 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_154 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_176 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_143 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_198 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_187 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_132 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_165 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_7 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_156 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_167 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_178 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_101 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_112 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_145 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_123 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_189 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_134 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_23 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_67 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_78 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_12 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_34 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_56 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_45 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_89 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_8 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_100 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_111 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_177 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_188 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_133 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_122 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_199 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_144 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_155 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_166 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_8 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_168 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_157 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_179 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_102 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_113 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_135 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_146 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_124 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_68 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_79 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_24 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_13 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_35 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_57 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_46 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_9 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_156 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_145 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_101 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_112 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_123 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_178 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_134 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_189 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_167 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_9 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_103 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_114 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_136 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_147 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_125 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_169 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_158 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_14 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_69 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_25 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_58 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_36 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_47 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_157 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_168 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_146 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_113 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_102 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_135 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_124 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_179 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_104 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_115 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_137 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_148 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_126 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_159 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_15 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_26 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_59 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_37 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_48 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_158 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_147 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_169 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_114 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_103 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_136 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_125 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_105 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_116 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_149 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_138 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_127 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_16 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_27 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_38 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_49 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_115 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_104 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_137 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_126 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_148 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_159 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_117 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_106 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_139 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_128 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_17 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_28 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_39 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_149 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_116 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_105 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_138 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_127 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_118 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_107 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_129 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_90 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_29 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_18 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_117 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_106 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_139 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_128 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_119 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_108 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_80 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_91 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_19 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_118 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_107 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_129 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_109 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_70 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_81 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_92 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_119 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_108 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_82 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_60 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_71 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_93 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_109 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_50 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_83 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_72 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_61 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_94 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_73 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_84 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_62 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_95 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_51 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_40 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_74 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_52 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_85 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_63 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_96 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_30 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_41 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_230 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_75 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_20 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_64 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_86 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_53 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_31 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_42 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_97 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_220 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_231 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_230 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_65 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_76 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_10 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_54 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_21 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_87 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_32 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_43 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_98 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_221 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_232 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_210 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_231 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_220 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_66 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_77 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_11 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_22 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_88 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_44 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_99 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_33 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_55 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_222 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_233 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_200 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_211 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_232 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_221 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_210 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_67 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_12 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_23 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_56 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_78 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_89 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_45 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_34 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_212 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_234 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_223 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_201 vss vdd VSUBS mim_cap_30_30
C0 vss vdd 0.196596p
C1 vdd VSUBS 4.633771p
C2 vss VSUBS 2.2518p
.ends

.subckt cap_mim_2p0fF_DMYL6H m4_n114303_n17580# m4_n114183_n17460# VSUBS
X0 m4_n114183_n17460# m4_n114303_n17580# cap_mim_2f0fF c_width=100u c_length=100u
C0 m4_n114183_n17460# m4_n114303_n17580# 8.5013f
C1 m4_n114183_n17460# VSUBS 85.381996f
C2 m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS cap_mim_2p0fF_DMYL6H
C0 cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt cap_mim_2p0fF_RCWXT2$2 m4_n3148_n3000# m4_n3268_n3120# VSUBS
X0 m4_n3148_n3000# m4_n3268_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3148_n3000# m4_n3268_n3120# 2.57661f
C1 m4_n3148_n3000# VSUBS 9.60519f
C2 m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30$1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_DMYL6H$1 m4_93823_n2660# m4_93943_n2540# VSUBS
X0 m4_93943_n2540# m4_93823_n2660# cap_mim_2f0fF c_width=100u c_length=100u
C0 m4_93943_n2540# m4_93823_n2660# 8.5013f
C1 m4_93943_n2540# VSUBS 85.381996f
C2 m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100$1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS cap_mim_2p0fF_DMYL6H$1
C0 cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap2 vdd vss VSUBS
Xmim_cap_100_100_0 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_1 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_2 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_20 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_0 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_3 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_21 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_22 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_1 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_10 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_11 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_4 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_23 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_2 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_12 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_24 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_3 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_13 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_4 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_14 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_5 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_6 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_15 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_16 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_7 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_8 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_17 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_9 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_18 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_19 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100$1_0 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_1 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_2 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_3 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_4 vss vdd VSUBS mim_cap_100_100$1
C0 vss vdd 0.263674p
C1 vdd VSUBS 1.472734p
C2 vss VSUBS 0.649945p
.ends

.subckt mim_cap_boss vss vdd VSUBS
Xmim_cap1_0 vss vdd VSUBS mim_cap1
Xmim_cap2_0 vdd vss VSUBS mim_cap2
C0 vdd vss 1.238065p
C1 vdd VSUBS 6.099724p
C2 vss VSUBS 3.300812p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VNW VPW VDD VSS a_36_472# a_572_375# a_124_375#
+ a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 a_124_375# a_572_375# 0.012222f
C1 a_36_472# VSS 0.151218f
C2 a_124_375# a_36_472# 0.285629f
C3 a_124_375# VSS 0.136476f
C4 a_484_472# VDD 0.179463f
C5 a_484_472# VNW 0.024396f
C6 VDD a_572_375# 0.129266f
C7 VNW a_572_375# 0.18122f
C8 a_36_472# VDD 0.093681f
C9 a_36_472# VNW 0.025611f
C10 VDD VSS 0.013184f
C11 VNW VSS 0.008822f
C12 a_124_375# VDD 0.12673f
C13 a_124_375# VNW 0.180172f
C14 a_484_472# a_572_375# 0.285629f
C15 a_484_472# a_36_472# 0.013276f
C16 a_484_472# VSS 0.148682f
C17 a_484_472# a_124_375# 0.086742f
C18 VDD VNW 0.11314f
C19 a_572_375# VSS 0.082563f
C20 VSS VSUBS 0.360066f
C21 VDD VSUBS 0.286281f
C22 VNW VSUBS 1.65967f
C23 a_484_472# VSUBS 0.345058f
C24 a_36_472# VSUBS 0.404746f
C25 a_572_375# VSUBS 0.232991f
C26 a_124_375# VSUBS 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VNW VPW VSS I VDD VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 I VDD 0.017439f
C1 VNW VDD 0.048519f
C2 I VNW 0.027206f
C3 VSS VDD 0.009725f
C4 I VSS 0.031625f
C5 VSS VNW 0.007461f
C6 VSS VSUBS 0.12617f
C7 VDD VSUBS 0.087026f
C8 I VSUBS 0.139667f
C9 VNW VSUBS 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VNW VPW VDD VSS ZN A1 A2 a_224_472# VSUBS
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 VNW VDD 0.093678f
C1 VNW A2 0.128798f
C2 a_224_472# VDD 0.013964f
C3 a_224_472# A2 0.008979f
C4 VSS VDD 0.023219f
C5 VSS A2 0.043352f
C6 VNW VSS 0.010571f
C7 A1 ZN 0.579732f
C8 A1 VDD 0.028041f
C9 A1 A2 0.037814f
C10 VNW A1 0.136915f
C11 ZN VDD 0.117921f
C12 ZN A2 0.378409f
C13 VNW ZN 0.019783f
C14 VSS A1 0.168633f
C15 a_224_472# ZN 0.023693f
C16 VSS ZN 0.08687f
C17 VDD A2 0.255318f
C18 VSS VSUBS 0.331491f
C19 ZN VSUBS 0.058886f
C20 VDD VSUBS 0.218051f
C21 A1 VSUBS 0.331856f
C22 A2 VSUBS 0.334514f
C23 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 VNW VPW D Q RN VSS CLK VDD a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_1456_156#
+ a_1288_156# a_2248_156# a_2560_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 a_36_151# a_2560_156# 0.003674f
C1 VSS VDD 0.01338f
C2 VDD a_1204_472# 0.282626f
C3 VNW a_2560_156# 0.020165f
C4 Q VDD 0.149344f
C5 CLK VDD 0.02303f
C6 VSS a_2665_112# 0.184997f
C7 RN VSS 0.441968f
C8 VDD a_36_151# 0.417088f
C9 RN a_1204_472# 0.021039f
C10 a_1000_472# VSS 0.04356f
C11 VNW VDD 0.503557f
C12 a_1000_472# a_1204_472# 0.66083f
C13 a_2248_156# VSS 0.030473f
C14 Q a_2665_112# 0.109436f
C15 VDD a_1308_423# 0.094185f
C16 a_448_472# a_1456_156# 0.00227f
C17 a_2248_156# Q 0.014355f
C18 D a_448_472# 0.328788f
C19 a_1000_472# a_796_472# 0.048436f
C20 a_36_151# a_2665_112# 0.019043f
C21 RN a_36_151# 0.080102f
C22 a_3041_156# a_2665_112# 0.001774f
C23 VNW a_2665_112# 0.354715f
C24 RN a_3041_156# 0.01068f
C25 a_1000_472# a_36_151# 0.08126f
C26 VNW RN 0.329494f
C27 a_1288_156# a_448_472# 0.002067f
C28 a_2248_156# a_36_151# 0.042802f
C29 VNW a_1000_472# 0.241357f
C30 RN a_1308_423# 0.079294f
C31 VDD a_2560_156# 0.00217f
C32 VNW a_2248_156# 0.212431f
C33 a_1000_472# a_1308_423# 0.934191f
C34 a_2248_156# a_1308_423# 0.056721f
C35 a_448_472# VSS 1.20207f
C36 a_448_472# a_1204_472# 0.008996f
C37 a_2560_156# a_2665_112# 0.116059f
C38 VSS a_1456_156# 0.001901f
C39 RN a_2560_156# 0.038779f
C40 D VSS 0.064618f
C41 a_448_472# a_796_472# 0.401636f
C42 a_2248_156# a_2560_156# 0.119687f
C43 a_448_472# CLK 0.002757f
C44 a_1288_156# VSS 0.001702f
C45 a_448_472# a_36_151# 0.536965f
C46 VNW a_448_472# 0.341284f
C47 D a_796_472# 0.082858f
C48 VDD a_2665_112# 0.102046f
C49 RN VDD 0.034984f
C50 a_448_472# a_1308_423# 0.882105f
C51 D a_36_151# 0.094113f
C52 a_1000_472# VDD 0.119211f
C53 a_2248_156# VDD 1.11667f
C54 VNW D 0.128231f
C55 Q VSS 0.113401f
C56 RN a_2665_112# 0.336469f
C57 a_448_472# a_2560_156# 0.277491f
C58 VSS a_796_472# 0.05215f
C59 CLK VSS 0.021952f
C60 a_1000_472# RN 0.0832f
C61 a_2248_156# a_2665_112# 0.633318f
C62 VSS a_36_151# 0.291264f
C63 a_2248_156# RN 0.094336f
C64 a_1204_472# a_36_151# 0.006996f
C65 a_1000_472# a_2248_156# 0.001232f
C66 VNW VSS 0.010602f
C67 VNW a_1204_472# 0.016269f
C68 VSS a_1308_423# 0.013866f
C69 a_1204_472# a_1308_423# 0.026665f
C70 VNW Q 0.034443f
C71 a_796_472# a_36_151# 0.011851f
C72 a_448_472# VDD 0.456269f
C73 CLK a_36_151# 0.669598f
C74 VNW a_796_472# 0.010232f
C75 VNW CLK 0.137037f
C76 VNW a_36_151# 1.28833f
C77 D VDD 0.009367f
C78 VSS a_2560_156# 0.128503f
C79 a_1308_423# a_36_151# 0.05539f
C80 a_448_472# a_2665_112# 0.020455f
C81 VNW a_1308_423# 0.149014f
C82 a_448_472# RN 0.078731f
C83 a_1000_472# a_448_472# 0.361958f
C84 a_2248_156# a_448_472# 0.510371f
C85 Q VSUBS 0.114762f
C86 VSS VSUBS 1.26186f
C87 RN VSUBS 1.36673f
C88 D VSUBS 0.253406f
C89 VDD VSUBS 0.79945f
C90 CLK VSUBS 0.291241f
C91 VNW VSUBS 6.1377f
C92 a_2560_156# VSUBS 0.016968f
C93 a_2665_112# VSUBS 0.62251f
C94 a_2248_156# VSUBS 0.371662f
C95 a_1204_472# VSUBS 0.012971f
C96 a_1000_472# VSUBS 0.291735f
C97 a_796_472# VSUBS 0.023206f
C98 a_1308_423# VSUBS 0.279043f
C99 a_448_472# VSUBS 0.684413f
C100 a_36_151# VSUBS 1.43589f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 VNW VPW A2 B1 B2 VDD VSS ZN A1 a_36_68# a_244_472#
+ a_692_472# VSUBS
X0 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 a_692_472# ZN 0.011665f
C1 VDD a_244_472# 0.00636f
C2 B1 VNW 0.125926f
C3 a_36_68# ZN 0.419486f
C4 ZN A2 0.390894f
C5 VDD VSS 0.011512f
C6 B1 B2 0.036483f
C7 VNW ZN 0.010694f
C8 VSS A1 0.084232f
C9 a_36_68# a_244_472# 0.027448f
C10 VSS a_36_68# 0.392965f
C11 B1 ZN 0.079f
C12 VSS A2 0.087422f
C13 a_244_472# B2 0.002003f
C14 VSS VNW 0.010714f
C15 B1 a_244_472# 0.003598f
C16 VSS B2 0.025295f
C17 VDD A1 0.014671f
C18 VDD a_692_472# 0.004194f
C19 B1 VSS 0.025138f
C20 VDD a_36_68# 0.787847f
C21 VDD A2 0.019572f
C22 VSS ZN 0.085273f
C23 VDD VNW 0.139306f
C24 a_36_68# A1 0.160084f
C25 A1 A2 0.038725f
C26 a_36_68# a_692_472# 0.015646f
C27 VDD B2 0.246452f
C28 a_36_68# A2 0.340509f
C29 VNW A1 0.115376f
C30 VDD B1 0.014643f
C31 VNW a_36_68# 0.040298f
C32 VNW A2 0.125671f
C33 B1 A1 0.163724f
C34 VDD ZN 0.004634f
C35 a_36_68# B2 0.369561f
C36 B1 a_36_68# 0.437534f
C37 VNW B2 0.133721f
C38 ZN A1 0.430191f
C39 VSS VSUBS 0.383233f
C40 ZN VSUBS 0.012598f
C41 VDD VSUBS 0.318857f
C42 A2 VSUBS 0.2826f
C43 A1 VSUBS 0.258579f
C44 B1 VSUBS 0.257485f
C45 B2 VSUBS 0.309037f
C46 VNW VSUBS 2.00777f
C47 a_36_68# VSUBS 0.150048f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 VNW VPW B1 B2 VDD VSS ZN A1 A2 a_49_472#
+ a_665_69# a_257_69# VSUBS
X0 ZN B1 a_257_69# VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
C0 a_49_472# B1 0.069833f
C1 ZN VNW 0.017894f
C2 a_49_472# B2 0.151151f
C3 VDD A1 0.013859f
C4 VSS B1 0.095385f
C5 VSS B2 0.06757f
C6 a_49_472# A1 0.021757f
C7 VSS a_665_69# 0.003829f
C8 VSS A1 0.087393f
C9 a_665_69# A2 0.006702f
C10 A2 A1 0.392541f
C11 a_49_472# VDD 0.887006f
C12 B1 VNW 0.109456f
C13 B2 VNW 0.129409f
C14 VDD VSS 0.00787f
C15 B1 ZN 0.367665f
C16 VDD A2 0.013575f
C17 B2 ZN 0.001886f
C18 a_49_472# VSS 0.02154f
C19 A1 VNW 0.10965f
C20 a_665_69# ZN 0.001059f
C21 a_49_472# A2 0.075759f
C22 A1 ZN 0.447732f
C23 VSS A2 0.150463f
C24 B1 a_257_69# 0.003901f
C25 B2 a_257_69# 0.003563f
C26 VDD VNW 0.112326f
C27 VDD ZN 0.004108f
C28 a_49_472# VNW 0.026629f
C29 B1 B2 0.18297f
C30 a_49_472# ZN 0.239204f
C31 VSS VNW 0.011011f
C32 A2 VNW 0.131727f
C33 VSS ZN 0.071892f
C34 B1 A1 0.041046f
C35 A2 ZN 0.102518f
C36 a_665_69# A1 0.002008f
C37 VDD B1 0.017923f
C38 VSS a_257_69# 0.00576f
C39 VDD B2 0.026097f
C40 VSS VSUBS 0.39457f
C41 ZN VSUBS 0.021794f
C42 VDD VSUBS 0.243433f
C43 A2 VSUBS 0.322629f
C44 A1 VSUBS 0.250967f
C45 B1 VSUBS 0.261124f
C46 B2 VSUBS 0.322244f
C47 VNW VSUBS 1.83372f
C48 a_49_472# VSUBS 0.054843f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VNW VPW VSS Z I VDD a_36_160# VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 a_36_160# VSS 0.074156f
C1 VDD VSS 0.009574f
C2 Z VNW 0.030347f
C3 I VSS 0.12329f
C4 VDD a_36_160# 0.2736f
C5 a_36_160# I 0.545454f
C6 VDD I 0.02612f
C7 VSS VNW 0.009324f
C8 a_36_160# VNW 0.170864f
C9 VDD VNW 0.087464f
C10 VSS Z 0.146199f
C11 I VNW 0.2276f
C12 a_36_160# Z 0.281838f
C13 VDD Z 0.128274f
C14 I Z 0.041707f
C15 VSS VSUBS 0.28275f
C16 Z VSUBS 0.10469f
C17 VDD VSUBS 0.178615f
C18 I VSUBS 0.323491f
C19 VNW VSUBS 1.31158f
C20 a_36_160# VSUBS 0.386641f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VNW VPW VDD VSS I ZN VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VNW ZN 0.031181f
C1 VNW VDD 0.076212f
C2 ZN VDD 0.098026f
C3 VNW VSS 0.011085f
C4 VSS ZN 0.077008f
C5 VNW I 0.135368f
C6 VSS VDD 0.025441f
C7 ZN I 0.47009f
C8 VDD I 0.157124f
C9 VSS I 0.058937f
C10 VSS VSUBS 0.242183f
C11 ZN VSUBS 0.095505f
C12 VDD VSUBS 0.182097f
C13 I VSUBS 0.355642f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VNW VPW VSS ZN I VDD VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VNW ZN 0.022202f
C1 VNW VDD 0.076257f
C2 ZN VDD 0.137375f
C3 VNW VSS 0.011339f
C4 VSS ZN 0.115297f
C5 VNW I 0.137757f
C6 VSS VDD 0.025626f
C7 ZN I 0.262199f
C8 VDD I 0.041847f
C9 VSS I 0.0533f
C10 VSS VSUBS 0.2316f
C11 ZN VSUBS 0.113404f
C12 VDD VSUBS 0.181139f
C13 I VSUBS 0.341982f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VNW VPW VDD VSS a_36_472# a_124_375# VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 a_124_375# VDD 0.126034f
C1 a_124_375# VNW 0.179924f
C2 VDD VNW 0.061035f
C3 a_124_375# VSS 0.082879f
C4 VSS VDD 0.006592f
C5 a_124_375# a_36_472# 0.285629f
C6 VSS VNW 0.004411f
C7 VDD a_36_472# 0.093681f
C8 VNW a_36_472# 0.025989f
C9 VSS a_36_472# 0.150876f
C10 VSS VSUBS 0.218985f
C11 VDD VSUBS 0.182777f
C12 VNW VSUBS 0.96348f
C13 a_36_472# VSUBS 0.417394f
C14 a_124_375# VSUBS 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 VNW VPW Z I VDD VSS a_224_472# VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 Z VSS 0.70427f
C1 a_224_472# VDD 0.74621f
C2 VSS VNW 0.01282f
C3 a_224_472# I 0.796069f
C4 VDD I 0.1311f
C5 a_224_472# Z 2.29481f
C6 Z VDD 0.819024f
C7 a_224_472# VNW 1.14633f
C8 Z I 0.001907f
C9 VDD VNW 0.305516f
C10 a_224_472# VSS 0.659695f
C11 I VNW 0.55539f
C12 VSS VDD 0.031131f
C13 VSS I 0.158668f
C14 Z VNW 0.038011f
C15 VSS VSUBS 0.910368f
C16 Z VSUBS 0.18914f
C17 VDD VSUBS 0.724491f
C18 I VSUBS 1.16773f
C19 VNW VSUBS 4.79254f
C20 a_224_472# VSUBS 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 VNW VPW B VDD VSS ZN A1 A2 a_36_472# a_244_68#
+ VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VSUBS nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
C0 VSS a_244_68# 0.00255f
C1 ZN B 0.00761f
C2 VSS VNW 0.009145f
C3 a_36_472# B 0.01027f
C4 ZN a_36_472# 0.088503f
C5 ZN A2 0.248411f
C6 A2 a_36_472# 0.10395f
C7 ZN A1 0.245346f
C8 A1 B 0.157699f
C9 A1 a_36_472# 0.104556f
C10 A1 A2 0.047589f
C11 VSS B 0.080416f
C12 ZN VSS 0.304078f
C13 VSS a_36_472# 0.004325f
C14 VNW VDD 0.11216f
C15 VSS A2 0.069479f
C16 A1 VSS 0.021732f
C17 VDD B 0.071777f
C18 ZN VDD 0.003129f
C19 ZN a_244_68# 0.008784f
C20 a_36_472# VDD 0.581285f
C21 VNW B 0.137038f
C22 ZN VNW 0.014655f
C23 A2 VDD 0.015143f
C24 a_36_472# VNW 0.013943f
C25 A2 VNW 0.128282f
C26 A1 VDD 0.0167f
C27 A1 VNW 0.122087f
C28 VSS VDD 0.01275f
C29 VSS VSUBS 0.361309f
C30 VDD VSUBS 0.259458f
C31 ZN VSUBS 0.040013f
C32 B VSUBS 0.378232f
C33 A1 VSUBS 0.264815f
C34 A2 VSUBS 0.3189f
C35 VNW VSUBS 1.65967f
C36 a_36_472# VSUBS 0.031137f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VNW VPW VSS Z I VDD a_36_113# VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VDD Z 0.085355f
C1 VDD VNW 0.088196f
C2 I VSS 0.070302f
C3 a_36_113# VSS 0.11114f
C4 VSS Z 0.136942f
C5 I a_36_113# 0.476912f
C6 VNW VSS 0.009307f
C7 VDD VSS 0.009561f
C8 I Z 0.031362f
C9 VNW I 0.152645f
C10 VDD I 0.028968f
C11 a_36_113# Z 0.191876f
C12 VNW a_36_113# 0.160792f
C13 VDD a_36_113# 0.278283f
C14 VNW Z 0.030118f
C15 VSS VSUBS 0.283681f
C16 Z VSUBS 0.117185f
C17 VDD VSUBS 0.180237f
C18 I VSUBS 0.336876f
C19 VNW VSUBS 1.31158f
C20 a_36_113# VSUBS 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VNW VPW VDD VSS a_1916_375# a_1380_472#
+ a_3260_375# a_36_472# a_932_472# a_2812_375# a_2276_472# a_1828_472# a_3172_472#
+ a_572_375# a_2724_472# a_124_375# a_1468_375# a_1020_375# a_484_472# a_2364_375#
+ VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_3260_375# a_3172_472# 0.285629f
C1 a_1380_472# VSS 0.142721f
C2 VNW a_3260_375# 0.18122f
C3 a_2276_472# VDD 0.179463f
C4 a_1468_375# a_1020_375# 0.013103f
C5 a_1020_375# a_572_375# 0.013103f
C6 VSS a_3260_375# 0.081304f
C7 a_2276_472# a_1828_472# 0.013276f
C8 a_1468_375# a_1916_375# 0.013103f
C9 a_2724_472# a_2364_375# 0.087174f
C10 a_1380_472# VDD 0.179463f
C11 a_484_472# a_36_472# 0.013276f
C12 a_2724_472# a_3172_472# 0.013276f
C13 VNW a_2724_472# 0.024018f
C14 a_484_472# a_572_375# 0.285629f
C15 VNW a_36_472# 0.025611f
C16 a_3260_375# VDD 0.129266f
C17 a_2364_375# a_2812_375# 0.013103f
C18 a_1380_472# a_1828_472# 0.013276f
C19 a_2724_472# VSS 0.142721f
C20 a_1468_375# VNW 0.181468f
C21 a_2812_375# a_3172_472# 0.087174f
C22 VNW a_572_375# 0.181468f
C23 VSS a_36_472# 0.142026f
C24 VNW a_2812_375# 0.181468f
C25 a_1380_472# a_932_472# 0.013276f
C26 a_1468_375# VSS 0.131736f
C27 VSS a_572_375# 0.131736f
C28 VSS a_2812_375# 0.131736f
C29 a_1916_375# a_2364_375# 0.013103f
C30 VNW a_1020_375# 0.181468f
C31 a_2724_472# VDD 0.179463f
C32 a_1916_375# VNW 0.181468f
C33 VSS a_1020_375# 0.131736f
C34 VDD a_36_472# 0.093681f
C35 a_1916_375# VSS 0.131736f
C36 a_1468_375# VDD 0.129962f
C37 VDD a_572_375# 0.129962f
C38 a_2812_375# VDD 0.129962f
C39 a_484_472# VNW 0.024018f
C40 VNW a_2364_375# 0.181468f
C41 a_124_375# a_36_472# 0.285629f
C42 a_1468_375# a_1828_472# 0.087174f
C43 VNW a_3172_472# 0.024396f
C44 a_2276_472# a_2724_472# 0.013276f
C45 a_484_472# VSS 0.142721f
C46 a_2364_375# VSS 0.131736f
C47 VDD a_1020_375# 0.129962f
C48 a_124_375# a_572_375# 0.013103f
C49 VSS a_3172_472# 0.139489f
C50 a_1916_375# VDD 0.129962f
C51 a_932_472# a_572_375# 0.087174f
C52 VNW VSS 0.035286f
C53 a_1916_375# a_1828_472# 0.285629f
C54 a_932_472# a_1020_375# 0.285629f
C55 a_484_472# VDD 0.179463f
C56 a_2364_375# VDD 0.129962f
C57 VDD a_3172_472# 0.179463f
C58 VNW VDD 0.425768f
C59 a_1916_375# a_2276_472# 0.087174f
C60 a_1380_472# a_1468_375# 0.285629f
C61 a_484_472# a_124_375# 0.087174f
C62 VSS VDD 0.052737f
C63 VNW a_1828_472# 0.024018f
C64 a_484_472# a_932_472# 0.013276f
C65 a_3260_375# a_2812_375# 0.013103f
C66 a_1380_472# a_1020_375# 0.087174f
C67 VNW a_124_375# 0.180172f
C68 a_2276_472# a_2364_375# 0.285629f
C69 a_1828_472# VSS 0.142721f
C70 VNW a_932_472# 0.024018f
C71 a_124_375# VSS 0.131736f
C72 a_2276_472# VNW 0.024018f
C73 a_932_472# VSS 0.142721f
C74 a_2276_472# VSS 0.142721f
C75 a_2724_472# a_2812_375# 0.285629f
C76 a_1828_472# VDD 0.179463f
C77 a_1380_472# VNW 0.024018f
C78 a_124_375# VDD 0.12673f
C79 a_932_472# VDD 0.179463f
C80 VSS VSUBS 1.20585f
C81 VDD VSUBS 0.907304f
C82 VNW VSUBS 5.83682f
C83 a_3172_472# VSUBS 0.345058f
C84 a_2724_472# VSUBS 0.33241f
C85 a_2276_472# VSUBS 0.33241f
C86 a_1828_472# VSUBS 0.33241f
C87 a_1380_472# VSUBS 0.33241f
C88 a_932_472# VSUBS 0.33241f
C89 a_484_472# VSUBS 0.33241f
C90 a_36_472# VSUBS 0.404746f
C91 a_3260_375# VSUBS 0.233093f
C92 a_2812_375# VSUBS 0.17167f
C93 a_2364_375# VSUBS 0.17167f
C94 a_1916_375# VSUBS 0.17167f
C95 a_1468_375# VSUBS 0.17167f
C96 a_1020_375# VSUBS 0.17167f
C97 a_572_375# VSUBS 0.17167f
C98 a_124_375# VSUBS 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 VNW VPW A3 VDD VSS ZN A1 A2 a_455_68# a_271_68#
+ VSUBS
X0 ZN A1 a_455_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 A2 VSS 0.104901f
C1 A2 a_455_68# 0.005127f
C2 A3 VNW 0.148237f
C3 a_271_68# ZN 0.001916f
C4 A3 VSS 0.07804f
C5 VNW ZN 0.034322f
C6 VSS ZN 0.064021f
C7 VNW VDD 0.112537f
C8 VSS VDD 0.008734f
C9 ZN a_455_68# 0.002926f
C10 A1 VNW 0.12917f
C11 A1 VSS 0.084906f
C12 A1 a_455_68# 0.004981f
C13 A2 A3 0.117566f
C14 A2 ZN 0.078589f
C15 a_271_68# VSS 0.006038f
C16 A2 VDD 0.023177f
C17 VSS VNW 0.008577f
C18 A3 ZN 0.008403f
C19 A1 A2 0.133044f
C20 A3 VDD 0.079999f
C21 VSS a_455_68# 0.006909f
C22 VDD ZN 0.33173f
C23 A2 a_271_68# 0.004027f
C24 A1 ZN 0.384588f
C25 A2 VNW 0.121191f
C26 A1 VDD 0.022021f
C27 VSS VSUBS 0.307914f
C28 ZN VSUBS 0.133449f
C29 VDD VSUBS 0.241872f
C30 A1 VSUBS 0.287469f
C31 A2 VSUBS 0.25736f
C32 A3 VSUBS 0.326833f
C33 VNW VSUBS 1.48562f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VNW VPW VDD VSS ZN A1 A2 a_245_68# VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
C0 A1 VDD 0.027485f
C1 A2 VNW 0.125396f
C2 VSS ZN 0.098328f
C3 A2 A1 0.226398f
C4 A1 VNW 0.119756f
C5 VSS VDD 0.017706f
C6 ZN VDD 0.240333f
C7 A1 a_245_68# 0.008831f
C8 A2 VSS 0.051087f
C9 VSS VNW 0.006174f
C10 A2 ZN 0.038658f
C11 ZN VNW 0.02653f
C12 VSS A1 0.131667f
C13 ZN A1 0.351362f
C14 A2 VDD 0.039698f
C15 VDD VNW 0.084263f
C16 VSS a_245_68# 0.002295f
C17 VSS VSUBS 0.238729f
C18 ZN VSUBS 0.105772f
C19 VDD VSUBS 0.243067f
C20 A1 VSUBS 0.290957f
C21 A2 VSUBS 0.314823f
C22 VNW VSUBS 1.13753f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VNW VPW VDD VSS Z A1 A2 a_255_603# a_67_603#
+ VSUBS
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 Z a_67_603# 0.181586f
C1 A1 a_67_603# 0.540888f
C2 A2 Z 0.027598f
C3 A1 A2 0.062395f
C4 VNW a_67_603# 0.157241f
C5 VNW A2 0.216313f
C6 VSS a_67_603# 0.250493f
C7 VDD a_67_603# 0.307039f
C8 a_67_603# a_255_603# 0.007617f
C9 A2 VSS 0.025748f
C10 A2 VDD 0.147628f
C11 A2 a_255_603# 0.001961f
C12 VNW Z 0.033884f
C13 A1 VNW 0.220003f
C14 Z VSS 0.158265f
C15 VDD Z 0.196046f
C16 A1 VSS 0.050738f
C17 A1 VDD 0.01431f
C18 VNW VSS 0.010039f
C19 VNW VDD 0.11771f
C20 VDD VSS 0.008648f
C21 VDD a_255_603# 0.005359f
C22 A2 a_67_603# 0.505374f
C23 VSS VSUBS 0.359722f
C24 Z VSUBS 0.102754f
C25 VDD VSUBS 0.233025f
C26 A2 VSUBS 0.313441f
C27 A1 VSUBS 0.39469f
C28 VNW VSUBS 1.65967f
C29 a_67_603# VSUBS 0.345683f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 VNW VPW B C VDD VSS ZN A1 A2 a_36_68# a_1612_497#
+ a_2124_68# a_244_497# a_2960_68# a_3368_68# a_2552_68# a_1164_497# a_716_497# VSUBS
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
C0 ZN a_36_68# 1.98502f
C1 B C 1.73339f
C2 C VDD 0.095093f
C3 ZN a_244_497# 0.009475f
C4 VSS B 0.072527f
C5 VSS VDD 0.005699f
C6 VNW B 0.600992f
C7 VNW VDD 0.366897f
C8 VSS A2 0.060501f
C9 a_36_68# a_2124_68# 0.012118f
C10 VSS A1 0.060963f
C11 VNW A2 0.590323f
C12 VSS a_2552_68# 0.002422f
C13 VNW A1 0.51833f
C14 ZN B 0.426118f
C15 ZN VDD 2.06829f
C16 ZN a_1164_497# 0.021094f
C17 ZN A2 1.2828f
C18 a_716_497# VDD 0.008599f
C19 ZN A1 1.37575f
C20 a_2960_68# VSS 0.002422f
C21 VSS a_3368_68# 0.004815f
C22 a_716_497# A2 0.00653f
C23 ZN a_1612_497# 0.024559f
C24 a_36_68# B 1.37417f
C25 a_36_68# VDD 0.021485f
C26 a_244_497# VDD 0.020528f
C27 A2 a_36_68# 0.108262f
C28 a_244_497# A2 0.01347f
C29 a_36_68# A1 0.065645f
C30 a_36_68# a_2552_68# 0.009506f
C31 B VDD 0.100578f
C32 a_1164_497# VDD 0.008664f
C33 VSS C 0.092809f
C34 a_2960_68# a_36_68# 0.009506f
C35 A2 B 0.037299f
C36 a_3368_68# a_36_68# 0.007478f
C37 A2 VDD 0.15752f
C38 VNW C 0.636287f
C39 a_1164_497# A2 0.009095f
C40 A1 VDD 0.078657f
C41 VSS VNW 0.004483f
C42 B a_2552_68# 0.002588f
C43 A2 A1 1.73987f
C44 a_1612_497# VDD 0.009792f
C45 ZN C 0.514613f
C46 ZN VSS 0.006216f
C47 A2 a_1612_497# 0.010709f
C48 a_2960_68# B 0.002626f
C49 ZN VNW 0.056895f
C50 VSS a_2124_68# 0.004133f
C51 a_36_68# C 0.105844f
C52 a_716_497# ZN 0.027752f
C53 VSS a_36_68# 3.64719f
C54 VNW a_36_68# 0.004654f
C55 VSS VSUBS 1.08055f
C56 ZN VSUBS 0.051826f
C57 VDD VSUBS 0.846798f
C58 C VSUBS 1.06351f
C59 B VSUBS 1.11555f
C60 A1 VSUBS 1.1956f
C61 A2 VSUBS 1.16629f
C62 VNW VSUBS 5.892971f
C63 a_36_68# VSUBS 0.063181f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 VNW VPW Z VSS VDD I a_36_160# VSUBS
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VSUBS nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VSUBS nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
C0 VNW VSS 0.00834f
C1 VNW a_36_160# 0.302514f
C2 Z VSS 0.111496f
C3 a_36_160# Z 0.426617f
C4 VNW VDD 0.111398f
C5 Z VDD 0.161733f
C6 I VSS 0.178818f
C7 I a_36_160# 0.564508f
C8 VNW Z 0.021185f
C9 a_36_160# VSS 0.114407f
C10 I VDD 0.028233f
C11 I VNW 0.1633f
C12 I Z 0.016176f
C13 VSS VDD 0.01316f
C14 a_36_160# VDD 0.31851f
C15 VSS VSUBS 0.397291f
C16 Z VSUBS 0.097163f
C17 VDD VSUBS 0.238155f
C18 I VSUBS 0.333888f
C19 VNW VSUBS 1.65967f
C20 a_36_160# VSUBS 0.696445f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VNW VPW VDD VSS a_1380_472# a_36_472#
+ a_932_472# a_572_375# a_124_375# a_1468_375# a_1020_375# a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 VSS a_1468_375# 0.082091f
C1 a_36_472# a_124_375# 0.285629f
C2 VNW a_124_375# 0.180172f
C3 VNW a_932_472# 0.024018f
C4 VDD a_124_375# 0.12673f
C5 VDD a_932_472# 0.179463f
C6 a_1380_472# a_1020_375# 0.086905f
C7 VNW a_1468_375# 0.18122f
C8 a_572_375# a_124_375# 0.012552f
C9 VDD a_1468_375# 0.129266f
C10 a_572_375# a_932_472# 0.086905f
C11 a_36_472# VSS 0.147381f
C12 VNW VSS 0.017643f
C13 VDD VSS 0.026369f
C14 a_572_375# VSS 0.134699f
C15 a_36_472# VNW 0.025611f
C16 a_36_472# VDD 0.093681f
C17 a_1380_472# a_932_472# 0.013276f
C18 VNW VDD 0.217349f
C19 a_1380_472# a_1468_375# 0.285629f
C20 a_572_375# VNW 0.181468f
C21 a_572_375# VDD 0.129962f
C22 a_1380_472# VSS 0.144845f
C23 a_484_472# a_124_375# 0.086905f
C24 a_484_472# a_932_472# 0.013276f
C25 VNW a_1380_472# 0.024396f
C26 a_1380_472# VDD 0.179463f
C27 VSS a_484_472# 0.148077f
C28 a_36_472# a_484_472# 0.013276f
C29 VNW a_484_472# 0.024018f
C30 VDD a_484_472# 0.179463f
C31 a_572_375# a_484_472# 0.285629f
C32 a_1020_375# a_932_472# 0.285629f
C33 a_1468_375# a_1020_375# 0.012552f
C34 VSS a_1020_375# 0.134699f
C35 VNW a_1020_375# 0.181468f
C36 VDD a_1020_375# 0.129962f
C37 a_572_375# a_1020_375# 0.012552f
C38 VSS a_124_375# 0.134699f
C39 VSS a_932_472# 0.148077f
C40 VSS VSUBS 0.642184f
C41 VDD VSUBS 0.493288f
C42 VNW VSUBS 3.05206f
C43 a_1380_472# VSUBS 0.345058f
C44 a_932_472# VSUBS 0.33241f
C45 a_484_472# VSUBS 0.33241f
C46 a_36_472# VSUBS 0.404746f
C47 a_1468_375# VSUBS 0.233029f
C48 a_1020_375# VSUBS 0.171606f
C49 a_572_375# VSUBS 0.171606f
C50 a_124_375# VSUBS 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VNW VPW VSS Z I VDD a_36_68# VSUBS
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VSUBS nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 a_36_68# VSS 0.156367f
C1 VDD I 0.029139f
C2 a_36_68# Z 0.432914f
C3 VNW VSS 0.009972f
C4 VNW Z 0.023138f
C5 VDD a_36_68# 0.271105f
C6 VDD VNW 0.114912f
C7 a_36_68# I 0.731677f
C8 VNW I 0.133333f
C9 a_36_68# VNW 0.296832f
C10 VSS Z 0.133443f
C11 VDD VSS 0.014283f
C12 VDD Z 0.172592f
C13 VSS I 0.128735f
C14 I Z 0.018906f
C15 VSS VSUBS 0.338876f
C16 Z VSUBS 0.103236f
C17 VDD VSUBS 0.234026f
C18 I VSUBS 0.298844f
C19 VNW VSUBS 1.65967f
C20 a_36_68# VSUBS 0.69549f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 VNW VPW S VDD VSS Z I0 I1 a_848_380# a_1084_68#
+ a_124_24# a_1152_472# a_692_472# VSUBS
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VSUBS nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VSUBS nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
C0 S a_848_380# 0.754833f
C1 a_692_68# VSS 0.001982f
C2 a_124_24# VNW 0.277682f
C3 I1 a_692_472# 0.001219f
C4 a_1084_68# S 0.001644f
C5 a_124_24# VDD 0.309232f
C6 a_124_24# a_1152_472# 0.00128f
C7 VDD VNW 0.182986f
C8 S I1 0.042269f
C9 I0 a_124_24# 0.004772f
C10 VSS a_124_24# 0.501844f
C11 I0 VNW 0.103064f
C12 a_124_24# Z 0.219295f
C13 S a_692_472# 0.002582f
C14 VSS VNW 0.009598f
C15 VDD a_1152_472# 0.00645f
C16 VNW Z 0.020389f
C17 I0 VDD 0.028914f
C18 a_124_24# a_848_380# 0.302602f
C19 VSS VDD 0.028952f
C20 VNW a_848_380# 0.174516f
C21 VDD Z 0.20273f
C22 I0 VSS 0.124513f
C23 a_1084_68# a_124_24# 0.002839f
C24 VDD a_848_380# 0.319708f
C25 VSS Z 0.129676f
C26 a_848_380# a_1152_472# 0.007362f
C27 a_124_24# I1 0.564972f
C28 I0 a_848_380# 0.082224f
C29 VNW I1 0.127749f
C30 VSS a_848_380# 0.130064f
C31 a_124_24# a_692_472# 0.033243f
C32 I0 a_1084_68# 0.00492f
C33 VDD I1 0.227359f
C34 a_1084_68# VSS 0.009508f
C35 S a_124_24# 0.245829f
C36 VDD a_692_472# 0.009663f
C37 S VNW 0.253706f
C38 VSS I1 0.026996f
C39 I1 Z 0.027341f
C40 S VDD 0.056165f
C41 a_692_68# a_124_24# 0.006853f
C42 I1 a_848_380# 0.013444f
C43 I0 S 0.533789f
C44 VSS S 0.081531f
C45 a_848_380# a_692_472# 0.003985f
C46 VSS VSUBS 0.565512f
C47 Z VSUBS 0.047467f
C48 VDD VSUBS 0.424967f
C49 I0 VSUBS 0.267152f
C50 S VSUBS 0.549493f
C51 I1 VSUBS 0.247562f
C52 VNW VSUBS 2.87801f
C53 a_848_380# VSUBS 0.40208f
C54 a_124_24# VSUBS 0.591898f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VNW VPW VDD B A2 ZN A1 VSS a_36_68# a_244_472#
+ VSUBS
X0 VSS B a_36_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 ZN VSS 0.088946f
C1 a_36_68# ZN 0.56857f
C2 a_244_472# VDD 0.004051f
C3 ZN A1 0.496662f
C4 VDD B 0.07579f
C5 ZN A2 0.400775f
C6 ZN VDD 0.006004f
C7 VSS VNW 0.0064f
C8 a_36_68# VNW 0.038286f
C9 a_36_68# VSS 0.117681f
C10 A1 VNW 0.117811f
C11 A1 VSS 0.090903f
C12 VNW A2 0.122386f
C13 VSS A2 0.083821f
C14 a_36_68# A1 0.292244f
C15 a_36_68# A2 0.489122f
C16 VNW VDD 0.117098f
C17 ZN a_244_472# 0.014146f
C18 VSS VDD 0.004855f
C19 A1 A2 0.038725f
C20 a_36_68# VDD 0.753239f
C21 A1 VDD 0.014914f
C22 VDD A2 0.017122f
C23 VNW B 0.163023f
C24 VSS B 0.198567f
C25 a_36_68# a_244_472# 0.013419f
C26 a_36_68# B 0.389329f
C27 ZN VNW 0.011308f
C28 A1 B 0.034707f
C29 VSS VSUBS 0.342662f
C30 ZN VSUBS 0.011384f
C31 VDD VSUBS 0.256635f
C32 B VSUBS 0.339176f
C33 A1 VSUBS 0.256004f
C34 A2 VSUBS 0.28395f
C35 VNW VSUBS 1.65967f
C36 a_36_68# VSUBS 0.112263f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 VNW VPW Z VSS VDD I a_224_552# VSUBS
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
C0 a_224_552# VDD 0.347549f
C1 a_224_552# I 0.421587f
C2 VDD Z 0.356369f
C3 Z I 0.002319f
C4 VDD VNW 0.176912f
C5 VNW I 0.376531f
C6 a_224_552# Z 1.17071f
C7 VSS VDD 0.030201f
C8 a_224_552# VNW 0.5926f
C9 VSS I 0.061715f
C10 Z VNW 0.027266f
C11 VSS a_224_552# 0.331404f
C12 VSS Z 0.275062f
C13 VDD I 0.069894f
C14 VSS VNW 0.009226f
C15 VSS VSUBS 0.628617f
C16 Z VSUBS 0.102362f
C17 VDD VSUBS 0.415149f
C18 I VSUBS 0.471574f
C19 VNW VSUBS 2.70396f
C20 a_224_552# VSUBS 1.31114f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VNW VPW VDD VSS ZN A1 A2 a_234_472# a_672_472#
+ VSUBS
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 A2 a_234_472# 0.018681f
C1 VNW VDD 0.137685f
C2 ZN a_234_472# 0.003154f
C3 A1 VDD 0.037494f
C4 VNW A1 0.25895f
C5 VDD A2 0.13595f
C6 a_672_472# VDD 0.005379f
C7 VNW A2 0.275679f
C8 A1 A2 0.636124f
C9 ZN VDD 0.517479f
C10 a_672_472# A2 0.0147f
C11 ZN VNW 0.03148f
C12 ZN A1 0.274601f
C13 VDD VSS 0.023993f
C14 VNW VSS 0.010681f
C15 A1 VSS 0.052992f
C16 ZN A2 0.509001f
C17 ZN a_672_472# 0.023475f
C18 A2 VSS 0.07211f
C19 ZN VSS 0.460527f
C20 VDD a_234_472# 0.0121f
C21 VSS VSUBS 0.451405f
C22 ZN VSUBS 0.138491f
C23 VDD VSUBS 0.322159f
C24 A1 VSUBS 0.557317f
C25 A2 VSUBS 0.617688f
C26 VNW VSUBS 2.00777f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 VNW VPW A3 VDD VSS ZN A1 A2 a_448_472# a_244_472#
+ VSUBS
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
C0 VNW ZN 0.040402f
C1 VDD A2 0.09496f
C2 VSS A2 0.027728f
C3 A1 A2 0.145555f
C4 VNW A3 0.136756f
C5 VDD a_244_472# 0.006513f
C6 a_448_472# A2 0.012315f
C7 A3 ZN 0.035547f
C8 VNW A2 0.116878f
C9 VSS VDD 0.01583f
C10 VDD A1 0.095023f
C11 VSS A1 0.025677f
C12 ZN A2 0.096665f
C13 a_448_472# VDD 0.013539f
C14 a_448_472# A1 0.012619f
C15 VDD VNW 0.11801f
C16 VSS VNW 0.008407f
C17 VNW A1 0.127941f
C18 a_244_472# ZN 0.001803f
C19 A3 A2 0.416588f
C20 a_244_472# A3 0.019089f
C21 VDD ZN 0.116419f
C22 VSS ZN 0.283414f
C23 A1 ZN 0.499849f
C24 a_448_472# ZN 0.006209f
C25 VDD A3 0.201466f
C26 VSS A3 0.058214f
C27 a_244_472# A2 0.003952f
C28 VSS VSUBS 0.367618f
C29 ZN VSUBS 0.134331f
C30 VDD VSUBS 0.264623f
C31 A1 VSUBS 0.311038f
C32 A2 VSUBS 0.285534f
C33 A3 VSUBS 0.334053f
C34 VNW VSUBS 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 VNW VPW A3 VDD VSS ZN A1 A2 a_36_68# a_1732_68#
+ a_244_68# a_1100_68# a_1528_68# a_672_68# VSUBS
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
C0 VDD A1 0.115489f
C1 a_36_68# VSS 2.77545f
C2 ZN A1 1.266f
C3 A3 A1 0.001696f
C4 VDD VSS 0.004708f
C5 VSS a_672_68# 0.003125f
C6 A3 a_1100_68# 0.003385f
C7 VSS ZN 0.00864f
C8 A3 VSS 0.09506f
C9 a_36_68# A2 0.223434f
C10 VNW A1 0.700258f
C11 VSS a_1528_68# 0.003775f
C12 VDD A2 0.124271f
C13 A2 ZN 1.77619f
C14 VNW VSS 0.003704f
C15 a_1732_68# VSS 0.002237f
C16 A3 A2 1.65768f
C17 VDD a_36_68# 0.029088f
C18 a_36_68# a_672_68# 0.012389f
C19 VSS A1 0.065524f
C20 VNW A2 0.630933f
C21 a_36_68# ZN 0.885472f
C22 a_244_68# VSS 0.006268f
C23 VSS a_1100_68# 0.003125f
C24 A3 a_36_68# 1.03106f
C25 VDD ZN 1.57207f
C26 a_36_68# a_1528_68# 0.012072f
C27 VDD A3 0.107959f
C28 A3 a_672_68# 0.003442f
C29 A2 A1 0.077487f
C30 A3 ZN 0.150755f
C31 VNW a_36_68# 0.007741f
C32 a_1732_68# a_36_68# 0.011094f
C33 VSS A2 0.070822f
C34 VNW VDD 0.292073f
C35 VNW ZN 0.095885f
C36 a_1732_68# ZN 0.002613f
C37 VNW A3 0.599629f
C38 a_36_68# A1 0.118844f
C39 a_244_68# a_36_68# 0.009768f
C40 a_36_68# a_1100_68# 0.012396f
C41 VSS VSUBS 0.861061f
C42 ZN VSUBS 0.103891f
C43 VDD VSUBS 0.701563f
C44 A1 VSUBS 1.27704f
C45 A3 VSUBS 1.11693f
C46 A2 VSUBS 1.08692f
C47 VNW VSUBS 4.73584f
C48 a_36_68# VSUBS 0.061249f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VNW VPW VDD VSS Z A1 A2 a_36_159# VSUBS
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VSUBS nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VSUBS nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
C0 a_36_159# a_244_159# 0.003343f
C1 VNW VSS 0.007925f
C2 VNW A2 0.20463f
C3 A1 VSS 0.010276f
C4 A2 A1 0.061431f
C5 a_36_159# VSS 0.244357f
C6 a_36_159# A2 0.472781f
C7 VDD Z 0.158212f
C8 VNW Z 0.032842f
C9 VDD VNW 0.125609f
C10 VDD A1 0.04397f
C11 a_36_159# Z 0.215269f
C12 a_244_159# VSS 0.001449f
C13 VDD a_36_159# 0.130189f
C14 A2 VSS 0.011099f
C15 VNW A1 0.206765f
C16 VNW a_36_159# 0.162496f
C17 a_36_159# A1 0.377122f
C18 Z VSS 0.102819f
C19 Z A2 0.020174f
C20 VDD VSS 0.014131f
C21 VDD A2 0.184025f
C22 VSS VSUBS 0.35312f
C23 Z VSUBS 0.096476f
C24 VDD VSUBS 0.251252f
C25 A2 VSUBS 0.262264f
C26 A1 VSUBS 0.321274f
C27 VNW VSUBS 1.65967f
C28 a_36_159# VSUBS 0.374116f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 VNW VPW A2 B C VDD VSS ZN A1 a_2590_472#
+ a_170_472# a_1602_69# a_786_69# a_3126_472# a_1194_69# a_3662_472# a_2034_472# a_358_69#
+ VSUBS
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VSUBS nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VSUBS nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VSUBS nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VSUBS nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
C0 VDD C 0.089678f
C1 B a_2034_472# 0.008709f
C2 VNW VSS 0.012025f
C3 ZN VDD 0.008843f
C4 ZN a_1602_69# 0.008113f
C5 a_2590_472# B 0.007345f
C6 VNW A1 0.480244f
C7 ZN A2 1.83822f
C8 ZN C 1.79111f
C9 ZN a_1194_69# 0.00847f
C10 a_358_69# VSS 0.005318f
C11 VNW VDD 0.393677f
C12 a_3126_472# a_170_472# 0.01307f
C13 VSS a_170_472# 0.00801f
C14 a_358_69# A1 0.001641f
C15 a_3662_472# VDD 0.007223f
C16 VNW A2 0.513788f
C17 a_170_472# A1 0.0698f
C18 VNW C 0.61926f
C19 a_3126_472# B 0.007345f
C20 B VSS 0.119454f
C21 ZN VNW 0.045695f
C22 B A1 0.001644f
C23 VDD a_170_472# 2.96356f
C24 A2 a_170_472# 0.109943f
C25 C a_170_472# 0.075372f
C26 VDD B 0.110239f
C27 VDD a_2034_472# 0.008673f
C28 ZN a_358_69# 0.011344f
C29 a_2590_472# VDD 0.007681f
C30 ZN a_170_472# 0.818521f
C31 A2 B 0.05388f
C32 a_786_69# VSS 0.003966f
C33 C B 1.34577f
C34 a_786_69# A1 0.001203f
C35 ZN B 0.231932f
C36 VSS A1 0.087217f
C37 VNW a_170_472# 0.018375f
C38 a_3662_472# a_170_472# 0.013628f
C39 a_3126_472# VDD 0.00779f
C40 VDD VSS 0.016824f
C41 VNW B 0.617219f
C42 a_1602_69# VSS 0.005669f
C43 VDD A1 0.051939f
C44 A2 VSS 0.104058f
C45 a_3662_472# B 0.007338f
C46 C VSS 0.088883f
C47 ZN a_786_69# 0.008749f
C48 A2 A1 1.72617f
C49 a_1194_69# VSS 0.005069f
C50 C A1 0.001754f
C51 ZN VSS 1.77446f
C52 ZN A1 1.40746f
C53 B a_170_472# 2.12702f
C54 a_170_472# a_2034_472# 0.020753f
C55 VDD A2 0.052548f
C56 a_2590_472# a_170_472# 0.013379f
C57 VSS VSUBS 1.33264f
C58 VDD VSUBS 0.809429f
C59 ZN VSUBS 0.171181f
C60 C VSUBS 1.26656f
C61 B VSUBS 1.19887f
C62 A1 VSUBS 1.12703f
C63 A2 VSUBS 1.09165f
C64 VNW VSUBS 6.53302f
C65 a_170_472# VSUBS 0.077257f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 VNW VPW A3 VDD VSS ZN A1 A2 a_1792_472# a_224_472#
+ a_1568_472# a_36_472# a_1120_472# a_672_472# VSUBS
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
C0 a_1568_472# A1 0.002055f
C1 ZN A2 0.250963f
C2 A3 VNW 0.478769f
C3 a_224_472# A2 0.002647f
C4 a_672_472# A2 0.002647f
C5 VDD VNW 0.286001f
C6 a_36_472# A2 0.993181f
C7 VDD A3 0.09322f
C8 ZN VNW 0.046016f
C9 a_1120_472# A2 0.002647f
C10 A1 A2 0.085569f
C11 a_36_472# VNW 0.031928f
C12 VSS A2 0.128956f
C13 ZN A3 1.42151f
C14 VDD ZN 0.005367f
C15 a_1568_472# A2 0.004974f
C16 a_224_472# VDD 0.010911f
C17 a_672_472# VDD 0.01105f
C18 a_1792_472# VDD 0.002998f
C19 A3 a_36_472# 0.100976f
C20 VDD a_36_472# 1.90933f
C21 VNW A1 0.520086f
C22 VSS VNW 0.009996f
C23 A3 A1 0.008795f
C24 a_1792_472# ZN 0.004144f
C25 a_1120_472# VDD 0.011157f
C26 VDD A1 0.054887f
C27 ZN a_36_472# 0.362263f
C28 a_224_472# a_36_472# 0.01823f
C29 a_672_472# a_36_472# 0.01823f
C30 a_1792_472# a_36_472# 0.022081f
C31 VSS A3 0.10353f
C32 VDD VSS 0.012739f
C33 VDD a_1568_472# 0.005385f
C34 ZN A1 1.56829f
C35 a_1792_472# A1 0.006624f
C36 VNW A2 0.539636f
C37 a_1120_472# a_36_472# 0.01951f
C38 a_36_472# A1 0.174868f
C39 VSS ZN 2.18568f
C40 VSS a_36_472# 0.020716f
C41 A3 A2 1.6562f
C42 VDD A2 0.082489f
C43 a_36_472# a_1568_472# 0.025433f
C44 VSS A1 0.115774f
C45 VSS VSUBS 0.918064f
C46 ZN VSUBS 0.159858f
C47 VDD VSUBS 0.61695f
C48 A1 VSUBS 1.35739f
C49 A3 VSUBS 1.33073f
C50 A2 VSUBS 1.29013f
C51 VNW VSUBS 4.79254f
C52 a_36_472# VSUBS 0.137725f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 VNW VPW A3 VDD VSS ZN A1 A2 a_468_472# a_244_472#
+ a_1130_472# a_906_472# VSUBS
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 ZN VSS 1.3936f
C1 A2 VSS 0.043139f
C2 A1 ZN 0.084783f
C3 a_244_472# VDD 0.00632f
C4 A2 A1 0.570018f
C5 a_906_472# VDD 0.011614f
C6 VNW VSS 0.007164f
C7 VNW A1 0.254404f
C8 a_1130_472# VDD 0.011629f
C9 A1 VSS 0.044587f
C10 A3 VDD 0.178286f
C11 A3 a_244_472# 0.010666f
C12 A3 a_906_472# 0.017829f
C13 ZN VDD 0.579119f
C14 A2 VDD 0.038421f
C15 VDD a_468_472# 0.00502f
C16 ZN a_244_472# 0.019831f
C17 a_906_472# ZN 0.002855f
C18 A3 a_1130_472# 0.016495f
C19 VNW VDD 0.178574f
C20 VDD VSS 0.009106f
C21 ZN a_1130_472# 0.001342f
C22 A3 ZN 1.03634f
C23 A3 A2 0.624599f
C24 A3 a_468_472# 0.010018f
C25 A1 VDD 0.038139f
C26 A3 VNW 0.28584f
C27 A2 ZN 0.694728f
C28 A3 VSS 0.0525f
C29 ZN a_468_472# 0.015602f
C30 A3 A1 0.292395f
C31 VNW ZN 0.031771f
C32 A2 VNW 0.241313f
C33 VSS VSUBS 0.509614f
C34 ZN VSUBS 0.172636f
C35 VDD VSUBS 0.441158f
C36 A1 VSUBS 0.622214f
C37 A2 VSUBS 0.627317f
C38 A3 VSUBS 0.692739f
C39 VNW VSUBS 2.70396f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 VNW VPW B C VDD VSS ZN A1 A2 a_1492_488#
+ a_244_68# a_1044_488# a_636_68# a_36_488# VSUBS
X0 VSS B ZN VSUBS nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VSUBS nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
C0 A2 ZN 0.752866f
C1 ZN a_244_68# 0.001328f
C2 A2 B 0.036672f
C3 A2 VNW 0.280457f
C4 A2 A1 0.652956f
C5 A1 a_244_68# 0.003444f
C6 a_1044_488# B 0.012375f
C7 VSS a_636_68# 0.002222f
C8 a_1492_488# VDD 0.00909f
C9 ZN VDD 0.004894f
C10 VDD VNW 0.191798f
C11 B VDD 0.04259f
C12 VSS a_36_488# 0.005331f
C13 A1 VDD 0.026261f
C14 B a_1492_488# 0.007233f
C15 C VDD 0.040747f
C16 ZN VNW 0.028815f
C17 ZN B 0.413891f
C18 A1 ZN 0.372797f
C19 ZN C 0.191881f
C20 B VNW 0.298561f
C21 A1 VNW 0.25321f
C22 A2 a_36_488# 0.076279f
C23 C B 0.560408f
C24 C VNW 0.268332f
C25 a_1044_488# a_36_488# 0.018358f
C26 ZN a_636_68# 0.00593f
C27 a_36_488# VDD 1.67897f
C28 A2 VSS 0.077665f
C29 VSS a_244_68# 0.004878f
C30 a_36_488# a_1492_488# 0.017313f
C31 ZN a_36_488# 0.459425f
C32 a_36_488# VNW 0.010653f
C33 B a_36_488# 0.80489f
C34 A1 a_36_488# 0.031215f
C35 C a_36_488# 0.041645f
C36 VSS VDD 0.009527f
C37 ZN VSS 0.708286f
C38 VSS B 0.089442f
C39 VSS VNW 0.008434f
C40 A1 VSS 0.090485f
C41 A2 VDD 0.02614f
C42 C VSS 0.05406f
C43 a_1044_488# VDD 0.004195f
C44 VSS VSUBS 0.653933f
C45 VDD VSUBS 0.406726f
C46 ZN VSUBS 0.089692f
C47 C VSUBS 0.626227f
C48 B VSUBS 0.654892f
C49 A1 VSUBS 0.552174f
C50 A2 VSUBS 0.559992f
C51 VNW VSUBS 3.2261f
C52 a_36_488# VSUBS 0.101145f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 VNW VPW A3 VDD VSS Z A1 A2 a_244_524# a_2215_68#
+ a_56_524# a_718_524# a_728_93# a_1936_472# a_1336_472# VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
C0 a_1336_472# VNW 0.144065f
C1 Z a_1336_472# 0.021039f
C2 a_728_93# VNW 0.346549f
C3 a_1936_472# VNW 0.004015f
C4 Z a_728_93# 0.402606f
C5 Z a_1936_472# 0.337902f
C6 a_952_93# a_728_93# 0.00421f
C7 A2 VSS 0.047538f
C8 a_718_524# A2 0.107911f
C9 A3 VSS 0.056027f
C10 VDD a_244_524# 0.004322f
C11 A2 VNW 0.369075f
C12 a_56_524# VDD 0.049641f
C13 A1 VSS 0.139902f
C14 a_1336_472# VDD 0.033982f
C15 A3 VNW 0.268193f
C16 Z A3 0.259021f
C17 A1 a_718_524# 0.026418f
C18 a_728_93# VDD 0.575073f
C19 a_1936_472# VDD 0.595117f
C20 a_56_524# a_728_93# 0.016741f
C21 A1 VNW 0.293766f
C22 a_728_93# a_1336_472# 0.62718f
C23 a_1936_472# a_1336_472# 0.004622f
C24 a_1936_472# a_728_93# 0.105997f
C25 A2 a_244_524# 0.004824f
C26 VSS VNW 0.007756f
C27 A2 VDD 0.208821f
C28 Z VSS 0.277351f
C29 a_56_524# A2 0.908796f
C30 a_2215_68# VSS 0.004309f
C31 a_718_524# VNW 0.020055f
C32 a_1336_472# A2 0.001757f
C33 A3 VDD 0.028848f
C34 a_728_93# A2 0.416172f
C35 Z VNW 0.028011f
C36 A3 a_1336_472# 0.490376f
C37 Z a_2215_68# 0.008507f
C38 A1 VDD 0.018915f
C39 A3 a_728_93# 0.720358f
C40 a_1936_472# A3 0.018144f
C41 a_56_524# A1 0.569057f
C42 a_1336_472# a_1524_472# 0.001046f
C43 VDD VSS 0.013872f
C44 a_728_93# A1 0.12992f
C45 a_56_524# VSS 0.214447f
C46 a_728_93# a_1524_472# 0.007139f
C47 a_718_524# VDD 0.554575f
C48 a_56_524# a_718_524# 0.009198f
C49 a_1336_472# VSS 0.326133f
C50 a_728_93# VSS 0.709567f
C51 VDD VNW 0.360391f
C52 Z VDD 0.01058f
C53 a_56_524# VNW 0.188846f
C54 a_728_93# a_718_524# 0.329834f
C55 A1 A2 0.321942f
C56 VSS VSUBS 0.861752f
C57 Z VSUBS 0.085787f
C58 A1 VSUBS 0.602985f
C59 A2 VSUBS 0.640744f
C60 VDD VSUBS 0.543474f
C61 A3 VSUBS 0.593976f
C62 VNW VSUBS 4.270391f
C63 a_1936_472# VSUBS 0.009918f
C64 a_718_524# VSUBS 0.005143f
C65 a_56_524# VSUBS 0.41096f
C66 a_728_93# VSUBS 0.654825f
C67 a_1336_472# VSUBS 0.316639f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VNW VPW VDD VSS ZN A1 A2 a_652_68# a_244_68#
+ VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
C0 a_244_68# A1 0.004867f
C1 a_652_68# VSS 0.003855f
C2 ZN A1 0.363066f
C3 A1 VDD 0.050088f
C4 A1 VSS 0.115936f
C5 ZN A2 0.891023f
C6 VDD A2 0.070487f
C7 A2 VSS 0.057292f
C8 A1 VNW 0.232646f
C9 a_244_68# ZN 0.001926f
C10 a_244_68# VSS 0.006834f
C11 VNW A2 0.277885f
C12 ZN VDD 0.409997f
C13 ZN VSS 0.2597f
C14 VDD VSS 0.020712f
C15 A1 A2 0.708017f
C16 ZN VNW 0.033841f
C17 VNW VDD 0.123338f
C18 VNW VSS 0.008805f
C19 ZN a_652_68# 0.008436f
C20 VSS VSUBS 0.385688f
C21 ZN VSUBS 0.120217f
C22 VDD VSUBS 0.305683f
C23 A1 VSUBS 0.522064f
C24 A2 VSUBS 0.568932f
C25 VNW VSUBS 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 VNW VPW A2 A3 B VDD VSS ZN A1 a_36_68# a_1612_497#
+ a_692_497# a_1388_497# a_960_497# VSUBS
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
C0 VSS a_36_68# 2.0408f
C1 a_960_497# ZN 0.012124f
C2 ZN a_36_68# 1.49222f
C3 VSS VDD 0.010407f
C4 VNW A2 0.281901f
C5 a_1612_497# A1 0.003158f
C6 ZN VDD 1.08837f
C7 A2 A3 1.11591f
C8 a_692_497# A3 0.019827f
C9 ZN VSS 0.006088f
C10 B a_36_68# 0.184521f
C11 A2 A1 0.703324f
C12 VNW a_36_68# 0.001442f
C13 B VDD 0.119783f
C14 a_960_497# A3 0.014254f
C15 VNW VDD 0.248379f
C16 a_36_68# A3 0.036843f
C17 B VSS 0.047409f
C18 a_1388_497# A2 0.008156f
C19 VDD A3 0.555327f
C20 a_1612_497# A2 0.006056f
C21 VNW VSS 0.008187f
C22 B ZN 0.244028f
C23 a_36_68# A1 0.158235f
C24 VNW ZN 0.025446f
C25 VSS A3 0.03178f
C26 VDD A1 0.091309f
C27 ZN A3 1.02771f
C28 a_692_497# A2 0.001398f
C29 VSS A1 0.032188f
C30 a_1388_497# VDD 0.005409f
C31 ZN A1 0.619225f
C32 VNW B 0.309147f
C33 a_1612_497# VDD 0.009412f
C34 B A3 0.036798f
C35 VNW A3 0.297068f
C36 a_960_497# A2 0.003506f
C37 a_1388_497# ZN 0.001168f
C38 a_36_68# A2 0.032025f
C39 VDD A2 0.030601f
C40 a_692_497# VDD 0.00542f
C41 VNW A1 0.279057f
C42 VSS A2 0.030287f
C43 A3 A1 0.206693f
C44 ZN A2 0.152712f
C45 a_692_497# ZN 0.018589f
C46 a_960_497# VDD 0.003264f
C47 VDD a_36_68# 0.001802f
C48 a_1388_497# A3 0.02079f
C49 a_1612_497# A3 0.030605f
C50 VSS VSUBS 0.663038f
C51 ZN VSUBS 0.080495f
C52 VDD VSUBS 0.512998f
C53 A1 VSUBS 0.643779f
C54 A2 VSUBS 0.561227f
C55 A3 VSUBS 0.573818f
C56 B VSUBS 0.585725f
C57 VNW VSUBS 3.48825f
C58 a_36_68# VSUBS 0.048026f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 VNW VPW D Q RN VDD VSS CLK a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_2248_156#
+ a_2560_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 RN a_2560_156# 0.038779f
C1 a_36_151# a_1204_472# 0.006996f
C2 RN a_1308_423# 0.079294f
C3 VDD a_1204_472# 0.282626f
C4 VSS a_3041_156# 0.004935f
C5 a_2560_156# a_2248_156# 0.119687f
C6 a_1000_472# a_1308_423# 0.934191f
C7 a_1308_423# a_2248_156# 0.056721f
C8 a_36_151# a_2665_112# 0.019033f
C9 RN a_1000_472# 0.0832f
C10 VDD Q 0.260055f
C11 RN a_2248_156# 0.080362f
C12 a_36_151# D 0.094113f
C13 VDD a_2665_112# 0.152571f
C14 VSS Q 0.170514f
C15 VSS a_2665_112# 0.21484f
C16 a_1000_472# a_2248_156# 0.001232f
C17 VDD D 0.009367f
C18 VSS a_1288_156# 0.001702f
C19 a_796_472# a_1000_472# 0.048436f
C20 VSS D 0.064618f
C21 VNW a_36_151# 1.28833f
C22 a_36_151# a_448_472# 0.536965f
C23 a_1308_423# a_1204_472# 0.026665f
C24 VNW VDD 0.546785f
C25 RN a_3041_156# 0.014924f
C26 VDD a_448_472# 0.456269f
C27 VSS VNW 0.012596f
C28 RN a_1204_472# 0.021039f
C29 VSS a_448_472# 1.20207f
C30 a_2560_156# a_2665_112# 0.116229f
C31 a_1000_472# a_1204_472# 0.66083f
C32 RN a_2665_112# 0.322698f
C33 Q a_2248_156# 0.013765f
C34 a_2665_112# a_2248_156# 0.63615f
C35 VNW a_2560_156# 0.019282f
C36 a_2560_156# a_448_472# 0.277491f
C37 VNW a_1308_423# 0.149014f
C38 a_1308_423# a_448_472# 0.882105f
C39 a_796_472# D 0.082858f
C40 RN VNW 0.304626f
C41 RN a_448_472# 0.078731f
C42 VNW a_1000_472# 0.241357f
C43 a_1000_472# a_448_472# 0.361958f
C44 VNW a_2248_156# 0.181292f
C45 VDD a_36_151# 0.417101f
C46 a_2665_112# a_3041_156# 0.001841f
C47 a_2248_156# a_448_472# 0.510371f
C48 VNW a_796_472# 0.010232f
C49 VSS a_36_151# 0.291264f
C50 a_796_472# a_448_472# 0.401636f
C51 VNW CLK 0.137037f
C52 a_448_472# CLK 0.002757f
C53 VSS VDD 0.02167f
C54 a_1456_156# a_448_472# 0.00227f
C55 Q a_2665_112# 0.263315f
C56 VNW a_1204_472# 0.016269f
C57 a_1204_472# a_448_472# 0.008996f
C58 a_36_151# a_2560_156# 0.003674f
C59 a_1308_423# a_36_151# 0.05539f
C60 VDD a_2560_156# 0.00302f
C61 VNW Q 0.026596f
C62 VNW a_2665_112# 0.486803f
C63 VDD a_1308_423# 0.094185f
C64 VSS a_2560_156# 0.128503f
C65 RN a_36_151# 0.080119f
C66 a_2665_112# a_448_472# 0.020455f
C67 VSS a_1308_423# 0.013866f
C68 VNW D 0.128231f
C69 a_1288_156# a_448_472# 0.002067f
C70 a_1000_472# a_36_151# 0.08126f
C71 RN VDD 0.035003f
C72 D a_448_472# 0.328788f
C73 a_36_151# a_2248_156# 0.042802f
C74 VSS RN 0.436942f
C75 VDD a_1000_472# 0.119211f
C76 a_796_472# a_36_151# 0.011851f
C77 VDD a_2248_156# 1.12036f
C78 VSS a_1000_472# 0.04356f
C79 a_36_151# CLK 0.669598f
C80 VSS a_2248_156# 0.030372f
C81 VSS a_796_472# 0.05215f
C82 VNW a_448_472# 0.341284f
C83 VDD CLK 0.02303f
C84 VSS CLK 0.021952f
C85 VSS a_1456_156# 0.001901f
C86 Q VSUBS 0.061347f
C87 VSS VSUBS 1.33519f
C88 RN VSUBS 1.37098f
C89 D VSUBS 0.253406f
C90 VDD VSUBS 0.859994f
C91 CLK VSUBS 0.291241f
C92 VNW VSUBS 6.48579f
C93 a_2560_156# VSUBS 0.016968f
C94 a_2665_112# VSUBS 0.91969f
C95 a_2248_156# VSUBS 0.30886f
C96 a_1204_472# VSUBS 0.012971f
C97 a_1000_472# VSUBS 0.291735f
C98 a_796_472# VSUBS 0.023206f
C99 a_1308_423# VSUBS 0.279043f
C100 a_448_472# VSUBS 0.684413f
C101 a_36_151# VSUBS 1.43587f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 VNW VPW A3 A4 VDD VSS ZN A1 A2 a_438_68#
+ a_244_68# a_1254_68# a_1060_68# a_632_68# a_1458_68# VSUBS
X0 a_1458_68# A3 a_1254_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
C0 ZN A2 0.068627f
C1 A1 ZN 0.071728f
C2 A4 VSS 0.056757f
C3 VDD VSS 0.004026f
C4 A1 VNW 0.345207f
C5 VNW A2 0.317841f
C6 A3 VSS 0.248503f
C7 a_1060_68# ZN 0.007219f
C8 a_1254_68# ZN 0.008913f
C9 A4 VDD 0.047422f
C10 ZN a_632_68# 0.001673f
C11 A4 A3 0.297972f
C12 a_438_68# VSS 0.00542f
C13 VDD A3 0.040467f
C14 A1 A2 0.516286f
C15 ZN VSS 0.89636f
C16 VNW VSS 0.006403f
C17 A4 ZN 1.94271f
C18 VDD ZN 1.39778f
C19 a_244_68# VSS 0.007139f
C20 a_438_68# A3 0.007312f
C21 A4 VNW 0.388525f
C22 a_1458_68# VSS 0.002548f
C23 VDD VNW 0.1769f
C24 A3 ZN 0.881941f
C25 A1 VSS 0.037456f
C26 A2 VSS 0.036637f
C27 A3 VNW 0.300046f
C28 a_1060_68# VSS 0.001868f
C29 a_244_68# A3 0.007f
C30 A1 A4 0.451294f
C31 A4 A2 0.762551f
C32 a_1254_68# VSS 0.002331f
C33 A1 VDD 0.044019f
C34 VDD A2 0.041932f
C35 a_632_68# VSS 0.005832f
C36 A1 A3 0.831807f
C37 A3 A2 0.40854f
C38 VNW ZN 0.062752f
C39 a_1060_68# A3 0.004303f
C40 a_1254_68# A3 0.004873f
C41 a_1458_68# ZN 0.01082f
C42 A3 a_632_68# 0.0083f
C43 VSS VSUBS 0.597574f
C44 VDD VSUBS 0.397078f
C45 ZN VSUBS 0.12583f
C46 A1 VSUBS 0.558392f
C47 A2 VSUBS 0.513744f
C48 A3 VSUBS 0.547819f
C49 A4 VSUBS 0.580825f
C50 VNW VSUBS 3.05206f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VNW VPW VDD VSS I ZN VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
C0 ZN I 0.614595f
C1 ZN VNW 0.025997f
C2 ZN VDD 0.24022f
C3 VSS ZN 0.15979f
C4 I VNW 0.283715f
C5 I VDD 0.164681f
C6 VSS I 0.071429f
C7 VNW VDD 0.103267f
C8 VSS VNW 0.01054f
C9 VSS VDD 0.022662f
C10 VSS VSUBS 0.345063f
C11 ZN VSUBS 0.094435f
C12 VDD VSUBS 0.235951f
C13 I VSUBS 0.642286f
C14 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 VNW VPW A3 B1 B2 VDD VSS ZN A1 A2 a_468_472#
+ a_224_472# a_244_68# a_916_472# VSUBS
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
C0 A3 a_224_472# 0.012212f
C1 B1 VDD 0.015317f
C2 a_244_68# a_468_472# 0.022611f
C3 VDD a_244_68# 0.520053f
C4 A2 A1 0.038953f
C5 A2 a_468_472# 0.002382f
C6 A1 a_468_472# 0.001494f
C7 a_244_68# a_224_472# 0.004752f
C8 A3 VSS 0.046517f
C9 A2 VDD 0.071137f
C10 A3 VNW 0.13805f
C11 VDD A1 0.015114f
C12 VDD a_468_472# 0.005594f
C13 B2 B1 0.038725f
C14 a_244_68# a_916_472# 0.018012f
C15 A2 a_224_472# 0.014544f
C16 B2 a_244_68# 0.29062f
C17 B1 VSS 0.072063f
C18 B1 VNW 0.116377f
C19 B1 ZN 0.457921f
C20 VSS a_244_68# 0.329999f
C21 VNW a_244_68# 0.043485f
C22 a_244_68# ZN 0.2576f
C23 VDD a_224_472# 0.016257f
C24 A2 VSS 0.030842f
C25 A2 VNW 0.121626f
C26 VSS A1 0.029231f
C27 VNW A1 0.125824f
C28 VDD a_916_472# 0.004169f
C29 ZN A1 0.164807f
C30 B2 VDD 0.018546f
C31 VDD VSS 0.027141f
C32 VNW VDD 0.158216f
C33 VDD ZN 0.006472f
C34 A3 a_244_68# 0.010697f
C35 VSS a_224_472# 0.00124f
C36 A2 A3 0.129823f
C37 B1 a_244_68# 0.212448f
C38 B2 VSS 0.072128f
C39 ZN a_916_472# 0.008827f
C40 B2 VNW 0.125762f
C41 B2 ZN 0.371232f
C42 A3 VDD 0.236688f
C43 VNW VSS 0.013582f
C44 B1 A1 0.13457f
C45 VSS ZN 0.069913f
C46 VNW ZN 0.012941f
C47 A2 a_244_68# 0.356992f
C48 a_244_68# A1 0.480797f
C49 VSS VSUBS 0.474343f
C50 ZN VSUBS 0.00986f
C51 VDD VSUBS 0.363224f
C52 B2 VSUBS 0.282623f
C53 B1 VSUBS 0.257203f
C54 A1 VSUBS 0.255736f
C55 A2 VSUBS 0.254473f
C56 A3 VSUBS 0.308666f
C57 VNW VSUBS 2.35586f
C58 a_244_68# VSUBS 0.138666f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 VNW VPW A3 VDD VSS ZN A1 A2 a_244_567# a_718_527#
+ a_2172_497# a_56_567# a_1948_68# a_728_93# a_1296_93# VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
C0 a_1948_68# ZN 0.381585f
C1 a_1296_93# ZN 0.029802f
C2 a_1504_93# a_1296_93# 0.003723f
C3 A1 A2 0.757944f
C4 a_1948_68# A3 0.069927f
C5 A3 a_1296_93# 0.356198f
C6 A2 VDD 0.210416f
C7 VSS a_56_567# 0.400197f
C8 a_728_93# A2 0.516752f
C9 ZN VSS 0.004739f
C10 a_1948_68# VDD 0.001604f
C11 a_1296_93# VDD 0.030892f
C12 a_718_527# A2 0.141128f
C13 A2 VNW 0.388997f
C14 a_1504_93# VSS 0.003902f
C15 a_1948_68# a_728_93# 0.02618f
C16 a_728_93# a_1296_93# 0.624643f
C17 a_244_567# A2 0.004089f
C18 a_1948_68# VNW 0.002346f
C19 a_1296_93# VNW 0.155715f
C20 A3 VSS 0.047056f
C21 VSS A1 0.0538f
C22 VSS VDD 0.011823f
C23 a_2172_497# ZN 0.03345f
C24 a_728_93# VSS 0.328386f
C25 A1 a_56_567# 0.368741f
C26 A3 ZN 0.033406f
C27 VSS VNW 0.009921f
C28 VSS a_952_93# 0.003841f
C29 a_56_567# VDD 0.056918f
C30 a_728_93# a_56_567# 0.070648f
C31 ZN VDD 0.47211f
C32 a_728_93# ZN 0.663929f
C33 a_56_567# a_718_527# 0.00772f
C34 a_56_567# VNW 0.187311f
C35 a_2172_497# VDD 0.010751f
C36 a_2172_497# a_728_93# 0.010602f
C37 a_56_567# a_244_567# 0.00105f
C38 ZN VNW 0.032895f
C39 a_1296_93# A2 0.002759f
C40 A3 VDD 0.022483f
C41 A1 VDD 0.022573f
C42 a_728_93# A3 0.721889f
C43 a_728_93# A1 0.281966f
C44 a_1948_68# a_1296_93# 0.005923f
C45 A3 VNW 0.298581f
C46 a_728_93# VDD 0.78216f
C47 A1 a_718_527# 0.023145f
C48 A1 VNW 0.342048f
C49 a_718_527# VDD 0.618394f
C50 VDD VNW 0.370487f
C51 VSS A2 0.051212f
C52 a_728_93# a_718_527# 0.21558f
C53 a_728_93# VNW 0.385878f
C54 a_244_567# VDD 0.006111f
C55 a_728_93# a_952_93# 0.003723f
C56 a_718_527# VNW 0.020227f
C57 a_1948_68# VSS 0.719859f
C58 a_1296_93# VSS 0.379749f
C59 a_56_567# A2 0.174541f
C60 VSS VSUBS 0.875791f
C61 ZN VSUBS 0.08517f
C62 A1 VSUBS 0.604039f
C63 A2 VSUBS 0.633287f
C64 VDD VSUBS 0.584594f
C65 A3 VSUBS 0.573218f
C66 VNW VSUBS 4.42794f
C67 a_1948_68# VSUBS 0.022025f
C68 a_718_527# VSUBS 0.001795f
C69 a_56_567# VSUBS 0.424713f
C70 a_728_93# VSUBS 0.65929f
C71 a_1296_93# VSUBS 0.317801f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 VNW VPW A2 ZN A1 B C VDD VSS a_36_68# a_244_497#
+ a_1657_68# a_1229_68# a_716_497# VSUBS
X0 a_1229_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
C0 B VSS 0.032629f
C1 VDD A1 0.033883f
C2 ZN A2 1.02528f
C3 ZN VSS 0.004788f
C4 VNW a_36_68# 0.00468f
C5 VNW B 0.311256f
C6 VNW ZN 0.042076f
C7 B a_36_68# 0.587375f
C8 a_716_497# A2 0.010693f
C9 ZN a_36_68# 0.528658f
C10 ZN B 0.3603f
C11 A2 a_244_497# 0.020646f
C12 VSS C 0.04168f
C13 A1 A2 0.722847f
C14 a_1229_68# VSS 0.002856f
C15 A1 VSS 0.031008f
C16 a_1657_68# VSS 0.002208f
C17 VNW C 0.309331f
C18 VDD A2 0.147417f
C19 ZN a_716_497# 0.025301f
C20 VNW A1 0.269127f
C21 VDD VSS 0.007619f
C22 ZN a_244_497# 0.006285f
C23 a_36_68# C 0.055076f
C24 B C 0.698524f
C25 a_1229_68# a_36_68# 0.011792f
C26 a_1229_68# B 0.003462f
C27 A1 a_36_68# 0.039393f
C28 ZN C 0.501479f
C29 a_1657_68# a_36_68# 0.009002f
C30 B a_1657_68# 0.002626f
C31 ZN A1 0.622246f
C32 VNW VDD 0.219901f
C33 VDD a_36_68# 0.019083f
C34 VDD B 0.089771f
C35 VDD ZN 0.761655f
C36 A2 VSS 0.030494f
C37 VDD a_716_497# 0.008883f
C38 VNW A2 0.30827f
C39 VDD a_244_497# 0.016799f
C40 VNW VSS 0.005994f
C41 A2 a_36_68# 0.091399f
C42 A2 B 0.037237f
C43 VDD C 0.056662f
C44 a_36_68# VSS 2.1107f
C45 VSS VSUBS 0.620026f
C46 ZN VSUBS 0.062404f
C47 VDD VSUBS 0.531064f
C48 C VSUBS 0.529789f
C49 B VSUBS 0.589191f
C50 A1 VSUBS 0.58772f
C51 A2 VSUBS 0.613706f
C52 VNW VSUBS 3.34705f
C53 a_36_68# VSUBS 0.052951f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 VNW VPW A3 VDD VSS Z A1 A2 a_428_148# a_36_148#
+ VSUBS
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VSUBS nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VSUBS nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VSUBS nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VSUBS nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
C0 a_36_148# A1 0.205722f
C1 a_36_148# A3 0.477475f
C2 VNW A1 0.214361f
C3 VNW A3 0.213241f
C4 VDD A2 0.022493f
C5 Z A3 0.001054f
C6 VNW a_36_148# 0.194548f
C7 VDD A1 0.021719f
C8 VDD A3 0.022574f
C9 Z a_36_148# 0.156534f
C10 A1 a_244_148# 0.002081f
C11 VSS A2 0.004456f
C12 VNW Z 0.033257f
C13 VDD a_36_148# 0.556761f
C14 VSS A1 0.00434f
C15 VNW VDD 0.134134f
C16 a_428_148# A3 0.001335f
C17 a_36_148# a_244_148# 0.004781f
C18 VSS A3 0.005273f
C19 VDD Z 0.164783f
C20 A1 A2 0.307806f
C21 a_428_148# a_36_148# 0.007047f
C22 VSS a_36_148# 0.798993f
C23 A2 A3 0.340591f
C24 VNW VSS 0.007319f
C25 VSS Z 0.093779f
C26 a_36_148# A2 0.141951f
C27 VNW A2 0.189332f
C28 VDD VSS 0.012823f
C29 VSS VSUBS 0.415001f
C30 Z VSUBS 0.095371f
C31 VDD VSUBS 0.277732f
C32 A3 VSUBS 0.275015f
C33 A2 VSUBS 0.257076f
C34 A1 VSUBS 0.330738f
C35 VNW VSUBS 2.00777f
C36 a_36_148# VSUBS 0.388358f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 VNW VPW A3 VDD VSS ZN A1 A2 a_1044_68# a_452_68#
+ a_276_68# a_860_68# VSUBS
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VSUBS nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 A3 A2 1.13496f
C1 VNW A2 0.279783f
C2 VDD A3 0.099291f
C3 a_276_68# ZN 0.007178f
C4 VDD VNW 0.172362f
C5 a_276_68# VSS 0.003438f
C6 A2 ZN 0.082264f
C7 VDD ZN 0.550625f
C8 A2 VSS 0.130985f
C9 a_1044_68# A2 0.006328f
C10 VDD VSS 0.009236f
C11 A2 A1 0.708241f
C12 ZN a_860_68# 0.001808f
C13 VDD A1 0.041745f
C14 a_860_68# VSS 0.005864f
C15 VNW A3 0.347673f
C16 a_452_68# ZN 0.007752f
C17 a_452_68# VSS 0.003244f
C18 A3 ZN 1.24554f
C19 VNW ZN 0.034063f
C20 a_452_68# A1 0.001247f
C21 A3 VSS 0.074424f
C22 VNW VSS 0.007349f
C23 VDD A2 0.041181f
C24 A3 A1 0.037905f
C25 VNW A1 0.280755f
C26 ZN VSS 0.476547f
C27 a_1044_68# ZN 0.001223f
C28 A2 a_860_68# 0.003842f
C29 a_1044_68# VSS 0.00861f
C30 A1 ZN 0.430404f
C31 A1 VSS 0.050488f
C32 VSS VSUBS 0.511432f
C33 ZN VSUBS 0.112753f
C34 VDD VSUBS 0.407724f
C35 A1 VSUBS 0.540441f
C36 A2 VSUBS 0.524145f
C37 A3 VSUBS 0.582222f
C38 VNW VSUBS 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 VNW VPW A3 A4 VDD VSS ZN A1 A2 a_692_473#
+ a_254_473# a_66_473# a_2700_473# a_1660_473# a_3220_473# a_1212_473# a_2180_473#
+ a_3740_473# a_1920_473# VSUBS
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
C0 a_66_473# A4 0.100571f
C1 a_66_473# a_3220_473# 0.021354f
C2 a_1920_473# ZN 0.017667f
C3 a_66_473# a_2180_473# 0.020817f
C4 a_66_473# a_1212_473# 0.018664f
C5 A3 VSS 0.078892f
C6 A2 VNW 0.584134f
C7 a_1660_473# VDD 0.008572f
C8 VDD VNW 0.394018f
C9 VDD a_254_473# 0.012952f
C10 a_66_473# a_3740_473# 0.028219f
C11 VDD a_692_473# 0.017923f
C12 A4 VSS 0.099821f
C13 A3 A4 1.96796f
C14 a_66_473# a_1660_473# 0.035002f
C15 a_66_473# VNW 0.040351f
C16 a_66_473# a_254_473# 0.016207f
C17 a_1920_473# VDD 0.004058f
C18 a_2700_473# ZN 0.019492f
C19 A2 ZN 2.14591f
C20 A1 VNW 0.553741f
C21 VDD ZN 0.007051f
C22 a_66_473# a_692_473# 0.022803f
C23 VNW VSS 0.006947f
C24 a_1660_473# A3 0.0054f
C25 a_66_473# a_1920_473# 0.023791f
C26 VNW A3 0.567739f
C27 a_66_473# ZN 0.956309f
C28 a_2700_473# VDD 0.003457f
C29 VNW A4 0.513548f
C30 A2 VDD 0.054912f
C31 A1 ZN 1.60655f
C32 ZN VSS 4.39577f
C33 A3 ZN 0.417545f
C34 a_2700_473# a_66_473# 0.021497f
C35 a_66_473# A2 0.182327f
C36 a_66_473# VDD 3.19476f
C37 A2 A1 2.13585f
C38 A4 ZN 1.44735f
C39 A1 VDD 0.055928f
C40 ZN a_3220_473# 0.019778f
C41 ZN a_2180_473# 0.018904f
C42 A2 VSS 0.076134f
C43 VDD VSS 0.009708f
C44 A2 A3 0.0303f
C45 VDD A3 0.086829f
C46 ZN a_3740_473# 0.004594f
C47 a_66_473# A1 0.077909f
C48 a_1660_473# ZN 0.00216f
C49 VNW ZN 0.038639f
C50 VDD A4 0.110338f
C51 VDD a_3220_473# 0.003326f
C52 a_66_473# VSS 0.01197f
C53 VDD a_2180_473# 0.00368f
C54 a_66_473# A3 1.66251f
C55 a_1212_473# VDD 0.014305f
C56 A1 VSS 0.093176f
C57 A2 a_3740_473# 0.010293f
C58 VDD a_3740_473# 0.003118f
C59 VSS VSUBS 1.3434f
C60 ZN VSUBS 0.240026f
C61 VDD VSUBS 0.844436f
C62 A1 VSUBS 1.40024f
C63 A2 VSUBS 1.30271f
C64 A4 VSUBS 1.33565f
C65 A3 VSUBS 1.29175f
C66 VNW VSUBS 6.70706f
C67 a_66_473# VSUBS 0.11665f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 VNW VPW B VDD VSS ZN A1 A2 a_49_472# a_1133_69#
+ a_741_69# VSUBS
X0 VSS A2 a_1133_69# VSUBS nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VSUBS nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VSUBS nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
C0 VDD A1 0.028601f
C1 a_49_472# VNW 0.012852f
C2 VDD A2 0.029358f
C3 A1 A2 0.809974f
C4 ZN VNW 0.025755f
C5 A2 a_741_69# 0.001142f
C6 ZN a_49_472# 0.475008f
C7 VDD B 0.045174f
C8 ZN a_1133_69# 0.001193f
C9 VDD VSS 0.009099f
C10 B A2 0.029994f
C11 A1 VSS 0.129775f
C12 VSS a_741_69# 0.002035f
C13 VSS A2 0.047574f
C14 B VSS 0.061328f
C15 VDD VNW 0.151549f
C16 A1 VNW 0.241301f
C17 VDD a_49_472# 1.09818f
C18 A1 a_49_472# 0.03417f
C19 A2 VNW 0.272677f
C20 ZN VDD 0.008463f
C21 ZN A1 0.182845f
C22 A1 a_1133_69# 0.003427f
C23 a_49_472# A2 0.086717f
C24 ZN a_741_69# 0.006341f
C25 B VNW 0.260678f
C26 ZN A2 0.800412f
C27 a_49_472# B 0.234399f
C28 VSS VNW 0.0086f
C29 ZN B 0.20884f
C30 a_49_472# VSS 0.01207f
C31 ZN VSS 0.784804f
C32 a_1133_69# VSS 0.00441f
C33 VSS VSUBS 0.510011f
C34 ZN VSUBS 0.070911f
C35 VDD VSUBS 0.327438f
C36 A1 VSUBS 0.556927f
C37 A2 VSUBS 0.56333f
C38 B VSUBS 0.662515f
C39 VNW VSUBS 2.52991f
C40 a_49_472# VSUBS 0.098072f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VNW VPW VSS ZN I VDD VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD I 0.074838f
C1 ZN I 0.58604f
C2 VNW VSS 0.010163f
C3 VDD VSS 0.023187f
C4 ZN VSS 0.179304f
C5 VNW VDD 0.097124f
C6 VNW ZN 0.027829f
C7 VDD ZN 0.266247f
C8 I VSS 0.091531f
C9 VNW I 0.285482f
C10 VSS VSUBS 0.308828f
C11 ZN VSUBS 0.100523f
C12 VDD VSUBS 0.240805f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VNW VPW VSS CLK VDD D Q SETN a_448_472#
+ a_36_151# a_1293_527# a_3081_151# a_1284_156# a_1040_527# a_1353_112# a_836_156#
+ a_1697_156# a_2449_156# a_3129_107# a_2225_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VSUBS nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VSUBS nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VSUBS nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VSUBS nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VSUBS nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VSUBS nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
C0 SETN a_1040_527# 0.063241f
C1 a_2225_156# a_1353_112# 0.152869f
C2 a_1353_112# a_448_472# 0.317251f
C3 a_2225_156# a_3081_151# 0.004129f
C4 a_1040_527# a_448_472# 0.869605f
C5 VDD D 0.004944f
C6 a_36_151# VDD 1.41468f
C7 a_1353_112# VNW 0.219511f
C8 VSS VDD 0.013814f
C9 VNW a_1040_527# 0.223863f
C10 D a_836_156# 0.108102f
C11 a_1284_156# a_448_472# 0.002691f
C12 a_36_151# a_836_156# 0.015697f
C13 VSS a_836_156# 0.050008f
C14 Q a_3129_107# 0.179468f
C15 a_1353_112# VDD 0.016257f
C16 a_36_151# D 0.092705f
C17 a_1040_527# VDD 0.039677f
C18 VSS D 0.067877f
C19 a_36_151# VSS 0.286331f
C20 Q VNW 0.031621f
C21 a_1040_527# a_836_156# 0.068207f
C22 SETN a_2449_156# 0.302222f
C23 a_448_472# a_1697_156# 0.007618f
C24 CLK a_448_472# 0.001313f
C25 a_2225_156# a_2449_156# 0.569174f
C26 a_2449_156# a_448_472# 0.056679f
C27 a_36_151# a_1353_112# 0.840879f
C28 a_3129_107# a_2449_156# 0.00955f
C29 VSS a_1353_112# 0.027348f
C30 Q VDD 0.282179f
C31 a_36_151# a_1040_527# 0.206392f
C32 VSS a_1040_527# 0.060221f
C33 CLK VNW 0.136589f
C34 VNW a_2449_156# 0.043816f
C35 VSS a_1284_156# 0.003637f
C36 a_1353_112# a_1040_527# 0.387423f
C37 a_2225_156# SETN 0.070597f
C38 SETN a_448_472# 0.083903f
C39 a_3129_107# SETN 0.089288f
C40 CLK VDD 0.022091f
C41 VDD a_2449_156# 0.208631f
C42 VSS Q 0.131272f
C43 a_2225_156# a_448_472# 0.153996f
C44 a_2225_156# a_3129_107# 0.514036f
C45 SETN VNW 0.811046f
C46 a_2225_156# VNW 0.209033f
C47 VNW a_448_472# 0.400964f
C48 a_3129_107# VNW 0.323464f
C49 a_36_151# a_1293_527# 0.008379f
C50 a_36_151# CLK 0.700974f
C51 a_36_151# a_2449_156# 0.005967f
C52 VSS CLK 0.021941f
C53 SETN VDD 0.127822f
C54 a_2225_156# VDD 0.073415f
C55 VDD a_448_472# 0.624585f
C56 a_3129_107# VDD 0.351307f
C57 a_1353_112# a_1697_156# 0.002752f
C58 VNW VDD 0.539099f
C59 a_448_472# a_836_156# 0.427756f
C60 a_1293_527# a_1040_527# 0.00215f
C61 a_2449_156# a_3081_151# 0.001203f
C62 a_36_151# SETN 0.077775f
C63 VSS SETN 0.008083f
C64 VNW a_836_156# 0.01368f
C65 a_448_472# D 0.400104f
C66 a_2225_156# a_36_151# 0.153684f
C67 a_36_151# a_448_472# 0.473132f
C68 a_2225_156# VSS 1.18908f
C69 VSS a_448_472# 1.07431f
C70 VSS a_3129_107# 0.136769f
C71 VNW D 0.1615f
C72 a_36_151# VNW 0.909435f
C73 VSS VNW 0.009462f
C74 SETN a_1353_112# 0.072983f
C75 Q VSUBS 0.105566f
C76 VSS VSUBS 1.35707f
C77 SETN VSUBS 0.710246f
C78 D VSUBS 0.247102f
C79 VDD VSUBS 0.833181f
C80 CLK VSUBS 0.290467f
C81 VNW VSUBS 6.44257f
C82 a_2449_156# VSUBS 0.049992f
C83 a_2225_156# VSUBS 0.434082f
C84 a_3129_107# VSUBS 0.58406f
C85 a_836_156# VSUBS 0.019766f
C86 a_1040_527# VSUBS 0.302082f
C87 a_1353_112# VSUBS 0.286513f
C88 a_448_472# VSUBS 1.21246f
C89 a_36_151# VSUBS 1.31409f
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[3] ctln[4] ctln[5] ctln[6] ctln[8] ctlp[0] ctlp[1]
+ ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8] ctlp[9] clk clkc comp en
+ result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7]
+ result[8] result[9] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0]
+ trimb[1] trimb[2] trimb[3] trimb[4] valid net10 output13/a_224_472# output23/a_224_472#
+ net59 net16 net27 output25/a_224_472# cal_itt\[1\] fanout65/a_36_113# ctln[2] ctln[7]
+ net15 ctln[9] output10/a_224_472# net26 net24 output11/a_224_472# output21/a_224_472#
+ net14 output12/a_224_472# output22/a_224_472# cal net62 net20 vss vdd
XFILLER_0_17_200 vdd FILLER_0_17_200/VPW vdd vss FILLER_0_17_200/a_36_472# FILLER_0_17_200/a_572_375#
+ FILLER_0_17_200/a_124_375# FILLER_0_17_200/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vdd ANTENNA_fanout56_I/VPW vss net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_294_ vdd _294_/VPW vdd vss _008_ _104_ _106_ _294_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_432_ vdd _432_/VPW _021_ mask\[3\] net63 vss net80 vdd _432_/a_2665_112# _432_/a_448_472#
+ _432_/a_796_472# _432_/a_36_151# _432_/a_1204_472# _432_/a_3041_156# _432_/a_1000_472#
+ _432_/a_1308_423# _432_/a_1456_156# _432_/a_1288_156# _432_/a_2248_156# _432_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_363_ vdd _363_/VPW _153_ _154_ _155_ vdd vss _028_ _151_ _363_/a_36_68# _363_/a_244_472#
+ _363_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ vdd _346_/VPW _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ _346_/a_49_472#
+ _346_/a_665_69# _346_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ vdd _415_/VPW _004_ net27 net58 vss net75 vdd _415_/a_2665_112# _415_/a_448_472#
+ _415_/a_796_472# _415_/a_36_151# _415_/a_1204_472# _415_/a_3041_156# _415_/a_1000_472#
+ _415_/a_1308_423# _415_/a_1456_156# _415_/a_1288_156# _415_/a_2248_156# _415_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vdd _277_/VPW vss _094_ _093_ vdd _277_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd _200_/VPW vdd vss net20 net10 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vdd _329_/VPW vss _133_ calibrate vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd FILLER_0_19_125/VPW vdd vss FILLER_0_19_125/a_36_472# FILLER_0_19_125/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vdd ANTENNA__392__A2/VPW vss _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd FILLER_0_15_150/VPW vdd vss FILLER_0_15_150/a_36_472# FILLER_0_15_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd FILLER_0_21_142/VPW vdd vss FILLER_0_21_142/a_36_472# FILLER_0_21_142/a_572_375#
+ FILLER_0_21_142/a_124_375# FILLER_0_21_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd FILLER_0_16_73/VPW vdd vss FILLER_0_16_73/a_36_472# FILLER_0_16_73/a_572_375#
+ FILLER_0_16_73/a_124_375# FILLER_0_16_73/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 vdd output20/VPW ctlp[3] net20 vdd vss output20/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 vdd output31/VPW result[4] net31 vdd vss output31/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 vdd output42/VPW trim[4] net42 vdd vss output42/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 vdd output7/VPW ctln[0] net7 vdd vss output7/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd FILLER_0_5_117/VPW vdd vss FILLER_0_5_117/a_36_472# FILLER_0_5_117/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd FILLER_0_5_128/VPW vdd vss FILLER_0_5_128/a_36_472# FILLER_0_5_128/a_572_375#
+ FILLER_0_5_128/a_124_375# FILLER_0_5_128/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_293_ vdd _293_/VPW net31 vdd vss _106_ mask\[4\] _105_ _293_/a_36_472# _293_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_431_ vdd _431_/VPW _020_ mask\[2\] net53 vss net70 vdd _431_/a_2665_112# _431_/a_448_472#
+ _431_/a_796_472# _431_/a_36_151# _431_/a_1204_472# _431_/a_3041_156# _431_/a_1000_472#
+ _431_/a_1308_423# _431_/a_1456_156# _431_/a_1288_156# _431_/a_2248_156# _431_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_362_ vdd _362_/VPW vdd vss trim_mask\[1\] _155_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_345_ vdd _345_/VPW vss _144_ _132_ vdd _345_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ vdd _276_/VPW vss _093_ _092_ vdd _276_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ vdd _414_/VPW _003_ cal_itt\[3\] net59 vss net76 vdd _414_/a_2665_112# _414_/a_448_472#
+ _414_/a_796_472# _414_/a_36_151# _414_/a_1204_472# _414_/a_3041_156# _414_/a_1000_472#
+ _414_/a_1308_423# _414_/a_1456_156# _414_/a_1288_156# _414_/a_2248_156# _414_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vdd _328_/VPW vss _132_ _114_ vdd _328_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd FILLER_0_9_28/VPW vdd vss FILLER_0_9_28/a_1916_375# FILLER_0_9_28/a_1380_472#
+ FILLER_0_9_28/a_3260_375# FILLER_0_9_28/a_36_472# FILLER_0_9_28/a_932_472# FILLER_0_9_28/a_2812_375#
+ FILLER_0_9_28/a_2276_472# FILLER_0_9_28/a_1828_472# FILLER_0_9_28/a_3172_472# FILLER_0_9_28/a_572_375#
+ FILLER_0_9_28/a_2724_472# FILLER_0_9_28/a_124_375# FILLER_0_9_28/a_1468_375# FILLER_0_9_28/a_1020_375#
+ FILLER_0_9_28/a_484_472# FILLER_0_9_28/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_204 vdd FILLER_0_3_204/VPW vdd vss FILLER_0_3_204/a_36_472# FILLER_0_3_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ vdd _259_/VPW _078_ vdd vss _080_ _073_ _076_ _259_/a_455_68# _259_/a_271_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd FILLER_0_16_107/VPW vdd vss FILLER_0_16_107/a_36_472# FILLER_0_16_107/a_572_375#
+ FILLER_0_16_107/a_124_375# FILLER_0_16_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vdd ANTENNA_fanout79_I/VPW vss net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vdd ANTENNA__358__I/VPW vss _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 vdd output21/VPW ctlp[4] net21 vdd vss output21/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 vdd output43/VPW trimb[0] net43 vdd vss output43/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 vdd output32/VPW result[5] net32 vdd vss output32/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 vdd output10/VPW ctln[3] net10 vdd vss output10/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 vdd output8/VPW ctln[1] net8 vdd vss output8/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vdd ANTENNA_input3_I/VPW vss comp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ vdd _292_/VPW vss _105_ _098_ vdd _292_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_430_ vdd _430_/VPW _019_ mask\[1\] net63 vss net80 vdd _430_/a_2665_112# _430_/a_448_472#
+ _430_/a_796_472# _430_/a_36_151# _430_/a_1204_472# _430_/a_3041_156# _430_/a_1000_472#
+ _430_/a_1308_423# _430_/a_1456_156# _430_/a_1288_156# _430_/a_2248_156# _430_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_361_ vdd _361_/VPW vdd vss _154_ _086_ _119_ _361_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd FILLER_0_7_72/VPW vdd vss FILLER_0_7_72/a_1916_375# FILLER_0_7_72/a_1380_472#
+ FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472# FILLER_0_7_72/a_932_472# FILLER_0_7_72/a_2812_375#
+ FILLER_0_7_72/a_2276_472# FILLER_0_7_72/a_1828_472# FILLER_0_7_72/a_3172_472# FILLER_0_7_72/a_572_375#
+ FILLER_0_7_72/a_2724_472# FILLER_0_7_72/a_124_375# FILLER_0_7_72/a_1468_375# FILLER_0_7_72/a_1020_375#
+ FILLER_0_7_72/a_484_472# FILLER_0_7_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd _344_/VPW vdd vss _143_ _021_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd _275_/VPW vdd vss _092_ _069_ _091_ _275_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__191__I vdd ANTENNA__191__I/VPW vss net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ vdd _413_/VPW _002_ cal_itt\[2\] net59 vss net76 vdd _413_/a_2665_112# _413_/a_448_472#
+ _413_/a_796_472# _413_/a_36_151# _413_/a_1204_472# _413_/a_3041_156# _413_/a_1000_472#
+ _413_/a_1308_423# _413_/a_1456_156# _413_/a_1288_156# _413_/a_2248_156# _413_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_96 vdd FILLER_0_24_96/VPW vdd vss FILLER_0_24_96/a_36_472# FILLER_0_24_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd FILLER_0_24_63/VPW vdd vss FILLER_0_24_63/a_36_472# FILLER_0_24_63/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ vdd _189_/VPW vdd vss _043_ net27 mask\[0\] _189_/a_255_603# _189_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_327_ vdd _327_/VPW _131_ vdd vss _016_ _127_ _130_ _327_/a_36_472# _327_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ vdd _258_/VPW vss _079_ _078_ vdd _258_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd FILLER_0_18_171/VPW vdd vss FILLER_0_18_171/a_36_472# FILLER_0_18_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd FILLER_0_24_130/VPW vdd vss FILLER_0_24_130/a_36_472# FILLER_0_24_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vdd ANTENNA__377__A1/VPW vss _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd FILLER_0_21_133/VPW vdd vss FILLER_0_21_133/a_36_472# FILLER_0_21_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd FILLER_0_8_138/VPW vdd vss FILLER_0_8_138/a_36_472# FILLER_0_8_138/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd FILLER_0_8_127/VPW vdd vss FILLER_0_8_127/a_36_472# FILLER_0_8_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 vdd output22/VPW ctlp[5] net22 vdd vss output22/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 vdd output33/VPW result[6] net33 vdd vss output33/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 vdd output44/VPW trimb[1] net44 vdd vss output44/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 vdd output11/VPW ctln[4] net11 vdd vss output11/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 vdd output9/VPW ctln[2] net9 vdd vss output9/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vdd ANTENNA__194__I/VPW vss net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vdd _291_/VPW vss _104_ _092_ vdd _291_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd FILLER_0_4_152/VPW vdd vss FILLER_0_4_152/a_36_472# FILLER_0_4_152/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd FILLER_0_4_185/VPW vdd vss FILLER_0_4_185/a_36_472# FILLER_0_4_185/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vdd _360_/VPW vss _153_ _152_ vdd _360_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd FILLER_0_13_65/VPW vdd vss FILLER_0_13_65/a_36_472# FILLER_0_13_65/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ vdd _343_/VPW _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ _343_/a_49_472#
+ _343_/a_665_69# _343_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_274_ vdd _274_/VPW _072_ _090_ vdd vss _091_ net4 _060_ _274_/a_36_68# _274_/a_1612_497#
+ _274_/a_2124_68# _274_/a_244_497# _274_/a_2960_68# _274_/a_3368_68# _274_/a_2552_68#
+ _274_/a_1164_497# _274_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_412_ vdd _412_/VPW _001_ cal_itt\[1\] net58 vss net75 vdd _412_/a_2665_112# _412_/a_448_472#
+ _412_/a_796_472# _412_/a_36_151# _412_/a_1204_472# _412_/a_3041_156# _412_/a_1000_472#
+ _412_/a_1308_423# _412_/a_1456_156# _412_/a_1288_156# _412_/a_2248_156# _412_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__292__I vdd ANTENNA__292__I/VPW vss _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ vdd _326_/VPW _131_ vss vdd _125_ _326_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ vdd _257_/VPW _077_ vdd vss _078_ _053_ _075_ _257_/a_36_472# _257_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vdd _309_/VPW vss _116_ net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vdd ANTENNA__197__I/VPW vss net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__301__A2 vdd ANTENNA__301__A2/VPW vss _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd FILLER_0_15_142/VPW vdd vss FILLER_0_15_142/a_36_472# FILLER_0_15_142/a_572_375#
+ FILLER_0_15_142/a_124_375# FILLER_0_15_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 vdd output23/VPW ctlp[6] net23 vdd vss output23/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 vdd output45/VPW trimb[2] net45 vdd vss output45/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 vdd output34/VPW result[7] net34 vdd vss output34/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 vdd output12/VPW ctln[5] net12 vdd vss output12/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd FILLER_0_5_109/VPW vdd vss FILLER_0_5_109/a_36_472# FILLER_0_5_109/a_572_375#
+ FILLER_0_5_109/a_124_375# FILLER_0_5_109/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd FILLER_0_17_226/VPW vdd vss FILLER_0_17_226/a_36_472# FILLER_0_17_226/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd FILLER_0_4_197/VPW vdd vss FILLER_0_4_197/a_1380_472# FILLER_0_4_197/a_36_472#
+ FILLER_0_4_197/a_932_472# FILLER_0_4_197/a_572_375# FILLER_0_4_197/a_124_375# FILLER_0_4_197/a_1468_375#
+ FILLER_0_4_197/a_1020_375# FILLER_0_4_197/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd _290_/VPW vdd vss _007_ _094_ _103_ _290_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd FILLER_0_9_223/VPW vdd vss FILLER_0_9_223/a_36_472# FILLER_0_9_223/a_572_375#
+ FILLER_0_9_223/a_124_375# FILLER_0_9_223/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd _342_/VPW vdd vss _142_ _020_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_273_ vdd _273_/VPW vss _090_ state\[0\] vdd _273_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_411_ vdd _411_/VPW _000_ cal_itt\[0\] net58 vss net75 vdd _411_/a_2665_112# _411_/a_448_472#
+ _411_/a_796_472# _411_/a_36_151# _411_/a_1204_472# _411_/a_3041_156# _411_/a_1000_472#
+ _411_/a_1308_423# _411_/a_1456_156# _411_/a_1288_156# _411_/a_2248_156# _411_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout80 vdd fanout80/VPW vss net80 net81 vdd fanout80/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_325_ vdd _325_/VPW vdd vss _130_ _118_ _129_ _325_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd FILLER_0_10_78/VPW vdd vss FILLER_0_10_78/a_1380_472# FILLER_0_10_78/a_36_472#
+ FILLER_0_10_78/a_932_472# FILLER_0_10_78/a_572_375# FILLER_0_10_78/a_124_375# FILLER_0_10_78/a_1468_375#
+ FILLER_0_10_78/a_1020_375# FILLER_0_10_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_256_ vdd _256_/VPW _056_ _068_ vdd vss _077_ net4 _076_ _256_/a_36_68# _256_/a_1612_497#
+ _256_/a_2124_68# _256_/a_244_497# _256_/a_2960_68# _256_/a_3368_68# _256_/a_2552_68#
+ _256_/a_1164_497# _256_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ vdd _308_/VPW _058_ vdd vss _115_ trim_mask\[0\] _114_ _308_/a_848_380# _308_/a_1084_68#
+ _308_/a_124_24# _308_/a_1152_472# _308_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd FILLER_0_1_98/VPW vdd vss FILLER_0_1_98/a_36_472# FILLER_0_1_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ vdd _239_/VPW net41 vss vdd _065_ _239_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd FILLER_0_12_124/VPW vdd vss FILLER_0_12_124/a_36_472# FILLER_0_12_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd FILLER_0_8_107/VPW vdd vss FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 vdd output24/VPW ctlp[7] net24 vdd vss output24/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 vdd output35/VPW result[8] net35 vdd vss output35/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 vdd output46/VPW trimb[3] net46 vdd vss output46/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd FILLER_0_18_2/VPW vdd vss FILLER_0_18_2/a_1916_375# FILLER_0_18_2/a_1380_472#
+ FILLER_0_18_2/a_3260_375# FILLER_0_18_2/a_36_472# FILLER_0_18_2/a_932_472# FILLER_0_18_2/a_2812_375#
+ FILLER_0_18_2/a_2276_472# FILLER_0_18_2/a_1828_472# FILLER_0_18_2/a_3172_472# FILLER_0_18_2/a_572_375#
+ FILLER_0_18_2/a_2724_472# FILLER_0_18_2/a_124_375# FILLER_0_18_2/a_1468_375# FILLER_0_18_2/a_1020_375#
+ FILLER_0_18_2/a_484_472# FILLER_0_18_2/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 vdd output13/VPW ctln[6] net13 vdd vss output13/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd FILLER_0_7_162/VPW vdd vss FILLER_0_7_162/a_36_472# FILLER_0_7_162/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd FILLER_0_7_195/VPW vdd vss FILLER_0_7_195/a_36_472# FILLER_0_7_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vdd ANTENNA_input1_I/VPW vss cal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vdd ANTENNA__414__RN/VPW vss net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ vdd _341_/VPW _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ _341_/a_49_472#
+ _341_/a_665_69# _341_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _410_/VPW vdd _188_ _187_ _042_ _120_ vss _410_/a_36_68# _410_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ vdd _272_/VPW _089_ vdd vss _003_ _079_ _087_ _272_/a_36_472# _272_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vdd fanout70/VPW vss net70 net73 vdd fanout70/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ vdd _255_/VPW _076_ vss vdd _057_ _255_/a_224_552# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_324_ vdd _324_/VPW vdd vss _129_ calibrate _062_ _324_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output40_I vdd ANTENNA_output40_I/VPW vss net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 vdd fanout81/VPW vss net81 net82 vdd fanout81/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_55 vdd FILLER_0_19_55/VPW vdd vss FILLER_0_19_55/a_36_472# FILLER_0_19_55/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A1 vdd ANTENNA__304__A1/VPW vss _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_307_ vdd _307_/VPW vdd vss _114_ _113_ _096_ _307_/a_234_472# _307_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd _238_/VPW vdd vss _065_ trim_mask\[3\] trim_val\[3\] _238_/a_255_603# _238_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd FILLER_0_21_125/VPW vdd vss FILLER_0_21_125/a_36_472# FILLER_0_21_125/a_572_375#
+ FILLER_0_21_125/a_124_375# FILLER_0_21_125/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd FILLER_0_16_89/VPW vdd vss FILLER_0_16_89/a_1380_472# FILLER_0_16_89/a_36_472#
+ FILLER_0_16_89/a_932_472# FILLER_0_16_89/a_572_375# FILLER_0_16_89/a_124_375# FILLER_0_16_89/a_1468_375#
+ FILLER_0_16_89/a_1020_375# FILLER_0_16_89/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd FILLER_0_12_136/VPW vdd vss FILLER_0_12_136/a_1380_472# FILLER_0_12_136/a_36_472#
+ FILLER_0_12_136/a_932_472# FILLER_0_12_136/a_572_375# FILLER_0_12_136/a_124_375#
+ FILLER_0_12_136/a_1468_375# FILLER_0_12_136/a_1020_375# FILLER_0_12_136/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 vdd output25/VPW ctlp[8] net25 vdd vss output25/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 vdd output47/VPW trimb[4] net47 vdd vss output47/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 vdd output36/VPW result[9] net36 vdd vss output36/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 vdd output14/VPW ctln[7] net14 vdd vss output14/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd FILLER_0_4_144/VPW vdd vss FILLER_0_4_144/a_36_472# FILLER_0_4_144/a_572_375#
+ FILLER_0_4_144/a_124_375# FILLER_0_4_144/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd FILLER_0_4_177/VPW vdd vss FILLER_0_4_177/a_36_472# FILLER_0_4_177/a_572_375#
+ FILLER_0_4_177/a_124_375# FILLER_0_4_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vdd _340_/VPW vss _141_ _140_ vdd _340_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd _271_/VPW vdd vss cal_itt\[3\] _089_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vdd ANTENNA__356__B/VPW vss _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd FILLER_0_10_256/VPW vdd vss FILLER_0_10_256/a_36_472# FILLER_0_10_256/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__200__I vdd ANTENNA__200__I/VPW vss net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vdd ANTENNA_fanout52_I/VPW vss net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_99 vdd FILLER_0_4_99/VPW vdd vss FILLER_0_4_99/a_36_472# FILLER_0_4_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd FILLER_0_6_239/VPW vdd vss FILLER_0_6_239/a_36_472# FILLER_0_6_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout71 vdd fanout71/VPW vss net71 net73 vdd fanout71/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 vdd fanout60/VPW net60 vss vdd net61 fanout60/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_323_ vdd _323_/VPW vss _015_ _128_ vdd _323_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vdd fanout82/VPW vss net82 net2 vdd fanout82/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ vdd _254_/VPW _074_ vdd vss _075_ cal_itt\[3\] _072_ _254_/a_448_472# _254_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_237_ vdd _237_/VPW vdd vss net40 net45 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_306_ vdd _306_/VPW vss _113_ _057_ vdd _306_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_57 vdd FILLER_0_16_57/VPW vdd vss FILLER_0_16_57/a_1380_472# FILLER_0_16_57/a_36_472#
+ FILLER_0_16_57/a_932_472# FILLER_0_16_57/a_572_375# FILLER_0_16_57/a_124_375# FILLER_0_16_57/a_1468_375#
+ FILLER_0_16_57/a_1020_375# FILLER_0_16_57/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 vdd output26/VPW ctlp[9] net26 vdd vss output26/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 vdd output15/VPW ctln[8] net15 vdd vss output15/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 vdd output48/VPW valid net48 vdd vss output48/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 vdd output37/VPW sample net37 vdd vss output37/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd FILLER_0_17_218/VPW vdd vss FILLER_0_17_218/a_36_472# FILLER_0_17_218/a_572_375#
+ FILLER_0_17_218/a_124_375# FILLER_0_17_218/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd FILLER_0_4_123/VPW vdd vss FILLER_0_4_123/a_36_472# FILLER_0_4_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vdd ANTENNA__203__I/VPW vss net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ vdd _270_/VPW _088_ vdd vss _002_ _079_ _087_ _270_/a_36_472# _270_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd _399_/VPW vdd vss _179_ cal_count\[1\] _178_ _399_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ vdd _322_/VPW _127_ vdd vss _128_ _068_ _124_ _322_/a_848_380# _322_/a_1084_68#
+ _322_/a_124_24# _322_/a_1152_472# _322_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vdd fanout61/VPW vss net61 net62 vdd fanout61/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vdd fanout72/VPW vss net72 net74 vdd fanout72/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd FILLER_0_10_37/VPW vdd vss FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 vdd fanout50/VPW net50 vss vdd net52 fanout50/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_253_ vdd _253_/VPW cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] _253_/a_36_68#
+ _253_/a_1732_68# _253_/a_244_68# _253_/a_1100_68# _253_/a_1528_68# _253_/a_672_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_305_ vdd _305_/VPW vdd vss _112_ net1 _081_ _305_/a_36_159# vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ vdd _236_/VPW net40 vss vdd _064_ _236_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vdd ANTENNA__206__I/VPW vss net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd FILLER_0_20_193/VPW vdd vss FILLER_0_20_193/a_36_472# FILLER_0_20_193/a_572_375#
+ FILLER_0_20_193/a_124_375# FILLER_0_20_193/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vdd _219_/VPW vss _053_ trim_mask\[0\] vdd _219_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 vdd output27/VPW result[0] net27 vdd vss output27/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 vdd output16/VPW ctln[9] net16 vdd vss output16/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 vdd output38/VPW trim[0] net38 vdd vss output38/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd FILLER_0_16_241/VPW vdd vss FILLER_0_16_241/a_36_472# FILLER_0_16_241/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vdd _398_/VPW vss _178_ net3 vdd _398_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd FILLER_0_10_247/VPW vdd vss FILLER_0_10_247/a_36_472# FILLER_0_10_247/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_214 vdd FILLER_0_10_214/VPW vdd vss FILLER_0_10_214/a_36_472# FILLER_0_10_214/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_91 vdd FILLER_0_14_91/VPW vdd vss FILLER_0_14_91/a_36_472# FILLER_0_14_91/a_572_375#
+ FILLER_0_14_91/a_124_375# FILLER_0_14_91/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__209__I vdd ANTENNA__209__I/VPW vss net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I vdd ANTENNA_output19_I/VPW vss net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd FILLER_0_19_47/VPW vdd vss FILLER_0_19_47/a_36_472# FILLER_0_19_47/a_572_375#
+ FILLER_0_19_47/a_124_375# FILLER_0_19_47/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vdd fanout73/VPW vss net73 net74 vdd fanout73/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 vdd fanout62/VPW net62 vss vdd net64 fanout62/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vdd fanout51/VPW vss net51 net52 vdd fanout51/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ vdd _321_/VPW _076_ _125_ _126_ vdd vss _127_ _069_ _321_/a_2590_472# _321_/a_170_472#
+ _321_/a_1602_69# _321_/a_786_69# _321_/a_3126_472# _321_/a_1194_69# _321_/a_3662_472#
+ _321_/a_2034_472# _321_/a_358_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_252_ vdd _252_/VPW vdd vss cal_itt\[0\] _073_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_100 vdd FILLER_0_18_100/VPW vdd vss FILLER_0_18_100/a_36_472# FILLER_0_18_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd FILLER_0_18_177/VPW vdd vss FILLER_0_18_177/a_1916_375# FILLER_0_18_177/a_1380_472#
+ FILLER_0_18_177/a_3260_375# FILLER_0_18_177/a_36_472# FILLER_0_18_177/a_932_472#
+ FILLER_0_18_177/a_2812_375# FILLER_0_18_177/a_2276_472# FILLER_0_18_177/a_1828_472#
+ FILLER_0_18_177/a_3172_472# FILLER_0_18_177/a_572_375# FILLER_0_18_177/a_2724_472#
+ FILLER_0_18_177/a_124_375# FILLER_0_18_177/a_1468_375# FILLER_0_18_177/a_1020_375#
+ FILLER_0_18_177/a_484_472# FILLER_0_18_177/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd _304_/VPW vdd vss _013_ _093_ _111_ _304_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd _235_/VPW vdd vss _064_ trim_mask\[2\] trim_val\[2\] _235_/a_255_603# _235_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vdd _218_/VPW vss net16 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd FILLER_0_16_37/VPW vdd vss FILLER_0_16_37/a_36_472# FILLER_0_16_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 vdd output17/VPW ctlp[0] net17 vdd vss output17/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 vdd output28/VPW result[1] net28 vdd vss output28/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 vdd output39/VPW trim[1] net39 vdd vss output39/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd FILLER_0_13_212/VPW vdd vss FILLER_0_13_212/a_1380_472# FILLER_0_13_212/a_36_472#
+ FILLER_0_13_212/a_932_472# FILLER_0_13_212/a_572_375# FILLER_0_13_212/a_124_375#
+ FILLER_0_13_212/a_1468_375# FILLER_0_13_212/a_1020_375# FILLER_0_13_212/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ vdd _397_/VPW _177_ vdd vss _040_ _131_ _175_ _397_/a_36_472# _397_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd FILLER_0_14_81/VPW vdd vss FILLER_0_14_81/a_36_472# FILLER_0_14_81/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout63 vdd fanout63/VPW net63 vss vdd net64 fanout63/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_320_ vdd _320_/VPW _096_ vdd vss _126_ mask\[0\] _113_ _320_/a_1792_472# _320_/a_224_472#
+ _320_/a_1568_472# _320_/a_36_472# _320_/a_1120_472# _320_/a_672_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_28 vdd FILLER_0_10_28/VPW vdd vss FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 vdd fanout74/VPW vss net74 net82 vdd fanout74/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 vdd fanout52/VPW net52 vss vdd net57 fanout52/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ vdd _251_/VPW _072_ vdd vss net48 _068_ _070_ _251_/a_468_472# _251_/a_244_472#
+ _251_/a_1130_472# _251_/a_906_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_449_ vdd _449_/VPW _038_ en_co_clk net55 vss net72 vdd _449_/a_2665_112# _449_/a_448_472#
+ _449_/a_796_472# _449_/a_36_151# _449_/a_1204_472# _449_/a_3041_156# _449_/a_1000_472#
+ _449_/a_1308_423# _449_/a_1456_156# _449_/a_1288_156# _449_/a_2248_156# _449_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ vdd _303_/VPW net36 vdd vss _111_ mask\[9\] _098_ _303_/a_36_472# _303_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vdd _234_/VPW vss net44 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_217_ vdd _217_/VPW vss net26 _052_ vdd _217_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_181 vdd FILLER_0_14_181/VPW vdd vss FILLER_0_14_181/a_36_472# FILLER_0_14_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 vdd output18/VPW ctlp[1] net18 vdd vss output18/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 vdd output29/VPW result[2] net29 vdd vss output29/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vdd ANTENNA_fanout80_I/VPW vss net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd _396_/VPW vdd vss _177_ cal_count\[1\] _176_ _396_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout53 vdd fanout53/VPW net53 vss vdd net56 fanout53/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_250_ vdd _250_/VPW vss _072_ _071_ vdd _250_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 vdd fanout75/VPW vss net75 net76 vdd fanout75/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vdd fanout64/VPW vss net64 net65 vdd fanout64/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ vdd _448_/VPW _037_ trim_val\[4\] net59 vss net76 vdd _448_/a_2665_112# _448_/a_448_472#
+ _448_/a_796_472# _448_/a_36_151# _448_/a_1204_472# _448_/a_3041_156# _448_/a_1000_472#
+ _448_/a_1308_423# _448_/a_1456_156# _448_/a_1288_156# _448_/a_2248_156# _448_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ vdd _379_/VPW trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ _379_/a_36_472#
+ _379_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_302_ vdd _302_/VPW vdd vss _012_ _093_ _110_ _302_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd FILLER_0_21_28/VPW vdd vss FILLER_0_21_28/a_1916_375# FILLER_0_21_28/a_1380_472#
+ FILLER_0_21_28/a_3260_375# FILLER_0_21_28/a_36_472# FILLER_0_21_28/a_932_472# FILLER_0_21_28/a_2812_375#
+ FILLER_0_21_28/a_2276_472# FILLER_0_21_28/a_1828_472# FILLER_0_21_28/a_3172_472#
+ FILLER_0_21_28/a_572_375# FILLER_0_21_28/a_2724_472# FILLER_0_21_28/a_124_375# FILLER_0_21_28/a_1468_375#
+ FILLER_0_21_28/a_1020_375# FILLER_0_21_28/a_484_472# FILLER_0_21_28/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__216__A2 vdd ANTENNA__216__A2/VPW vss net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ vdd _233_/VPW vss net39 _063_ vdd _233_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd FILLER_0_15_116/VPW vdd vss FILLER_0_15_116/a_36_472# FILLER_0_15_116/a_572_375#
+ FILLER_0_15_116/a_124_375# FILLER_0_15_116/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vdd ANTENNA__373__A1/VPW vss cal_count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_216_ vdd _216_/VPW vdd vss _052_ mask\[9\] net36 _216_/a_255_603# _216_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_146 vdd FILLER_0_7_146/VPW vdd vss FILLER_0_7_146/a_36_472# FILLER_0_7_146/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 vdd output19/VPW ctlp[2] net19 vdd vss output19/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd FILLER_0_7_59/VPW vdd vss FILLER_0_7_59/a_36_472# FILLER_0_7_59/a_572_375#
+ FILLER_0_7_59/a_124_375# FILLER_0_7_59/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd FILLER_0_16_255/VPW vdd vss FILLER_0_16_255/a_36_472# FILLER_0_16_255/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd FILLER_0_0_130/VPW vdd vss FILLER_0_0_130/a_36_472# FILLER_0_0_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd FILLER_0_8_263/VPW vdd vss FILLER_0_8_263/a_36_472# FILLER_0_8_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd FILLER_0_14_50/VPW vdd vss FILLER_0_14_50/a_36_472# FILLER_0_14_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ vdd _395_/VPW _070_ _085_ vdd vss _176_ _116_ _072_ _395_/a_1492_488# _395_/a_244_68#
+ _395_/a_1044_488# _395_/a_636_68# _395_/a_36_488# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd FILLER_0_4_49/VPW vdd vss FILLER_0_4_49/a_36_472# FILLER_0_4_49/a_572_375#
+ FILLER_0_4_49/a_124_375# FILLER_0_4_49/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 vdd fanout54/VPW net54 vss vdd net56 fanout54/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vdd fanout76/VPW vss net76 net81 vdd fanout76/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vdd fanout65/VPW vss net65 net5 vdd fanout65/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd FILLER_0_19_28/VPW vdd vss FILLER_0_19_28/a_36_472# FILLER_0_19_28/a_572_375#
+ FILLER_0_19_28/a_124_375# FILLER_0_19_28/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ vdd _447_/VPW _036_ trim_val\[3\] net50 vss net68 vdd _447_/a_2665_112# _447_/a_448_472#
+ _447_/a_796_472# _447_/a_36_151# _447_/a_1204_472# _447_/a_3041_156# _447_/a_1000_472#
+ _447_/a_1308_423# _447_/a_1456_156# _447_/a_1288_156# _447_/a_2248_156# _447_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_2 vdd FILLER_0_3_2/VPW vdd vss FILLER_0_3_2/a_36_472# FILLER_0_3_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ vdd _378_/VPW vdd vss _033_ _160_ _165_ _378_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ vdd _301_/VPW net35 vdd vss _110_ mask\[8\] _098_ _301_/a_36_472# _301_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vdd ANTENNA_output17_I/VPW vss net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd _232_/VPW vdd vss _063_ trim_mask\[1\] trim_val\[1\] _232_/a_255_603# _232_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vdd _215_/VPW vss net15 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd FILLER_0_11_142/VPW vdd vss FILLER_0_11_142/a_36_472# FILLER_0_11_142/a_572_375#
+ FILLER_0_11_142/a_124_375# FILLER_0_11_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd FILLER_0_2_93/VPW vdd vss FILLER_0_2_93/a_36_472# FILLER_0_2_93/a_572_375#
+ FILLER_0_2_93/a_124_375# FILLER_0_2_93/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd FILLER_0_17_72/VPW vdd vss FILLER_0_17_72/a_1916_375# FILLER_0_17_72/a_1380_472#
+ FILLER_0_17_72/a_3260_375# FILLER_0_17_72/a_36_472# FILLER_0_17_72/a_932_472# FILLER_0_17_72/a_2812_375#
+ FILLER_0_17_72/a_2276_472# FILLER_0_17_72/a_1828_472# FILLER_0_17_72/a_3172_472#
+ FILLER_0_17_72/a_572_375# FILLER_0_17_72/a_2724_472# FILLER_0_17_72/a_124_375# FILLER_0_17_72/a_1468_375#
+ FILLER_0_17_72/a_1020_375# FILLER_0_17_72/a_484_472# FILLER_0_17_72/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd FILLER_0_3_172/VPW vdd vss FILLER_0_3_172/a_1916_375# FILLER_0_3_172/a_1380_472#
+ FILLER_0_3_172/a_3260_375# FILLER_0_3_172/a_36_472# FILLER_0_3_172/a_932_472# FILLER_0_3_172/a_2812_375#
+ FILLER_0_3_172/a_2276_472# FILLER_0_3_172/a_1828_472# FILLER_0_3_172/a_3172_472#
+ FILLER_0_3_172/a_572_375# FILLER_0_3_172/a_2724_472# FILLER_0_3_172/a_124_375# FILLER_0_3_172/a_1468_375#
+ FILLER_0_3_172/a_1020_375# FILLER_0_3_172/a_484_472# FILLER_0_3_172/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vdd ANTENNA_output47_I/VPW vss net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ vdd _394_/VPW _095_ vdd vss _175_ _174_ cal_count\[1\] _394_/a_244_524# _394_/a_2215_68#
+ _394_/a_56_524# _394_/a_718_524# _394_/a_728_93# _394_/a_1936_472# _394_/a_1336_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 vdd fanout55/VPW net55 vss vdd net57 fanout55/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd FILLER_0_5_212/VPW vdd vss FILLER_0_5_212/a_36_472# FILLER_0_5_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vdd fanout77/VPW vss net77 net78 vdd fanout77/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ vdd _446_/VPW _035_ trim_val\[2\] net49 vss net66 vdd _446_/a_2665_112# _446_/a_448_472#
+ _446_/a_796_472# _446_/a_36_151# _446_/a_1204_472# _446_/a_3041_156# _446_/a_1000_472#
+ _446_/a_1308_423# _446_/a_1456_156# _446_/a_1288_156# _446_/a_2248_156# _446_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout66 vdd fanout66/VPW vss net66 net68 vdd fanout66/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ vdd _377_/VPW trim_val\[0\] vdd vss _165_ _053_ _164_ _377_/a_36_472# _377_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd _300_/VPW vdd vss _011_ _104_ _109_ _300_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd _231_/VPW vdd vss net37 _059_ _062_ _231_/a_652_68# _231_/a_244_68# vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ vdd _429_/VPW _018_ mask\[0\] net62 vss net79 vdd _429_/a_2665_112# _429_/a_448_472#
+ _429_/a_796_472# _429_/a_36_151# _429_/a_1204_472# _429_/a_3041_156# _429_/a_1000_472#
+ _429_/a_1308_423# _429_/a_1456_156# _429_/a_1288_156# _429_/a_2248_156# _429_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vdd input1/VPW vss net1 cal vdd input1/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vdd _214_/VPW vss net25 _051_ vdd _214_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd FILLER_0_7_104/VPW vdd vss FILLER_0_7_104/a_1380_472# FILLER_0_7_104/a_36_472#
+ FILLER_0_7_104/a_932_472# FILLER_0_7_104/a_572_375# FILLER_0_7_104/a_124_375# FILLER_0_7_104/a_1468_375#
+ FILLER_0_7_104/a_1020_375# FILLER_0_7_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd FILLER_0_4_107/VPW vdd vss FILLER_0_4_107/a_1380_472# FILLER_0_4_107/a_36_472#
+ FILLER_0_4_107/a_932_472# FILLER_0_4_107/a_572_375# FILLER_0_4_107/a_124_375# FILLER_0_4_107/a_1468_375#
+ FILLER_0_4_107/a_1020_375# FILLER_0_4_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd FILLER_0_24_290/VPW vdd vss FILLER_0_24_290/a_36_472# FILLER_0_24_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd FILLER_0_15_290/VPW vdd vss FILLER_0_15_290/a_36_472# FILLER_0_15_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd FILLER_0_0_198/VPW vdd vss FILLER_0_0_198/a_36_472# FILLER_0_0_198/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd _393_/VPW vdd vss cal_count\[0\] _174_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vdd fanout78/VPW vss net78 net79 vdd fanout78/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vdd fanout56/VPW vss net56 net57 vdd fanout56/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vdd fanout67/VPW vss net67 net68 vdd fanout67/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ vdd _445_/VPW _034_ trim_val\[1\] net49 vss net66 vdd _445_/a_2665_112# _445_/a_448_472#
+ _445_/a_796_472# _445_/a_36_151# _445_/a_1204_472# _445_/a_3041_156# _445_/a_1000_472#
+ _445_/a_1308_423# _445_/a_1456_156# _445_/a_1288_156# _445_/a_2248_156# _445_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vdd _376_/VPW vss _164_ _163_ vdd _376_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd _230_/VPW vdd vss _062_ _060_ _061_ _230_/a_652_68# _230_/a_244_68# vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd FILLER_0_5_72/VPW vdd vss FILLER_0_5_72/a_1380_472# FILLER_0_5_72/a_36_472#
+ FILLER_0_5_72/a_932_472# FILLER_0_5_72/a_572_375# FILLER_0_5_72/a_124_375# FILLER_0_5_72/a_1468_375#
+ FILLER_0_5_72/a_1020_375# FILLER_0_5_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ vdd _428_/VPW _017_ state\[2\] net53 vss net70 vdd _428_/a_2665_112# _428_/a_448_472#
+ _428_/a_796_472# _428_/a_36_151# _428_/a_1204_472# _428_/a_3041_156# _428_/a_1000_472#
+ _428_/a_1308_423# _428_/a_1456_156# _428_/a_1288_156# _428_/a_2248_156# _428_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd FILLER_0_11_64/VPW vdd vss FILLER_0_11_64/a_36_472# FILLER_0_11_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ vdd _359_/VPW _131_ _129_ vdd vss _152_ _059_ _062_ _359_/a_1492_488# _359_/a_244_68#
+ _359_/a_1044_488# _359_/a_636_68# _359_/a_36_488# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vdd input2/VPW vss net2 clk vdd input2/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output22_I vdd ANTENNA_output22_I/VPW vss net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd _213_/VPW vdd vss _051_ mask\[8\] net35 _213_/a_255_603# _213_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_177 vdd FILLER_0_20_177/VPW vdd vss FILLER_0_20_177/a_1380_472# FILLER_0_20_177/a_36_472#
+ FILLER_0_20_177/a_932_472# FILLER_0_20_177/a_572_375# FILLER_0_20_177/a_124_375#
+ FILLER_0_20_177/a_1468_375# FILLER_0_20_177/a_1020_375# FILLER_0_20_177/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_206 vdd FILLER_0_13_206/VPW vdd vss FILLER_0_13_206/a_36_472# FILLER_0_13_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd FILLER_0_13_228/VPW vdd vss FILLER_0_13_228/a_36_472# FILLER_0_13_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _392_/VPW vdd _173_ _077_ _039_ cal_count\[0\] vss _392_/a_36_68# _392_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__282__I vdd ANTENNA__282__I/VPW vss _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 vdd fanout79/VPW vss net79 net81 vdd fanout79/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_2 vdd FILLER_0_12_2/VPW vdd vss FILLER_0_12_2/a_36_472# FILLER_0_12_2/a_572_375#
+ FILLER_0_12_2/a_124_375# FILLER_0_12_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout68 vdd fanout68/VPW vss net68 net69 vdd fanout68/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 vdd fanout57/VPW vss net57 net65 vdd fanout57/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ vdd _444_/VPW _033_ trim_val\[0\] net50 vss net67 vdd _444_/a_2665_112# _444_/a_448_472#
+ _444_/a_796_472# _444_/a_36_151# _444_/a_1204_472# _444_/a_3041_156# _444_/a_1000_472#
+ _444_/a_1308_423# _444_/a_1456_156# _444_/a_1288_156# _444_/a_2248_156# _444_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ vdd _375_/VPW _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] _375_/a_36_68# _375_/a_1612_497#
+ _375_/a_692_497# _375_/a_1388_497# _375_/a_960_497# vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__277__I vdd ANTENNA__277__I/VPW vss _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd FILLER_0_18_139/VPW vdd vss FILLER_0_18_139/a_1380_472# FILLER_0_18_139/a_36_472#
+ FILLER_0_18_139/a_932_472# FILLER_0_18_139/a_572_375# FILLER_0_18_139/a_124_375#
+ FILLER_0_18_139/a_1468_375# FILLER_0_18_139/a_1020_375# FILLER_0_18_139/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_161 vdd FILLER_0_17_161/VPW vdd vss FILLER_0_17_161/a_36_472# FILLER_0_17_161/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ vdd _427_/VPW _016_ state\[1\] net53 vdd vss net70 _427_/a_2665_112# _427_/a_448_472#
+ _427_/a_796_472# _427_/a_36_151# _427_/a_1204_472# _427_/a_3041_156# _427_/a_1000_472#
+ _427_/a_1308_423# _427_/a_2248_156# _427_/a_2560_156# vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_358_ vdd _358_/VPW vdd vss _053_ _151_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vdd ANTENNA__385__A2/VPW vss net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ vdd _289_/VPW net30 vdd vss _103_ mask\[3\] _099_ _289_/a_36_472# _289_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vdd input3/VPW vss net3 comp vdd input3/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vdd _212_/VPW vss net14 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vdd ANTENNA_output15_I/VPW vss net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd FILLER_0_22_86/VPW vdd vss FILLER_0_22_86/a_1380_472# FILLER_0_22_86/a_36_472#
+ FILLER_0_22_86/a_932_472# FILLER_0_22_86/a_572_375# FILLER_0_22_86/a_124_375# FILLER_0_22_86/a_1468_375#
+ FILLER_0_22_86/a_1020_375# FILLER_0_22_86/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd FILLER_0_11_101/VPW vdd vss FILLER_0_11_101/a_36_472# FILLER_0_11_101/a_572_375#
+ FILLER_0_11_101/a_124_375# FILLER_0_11_101/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd FILLER_0_17_64/VPW vdd vss FILLER_0_17_64/a_36_472# FILLER_0_17_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd FILLER_0_3_142/VPW vdd vss FILLER_0_3_142/a_36_472# FILLER_0_3_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd _391_/VPW vdd vss _173_ cal_count\[0\] _120_ _391_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 vdd fanout69/VPW vss net69 net74 vdd fanout69/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 vdd fanout58/VPW net58 vss vdd net59 fanout58/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_374_ vdd _374_/VPW vdd _061_ _056_ _162_ calibrate vss _374_/a_36_68# _374_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_443_ vdd _443_/VPW _032_ trim_mask\[4\] net52 vss net69 vdd _443_/a_2665_112# _443_/a_448_472#
+ _443_/a_796_472# _443_/a_36_151# _443_/a_1204_472# _443_/a_3041_156# _443_/a_1000_472#
+ _443_/a_1308_423# _443_/a_1456_156# _443_/a_1288_156# _443_/a_2248_156# _443_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_107 vdd FILLER_0_18_107/VPW vdd vss FILLER_0_18_107/a_1916_375# FILLER_0_18_107/a_1380_472#
+ FILLER_0_18_107/a_3260_375# FILLER_0_18_107/a_36_472# FILLER_0_18_107/a_932_472#
+ FILLER_0_18_107/a_2812_375# FILLER_0_18_107/a_2276_472# FILLER_0_18_107/a_1828_472#
+ FILLER_0_18_107/a_3172_472# FILLER_0_18_107/a_572_375# FILLER_0_18_107/a_2724_472#
+ FILLER_0_18_107/a_124_375# FILLER_0_18_107/a_1468_375# FILLER_0_18_107/a_1020_375#
+ FILLER_0_18_107/a_484_472# FILLER_0_18_107/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vdd ANTENNA__394__A3/VPW vss _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd _288_/VPW vdd vss _006_ _094_ _102_ _288_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd _357_/VPW vdd vss _150_ _027_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ vdd _426_/VPW _015_ state\[0\] net64 vss net81 vdd _426_/a_2665_112# _426_/a_448_472#
+ _426_/a_796_472# _426_/a_36_151# _426_/a_1204_472# _426_/a_3041_156# _426_/a_1000_472#
+ _426_/a_1308_423# _426_/a_1456_156# _426_/a_1288_156# _426_/a_2248_156# _426_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 vdd input4/VPW vss net4 en vdd input4/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_211_ vdd _211_/VPW vss net24 _050_ vdd _211_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd _409_/VPW vdd vss _188_ cal_count\[3\] _077_ _409_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd FILLER_0_11_135/VPW vdd vss FILLER_0_11_135/a_36_472# FILLER_0_11_135/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd FILLER_0_11_124/VPW vdd vss FILLER_0_11_124/a_36_472# FILLER_0_11_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd FILLER_0_15_282/VPW vdd vss FILLER_0_15_282/a_36_472# FILLER_0_15_282/a_572_375#
+ FILLER_0_15_282/a_124_375# FILLER_0_15_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vdd ANTENNA__413__RN/VPW vss net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ vdd _390_/VPW _136_ _172_ _067_ vdd vss _038_ _070_ _390_/a_36_68# _390_/a_244_472#
+ _390_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd FILLER_0_14_99/VPW vdd vss FILLER_0_14_99/a_36_472# FILLER_0_14_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 vdd fanout59/VPW net59 vss vdd net64 fanout59/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ vdd _373_/VPW _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ _373_/a_438_68#
+ _373_/a_244_68# _373_/a_1254_68# _373_/a_1060_68# _373_/a_632_68# _373_/a_1458_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ vdd _442_/VPW _031_ trim_mask\[3\] net52 vss net69 vdd _442_/a_2665_112# _442_/a_448_472#
+ _442_/a_796_472# _442_/a_36_151# _442_/a_1204_472# _442_/a_3041_156# _442_/a_1000_472#
+ _442_/a_1308_423# _442_/a_1456_156# _442_/a_1288_156# _442_/a_2248_156# _442_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_356_ vdd _356_/VPW _093_ vdd vss _150_ mask\[9\] _136_ _356_/a_36_472# _356_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_287_ vdd _287_/VPW net29 vdd vss _102_ mask\[2\] _099_ _287_/a_36_472# _287_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd FILLER_0_11_78/VPW vdd vss FILLER_0_11_78/a_36_472# FILLER_0_11_78/a_572_375#
+ FILLER_0_11_78/a_124_375# FILLER_0_11_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vdd input5/VPW vss net5 rstn vdd input5/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ vdd _425_/VPW _014_ calibrate net58 vss net75 vdd _425_/a_2665_112# _425_/a_448_472#
+ _425_/a_796_472# _425_/a_36_151# _425_/a_1204_472# _425_/a_3041_156# _425_/a_1000_472#
+ _425_/a_1308_423# _425_/a_1456_156# _425_/a_1288_156# _425_/a_2248_156# _425_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd _210_/VPW vdd vss _050_ mask\[7\] net34 _210_/a_255_603# _210_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd FILLER_0_20_169/VPW vdd vss FILLER_0_20_169/a_36_472# FILLER_0_20_169/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ vdd _408_/VPW _186_ vdd vss _187_ _095_ cal_count\[3\] _408_/a_244_524# _408_/a_2215_68#
+ _408_/a_56_524# _408_/a_718_524# _408_/a_728_93# _408_/a_1936_472# _408_/a_1336_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vdd _339_/VPW vss _140_ _091_ vdd _339_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vdd ANTENNA_output20_I/VPW vss net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd FILLER_0_21_286/VPW vdd vss FILLER_0_21_286/a_36_472# FILLER_0_21_286/a_572_375#
+ FILLER_0_21_286/a_124_375# FILLER_0_21_286/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd FILLER_0_12_220/VPW vdd vss FILLER_0_12_220/a_1380_472# FILLER_0_12_220/a_36_472#
+ FILLER_0_12_220/a_932_472# FILLER_0_12_220/a_572_375# FILLER_0_12_220/a_124_375#
+ FILLER_0_12_220/a_1468_375# FILLER_0_12_220/a_1020_375# FILLER_0_12_220/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd FILLER_0_8_247/VPW vdd vss FILLER_0_8_247/a_1380_472# FILLER_0_8_247/a_36_472#
+ FILLER_0_8_247/a_932_472# FILLER_0_8_247/a_572_375# FILLER_0_8_247/a_124_375# FILLER_0_8_247/a_1468_375#
+ FILLER_0_8_247/a_1020_375# FILLER_0_8_247/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 vdd fanout49/VPW net49 vss vdd net50 fanout49/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_206 vdd FILLER_0_5_206/VPW vdd vss FILLER_0_5_206/a_36_472# FILLER_0_5_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ vdd _441_/VPW _030_ trim_mask\[2\] net49 vss net66 vdd _441_/a_2665_112# _441_/a_448_472#
+ _441_/a_796_472# _441_/a_36_151# _441_/a_1204_472# _441_/a_3041_156# _441_/a_1000_472#
+ _441_/a_1308_423# _441_/a_1456_156# _441_/a_1288_156# _441_/a_2248_156# _441_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_372_ vdd _372_/VPW _070_ _076_ _068_ vdd vss _160_ _133_ _372_/a_2590_472# _372_/a_170_472#
+ _372_/a_1602_69# _372_/a_786_69# _372_/a_3126_472# _372_/a_1194_69# _372_/a_3662_472#
+ _372_/a_2034_472# _372_/a_358_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__303__A2 vdd ANTENNA__303__A2/VPW vss _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd FILLER_0_17_142/VPW vdd vss FILLER_0_17_142/a_36_472# FILLER_0_17_142/a_572_375#
+ FILLER_0_17_142/a_124_375# FILLER_0_17_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_54 vdd FILLER_0_5_54/VPW vdd vss FILLER_0_5_54/a_1380_472# FILLER_0_5_54/a_36_472#
+ FILLER_0_5_54/a_932_472# FILLER_0_5_54/a_572_375# FILLER_0_5_54/a_124_375# FILLER_0_5_54/a_1468_375#
+ FILLER_0_5_54/a_1020_375# FILLER_0_5_54/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_355_ vdd _355_/VPW vdd vss _149_ _026_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ vdd _424_/VPW _013_ net36 net55 vss net72 vdd _424_/a_2665_112# _424_/a_448_472#
+ _424_/a_796_472# _424_/a_36_151# _424_/a_1204_472# _424_/a_3041_156# _424_/a_1000_472#
+ _424_/a_1308_423# _424_/a_1456_156# _424_/a_1288_156# _424_/a_2248_156# _424_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ vdd _286_/VPW vdd vss _005_ _094_ _101_ _286_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_123 vdd FILLER_0_14_123/VPW vdd vss FILLER_0_14_123/a_36_472# FILLER_0_14_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd _338_/VPW vdd vss _139_ _019_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ vdd _407_/VPW _185_ vdd vss _186_ _181_ _184_ _407_/a_36_472# _407_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ vdd _269_/VPW cal_itt\[2\] vdd vss _088_ _083_ _078_ _269_/a_36_472# _269_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd FILLER_0_17_56/VPW vdd vss FILLER_0_17_56/a_36_472# FILLER_0_17_56/a_572_375#
+ FILLER_0_17_56/a_124_375# FILLER_0_17_56/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vdd ANTENNA_input4_I/VPW vss en vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vdd _371_/VPW vss _032_ _159_ vdd _371_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ vdd _440_/VPW _029_ trim_mask\[1\] net49 vss net66 vdd _440_/a_2665_112# _440_/a_448_472#
+ _440_/a_796_472# _440_/a_36_151# _440_/a_1204_472# _440_/a_3041_156# _440_/a_1000_472#
+ _440_/a_1308_423# _440_/a_1456_156# _440_/a_1288_156# _440_/a_2248_156# _440_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd FILLER_0_5_88/VPW vdd vss FILLER_0_5_88/a_36_472# FILLER_0_5_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ vdd _423_/VPW _012_ net35 net55 vss net72 vdd _423_/a_2665_112# _423_/a_448_472#
+ _423_/a_796_472# _423_/a_36_151# _423_/a_1204_472# _423_/a_3041_156# _423_/a_1000_472#
+ _423_/a_1308_423# _423_/a_1456_156# _423_/a_1288_156# _423_/a_2248_156# _423_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ vdd _354_/VPW _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ _354_/a_49_472#
+ _354_/a_665_69# _354_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_285_ vdd _285_/VPW net28 vdd vss _101_ mask\[1\] _099_ _285_/a_36_472# _285_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_199_ vdd _199_/VPW net20 vss vdd _046_ _199_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ vdd _337_/VPW _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ _337_/a_49_472#
+ _337_/a_665_69# _337_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd _406_/VPW vdd vss _185_ _178_ cal_count\[2\] _406_/a_36_159# vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd _268_/VPW vdd vss _087_ _086_ _074_ _268_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd FILLER_0_24_274/VPW vdd vss FILLER_0_24_274/a_1380_472# FILLER_0_24_274/a_36_472#
+ FILLER_0_24_274/a_932_472# FILLER_0_24_274/a_572_375# FILLER_0_24_274/a_124_375#
+ FILLER_0_24_274/a_1468_375# FILLER_0_24_274/a_1020_375# FILLER_0_24_274/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ vdd _370_/VPW _152_ vdd vss _159_ trim_mask\[4\] _081_ _370_/a_848_380# _370_/a_1084_68#
+ _370_/a_124_24# _370_/a_1152_472# _370_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vdd ANTENNA_fanout55_I/VPW vss net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd FILLER_0_1_266/VPW vdd vss FILLER_0_1_266/a_36_472# FILLER_0_1_266/a_572_375#
+ FILLER_0_1_266/a_124_375# FILLER_0_1_266/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_422_ vdd _422_/VPW _011_ net34 net61 vss net78 vdd _422_/a_2665_112# _422_/a_448_472#
+ _422_/a_796_472# _422_/a_36_151# _422_/a_1204_472# _422_/a_3041_156# _422_/a_1000_472#
+ _422_/a_1308_423# _422_/a_1456_156# _422_/a_1288_156# _422_/a_2248_156# _422_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_353_ vdd _353_/VPW vdd vss _148_ _025_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd FILLER_0_17_133/VPW vdd vss FILLER_0_17_133/a_36_472# FILLER_0_17_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output36_I vdd ANTENNA_output36_I/VPW vss net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_284_ vdd _284_/VPW vdd vss _004_ _094_ _100_ _284_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_198_ vdd _198_/VPW vdd vss _046_ mask\[3\] net30 _198_/a_255_603# _198_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_336_ vdd _336_/VPW vdd vss _138_ _018_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_405_ vdd _405_/VPW vdd vss _184_ _178_ cal_count\[2\] _405_/a_255_603# _405_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ vdd _267_/VPW _071_ vdd vss _086_ _085_ state\[1\] _267_/a_1792_472# _267_/a_224_472#
+ _267_/a_1568_472# _267_/a_36_472# _267_/a_1120_472# _267_/a_672_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd FILLER_0_6_177/VPW vdd vss FILLER_0_6_177/a_36_472# FILLER_0_6_177/a_572_375#
+ FILLER_0_6_177/a_124_375# FILLER_0_6_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd _319_/VPW vdd vss _125_ _058_ _119_ _319_/a_234_472# _319_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd FILLER_0_8_239/VPW vdd vss FILLER_0_8_239/a_36_472# FILLER_0_8_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd FILLER_0_1_212/VPW vdd vss FILLER_0_1_212/a_36_472# FILLER_0_1_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ vdd _421_/VPW _010_ net33 net60 vss net77 vdd _421_/a_2665_112# _421_/a_448_472#
+ _421_/a_796_472# _421_/a_36_151# _421_/a_1204_472# _421_/a_3041_156# _421_/a_1000_472#
+ _421_/a_1308_423# _421_/a_1456_156# _421_/a_1288_156# _421_/a_2248_156# _421_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_352_ vdd _352_/VPW _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ _352_/a_49_472#
+ _352_/a_665_69# _352_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_283_ vdd _283_/VPW net27 vdd vss _100_ mask\[0\] _099_ _283_/a_36_472# _283_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vdd FILLER_0_9_142/VPW vdd vss FILLER_0_9_142/a_36_472# FILLER_0_9_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd FILLER_0_20_107/VPW vdd vss FILLER_0_20_107/a_36_472# FILLER_0_20_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ vdd _404_/VPW _183_ vdd vss _041_ _131_ _182_ _404_/a_36_472# _404_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_335_ vdd _335_/VPW _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ _335_/a_49_472#
+ _335_/a_665_69# _335_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_266_ vdd _266_/VPW vdd vss _055_ _085_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_197_ vdd _197_/VPW vdd vss net19 net9 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vdd _249_/VPW vss _071_ state\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vdd ANTENNA__409__A1/VPW vss cal_count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd _318_/VPW vdd vss _124_ _115_ _118_ _318_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd FILLER_0_8_24/VPW vdd vss FILLER_0_8_24/a_36_472# FILLER_0_8_24/a_572_375#
+ FILLER_0_8_24/a_124_375# FILLER_0_8_24/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vdd ANTENNA__251__A2/VPW vss _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd FILLER_0_8_2/VPW vdd vss FILLER_0_8_2/a_36_472# FILLER_0_8_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vdd ANTENNA_input2_I/VPW vss clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ vdd _420_/VPW _009_ net32 net60 vss net77 vdd _420_/a_2665_112# _420_/a_448_472#
+ _420_/a_796_472# _420_/a_36_151# _420_/a_1204_472# _420_/a_3041_156# _420_/a_1000_472#
+ _420_/a_1308_423# _420_/a_1456_156# _420_/a_1288_156# _420_/a_2248_156# _420_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd _351_/VPW vdd vss _147_ _024_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vdd _282_/VPW vss _099_ _098_ vdd _282_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vdd ANTENNA__390__A1/VPW vss _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_334_ vdd _334_/VPW vss _137_ _132_ vdd _334_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_403_ vdd _403_/VPW vdd vss _183_ cal_count\[2\] _176_ _403_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vdd ANTENNA_output41_I/VPW vss net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd FILLER_0_6_90/VPW vdd vss FILLER_0_6_90/a_36_472# FILLER_0_6_90/a_572_375#
+ FILLER_0_6_90/a_124_375# FILLER_0_6_90/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ vdd _196_/VPW net19 vss vdd _045_ _196_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ vdd _265_/VPW _084_ _079_ _082_ vdd vss _001_ _081_ _083_ _265_/a_468_472#
+ _265_/a_224_472# _265_/a_244_68# _265_/a_916_472# vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vdd ANTENNA__395__B/VPW vss _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd FILLER_0_17_38/VPW vdd vss FILLER_0_17_38/a_36_472# FILLER_0_17_38/a_572_375#
+ FILLER_0_17_38/a_124_375# FILLER_0_17_38/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_248_ vdd _248_/VPW vss _070_ _069_ vdd _248_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__409__A2 vdd ANTENNA__409__A2/VPW vss _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vdd _317_/VPW vss _014_ _123_ vdd _317_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd FILLER_0_2_171/VPW vdd vss FILLER_0_2_171/a_36_472# FILLER_0_2_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd FILLER_0_12_236/VPW vdd vss FILLER_0_12_236/a_36_472# FILLER_0_12_236/a_572_375#
+ FILLER_0_12_236/a_124_375# FILLER_0_12_236/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ vdd _350_/VPW _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ _350_/a_49_472#
+ _350_/a_665_69# _350_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd _281_/VPW vdd vss _098_ _091_ _097_ _281_/a_234_472# _281_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vdd ANTENNA__237__I/VPW vss net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vdd _333_/VPW vss _136_ _091_ vdd _333_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd _195_/VPW vdd vss _045_ mask\[2\] net29 _195_/a_255_603# _195_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ vdd _402_/VPW _181_ vdd vss _182_ _095_ cal_count\[2\] _402_/a_244_567# _402_/a_718_527#
+ _402_/a_2172_497# _402_/a_56_567# _402_/a_1948_68# _402_/a_728_93# _402_/a_1296_93#
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd FILLER_0_11_109/VPW vdd vss FILLER_0_11_109/a_36_472# FILLER_0_11_109/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd _264_/VPW vdd vss _084_ cal_itt\[0\] cal_itt\[1\] _264_/a_224_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vdd ANTENNA__372__A2/VPW vss _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd FILLER_0_12_50/VPW vdd vss FILLER_0_12_50/a_36_472# FILLER_0_12_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ vdd _247_/VPW _069_ vss vdd _060_ _247_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ vdd _316_/VPW _122_ vdd vss _123_ _112_ calibrate _316_/a_848_380# _316_/a_1084_68#
+ _316_/a_124_24# _316_/a_1152_472# _316_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_60 vdd FILLER_0_23_60/VPW vdd vss FILLER_0_23_60/a_36_472# FILLER_0_23_60/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd FILLER_0_15_212/VPW vdd vss FILLER_0_15_212/a_1380_472# FILLER_0_15_212/a_36_472#
+ FILLER_0_15_212/a_932_472# FILLER_0_15_212/a_572_375# FILLER_0_15_212/a_124_375#
+ FILLER_0_15_212/a_1468_375# FILLER_0_15_212/a_1020_375# FILLER_0_15_212/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd FILLER_0_8_37/VPW vdd vss FILLER_0_8_37/a_36_472# FILLER_0_8_37/a_572_375#
+ FILLER_0_8_37/a_124_375# FILLER_0_8_37/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd FILLER_0_17_104/VPW vdd vss FILLER_0_17_104/a_1380_472# FILLER_0_17_104/a_36_472#
+ FILLER_0_17_104/a_932_472# FILLER_0_17_104/a_572_375# FILLER_0_17_104/a_124_375#
+ FILLER_0_17_104/a_1468_375# FILLER_0_17_104/a_1020_375# FILLER_0_17_104/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_72 vdd FILLER_0_15_72/VPW vdd vss FILLER_0_15_72/a_36_472# FILLER_0_15_72/a_572_375#
+ FILLER_0_15_72/a_124_375# FILLER_0_15_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd FILLER_0_1_204/VPW vdd vss FILLER_0_1_204/a_36_472# FILLER_0_1_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd _280_/VPW vdd vss _097_ _095_ _096_ _280_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd FILLER_0_14_107/VPW vdd vss FILLER_0_14_107/a_1380_472# FILLER_0_14_107/a_36_472#
+ FILLER_0_14_107/a_932_472# FILLER_0_14_107/a_572_375# FILLER_0_14_107/a_124_375#
+ FILLER_0_14_107/a_1468_375# FILLER_0_14_107/a_1020_375# FILLER_0_14_107/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ vdd _401_/VPW vdd _180_ _179_ _181_ _174_ vss _401_/a_36_68# _401_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_332_ vdd _332_/VPW _126_ vdd vss _017_ _127_ _135_ _332_/a_36_472# _332_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_194_ vdd _194_/VPW vss net8 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd _263_/VPW vdd vss _083_ _073_ _082_ _263_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd FILLER_0_5_181/VPW vdd vss FILLER_0_5_181/a_36_472# FILLER_0_5_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_246_ vdd _246_/VPW vss _068_ _055_ vdd _246_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_315_ vdd _315_/VPW _118_ _122_ _115_ _120_ _121_ vdd vss _315_/a_36_68# _315_/a_244_497#
+ _315_/a_1657_68# _315_/a_1229_68# _315_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_290 vdd FILLER_0_23_290/VPW vdd vss FILLER_0_23_290/a_36_472# FILLER_0_23_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd FILLER_0_15_235/VPW vdd vss FILLER_0_15_235/a_36_472# FILLER_0_15_235/a_572_375#
+ FILLER_0_15_235/a_124_375# FILLER_0_15_235/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd _229_/VPW vdd vss _061_ _055_ _057_ _229_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd FILLER_0_18_61/VPW vdd vss FILLER_0_18_61/a_36_472# FILLER_0_18_61/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd FILLER_0_11_282/VPW vdd vss FILLER_0_11_282/a_36_472# FILLER_0_11_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vdd ANTENNA_fanout76_I/VPW vss net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd FILLER_0_4_213/VPW vdd vss FILLER_0_4_213/a_36_472# FILLER_0_4_213/a_572_375#
+ FILLER_0_4_213/a_124_375# FILLER_0_4_213/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ vdd _400_/VPW vdd vss _180_ cal_count\[1\] _178_ _400_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_193_ vdd _193_/VPW net18 vss vdd _044_ _193_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_331_ vdd _331_/VPW _134_ vdd vss _135_ _086_ _132_ _331_/a_448_472# _331_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd _262_/VPW vdd vss cal_itt\[1\] _082_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vdd ANTENNA__303__B/VPW vss net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ vdd _314_/VPW vdd vss _121_ _085_ _069_ _314_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_245_ vdd _245_/VPW vdd vss net6 _067_ net67 _245_/a_234_472# _245_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_206 vdd FILLER_0_21_206/VPW vdd vss FILLER_0_21_206/a_36_472# FILLER_0_21_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vdd _228_/VPW vss _060_ state\[1\] vdd _228_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd FILLER_0_7_233/VPW vdd vss FILLER_0_7_233/a_36_472# FILLER_0_7_233/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd FILLER_0_9_60/VPW vdd vss FILLER_0_9_60/a_36_472# FILLER_0_9_60/a_572_375#
+ FILLER_0_9_60/a_124_375# FILLER_0_9_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd FILLER_0_13_142/VPW vdd vss FILLER_0_13_142/a_1380_472# FILLER_0_13_142/a_36_472#
+ FILLER_0_13_142/a_932_472# FILLER_0_13_142/a_572_375# FILLER_0_13_142/a_124_375#
+ FILLER_0_13_142/a_1468_375# FILLER_0_13_142/a_1020_375# FILLER_0_13_142/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ vdd _192_/VPW vdd vss _044_ mask\[1\] net28 _192_/a_255_603# _192_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_261_ vdd _261_/VPW vss _081_ _059_ vdd _261_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_330_ vdd _330_/VPW vdd vss _134_ _133_ _062_ _330_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd FILLER_0_12_20/VPW vdd vss FILLER_0_12_20/a_36_472# FILLER_0_12_20/a_572_375#
+ FILLER_0_12_20/a_124_375# FILLER_0_12_20/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd FILLER_0_5_172/VPW vdd vss FILLER_0_5_172/a_36_472# FILLER_0_5_172/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ vdd _244_/VPW vdd vss en_co_clk _067_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__190__I vdd ANTENNA__190__I/VPW vss _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_313_ vdd _313_/VPW vdd vss _120_ _059_ _119_ _313_/a_255_603# _313_/a_67_603# vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__257__A1 vdd ANTENNA__257__A1/VPW vss _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vdd _227_/VPW vss _059_ _058_ vdd _227_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vdd ANTENNA__402__A1/VPW vss _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd FILLER_0_20_31/VPW vdd vss FILLER_0_20_31/a_36_472# FILLER_0_20_31/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd FILLER_0_9_72/VPW vdd vss FILLER_0_9_72/a_1380_472# FILLER_0_9_72/a_36_472#
+ FILLER_0_9_72/a_932_472# FILLER_0_9_72/a_572_375# FILLER_0_9_72/a_124_375# FILLER_0_9_72/a_1468_375#
+ FILLER_0_9_72/a_1020_375# FILLER_0_9_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd FILLER_0_0_96/VPW vdd vss FILLER_0_0_96/a_36_472# FILLER_0_0_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _260_/VPW vdd _080_ _079_ _000_ _073_ vss _260_/a_36_68# _260_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ vdd _389_/VPW _171_ vdd vss _172_ _115_ _120_ _389_/a_428_148# _389_/a_36_148#
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd _191_/VPW vdd vss net17 net7 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd _312_/VPW vdd vss _119_ cal_itt\[3\] _074_ _312_/a_234_472# _312_/a_672_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd _243_/VPW vdd vss net47 net42 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd FILLER_0_23_282/VPW vdd vss FILLER_0_23_282/a_36_472# FILLER_0_23_282/a_572_375#
+ FILLER_0_23_282/a_124_375# FILLER_0_23_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd FILLER_0_15_205/VPW vdd vss FILLER_0_15_205/a_36_472# FILLER_0_15_205/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd FILLER_0_2_165/VPW vdd vss FILLER_0_2_165/a_36_472# FILLER_0_2_165/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd FILLER_0_18_53/VPW vdd vss FILLER_0_18_53/a_36_472# FILLER_0_18_53/a_572_375#
+ FILLER_0_18_53/a_124_375# FILLER_0_18_53/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ vdd _226_/VPW _057_ vdd vss _058_ _055_ _056_ _226_/a_1044_68# _226_/a_452_68#
+ _226_/a_276_68# _226_/a_860_68# vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vdd ANTENNA__426__CLK/VPW vss net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_98 vdd FILLER_0_20_98/VPW vdd vss FILLER_0_20_98/a_36_472# FILLER_0_20_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_87 vdd FILLER_0_20_87/VPW vdd vss FILLER_0_20_87/a_36_472# FILLER_0_20_87/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd _209_/VPW vdd vss net23 net13 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd FILLER_0_19_171/VPW vdd vss FILLER_0_19_171/a_1380_472# FILLER_0_19_171/a_36_472#
+ FILLER_0_19_171/a_932_472# FILLER_0_19_171/a_572_375# FILLER_0_19_171/a_124_375#
+ FILLER_0_19_171/a_1468_375# FILLER_0_19_171/a_1020_375# FILLER_0_19_171/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vdd ANTENNA__302__A1/VPW vss _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd FILLER_0_15_10/VPW vdd vss FILLER_0_15_10/a_36_472# FILLER_0_15_10/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd FILLER_0_15_2/VPW vdd vss FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_572_375#
+ FILLER_0_15_2/a_124_375# FILLER_0_15_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd FILLER_0_22_177/VPW vdd vss FILLER_0_22_177/a_1380_472# FILLER_0_22_177/a_36_472#
+ FILLER_0_22_177/a_932_472# FILLER_0_22_177/a_572_375# FILLER_0_22_177/a_124_375#
+ FILLER_0_22_177/a_1468_375# FILLER_0_22_177/a_1020_375# FILLER_0_22_177/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd FILLER_0_13_100/VPW vdd vss FILLER_0_13_100/a_36_472# FILLER_0_13_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd FILLER_0_9_105/VPW vdd vss FILLER_0_9_105/a_36_472# FILLER_0_9_105/a_572_375#
+ FILLER_0_9_105/a_124_375# FILLER_0_9_105/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ vdd _190_/VPW net17 vss vdd _043_ _190_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd _388_/VPW vdd vss _126_ _171_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vdd ANTENNA_output18_I/VPW vss net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ vdd _311_/VPW _114_ _117_ vdd vss _118_ _116_ _086_ _311_/a_692_473# _311_/a_254_473#
+ _311_/a_66_473# _311_/a_2700_473# _311_/a_1660_473# _311_/a_3220_473# _311_/a_1212_473#
+ _311_/a_2180_473# _311_/a_3740_473# _311_/a_1920_473# vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_242_ vdd _242_/VPW net47 vss vdd _066_ _242_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_228 vdd FILLER_0_15_228/VPW vdd vss FILLER_0_15_228/a_36_472# FILLER_0_15_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd FILLER_0_2_111/VPW vdd vss FILLER_0_2_111/a_1380_472# FILLER_0_2_111/a_36_472#
+ FILLER_0_2_111/a_932_472# FILLER_0_2_111/a_572_375# FILLER_0_2_111/a_124_375# FILLER_0_2_111/a_1468_375#
+ FILLER_0_2_111/a_1020_375# FILLER_0_2_111/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd FILLER_0_2_177/VPW vdd vss FILLER_0_2_177/a_36_472# FILLER_0_2_177/a_572_375#
+ FILLER_0_2_177/a_124_375# FILLER_0_2_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vdd _225_/VPW vss _057_ state\[2\] vdd _225_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd FILLER_0_18_76/VPW vdd vss FILLER_0_18_76/a_36_472# FILLER_0_18_76/a_572_375#
+ FILLER_0_18_76/a_124_375# FILLER_0_18_76/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ vdd _208_/VPW net23 vss vdd _049_ _208_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vdd _387_/VPW vss _037_ _170_ vdd _387_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_310_ vdd _310_/VPW _090_ vdd vss _117_ _060_ _113_ _310_/a_49_472# _310_/a_1133_69#
+ _310_/a_741_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_164 vdd FILLER_0_5_164/VPW vdd vss FILLER_0_5_164/a_36_472# FILLER_0_5_164/a_572_375#
+ FILLER_0_5_164/a_124_375# FILLER_0_5_164/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd FILLER_0_23_88/VPW vdd vss FILLER_0_23_88/a_36_472# FILLER_0_23_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd FILLER_0_23_44/VPW vdd vss FILLER_0_23_44/a_1380_472# FILLER_0_23_44/a_36_472#
+ FILLER_0_23_44/a_932_472# FILLER_0_23_44/a_572_375# FILLER_0_23_44/a_124_375# FILLER_0_23_44/a_1468_375#
+ FILLER_0_23_44/a_1020_375# FILLER_0_23_44/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd _241_/VPW vdd vss _066_ trim_mask\[4\] trim_val\[4\] _241_/a_224_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ vdd _439_/VPW _028_ trim_mask\[0\] net50 vss net67 vdd _439_/a_2665_112# _439_/a_448_472#
+ _439_/a_796_472# _439_/a_36_151# _439_/a_1204_472# _439_/a_3041_156# _439_/a_1000_472#
+ _439_/a_1308_423# _439_/a_1456_156# _439_/a_1288_156# _439_/a_2248_156# _439_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd FILLER_0_2_101/VPW vdd vss FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd FILLER_0_3_54/VPW vdd vss FILLER_0_3_54/a_36_472# FILLER_0_3_54/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vdd _224_/VPW vss _056_ state\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd _207_/VPW vdd vss _049_ mask\[6\] net33 _207_/a_255_603# _207_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd FILLER_0_19_195/VPW vdd vss FILLER_0_19_195/a_36_472# FILLER_0_19_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd FILLER_0_0_232/VPW vdd vss FILLER_0_0_232/a_36_472# FILLER_0_0_232/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd FILLER_0_16_154/VPW vdd vss FILLER_0_16_154/a_1380_472# FILLER_0_16_154/a_36_472#
+ FILLER_0_16_154/a_932_472# FILLER_0_16_154/a_572_375# FILLER_0_16_154/a_124_375#
+ FILLER_0_16_154/a_1468_375# FILLER_0_16_154/a_1020_375# FILLER_0_16_154/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vdd ANTENNA__257__B/VPW vss _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vdd ANTENNA__220__A2/VPW vss _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd FILLER_0_20_2/VPW vdd vss FILLER_0_20_2/a_36_472# FILLER_0_20_2/a_572_375#
+ FILLER_0_20_2/a_124_375# FILLER_0_20_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ vdd _386_/VPW _163_ vdd vss _170_ trim_val\[4\] _169_ _386_/a_848_380# _386_/a_1084_68#
+ _386_/a_124_24# _386_/a_1152_472# _386_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd FILLER_0_5_198/VPW vdd vss FILLER_0_5_198/a_36_472# FILLER_0_5_198/a_572_375#
+ FILLER_0_5_198/a_124_375# FILLER_0_5_198/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_240_ vdd _240_/VPW vdd vss net41 net46 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_282 vdd FILLER_0_17_282/VPW vdd vss FILLER_0_17_282/a_36_472# FILLER_0_17_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_274 vdd FILLER_0_23_274/VPW vdd vss FILLER_0_23_274/a_36_472# FILLER_0_23_274/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ vdd _438_/VPW _027_ mask\[9\] net54 vss net71 vdd _438_/a_2665_112# _438_/a_448_472#
+ _438_/a_796_472# _438_/a_36_151# _438_/a_1204_472# _438_/a_3041_156# _438_/a_1000_472#
+ _438_/a_1308_423# _438_/a_1456_156# _438_/a_1288_156# _438_/a_2248_156# _438_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ vdd _369_/VPW _153_ _154_ _158_ vdd vss _031_ _157_ _369_/a_36_68# _369_/a_244_472#
+ _369_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vdd ANTENNA_output23_I/VPW vss net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd FILLER_0_14_263/VPW vdd vss FILLER_0_14_263/a_36_472# FILLER_0_14_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ vdd _223_/VPW _055_ vss vdd state\[0\] _223_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd FILLER_0_9_290/VPW vdd vss FILLER_0_9_290/a_36_472# FILLER_0_9_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd _206_/VPW vdd vss net22 net12 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd FILLER_0_0_266/VPW vdd vss FILLER_0_0_266/a_36_472# FILLER_0_0_266/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd _385_/VPW vdd net37 net47 _169_ _081_ vss _385_/a_36_68# _385_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ vdd _299_/VPW net34 vdd vss _109_ mask\[7\] _105_ _299_/a_36_472# _299_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ vdd _437_/VPW _026_ mask\[8\] net54 vss net71 vdd _437_/a_2665_112# _437_/a_448_472#
+ _437_/a_796_472# _437_/a_36_151# _437_/a_1204_472# _437_/a_3041_156# _437_/a_1000_472#
+ _437_/a_1308_423# _437_/a_1456_156# _437_/a_1288_156# _437_/a_2248_156# _437_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_78 vdd FILLER_0_3_78/VPW vdd vss FILLER_0_3_78/a_36_472# FILLER_0_3_78/a_572_375#
+ FILLER_0_3_78/a_124_375# FILLER_0_3_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_368_ vdd _368_/VPW vdd vss trim_mask\[4\] _158_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_222_ vdd _222_/VPW vdd vss net38 net43 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ vdd _205_/VPW net22 vss vdd _048_ _205_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd FILLER_0_19_142/VPW vdd vss FILLER_0_19_142/a_36_472# FILLER_0_19_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ vdd _453_/VPW _042_ cal_count\[3\] net51 vss net68 vdd _453_/a_2665_112# _453_/a_448_472#
+ _453_/a_796_472# _453_/a_36_151# _453_/a_1204_472# _453_/a_3041_156# _453_/a_1000_472#
+ _453_/a_1308_423# _453_/a_1456_156# _453_/a_1288_156# _453_/a_2248_156# _453_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd _384_/VPW vdd vss _036_ _160_ _168_ _384_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd FILLER_0_10_107/VPW vdd vss FILLER_0_10_107/a_36_472# FILLER_0_10_107/a_572_375#
+ FILLER_0_10_107/a_124_375# FILLER_0_10_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd _298_/VPW vdd vss _010_ _104_ _108_ _298_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ vdd _436_/VPW _025_ mask\[7\] net54 vss net71 vdd _436_/a_2665_112# _436_/a_448_472#
+ _436_/a_796_472# _436_/a_36_151# _436_/a_1204_472# _436_/a_3041_156# _436_/a_1000_472#
+ _436_/a_1308_423# _436_/a_1456_156# _436_/a_1288_156# _436_/a_2248_156# _436_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vdd ANTENNA__408__A1/VPW vss _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ vdd _367_/VPW _153_ _154_ _157_ vdd vss _030_ _156_ _367_/a_36_68# _367_/a_244_472#
+ _367_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd FILLER_0_13_80/VPW vdd vss FILLER_0_13_80/a_36_472# FILLER_0_13_80/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd FILLER_0_1_192/VPW vdd vss FILLER_0_1_192/a_36_472# FILLER_0_1_192/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd FILLER_0_9_270/VPW vdd vss FILLER_0_9_270/a_36_472# FILLER_0_9_270/a_572_375#
+ FILLER_0_9_270/a_124_375# FILLER_0_9_270/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vdd _221_/VPW vss net38 _054_ vdd _221_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ vdd _419_/VPW _008_ net31 net60 vss net77 vdd _419_/a_2665_112# _419_/a_448_472#
+ _419_/a_796_472# _419_/a_36_151# _419_/a_1204_472# _419_/a_3041_156# _419_/a_1000_472#
+ _419_/a_1308_423# _419_/a_1456_156# _419_/a_1288_156# _419_/a_2248_156# _419_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd _204_/VPW vdd vss _048_ mask\[5\] net32 _204_/a_255_603# _204_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd FILLER_0_20_15/VPW vdd vss FILLER_0_20_15/a_1380_472# FILLER_0_20_15/a_36_472#
+ FILLER_0_20_15/a_932_472# FILLER_0_20_15/a_572_375# FILLER_0_20_15/a_124_375# FILLER_0_20_15/a_1468_375#
+ FILLER_0_20_15/a_1020_375# FILLER_0_20_15/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd FILLER_0_19_187/VPW vdd vss FILLER_0_19_187/a_36_472# FILLER_0_19_187/a_572_375#
+ FILLER_0_19_187/a_124_375# FILLER_0_19_187/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd FILLER_0_3_221/VPW vdd vss FILLER_0_3_221/a_1380_472# FILLER_0_3_221/a_36_472#
+ FILLER_0_3_221/a_932_472# FILLER_0_3_221/a_572_375# FILLER_0_3_221/a_124_375# FILLER_0_3_221/a_1468_375#
+ FILLER_0_3_221/a_1020_375# FILLER_0_3_221/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd FILLER_0_15_59/VPW vdd vss FILLER_0_15_59/a_36_472# FILLER_0_15_59/a_572_375#
+ FILLER_0_15_59/a_124_375# FILLER_0_15_59/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vdd ANTENNA_fanout58_I/VPW vss net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd FILLER_0_6_79/VPW vdd vss FILLER_0_6_79/a_36_472# FILLER_0_6_79/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vdd _452_/VPW vss net72 vdd _041_ cal_count\[2\] net55 _452_/a_448_472# _452_/a_36_151#
+ _452_/a_1293_527# _452_/a_3081_151# _452_/a_1284_156# _452_/a_1040_527# _452_/a_1353_112#
+ _452_/a_836_156# _452_/a_1697_156# _452_/a_2449_156# _452_/a_3129_107# _452_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ vdd _383_/VPW trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ _383_/a_36_472#
+ _383_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_297_ vdd _297_/VPW net33 vdd vss _108_ mask\[6\] _105_ _297_/a_36_472# _297_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ vdd _435_/VPW _024_ mask\[6\] net63 vss net80 vdd _435_/a_2665_112# _435_/a_448_472#
+ _435_/a_796_472# _435_/a_36_151# _435_/a_1204_472# _435_/a_3041_156# _435_/a_1000_472#
+ _435_/a_1308_423# _435_/a_1456_156# _435_/a_1288_156# _435_/a_2248_156# _435_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A2 vdd ANTENNA__408__A2/VPW vss cal_count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ vdd _366_/VPW vdd vss trim_mask\[3\] _157_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_127 vdd FILLER_0_2_127/VPW vdd vss FILLER_0_2_127/a_36_472# FILLER_0_2_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd FILLER_0_18_37/VPW vdd vss FILLER_0_18_37/a_1380_472# FILLER_0_18_37/a_36_472#
+ FILLER_0_18_37/a_932_472# FILLER_0_18_37/a_572_375# FILLER_0_18_37/a_124_375# FILLER_0_18_37/a_1468_375#
+ FILLER_0_18_37/a_1020_375# FILLER_0_18_37/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd FILLER_0_9_282/VPW vdd vss FILLER_0_9_282/a_36_472# FILLER_0_9_282/a_572_375#
+ FILLER_0_9_282/a_124_375# FILLER_0_9_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd _220_/VPW vdd vss _054_ trim_val\[0\] _053_ _220_/a_255_603# _220_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_349_ vdd _349_/VPW vdd vss _146_ _023_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ vdd _418_/VPW _007_ net30 net60 vss net77 vdd _418_/a_2665_112# _418_/a_448_472#
+ _418_/a_796_472# _418_/a_36_151# _418_/a_1204_472# _418_/a_3041_156# _418_/a_1000_472#
+ _418_/a_1308_423# _418_/a_1456_156# _418_/a_1288_156# _418_/a_2248_156# _418_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output21_I vdd ANTENNA_output21_I/VPW vss net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd _203_/VPW vdd vss net21 net11 vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd FILLER_0_19_155/VPW vdd vss FILLER_0_19_155/a_36_472# FILLER_0_19_155/a_572_375#
+ FILLER_0_19_155/a_124_375# FILLER_0_19_155/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd FILLER_0_19_111/VPW vdd vss FILLER_0_19_111/a_36_472# FILLER_0_19_111/a_572_375#
+ FILLER_0_19_111/a_124_375# FILLER_0_19_111/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd FILLER_0_22_128/VPW vdd vss FILLER_0_22_128/a_1916_375# FILLER_0_22_128/a_1380_472#
+ FILLER_0_22_128/a_3260_375# FILLER_0_22_128/a_36_472# FILLER_0_22_128/a_932_472#
+ FILLER_0_22_128/a_2812_375# FILLER_0_22_128/a_2276_472# FILLER_0_22_128/a_1828_472#
+ FILLER_0_22_128/a_3172_472# FILLER_0_22_128/a_572_375# FILLER_0_22_128/a_2724_472#
+ FILLER_0_22_128/a_124_375# FILLER_0_22_128/a_1468_375# FILLER_0_22_128/a_1020_375#
+ FILLER_0_22_128/a_484_472# FILLER_0_22_128/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd FILLER_0_15_180/VPW vdd vss FILLER_0_15_180/a_36_472# FILLER_0_15_180/a_572_375#
+ FILLER_0_15_180/a_124_375# FILLER_0_15_180/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd FILLER_0_21_150/VPW vdd vss FILLER_0_21_150/a_36_472# FILLER_0_21_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd FILLER_0_6_47/VPW vdd vss FILLER_0_6_47/a_1916_375# FILLER_0_6_47/a_1380_472#
+ FILLER_0_6_47/a_3260_375# FILLER_0_6_47/a_36_472# FILLER_0_6_47/a_932_472# FILLER_0_6_47/a_2812_375#
+ FILLER_0_6_47/a_2276_472# FILLER_0_6_47/a_1828_472# FILLER_0_6_47/a_3172_472# FILLER_0_6_47/a_572_375#
+ FILLER_0_6_47/a_2724_472# FILLER_0_6_47/a_124_375# FILLER_0_6_47/a_1468_375# FILLER_0_6_47/a_1020_375#
+ FILLER_0_6_47/a_484_472# FILLER_0_6_47/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_451_ vdd _451_/VPW vss net70 vdd _040_ cal_count\[1\] net53 _451_/a_448_472# _451_/a_36_151#
+ _451_/a_1293_527# _451_/a_3081_151# _451_/a_1284_156# _451_/a_1040_527# _451_/a_1353_112#
+ _451_/a_836_156# _451_/a_1697_156# _451_/a_2449_156# _451_/a_3129_107# _451_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_28 vdd FILLER_0_12_28/VPW vdd vss FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd _382_/VPW vdd vss _035_ _160_ _167_ _382_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd FILLER_0_18_209/VPW vdd vss FILLER_0_18_209/a_36_472# FILLER_0_18_209/a_572_375#
+ FILLER_0_18_209/a_124_375# FILLER_0_18_209/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd FILLER_0_5_136/VPW vdd vss FILLER_0_5_136/a_36_472# FILLER_0_5_136/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd _296_/VPW vdd vss _009_ _104_ _107_ _296_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ vdd _434_/VPW _023_ mask\[5\] net63 vss net80 vdd _434_/a_2665_112# _434_/a_448_472#
+ _434_/a_796_472# _434_/a_36_151# _434_/a_1204_472# _434_/a_3041_156# _434_/a_1000_472#
+ _434_/a_1308_423# _434_/a_1456_156# _434_/a_1288_156# _434_/a_2248_156# _434_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ vdd _365_/VPW _153_ _154_ _156_ vdd vss _029_ _155_ _365_/a_36_68# _365_/a_244_472#
+ _365_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vdd ANTENNA__280__A1/VPW vss _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vdd ANTENNA__240__I/VPW vss net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ vdd _348_/VPW _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ _348_/a_49_472#
+ _348_/a_665_69# _348_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ vdd _417_/VPW _006_ net29 net62 vss net79 vdd _417_/a_2665_112# _417_/a_448_472#
+ _417_/a_796_472# _417_/a_36_151# _417_/a_1204_472# _417_/a_3041_156# _417_/a_1000_472#
+ _417_/a_1308_423# _417_/a_1456_156# _417_/a_1288_156# _417_/a_2248_156# _417_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_279_ vdd _279_/VPW vdd vss _096_ _090_ state\[1\] _279_/a_652_68# _279_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_231 vdd FILLER_0_6_231/VPW vdd vss FILLER_0_6_231/a_36_472# FILLER_0_6_231/a_572_375#
+ FILLER_0_6_231/a_124_375# FILLER_0_6_231/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ vdd _202_/VPW net21 vss vdd _047_ _202_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output14_I vdd ANTENNA_output14_I/VPW vss net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd FILLER_0_4_91/VPW vdd vss FILLER_0_4_91/a_36_472# FILLER_0_4_91/a_572_375#
+ FILLER_0_4_91/a_124_375# FILLER_0_4_91/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_94 vdd FILLER_0_10_94/VPW vdd vss FILLER_0_10_94/a_36_472# FILLER_0_10_94/a_572_375#
+ FILLER_0_10_94/a_124_375# FILLER_0_10_94/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd FILLER_0_3_212/VPW vdd vss FILLER_0_3_212/a_36_472# FILLER_0_3_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd FILLER_0_19_134/VPW vdd vss FILLER_0_19_134/a_36_472# FILLER_0_19_134/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd FILLER_0_16_115/VPW vdd vss FILLER_0_16_115/a_36_472# FILLER_0_16_115/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd FILLER_0_22_107/VPW vdd vss FILLER_0_22_107/a_36_472# FILLER_0_22_107/a_572_375#
+ FILLER_0_22_107/a_124_375# FILLER_0_22_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd FILLER_0_21_60/VPW vdd vss FILLER_0_21_60/a_36_472# FILLER_0_21_60/a_572_375#
+ FILLER_0_21_60/a_124_375# FILLER_0_21_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd FILLER_0_6_37/VPW vdd vss FILLER_0_6_37/a_36_472# FILLER_0_6_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd FILLER_0_8_156/VPW vdd vss FILLER_0_8_156/a_36_472# FILLER_0_8_156/a_572_375#
+ FILLER_0_8_156/a_124_375# FILLER_0_8_156/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I vdd ANTENNA_input5_I/VPW vss rstn vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__243__I vdd ANTENNA__243__I/VPW vss net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_450_ vdd _450_/VPW vss net67 vdd _039_ cal_count\[0\] net51 _450_/a_448_472# _450_/a_36_151#
+ _450_/a_1293_527# _450_/a_3081_151# _450_/a_1284_156# _450_/a_1040_527# _450_/a_1353_112#
+ _450_/a_836_156# _450_/a_1697_156# _450_/a_2449_156# _450_/a_3129_107# _450_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xoutput40 vdd output40/VPW trim[2] net40 vdd vss output40/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_381_ vdd _381_/VPW trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ _381_/a_36_472#
+ _381_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_148 vdd FILLER_0_5_148/VPW vdd vss FILLER_0_5_148/a_36_472# FILLER_0_5_148/a_572_375#
+ FILLER_0_5_148/a_124_375# FILLER_0_5_148/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ vdd _433_/VPW _022_ mask\[4\] net54 vss net71 vdd _433_/a_2665_112# _433_/a_448_472#
+ _433_/a_796_472# _433_/a_36_151# _433_/a_1204_472# _433_/a_3041_156# _433_/a_1000_472#
+ _433_/a_1308_423# _433_/a_1456_156# _433_/a_1288_156# _433_/a_2248_156# _433_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ vdd _295_/VPW net32 vdd vss _107_ mask\[5\] _105_ _295_/a_36_472# _295_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd _364_/VPW vdd vss trim_mask\[2\] _156_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd FILLER_0_14_235/VPW vdd vss FILLER_0_14_235/a_36_472# FILLER_0_14_235/a_572_375#
+ FILLER_0_14_235/a_124_375# FILLER_0_14_235/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd FILLER_0_13_72/VPW vdd vss FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_572_375#
+ FILLER_0_13_72/a_124_375# FILLER_0_13_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_347_ vdd _347_/VPW vdd vss _145_ _022_ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ vdd _278_/VPW _095_ vss vdd net3 _278_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_290 vdd FILLER_0_13_290/VPW vdd vss FILLER_0_13_290/a_36_472# FILLER_0_13_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ vdd _416_/VPW _005_ net28 net62 vss net79 vdd _416_/a_2665_112# _416_/a_448_472#
+ _416_/a_796_472# _416_/a_36_151# _416_/a_1204_472# _416_/a_3041_156# _416_/a_1000_472#
+ _416_/a_1308_423# _416_/a_1456_156# _416_/a_1288_156# _416_/a_2248_156# _416_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_201_ vdd _201_/VPW vdd vss _047_ mask\[4\] net31 _201_/a_255_603# _201_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vdd ANTENNA__448__RN/VPW vss net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 vdd output30/VPW result[3] net30 vdd vss output30/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_196 vdd FILLER_0_12_196/VPW vdd vss FILLER_0_12_196/a_36_472# FILLER_0_12_196/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 vdd output6/VPW clkc net6 vdd vss output6/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 vdd output41/VPW trim[3] net41 vdd vss output41/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd _380_/VPW vdd vss _034_ _160_ _166_ _380_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
C0 output42/a_224_472# net6 0.010571f
C1 net17 FILLER_0_20_15/a_1020_375# 0.039975f
C2 net73 FILLER_0_18_107/a_36_472# 0.002425f
C3 _370_/a_848_380# vss 0.051599f
C4 _163_ FILLER_0_5_148/a_572_375# 0.001706f
C5 _131_ _124_ 0.002448f
C6 mask\[7\] FILLER_0_22_128/a_1916_375# 0.007718f
C7 trim_val\[3\] net14 0.01035f
C8 FILLER_0_17_72/a_1020_375# _175_ 0.028592f
C9 cal_count\[2\] FILLER_0_15_10/a_124_375# 0.017594f
C10 FILLER_0_18_177/a_3260_375# _047_ 0.030543f
C11 _070_ _389_/a_36_148# 0.010534f
C12 _255_/a_224_552# vss 0.001019f
C13 output27/a_224_472# net65 0.019729f
C14 net38 FILLER_0_12_2/a_572_375# 0.00609f
C15 FILLER_0_14_50/a_36_472# cal_count\[3\] 0.005814f
C16 FILLER_0_21_28/a_3172_472# _424_/a_36_151# 0.001723f
C17 trim_val\[3\] _164_ 0.018411f
C18 net61 output18/a_224_472# 0.059062f
C19 cal_itt\[2\] FILLER_0_3_221/a_572_375# 0.060779f
C20 net52 _439_/a_36_151# 0.01388f
C21 _335_/a_49_472# mask\[1\] 0.032497f
C22 FILLER_0_5_109/a_36_472# _163_ 0.00319f
C23 _096_ _085_ 0.0099f
C24 FILLER_0_16_57/a_484_472# FILLER_0_15_59/a_124_375# 0.001543f
C25 cal_itt\[2\] _000_ 0.042235f
C26 FILLER_0_9_28/a_1828_472# _054_ 0.003145f
C27 _394_/a_728_93# _043_ 0.00355f
C28 FILLER_0_4_152/a_36_472# net23 0.047194f
C29 _136_ net21 0.022198f
C30 _024_ vss 0.132549f
C31 result[9] result[5] 0.064058f
C32 mask\[4\] _091_ 0.071954f
C33 ctln[7] FILLER_0_0_96/a_36_472# 0.01317f
C34 _128_ _090_ 0.018296f
C35 _136_ _333_/a_36_160# 0.00842f
C36 cal_count\[1\] vss 0.307993f
C37 _428_/a_796_472# _095_ 0.00117f
C38 _178_ cal_count\[1\] 0.470244f
C39 _443_/a_2248_156# _170_ 0.068179f
C40 net15 _440_/a_796_472# 0.005848f
C41 _061_ _060_ 0.066418f
C42 state\[2\] FILLER_0_13_142/a_36_472# 0.022678f
C43 net53 FILLER_0_13_142/a_932_472# 0.059367f
C44 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_484_472# 0.026657f
C45 net63 _434_/a_2560_156# 0.014333f
C46 _091_ FILLER_0_13_212/a_1020_375# 0.00799f
C47 _015_ FILLER_0_8_247/a_124_375# 0.00706f
C48 FILLER_0_3_78/a_124_375# vdd 0.002419f
C49 _430_/a_448_472# _019_ 0.019666f
C50 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_36_472# 0.001723f
C51 _367_/a_36_68# net14 0.055776f
C52 _448_/a_2665_112# _037_ 0.042225f
C53 _091_ FILLER_0_10_214/a_36_472# 0.001357f
C54 net44 net40 0.003336f
C55 _161_ _062_ 0.046903f
C56 vdd trim[2] 0.166648f
C57 _345_/a_36_160# FILLER_0_19_125/a_124_375# 0.005398f
C58 FILLER_0_22_128/a_2812_375# vss 0.004347f
C59 FILLER_0_22_128/a_3260_375# vdd 0.005207f
C60 _100_ _094_ 0.031066f
C61 net71 FILLER_0_22_107/a_484_472# 0.00689f
C62 FILLER_0_9_28/a_1828_472# vss 0.001663f
C63 net33 vdd 0.42212f
C64 output15/a_224_472# FILLER_0_0_96/a_124_375# 0.00515f
C65 FILLER_0_3_78/a_36_472# _168_ 0.063262f
C66 FILLER_0_20_15/a_1380_472# net40 0.014911f
C67 _028_ _439_/a_1000_472# 0.003267f
C68 FILLER_0_6_79/a_36_472# vss 0.008693f
C69 result[9] output20/a_224_472# 0.001884f
C70 _129_ _062_ 0.20212f
C71 net31 _277_/a_36_160# 0.053915f
C72 _079_ FILLER_0_3_172/a_1828_472# 0.001638f
C73 _065_ fanout50/a_36_160# 0.022932f
C74 _425_/a_36_151# net19 0.009499f
C75 _115_ _070_ 0.890903f
C76 net76 _078_ 0.029213f
C77 _406_/a_36_159# _402_/a_56_567# 0.001025f
C78 net82 FILLER_0_3_172/a_1468_375# 0.010439f
C79 _008_ _094_ 0.234346f
C80 FILLER_0_21_206/a_124_375# _048_ 0.018458f
C81 _105_ _104_ 0.931514f
C82 FILLER_0_13_228/a_124_375# _043_ 0.133079f
C83 _114_ FILLER_0_11_101/a_124_375# 0.013348f
C84 FILLER_0_15_282/a_484_472# vss 0.005507f
C85 trim_val\[0\] _164_ 0.133785f
C86 FILLER_0_17_38/a_484_472# vdd 0.009211f
C87 _114_ _076_ 0.088609f
C88 _072_ _060_ 0.080908f
C89 FILLER_0_3_172/a_572_375# net65 0.008318f
C90 FILLER_0_3_2/a_124_375# output41/a_224_472# 0.030009f
C91 _105_ vss 0.485198f
C92 net79 _418_/a_36_151# 0.059124f
C93 _142_ mask\[2\] 0.093231f
C94 _392_/a_36_68# vss 0.002019f
C95 vss FILLER_0_3_212/a_124_375# 0.009048f
C96 vdd FILLER_0_3_212/a_36_472# 0.110132f
C97 FILLER_0_6_177/a_572_375# _163_ 0.001839f
C98 _116_ _061_ 0.04837f
C99 FILLER_0_17_282/a_124_375# vdd 0.004586f
C100 _152_ _261_/a_36_160# 0.001102f
C101 _414_/a_36_151# FILLER_0_6_177/a_484_472# 0.006095f
C102 _316_/a_848_380# calibrate 0.012121f
C103 _316_/a_124_24# _122_ 0.040082f
C104 _116_ _311_/a_66_473# 0.001527f
C105 _431_/a_2560_156# vss 0.004767f
C106 _149_ _098_ 0.398643f
C107 _131_ _041_ 0.035642f
C108 _028_ _086_ 0.011526f
C109 _306_/a_36_68# vdd 0.044152f
C110 net62 FILLER_0_21_286/a_572_375# 0.003744f
C111 FILLER_0_21_125/a_36_472# _436_/a_36_151# 0.001695f
C112 output36/a_224_472# net19 0.106928f
C113 FILLER_0_5_109/a_484_472# net47 0.002299f
C114 net20 _282_/a_36_160# 0.016884f
C115 _449_/a_36_151# _394_/a_1336_472# 0.001582f
C116 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_484_472# 0.001963f
C117 _415_/a_1000_472# _004_ 0.005004f
C118 net31 FILLER_0_16_255/a_124_375# 0.029277f
C119 net52 FILLER_0_6_47/a_3260_375# 0.040612f
C120 FILLER_0_23_60/a_124_375# vdd 0.031398f
C121 mask\[9\] FILLER_0_20_98/a_124_375# 0.003444f
C122 net55 FILLER_0_19_28/a_572_375# 0.002115f
C123 trimb[1] FILLER_0_18_2/a_1916_375# 0.001855f
C124 net20 FILLER_0_6_231/a_484_472# 0.017025f
C125 net20 _421_/a_448_472# 0.015767f
C126 _440_/a_2665_112# FILLER_0_4_91/a_124_375# 0.006271f
C127 FILLER_0_12_2/a_36_472# clkc 0.004826f
C128 _411_/a_2248_156# net10 0.002419f
C129 _432_/a_796_472# _093_ 0.002586f
C130 FILLER_0_4_144/a_36_472# vss 0.008308f
C131 FILLER_0_4_144/a_484_472# vdd 0.004027f
C132 FILLER_0_18_100/a_124_375# vdd 0.044014f
C133 _066_ net37 0.006164f
C134 _379_/a_36_472# _166_ 0.038062f
C135 _061_ _118_ 0.268815f
C136 _443_/a_1204_472# net69 0.002642f
C137 _257_/a_36_472# _070_ 0.002295f
C138 net54 FILLER_0_22_107/a_36_472# 0.043792f
C139 _426_/a_2665_112# FILLER_0_8_239/a_124_375# 0.010736f
C140 net63 FILLER_0_20_193/a_36_472# 0.048818f
C141 _433_/a_1308_423# _145_ 0.026613f
C142 net72 _403_/a_224_472# 0.002276f
C143 net74 _372_/a_170_472# 0.079123f
C144 _176_ _076_ 0.046873f
C145 _118_ _311_/a_66_473# 0.008528f
C146 _431_/a_448_472# net70 0.002293f
C147 _104_ output19/a_224_472# 0.064818f
C148 _105_ _107_ 0.020727f
C149 _072_ _116_ 0.283323f
C150 ctlp[3] result[8] 0.278543f
C151 _236_/a_36_160# net39 0.052649f
C152 _132_ _126_ 0.247838f
C153 net35 net22 0.001381f
C154 net23 FILLER_0_19_155/a_124_375# 0.001347f
C155 FILLER_0_17_72/a_124_375# vss 0.048053f
C156 FILLER_0_17_72/a_572_375# vdd 0.002455f
C157 FILLER_0_1_98/a_36_472# FILLER_0_0_96/a_124_375# 0.001684f
C158 _008_ net78 0.032202f
C159 net80 _136_ 0.034194f
C160 FILLER_0_18_2/a_484_472# vss 0.001228f
C161 cal_count\[3\] _121_ 0.011368f
C162 output19/a_224_472# vss 0.048948f
C163 FILLER_0_17_161/a_124_375# _137_ 0.016092f
C164 net81 _426_/a_448_472# 0.003907f
C165 net7 output41/a_224_472# 0.019483f
C166 net23 net37 0.01763f
C167 net4 calibrate 0.04302f
C168 FILLER_0_16_89/a_484_472# _451_/a_448_472# 0.059367f
C169 FILLER_0_4_107/a_124_375# vss 0.00322f
C170 FILLER_0_4_107/a_572_375# vdd 0.034678f
C171 FILLER_0_7_195/a_36_472# _055_ 0.03271f
C172 _077_ FILLER_0_12_50/a_36_472# 0.177624f
C173 FILLER_0_9_270/a_124_375# vdd 0.013312f
C174 _445_/a_2560_156# net47 0.014069f
C175 FILLER_0_9_28/a_1380_472# _120_ 0.00154f
C176 net38 FILLER_0_20_2/a_572_375# 0.004413f
C177 _065_ net14 0.005438f
C178 _413_/a_36_151# FILLER_0_4_197/a_36_472# 0.001512f
C179 _091_ _429_/a_448_472# 0.034713f
C180 ctlp[2] _422_/a_36_151# 0.068086f
C181 _395_/a_36_488# vdd 0.066813f
C182 trimb[0] net17 0.006176f
C183 fanout63/a_36_160# net64 0.016132f
C184 FILLER_0_17_200/a_484_472# net21 0.017997f
C185 net54 FILLER_0_20_98/a_36_472# 0.059367f
C186 net63 FILLER_0_18_177/a_1916_375# 0.040551f
C187 net57 FILLER_0_16_154/a_932_472# 0.003453f
C188 cal_count\[2\] _180_ 0.153207f
C189 _120_ vss 0.42505f
C190 _072_ _118_ 0.120452f
C191 _038_ vss 0.373776f
C192 net60 _421_/a_1308_423# 0.020693f
C193 _136_ mask\[1\] 0.407932f
C194 net48 cal_itt\[0\] 0.006171f
C195 _449_/a_2248_156# net74 0.004565f
C196 en_co_clk _176_ 0.099475f
C197 _401_/a_36_68# cal_count\[1\] 0.006747f
C198 _065_ _164_ 0.006953f
C199 FILLER_0_16_89/a_1468_375# _131_ 0.016581f
C200 output8/a_224_472# net4 0.015359f
C201 FILLER_0_12_136/a_932_472# _069_ 0.002161f
C202 FILLER_0_12_136/a_36_472# _126_ 0.014981f
C203 _009_ net77 0.001183f
C204 FILLER_0_23_282/a_124_375# vss 0.005048f
C205 FILLER_0_23_282/a_572_375# vdd -0.013698f
C206 net62 mask\[1\] 0.227329f
C207 net76 _263_/a_224_472# 0.00132f
C208 FILLER_0_13_142/a_1468_375# vdd 0.028002f
C209 _438_/a_2248_156# vss 0.002607f
C210 _438_/a_2665_112# vdd 0.00587f
C211 FILLER_0_13_142/a_1020_375# vss 0.005307f
C212 _030_ _440_/a_36_151# 0.001187f
C213 FILLER_0_5_172/a_36_472# net37 0.013857f
C214 _098_ FILLER_0_18_209/a_572_375# 0.001352f
C215 net52 FILLER_0_5_72/a_484_472# 0.050714f
C216 net50 FILLER_0_5_72/a_1468_375# 0.001777f
C217 _131_ FILLER_0_17_64/a_124_375# 0.005913f
C218 _056_ _062_ 0.320621f
C219 output19/a_224_472# _107_ 0.005034f
C220 state\[0\] _055_ 0.042917f
C221 net75 net59 0.06935f
C222 _087_ FILLER_0_5_172/a_124_375# 0.003043f
C223 net15 FILLER_0_9_72/a_124_375# 0.006492f
C224 _390_/a_36_68# _067_ 0.029588f
C225 net19 FILLER_0_14_263/a_36_472# 0.135429f
C226 output29/a_224_472# net18 0.010345f
C227 cal FILLER_0_1_266/a_572_375# 0.001707f
C228 FILLER_0_4_152/a_36_472# net57 0.015332f
C229 net44 FILLER_0_15_2/a_484_472# 0.047161f
C230 net52 _160_ 0.133292f
C231 _152_ FILLER_0_5_136/a_124_375# 0.039558f
C232 _081_ FILLER_0_5_136/a_36_472# 0.0028f
C233 net17 _190_/a_36_160# 0.04702f
C234 net73 net74 0.016949f
C235 _164_ FILLER_0_6_47/a_484_472# 0.012286f
C236 net54 _433_/a_36_151# 0.00661f
C237 fanout66/a_36_113# net15 0.024302f
C238 _050_ _210_/a_67_603# 0.006444f
C239 net68 FILLER_0_5_54/a_932_472# 0.013043f
C240 fanout72/a_36_113# _174_ 0.026207f
C241 FILLER_0_20_107/a_124_375# _098_ 0.01186f
C242 net32 ctlp[1] 0.032275f
C243 FILLER_0_11_282/a_36_472# vdd 0.106843f
C244 FILLER_0_11_282/a_124_375# vss 0.005415f
C245 net15 _453_/a_1308_423# 0.00293f
C246 net49 _160_ 1.243817f
C247 FILLER_0_15_142/a_572_375# vss 0.095176f
C248 _447_/a_2560_156# net69 0.001774f
C249 FILLER_0_14_81/a_124_375# _394_/a_728_93# 0.004587f
C250 FILLER_0_4_197/a_572_375# net21 0.041173f
C251 _068_ _062_ 0.089152f
C252 _070_ _134_ 0.087767f
C253 net64 _005_ 0.006192f
C254 _057_ _043_ 0.02152f
C255 _415_/a_36_151# net75 0.024047f
C256 _144_ FILLER_0_19_155/a_572_375# 0.003611f
C257 net73 _144_ 0.003657f
C258 mask\[8\] vss 0.378558f
C259 net35 vdd 1.0365f
C260 mask\[6\] vss 0.348967f
C261 _417_/a_2665_112# _006_ 0.023025f
C262 FILLER_0_7_104/a_1380_472# _131_ 0.043557f
C263 FILLER_0_9_223/a_484_472# net4 0.047334f
C264 ctlp[5] net23 0.025206f
C265 _086_ FILLER_0_5_172/a_124_375# 0.007355f
C266 FILLER_0_7_72/a_1020_375# _053_ 0.014569f
C267 _320_/a_36_472# _113_ 0.030365f
C268 net56 FILLER_0_17_142/a_572_375# 0.014948f
C269 FILLER_0_5_109/a_484_472# _154_ 0.039428f
C270 net75 _122_ 0.052177f
C271 _014_ _123_ 0.050082f
C272 FILLER_0_10_78/a_484_472# _439_/a_36_151# 0.00271f
C273 _429_/a_2665_112# mask\[1\] 0.001022f
C274 _411_/a_2665_112# _073_ 0.009313f
C275 _367_/a_36_68# _153_ 0.019803f
C276 _119_ FILLER_0_8_156/a_124_375# 0.025304f
C277 FILLER_0_17_56/a_484_472# vss 0.006298f
C278 net63 net33 0.048496f
C279 _025_ _436_/a_36_151# 0.026707f
C280 _449_/a_36_151# net72 0.039436f
C281 fanout52/a_36_160# vss 0.010082f
C282 FILLER_0_5_117/a_124_375# _163_ 0.003096f
C283 net75 FILLER_0_10_256/a_36_472# 0.010024f
C284 net80 FILLER_0_19_171/a_124_375# 0.024758f
C285 net79 _416_/a_2665_112# 0.035115f
C286 _093_ _094_ 0.003586f
C287 _093_ FILLER_0_17_218/a_572_375# 0.0029f
C288 net55 FILLER_0_18_76/a_36_472# 0.003695f
C289 net75 net64 0.037337f
C290 net62 _416_/a_2560_156# 0.010748f
C291 _132_ _436_/a_36_151# 0.00162f
C292 _424_/a_448_472# FILLER_0_18_37/a_1020_375# 0.001674f
C293 _430_/a_36_151# _019_ 0.019296f
C294 vss FILLER_0_13_290/a_36_472# 0.009561f
C295 output14/a_224_472# vdd 0.054725f
C296 cal_count\[3\] _408_/a_728_93# 0.040643f
C297 _432_/a_2665_112# _093_ 0.02266f
C298 _128_ _117_ 0.045015f
C299 FILLER_0_2_111/a_124_375# trim_mask\[3\] 0.004993f
C300 output44/a_224_472# vdd 0.043902f
C301 output31/a_224_472# _418_/a_2248_156# 0.023576f
C302 FILLER_0_8_127/a_124_375# net74 0.026604f
C303 state\[2\] vss 0.185787f
C304 _453_/a_796_472# _042_ 0.005463f
C305 _453_/a_1308_423# net51 0.001804f
C306 _136_ _171_ 0.008792f
C307 _095_ cal_count\[1\] 0.853949f
C308 output25/a_224_472# ctlp[7] 0.002088f
C309 net41 _233_/a_36_160# 0.053625f
C310 _058_ FILLER_0_10_94/a_36_472# 0.009346f
C311 _086_ net74 0.058077f
C312 _440_/a_448_472# _164_ 0.0036f
C313 FILLER_0_20_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001543f
C314 output44/a_224_472# FILLER_0_20_15/a_484_472# 0.0323f
C315 _102_ net30 0.043037f
C316 _448_/a_36_151# net76 0.03831f
C317 _175_ vss 0.162988f
C318 _010_ _420_/a_448_472# 0.027802f
C319 vdd _167_ 0.012869f
C320 FILLER_0_19_171/a_1468_375# vdd 0.064097f
C321 FILLER_0_15_150/a_36_472# fanout53/a_36_160# 0.002059f
C322 FILLER_0_22_86/a_932_472# net71 0.005789f
C323 net15 FILLER_0_13_72/a_484_472# 0.002925f
C324 _414_/a_1000_472# _003_ 0.002053f
C325 _114_ _090_ 0.001909f
C326 _451_/a_836_156# net14 0.00174f
C327 FILLER_0_5_72/a_1380_472# _164_ 0.049427f
C328 _412_/a_36_151# output37/a_224_472# 0.006358f
C329 net61 net18 0.71051f
C330 _088_ FILLER_0_4_213/a_36_472# 0.01735f
C331 net55 FILLER_0_21_28/a_3260_375# 0.006399f
C332 net72 FILLER_0_21_28/a_932_472# 0.015756f
C333 _058_ calibrate 0.075294f
C334 mask\[0\] _136_ 0.025838f
C335 net21 _047_ 0.048701f
C336 _091_ FILLER_0_15_180/a_484_472# 0.001757f
C337 _235_/a_67_603# vdd 0.026582f
C338 _242_/a_36_160# FILLER_0_5_148/a_484_472# 0.003699f
C339 _136_ FILLER_0_13_100/a_36_472# 0.005029f
C340 result[6] net19 0.834308f
C341 FILLER_0_24_96/a_36_472# vss 0.003218f
C342 trim_mask\[4\] FILLER_0_2_111/a_1468_375# 0.001226f
C343 net62 mask\[0\] 0.552008f
C344 _359_/a_36_488# _131_ 0.006398f
C345 FILLER_0_10_37/a_124_375# _173_ 0.00262f
C346 _053_ _077_ 0.123663f
C347 net20 FILLER_0_13_228/a_36_472# 0.020589f
C348 _414_/a_2665_112# _074_ 0.004912f
C349 _352_/a_49_472# mask\[7\] 0.001066f
C350 _058_ net21 0.004383f
C351 FILLER_0_4_185/a_36_472# _087_ 0.008805f
C352 FILLER_0_18_100/a_36_472# FILLER_0_17_72/a_3172_472# 0.05841f
C353 _033_ net67 0.148585f
C354 net22 vdd 1.920713f
C355 _440_/a_796_472# net47 0.002508f
C356 FILLER_0_18_61/a_124_375# FILLER_0_18_53/a_572_375# 0.012001f
C357 FILLER_0_18_2/a_2812_375# vdd 0.021655f
C358 output22/a_224_472# _435_/a_448_472# 0.010723f
C359 FILLER_0_4_177/a_124_375# net37 0.00459f
C360 _341_/a_49_472# mask\[2\] 0.026222f
C361 FILLER_0_14_107/a_1468_375# vdd 0.007687f
C362 _119_ _153_ 0.001741f
C363 _152_ _062_ 0.097086f
C364 net57 net37 0.091923f
C365 FILLER_0_8_138/a_36_472# _120_ 0.006759f
C366 FILLER_0_9_72/a_932_472# vss 0.007033f
C367 FILLER_0_9_72/a_1380_472# vdd 0.007659f
C368 _448_/a_36_151# FILLER_0_2_177/a_124_375# 0.001597f
C369 _420_/a_36_151# FILLER_0_23_282/a_484_472# 0.001723f
C370 cal_itt\[2\] ctln[1] 0.053339f
C371 FILLER_0_8_107/a_36_472# vss 0.006371f
C372 _389_/a_36_148# FILLER_0_10_94/a_36_472# 0.001723f
C373 FILLER_0_22_177/a_124_375# net33 0.013581f
C374 _431_/a_1204_472# _137_ 0.005886f
C375 net41 net49 0.392356f
C376 cal_itt\[3\] _375_/a_1612_497# 0.003901f
C377 ctlp[3] _109_ 0.001371f
C378 net15 FILLER_0_9_60/a_572_375# 0.047331f
C379 net1 vss 0.161208f
C380 _085_ _113_ 0.084246f
C381 _091_ FILLER_0_20_169/a_124_375# 0.003958f
C382 _187_ _181_ 0.001158f
C383 output24/a_224_472# ctlp[7] 0.060657f
C384 _453_/a_2560_156# vss 0.00337f
C385 _432_/a_2665_112# _337_/a_49_472# 0.001051f
C386 _016_ _043_ 0.030341f
C387 _122_ _059_ 0.190023f
C388 _430_/a_1308_423# net22 0.035518f
C389 FILLER_0_9_28/a_1468_375# _444_/a_2248_156# 0.001074f
C390 _015_ _426_/a_2560_156# 0.024461f
C391 _086_ _154_ 0.102849f
C392 input5/a_36_113# net5 0.061819f
C393 net2 input4/a_36_68# 0.031809f
C394 FILLER_0_7_72/a_2276_472# vdd 0.004035f
C395 net33 _435_/a_2665_112# 0.005831f
C396 FILLER_0_16_107/a_36_472# _040_ 0.015026f
C397 _089_ _122_ 0.006163f
C398 net78 _109_ 0.001432f
C399 _402_/a_1296_93# cal_count\[1\] 0.004472f
C400 _221_/a_36_160# _054_ 0.02124f
C401 output21/a_224_472# _104_ 0.002459f
C402 _136_ FILLER_0_16_154/a_36_472# 0.00615f
C403 _059_ _227_/a_36_160# 0.099735f
C404 _428_/a_448_472# _131_ 0.041178f
C405 _443_/a_2665_112# net59 0.0434f
C406 net62 _099_ 0.062012f
C407 net20 _083_ 0.230786f
C408 trimb[1] FILLER_0_20_2/a_484_472# 0.003628f
C409 _091_ FILLER_0_18_177/a_932_472# 0.002113f
C410 output21/a_224_472# vss 0.082781f
C411 net32 _421_/a_2560_156# 0.049213f
C412 _072_ _228_/a_36_68# 0.005788f
C413 vss _433_/a_2248_156# 0.034403f
C414 vdd _433_/a_2665_112# 0.002569f
C415 mask\[0\] _429_/a_2665_112# 0.016053f
C416 _087_ _079_ 0.251042f
C417 net74 FILLER_0_2_111/a_1468_375# 0.003854f
C418 _111_ FILLER_0_18_76/a_36_472# 0.006706f
C419 FILLER_0_3_172/a_2812_375# net22 0.013048f
C420 FILLER_0_18_53/a_484_472# vss 0.003579f
C421 FILLER_0_9_28/a_2364_375# net68 0.019969f
C422 _094_ _418_/a_1204_472# 0.009231f
C423 _057_ _267_/a_1568_472# 0.002083f
C424 FILLER_0_17_133/a_36_472# vss 0.006791f
C425 net54 _050_ 0.040506f
C426 _422_/a_36_151# mask\[7\] 0.043316f
C427 FILLER_0_17_72/a_932_472# net71 0.001418f
C428 cal_itt\[2\] _074_ 0.082824f
C429 _285_/a_36_472# _045_ 0.00269f
C430 result[6] _420_/a_36_151# 0.011901f
C431 _052_ FILLER_0_21_60/a_124_375# 0.002308f
C432 FILLER_0_16_57/a_932_472# _131_ 0.007885f
C433 _221_/a_36_160# vss 0.037067f
C434 FILLER_0_9_60/a_572_375# net51 0.002279f
C435 net34 FILLER_0_22_177/a_484_472# 0.003953f
C436 _078_ FILLER_0_6_231/a_36_472# 0.013046f
C437 FILLER_0_12_124/a_36_472# _131_ 0.028609f
C438 result[7] _108_ 0.063624f
C439 trim[4] output6/a_224_472# 0.004337f
C440 _115_ FILLER_0_10_94/a_36_472# 0.014605f
C441 net36 FILLER_0_16_115/a_36_472# 0.003805f
C442 _379_/a_36_472# trim_val\[1\] 0.00909f
C443 _321_/a_2034_472# _176_ 0.002722f
C444 _069_ _395_/a_36_488# 0.042974f
C445 result[7] net19 0.087363f
C446 _445_/a_1000_472# net40 0.015508f
C447 FILLER_0_21_142/a_124_375# FILLER_0_22_128/a_1828_472# 0.001543f
C448 _053_ FILLER_0_6_47/a_1468_375# 0.008103f
C449 net2 _001_ 0.081616f
C450 _093_ FILLER_0_17_72/a_484_472# 0.008637f
C451 FILLER_0_7_72/a_2724_472# _077_ 0.004635f
C452 FILLER_0_10_28/a_36_472# vss 0.001102f
C453 _008_ _418_/a_2248_156# 0.047066f
C454 FILLER_0_15_235/a_124_375# vss 0.001993f
C455 FILLER_0_15_235/a_572_375# vdd -0.005887f
C456 result[0] vss 0.291352f
C457 fanout63/a_36_160# mask\[2\] 0.026642f
C458 FILLER_0_9_105/a_36_472# vdd 0.009746f
C459 FILLER_0_9_105/a_572_375# vss 0.020145f
C460 FILLER_0_13_142/a_36_472# _043_ 0.011974f
C461 FILLER_0_20_177/a_36_472# vss 0.003944f
C462 FILLER_0_20_177/a_484_472# vdd 0.010805f
C463 _126_ net79 0.085443f
C464 FILLER_0_21_125/a_484_472# _098_ 0.002964f
C465 FILLER_0_5_54/a_124_375# FILLER_0_6_47/a_932_472# 0.001597f
C466 result[9] _418_/a_2665_112# 0.053489f
C467 _432_/a_1308_423# FILLER_0_18_177/a_36_472# 0.009119f
C468 _411_/a_36_151# vss 0.035447f
C469 FILLER_0_16_57/a_124_375# FILLER_0_17_56/a_124_375# 0.026339f
C470 output9/a_224_472# net18 0.114757f
C471 _192_/a_67_603# vdd 0.027014f
C472 output16/a_224_472# _447_/a_2248_156# 0.001937f
C473 net16 _447_/a_1000_472# 0.003207f
C474 output21/a_224_472# _107_ 0.086601f
C475 _013_ FILLER_0_21_28/a_1916_375# 0.006025f
C476 net36 FILLER_0_15_212/a_1020_375# 0.004863f
C477 FILLER_0_21_142/a_484_472# net23 0.005353f
C478 _414_/a_2665_112# _081_ 0.00247f
C479 _414_/a_2248_156# vss 0.00384f
C480 _176_ _318_/a_224_472# 0.003019f
C481 state\[0\] _426_/a_2665_112# 0.017088f
C482 net63 net35 0.126544f
C483 FILLER_0_2_165/a_124_375# net22 0.206491f
C484 ctln[3] net19 0.003077f
C485 FILLER_0_10_78/a_572_375# _120_ 0.006134f
C486 FILLER_0_18_107/a_572_375# vdd 0.00419f
C487 FILLER_0_18_107/a_124_375# vss 0.003425f
C488 _053_ net50 0.711279f
C489 FILLER_0_9_28/a_1468_375# net51 0.00111f
C490 _434_/a_36_151# _348_/a_49_472# 0.017459f
C491 _267_/a_224_472# _121_ 0.0029f
C492 _422_/a_796_472# vdd 0.003546f
C493 _021_ net80 0.254353f
C494 cal_count\[2\] _452_/a_3129_107# 0.008853f
C495 _062_ _113_ 0.020368f
C496 state\[2\] _071_ 0.04575f
C497 net79 FILLER_0_12_220/a_572_375# 0.010889f
C498 fanout80/a_36_113# net36 0.007625f
C499 _441_/a_1000_472# vss 0.01858f
C500 _242_/a_36_160# _386_/a_124_24# 0.031797f
C501 _232_/a_67_603# _164_ 0.076123f
C502 FILLER_0_7_162/a_124_375# _169_ 0.00336f
C503 _430_/a_1308_423# vdd 0.00218f
C504 output23/a_224_472# FILLER_0_22_128/a_2364_375# 0.002439f
C505 net55 _424_/a_1000_472# 0.001357f
C506 mask\[4\] FILLER_0_18_177/a_124_375# 0.016093f
C507 _064_ _446_/a_2560_156# 0.029586f
C508 _414_/a_2248_156# _075_ 0.044302f
C509 _415_/a_2248_156# net64 0.051575f
C510 net76 _080_ 0.03728f
C511 _447_/a_36_151# net68 0.040925f
C512 _372_/a_358_69# _160_ 0.001562f
C513 _412_/a_2665_112# fanout58/a_36_160# 0.001221f
C514 net53 FILLER_0_16_154/a_36_472# 0.006261f
C515 _125_ vss 0.149512f
C516 _024_ _147_ 0.006801f
C517 _093_ mask\[9\] 0.460108f
C518 FILLER_0_15_142/a_572_375# _095_ 0.003935f
C519 _318_/a_224_472# _124_ 0.001288f
C520 _430_/a_1000_472# mask\[2\] 0.00785f
C521 _131_ FILLER_0_17_104/a_1020_375# 0.006574f
C522 FILLER_0_6_239/a_36_472# vss 0.003177f
C523 ctlp[1] _421_/a_2665_112# 0.008695f
C524 _411_/a_2248_156# net8 0.06032f
C525 net15 _423_/a_448_472# 0.004833f
C526 FILLER_0_21_28/a_1468_375# _423_/a_36_151# 0.001543f
C527 _226_/a_860_68# net21 0.00107f
C528 _101_ _045_ 0.001111f
C529 _449_/a_448_472# _038_ 0.064169f
C530 FILLER_0_3_172/a_2812_375# vdd -0.012025f
C531 FILLER_0_5_54/a_1020_375# _440_/a_36_151# 0.059049f
C532 _359_/a_1044_488# _133_ 0.001894f
C533 _359_/a_1492_488# _070_ 0.0043f
C534 _359_/a_36_488# _076_ 0.005184f
C535 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_124_375# 0.012001f
C536 result[7] _420_/a_36_151# 0.006868f
C537 net63 FILLER_0_19_171/a_1468_375# 0.006671f
C538 FILLER_0_7_104/a_124_375# _058_ 0.006125f
C539 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1380_472# 0.013276f
C540 FILLER_0_9_28/a_2724_472# _453_/a_448_472# 0.008036f
C541 _052_ FILLER_0_18_37/a_124_375# 0.03242f
C542 _251_/a_906_472# vss 0.0016f
C543 _105_ _106_ 0.038327f
C544 _163_ FILLER_0_5_136/a_36_472# 0.007779f
C545 _267_/a_36_472# _090_ 0.001109f
C546 FILLER_0_21_286/a_124_375# _420_/a_36_151# 0.001597f
C547 output33/a_224_472# ctlp[1] 0.018552f
C548 net9 vdd 0.190349f
C549 result[1] net79 0.25261f
C550 net36 FILLER_0_15_205/a_36_472# 0.005101f
C551 _127_ net23 0.069001f
C552 net15 FILLER_0_17_72/a_484_472# 0.002925f
C553 output17/a_224_472# vdd 0.026649f
C554 cal_itt\[2\] _081_ 0.003204f
C555 vss _416_/a_1000_472# 0.001784f
C556 _422_/a_1204_472# _108_ 0.015401f
C557 _135_ vdd 0.018662f
C558 net57 _390_/a_36_68# 0.001112f
C559 _091_ _113_ 0.006236f
C560 net13 _170_ 0.001668f
C561 state\[2\] _095_ 0.001426f
C562 FILLER_0_11_142/a_572_375# cal_count\[3\] 0.014082f
C563 FILLER_0_22_177/a_572_375# mask\[6\] 0.002657f
C564 net35 FILLER_0_22_177/a_124_375# 0.0073f
C565 _098_ _434_/a_2665_112# 0.013854f
C566 net15 trim_mask\[1\] 0.042093f
C567 net63 net22 0.223664f
C568 net15 output16/a_224_472# 0.013768f
C569 net20 FILLER_0_17_226/a_124_375# 0.001895f
C570 _430_/a_2665_112# vdd 0.021353f
C571 FILLER_0_6_79/a_124_375# FILLER_0_6_47/a_3260_375# 0.012001f
C572 _176_ FILLER_0_11_78/a_124_375# 0.004803f
C573 net79 FILLER_0_12_236/a_484_472# 0.009305f
C574 net54 mask\[9\] 0.094381f
C575 _175_ _095_ 0.041931f
C576 _434_/a_796_472# _023_ 0.002118f
C577 _292_/a_36_160# _201_/a_67_603# 0.003917f
C578 FILLER_0_2_165/a_124_375# vdd 0.020315f
C579 cal_itt\[2\] net65 0.514538f
C580 FILLER_0_7_72/a_2724_472# net50 0.007192f
C581 FILLER_0_4_49/a_124_375# net49 0.005427f
C582 FILLER_0_4_49/a_484_472# net66 0.015555f
C583 _114_ _117_ 0.008886f
C584 net75 FILLER_0_8_247/a_572_375# 0.003962f
C585 FILLER_0_5_198/a_572_375# net22 0.029657f
C586 _140_ FILLER_0_22_128/a_3260_375# 0.003524f
C587 mask\[3\] _019_ 0.001403f
C588 _140_ net33 0.026401f
C589 fanout67/a_36_160# vdd 0.018829f
C590 result[7] _419_/a_448_472# 0.021809f
C591 _174_ cal_count\[3\] 0.053844f
C592 net35 _435_/a_2665_112# 0.007912f
C593 _412_/a_1456_156# net58 0.001045f
C594 trim_mask\[1\] FILLER_0_6_90/a_572_375# 0.001263f
C595 ctln[7] FILLER_0_0_130/a_124_375# 0.002726f
C596 FILLER_0_17_161/a_36_472# vss 0.003343f
C597 net69 net14 0.056927f
C598 cal_count\[2\] _278_/a_36_160# 0.023061f
C599 _018_ _043_ 0.0022f
C600 FILLER_0_15_290/a_36_472# _417_/a_36_151# 0.027236f
C601 net15 _447_/a_2665_112# 0.063341f
C602 _323_/a_36_113# FILLER_0_10_247/a_124_375# 0.001846f
C603 FILLER_0_14_107/a_36_472# _043_ 0.001661f
C604 net79 state\[1\] 0.005861f
C605 net41 _052_ 0.001927f
C606 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_36_472# 0.086635f
C607 _370_/a_124_24# _160_ 0.001126f
C608 _165_ _160_ 0.008705f
C609 net15 mask\[9\] 0.128816f
C610 _069_ net22 0.327999f
C611 _053_ cal_itt\[3\] 0.471909f
C612 cal_count\[2\] vss 0.361185f
C613 FILLER_0_24_63/a_36_472# output25/a_224_472# 0.002338f
C614 _178_ cal_count\[2\] 0.119443f
C615 net69 _164_ 0.040362f
C616 FILLER_0_7_72/a_36_472# net50 0.011974f
C617 net79 _007_ 0.096772f
C618 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_36_472# 0.086635f
C619 FILLER_0_4_197/a_932_472# FILLER_0_3_204/a_36_472# 0.026657f
C620 _255_/a_224_552# _375_/a_36_68# 0.00229f
C621 _013_ _424_/a_448_472# 0.043803f
C622 net72 FILLER_0_12_50/a_36_472# 0.002007f
C623 _420_/a_1308_423# vdd 0.00284f
C624 _420_/a_448_472# vss 0.007371f
C625 _095_ FILLER_0_14_107/a_1020_375# 0.014156f
C626 _094_ _045_ 0.102437f
C627 net19 _416_/a_2665_112# 0.059453f
C628 mask\[5\] net32 0.304094f
C629 net4 FILLER_0_12_220/a_1020_375# 0.020782f
C630 _141_ FILLER_0_19_155/a_124_375# 0.029562f
C631 input3/a_36_113# vss 0.043862f
C632 FILLER_0_19_47/a_36_472# _052_ 0.015772f
C633 FILLER_0_9_28/a_1916_375# vdd 0.01295f
C634 state\[0\] _223_/a_36_160# 0.070065f
C635 _398_/a_36_113# net3 0.099638f
C636 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3172_472# 0.013276f
C637 _444_/a_36_151# net67 0.055072f
C638 _177_ _451_/a_3129_107# 0.043731f
C639 net72 _394_/a_56_524# 0.066156f
C640 mask\[4\] _143_ 0.352305f
C641 FILLER_0_19_28/a_484_472# vss 0.001207f
C642 net52 _443_/a_36_151# 0.020518f
C643 valid _425_/a_2248_156# 0.00154f
C644 net47 _365_/a_692_472# 0.002051f
C645 _446_/a_2248_156# net66 0.002766f
C646 net76 vss 0.436111f
C647 net44 _450_/a_36_151# 0.026203f
C648 FILLER_0_10_78/a_36_472# _115_ 0.002611f
C649 vss _450_/a_448_472# -0.001661f
C650 cal_count\[3\] _373_/a_1254_68# 0.001391f
C651 FILLER_0_16_241/a_124_375# net30 0.028559f
C652 FILLER_0_7_72/a_572_375# vss 0.006884f
C653 _087_ FILLER_0_6_177/a_124_375# 0.001151f
C654 _322_/a_124_24# _070_ 0.033355f
C655 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1380_472# 0.026657f
C656 _423_/a_2665_112# vss 0.016881f
C657 net63 FILLER_0_20_177/a_484_472# 0.002172f
C658 _283_/a_36_472# vdd 0.092097f
C659 net40 _160_ 0.152292f
C660 trim_mask\[4\] _031_ 0.001262f
C661 _074_ _265_/a_224_472# 0.001223f
C662 _076_ FILLER_0_8_156/a_572_375# 0.010751f
C663 FILLER_0_20_193/a_572_375# _098_ 0.078973f
C664 FILLER_0_20_177/a_124_375# _434_/a_36_151# 0.059049f
C665 _412_/a_2665_112# net18 0.001321f
C666 _185_ cal_count\[1\] 0.001949f
C667 FILLER_0_16_154/a_124_375# vss 0.004317f
C668 FILLER_0_16_154/a_572_375# vdd 0.004706f
C669 _448_/a_36_151# FILLER_0_1_192/a_36_472# 0.008172f
C670 net63 vdd 1.002883f
C671 _253_/a_1100_68# _074_ 0.001563f
C672 net73 net70 0.040702f
C673 _150_ vss 0.016993f
C674 _424_/a_36_151# _423_/a_36_151# 0.006746f
C675 FILLER_0_20_193/a_572_375# _205_/a_36_160# 0.002828f
C676 FILLER_0_4_49/a_36_472# _164_ 0.033727f
C677 _440_/a_36_151# FILLER_0_6_47/a_3172_472# 0.001653f
C678 FILLER_0_21_142/a_572_375# net54 0.043619f
C679 _083_ _265_/a_244_68# 0.004022f
C680 FILLER_0_17_72/a_3172_472# vss 0.001338f
C681 _421_/a_36_151# _010_ 0.015107f
C682 _389_/a_36_148# _171_ 0.023988f
C683 net22 _435_/a_2665_112# 0.004214f
C684 FILLER_0_5_198/a_572_375# vdd 0.005402f
C685 FILLER_0_22_86/a_1468_375# net14 0.024975f
C686 _144_ _433_/a_36_151# 0.086558f
C687 FILLER_0_16_89/a_932_472# _040_ 0.00702f
C688 _043_ _278_/a_36_160# 0.004357f
C689 output32/a_224_472# _010_ 0.001508f
C690 _086_ FILLER_0_6_177/a_124_375# 0.043788f
C691 FILLER_0_4_123/a_36_472# _153_ 0.001419f
C692 FILLER_0_18_2/a_3172_472# FILLER_0_19_28/a_124_375# 0.001684f
C693 _430_/a_1308_423# net63 0.01125f
C694 FILLER_0_2_177/a_124_375# vss 0.00252f
C695 FILLER_0_2_177/a_572_375# vdd 0.022268f
C696 net19 _420_/a_1000_472# 0.006558f
C697 FILLER_0_16_89/a_572_375# _093_ 0.002889f
C698 FILLER_0_12_136/a_572_375# _127_ 0.00116f
C699 FILLER_0_15_150/a_124_375# net56 0.011873f
C700 _372_/a_3126_472# _068_ 0.005304f
C701 net74 FILLER_0_13_72/a_484_472# 0.007142f
C702 _043_ vss 1.362912f
C703 _178_ _043_ 0.130207f
C704 _211_/a_36_160# net14 0.005761f
C705 _000_ _260_/a_36_68# 0.004354f
C706 net68 _054_ 0.08092f
C707 _449_/a_1308_423# _453_/a_2665_112# 0.001066f
C708 net7 net17 0.050676f
C709 _069_ vdd 0.985405f
C710 FILLER_0_8_138/a_124_375# _070_ 0.002997f
C711 _139_ net36 0.024268f
C712 sample en 0.001572f
C713 FILLER_0_13_212/a_124_375# net79 0.007396f
C714 ctln[4] net75 0.00718f
C715 net62 FILLER_0_13_212/a_572_375# 0.001597f
C716 _239_/a_36_160# net40 0.010925f
C717 net76 fanout76/a_36_160# 0.004503f
C718 _430_/a_36_151# FILLER_0_18_177/a_2276_472# 0.001793f
C719 FILLER_0_9_28/a_1380_472# net68 0.008573f
C720 net4 FILLER_0_3_221/a_572_375# 0.030599f
C721 net46 vss 0.110452f
C722 output9/a_224_472# net65 0.095296f
C723 mask\[7\] _435_/a_1000_472# 0.024725f
C724 _147_ mask\[6\] 0.103475f
C725 _000_ net4 0.036895f
C726 _131_ FILLER_0_14_123/a_36_472# 0.029747f
C727 mask\[5\] FILLER_0_19_155/a_572_375# 0.007026f
C728 net68 vss 0.635359f
C729 net25 FILLER_0_22_86/a_36_472# 0.001265f
C730 _430_/a_1308_423# _069_ 0.024499f
C731 cal_itt\[0\] net8 0.026229f
C732 output47/a_224_472# net40 0.002339f
C733 _110_ net71 0.004816f
C734 _273_/a_36_68# _091_ 0.00155f
C735 _026_ vss 0.005992f
C736 net23 FILLER_0_22_128/a_2724_472# 0.054521f
C737 net50 _447_/a_448_472# 0.001219f
C738 _115_ _171_ 0.033359f
C739 net80 _435_/a_1000_472# 0.001079f
C740 _426_/a_1308_423# calibrate 0.001708f
C741 FILLER_0_18_139/a_1468_375# vss 0.009191f
C742 FILLER_0_18_139/a_36_472# vdd 0.089771f
C743 FILLER_0_16_107/a_484_472# net14 0.001528f
C744 _408_/a_718_524# _067_ 0.006516f
C745 _028_ trim_mask\[1\] 0.148182f
C746 _377_/a_36_472# _164_ 0.03259f
C747 FILLER_0_9_72/a_484_472# _439_/a_36_151# 0.001723f
C748 net54 _022_ 0.004106f
C749 _093_ FILLER_0_18_107/a_484_472# 0.008683f
C750 FILLER_0_15_282/a_572_375# net18 0.00298f
C751 FILLER_0_22_177/a_124_375# vdd 0.001293f
C752 FILLER_0_18_107/a_36_472# mask\[9\] 0.005458f
C753 FILLER_0_15_282/a_36_472# net30 0.001692f
C754 FILLER_0_15_282/a_124_375# result[3] 0.004601f
C755 output11/a_224_472# ctln[3] 0.068614f
C756 cal_count\[2\] _184_ 0.033241f
C757 _390_/a_244_472# _136_ 0.001777f
C758 _114_ _172_ 0.045798f
C759 net20 result[6] 0.026511f
C760 trim_val\[3\] _441_/a_448_472# 0.00469f
C761 FILLER_0_4_177/a_36_472# _074_ 0.002603f
C762 cal_count\[2\] _401_/a_36_68# 0.008136f
C763 vss _156_ 0.089339f
C764 _426_/a_448_472# net64 0.054931f
C765 _198_/a_67_603# net30 0.017304f
C766 _064_ trim[1] 0.166575f
C767 net67 _054_ 0.391592f
C768 _439_/a_36_151# _453_/a_2665_112# 0.001738f
C769 _430_/a_2665_112# net63 0.075661f
C770 _095_ _280_/a_224_472# 0.001416f
C771 net35 _140_ 0.12583f
C772 net71 _437_/a_2665_112# 0.039687f
C773 _081_ _265_/a_224_472# 0.008598f
C774 net41 net40 2.687418f
C775 _435_/a_2665_112# vdd 0.01769f
C776 FILLER_0_21_142/a_36_472# FILLER_0_22_128/a_1468_375# 0.001543f
C777 FILLER_0_17_72/a_3260_375# net14 0.040606f
C778 _136_ _451_/a_1040_527# 0.00497f
C779 net27 _323_/a_36_113# 0.010949f
C780 _449_/a_36_151# vdd 0.09324f
C781 _210_/a_67_603# net23 0.005398f
C782 _303_/a_36_472# FILLER_0_20_87/a_36_472# 0.005725f
C783 _079_ _001_ 0.082209f
C784 net81 net79 0.178225f
C785 fanout65/a_36_113# vss 0.053899f
C786 _443_/a_796_472# net23 0.002306f
C787 _443_/a_448_472# net13 0.002263f
C788 net28 vdd 0.489756f
C789 net28 _192_/a_67_603# 0.119061f
C790 FILLER_0_9_223/a_572_375# vdd 0.007158f
C791 _431_/a_448_472# FILLER_0_17_142/a_124_375# 0.006782f
C792 _149_ _437_/a_448_472# 0.009274f
C793 _392_/a_36_68# cal_count\[0\] 0.038691f
C794 _053_ FILLER_0_5_54/a_484_472# 0.001135f
C795 net67 vss 0.435869f
C796 FILLER_0_11_124/a_36_472# _120_ 0.014712f
C797 _131_ _136_ 1.42765f
C798 trim_val\[4\] _443_/a_2665_112# 0.018733f
C799 net21 FILLER_0_12_196/a_124_375# 0.005374f
C800 _412_/a_2248_156# fanout58/a_36_160# 0.005856f
C801 _176_ _172_ 0.043154f
C802 _031_ _154_ 0.037238f
C803 net69 _153_ 0.003678f
C804 _255_/a_224_552# _070_ 0.001333f
C805 FILLER_0_20_193/a_484_472# FILLER_0_18_177/a_2364_375# 0.0027f
C806 sample output27/a_224_472# 0.006116f
C807 ctln[7] net52 0.06558f
C808 _415_/a_448_472# net18 0.057688f
C809 _105_ _098_ 0.055065f
C810 FILLER_0_21_133/a_36_472# vdd 0.092168f
C811 net72 _182_ 0.044895f
C812 net50 FILLER_0_8_24/a_124_375# 0.001597f
C813 FILLER_0_11_64/a_36_472# vss 0.006069f
C814 FILLER_0_24_290/a_36_472# FILLER_0_23_290/a_36_472# 0.05841f
C815 FILLER_0_12_236/a_572_375# vdd 0.024713f
C816 FILLER_0_12_236/a_124_375# vss 0.001024f
C817 _412_/a_36_151# net58 0.010226f
C818 _415_/a_2665_112# net64 0.074373f
C819 net71 net14 0.147175f
C820 _376_/a_36_160# FILLER_0_5_72/a_1380_472# 0.035111f
C821 FILLER_0_14_91/a_572_375# vdd -0.011429f
C822 _105_ _205_/a_36_160# 0.001167f
C823 _442_/a_448_472# _031_ 0.019293f
C824 _445_/a_1308_423# vdd 0.001478f
C825 FILLER_0_21_28/a_932_472# vdd 0.04815f
C826 FILLER_0_18_209/a_484_472# vss 0.005794f
C827 net52 FILLER_0_2_93/a_484_472# 0.009006f
C828 net50 FILLER_0_2_93/a_572_375# 0.00275f
C829 _246_/a_36_68# _090_ 0.001712f
C830 _423_/a_448_472# _012_ 0.038928f
C831 _429_/a_36_151# _136_ 0.001188f
C832 _144_ FILLER_0_19_125/a_124_375# 0.012834f
C833 _144_ FILLER_0_22_128/a_3172_472# 0.001287f
C834 _001_ cal_itt\[1\] 0.057933f
C835 ctlp[7] _211_/a_36_160# 0.003488f
C836 _152_ _153_ 0.002954f
C837 _074_ _084_ 0.110937f
C838 FILLER_0_8_239/a_36_472# calibrate 0.008683f
C839 net54 _437_/a_2248_156# 0.046559f
C840 _013_ _217_/a_36_160# 0.001614f
C841 net20 result[7] 0.134149f
C842 FILLER_0_21_28/a_1020_375# _424_/a_36_151# 0.001252f
C843 fanout70/a_36_113# _131_ 0.003364f
C844 net34 _023_ 0.00872f
C845 net76 FILLER_0_5_198/a_36_472# 0.003987f
C846 comp vss 0.148428f
C847 net62 net18 0.089041f
C848 net31 _104_ 0.102776f
C849 mask\[4\] _291_/a_36_160# 0.00591f
C850 net81 _429_/a_2560_156# 0.003888f
C851 net15 net66 0.006618f
C852 _430_/a_448_472# _091_ 0.065306f
C853 FILLER_0_14_50/a_124_375# cal_count\[1\] 0.023752f
C854 net56 _136_ 0.462275f
C855 _068_ _315_/a_716_497# 0.00217f
C856 _076_ _315_/a_36_68# 0.001568f
C857 _070_ _315_/a_1657_68# 0.001601f
C858 net3 _190_/a_36_160# 0.013324f
C859 _095_ cal_count\[2\] 0.270066f
C860 _412_/a_36_151# _082_ 0.016538f
C861 output38/a_224_472# trim[1] 0.003114f
C862 net38 net39 0.066083f
C863 output42/a_224_472# FILLER_0_9_28/a_36_472# 0.010684f
C864 result[1] net19 0.084617f
C865 net15 _067_ 0.042278f
C866 trim_mask\[1\] net47 0.306848f
C867 _412_/a_36_151# net82 0.064296f
C868 FILLER_0_12_20/a_484_472# net17 0.05005f
C869 net77 vdd 0.526632f
C870 net31 vss 0.562041f
C871 net62 _196_/a_36_160# 0.029171f
C872 trim_val\[2\] net49 0.00301f
C873 net76 FILLER_0_2_177/a_36_472# 0.003526f
C874 _009_ FILLER_0_23_282/a_484_472# 0.009744f
C875 ctln[0] net40 0.001334f
C876 output28/a_224_472# _416_/a_2665_112# 0.008243f
C877 _150_ _027_ 0.006689f
C878 net16 _450_/a_2225_156# 0.001015f
C879 _112_ _425_/a_448_472# 0.002335f
C880 result[9] FILLER_0_23_274/a_124_375# 0.003102f
C881 net55 cal_count\[1\] 0.204733f
C882 FILLER_0_16_57/a_572_375# _176_ 0.006422f
C883 net53 _451_/a_1040_527# 0.023651f
C884 _120_ cal_count\[0\] 0.014209f
C885 _131_ FILLER_0_17_56/a_572_375# 0.006224f
C886 net16 _183_ 0.001103f
C887 FILLER_0_15_116/a_36_472# FILLER_0_17_104/a_1468_375# 0.001512f
C888 _425_/a_2560_156# net37 0.002508f
C889 _102_ _006_ 0.006115f
C890 _176_ _183_ 0.024038f
C891 _412_/a_1000_472# cal_itt\[1\] 0.012926f
C892 ctlp[6] vss 0.115894f
C893 _095_ _450_/a_448_472# 0.001393f
C894 mask\[5\] FILLER_0_19_187/a_36_472# 0.007596f
C895 _093_ net23 0.042838f
C896 _256_/a_36_68# net4 0.017783f
C897 _118_ net23 0.108864f
C898 net35 FILLER_0_21_150/a_36_472# 0.004456f
C899 _103_ _102_ 0.392644f
C900 output47/a_224_472# FILLER_0_15_2/a_484_472# 0.038484f
C901 _413_/a_2248_156# net82 0.009308f
C902 FILLER_0_10_78/a_932_472# vdd 0.005517f
C903 _132_ FILLER_0_15_116/a_36_472# 0.020589f
C904 FILLER_0_9_142/a_124_375# _313_/a_67_603# 0.029786f
C905 mask\[5\] output33/a_224_472# 0.0238f
C906 net53 _131_ 0.059223f
C907 FILLER_0_14_81/a_124_375# vss 0.03341f
C908 FILLER_0_14_81/a_36_472# vdd 0.00958f
C909 net60 _418_/a_448_472# 0.055895f
C910 net63 _069_ 0.04528f
C911 result[2] vss 0.327009f
C912 net29 mask\[1\] 0.023266f
C913 output44/a_224_472# net43 0.001041f
C914 FILLER_0_7_162/a_36_472# _119_ 0.005739f
C915 _426_/a_1204_472# vdd 0.003412f
C916 _028_ FILLER_0_6_90/a_36_472# 0.013106f
C917 net82 _370_/a_848_380# 0.014538f
C918 _439_/a_2248_156# trim_mask\[0\] 0.005416f
C919 _140_ _433_/a_2665_112# 0.001108f
C920 _098_ _438_/a_2248_156# 0.002798f
C921 FILLER_0_9_290/a_124_375# vss 0.033914f
C922 FILLER_0_9_290/a_36_472# vdd 0.094552f
C923 FILLER_0_12_220/a_1380_472# _060_ 0.01563f
C924 net61 FILLER_0_21_286/a_484_472# 0.001829f
C925 _176_ FILLER_0_15_59/a_572_375# 0.007169f
C926 FILLER_0_16_89/a_1380_472# vss 0.005351f
C927 _065_ _441_/a_448_472# 0.001973f
C928 mask\[9\] _012_ 0.008145f
C929 net79 _417_/a_36_151# 0.082646f
C930 output27/a_224_472# FILLER_0_9_282/a_572_375# 0.029138f
C931 _427_/a_1000_472# net74 0.009646f
C932 net55 FILLER_0_17_38/a_36_472# 0.010728f
C933 net62 _417_/a_448_472# 0.011318f
C934 result[6] _009_ 0.095754f
C935 _057_ _250_/a_36_68# 0.014333f
C936 FILLER_0_6_47/a_2364_375# vdd 0.015888f
C937 FILLER_0_6_47/a_1916_375# vss 0.005279f
C938 _187_ net51 0.04894f
C939 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_36_472# 0.016748f
C940 FILLER_0_4_197/a_36_472# net22 0.003404f
C941 _321_/a_3662_472# net74 0.00253f
C942 ctlp[1] net78 0.025929f
C943 _431_/a_2665_112# FILLER_0_17_142/a_124_375# 0.004834f
C944 _068_ FILLER_0_5_148/a_36_472# 0.003015f
C945 _095_ _043_ 2.807456f
C946 net60 mask\[7\] 0.001053f
C947 output15/a_224_472# trim_mask\[3\] 0.024718f
C948 cal_count\[2\] _402_/a_1296_93# 0.022009f
C949 FILLER_0_17_38/a_484_472# _182_ 0.00527f
C950 _431_/a_1000_472# net36 0.001771f
C951 _320_/a_36_472# FILLER_0_13_206/a_36_472# 0.038251f
C952 net54 net23 0.084191f
C953 cal net8 0.271166f
C954 FILLER_0_8_107/a_124_375# _219_/a_36_160# 0.002515f
C955 _119_ _059_ 0.039711f
C956 _432_/a_2665_112# _019_ 0.002852f
C957 _428_/a_2665_112# state\[2\] 0.001746f
C958 _140_ vdd 0.598538f
C959 _282_/a_36_160# vdd 0.010099f
C960 net56 net53 0.053535f
C961 _412_/a_2248_156# net18 0.05155f
C962 FILLER_0_6_90/a_124_375# net14 0.005361f
C963 _050_ _436_/a_1204_472# 0.006724f
C964 _081_ _084_ 0.016804f
C965 net27 FILLER_0_9_282/a_36_472# 0.002962f
C966 _161_ _311_/a_1212_473# 0.004138f
C967 _098_ mask\[6\] 0.297837f
C968 mask\[8\] _098_ 0.096999f
C969 vss FILLER_0_6_231/a_36_472# 0.0048f
C970 vdd FILLER_0_6_231/a_484_472# 0.004642f
C971 _086_ _331_/a_448_472# 0.004356f
C972 _421_/a_36_151# vss 0.021759f
C973 _421_/a_448_472# vdd 0.030898f
C974 _070_ _120_ 0.838223f
C975 net63 _435_/a_2665_112# 0.039512f
C976 result[9] FILLER_0_24_274/a_1020_375# 0.001657f
C977 net67 _450_/a_1040_527# 0.032098f
C978 _038_ _070_ 0.075667f
C979 FILLER_0_18_107/a_3172_472# vss 0.006614f
C980 ctln[2] net19 0.073057f
C981 _136_ FILLER_0_15_180/a_36_472# 0.006924f
C982 _435_/a_36_151# _434_/a_1308_423# 0.001518f
C983 result[8] FILLER_0_24_274/a_572_375# 0.00726f
C984 output32/a_224_472# vss -0.003023f
C985 _424_/a_2665_112# vdd 0.013636f
C986 _424_/a_2248_156# vss 0.004855f
C987 net26 FILLER_0_23_44/a_572_375# 0.003172f
C988 FILLER_0_1_192/a_36_472# vss 0.004422f
C989 _320_/a_1568_472# state\[1\] 0.001531f
C990 net4 net18 0.034592f
C991 result[2] _416_/a_2248_156# 0.001396f
C992 net55 FILLER_0_17_72/a_124_375# 0.019544f
C993 net15 net25 0.013745f
C994 net65 _084_ 0.031674f
C995 mask\[4\] FILLER_0_18_177/a_3172_472# 0.014657f
C996 _093_ FILLER_0_17_104/a_124_375# 0.01418f
C997 _105_ output35/a_224_472# 0.013092f
C998 _144_ mask\[9\] 0.001909f
C999 net50 _441_/a_2665_112# 0.056602f
C1000 output37/a_224_472# net76 0.004028f
C1001 mask\[3\] FILLER_0_18_177/a_2276_472# 0.01204f
C1002 net68 _036_ 0.168017f
C1003 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_484_472# 0.013276f
C1004 _277_/a_36_160# vss 0.030147f
C1005 net82 FILLER_0_3_212/a_124_375# 0.015932f
C1006 trim_mask\[1\] _154_ 0.004835f
C1007 FILLER_0_8_37/a_124_375# vdd 0.029725f
C1008 _049_ FILLER_0_22_128/a_3260_375# 0.16381f
C1009 net25 FILLER_0_23_44/a_1380_472# 0.0014f
C1010 result[9] FILLER_0_15_282/a_124_375# 0.001233f
C1011 _269_/a_36_472# net59 0.011985f
C1012 _340_/a_36_160# FILLER_0_20_169/a_36_472# 0.195478f
C1013 output25/a_224_472# _213_/a_67_603# 0.032497f
C1014 FILLER_0_21_125/a_484_472# mask\[7\] 0.003404f
C1015 FILLER_0_21_28/a_1468_375# _012_ 0.00351f
C1016 net34 _297_/a_36_472# 0.005603f
C1017 _074_ FILLER_0_6_177/a_484_472# 0.002068f
C1018 mask\[3\] FILLER_0_17_218/a_36_472# 0.015535f
C1019 _411_/a_2248_156# _073_ 0.003809f
C1020 FILLER_0_5_72/a_1020_375# vss 0.004157f
C1021 FILLER_0_5_72/a_1468_375# vdd 0.001826f
C1022 net21 _434_/a_2665_112# 0.004945f
C1023 _397_/a_36_472# net36 0.010045f
C1024 net69 FILLER_0_2_111/a_932_472# 0.011453f
C1025 net14 FILLER_0_4_91/a_484_472# 0.020589f
C1026 _031_ FILLER_0_2_111/a_36_472# 0.034656f
C1027 net55 _120_ 0.001054f
C1028 net55 _038_ 0.05656f
C1029 en_co_clk _136_ 0.034892f
C1030 _050_ FILLER_0_22_128/a_572_375# 0.002607f
C1031 net61 _422_/a_2560_156# 0.010748f
C1032 net20 _259_/a_455_68# 0.001427f
C1033 _289_/a_36_472# net30 0.009623f
C1034 FILLER_0_5_54/a_1020_375# _029_ 0.024737f
C1035 FILLER_0_4_144/a_124_375# _081_ 0.004558f
C1036 _122_ FILLER_0_8_156/a_36_472# 0.047846f
C1037 _057_ _310_/a_49_472# 0.015839f
C1038 result[7] _009_ 0.697145f
C1039 _315_/a_1229_68# _121_ 0.003401f
C1040 _183_ _041_ 0.001931f
C1041 _441_/a_36_151# _440_/a_1308_423# 0.001736f
C1042 net38 clkc 0.088241f
C1043 FILLER_0_7_72/a_1828_472# net52 0.00159f
C1044 _119_ FILLER_0_7_162/a_124_375# 0.059009f
C1045 _451_/a_36_151# vdd 0.088651f
C1046 _154_ _157_ 0.447829f
C1047 FILLER_0_21_286/a_124_375# _009_ 0.001024f
C1048 FILLER_0_9_223/a_124_375# _068_ 0.010485f
C1049 _446_/a_796_472# net40 0.001504f
C1050 _028_ FILLER_0_7_104/a_484_472# 0.00499f
C1051 FILLER_0_1_98/a_36_472# trim_mask\[3\] 0.106084f
C1052 _426_/a_36_151# FILLER_0_8_247/a_1020_375# 0.059049f
C1053 FILLER_0_4_197/a_36_472# vdd 0.042721f
C1054 _227_/a_36_160# FILLER_0_8_156/a_36_472# 0.006647f
C1055 FILLER_0_16_255/a_36_472# vdd 0.044615f
C1056 _081_ FILLER_0_5_148/a_484_472# 0.016132f
C1057 _274_/a_1164_497# net64 0.002049f
C1058 _421_/a_796_472# net19 0.009462f
C1059 _415_/a_2560_156# net27 0.008433f
C1060 ctln[1] net4 0.009703f
C1061 net57 _116_ 0.069858f
C1062 output12/a_224_472# net12 0.007193f
C1063 _093_ FILLER_0_19_134/a_124_375# 0.003473f
C1064 _363_/a_36_68# vdd 0.04306f
C1065 _077_ _055_ 0.083808f
C1066 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_36_472# 0.086635f
C1067 net27 fanout62/a_36_160# 0.005558f
C1068 net34 result[8] 0.076645f
C1069 _253_/a_244_68# _073_ 0.002878f
C1070 _256_/a_36_68# _058_ 0.001402f
C1071 output35/a_224_472# output19/a_224_472# 0.015892f
C1072 _186_ _402_/a_728_93# 0.002381f
C1073 FILLER_0_14_91/a_36_472# _043_ 0.001779f
C1074 FILLER_0_11_124/a_124_375# vdd 0.016626f
C1075 _168_ _160_ 0.03261f
C1076 _170_ _386_/a_124_24# 0.008511f
C1077 net16 _445_/a_2665_112# 0.061595f
C1078 net50 FILLER_0_5_88/a_36_472# 0.00867f
C1079 FILLER_0_22_177/a_1380_472# _435_/a_36_151# 0.001723f
C1080 _091_ FILLER_0_15_212/a_1468_375# 0.002531f
C1081 _002_ net59 0.016205f
C1082 _408_/a_56_524# FILLER_0_12_20/a_572_375# 0.009967f
C1083 _431_/a_36_151# net36 0.006618f
C1084 net43 vdd 0.210686f
C1085 net34 FILLER_0_22_128/a_2724_472# 0.004465f
C1086 net73 FILLER_0_15_142/a_36_472# 0.001893f
C1087 _091_ FILLER_0_16_154/a_1380_472# 0.00133f
C1088 _372_/a_170_472# _062_ 0.014919f
C1089 FILLER_0_8_138/a_124_375# calibrate 0.013177f
C1090 net70 FILLER_0_11_101/a_484_472# 0.001474f
C1091 FILLER_0_14_91/a_124_375# _095_ 0.01418f
C1092 FILLER_0_15_150/a_124_375# _427_/a_448_472# 0.008952f
C1093 _350_/a_49_472# net23 0.002397f
C1094 _127_ FILLER_0_9_142/a_36_472# 0.004721f
C1095 net43 FILLER_0_20_15/a_484_472# 0.001534f
C1096 FILLER_0_5_109/a_124_375# vdd 0.060786f
C1097 fanout79/a_36_160# _094_ 0.008308f
C1098 _419_/a_796_472# net77 0.001053f
C1099 _102_ mask\[2\] 0.036292f
C1100 _198_/a_67_603# _046_ 0.007349f
C1101 net57 _118_ 0.036179f
C1102 net2 rstn 0.002598f
C1103 FILLER_0_21_150/a_36_472# vdd 0.092128f
C1104 FILLER_0_21_150/a_124_375# vss 0.013882f
C1105 _162_ _058_ 0.015239f
C1106 mask\[0\] FILLER_0_12_196/a_124_375# 0.034009f
C1107 _430_/a_36_151# _091_ 0.02228f
C1108 fanout50/a_36_160# _383_/a_36_472# 0.096296f
C1109 _093_ FILLER_0_19_155/a_484_472# 0.001236f
C1110 _078_ _080_ 0.030094f
C1111 _412_/a_448_472# net81 0.047334f
C1112 net26 vss 0.263774f
C1113 _101_ _285_/a_244_68# 0.001153f
C1114 _035_ _446_/a_1000_472# 0.00349f
C1115 net29 _099_ 0.358926f
C1116 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2812_375# 0.001597f
C1117 FILLER_0_11_101/a_572_375# FILLER_0_10_107/a_36_472# 0.001684f
C1118 FILLER_0_7_72/a_932_472# net52 0.008749f
C1119 _127_ _128_ 0.257374f
C1120 net55 FILLER_0_17_56/a_484_472# 0.023554f
C1121 vdd output30/a_224_472# 0.068123f
C1122 _074_ net4 0.088616f
C1123 _131_ _058_ 0.031061f
C1124 FILLER_0_18_2/a_1828_472# _452_/a_448_472# 0.005748f
C1125 net34 _210_/a_67_603# 0.01049f
C1126 net81 net19 0.786284f
C1127 net54 FILLER_0_19_134/a_124_375# 0.002681f
C1128 FILLER_0_12_50/a_124_375# vss 0.004123f
C1129 FILLER_0_12_50/a_36_472# vdd 0.012805f
C1130 net38 net47 0.352245f
C1131 output28/a_224_472# result[1] 0.054333f
C1132 output31/a_224_472# _417_/a_2248_156# 0.024448f
C1133 _428_/a_2248_156# vdd 0.006977f
C1134 _098_ _433_/a_2248_156# 0.034774f
C1135 FILLER_0_20_193/a_572_375# net21 0.002103f
C1136 net38 _450_/a_1284_156# 0.001291f
C1137 FILLER_0_17_64/a_124_375# _183_ 0.001236f
C1138 net4 _076_ 1.140706f
C1139 _086_ _085_ 0.374127f
C1140 _437_/a_1000_472# net14 0.028506f
C1141 en_co_clk net53 0.001712f
C1142 _432_/a_448_472# _139_ 0.001772f
C1143 trim_mask\[4\] _158_ 0.022724f
C1144 _130_ cal_count\[3\] 0.037708f
C1145 _394_/a_56_524# vdd 0.010692f
C1146 _394_/a_728_93# vss 0.024106f
C1147 _161_ cal_count\[3\] 0.047389f
C1148 _432_/a_2248_156# mask\[3\] 0.002775f
C1149 _449_/a_448_472# FILLER_0_11_64/a_36_472# 0.001462f
C1150 net55 _175_ 0.142124f
C1151 net52 _032_ 0.009879f
C1152 _081_ FILLER_0_6_177/a_484_472# 0.010037f
C1153 _408_/a_728_93# net40 0.084147f
C1154 _105_ ctlp[2] 0.223601f
C1155 _422_/a_1204_472# _009_ 0.009783f
C1156 net44 _039_ 0.15647f
C1157 _132_ FILLER_0_14_107/a_1380_472# 0.049391f
C1158 _112_ calibrate 0.024557f
C1159 FILLER_0_8_107/a_36_472# _070_ 0.001287f
C1160 net41 FILLER_0_10_28/a_124_375# 0.003909f
C1161 output37/a_224_472# fanout65/a_36_113# 0.013171f
C1162 FILLER_0_11_124/a_124_375# _135_ 0.004831f
C1163 _098_ FILLER_0_15_235/a_124_375# 0.012702f
C1164 output17/a_224_472# net43 0.006661f
C1165 net52 trim_val\[4\] 0.21532f
C1166 _129_ cal_count\[3\] 0.005967f
C1167 _091_ FILLER_0_12_220/a_484_472# 0.001453f
C1168 _413_/a_1308_423# vdd 0.002686f
C1169 FILLER_0_20_177/a_36_472# _098_ 0.015061f
C1170 fanout78/a_36_113# net79 0.029496f
C1171 net20 _055_ 0.203142f
C1172 output35/a_224_472# mask\[6\] 0.069819f
C1173 result[7] FILLER_0_23_290/a_36_472# 0.013403f
C1174 net55 _452_/a_836_156# 0.010887f
C1175 _413_/a_36_151# FILLER_0_2_177/a_484_472# 0.006095f
C1176 FILLER_0_5_164/a_36_472# _386_/a_848_380# 0.001177f
C1177 _052_ FILLER_0_18_61/a_36_472# 0.001508f
C1178 _129_ _059_ 0.005414f
C1179 FILLER_0_14_81/a_124_375# _095_ 0.009791f
C1180 net66 net47 0.238874f
C1181 _068_ _311_/a_1212_473# 0.002835f
C1182 fanout77/a_36_113# net18 0.060158f
C1183 _111_ _303_/a_244_68# 0.001153f
C1184 _091_ _323_/a_36_113# 0.001651f
C1185 net20 _419_/a_1204_472# 0.006482f
C1186 mask\[5\] FILLER_0_19_195/a_124_375# 0.007169f
C1187 output42/a_224_472# net39 0.027208f
C1188 FILLER_0_4_177/a_36_472# _163_ 0.002787f
C1189 net54 _436_/a_2248_156# 0.043158f
C1190 _067_ net47 0.0609f
C1191 trim_mask\[1\] FILLER_0_6_47/a_1828_472# 0.007542f
C1192 _149_ _354_/a_49_472# 0.017453f
C1193 _424_/a_36_151# _012_ 0.005964f
C1194 _413_/a_2248_156# net21 0.009186f
C1195 _033_ _444_/a_36_151# 0.014843f
C1196 FILLER_0_18_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001684f
C1197 _360_/a_36_160# vss 0.028817f
C1198 _118_ _315_/a_244_497# 0.003007f
C1199 FILLER_0_8_2/a_124_375# vdd 0.016103f
C1200 _053_ net22 0.039386f
C1201 _144_ _022_ 0.139742f
C1202 FILLER_0_15_116/a_484_472# _136_ 0.002712f
C1203 net82 fanout52/a_36_160# 0.026154f
C1204 state\[0\] net64 0.01679f
C1205 net19 net30 0.311153f
C1206 FILLER_0_13_228/a_36_472# vdd 0.085375f
C1207 FILLER_0_13_228/a_124_375# vss 0.007465f
C1208 _088_ _073_ 0.001254f
C1209 FILLER_0_19_47/a_124_375# vdd 0.025971f
C1210 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001723f
C1211 _286_/a_224_472# _005_ 0.001254f
C1212 net18 _416_/a_1308_423# 0.021956f
C1213 _301_/a_36_472# FILLER_0_22_86/a_36_472# 0.010679f
C1214 mask\[8\] FILLER_0_22_86/a_124_375# 0.014263f
C1215 FILLER_0_15_10/a_36_472# vdd 0.086171f
C1216 FILLER_0_15_10/a_124_375# vss 0.002173f
C1217 _178_ FILLER_0_15_10/a_124_375# 0.002355f
C1218 net35 FILLER_0_22_128/a_484_472# 0.004578f
C1219 output19/a_224_472# ctlp[2] 0.04607f
C1220 net17 _452_/a_836_156# 0.002817f
C1221 _048_ _047_ 0.007849f
C1222 net35 _049_ 0.022439f
C1223 result[6] net33 0.363421f
C1224 _053_ FILLER_0_7_72/a_2276_472# 0.016004f
C1225 net20 FILLER_0_1_212/a_124_375# 0.084041f
C1226 FILLER_0_18_177/a_2812_375# net22 0.010501f
C1227 _096_ cal_count\[3\] 0.016393f
C1228 _185_ cal_count\[2\] 0.205002f
C1229 net41 FILLER_0_20_31/a_36_472# 0.030033f
C1230 _281_/a_672_472# _097_ 0.002131f
C1231 net60 _419_/a_2248_156# 0.047724f
C1232 net61 _419_/a_2560_156# 0.008214f
C1233 mask\[5\] FILLER_0_18_177/a_1828_472# 0.001038f
C1234 FILLER_0_8_127/a_124_375# _062_ 0.046401f
C1235 net20 FILLER_0_12_220/a_572_375# 0.007386f
C1236 net54 FILLER_0_22_128/a_1020_375# 0.010068f
C1237 FILLER_0_17_104/a_1380_472# vdd 0.010877f
C1238 _412_/a_2248_156# net65 0.039861f
C1239 _444_/a_796_472# net40 0.005776f
C1240 net4 _081_ 0.02226f
C1241 _070_ FILLER_0_9_105/a_572_375# 0.017191f
C1242 _013_ FILLER_0_18_37/a_1380_472# 0.01384f
C1243 FILLER_0_17_72/a_2812_375# _136_ 0.017702f
C1244 net58 net1 0.626432f
C1245 net34 _093_ 0.005701f
C1246 fanout70/a_36_113# FILLER_0_15_116/a_484_472# 0.002001f
C1247 _077_ _439_/a_36_151# 0.035432f
C1248 _086_ _062_ 0.066419f
C1249 _013_ FILLER_0_17_56/a_124_375# 0.001047f
C1250 net74 _067_ 0.674895f
C1251 _083_ vdd 0.157549f
C1252 _078_ vss 0.367953f
C1253 _115_ _131_ 0.410424f
C1254 FILLER_0_18_2/a_1916_375# net38 0.006403f
C1255 output10/a_224_472# vdd 0.107357f
C1256 FILLER_0_7_146/a_124_375# vdd 0.034288f
C1257 net52 trim_val\[3\] 0.082691f
C1258 _073_ cal_itt\[0\] 0.211566f
C1259 net24 _436_/a_36_151# 0.075327f
C1260 net55 FILLER_0_18_53/a_484_472# 0.012319f
C1261 FILLER_0_10_78/a_1020_375# net52 0.001158f
C1262 net65 net4 0.614946f
C1263 FILLER_0_2_111/a_36_472# _157_ 0.104961f
C1264 _176_ _390_/a_36_68# 0.005007f
C1265 _132_ FILLER_0_18_107/a_2364_375# 0.006403f
C1266 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_36_472# 0.001723f
C1267 trim_val\[3\] net49 0.009336f
C1268 _075_ _078_ 0.001896f
C1269 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1380_472# 0.013276f
C1270 _096_ _320_/a_672_472# 0.0082f
C1271 FILLER_0_13_65/a_36_472# fanout72/a_36_113# 0.193651f
C1272 trim_mask\[4\] _066_ 0.396509f
C1273 net34 _109_ 0.001298f
C1274 FILLER_0_8_107/a_124_375# _058_ 0.01823f
C1275 net1 _082_ 0.033169f
C1276 trim_val\[2\] net40 0.06019f
C1277 net82 net1 0.029512f
C1278 FILLER_0_20_193/a_484_472# vss 0.002439f
C1279 net47 _066_ 0.096823f
C1280 result[9] _417_/a_2665_112# 0.060365f
C1281 FILLER_0_17_72/a_2276_472# _131_ 0.004125f
C1282 trim_val\[0\] FILLER_0_6_47/a_572_375# 0.03235f
C1283 trim[0] trim[3] 0.012429f
C1284 FILLER_0_4_185/a_124_375# FILLER_0_4_177/a_572_375# 0.012001f
C1285 _420_/a_1000_472# _009_ 0.019219f
C1286 _141_ _343_/a_49_472# 0.04106f
C1287 FILLER_0_11_101/a_124_375# _058_ 0.002209f
C1288 _173_ _067_ 0.011854f
C1289 _158_ _154_ 0.008872f
C1290 _369_/a_36_68# _153_ 0.008048f
C1291 _053_ vdd 1.467835f
C1292 _056_ cal_count\[3\] 0.186969f
C1293 FILLER_0_12_136/a_1380_472# vss 0.031524f
C1294 FILLER_0_15_116/a_484_472# net53 0.002804f
C1295 _070_ _125_ 0.125523f
C1296 _076_ _058_ 0.912225f
C1297 FILLER_0_7_72/a_1380_472# net52 0.003507f
C1298 net68 FILLER_0_8_37/a_572_375# 0.011704f
C1299 net46 output46/a_224_472# 0.008691f
C1300 _438_/a_796_472# net71 0.00514f
C1301 cal_count\[3\] _453_/a_36_151# 0.023915f
C1302 net34 net54 0.003682f
C1303 net31 _106_ 0.035117f
C1304 result[7] FILLER_0_24_274/a_932_472# 0.006454f
C1305 trim_mask\[4\] net23 0.180803f
C1306 FILLER_0_12_136/a_1020_375# FILLER_0_11_142/a_484_472# 0.001543f
C1307 FILLER_0_18_177/a_2276_472# FILLER_0_19_195/a_124_375# 0.001684f
C1308 net73 FILLER_0_17_142/a_124_375# 0.003021f
C1309 FILLER_0_15_72/a_124_375# FILLER_0_15_59/a_572_375# 0.003228f
C1310 _233_/a_36_160# _445_/a_2248_156# 0.00136f
C1311 FILLER_0_5_54/a_932_472# vss 0.003426f
C1312 FILLER_0_5_54/a_1380_472# vdd 0.008983f
C1313 net23 net47 0.090948f
C1314 output21/a_224_472# output35/a_224_472# 0.001374f
C1315 _292_/a_36_160# net32 0.011466f
C1316 FILLER_0_17_72/a_36_472# net36 0.001121f
C1317 _077_ _426_/a_2665_112# 0.001392f
C1318 net58 result[0] 0.443436f
C1319 cal_count\[3\] FILLER_0_11_135/a_124_375# 0.004365f
C1320 _187_ _173_ 0.03421f
C1321 _093_ _438_/a_1308_423# 0.001057f
C1322 mask\[9\] _438_/a_448_472# 0.046823f
C1323 FILLER_0_5_164/a_124_375# vdd 0.00419f
C1324 _328_/a_36_113# _126_ 0.023932f
C1325 _026_ FILLER_0_20_87/a_124_375# 0.031902f
C1326 _251_/a_906_472# _070_ 0.002124f
C1327 _033_ _054_ 0.003394f
C1328 net15 FILLER_0_6_47/a_2276_472# 0.049487f
C1329 _182_ vdd 0.161134f
C1330 FILLER_0_10_28/a_36_472# net17 0.012954f
C1331 net25 _012_ 0.001747f
C1332 cal_itt\[3\] _055_ 0.007428f
C1333 FILLER_0_6_239/a_124_375# _317_/a_36_113# 0.002437f
C1334 _077_ _308_/a_692_472# 0.002268f
C1335 mask\[7\] _024_ 0.122185f
C1336 FILLER_0_18_177/a_2812_375# vdd 0.003766f
C1337 output10/a_224_472# net9 0.003212f
C1338 _449_/a_2665_112# _067_ 0.03661f
C1339 FILLER_0_21_133/a_36_472# _140_ 0.008378f
C1340 ctln[6] net13 0.065837f
C1341 _450_/a_836_156# _039_ 0.019042f
C1342 FILLER_0_11_101/a_572_375# cal_count\[3\] 0.002017f
C1343 net18 _419_/a_36_151# 0.021491f
C1344 net69 _384_/a_224_472# 0.002407f
C1345 net75 _425_/a_1000_472# 0.038919f
C1346 mask\[4\] FILLER_0_18_209/a_124_375# 0.020811f
C1347 net16 FILLER_0_18_37/a_1468_375# 0.002269f
C1348 FILLER_0_15_282/a_36_472# _006_ 0.003055f
C1349 net69 _441_/a_448_472# 0.028545f
C1350 _068_ _059_ 0.255081f
C1351 state\[1\] _225_/a_36_160# 0.0535f
C1352 output42/a_224_472# clkc 0.004924f
C1353 result[5] _094_ 0.065897f
C1354 _425_/a_36_151# vdd 0.078723f
C1355 FILLER_0_16_73/a_36_472# _176_ 0.013449f
C1356 net80 _024_ 0.064854f
C1357 FILLER_0_5_172/a_36_472# net47 0.0015f
C1358 net17 FILLER_0_20_15/a_36_472# 0.004375f
C1359 net73 FILLER_0_18_107/a_932_472# 0.016711f
C1360 _163_ FILLER_0_5_148/a_484_472# 0.002734f
C1361 _033_ vss 0.019158f
C1362 mask\[7\] FILLER_0_22_128/a_2812_375# 0.001476f
C1363 FILLER_0_24_96/a_124_375# net24 0.040364f
C1364 FILLER_0_15_142/a_124_375# net23 0.002212f
C1365 net4 _090_ 0.06324f
C1366 _415_/a_36_151# net79 0.001156f
C1367 FILLER_0_24_290/a_124_375# vss 0.034103f
C1368 FILLER_0_24_290/a_36_472# vdd 0.089567f
C1369 net53 _427_/a_448_472# 0.047356f
C1370 calibrate _120_ 0.001106f
C1371 _103_ _198_/a_67_603# 0.005362f
C1372 _057_ vss 0.169369f
C1373 state\[1\] FILLER_0_12_196/a_36_472# 0.030132f
C1374 _141_ _093_ 0.396041f
C1375 _448_/a_448_472# net22 0.085004f
C1376 net38 FILLER_0_12_2/a_484_472# 0.002706f
C1377 _428_/a_2665_112# _043_ 0.021483f
C1378 fanout74/a_36_113# vss 0.048756f
C1379 cal_itt\[2\] FILLER_0_3_221/a_1468_375# 0.016021f
C1380 net32 _011_ 0.072502f
C1381 net60 output18/a_224_472# 0.001518f
C1382 net50 _439_/a_36_151# 0.009774f
C1383 net52 _439_/a_1308_423# 0.033366f
C1384 _445_/a_2248_156# net49 0.029744f
C1385 _137_ vdd 0.945976f
C1386 fanout51/a_36_113# cal_count\[3\] 0.054567f
C1387 FILLER_0_24_130/a_36_472# ctlp[6] 0.005932f
C1388 _093_ net36 0.214976f
C1389 net74 net23 0.0064f
C1390 net81 output28/a_224_472# 0.01335f
C1391 FILLER_0_16_57/a_932_472# FILLER_0_15_59/a_572_375# 0.001543f
C1392 net27 _425_/a_2248_156# 0.027078f
C1393 _250_/a_36_68# vss 0.005108f
C1394 output36/a_224_472# vdd 0.145046f
C1395 _128_ _060_ 0.022833f
C1396 net79 net64 0.049663f
C1397 _013_ FILLER_0_18_53/a_124_375# 0.015996f
C1398 _180_ vss 0.106022f
C1399 _178_ _180_ 0.004668f
C1400 _432_/a_36_151# FILLER_0_17_161/a_36_472# 0.004847f
C1401 output26/a_224_472# net26 0.047008f
C1402 _443_/a_2248_156# _037_ 0.005717f
C1403 _443_/a_2560_156# _170_ 0.00758f
C1404 net15 _440_/a_1204_472# 0.01349f
C1405 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_932_472# 0.026657f
C1406 state\[2\] FILLER_0_13_142/a_932_472# 0.004118f
C1407 _105_ mask\[7\] 0.486236f
C1408 _091_ mask\[3\] 0.044304f
C1409 net16 _181_ 0.48682f
C1410 _091_ FILLER_0_13_212/a_36_472# 0.007355f
C1411 FILLER_0_7_72/a_2724_472# vdd 0.007669f
C1412 _114_ _127_ 0.006414f
C1413 _015_ FILLER_0_8_247/a_1020_375# 0.006994f
C1414 FILLER_0_18_2/a_1468_375# net55 0.007169f
C1415 _043_ cal_count\[0\] 0.019077f
C1416 _421_/a_448_472# net77 0.003958f
C1417 _432_/a_2665_112# FILLER_0_18_177/a_2276_472# 0.021761f
C1418 FILLER_0_3_78/a_36_472# vdd 0.082597f
C1419 FILLER_0_3_78/a_572_375# vss 0.04008f
C1420 FILLER_0_2_127/a_124_375# vss 0.008566f
C1421 FILLER_0_2_127/a_36_472# vdd 0.08468f
C1422 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_124_375# 0.012222f
C1423 _394_/a_728_93# _095_ 0.035417f
C1424 FILLER_0_24_274/a_1380_472# vss 0.005744f
C1425 _144_ net23 0.091811f
C1426 FILLER_0_17_104/a_1468_375# FILLER_0_16_115/a_124_375# 0.026339f
C1427 en_co_clk _389_/a_36_148# 0.001249f
C1428 FILLER_0_22_128/a_484_472# vdd 0.002467f
C1429 _297_/a_36_472# _295_/a_36_472# 0.004259f
C1430 FILLER_0_22_128/a_36_472# vss 0.001309f
C1431 _449_/a_2248_156# fanout55/a_36_160# 0.027388f
C1432 _186_ _407_/a_244_68# 0.001153f
C1433 FILLER_0_17_226/a_124_375# vdd 0.026497f
C1434 _049_ vdd 0.199608f
C1435 _020_ _131_ 0.011012f
C1436 _098_ _043_ 0.032706f
C1437 net20 _426_/a_2665_112# 0.018602f
C1438 _412_/a_36_151# output48/a_224_472# 0.229574f
C1439 _053_ fanout67/a_36_160# 0.05724f
C1440 net56 FILLER_0_18_139/a_572_375# 0.005919f
C1441 output27/a_224_472# FILLER_0_8_263/a_124_375# 0.011584f
C1442 result[5] net78 0.020038f
C1443 _441_/a_2248_156# FILLER_0_3_78/a_572_375# 0.001068f
C1444 _131_ _134_ 0.887647f
C1445 _410_/a_36_68# _120_ 0.073688f
C1446 _132_ FILLER_0_16_115/a_124_375# 0.033245f
C1447 _088_ FILLER_0_3_172/a_2276_472# 0.024532f
C1448 net34 _350_/a_49_472# 0.008001f
C1449 _086_ FILLER_0_7_104/a_932_472# 0.001786f
C1450 _425_/a_1308_423# net19 0.058462f
C1451 FILLER_0_9_28/a_3260_375# net68 0.009969f
C1452 _304_/a_224_472# vss 0.001746f
C1453 _065_ net52 0.017184f
C1454 _115_ _076_ 0.051404f
C1455 FILLER_0_16_241/a_124_375# mask\[2\] 0.027201f
C1456 net41 _186_ 0.054661f
C1457 ctlp[3] output20/a_224_472# 0.023589f
C1458 net82 FILLER_0_3_172/a_2364_375# 0.010439f
C1459 FILLER_0_7_72/a_36_472# vdd 0.106377f
C1460 output42/a_224_472# net47 0.083794f
C1461 _276_/a_36_160# vdd 0.010213f
C1462 _114_ FILLER_0_11_101/a_36_472# 0.00501f
C1463 net54 net36 0.005827f
C1464 FILLER_0_18_2/a_1468_375# net17 0.004803f
C1465 _065_ net49 0.001576f
C1466 _446_/a_448_472# vdd 0.006805f
C1467 _128_ _116_ 0.069335f
C1468 _127_ _176_ 0.319517f
C1469 net55 cal_count\[2\] 0.022989f
C1470 net79 _006_ 0.050445f
C1471 FILLER_0_6_177/a_484_472# _163_ 0.002256f
C1472 output48/a_224_472# _112_ 0.027383f
C1473 _322_/a_848_380# _126_ 0.002519f
C1474 _449_/a_36_151# FILLER_0_12_50/a_36_472# 0.003462f
C1475 net21 mask\[6\] 0.634881f
C1476 result[7] FILLER_0_23_282/a_572_375# 0.015853f
C1477 _152_ _059_ 0.038141f
C1478 FILLER_0_17_282/a_36_472# vss 0.007765f
C1479 output19/a_224_472# mask\[7\] 0.001181f
C1480 _316_/a_692_472# _122_ 0.002929f
C1481 _316_/a_1152_472# calibrate 0.001604f
C1482 FILLER_0_18_2/a_124_375# vss 0.003207f
C1483 FILLER_0_15_116/a_124_375# vdd 0.012886f
C1484 _026_ _098_ 0.197713f
C1485 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_36_472# 0.012267f
C1486 FILLER_0_9_142/a_36_472# _118_ 0.01533f
C1487 output20/a_224_472# net78 0.001495f
C1488 FILLER_0_18_2/a_3172_472# net40 0.046864f
C1489 _076_ _226_/a_860_68# 0.001752f
C1490 net27 FILLER_0_8_263/a_36_472# 0.003956f
C1491 _095_ FILLER_0_15_10/a_124_375# 0.023187f
C1492 _132_ FILLER_0_19_111/a_572_375# 0.01675f
C1493 _448_/a_448_472# vdd 0.02042f
C1494 net27 FILLER_0_14_235/a_572_375# 0.006429f
C1495 mask\[4\] _339_/a_36_160# 0.003234f
C1496 FILLER_0_3_142/a_124_375# net23 0.25251f
C1497 _413_/a_3041_156# net59 0.001022f
C1498 _257_/a_36_472# _074_ 0.011352f
C1499 FILLER_0_23_60/a_36_472# vss 0.006794f
C1500 net55 FILLER_0_19_28/a_484_472# 0.001426f
C1501 FILLER_0_3_142/a_36_472# trim_mask\[4\] 0.008297f
C1502 net15 net36 0.265646f
C1503 _440_/a_2665_112# FILLER_0_4_91/a_36_472# 0.007491f
C1504 FILLER_0_12_136/a_1380_472# _071_ 0.004003f
C1505 _128_ _118_ 0.58787f
C1506 _127_ _124_ 0.035569f
C1507 FILLER_0_18_100/a_36_472# vss 0.002412f
C1508 _104_ _010_ 0.252687f
C1509 FILLER_0_7_59/a_124_375# net68 0.019553f
C1510 _041_ FILLER_0_18_37/a_1468_375# 0.001032f
C1511 _016_ vss 0.069165f
C1512 FILLER_0_4_152/a_124_375# _170_ 0.029927f
C1513 _379_/a_244_68# _160_ 0.001202f
C1514 FILLER_0_5_54/a_124_375# net47 0.012889f
C1515 net55 _423_/a_2665_112# 0.002379f
C1516 net26 FILLER_0_21_28/a_1380_472# 0.035291f
C1517 _433_/a_1000_472# _145_ 0.004227f
C1518 _432_/a_2560_156# _139_ 0.002737f
C1519 FILLER_0_14_99/a_36_472# net14 0.036527f
C1520 FILLER_0_7_72/a_484_472# vss 0.003793f
C1521 cal_count\[2\] net17 0.074204f
C1522 _376_/a_36_160# FILLER_0_6_90/a_124_375# 0.005705f
C1523 FILLER_0_14_263/a_124_375# vss 0.007923f
C1524 FILLER_0_14_263/a_36_472# vdd 0.02759f
C1525 _028_ FILLER_0_7_72/a_124_375# 0.017052f
C1526 _043_ FILLER_0_15_180/a_124_375# 0.003099f
C1527 _010_ vss 0.064717f
C1528 net57 trim_mask\[4\] 0.259381f
C1529 _072_ _085_ 0.408915f
C1530 ctln[2] fanout81/a_36_160# 0.003798f
C1531 _386_/a_848_380# _169_ 0.001355f
C1532 _386_/a_124_24# _163_ 0.001234f
C1533 _236_/a_36_160# trim[1] 0.003604f
C1534 net23 FILLER_0_19_155/a_36_472# 0.019429f
C1535 _432_/a_2248_156# FILLER_0_18_177/a_1828_472# 0.035805f
C1536 FILLER_0_17_72/a_1020_375# vss 0.005441f
C1537 FILLER_0_17_72/a_1468_375# vdd 0.003316f
C1538 net57 net47 0.279638f
C1539 net58 net76 0.700034f
C1540 fanout49/a_36_160# _156_ 0.002871f
C1541 mask\[0\] _335_/a_665_69# 0.001711f
C1542 FILLER_0_4_107/a_1468_375# vdd 0.023541f
C1543 FILLER_0_15_142/a_124_375# fanout73/a_36_113# 0.00146f
C1544 _028_ FILLER_0_6_47/a_2276_472# 0.002066f
C1545 net4 FILLER_0_7_233/a_36_472# 0.036721f
C1546 FILLER_0_9_270/a_36_472# vdd 0.008742f
C1547 FILLER_0_9_270/a_572_375# vss 0.017196f
C1548 _032_ _370_/a_124_24# 0.007035f
C1549 net38 FILLER_0_20_2/a_484_472# 0.006727f
C1550 net17 _450_/a_448_472# 0.017832f
C1551 FILLER_0_16_241/a_36_472# _099_ 0.158391f
C1552 net52 FILLER_0_2_111/a_572_375# 0.00245f
C1553 _343_/a_257_69# _141_ 0.001515f
C1554 output19/a_224_472# _422_/a_2248_156# 0.011418f
C1555 _063_ _160_ 0.091185f
C1556 _105_ output34/a_224_472# 0.007506f
C1557 net52 _440_/a_448_472# 0.067294f
C1558 net60 _421_/a_1000_472# 0.035511f
C1559 net55 _043_ 0.053191f
C1560 fanout73/a_36_113# net74 0.04136f
C1561 input5/a_36_113# net59 0.257143f
C1562 FILLER_0_10_78/a_36_472# _120_ 0.004669f
C1563 _401_/a_36_68# _180_ 0.051459f
C1564 _179_ cal_count\[1\] 0.088667f
C1565 net20 net81 0.036173f
C1566 FILLER_0_16_89/a_484_472# _131_ 0.01075f
C1567 FILLER_0_10_78/a_1468_375# vdd 0.001778f
C1568 FILLER_0_16_107/a_572_375# _093_ 0.002827f
C1569 net50 FILLER_0_8_37/a_36_472# 0.059367f
C1570 FILLER_0_12_136/a_932_472# _126_ 0.014483f
C1571 FILLER_0_11_142/a_124_375# _120_ 0.036088f
C1572 _057_ _071_ 0.139904f
C1573 FILLER_0_23_282/a_36_472# vss 0.003317f
C1574 fanout64/a_36_160# fanout65/a_36_113# 0.001627f
C1575 _198_/a_67_603# mask\[2\] 0.005143f
C1576 FILLER_0_3_142/a_36_472# net74 0.001098f
C1577 mask\[7\] mask\[6\] 0.227476f
C1578 FILLER_0_13_142/a_36_472# vss 0.005768f
C1579 net49 _440_/a_448_472# 0.049861f
C1580 mask\[8\] mask\[7\] 0.021731f
C1581 net82 net76 0.061682f
C1582 net52 FILLER_0_5_72/a_1380_472# 0.001523f
C1583 FILLER_0_7_59/a_124_375# net67 0.036499f
C1584 FILLER_0_7_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001723f
C1585 _114_ trim_mask\[0\] 0.021887f
C1586 _061_ _062_ 0.344031f
C1587 FILLER_0_19_142/a_36_472# vdd 0.107105f
C1588 FILLER_0_19_142/a_124_375# vss 0.032026f
C1589 _040_ vdd 0.065702f
C1590 net74 _442_/a_1308_423# 0.001618f
C1591 FILLER_0_11_142/a_36_472# FILLER_0_13_142/a_124_375# 0.0027f
C1592 _062_ _311_/a_66_473# 0.027039f
C1593 _447_/a_448_472# vdd 0.014537f
C1594 _447_/a_36_151# vss 0.001541f
C1595 _250_/a_36_68# _071_ 0.199512f
C1596 cal_count\[3\] _113_ 0.093684f
C1597 FILLER_0_16_89/a_124_375# net36 0.011956f
C1598 FILLER_0_5_72/a_1380_472# net49 0.002057f
C1599 output45/a_224_472# trimb[2] 0.045907f
C1600 _413_/a_2665_112# FILLER_0_3_212/a_124_375# 0.001077f
C1601 net57 net74 2.360287f
C1602 net80 mask\[6\] 0.080689f
C1603 net20 _223_/a_36_160# 0.066119f
C1604 net50 _160_ 0.048787f
C1605 _137_ FILLER_0_16_154/a_572_375# 0.010132f
C1606 net63 _137_ 0.006317f
C1607 _089_ _272_/a_36_472# 0.003862f
C1608 net17 _043_ 0.571818f
C1609 _028_ FILLER_0_7_72/a_1468_375# 0.003785f
C1610 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_36_472# 0.086905f
C1611 FILLER_0_8_107/a_124_375# _134_ 0.007753f
C1612 FILLER_0_5_72/a_124_375# _440_/a_36_151# 0.059049f
C1613 net54 _433_/a_1308_423# 0.004372f
C1614 fanout54/a_36_160# _433_/a_2248_156# 0.012122f
C1615 net29 _196_/a_36_160# 0.073294f
C1616 FILLER_0_12_28/a_36_472# _450_/a_3129_107# 0.009814f
C1617 _450_/a_3129_107# net40 0.034729f
C1618 mask\[4\] FILLER_0_17_200/a_36_472# 0.001242f
C1619 _447_/a_2248_156# _441_/a_36_151# 0.035837f
C1620 net49 _034_ 0.031359f
C1621 output21/a_224_472# net21 0.011791f
C1622 net22 net12 0.032084f
C1623 _077_ _374_/a_36_68# 0.012411f
C1624 vdd FILLER_0_10_94/a_572_375# 0.02784f
C1625 _444_/a_36_151# _054_ 0.011342f
C1626 net46 net17 0.791341f
C1627 _144_ FILLER_0_19_155/a_484_472# 0.006137f
C1628 _072_ _062_ 0.025795f
C1629 net82 FILLER_0_2_177/a_124_375# 0.003837f
C1630 result[6] vdd 0.513079f
C1631 _093_ FILLER_0_18_177/a_2724_472# 0.003036f
C1632 _413_/a_2248_156# FILLER_0_1_212/a_36_472# 0.035805f
C1633 FILLER_0_5_109/a_484_472# _153_ 0.071582f
C1634 _320_/a_1120_472# _090_ 0.001215f
C1635 _140_ FILLER_0_21_150/a_36_472# 0.015502f
C1636 net56 FILLER_0_17_142/a_484_472# 0.008895f
C1637 _274_/a_36_68# _060_ 0.02117f
C1638 net20 net30 0.033149f
C1639 result[0] calibrate 0.00287f
C1640 FILLER_0_17_226/a_124_375# net63 0.00507f
C1641 net68 net17 0.601273f
C1642 _028_ FILLER_0_7_72/a_3260_375# 0.003505f
C1643 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_124_375# 0.003228f
C1644 _119_ FILLER_0_8_156/a_36_472# 0.010504f
C1645 _025_ _436_/a_1308_423# 0.006243f
C1646 _057_ _095_ 0.001346f
C1647 _432_/a_796_472# _091_ 0.018082f
C1648 net68 trim_val\[1\] 0.006974f
C1649 net75 FILLER_0_0_232/a_36_472# 0.001514f
C1650 FILLER_0_15_142/a_484_472# net56 0.003214f
C1651 FILLER_0_12_124/a_124_375# _131_ 0.07304f
C1652 _093_ FILLER_0_17_218/a_484_472# 0.004665f
C1653 _444_/a_36_151# vss 0.003795f
C1654 _444_/a_448_472# vdd 0.03285f
C1655 fanout81/a_36_160# net81 0.025745f
C1656 _448_/a_2248_156# _443_/a_2248_156# 0.006556f
C1657 FILLER_0_3_172/a_1916_375# net59 0.001221f
C1658 _412_/a_448_472# net59 0.001462f
C1659 output44/a_224_472# net44 0.051347f
C1660 FILLER_0_8_24/a_124_375# vdd 0.01166f
C1661 _077_ _133_ 0.003921f
C1662 fanout59/a_36_160# vdd 0.02169f
C1663 _095_ _180_ 0.013383f
C1664 _453_/a_1204_472# _042_ 0.002408f
C1665 _120_ _171_ 0.414533f
C1666 _136_ _172_ 0.024344f
C1667 net41 _063_ 0.105528f
C1668 cal_itt\[2\] net8 0.057335f
C1669 net19 net59 0.0206f
C1670 _414_/a_2248_156# net21 0.00415f
C1671 FILLER_0_12_136/a_124_375# net57 0.001727f
C1672 FILLER_0_2_93/a_572_375# vdd 0.022073f
C1673 _438_/a_36_151# net14 0.008367f
C1674 _080_ vss 0.012982f
C1675 output8/a_224_472# _411_/a_36_151# 0.12978f
C1676 FILLER_0_19_171/a_484_472# vdd 0.009225f
C1677 FILLER_0_19_171/a_36_472# vss 0.001338f
C1678 FILLER_0_15_150/a_36_472# net56 0.011741f
C1679 mask\[8\] _437_/a_448_472# 0.008198f
C1680 net57 FILLER_0_3_142/a_124_375# 0.003738f
C1681 _114_ _060_ 0.003352f
C1682 _053_ _385_/a_244_472# 0.00134f
C1683 net23 FILLER_0_5_148/a_124_375# 0.01836f
C1684 net60 net18 0.949607f
C1685 _306_/a_36_68# _055_ 0.006686f
C1686 _452_/a_3129_107# vss 0.00145f
C1687 _452_/a_2225_156# vdd 0.005612f
C1688 fanout56/a_36_113# vdd 0.078814f
C1689 _091_ _072_ 0.162027f
C1690 FILLER_0_6_239/a_124_375# _122_ 0.01772f
C1691 net47 FILLER_0_5_148/a_572_375# 0.062581f
C1692 output35/a_224_472# _435_/a_2248_156# 0.019736f
C1693 net16 _446_/a_2248_156# 0.010032f
C1694 FILLER_0_22_86/a_124_375# _026_ 0.001024f
C1695 _253_/a_36_68# cal_itt\[0\] 0.001495f
C1696 net67 net17 0.04175f
C1697 _359_/a_1044_488# _129_ 0.001111f
C1698 FILLER_0_23_44/a_1020_375# vdd -0.014642f
C1699 net15 _441_/a_36_151# 0.01821f
C1700 _415_/a_36_151# net19 0.05689f
C1701 _002_ _270_/a_244_68# 0.001153f
C1702 cal net2 0.081236f
C1703 net41 net50 0.002438f
C1704 output21/a_224_472# mask\[7\] 0.032297f
C1705 net12 vdd 0.082923f
C1706 _165_ trim_val\[0\] 0.164683f
C1707 _018_ vss 0.022336f
C1708 _440_/a_1204_472# net47 0.006257f
C1709 FILLER_0_5_109/a_36_472# net47 0.005565f
C1710 result[5] _418_/a_2248_156# 0.001309f
C1711 _418_/a_36_151# vdd 0.155643f
C1712 FILLER_0_4_177/a_36_472# net37 0.004017f
C1713 FILLER_0_14_107/a_36_472# vss 0.003706f
C1714 FILLER_0_14_107/a_484_472# vdd 0.030114f
C1715 result[7] vdd 0.500292f
C1716 _136_ FILLER_0_16_115/a_36_472# 0.013477f
C1717 _448_/a_36_151# FILLER_0_2_177/a_36_472# 0.04556f
C1718 FILLER_0_3_172/a_2364_375# net21 0.004803f
C1719 _306_/a_36_68# _126_ 0.01893f
C1720 FILLER_0_22_177/a_1020_375# net33 0.013731f
C1721 _433_/a_448_472# _022_ 0.074451f
C1722 _142_ net73 0.090025f
C1723 net36 _045_ 0.091033f
C1724 FILLER_0_18_2/a_2812_375# FILLER_0_20_15/a_1380_472# 0.001338f
C1725 net15 FILLER_0_9_60/a_484_472# 0.020589f
C1726 _395_/a_1044_488# _071_ 0.001198f
C1727 FILLER_0_21_286/a_124_375# vdd 0.026138f
C1728 _010_ _419_/a_1000_472# 0.001598f
C1729 _445_/a_448_472# net17 0.038794f
C1730 net64 net19 0.029763f
C1731 FILLER_0_4_177/a_572_375# _087_ 0.006527f
C1732 _114_ _116_ 0.038641f
C1733 _275_/a_224_472# mask\[3\] 0.002528f
C1734 _086_ _153_ 0.017325f
C1735 net2 en 0.067828f
C1736 net50 FILLER_0_7_59/a_572_375# 0.009554f
C1737 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_124_375# 0.001597f
C1738 net33 _204_/a_67_603# 0.022193f
C1739 mask\[4\] _202_/a_36_160# 0.007912f
C1740 ctln[3] vdd 0.167569f
C1741 output24/a_224_472# _025_ 0.010601f
C1742 net34 _144_ 0.029247f
C1743 net54 FILLER_0_22_86/a_1380_472# 0.059367f
C1744 _136_ FILLER_0_16_154/a_932_472# 0.008185f
C1745 _395_/a_36_488# _055_ 0.002775f
C1746 _334_/a_36_160# vdd 0.041716f
C1747 _016_ _095_ 0.034744f
C1748 _088_ FILLER_0_3_221/a_484_472# 0.002245f
C1749 comp net17 0.02802f
C1750 net48 _316_/a_848_380# 0.026413f
C1751 net35 _051_ 0.019252f
C1752 FILLER_0_14_81/a_124_375# net55 0.038949f
C1753 fanout80/a_36_113# _136_ 0.006151f
C1754 output26/a_224_472# FILLER_0_23_60/a_36_472# 0.003292f
C1755 _414_/a_1456_156# cal_itt\[3\] 0.001134f
C1756 _074_ FILLER_0_6_231/a_124_375# 0.006087f
C1757 vss _433_/a_2560_156# 0.003477f
C1758 _079_ _088_ 0.012529f
C1759 net16 FILLER_0_6_37/a_36_472# 0.013074f
C1760 FILLER_0_9_28/a_1380_472# _054_ 0.004017f
C1761 cal_count\[3\] FILLER_0_11_78/a_572_375# 0.010243f
C1762 ctlp[1] FILLER_0_24_274/a_572_375# 0.002408f
C1763 _005_ _044_ 0.50767f
C1764 input1/a_36_113# net2 0.018839f
C1765 FILLER_0_4_197/a_1380_472# net59 0.022002f
C1766 FILLER_0_3_172/a_36_472# net22 0.012287f
C1767 output7/a_224_472# ctln[9] 0.001987f
C1768 _114_ _118_ 0.074399f
C1769 _094_ _418_/a_2665_112# 0.035668f
C1770 _105_ _204_/a_255_603# 0.002146f
C1771 _422_/a_1308_423# mask\[7\] 0.045368f
C1772 FILLER_0_16_107/a_124_375# vdd 0.026251f
C1773 net5 vdd 0.516129f
C1774 result[6] _420_/a_1308_423# 0.008756f
C1775 cal valid 0.06045f
C1776 net34 FILLER_0_22_177/a_1380_472# 0.003953f
C1777 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_484_472# 0.026657f
C1778 _054_ vss 0.176655f
C1779 FILLER_0_9_60/a_484_472# net51 0.061362f
C1780 _070_ FILLER_0_6_231/a_36_472# 0.001096f
C1781 _076_ FILLER_0_6_231/a_124_375# 0.001382f
C1782 _091_ FILLER_0_17_218/a_572_375# 0.001927f
C1783 net20 _317_/a_36_113# 0.00189f
C1784 _058_ _117_ 0.003932f
C1785 _116_ _176_ 0.067051f
C1786 trim[4] net6 0.002404f
C1787 _432_/a_2665_112# _091_ 0.002978f
C1788 net19 _006_ 0.090449f
C1789 _445_/a_2248_156# net40 0.004545f
C1790 _321_/a_3126_472# _176_ 0.001932f
C1791 _069_ _395_/a_1492_488# 0.002565f
C1792 FILLER_0_16_37/a_124_375# cal_count\[2\] 0.008393f
C1793 _053_ FILLER_0_6_47/a_2364_375# 0.007053f
C1794 _093_ FILLER_0_17_72/a_1380_472# 0.008517f
C1795 _446_/a_36_151# output41/a_224_472# 0.135198f
C1796 _008_ _418_/a_2560_156# 0.006651f
C1797 _408_/a_56_524# _190_/a_36_160# 0.004025f
C1798 _408_/a_1336_472# _043_ 0.023648f
C1799 FILLER_0_15_235/a_484_472# vdd 0.006f
C1800 FILLER_0_15_235/a_36_472# vss 0.003138f
C1801 _436_/a_2665_112# FILLER_0_22_128/a_124_375# 0.004834f
C1802 _436_/a_2248_156# FILLER_0_22_128/a_572_375# 0.006739f
C1803 FILLER_0_15_235/a_124_375# mask\[1\] 0.013103f
C1804 FILLER_0_9_105/a_484_472# vss 0.004412f
C1805 FILLER_0_13_142/a_932_472# _043_ 0.011974f
C1806 _104_ vss 0.564464f
C1807 FILLER_0_20_177/a_1380_472# vdd 0.009871f
C1808 FILLER_0_20_177/a_932_472# vss 0.001272f
C1809 _178_ _278_/a_36_160# 0.269109f
C1810 net58 FILLER_0_9_290/a_124_375# 0.001157f
C1811 _103_ net19 0.047895f
C1812 _144_ _340_/a_36_160# 0.008886f
C1813 FILLER_0_1_266/a_124_375# net19 0.007016f
C1814 FILLER_0_5_54/a_572_375# FILLER_0_6_47/a_1380_472# 0.001597f
C1815 net44 vdd 0.897202f
C1816 output9/a_224_472# net8 0.020421f
C1817 _012_ net36 0.053654f
C1818 FILLER_0_16_57/a_572_375# FILLER_0_17_56/a_572_375# 0.026339f
C1819 fanout66/a_36_113# FILLER_0_3_54/a_36_472# 0.001645f
C1820 valid en 0.026142f
C1821 net48 net4 0.099614f
C1822 _105_ output18/a_224_472# 0.105478f
C1823 _178_ vss 0.150839f
C1824 _408_/a_728_93# _186_ 0.003815f
C1825 _432_/a_448_472# _093_ 0.048289f
C1826 net36 FILLER_0_15_212/a_36_472# 0.005396f
C1827 net52 fanout51/a_36_113# 0.036773f
C1828 _095_ FILLER_0_13_142/a_36_472# 0.001782f
C1829 FILLER_0_17_56/a_572_375# _183_ 0.002605f
C1830 _429_/a_2248_156# FILLER_0_15_212/a_1468_375# 0.001068f
C1831 cal_count\[3\] _042_ 0.001716f
C1832 _176_ _118_ 0.392531f
C1833 FILLER_0_20_98/a_36_472# net14 0.024154f
C1834 FILLER_0_20_15/a_1380_472# vdd 0.007068f
C1835 _189_/a_255_603# net64 0.002455f
C1836 _079_ cal_itt\[0\] 0.018495f
C1837 _092_ FILLER_0_17_218/a_124_375# 0.020704f
C1838 FILLER_0_18_107/a_1468_375# vdd 0.004726f
C1839 _098_ FILLER_0_21_150/a_124_375# 0.006526f
C1840 FILLER_0_4_107/a_36_472# _156_ 0.005297f
C1841 _076_ FILLER_0_8_239/a_36_472# 0.029514f
C1842 _289_/a_36_472# mask\[2\] 0.006392f
C1843 _321_/a_3126_472# _124_ 0.001072f
C1844 FILLER_0_12_50/a_124_375# cal_count\[0\] 0.002359f
C1845 _422_/a_1204_472# vdd 0.001062f
C1846 _075_ vss 0.046342f
C1847 FILLER_0_18_139/a_572_375# _145_ 0.00346f
C1848 net79 FILLER_0_12_220/a_1468_375# 0.012754f
C1849 _441_/a_2248_156# vss 0.005663f
C1850 _441_/a_2665_112# vdd 0.012404f
C1851 net76 net21 0.041873f
C1852 _430_/a_2248_156# mask\[2\] 0.009336f
C1853 _074_ _375_/a_692_497# 0.004556f
C1854 FILLER_0_15_142/a_124_375# net36 0.006533f
C1855 net34 ctlp[1] 0.127025f
C1856 net55 _424_/a_2248_156# 0.057967f
C1857 mask\[4\] FILLER_0_18_177/a_1020_375# 0.015941f
C1858 output48/a_224_472# net1 0.006536f
C1859 trim_val\[4\] _386_/a_848_380# 0.007605f
C1860 _412_/a_1204_472# net58 0.018724f
C1861 mask\[3\] FILLER_0_18_177/a_124_375# 0.002924f
C1862 _447_/a_1308_423# net68 0.006686f
C1863 _447_/a_36_151# _036_ 0.007244f
C1864 _414_/a_36_151# net76 0.037157f
C1865 net52 net69 0.372114f
C1866 _414_/a_2560_156# cal_itt\[3\] 0.007141f
C1867 fanout66/a_36_113# _164_ 0.010496f
C1868 _104_ _107_ 0.021508f
C1869 result[5] fanout60/a_36_160# 0.001585f
C1870 FILLER_0_18_139/a_484_472# FILLER_0_19_142/a_124_375# 0.001723f
C1871 FILLER_0_19_125/a_36_472# vss 0.001056f
C1872 FILLER_0_5_109/a_36_472# _154_ 0.070958f
C1873 net47 _452_/a_36_151# 0.021978f
C1874 _131_ FILLER_0_17_104/a_36_472# 0.004125f
C1875 _118_ _124_ 0.652002f
C1876 vss _107_ 0.186994f
C1877 net74 net36 0.012494f
C1878 net69 net49 0.051235f
C1879 _437_/a_36_151# vdd 0.115376f
C1880 FILLER_0_19_55/a_36_472# _013_ 0.005889f
C1881 FILLER_0_3_172/a_124_375# FILLER_0_2_171/a_124_375# 0.026339f
C1882 cal_itt\[3\] _374_/a_36_68# 0.001569f
C1883 _449_/a_796_472# _038_ 0.018626f
C1884 FILLER_0_3_172/a_36_472# vdd 0.006145f
C1885 FILLER_0_3_172/a_3260_375# vss 0.054783f
C1886 _306_/a_36_68# state\[1\] 0.028553f
C1887 FILLER_0_5_198/a_124_375# net21 0.029659f
C1888 FILLER_0_21_125/a_124_375# _433_/a_36_151# 0.059049f
C1889 output18/a_224_472# output19/a_224_472# 0.00124f
C1890 _141_ _144_ 0.095441f
C1891 FILLER_0_15_290/a_36_472# result[3] 0.014709f
C1892 FILLER_0_21_133/a_124_375# FILLER_0_21_125/a_572_375# 0.012001f
C1893 net41 _039_ 0.030362f
C1894 trimb[1] FILLER_0_18_2/a_36_472# 0.010728f
C1895 net16 _444_/a_2248_156# 0.065914f
C1896 _144_ _348_/a_49_472# 0.037768f
C1897 _264_/a_224_472# _084_ 0.007508f
C1898 cal_itt\[1\] cal_itt\[0\] 0.055355f
C1899 mask\[5\] net23 0.002188f
C1900 _052_ FILLER_0_18_37/a_1020_375# 0.001287f
C1901 FILLER_0_18_2/a_2724_472# _452_/a_448_472# 0.008967f
C1902 FILLER_0_10_28/a_36_472# output6/a_224_472# 0.010475f
C1903 FILLER_0_21_286/a_36_472# _420_/a_36_151# 0.059367f
C1904 net37 FILLER_0_5_148/a_484_472# 0.001212f
C1905 fanout76/a_36_160# vss 0.028897f
C1906 _414_/a_448_472# net76 0.002346f
C1907 FILLER_0_18_76/a_572_375# net71 0.006025f
C1908 vdd _416_/a_2665_112# 0.027256f
C1909 _043_ net21 0.033824f
C1910 _192_/a_67_603# _416_/a_2665_112# 0.012638f
C1911 FILLER_0_16_73/a_484_472# cal_count\[1\] 0.001135f
C1912 FILLER_0_12_136/a_36_472# _130_ 0.082451f
C1913 _422_/a_2665_112# _108_ 0.023365f
C1914 FILLER_0_5_88/a_124_375# vss 0.015423f
C1915 FILLER_0_5_88/a_36_472# vdd 0.090268f
C1916 FILLER_0_8_263/a_124_375# _426_/a_36_151# 0.001252f
C1917 FILLER_0_4_152/a_36_472# _386_/a_124_24# 0.004755f
C1918 _422_/a_2665_112# net19 0.006987f
C1919 _363_/a_36_68# _053_ 0.021227f
C1920 FILLER_0_10_214/a_36_472# _247_/a_36_160# 0.004828f
C1921 FILLER_0_7_195/a_36_472# _161_ 0.015074f
C1922 FILLER_0_11_142/a_484_472# cal_count\[3\] 0.014314f
C1923 FILLER_0_12_124/a_36_472# _127_ 0.01468f
C1924 FILLER_0_22_177/a_1468_375# mask\[6\] 0.002149f
C1925 net35 FILLER_0_22_177/a_1020_375# 0.008333f
C1926 _093_ FILLER_0_18_76/a_124_375# 0.061549f
C1927 _195_/a_67_603# vss 0.002638f
C1928 result[4] FILLER_0_15_290/a_36_472# 0.001422f
C1929 net80 FILLER_0_17_161/a_36_472# 0.003342f
C1930 ctln[8] output16/a_224_472# 0.006971f
C1931 _013_ FILLER_0_17_64/a_36_472# 0.001991f
C1932 FILLER_0_15_72/a_124_375# FILLER_0_13_72/a_36_472# 0.001418f
C1933 net15 _176_ 0.038396f
C1934 _055_ net22 0.084669f
C1935 _176_ FILLER_0_11_78/a_36_472# 0.003603f
C1936 FILLER_0_2_165/a_36_472# vss 0.001099f
C1937 FILLER_0_4_49/a_36_472# net49 0.010951f
C1938 net75 FILLER_0_8_247/a_1468_375# 0.047331f
C1939 FILLER_0_5_198/a_484_472# net22 0.012457f
C1940 result[1] FILLER_0_11_282/a_36_472# 0.01775f
C1941 _140_ _049_ 0.003069f
C1942 mask\[4\] FILLER_0_18_171/a_124_375# 0.008445f
C1943 _132_ _428_/a_1456_156# 0.001009f
C1944 FILLER_0_9_223/a_36_472# _128_ 0.00702f
C1945 _008_ net61 0.004059f
C1946 _395_/a_36_488# state\[1\] 0.002702f
C1947 _116_ _267_/a_36_472# 0.029316f
C1948 _025_ FILLER_0_22_107/a_124_375# 0.001891f
C1949 fanout71/a_36_113# net54 0.001194f
C1950 trim_mask\[1\] FILLER_0_6_90/a_484_472# 0.014443f
C1951 FILLER_0_2_177/a_484_472# net22 0.001324f
C1952 _031_ net14 0.00913f
C1953 output11/a_224_472# net59 0.002364f
C1954 _103_ _419_/a_448_472# 0.001207f
C1955 net72 FILLER_0_18_37/a_124_375# 0.05632f
C1956 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_36_472# 0.086635f
C1957 ctln[8] _447_/a_2665_112# 0.001271f
C1958 net20 _046_ 0.194455f
C1959 FILLER_0_14_107/a_932_472# _043_ 0.0017f
C1960 FILLER_0_13_100/a_124_375# vdd 0.039324f
C1961 _051_ vdd 0.036931f
C1962 net26 net55 0.002901f
C1963 output11/a_224_472# FILLER_0_0_198/a_124_375# 0.00363f
C1964 _033_ _166_ 0.004448f
C1965 _136_ FILLER_0_14_99/a_124_375# 0.007209f
C1966 result[8] net61 0.001106f
C1967 FILLER_0_5_117/a_124_375# net47 0.011773f
C1968 _415_/a_36_151# output28/a_224_472# 0.229574f
C1969 _184_ vss 0.068129f
C1970 state\[1\] FILLER_0_13_142/a_1468_375# 0.010245f
C1971 _178_ _184_ 0.436202f
C1972 trim_mask\[2\] net68 0.099597f
C1973 _128_ net74 0.121254f
C1974 _412_/a_36_151# net18 0.011383f
C1975 FILLER_0_11_101/a_484_472# FILLER_0_11_109/a_36_472# 0.013276f
C1976 _255_/a_224_552# _162_ 0.010564f
C1977 _057_ _375_/a_36_68# 0.003063f
C1978 _013_ _424_/a_796_472# 0.032857f
C1979 _095_ FILLER_0_14_107/a_36_472# 0.011439f
C1980 _420_/a_796_472# vss 0.001659f
C1981 net16 net51 0.035455f
C1982 output22/a_224_472# ctlp[4] 0.008275f
C1983 fanout73/a_36_113# net70 0.00238f
C1984 _435_/a_2248_156# net21 0.012406f
C1985 _141_ FILLER_0_19_155/a_36_472# 0.05777f
C1986 _359_/a_1044_488# _152_ 0.001339f
C1987 net4 FILLER_0_12_220/a_36_472# 0.019348f
C1988 FILLER_0_8_138/a_36_472# vss 0.008189f
C1989 FILLER_0_10_28/a_124_375# _450_/a_3129_107# 0.010735f
C1990 _444_/a_1308_423# net67 0.021684f
C1991 _177_ _451_/a_2449_156# 0.002085f
C1992 _360_/a_36_160# _070_ 0.012463f
C1993 net72 _394_/a_718_524# 0.001558f
C1994 net55 _394_/a_728_93# 0.0026f
C1995 _136_ _139_ 0.394888f
C1996 net52 _443_/a_1308_423# 0.02003f
C1997 trim_mask\[2\] _156_ 0.018332f
C1998 _446_/a_2560_156# net66 0.002649f
C1999 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_124_375# 0.009654f
C2000 _071_ vss 0.126519f
C2001 net35 _436_/a_36_151# 0.014669f
C2002 _143_ mask\[3\] 0.023322f
C2003 net63 _430_/a_796_472# 0.002914f
C2004 _305_/a_36_159# _316_/a_124_24# 0.003478f
C2005 FILLER_0_3_78/a_124_375# _160_ 0.003276f
C2006 net48 _251_/a_244_472# 0.001259f
C2007 _322_/a_692_472# _070_ 0.002328f
C2008 _233_/a_36_160# FILLER_0_6_37/a_124_375# 0.001713f
C2009 net26 net17 0.132516f
C2010 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_36_472# 0.026657f
C2011 _077_ FILLER_0_10_94/a_484_472# 0.001548f
C2012 net63 FILLER_0_20_177/a_1380_472# 0.011079f
C2013 ctln[5] FILLER_0_1_192/a_124_375# 0.001391f
C2014 net40 _034_ 0.04333f
C2015 _076_ FILLER_0_8_156/a_484_472# 0.008487f
C2016 net57 net70 0.012088f
C2017 FILLER_0_16_89/a_124_375# _176_ 0.002781f
C2018 _131_ cal_count\[1\] 0.001497f
C2019 _316_/a_848_380# net37 0.01216f
C2020 FILLER_0_20_193/a_484_472# _098_ 0.012457f
C2021 FILLER_0_21_142/a_124_375# net54 0.027551f
C2022 FILLER_0_20_177/a_1020_375# _434_/a_36_151# 0.059049f
C2023 FILLER_0_4_99/a_124_375# vdd 0.029154f
C2024 _185_ _180_ 0.001053f
C2025 FILLER_0_16_154/a_1468_375# vdd 0.017574f
C2026 FILLER_0_16_154/a_1020_375# vss 0.001453f
C2027 _068_ _229_/a_224_472# 0.002601f
C2028 net41 net72 0.319547f
C2029 _027_ vss 0.011873f
C2030 _055_ vdd 0.406945f
C2031 _424_/a_36_151# _423_/a_1308_423# 0.001722f
C2032 FILLER_0_20_193/a_484_472# _205_/a_36_160# 0.001684f
C2033 net22 _204_/a_67_603# 0.006495f
C2034 _389_/a_36_148# _172_ 0.039684f
C2035 result[6] net77 0.111093f
C2036 FILLER_0_22_86/a_484_472# net14 0.006746f
C2037 _077_ _122_ 0.144611f
C2038 _144_ _433_/a_1308_423# 0.027969f
C2039 _386_/a_124_24# net37 0.00431f
C2040 _420_/a_2248_156# _108_ 0.021735f
C2041 _177_ net36 0.371814f
C2042 _086_ FILLER_0_6_177/a_36_472# 0.064045f
C2043 _004_ _101_ 0.001514f
C2044 _092_ _093_ 0.287983f
C2045 FILLER_0_17_161/a_124_375# mask\[2\] 0.00227f
C2046 FILLER_0_2_177/a_484_472# vdd 0.008489f
C2047 _077_ _227_/a_36_160# 0.012587f
C2048 net19 _420_/a_2248_156# 0.058662f
C2049 FILLER_0_16_89/a_1468_375# _093_ 0.003988f
C2050 FILLER_0_13_142/a_1380_472# _225_/a_36_160# 0.004111f
C2051 FILLER_0_9_28/a_2276_472# _453_/a_36_151# 0.059367f
C2052 FILLER_0_15_116/a_124_375# _451_/a_36_151# 0.006111f
C2053 mask\[1\] _043_ 0.027561f
C2054 output36/a_224_472# output30/a_224_472# 0.003578f
C2055 net76 FILLER_0_3_172/a_484_472# 0.002542f
C2056 _050_ net14 0.001835f
C2057 _095_ _278_/a_36_160# 0.030448f
C2058 mask\[8\] _354_/a_49_472# 0.105272f
C2059 _413_/a_36_151# net59 0.02781f
C2060 FILLER_0_8_138/a_124_375# _076_ 0.031436f
C2061 _126_ vdd 0.682779f
C2062 net20 _256_/a_716_497# 0.007413f
C2063 _093_ FILLER_0_17_142/a_572_375# 0.009547f
C2064 _019_ net36 0.309649f
C2065 _096_ _335_/a_257_69# 0.001084f
C2066 FILLER_0_13_206/a_124_375# net4 0.031251f
C2067 net53 FILLER_0_14_99/a_124_375# 0.00494f
C2068 FILLER_0_13_212/a_1020_375# net79 0.009597f
C2069 net62 FILLER_0_13_212/a_1468_375# 0.003327f
C2070 net4 net37 0.021795f
C2071 _095_ vss 1.465527f
C2072 _178_ _095_ 0.839141f
C2073 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_124_375# 0.001597f
C2074 _430_/a_36_151# FILLER_0_18_177/a_3172_472# 0.001512f
C2075 FILLER_0_19_47/a_124_375# _182_ 0.001771f
C2076 net4 FILLER_0_3_221/a_1468_375# 0.006974f
C2077 _261_/a_36_160# net23 0.005015f
C2078 mask\[7\] _435_/a_2248_156# 0.026974f
C2079 net27 _274_/a_244_497# 0.010334f
C2080 net76 FILLER_0_5_181/a_124_375# 0.031324f
C2081 net20 net59 0.045227f
C2082 FILLER_0_1_212/a_124_375# vdd 0.020159f
C2083 mask\[5\] FILLER_0_19_155/a_484_472# 0.043011f
C2084 _011_ net78 0.002956f
C2085 _036_ vss 0.161195f
C2086 FILLER_0_10_78/a_572_375# vss 0.004588f
C2087 cal_count\[1\] FILLER_0_13_80/a_36_472# 0.001559f
C2088 FILLER_0_21_142/a_484_472# FILLER_0_22_128/a_1916_375# 0.001543f
C2089 _084_ net8 0.001821f
C2090 output26/a_224_472# vss 0.0137f
C2091 FILLER_0_12_220/a_572_375# vdd -0.014642f
C2092 FILLER_0_24_96/a_124_375# net35 0.001886f
C2093 FILLER_0_12_220/a_124_375# vss 0.040895f
C2094 FILLER_0_12_136/a_484_472# _076_ 0.001683f
C2095 fanout50/a_36_160# _447_/a_2665_112# 0.002885f
C2096 _426_/a_1000_472# calibrate 0.002865f
C2097 FILLER_0_18_139/a_932_472# vdd 0.002904f
C2098 FILLER_0_18_139/a_484_472# vss 0.006719f
C2099 FILLER_0_4_123/a_36_472# _370_/a_124_24# 0.003595f
C2100 _053_ FILLER_0_7_146/a_124_375# 0.005844f
C2101 _408_/a_1936_472# _067_ 0.003007f
C2102 FILLER_0_9_72/a_1380_472# _439_/a_36_151# 0.001723f
C2103 _093_ FILLER_0_18_107/a_1380_472# 0.001782f
C2104 FILLER_0_15_282/a_484_472# net18 0.018113f
C2105 trim_val\[3\] _168_ 0.271475f
C2106 FILLER_0_5_72/a_124_375# _029_ 0.010208f
C2107 FILLER_0_5_117/a_124_375# _154_ 0.005866f
C2108 FILLER_0_22_177/a_1020_375# vdd 0.001695f
C2109 FILLER_0_18_107/a_932_472# mask\[9\] 0.005296f
C2110 _415_/a_1000_472# net19 0.001125f
C2111 net19 _419_/a_2665_112# 0.00276f
C2112 output48/a_224_472# net76 0.069862f
C2113 state\[1\] net22 0.007096f
C2114 _110_ mask\[9\] 0.00319f
C2115 cal cal_itt\[1\] 0.036277f
C2116 _390_/a_244_472# _038_ 0.001278f
C2117 _390_/a_36_68# _136_ 0.032598f
C2118 _447_/a_2248_156# _030_ 0.001588f
C2119 FILLER_0_18_139/a_124_375# FILLER_0_18_107/a_3260_375# 0.012552f
C2120 cal_count\[2\] _179_ 0.404284f
C2121 _081_ FILLER_0_8_156/a_484_472# 0.001772f
C2122 _426_/a_796_472# net64 0.006933f
C2123 net81 FILLER_0_9_270/a_124_375# 0.014206f
C2124 FILLER_0_4_107/a_572_375# _160_ 0.008945f
C2125 FILLER_0_17_282/a_124_375# net30 0.001288f
C2126 mask\[3\] _341_/a_49_472# 0.00631f
C2127 FILLER_0_1_192/a_124_375# net59 0.014491f
C2128 _187_ _408_/a_1936_472# 0.017573f
C2129 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_124_375# 0.003732f
C2130 _418_/a_36_151# net77 0.019316f
C2131 net3 cal_count\[2\] 0.119728f
C2132 result[7] net77 0.005269f
C2133 FILLER_0_17_72/a_124_375# _131_ 0.006224f
C2134 _081_ _265_/a_916_472# 0.002264f
C2135 _204_/a_67_603# vdd 0.039556f
C2136 _435_/a_1288_156# vdd 0.001119f
C2137 net20 _122_ 0.046817f
C2138 _431_/a_796_472# _137_ 0.002195f
C2139 _367_/a_244_472# vdd 0.001113f
C2140 _449_/a_1308_423# vdd 0.002584f
C2141 _449_/a_448_472# vss 0.032274f
C2142 _405_/a_67_603# net47 0.004116f
C2143 _431_/a_2560_156# net56 0.001258f
C2144 _153_ _365_/a_692_472# 0.002377f
C2145 FILLER_0_21_286/a_124_375# net77 0.00301f
C2146 net20 FILLER_0_7_233/a_124_375# 0.017217f
C2147 result[6] _421_/a_448_472# 0.038671f
C2148 _410_/a_244_472# _042_ 0.003902f
C2149 _443_/a_1204_472# net23 0.026261f
C2150 result[1] vdd 0.221634f
C2151 _431_/a_2248_156# vdd 0.00968f
C2152 net4 _264_/a_224_472# 0.001408f
C2153 en cal_itt\[1\] 0.028447f
C2154 input3/a_36_113# net3 0.015124f
C2155 _443_/a_2248_156# trim_mask\[4\] 0.002315f
C2156 _255_/a_224_552# _074_ 0.005907f
C2157 _004_ _094_ 0.213913f
C2158 _126_ _135_ 0.011447f
C2159 mask\[9\] _437_/a_2665_112# 0.014146f
C2160 _026_ _437_/a_448_472# 0.026072f
C2161 net20 net64 0.374636f
C2162 vss output41/a_224_472# -0.007739f
C2163 FILLER_0_9_28/a_484_472# net40 0.020293f
C2164 fanout49/a_36_160# FILLER_0_3_78/a_572_375# 0.00805f
C2165 _451_/a_36_151# _040_ 0.018648f
C2166 trim_mask\[1\] net14 0.024935f
C2167 _053_ FILLER_0_5_54/a_1380_472# 0.00114f
C2168 net15 FILLER_0_17_64/a_124_375# 0.047331f
C2169 _122_ FILLER_0_6_231/a_572_375# 0.016091f
C2170 net75 _305_/a_36_159# 0.049563f
C2171 _346_/a_49_472# vss 0.0031f
C2172 _131_ _120_ 0.191602f
C2173 FILLER_0_14_263/a_36_472# output30/a_224_472# 0.002002f
C2174 _031_ _153_ 0.009316f
C2175 _255_/a_224_552# _076_ 0.081663f
C2176 _057_ _070_ 0.033401f
C2177 _016_ _428_/a_2665_112# 0.050481f
C2178 FILLER_0_16_73/a_484_472# _175_ 0.036868f
C2179 _402_/a_728_93# vdd 0.050988f
C2180 _178_ _402_/a_1296_93# 0.062418f
C2181 FILLER_0_7_233/a_36_472# FILLER_0_6_231/a_124_375# 0.001684f
C2182 _432_/a_2560_156# _093_ 0.007613f
C2183 trim_mask\[1\] _164_ 0.195956f
C2184 net82 _078_ 0.00197f
C2185 net50 FILLER_0_8_24/a_36_472# 0.015187f
C2186 mask\[4\] FILLER_0_19_171/a_572_375# 0.006277f
C2187 ctln[5] output12/a_224_472# 0.069673f
C2188 _068_ _247_/a_36_160# 0.003213f
C2189 FILLER_0_12_236/a_36_472# vss 0.001526f
C2190 FILLER_0_12_236/a_484_472# vdd 0.00923f
C2191 cal_itt\[2\] _073_ 0.202415f
C2192 output37/a_224_472# vss 0.026983f
C2193 FILLER_0_15_282/a_36_472# _417_/a_1308_423# 0.001295f
C2194 FILLER_0_14_91/a_36_472# vss 0.001729f
C2195 FILLER_0_14_91/a_484_472# vdd 0.00605f
C2196 _157_ net14 0.026868f
C2197 _105_ _048_ 0.02699f
C2198 _385_/a_36_68# vss 0.002408f
C2199 _442_/a_796_472# _031_ 0.013039f
C2200 _372_/a_170_472# _059_ 0.033956f
C2201 FILLER_0_21_28/a_1828_472# vdd 0.004227f
C2202 FILLER_0_21_28/a_1380_472# vss 0.001688f
C2203 _436_/a_36_151# vdd 0.078019f
C2204 mask\[0\] _043_ 0.929722f
C2205 net50 FILLER_0_2_93/a_484_472# 0.002377f
C2206 FILLER_0_3_221/a_124_375# vdd 0.008869f
C2207 trimb[1] FILLER_0_19_28/a_124_375# 0.00285f
C2208 _423_/a_796_472# _012_ 0.015809f
C2209 ctlp[6] mask\[7\] 0.011418f
C2210 FILLER_0_17_282/a_124_375# _417_/a_36_151# 0.059049f
C2211 FILLER_0_1_192/a_36_472# net21 0.016033f
C2212 FILLER_0_13_100/a_36_472# _043_ 0.012726f
C2213 _411_/a_36_151# _000_ 0.023297f
C2214 net36 _438_/a_448_472# 0.034338f
C2215 ctlp[7] _050_ 0.153673f
C2216 mask\[9\] net14 0.090939f
C2217 _439_/a_36_151# vdd 0.095368f
C2218 net36 _451_/a_2225_156# 0.044144f
C2219 net54 _437_/a_2560_156# 0.009745f
C2220 _013_ _052_ 0.284735f
C2221 net20 _006_ 0.014721f
C2222 mask\[3\] fanout63/a_36_160# 0.002585f
C2223 net47 FILLER_0_5_136/a_36_472# 0.006139f
C2224 FILLER_0_21_28/a_1916_375# _424_/a_36_151# 0.059049f
C2225 _256_/a_244_497# _128_ 0.002372f
C2226 net79 result[3] 0.138076f
C2227 state\[1\] vdd 0.544231f
C2228 net15 _030_ 0.355335f
C2229 FILLER_0_14_50/a_124_375# _180_ 0.022435f
C2230 _050_ _148_ 0.002456f
C2231 net1 fanout58/a_36_160# 0.060243f
C2232 _085_ net23 0.020463f
C2233 net3 _043_ 0.004313f
C2234 _095_ _184_ 0.265966f
C2235 net34 mask\[5\] 0.041303f
C2236 net69 _370_/a_124_24# 0.001491f
C2237 _095_ _401_/a_36_68# 0.001398f
C2238 net20 _103_ 0.261438f
C2239 _007_ vdd 0.129966f
C2240 _064_ net49 0.377675f
C2241 _321_/a_358_69# net23 0.001718f
C2242 _449_/a_2248_156# cal_count\[3\] 0.002041f
C2243 net16 net47 0.089651f
C2244 net28 _416_/a_2665_112# 0.008877f
C2245 _104_ _106_ 0.17237f
C2246 _428_/a_2665_112# FILLER_0_13_142/a_36_472# 0.003706f
C2247 ctln[0] trim[2] 0.011834f
C2248 FILLER_0_0_266/a_124_375# vdd 0.006328f
C2249 fanout75/a_36_113# net1 0.011428f
C2250 _274_/a_36_68# FILLER_0_12_220/a_932_472# 0.001237f
C2251 _096_ net79 0.015605f
C2252 output23/a_224_472# vdd 0.033718f
C2253 _412_/a_36_151# net65 0.015454f
C2254 _112_ _081_ 0.037903f
C2255 FILLER_0_16_57/a_1468_375# _176_ 0.006445f
C2256 FILLER_0_7_72/a_2724_472# _053_ 0.016187f
C2257 result[7] _421_/a_448_472# 0.018021f
C2258 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_36_472# 0.001723f
C2259 _106_ vss 0.180823f
C2260 output7/a_224_472# net7 0.01565f
C2261 cal_itt\[3\] net59 0.018616f
C2262 result[8] FILLER_0_23_274/a_36_472# 0.001908f
C2263 _431_/a_1000_472# _136_ 0.024253f
C2264 _131_ FILLER_0_17_56/a_484_472# 0.002672f
C2265 FILLER_0_3_142/a_36_472# _261_/a_36_160# 0.001542f
C2266 net67 output6/a_224_472# 0.070024f
C2267 _114_ net74 0.559239f
C2268 _033_ net17 0.028529f
C2269 output32/a_224_472# _418_/a_448_472# 0.008149f
C2270 result[4] net79 0.048452f
C2271 net18 FILLER_0_11_282/a_124_375# 0.042342f
C2272 _256_/a_1164_497# _076_ 0.001871f
C2273 _370_/a_124_24# _152_ 0.069015f
C2274 _370_/a_848_380# _081_ 0.035068f
C2275 FILLER_0_13_65/a_124_375# _043_ 0.013045f
C2276 _167_ _160_ 0.157458f
C2277 FILLER_0_21_125/a_572_375# net54 0.024701f
C2278 ctln[2] vdd 0.245598f
C2279 net60 _418_/a_796_472# 0.008602f
C2280 trim[1] net66 0.007756f
C2281 _413_/a_2248_156# net65 0.036792f
C2282 net24 FILLER_0_23_88/a_124_375# 0.020193f
C2283 FILLER_0_24_130/a_124_375# net54 0.001269f
C2284 FILLER_0_15_142/a_572_375# net56 0.001809f
C2285 _069_ _055_ 0.741952f
C2286 _426_/a_2248_156# vss 0.002303f
C2287 _426_/a_2665_112# vdd 0.008893f
C2288 _070_ _310_/a_49_472# 0.00564f
C2289 _147_ vss 0.006333f
C2290 FILLER_0_16_107/a_484_472# _132_ 0.005391f
C2291 _065_ _168_ 0.020406f
C2292 net74 FILLER_0_5_136/a_36_472# 0.003704f
C2293 mask\[5\] _340_/a_36_160# 0.031249f
C2294 _175_ _131_ 0.050098f
C2295 _432_/a_1000_472# vdd 0.010431f
C2296 _444_/a_2665_112# _164_ 0.015644f
C2297 FILLER_0_7_72/a_36_472# _053_ 0.01287f
C2298 _176_ FILLER_0_15_59/a_484_472# 0.007596f
C2299 output27/a_224_472# FILLER_0_9_282/a_484_472# 0.001711f
C2300 net50 FILLER_0_4_91/a_572_375# 0.007234f
C2301 FILLER_0_24_96/a_124_375# vdd 0.029269f
C2302 net29 _287_/a_36_472# 0.002936f
C2303 output12/a_224_472# net59 0.015069f
C2304 net70 net36 0.066607f
C2305 FILLER_0_24_130/a_36_472# vss 0.001687f
C2306 _430_/a_1204_472# _091_ 0.007301f
C2307 fanout74/a_36_113# net82 0.018392f
C2308 cal_itt\[3\] _122_ 0.03282f
C2309 _176_ net74 0.067915f
C2310 net81 net22 0.064261f
C2311 output12/a_224_472# FILLER_0_0_198/a_124_375# 0.00515f
C2312 FILLER_0_6_47/a_2812_375# vss 0.035758f
C2313 FILLER_0_6_47/a_3260_375# vdd 0.003435f
C2314 FILLER_0_14_107/a_484_472# _451_/a_36_151# 0.001723f
C2315 net79 _056_ 0.022406f
C2316 net15 FILLER_0_15_72/a_124_375# 0.006566f
C2317 net18 FILLER_0_13_290/a_36_472# 0.079901f
C2318 _332_/a_244_68# _135_ 0.001325f
C2319 ctln[6] FILLER_0_0_130/a_36_472# 0.023355f
C2320 net31 output34/a_224_472# 0.165772f
C2321 net63 FILLER_0_22_177/a_1020_375# 0.003419f
C2322 cal_count\[2\] _402_/a_56_567# 0.07745f
C2323 _089_ _087_ 0.002217f
C2324 _402_/a_1296_93# _401_/a_36_68# 0.001523f
C2325 net36 FILLER_0_15_228/a_124_375# 0.00167f
C2326 FILLER_0_4_99/a_36_472# _156_ 0.0255f
C2327 FILLER_0_13_212/a_124_375# vdd 0.010978f
C2328 _104_ _421_/a_1308_423# 0.001621f
C2329 output31/a_224_472# net62 0.030092f
C2330 FILLER_0_4_197/a_124_375# net76 0.00811f
C2331 FILLER_0_6_90/a_36_472# net14 0.002705f
C2332 fanout67/a_36_160# _439_/a_36_151# 0.00246f
C2333 _050_ _436_/a_2665_112# 0.030939f
C2334 _062_ net23 0.061239f
C2335 FILLER_0_12_136/a_124_375# _114_ 0.006974f
C2336 output38/a_224_472# net49 0.002434f
C2337 FILLER_0_11_101/a_124_375# _120_ 0.008016f
C2338 _086_ cal_count\[3\] 0.259095f
C2339 net74 _124_ 0.180235f
C2340 result[9] FILLER_0_24_274/a_36_472# 0.009425f
C2341 _446_/a_36_151# net17 0.006518f
C2342 FILLER_0_7_72/a_932_472# _077_ 0.001315f
C2343 _076_ _120_ 0.736844f
C2344 net16 _173_ 0.029412f
C2345 ctln[2] net9 0.022757f
C2346 net79 _286_/a_224_472# 0.001276f
C2347 _025_ net71 0.030824f
C2348 FILLER_0_17_226/a_36_472# mask\[3\] 0.011509f
C2349 FILLER_0_8_37/a_572_375# _054_ 0.137749f
C2350 result[8] FILLER_0_24_274/a_1468_375# 0.00726f
C2351 mask\[5\] _141_ 0.241158f
C2352 _424_/a_2560_156# vss 0.001554f
C2353 vdd FILLER_0_21_60/a_124_375# 0.014029f
C2354 trimb[4] FILLER_0_18_2/a_36_472# 0.001673f
C2355 net4 net8 0.00647f
C2356 _265_/a_244_68# net59 0.001147f
C2357 mask\[5\] _348_/a_49_472# 0.025962f
C2358 net55 FILLER_0_17_72/a_1020_375# 0.049648f
C2359 _422_/a_36_151# _421_/a_2248_156# 0.001189f
C2360 mask\[4\] _293_/a_36_472# 0.023203f
C2361 _093_ FILLER_0_17_104/a_1020_375# 0.01418f
C2362 _132_ net71 0.099427f
C2363 _431_/a_36_151# _136_ 0.03371f
C2364 FILLER_0_9_223/a_572_375# _055_ 0.022619f
C2365 FILLER_0_16_107/a_124_375# _451_/a_36_151# 0.001597f
C2366 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_124_375# 0.026339f
C2367 _377_/a_36_472# _165_ 0.025689f
C2368 mask\[9\] _148_ 0.01635f
C2369 FILLER_0_5_109/a_36_472# _365_/a_36_68# 0.07596f
C2370 output29/a_224_472# _045_ 0.002303f
C2371 FILLER_0_6_239/a_36_472# fanout75/a_36_113# 0.00191f
C2372 FILLER_0_16_57/a_932_472# net15 0.037807f
C2373 _207_/a_67_603# FILLER_0_22_128/a_3172_472# 0.005759f
C2374 FILLER_0_8_37/a_572_375# vss 0.00282f
C2375 FILLER_0_8_37/a_36_472# vdd 0.135405f
C2376 result[9] FILLER_0_15_282/a_36_472# 0.003213f
C2377 net65 FILLER_0_3_212/a_124_375# 0.003807f
C2378 _449_/a_2665_112# _176_ 0.048319f
C2379 FILLER_0_21_28/a_2364_375# _012_ 0.017669f
C2380 comp net3 0.05248f
C2381 net1 net18 0.047886f
C2382 FILLER_0_5_72/a_36_472# vss 0.031034f
C2383 FILLER_0_5_72/a_484_472# vdd 0.002735f
C2384 _031_ FILLER_0_2_111/a_932_472# 0.017509f
C2385 _270_/a_36_472# net76 0.009569f
C2386 en_co_clk _038_ 0.014475f
C2387 en_co_clk _120_ 0.008507f
C2388 _050_ FILLER_0_22_128/a_1468_375# 0.001661f
C2389 _098_ FILLER_0_19_171/a_36_472# 0.021559f
C2390 net81 FILLER_0_15_235/a_572_375# 0.009675f
C2391 FILLER_0_5_54/a_572_375# trim_mask\[1\] 0.011664f
C2392 output46/a_224_472# vss 0.00432f
C2393 FILLER_0_16_89/a_572_375# net14 0.00106f
C2394 FILLER_0_4_144/a_36_472# _081_ 0.003547f
C2395 _255_/a_224_552# _090_ 0.001598f
C2396 FILLER_0_21_125/a_124_375# _022_ 0.007023f
C2397 output45/a_224_472# net40 0.001284f
C2398 FILLER_0_20_87/a_124_375# vss 0.00279f
C2399 FILLER_0_20_87/a_36_472# vdd 0.006784f
C2400 FILLER_0_15_142/a_36_472# fanout73/a_36_113# 0.009544f
C2401 _127_ net53 0.00917f
C2402 FILLER_0_7_72/a_1828_472# net50 0.094122f
C2403 fanout52/a_36_160# _170_ 0.024724f
C2404 net58 FILLER_0_9_270/a_572_375# 0.006256f
C2405 _451_/a_1353_112# vdd 0.009693f
C2406 _153_ _157_ 0.050552f
C2407 _308_/a_1084_68# trim_mask\[0\] 0.001592f
C2408 FILLER_0_21_286/a_36_472# _009_ 0.003266f
C2409 net81 vdd 1.658963f
C2410 _446_/a_1204_472# net40 0.026414f
C2411 _070_ FILLER_0_10_94/a_124_375# 0.008294f
C2412 _426_/a_36_151# FILLER_0_8_247/a_36_472# 0.001723f
C2413 _304_/a_224_472# _111_ 0.003461f
C2414 vss _166_ 0.011302f
C2415 vdd _160_ 0.606139f
C2416 _431_/a_36_151# fanout70/a_36_113# 0.016241f
C2417 _375_/a_36_68# vss 0.02182f
C2418 net20 mask\[2\] 0.050364f
C2419 FILLER_0_12_2/a_124_375# _450_/a_36_151# 0.001543f
C2420 net57 _085_ 0.211414f
C2421 net41 FILLER_0_23_44/a_124_375# 0.001526f
C2422 _131_ FILLER_0_9_105/a_572_375# 0.031928f
C2423 FILLER_0_2_93/a_484_472# FILLER_0_2_101/a_36_472# 0.013277f
C2424 output9/a_224_472# FILLER_0_1_266/a_484_472# 0.0323f
C2425 FILLER_0_9_28/a_932_472# net16 0.017841f
C2426 _185_ _278_/a_36_160# 0.001237f
C2427 net31 _099_ 0.01086f
C2428 _165_ FILLER_0_6_37/a_124_375# 0.002884f
C2429 FILLER_0_11_124/a_36_472# vss 0.002545f
C2430 _267_/a_1792_472# _055_ 0.003058f
C2431 _016_ _327_/a_36_472# 0.04536f
C2432 _091_ FILLER_0_15_212/a_484_472# 0.049391f
C2433 net34 _199_/a_36_160# 0.026709f
C2434 output34/a_224_472# output32/a_224_472# 0.001691f
C2435 output36/a_224_472# FILLER_0_14_263/a_36_472# 0.001711f
C2436 _223_/a_36_160# vdd 0.018653f
C2437 _185_ vss 0.021437f
C2438 fanout82/a_36_113# net19 0.021188f
C2439 _178_ _185_ 0.979797f
C2440 net66 FILLER_0_3_54/a_36_472# 0.008174f
C2441 _414_/a_2560_156# net22 0.00603f
C2442 _372_/a_2590_472# _062_ 0.0012f
C2443 FILLER_0_14_91/a_36_472# _095_ 0.014431f
C2444 _350_/a_665_69# net23 0.001468f
C2445 ctln[1] net1 0.003756f
C2446 output11/a_224_472# ctln[4] 0.072677f
C2447 _128_ FILLER_0_9_142/a_124_375# 0.004439f
C2448 net31 _419_/a_2248_156# 0.001521f
C2449 FILLER_0_18_107/a_484_472# net14 0.002472f
C2450 net62 _100_ 0.006742f
C2451 output34/a_224_472# _277_/a_36_160# 0.014508f
C2452 _219_/a_36_160# trim_mask\[0\] 0.395762f
C2453 _372_/a_786_69# _163_ 0.001179f
C2454 _414_/a_796_472# _081_ 0.003538f
C2455 FILLER_0_18_37/a_124_375# vdd 0.024546f
C2456 _432_/a_1204_472# net80 0.009362f
C2457 FILLER_0_0_130/a_124_375# _442_/a_36_151# 0.059049f
C2458 result[0] net18 0.085445f
C2459 _447_/a_36_151# net17 0.001448f
C2460 FILLER_0_16_107/a_572_375# net70 0.002193f
C2461 _431_/a_36_151# net53 0.001579f
C2462 output8/a_224_472# _078_ 0.001267f
C2463 _069_ state\[1\] 0.003884f
C2464 _431_/a_448_472# _132_ 0.003024f
C2465 _413_/a_448_472# net59 0.059041f
C2466 _239_/a_36_160# vdd 0.042369f
C2467 FILLER_0_7_72/a_932_472# net50 0.074005f
C2468 net20 _420_/a_2248_156# 0.003737f
C2469 net79 _138_ 0.024731f
C2470 fanout55/a_36_160# _067_ 0.126784f
C2471 vdd net30 0.636147f
C2472 _131_ _125_ 0.013932f
C2473 _177_ _176_ 0.226424f
C2474 net66 _164_ 0.093385f
C2475 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_36_472# 0.086635f
C2476 _059_ _313_/a_67_603# 0.061666f
C2477 FILLER_0_10_37/a_36_472# net16 0.012905f
C2478 FILLER_0_16_37/a_36_472# net72 0.005134f
C2479 _098_ _433_/a_2560_156# 0.004273f
C2480 fanout53/a_36_160# vss 0.006674f
C2481 _428_/a_2665_112# vss 0.005991f
C2482 FILLER_0_20_193/a_484_472# net21 0.00371f
C2483 _077_ FILLER_0_10_78/a_1020_375# 0.001131f
C2484 output47/a_224_472# vdd 0.028666f
C2485 _437_/a_2248_156# net14 0.023718f
C2486 FILLER_0_4_144/a_484_472# _443_/a_36_151# 0.002841f
C2487 _072_ _248_/a_36_68# 0.001683f
C2488 fanout75/a_36_113# net76 0.040306f
C2489 _074_ net1 0.128466f
C2490 _395_/a_36_488# _121_ 0.009689f
C2491 FILLER_0_9_28/a_3260_375# vss 0.05542f
C2492 _408_/a_718_524# FILLER_0_12_28/a_124_375# 0.001192f
C2493 FILLER_0_13_80/a_124_375# vdd 0.018971f
C2494 _422_/a_2665_112# _009_ 0.061508f
C2495 ctln[7] _442_/a_2665_112# 0.01075f
C2496 vss cal_count\[0\] 0.160743f
C2497 _178_ _407_/a_36_472# 0.001699f
C2498 _178_ cal_count\[0\] 0.011488f
C2499 _098_ FILLER_0_15_235/a_36_472# 0.093007f
C2500 FILLER_0_20_177/a_932_472# _098_ 0.008366f
C2501 FILLER_0_17_64/a_124_375# FILLER_0_15_59/a_484_472# 0.001188f
C2502 net27 FILLER_0_10_247/a_36_472# 0.016681f
C2503 net57 _062_ 0.067654f
C2504 FILLER_0_7_72/a_1380_472# _077_ 0.001315f
C2505 net55 _452_/a_3129_107# 0.006395f
C2506 _444_/a_36_151# net17 0.001435f
C2507 _068_ _311_/a_1920_473# 0.001498f
C2508 net60 _420_/a_2665_112# 0.038894f
C2509 net41 vdd 1.983262f
C2510 FILLER_0_18_177/a_2364_375# net21 0.018463f
C2511 ctln[1] _411_/a_36_151# 0.018351f
C2512 _098_ vss 0.958032f
C2513 net15 FILLER_0_5_54/a_1020_375# 0.015944f
C2514 FILLER_0_3_54/a_124_375# _164_ 0.008654f
C2515 _334_/a_36_160# FILLER_0_17_104/a_1380_472# 0.004111f
C2516 net54 _436_/a_2560_156# 0.010748f
C2517 FILLER_0_21_286/a_484_472# FILLER_0_23_290/a_124_375# 0.001404f
C2518 trim_mask\[1\] FILLER_0_6_47/a_2724_472# 0.003645f
C2519 _424_/a_1308_423# _012_ 0.007041f
C2520 net62 FILLER_0_14_235/a_124_375# 0.015659f
C2521 mask\[5\] FILLER_0_20_177/a_124_375# 0.013531f
C2522 _033_ _444_/a_1308_423# 0.002877f
C2523 net44 FILLER_0_8_2/a_124_375# 0.083677f
C2524 FILLER_0_18_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001684f
C2525 FILLER_0_8_2/a_36_472# vss 0.004429f
C2526 _118_ _315_/a_36_68# 0.005792f
C2527 _205_/a_36_160# vss 0.003612f
C2528 ctln[3] output10/a_224_472# 0.064347f
C2529 output9/a_224_472# net2 0.003405f
C2530 _057_ calibrate 0.002047f
C2531 _417_/a_36_151# vdd 0.140703f
C2532 FILLER_0_19_47/a_572_375# vss 0.055293f
C2533 FILLER_0_19_47/a_36_472# vdd 0.072773f
C2534 net18 _416_/a_1000_472# 0.046085f
C2535 _101_ _005_ 0.003946f
C2536 _421_/a_36_151# _419_/a_2248_156# 0.001203f
C2537 _374_/a_36_68# vdd 0.075685f
C2538 net35 FILLER_0_22_86/a_572_375# 0.010986f
C2539 mask\[8\] FILLER_0_22_86/a_1020_375# 0.009431f
C2540 net44 FILLER_0_15_10/a_36_472# 0.012286f
C2541 fanout49/a_36_160# vss 0.025717f
C2542 _057_ net21 0.143214f
C2543 FILLER_0_7_59/a_572_375# vdd 0.005991f
C2544 FILLER_0_7_59/a_124_375# vss 0.002006f
C2545 _277_/a_36_160# _099_ 0.001628f
C2546 FILLER_0_13_212/a_572_375# _043_ 0.01418f
C2547 state\[0\] _273_/a_36_68# 0.012187f
C2548 FILLER_0_9_28/a_2276_472# _042_ 0.002496f
C2549 FILLER_0_22_128/a_3260_375# _146_ 0.004692f
C2550 net75 _001_ 0.056236f
C2551 _255_/a_224_552# _163_ 0.002169f
C2552 net35 FILLER_0_22_128/a_1380_472# 0.016004f
C2553 net79 _113_ 0.002432f
C2554 fanout64/a_36_160# vss 0.007097f
C2555 net33 _146_ 0.306187f
C2556 _069_ FILLER_0_13_212/a_124_375# 0.070185f
C2557 _414_/a_36_151# _057_ 0.003902f
C2558 net59 FILLER_0_3_212/a_36_472# 0.058623f
C2559 _387_/a_36_113# vss 0.047621f
C2560 _131_ cal_count\[2\] 0.044147f
C2561 net20 ctln[4] 0.00225f
C2562 net68 FILLER_0_6_47/a_36_472# 0.001248f
C2563 _415_/a_2248_156# fanout62/a_36_160# 0.007753f
C2564 _185_ _184_ 0.047803f
C2565 net17 FILLER_0_23_44/a_572_375# 0.001332f
C2566 net31 output18/a_224_472# 0.04975f
C2567 fanout49/a_36_160# _441_/a_2248_156# 0.027388f
C2568 result[4] net19 0.015095f
C2569 FILLER_0_4_49/a_124_375# _167_ 0.009437f
C2570 net60 _419_/a_2560_156# 0.006989f
C2571 net20 FILLER_0_12_220/a_1468_375# 0.016974f
C2572 net54 FILLER_0_22_128/a_1916_375# 0.001933f
C2573 _444_/a_1204_472# net40 0.017496f
C2574 _070_ FILLER_0_9_105/a_484_472# 0.020248f
C2575 _091_ net57 0.006076f
C2576 FILLER_0_5_128/a_484_472# _370_/a_124_24# 0.00171f
C2577 _414_/a_2248_156# _074_ 0.013023f
C2578 _077_ _439_/a_1308_423# 0.022235f
C2579 net81 _283_/a_36_472# 0.032292f
C2580 _013_ FILLER_0_17_56/a_36_472# 0.002659f
C2581 mask\[5\] _295_/a_36_472# 0.034027f
C2582 _440_/a_2248_156# trim_mask\[1\] 0.004408f
C2583 _133_ vdd 0.27652f
C2584 _070_ vss 1.363355f
C2585 net32 _102_ 0.038622f
C2586 _217_/a_36_160# _424_/a_36_151# 0.035111f
C2587 _432_/a_36_151# vss 0.003647f
C2588 FILLER_0_17_72/a_1828_472# _438_/a_36_151# 0.001221f
C2589 cal_itt\[2\] _253_/a_36_68# 0.010756f
C2590 _406_/a_36_159# net47 0.034933f
C2591 _429_/a_2665_112# FILLER_0_14_235/a_124_375# 0.006271f
C2592 FILLER_0_15_180/a_572_375# vdd 0.068901f
C2593 _073_ _084_ 0.048469f
C2594 FILLER_0_7_146/a_36_472# vss 0.029149f
C2595 net50 trim_val\[3\] 0.111824f
C2596 FILLER_0_9_223/a_572_375# _426_/a_2665_112# 0.005202f
C2597 _411_/a_2665_112# net75 0.005223f
C2598 _119_ _077_ 2.584241f
C2599 result[7] FILLER_0_24_290/a_36_472# 0.005185f
C2600 FILLER_0_4_185/a_124_375# _002_ 0.013895f
C2601 net75 _014_ 0.204357f
C2602 net1 _081_ 0.111227f
C2603 _321_/a_170_472# _395_/a_36_488# 0.007047f
C2604 FILLER_0_21_28/a_572_375# net40 0.001406f
C2605 _163_ FILLER_0_6_79/a_36_472# 0.001789f
C2606 ctln[0] vdd 0.051631f
C2607 trim_mask\[2\] FILLER_0_3_78/a_572_375# 0.011713f
C2608 _075_ _070_ 0.009314f
C2609 _321_/a_2034_472# _120_ 0.002489f
C2610 _300_/a_224_472# _009_ 0.001405f
C2611 _096_ _320_/a_1568_472# 0.001632f
C2612 _317_/a_36_113# vdd 0.054289f
C2613 _063_ trim_val\[0\] 0.001978f
C2614 FILLER_0_14_50/a_36_472# vdd 0.081414f
C2615 FILLER_0_14_50/a_124_375# vss 0.002412f
C2616 net34 _435_/a_448_472# 0.013341f
C2617 _064_ net40 0.141744f
C2618 _308_/a_124_24# _070_ 0.001465f
C2619 _326_/a_36_160# _077_ 0.00419f
C2620 FILLER_0_6_239/a_36_472# _074_ 0.004715f
C2621 net77 _007_ 0.002591f
C2622 net68 _440_/a_36_151# 0.080854f
C2623 _176_ _451_/a_2225_156# 0.030788f
C2624 FILLER_0_17_72/a_3172_472# _131_ 0.003717f
C2625 net67 FILLER_0_6_47/a_36_472# 0.004607f
C2626 _420_/a_2248_156# _009_ 0.00681f
C2627 _086_ _267_/a_224_472# 0.004041f
C2628 net1 net65 0.035488f
C2629 _061_ cal_count\[3\] 0.003415f
C2630 net81 _069_ 0.034401f
C2631 net76 net18 0.002264f
C2632 net68 FILLER_0_8_37/a_484_472# 0.002696f
C2633 _076_ _125_ 0.009254f
C2634 net55 vss 0.947665f
C2635 FILLER_0_7_72/a_1380_472# net50 0.077411f
C2636 ctlp[4] net32 0.001413f
C2637 fanout49/a_36_160# FILLER_0_5_88/a_124_375# 0.001154f
C2638 _155_ FILLER_0_4_107/a_124_375# 0.00162f
C2639 _188_ _453_/a_36_151# 0.03354f
C2640 output25/a_224_472# net24 0.002325f
C2641 _407_/a_36_472# _184_ 0.004667f
C2642 _093_ _136_ 0.226819f
C2643 _095_ _451_/a_448_472# 0.002474f
C2644 net42 net40 0.007686f
C2645 net27 output27/a_224_472# 0.046353f
C2646 FILLER_0_17_200/a_36_472# _430_/a_36_151# 0.001723f
C2647 _005_ _094_ 0.162984f
C2648 _074_ _251_/a_906_472# 0.002887f
C2649 net73 FILLER_0_17_142/a_36_472# 0.002925f
C2650 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_572_375# 0.007947f
C2651 _063_ _445_/a_2248_156# 0.008121f
C2652 net17 _054_ 0.034759f
C2653 ctlp[2] _299_/a_36_472# 0.012937f
C2654 _131_ _043_ 0.047425f
C2655 FILLER_0_17_72/a_932_472# net36 0.00356f
C2656 FILLER_0_7_104/a_1380_472# _154_ 0.002799f
C2657 _359_/a_36_488# net74 0.037211f
C2658 _137_ _334_/a_36_160# 0.015722f
C2659 _093_ _438_/a_1000_472# 0.001556f
C2660 _442_/a_3041_156# vdd 0.001178f
C2661 mask\[9\] _438_/a_796_472# 0.004751f
C2662 _030_ _154_ 0.004803f
C2663 FILLER_0_5_164/a_572_375# vss 0.055055f
C2664 FILLER_0_5_164/a_36_472# vdd 0.004144f
C2665 _126_ FILLER_0_11_124/a_124_375# 0.038971f
C2666 _376_/a_36_160# trim_mask\[1\] 0.003111f
C2667 FILLER_0_18_171/a_36_472# vdd 0.010704f
C2668 net50 trim_val\[0\] 0.390586f
C2669 net58 vss 0.589419f
C2670 net52 _442_/a_36_151# 0.029373f
C2671 FILLER_0_18_177/a_3260_375# vss 0.055219f
C2672 FILLER_0_18_177/a_36_472# vdd 0.110153f
C2673 net72 _174_ 0.199504f
C2674 net20 FILLER_0_3_221/a_1020_375# 0.025371f
C2675 net66 FILLER_0_5_54/a_572_375# 0.002203f
C2676 _339_/a_36_160# FILLER_0_19_155/a_572_375# 0.003589f
C2677 _450_/a_3129_107# _039_ 0.012762f
C2678 FILLER_0_11_101/a_484_472# cal_count\[3\] 0.00702f
C2679 net18 _419_/a_1308_423# 0.013637f
C2680 _095_ _185_ 0.034457f
C2681 net69 _168_ 0.035976f
C2682 _439_/a_36_151# FILLER_0_6_47/a_2364_375# 0.002807f
C2683 output27/a_224_472# _425_/a_2665_112# 0.021504f
C2684 mask\[4\] FILLER_0_18_209/a_36_472# 0.018888f
C2685 net16 FILLER_0_18_37/a_484_472# 0.054878f
C2686 net17 vss 0.940703f
C2687 net69 _441_/a_796_472# 0.002057f
C2688 FILLER_0_17_104/a_124_375# net14 0.010099f
C2689 _178_ net17 0.115251f
C2690 _429_/a_36_151# _043_ 0.002771f
C2691 _072_ cal_count\[3\] 0.028346f
C2692 trim_val\[1\] vss 0.029927f
C2693 _114_ FILLER_0_10_107/a_124_375# 0.004825f
C2694 _140_ _436_/a_36_151# 0.031519f
C2695 FILLER_0_21_125/a_572_375# _144_ 0.003787f
C2696 _425_/a_1308_423# vdd 0.021703f
C2697 FILLER_0_17_282/a_36_472# _418_/a_448_472# 0.011962f
C2698 net17 FILLER_0_20_15/a_932_472# 0.047256f
C2699 net73 FILLER_0_18_107/a_1828_472# 0.01544f
C2700 net37 FILLER_0_6_231/a_124_375# 0.001989f
C2701 mask\[7\] FILLER_0_22_128/a_36_472# 0.013408f
C2702 FILLER_0_17_282/a_124_375# _006_ 0.004694f
C2703 FILLER_0_15_142/a_36_472# net36 0.015456f
C2704 net4 _060_ 0.327437f
C2705 ctln[5] net22 0.072969f
C2706 net64 FILLER_0_9_270/a_124_375# 0.013532f
C2707 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1468_375# 0.086635f
C2708 state\[2\] _427_/a_448_472# 0.00237f
C2709 net53 _427_/a_796_472# 0.001983f
C2710 _414_/a_2248_156# _081_ 0.002027f
C2711 output35/a_224_472# vss 0.01667f
C2712 _002_ FILLER_0_3_172/a_1828_472# 0.016749f
C2713 _067_ FILLER_0_12_20/a_124_375# 0.017026f
C2714 _082_ vss 0.053349f
C2715 result[0] net65 0.011634f
C2716 net82 vss 0.550252f
C2717 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_572_375# 0.086635f
C2718 FILLER_0_18_76/a_572_375# _438_/a_36_151# 0.059049f
C2719 cal_itt\[2\] FILLER_0_3_221/a_484_472# 0.016997f
C2720 _428_/a_448_472# net74 0.019814f
C2721 net61 ctlp[1] 2.770871f
C2722 FILLER_0_16_107/a_484_472# FILLER_0_14_107/a_572_375# 0.001404f
C2723 _445_/a_2560_156# net49 0.001208f
C2724 net50 _439_/a_1308_423# 0.008832f
C2725 net52 _439_/a_1000_472# 0.03537f
C2726 net3 FILLER_0_15_10/a_124_375# 0.035504f
C2727 output24/a_224_472# net24 0.005559f
C2728 FILLER_0_4_49/a_124_375# vdd 0.008637f
C2729 _126_ _428_/a_2248_156# 0.001131f
C2730 _115_ _127_ 0.042389f
C2731 _411_/a_36_151# net65 0.001415f
C2732 FILLER_0_9_223/a_36_472# _246_/a_36_68# 0.006596f
C2733 _098_ FILLER_0_16_154/a_1020_375# 0.003386f
C2734 net81 net28 0.034606f
C2735 fanout57/a_36_113# vss 0.046378f
C2736 fanout54/a_36_160# FILLER_0_19_142/a_124_375# 0.005489f
C2737 output38/a_224_472# net40 0.072234f
C2738 cal_itt\[2\] _079_ 0.017071f
C2739 _013_ FILLER_0_18_53/a_36_472# 0.013138f
C2740 _428_/a_2665_112# _095_ 0.001471f
C2741 ctlp[7] net25 0.003141f
C2742 fanout53/a_36_160# _095_ 0.007436f
C2743 _238_/a_67_603# vss 0.008203f
C2744 _043_ FILLER_0_13_80/a_36_472# 0.016194f
C2745 _136_ _337_/a_49_472# 0.058704f
C2746 _091_ FILLER_0_13_212/a_932_472# 0.008749f
C2747 FILLER_0_5_54/a_124_375# FILLER_0_3_54/a_36_472# 0.001512f
C2748 _015_ FILLER_0_8_247/a_36_472# 0.005458f
C2749 FILLER_0_3_78/a_484_472# vss 0.005811f
C2750 _176_ FILLER_0_10_107/a_124_375# 0.013408f
C2751 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_36_472# 0.086743f
C2752 FILLER_0_12_124/a_36_472# net74 0.021369f
C2753 FILLER_0_22_86/a_124_375# vss 0.00285f
C2754 FILLER_0_22_86/a_572_375# vdd 0.017472f
C2755 FILLER_0_11_78/a_124_375# _120_ 0.014367f
C2756 net68 fanout68/a_36_113# 0.027807f
C2757 net58 fanout76/a_36_160# 0.055026f
C2758 FILLER_0_22_128/a_1380_472# vdd 0.005746f
C2759 FILLER_0_22_128/a_932_472# vss 0.003452f
C2760 _058_ trim_mask\[0\] 0.076069f
C2761 net35 _146_ 0.096468f
C2762 _216_/a_67_603# vss 0.012211f
C2763 FILLER_0_4_197/a_932_472# _088_ 0.014643f
C2764 net81 FILLER_0_12_236/a_572_375# 0.021025f
C2765 _095_ cal_count\[0\] 0.005211f
C2766 result[8] _422_/a_36_151# 0.001488f
C2767 _074_ net76 0.026801f
C2768 ctln[8] FILLER_0_0_96/a_124_375# 0.002726f
C2769 FILLER_0_9_223/a_572_375# _223_/a_36_160# 0.001177f
C2770 _116_ net4 0.00603f
C2771 _056_ _226_/a_1044_68# 0.002852f
C2772 FILLER_0_8_138/a_36_472# _070_ 0.001342f
C2773 net45 net40 0.029947f
C2774 _412_/a_36_151# net48 0.001091f
C2775 _121_ vdd 0.106437f
C2776 net56 FILLER_0_18_139/a_1468_375# 0.065206f
C2777 net75 FILLER_0_8_263/a_36_472# 0.020293f
C2778 fanout78/a_36_113# vdd 0.061637f
C2779 _088_ FILLER_0_3_172/a_3172_472# 0.004381f
C2780 _425_/a_1000_472# net19 0.020388f
C2781 _111_ vss 0.233815f
C2782 _065_ net50 0.123581f
C2783 _445_/a_36_151# _034_ 0.005488f
C2784 net64 FILLER_0_11_282/a_36_472# 0.003938f
C2785 net76 _076_ 0.003124f
C2786 _185_ _402_/a_1296_93# 0.001714f
C2787 ctln[4] output12/a_224_472# 0.041517f
C2788 net82 FILLER_0_3_172/a_3260_375# 0.007693f
C2789 _070_ _071_ 0.001757f
C2790 FILLER_0_14_50/a_124_375# _401_/a_36_68# 0.001129f
C2791 FILLER_0_5_54/a_124_375# _164_ 0.004076f
C2792 _095_ _098_ 0.057687f
C2793 net57 net14 0.05113f
C2794 trim_mask\[2\] _447_/a_36_151# 0.022881f
C2795 FILLER_0_3_172/a_2364_375# net65 0.003745f
C2796 cal_itt\[2\] cal_itt\[1\] 0.057194f
C2797 mask\[5\] FILLER_0_21_206/a_124_375# 0.011644f
C2798 _256_/a_1612_497# net4 0.002497f
C2799 _128_ _085_ 0.004532f
C2800 net57 fanout55/a_36_160# 0.017476f
C2801 _077_ _161_ 0.023053f
C2802 FILLER_0_8_127/a_36_472# net74 0.063481f
C2803 _046_ vdd 0.041841f
C2804 net48 _112_ 0.284235f
C2805 result[7] FILLER_0_23_282/a_484_472# 0.013947f
C2806 net82 fanout76/a_36_160# 0.001033f
C2807 result[9] _108_ 0.015443f
C2808 _316_/a_848_380# _123_ 0.0018f
C2809 FILLER_0_17_200/a_484_472# _093_ 0.007492f
C2810 FILLER_0_15_116/a_36_472# vdd 0.013454f
C2811 _443_/a_36_151# vdd 0.175472f
C2812 _274_/a_36_68# net27 0.027359f
C2813 result[9] net19 0.540761f
C2814 ctln[5] vdd 0.256793f
C2815 FILLER_0_12_136/a_1020_375# net23 0.005919f
C2816 net20 FILLER_0_13_212/a_1020_375# 0.003962f
C2817 _077_ _129_ 0.08682f
C2818 _409_/a_245_68# cal_count\[3\] 0.001164f
C2819 _132_ FILLER_0_19_111/a_484_472# 0.004619f
C2820 _448_/a_796_472# vdd 0.002153f
C2821 _439_/a_2248_156# net14 0.001279f
C2822 net27 FILLER_0_14_235/a_484_472# 0.010072f
C2823 output14/a_224_472# ctln[7] 0.076006f
C2824 net22 net59 0.195226f
C2825 net68 _220_/a_67_603# 0.030878f
C2826 _149_ FILLER_0_20_98/a_124_375# 0.020028f
C2827 FILLER_0_13_228/a_124_375# FILLER_0_12_220/a_1020_375# 0.05841f
C2828 net20 _421_/a_1204_472# 0.019627f
C2829 FILLER_0_16_57/a_124_375# net72 0.052543f
C2830 net15 FILLER_0_17_56/a_572_375# 0.007386f
C2831 FILLER_0_7_59/a_36_472# net68 0.050931f
C2832 FILLER_0_5_54/a_1020_375# net47 0.005159f
C2833 net26 FILLER_0_21_28/a_2276_472# 0.001561f
C2834 net57 _428_/a_36_151# 0.023215f
C2835 _184_ net17 0.007958f
C2836 _433_/a_2248_156# _145_ 0.009108f
C2837 _073_ _260_/a_36_68# 0.079772f
C2838 FILLER_0_16_89/a_124_375# _136_ 0.011795f
C2839 _376_/a_36_160# FILLER_0_6_90/a_36_472# 0.195478f
C2840 FILLER_0_8_107/a_36_472# _155_ 0.002068f
C2841 _043_ FILLER_0_15_180/a_36_472# 0.001219f
C2842 _104_ ctlp[2] 1.420577f
C2843 _431_/a_1000_472# _020_ 0.009685f
C2844 mask\[3\] _102_ 0.142836f
C2845 FILLER_0_17_72/a_2364_375# vdd 0.002455f
C2846 FILLER_0_17_72/a_1916_375# vss 0.001345f
C2847 FILLER_0_12_20/a_572_375# net47 0.00139f
C2848 net55 _027_ 0.002104f
C2849 ctlp[2] vss 0.131085f
C2850 _091_ _141_ 0.010074f
C2851 _142_ net23 0.037306f
C2852 result[7] result[6] 0.119475f
C2853 net7 trim[3] 0.044017f
C2854 FILLER_0_4_107/a_36_472# vss 0.002634f
C2855 FILLER_0_2_111/a_932_472# _158_ 0.00264f
C2856 FILLER_0_4_107/a_484_472# vdd 0.03151f
C2857 _028_ FILLER_0_6_47/a_3172_472# 0.015585f
C2858 output8/a_224_472# _080_ 0.001971f
C2859 FILLER_0_18_2/a_3260_375# _452_/a_36_151# 0.001597f
C2860 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001597f
C2861 _073_ net4 0.076114f
C2862 _091_ net36 0.067629f
C2863 FILLER_0_9_28/a_3172_472# net51 0.047897f
C2864 result[6] FILLER_0_21_286/a_124_375# 0.019179f
C2865 FILLER_0_16_107/a_124_375# _040_ 0.008721f
C2866 _427_/a_36_151# vdd 0.107344f
C2867 net72 FILLER_0_15_59/a_124_375# 0.022905f
C2868 _346_/a_49_472# _098_ 0.028579f
C2869 _119_ cal_itt\[3\] 0.010152f
C2870 _122_ net22 0.024638f
C2871 _043_ FILLER_0_13_72/a_124_375# 0.013517f
C2872 _091_ _429_/a_1204_472# 0.024554f
C2873 net31 net18 0.114197f
C2874 _424_/a_2248_156# FILLER_0_21_60/a_572_375# 0.030666f
C2875 _424_/a_2665_112# FILLER_0_21_60/a_124_375# 0.010688f
C2876 FILLER_0_12_220/a_124_375# _070_ 0.007554f
C2877 trim_val\[2\] _167_ 0.011787f
C2878 trim_mask\[2\] FILLER_0_2_93/a_124_375# 0.046032f
C2879 net63 FILLER_0_18_177/a_36_472# 0.015187f
C2880 net76 _081_ 0.706096f
C2881 net60 _421_/a_2248_156# 0.036944f
C2882 _321_/a_170_472# vdd 0.060585f
C2883 en_co_clk _043_ 0.041355f
C2884 FILLER_0_14_50/a_124_375# _095_ 0.052375f
C2885 _115_ trim_mask\[0\] 0.008966f
C2886 _179_ _180_ 0.018662f
C2887 FILLER_0_16_89/a_1380_472# _131_ 0.004201f
C2888 _018_ net21 0.077174f
C2889 net79 _044_ 0.013636f
C2890 FILLER_0_11_142/a_36_472# _120_ 0.040786f
C2891 _408_/a_1336_472# vss 0.001022f
C2892 _408_/a_728_93# vdd 0.024163f
C2893 net41 FILLER_0_21_28/a_932_472# 0.014034f
C2894 FILLER_0_13_142/a_932_472# vss 0.005192f
C2895 FILLER_0_13_142/a_1380_472# vdd 0.001977f
C2896 net49 _440_/a_796_472# 0.003597f
C2897 _128_ _062_ 0.025708f
C2898 mask\[7\] _299_/a_36_472# 0.033949f
C2899 net50 FILLER_0_5_72/a_1380_472# 0.002431f
C2900 FILLER_0_7_59/a_36_472# net67 0.021549f
C2901 net38 FILLER_0_15_2/a_572_375# 0.007477f
C2902 _235_/a_255_603# trim_mask\[2\] 0.001488f
C2903 _235_/a_67_603# trim_val\[2\] 0.00747f
C2904 net55 _095_ 0.055644f
C2905 _415_/a_2665_112# fanout62/a_36_160# 0.016426f
C2906 FILLER_0_11_142/a_484_472# FILLER_0_13_142/a_572_375# 0.0027f
C2907 net76 net65 0.14935f
C2908 _062_ _311_/a_692_473# 0.008632f
C2909 _447_/a_796_472# vdd 0.001959f
C2910 net57 FILLER_0_8_156/a_124_375# 0.001628f
C2911 net24 FILLER_0_22_107/a_124_375# 0.001023f
C2912 net15 FILLER_0_9_72/a_36_472# 0.006905f
C2913 _356_/a_36_472# vdd 0.016338f
C2914 result[2] net18 0.086474f
C2915 FILLER_0_11_64/a_124_375# _453_/a_36_151# 0.005577f
C2916 net23 FILLER_0_22_128/a_1468_375# 0.001866f
C2917 net54 _352_/a_49_472# 0.003941f
C2918 net59 vdd 2.180407f
C2919 _137_ FILLER_0_16_154/a_1468_375# 0.014214f
C2920 net23 _207_/a_67_603# 0.002734f
C2921 _189_/a_67_603# net62 0.001695f
C2922 _315_/a_716_497# net23 0.004725f
C2923 fanout72/a_36_113# _067_ 0.005796f
C2924 net54 _433_/a_1000_472# 0.0025f
C2925 FILLER_0_0_198/a_124_375# vdd 0.04491f
C2926 output37/a_224_472# fanout64/a_36_160# 0.017421f
C2927 _450_/a_2449_156# net40 0.010265f
C2928 net15 _453_/a_2248_156# 0.044493f
C2929 _008_ _419_/a_36_151# 0.014476f
C2930 FILLER_0_17_200/a_36_472# mask\[3\] 0.27914f
C2931 _214_/a_36_160# _213_/a_67_603# 0.002505f
C2932 _077_ _056_ 1.777574f
C2933 FILLER_0_16_89/a_124_375# net53 0.001032f
C2934 _095_ net17 0.172789f
C2935 net20 _429_/a_448_472# 0.002244f
C2936 _444_/a_1308_423# _054_ 0.005457f
C2937 vdd FILLER_0_10_94/a_484_472# 0.008627f
C2938 _077_ FILLER_0_7_59/a_484_472# 0.001371f
C2939 net73 FILLER_0_17_104/a_1468_375# 0.002342f
C2940 trim[4] net39 0.004535f
C2941 _077_ _453_/a_36_151# 0.042928f
C2942 FILLER_0_20_107/a_124_375# FILLER_0_20_98/a_124_375# 0.003228f
C2943 _146_ vdd 0.031209f
C2944 _105_ _420_/a_2665_112# 0.001159f
C2945 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_124_375# 0.001597f
C2946 result[9] _419_/a_448_472# 0.015767f
C2947 FILLER_0_18_2/a_2724_472# net40 0.011079f
C2948 _413_/a_448_472# ctln[4] 0.001072f
C2949 net82 FILLER_0_2_177/a_36_472# 0.001777f
C2950 trimb[1] net40 0.00126f
C2951 fanout59/a_36_160# net5 0.05829f
C2952 FILLER_0_8_24/a_572_375# _054_ 0.004858f
C2953 _261_/a_36_160# FILLER_0_5_136/a_36_472# 0.00304f
C2954 _431_/a_36_151# _020_ 0.023081f
C2955 cal_count\[1\] FILLER_0_15_59/a_572_375# 0.008797f
C2956 _415_/a_36_151# vdd 0.115639f
C2957 FILLER_0_21_142/a_124_375# _433_/a_448_472# 0.006782f
C2958 FILLER_0_0_130/a_124_375# _031_ 0.001861f
C2959 net65 FILLER_0_2_177/a_124_375# 0.018094f
C2960 _036_ net17 0.153479f
C2961 _058_ _118_ 0.001451f
C2962 _449_/a_1000_472# net72 0.001247f
C2963 _449_/a_448_472# net55 0.004439f
C2964 output26/a_224_472# net17 0.004277f
C2965 _025_ _436_/a_1000_472# 0.061189f
C2966 _021_ _093_ 0.049589f
C2967 _070_ _385_/a_36_68# 0.049178f
C2968 _091_ _128_ 0.003717f
C2969 _132_ net73 0.460325f
C2970 _422_/a_36_151# _109_ 0.036674f
C2971 _096_ _225_/a_36_160# 0.004807f
C2972 FILLER_0_5_206/a_124_375# net22 0.019537f
C2973 calibrate vss 1.140031f
C2974 _122_ vdd 0.379907f
C2975 net80 FILLER_0_19_171/a_36_472# 0.040915f
C2976 trimb[3] FILLER_0_20_2/a_484_472# 0.001829f
C2977 _110_ net36 0.002287f
C2978 fanout54/a_36_160# vss 0.061573f
C2979 net64 FILLER_0_15_235/a_572_375# 0.007219f
C2980 FILLER_0_16_37/a_124_375# vss 0.021237f
C2981 FILLER_0_16_37/a_36_472# vdd 0.142203f
C2982 _178_ FILLER_0_16_37/a_124_375# 0.036901f
C2983 FILLER_0_7_233/a_124_375# vdd 0.03915f
C2984 _308_/a_124_24# FILLER_0_10_94/a_36_472# 0.001811f
C2985 _044_ FILLER_0_13_290/a_124_375# 0.001855f
C2986 ctln[7] vdd 0.359832f
C2987 _411_/a_36_151# FILLER_0_0_232/a_124_375# 0.059049f
C2988 FILLER_0_10_256/a_124_375# vss 0.006036f
C2989 FILLER_0_10_256/a_36_472# vdd 0.025204f
C2990 FILLER_0_2_111/a_36_472# trim_mask\[3\] 0.007915f
C2991 _421_/a_36_151# net18 0.00659f
C2992 FILLER_0_8_24/a_572_375# vss 0.012859f
C2993 FILLER_0_8_24/a_36_472# vdd 0.007423f
C2994 _077_ _068_ 0.601166f
C2995 _035_ net47 0.101683f
C2996 _227_/a_36_160# vdd 0.007828f
C2997 state\[0\] _323_/a_36_113# 0.016796f
C2998 net64 vdd 1.155692f
C2999 _453_/a_2248_156# net51 0.05329f
C3000 _120_ _172_ 0.010275f
C3001 _038_ _172_ 0.050158f
C3002 net21 vss 1.123312f
C3003 net35 FILLER_0_23_88/a_124_375# 0.009071f
C3004 fanout51/a_36_113# FILLER_0_11_64/a_124_375# 0.002335f
C3005 net62 _045_ 0.029263f
C3006 FILLER_0_7_72/a_1468_375# _164_ 0.003223f
C3007 output32/a_224_472# net18 0.022521f
C3008 _333_/a_36_160# vss 0.030799f
C3009 FILLER_0_4_144/a_124_375# trim_mask\[4\] 0.014395f
C3010 _169_ vdd 0.055642f
C3011 _075_ calibrate 0.022901f
C3012 net38 _452_/a_448_472# 0.016895f
C3013 _189_/a_67_603# _429_/a_2665_112# 0.015187f
C3014 FILLER_0_4_49/a_572_375# net68 0.023227f
C3015 net20 result[4] 0.001673f
C3016 net70 FILLER_0_18_107/a_1380_472# 0.00116f
C3017 FILLER_0_2_93/a_484_472# vdd 0.005163f
C3018 _414_/a_36_151# vss 0.002101f
C3019 _072_ _267_/a_224_472# 0.004269f
C3020 _438_/a_1308_423# net14 0.005201f
C3021 FILLER_0_0_96/a_124_375# net14 0.077876f
C3022 FILLER_0_4_144/a_124_375# net47 0.012023f
C3023 FILLER_0_19_171/a_932_472# vss 0.001256f
C3024 FILLER_0_19_171/a_1380_472# vdd 0.03086f
C3025 output8/a_224_472# vss 0.076244f
C3026 _063_ _232_/a_67_603# 0.005404f
C3027 FILLER_0_14_91/a_124_375# en_co_clk 0.006788f
C3028 _069_ _121_ 0.137961f
C3029 net23 FILLER_0_5_148/a_36_472# 0.011079f
C3030 FILLER_0_7_72/a_3260_375# net14 0.025344f
C3031 FILLER_0_15_72/a_572_375# _451_/a_3129_107# 0.007026f
C3032 _075_ net21 0.012335f
C3033 output10/a_224_472# FILLER_0_0_266/a_124_375# 0.00515f
C3034 net44 _452_/a_2225_156# 0.044858f
C3035 _412_/a_2560_156# en 0.049213f
C3036 _402_/a_728_93# _182_ 0.00263f
C3037 trim_val\[2\] vdd 0.160419f
C3038 trim_mask\[2\] vss 0.182675f
C3039 net47 FILLER_0_5_148/a_484_472# 0.009741f
C3040 net17 output41/a_224_472# 0.030456f
C3041 FILLER_0_22_86/a_1020_375# _026_ 0.001032f
C3042 _253_/a_36_68# _084_ 0.029805f
C3043 FILLER_0_2_165/a_124_375# net59 0.00999f
C3044 _230_/a_652_68# _062_ 0.001144f
C3045 _410_/a_36_68# vss 0.02717f
C3046 _086_ _132_ 0.014693f
C3047 FILLER_0_23_44/a_36_472# vdd 0.01833f
C3048 FILLER_0_23_44/a_1468_375# vss 0.055902f
C3049 net15 _441_/a_1308_423# 0.009697f
C3050 _173_ FILLER_0_12_28/a_124_375# 0.009218f
C3051 _002_ _087_ 0.00636f
C3052 net58 output37/a_224_472# 0.099539f
C3053 _408_/a_1336_472# _184_ 0.003286f
C3054 _018_ mask\[1\] 0.001206f
C3055 _440_/a_2665_112# net47 0.014066f
C3056 FILLER_0_4_197/a_484_472# _088_ 0.014756f
C3057 _418_/a_448_472# vss 0.005772f
C3058 _418_/a_1308_423# vdd 0.002258f
C3059 _006_ vdd 0.632993f
C3060 FILLER_0_14_107/a_1380_472# vdd 0.002511f
C3061 _112_ net37 0.070289f
C3062 ctln[2] output10/a_224_472# 0.024524f
C3063 FILLER_0_3_172/a_3260_375# net21 0.049606f
C3064 _431_/a_2248_156# _137_ 0.01617f
C3065 clk vss 0.210484f
C3066 _056_ FILLER_0_12_196/a_36_472# 0.039555f
C3067 FILLER_0_22_177/a_36_472# net33 0.013661f
C3068 _433_/a_796_472# _022_ 0.025882f
C3069 cal_itt\[3\] _161_ 0.20195f
C3070 fanout65/a_36_113# net65 0.019148f
C3071 net52 FILLER_0_9_72/a_124_375# 0.029702f
C3072 _043_ _090_ 0.001578f
C3073 FILLER_0_21_286/a_572_375# vss 0.031895f
C3074 FILLER_0_21_286/a_36_472# vdd 0.008714f
C3075 FILLER_0_16_255/a_36_472# net30 0.00209f
C3076 FILLER_0_15_116/a_572_375# _095_ 0.00152f
C3077 _103_ vdd 0.590261f
C3078 net36 net14 0.037175f
C3079 FILLER_0_3_204/a_124_375# FILLER_0_4_197/a_932_472# 0.001597f
C3080 FILLER_0_21_28/a_1380_472# net17 0.001709f
C3081 FILLER_0_1_266/a_124_375# vdd -0.002281f
C3082 FILLER_0_4_177/a_484_472# _087_ 0.005486f
C3083 FILLER_0_9_223/a_484_472# vss 0.006102f
C3084 _114_ _085_ 0.056448f
C3085 _075_ _414_/a_448_472# 0.020304f
C3086 FILLER_0_5_206/a_124_375# vdd 0.038311f
C3087 net2 net4 0.854661f
C3088 net50 FILLER_0_7_59/a_484_472# 0.011974f
C3089 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_36_472# 0.026657f
C3090 _104_ mask\[7\] 0.069172f
C3091 FILLER_0_18_61/a_124_375# vss 0.021307f
C3092 FILLER_0_18_61/a_36_472# vdd 0.08828f
C3093 _428_/a_1204_472# _131_ 0.012968f
C3094 fanout66/a_36_113# net49 0.001044f
C3095 mask\[7\] vss 0.85153f
C3096 _115_ _118_ 1.045555f
C3097 _411_/a_448_472# vss 0.009447f
C3098 net26 FILLER_0_18_37/a_572_375# 0.00109f
C3099 FILLER_0_12_124/a_124_375# _127_ 0.003767f
C3100 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_124_375# 0.001597f
C3101 vdd FILLER_0_4_91/a_572_375# 0.019853f
C3102 _074_ FILLER_0_6_231/a_36_472# 0.004325f
C3103 _098_ FILLER_0_20_87/a_124_375# 0.019333f
C3104 FILLER_0_15_142/a_124_375# _136_ 0.001706f
C3105 cal_count\[3\] FILLER_0_11_78/a_484_472# 0.011737f
C3106 ctlp[1] FILLER_0_24_274/a_1468_375# 0.01305f
C3107 FILLER_0_3_172/a_932_472# net22 0.012284f
C3108 _427_/a_448_472# _043_ 0.002896f
C3109 _422_/a_1000_472# mask\[7\] 0.039617f
C3110 FILLER_0_5_109/a_572_375# FILLER_0_5_117/a_124_375# 0.012001f
C3111 result[6] _420_/a_1000_472# 0.007761f
C3112 _341_/a_49_472# net23 0.031763f
C3113 net80 vss 0.347557f
C3114 FILLER_0_18_177/a_1468_375# _139_ 0.001359f
C3115 _076_ FILLER_0_6_231/a_36_472# 0.005517f
C3116 _407_/a_36_472# _185_ 0.009281f
C3117 _085_ _176_ 0.024708f
C3118 _185_ cal_count\[0\] 0.008096f
C3119 trim[4] clkc 0.005f
C3120 output30/a_224_472# net30 0.043557f
C3121 output31/a_224_472# net60 0.216716f
C3122 FILLER_0_18_107/a_2812_375# FILLER_0_17_133/a_36_472# 0.001543f
C3123 net74 _136_ 0.042043f
C3124 net27 _426_/a_36_151# 0.008613f
C3125 _053_ FILLER_0_6_47/a_3260_375# 0.002746f
C3126 _093_ FILLER_0_17_72/a_2276_472# 0.017114f
C3127 net16 _408_/a_1936_472# 0.022235f
C3128 _321_/a_170_472# _069_ 0.025551f
C3129 _408_/a_56_524# _043_ 0.10151f
C3130 _436_/a_2665_112# FILLER_0_22_128/a_1020_375# 0.029834f
C3131 FILLER_0_15_235/a_36_472# mask\[1\] 0.009316f
C3132 net74 FILLER_0_13_142/a_124_375# 0.002722f
C3133 FILLER_0_5_198/a_572_375# net59 0.00183f
C3134 FILLER_0_8_138/a_36_472# calibrate 0.047835f
C3135 _431_/a_36_151# FILLER_0_18_107/a_2276_472# 0.002799f
C3136 FILLER_0_1_266/a_36_472# net19 0.07227f
C3137 FILLER_0_5_54/a_36_472# FILLER_0_6_47/a_932_472# 0.026657f
C3138 FILLER_0_5_54/a_1020_375# FILLER_0_6_47/a_1828_472# 0.001597f
C3139 mask\[7\] _107_ 0.13732f
C3140 _428_/a_448_472# net70 0.007116f
C3141 mask\[2\] net22 0.034216f
C3142 _412_/a_2665_112# cal_itt\[1\] 0.015571f
C3143 net68 _029_ 0.094915f
C3144 _369_/a_244_472# vdd 0.001255f
C3145 FILLER_0_16_57/a_36_472# FILLER_0_17_56/a_124_375# 0.001723f
C3146 mask\[1\] vss 0.46268f
C3147 _192_/a_255_603# mask\[1\] 0.001059f
C3148 FILLER_0_10_78/a_36_472# vss 0.008832f
C3149 net36 FILLER_0_15_212/a_932_472# 0.008239f
C3150 _408_/a_1336_472# _095_ 0.011305f
C3151 _104_ _422_/a_2248_156# 0.041703f
C3152 _095_ FILLER_0_13_142/a_932_472# 0.001782f
C3153 FILLER_0_2_177/a_572_375# net59 0.005397f
C3154 FILLER_0_11_142/a_572_375# vdd 0.014107f
C3155 FILLER_0_11_142/a_124_375# vss 0.008766f
C3156 _188_ _042_ 0.015684f
C3157 _079_ _084_ 0.046584f
C3158 _322_/a_848_380# _129_ 0.048486f
C3159 _092_ FILLER_0_17_218/a_36_472# 0.033277f
C3160 FILLER_0_18_107/a_2364_375# vdd 0.017472f
C3161 _434_/a_36_151# mask\[6\] 0.048644f
C3162 net24 FILLER_0_22_86/a_1468_375# 0.008075f
C3163 _422_/a_2248_156# vss 0.001755f
C3164 _422_/a_2665_112# vdd 0.008306f
C3165 trim_mask\[4\] _386_/a_124_24# 0.040347f
C3166 FILLER_0_7_104/a_572_375# vdd 0.038253f
C3167 FILLER_0_7_72/a_36_472# _439_/a_36_151# 0.013806f
C3168 FILLER_0_18_139/a_1468_375# _145_ 0.002318f
C3169 net79 FILLER_0_12_220/a_484_472# 0.005464f
C3170 _441_/a_2560_156# vss 0.001374f
C3171 net47 _386_/a_124_24# 0.024696f
C3172 _029_ _156_ 0.018258f
C3173 fanout70/a_36_113# net74 0.002663f
C3174 _074_ _375_/a_1388_497# 0.005488f
C3175 _114_ _062_ 0.028432f
C3176 net55 _424_/a_2560_156# 0.003707f
C3177 mask\[4\] FILLER_0_18_177/a_1916_375# 0.013466f
C3178 net48 net1 0.006424f
C3179 fanout78/a_36_113# net77 0.036366f
C3180 output23/a_224_472# _049_ 0.001034f
C3181 _174_ vdd 0.18623f
C3182 mask\[0\] _018_ 0.328328f
C3183 mask\[3\] FILLER_0_16_241/a_124_375# 0.006824f
C3184 mask\[3\] FILLER_0_18_177/a_1020_375# 0.002924f
C3185 _447_/a_1000_472# net68 0.006223f
C3186 _447_/a_1308_423# _036_ 0.003079f
C3187 net50 net69 0.634381f
C3188 net52 _031_ 0.633473f
C3189 FILLER_0_23_88/a_124_375# vdd 0.03583f
C3190 _432_/a_1000_472# _137_ 0.008914f
C3191 _033_ FILLER_0_6_47/a_36_472# 0.001185f
C3192 _325_/a_224_472# _130_ 0.001685f
C3193 result[5] net61 0.092275f
C3194 net24 _211_/a_36_160# 0.021941f
C3195 input2/a_36_113# vss 0.055539f
C3196 _122_ FILLER_0_5_198/a_572_375# 0.001352f
C3197 FILLER_0_5_109/a_36_472# _153_ 0.034328f
C3198 _431_/a_1456_156# net73 0.001304f
C3199 net47 _452_/a_1353_112# 0.003681f
C3200 _417_/a_36_151# output30/a_224_472# 0.004902f
C3201 _126_ FILLER_0_10_94/a_572_375# 0.027249f
C3202 _091_ _274_/a_36_68# 0.025773f
C3203 _208_/a_36_160# FILLER_0_22_128/a_3260_375# 0.001948f
C3204 net63 net64 0.002181f
C3205 _131_ FILLER_0_17_104/a_932_472# 0.002988f
C3206 _062_ _226_/a_276_68# 0.001286f
C3207 _441_/a_448_472# net66 0.023761f
C3208 ctlp[5] _024_ 0.022549f
C3209 FILLER_0_18_2/a_3172_472# vdd 0.011201f
C3210 _093_ FILLER_0_18_139/a_572_375# 0.008393f
C3211 _097_ vdd 0.191424f
C3212 _053_ FILLER_0_8_37/a_36_472# 0.001011f
C3213 _324_/a_224_472# net74 0.001704f
C3214 _437_/a_448_472# vss 0.001524f
C3215 _437_/a_1308_423# vdd 0.005139f
C3216 trim[4] net47 0.009333f
C3217 FILLER_0_19_125/a_36_472# FILLER_0_18_107/a_1916_375# 0.001684f
C3218 FILLER_0_15_142/a_124_375# net53 0.033224f
C3219 cal_itt\[3\] _056_ 0.023192f
C3220 _449_/a_1204_472# _038_ 0.005899f
C3221 FILLER_0_18_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001684f
C3222 FILLER_0_3_172/a_932_472# vdd 0.009887f
C3223 _062_ FILLER_0_5_136/a_36_472# 0.001404f
C3224 FILLER_0_5_54/a_932_472# _440_/a_36_151# 0.001723f
C3225 FILLER_0_5_198/a_36_472# net21 0.014911f
C3226 _325_/a_224_472# _129_ 0.003137f
C3227 net63 FILLER_0_19_171/a_1380_472# 0.003014f
C3228 FILLER_0_21_125/a_36_472# _433_/a_36_151# 0.001723f
C3229 net38 cal_count\[3\] 0.002225f
C3230 output13/a_224_472# vss 0.108144f
C3231 FILLER_0_7_104/a_36_472# _058_ 0.006613f
C3232 FILLER_0_14_107/a_1020_375# FILLER_0_16_115/a_36_472# 0.001512f
C3233 net16 _444_/a_2560_156# 0.010829f
C3234 _413_/a_36_151# FILLER_0_3_204/a_36_472# 0.001723f
C3235 cal_itt\[1\] _084_ 0.495918f
C3236 FILLER_0_18_2/a_2724_472# _452_/a_1040_527# 0.001138f
C3237 output34/a_224_472# _104_ 0.112239f
C3238 FILLER_0_10_28/a_36_472# net6 0.038613f
C3239 _069_ _122_ 0.002164f
C3240 net19 _044_ 0.138869f
C3241 _414_/a_796_472# _003_ 0.006511f
C3242 trim_val\[4\] net22 0.144267f
C3243 output20/a_224_472# net61 0.177946f
C3244 net20 result[9] 1.593573f
C3245 output47/a_224_472# FILLER_0_15_10/a_36_472# 0.038484f
C3246 ctlp[0] vdd 0.08832f
C3247 _102_ _094_ 0.727442f
C3248 FILLER_0_18_76/a_484_472# net71 0.004649f
C3249 net53 net74 0.164124f
C3250 FILLER_0_16_107/a_572_375# net14 0.002308f
C3251 output34/a_224_472# vss 0.011966f
C3252 _053_ _160_ 0.0539f
C3253 mask\[2\] FILLER_0_15_235/a_572_375# 0.003879f
C3254 _412_/a_1204_472# net65 0.001629f
C3255 FILLER_0_5_181/a_124_375# vss 0.011456f
C3256 FILLER_0_5_181/a_36_472# vdd 0.081434f
C3257 _155_ _156_ 0.037229f
C3258 vss output6/a_224_472# 0.004205f
C3259 FILLER_0_24_63/a_124_375# vdd 0.029514f
C3260 FILLER_0_9_223/a_36_472# net4 0.014911f
C3261 FILLER_0_22_177/a_484_472# mask\[6\] 0.006573f
C3262 FILLER_0_22_177/a_124_375# _146_ 0.001864f
C3263 net35 FILLER_0_22_177/a_36_472# 0.005721f
C3264 _093_ FILLER_0_18_76/a_36_472# 0.129892f
C3265 mask\[2\] vdd 0.433058f
C3266 _098_ _205_/a_36_160# 0.033853f
C3267 mask\[9\] FILLER_0_18_76/a_572_375# 0.006158f
C3268 _195_/a_67_603# mask\[1\] 0.016836f
C3269 _028_ _058_ 0.041158f
C3270 net15 ctln[9] 0.01475f
C3271 net70 FILLER_0_17_104/a_1020_375# 0.001894f
C3272 net76 FILLER_0_5_206/a_36_472# 0.00169f
C3273 _171_ vss 0.004501f
C3274 net34 FILLER_0_22_128/a_1468_375# 0.003214f
C3275 _020_ _093_ 0.015474f
C3276 FILLER_0_13_206/a_36_472# net79 0.00402f
C3277 net54 _149_ 0.212511f
C3278 net34 _207_/a_67_603# 0.008585f
C3279 net75 FILLER_0_8_247/a_484_472# 0.003007f
C3280 output46/a_224_472# net17 0.082914f
C3281 _104_ _298_/a_224_472# 0.001731f
C3282 net54 FILLER_0_18_139/a_572_375# 0.00217f
C3283 output48/a_224_472# vss 0.006655f
C3284 cal_count\[3\] _067_ 0.478427f
C3285 _360_/a_36_160# FILLER_0_4_123/a_124_375# 0.013555f
C3286 _004_ FILLER_0_10_247/a_36_472# 0.001551f
C3287 result[7] _419_/a_1204_472# 0.018181f
C3288 _008_ net60 0.314106f
C3289 _413_/a_2665_112# vss 0.012213f
C3290 FILLER_0_8_247/a_124_375# vss 0.002674f
C3291 FILLER_0_8_247/a_572_375# vdd -0.007963f
C3292 net46 FILLER_0_21_28/a_124_375# 0.011995f
C3293 _430_/a_1308_423# mask\[2\] 0.020226f
C3294 FILLER_0_18_171/a_124_375# mask\[3\] 0.001156f
C3295 _085_ _267_/a_36_472# 0.034055f
C3296 net81 _425_/a_36_151# 0.014663f
C3297 mask\[0\] vss 0.694674f
C3298 trim_val\[1\] _166_ 0.06773f
C3299 _399_/a_224_472# net72 0.002538f
C3300 _015_ FILLER_0_10_247/a_124_375# 0.001261f
C3301 _300_/a_224_472# vdd 0.001344f
C3302 FILLER_0_13_100/a_36_472# vss 0.003094f
C3303 _187_ cal_count\[3\] 0.031898f
C3304 _093_ FILLER_0_18_209/a_572_375# 0.064723f
C3305 FILLER_0_9_28/a_2812_375# _077_ 0.006629f
C3306 _432_/a_448_472# _091_ 0.050539f
C3307 FILLER_0_5_206/a_124_375# FILLER_0_5_198/a_572_375# 0.012001f
C3308 _415_/a_36_151# net28 0.001195f
C3309 _441_/a_36_151# _164_ 0.008955f
C3310 trim_mask\[2\] _036_ 0.466145f
C3311 FILLER_0_16_73/a_572_375# _176_ 0.006454f
C3312 _179_ vss 0.089947f
C3313 _163_ _156_ 0.001616f
C3314 net3 _278_/a_36_160# 0.014154f
C3315 _178_ _179_ 0.063494f
C3316 _046_ _282_/a_36_160# 0.005584f
C3317 mask\[3\] _198_/a_67_603# 0.024102f
C3318 FILLER_0_20_107/a_36_472# net71 0.004375f
C3319 _185_ net17 0.270086f
C3320 _095_ FILLER_0_14_107/a_932_472# 0.014431f
C3321 _420_/a_2248_156# vdd 0.00331f
C3322 output17/a_224_472# ctlp[0] 0.018696f
C3323 FILLER_0_15_205/a_124_375# net22 0.049201f
C3324 net4 FILLER_0_12_220/a_932_472# 0.050731f
C3325 net3 vss 0.02666f
C3326 net24 net71 0.015101f
C3327 _432_/a_36_151# _098_ 0.00957f
C3328 vdd FILLER_0_16_115/a_124_375# 0.020393f
C3329 _032_ vdd 0.174834f
C3330 _178_ net3 0.257606f
C3331 FILLER_0_10_256/a_36_472# net28 0.00136f
C3332 _098_ FILLER_0_15_180/a_124_375# 0.019007f
C3333 _142_ _141_ 0.200324f
C3334 _242_/a_36_160# vss 0.032884f
C3335 _444_/a_1000_472# net67 0.025169f
C3336 ctlp[3] ctlp[4] 0.027598f
C3337 _113_ FILLER_0_12_196/a_36_472# 0.002495f
C3338 _136_ _019_ 0.049263f
C3339 net52 _443_/a_1000_472# 0.016322f
C3340 _308_/a_848_380# _114_ 0.005266f
C3341 FILLER_0_17_200/a_36_472# _432_/a_2665_112# 0.007491f
C3342 _446_/a_2665_112# net49 0.006979f
C3343 trim_val\[4\] vdd 0.245329f
C3344 net44 _450_/a_836_156# 0.006278f
C3345 FILLER_0_16_57/a_124_375# vdd 0.008567f
C3346 net67 FILLER_0_8_24/a_484_472# 0.001065f
C3347 vdd _450_/a_3129_107# 0.039939f
C3348 net35 _436_/a_1308_423# 0.008773f
C3349 FILLER_0_3_78/a_36_472# _160_ 0.006564f
C3350 _330_/a_224_472# _134_ 0.007508f
C3351 _174_ _401_/a_244_472# 0.001957f
C3352 net48 _251_/a_906_472# 0.001362f
C3353 _322_/a_848_380# _068_ 0.009682f
C3354 _063_ FILLER_0_6_37/a_124_375# 0.012149f
C3355 net52 _448_/a_2665_112# 0.039348f
C3356 output37/a_224_472# calibrate 0.013149f
C3357 FILLER_0_15_212/a_124_375# vss 0.005813f
C3358 FILLER_0_15_212/a_572_375# vdd -0.014642f
C3359 _099_ vss 0.255039f
C3360 output11/a_224_472# FILLER_0_0_232/a_36_472# 0.023414f
C3361 net57 _017_ 0.045694f
C3362 net15 FILLER_0_18_76/a_36_472# 0.001341f
C3363 _131_ _180_ 0.016104f
C3364 FILLER_0_18_2/a_932_472# net55 0.012117f
C3365 calibrate _385_/a_36_68# 0.001996f
C3366 FILLER_0_20_177/a_36_472# _434_/a_36_151# 0.001723f
C3367 FILLER_0_20_177/a_1468_375# _434_/a_448_472# 0.008952f
C3368 FILLER_0_4_99/a_36_472# vss 0.002273f
C3369 FILLER_0_16_154/a_36_472# vss 0.005098f
C3370 FILLER_0_16_154/a_484_472# vdd 0.001006f
C3371 FILLER_0_13_65/a_124_375# vss 0.030194f
C3372 _104_ _294_/a_224_472# 0.003008f
C3373 _430_/a_2665_112# mask\[2\] 0.028551f
C3374 net64 FILLER_0_12_236/a_572_375# 0.005704f
C3375 _144_ _352_/a_49_472# 0.00176f
C3376 _411_/a_2248_156# net75 0.032114f
C3377 trim_mask\[1\] FILLER_0_6_47/a_572_375# 0.007164f
C3378 FILLER_0_19_111/a_572_375# vdd -0.008314f
C3379 _236_/a_36_160# net40 0.035082f
C3380 _421_/a_1000_472# _010_ 0.01379f
C3381 FILLER_0_22_86/a_1380_472# net14 0.039176f
C3382 _294_/a_224_472# vss 0.001022f
C3383 _414_/a_2560_156# _053_ 0.008732f
C3384 _415_/a_1000_472# vdd 0.002497f
C3385 _419_/a_2665_112# vdd 0.030085f
C3386 _144_ _433_/a_1000_472# 0.029564f
C3387 _074_ _078_ 0.003088f
C3388 FILLER_0_15_59/a_124_375# vdd 0.017243f
C3389 output25/a_224_472# net35 0.016177f
C3390 FILLER_0_18_2/a_3260_375# _041_ 0.001024f
C3391 _143_ _340_/a_36_160# 0.001064f
C3392 _057_ net56 0.002158f
C3393 FILLER_0_19_47/a_572_375# net55 0.003447f
C3394 _116_ FILLER_0_12_196/a_124_375# 0.005332f
C3395 FILLER_0_12_136/a_484_472# _127_ 0.005549f
C3396 net19 _420_/a_2560_156# 0.010978f
C3397 FILLER_0_16_89/a_484_472# _093_ 0.001526f
C3398 _132_ _433_/a_36_151# 0.024768f
C3399 _076_ _078_ 0.012626f
C3400 net50 FILLER_0_6_37/a_124_375# 0.003821f
C3401 net54 FILLER_0_20_107/a_124_375# 0.072539f
C3402 mask\[7\] FILLER_0_22_177/a_572_375# 0.001315f
C3403 FILLER_0_15_116/a_36_472# _451_/a_36_151# 0.096503f
C3404 FILLER_0_19_195/a_124_375# _202_/a_36_160# 0.005489f
C3405 output36/a_224_472# net30 0.083671f
C3406 net76 FILLER_0_3_172/a_1380_472# 0.015215f
C3407 _053_ FILLER_0_7_59/a_572_375# 0.014569f
C3408 _000_ _080_ 0.002867f
C3409 FILLER_0_7_146/a_124_375# _133_ 0.001577f
C3410 net52 trim_mask\[1\] 0.04149f
C3411 net72 _453_/a_36_151# 0.001607f
C3412 FILLER_0_17_200/a_572_375# vss 0.017327f
C3413 _079_ _260_/a_36_68# 0.043596f
C3414 _093_ FILLER_0_17_142/a_484_472# 0.011974f
C3415 _064_ _445_/a_36_151# 0.03209f
C3416 FILLER_0_13_212/a_36_472# net79 0.006158f
C3417 cal_count\[3\] net23 0.045417f
C3418 FILLER_0_18_177/a_3260_375# _205_/a_36_160# 0.001313f
C3419 result[9] _009_ 0.19745f
C3420 net62 FILLER_0_13_212/a_484_472# 0.059367f
C3421 _069_ FILLER_0_11_142/a_572_375# 0.020472f
C3422 _095_ mask\[1\] 0.001297f
C3423 net49 trim_mask\[1\] 0.003402f
C3424 output39/a_224_472# net67 0.008957f
C3425 mask\[5\] FILLER_0_18_177/a_572_375# 0.002653f
C3426 FILLER_0_18_107/a_3172_472# _145_ 0.002415f
C3427 net4 FILLER_0_3_221/a_484_472# 0.043027f
C3428 _059_ net23 0.265909f
C3429 net80 FILLER_0_22_177/a_572_375# 0.005202f
C3430 mask\[7\] _435_/a_2560_156# 0.011544f
C3431 net69 FILLER_0_2_101/a_36_472# 0.00845f
C3432 FILLER_0_15_205/a_124_375# vdd 0.015886f
C3433 ctln[4] vdd 0.210384f
C3434 FILLER_0_1_212/a_36_472# vss 0.00858f
C3435 _450_/a_1040_527# output6/a_224_472# 0.005581f
C3436 _450_/a_448_472# net6 0.041113f
C3437 net52 _157_ 0.005889f
C3438 trim_val\[3\] vdd 0.211478f
C3439 _079_ net4 0.023763f
C3440 output35/a_224_472# _098_ 0.003653f
C3441 _181_ cal_count\[1\] 0.186904f
C3442 FILLER_0_10_78/a_1020_375# vdd 0.002901f
C3443 FILLER_0_12_220/a_1020_375# vss 0.004698f
C3444 FILLER_0_12_220/a_1468_375# vdd 0.002801f
C3445 _411_/a_36_151# net10 0.127193f
C3446 _053_ _133_ 0.288819f
C3447 net58 fanout64/a_36_160# 0.002438f
C3448 FILLER_0_12_136/a_1380_472# _076_ 0.001809f
C3449 net1 net37 0.00519f
C3450 _426_/a_2248_156# calibrate 0.004597f
C3451 cal_count\[3\] FILLER_0_11_109/a_124_375# 0.004618f
C3452 output35/a_224_472# _205_/a_36_160# 0.002043f
C3453 FILLER_0_18_139/a_1380_472# vss 0.009272f
C3454 net74 _058_ 0.026905f
C3455 FILLER_0_9_72/a_1468_375# _439_/a_2248_156# 0.001901f
C3456 trim_val\[4\] FILLER_0_2_165/a_124_375# 0.009193f
C3457 output39/a_224_472# _445_/a_448_472# 0.009352f
C3458 _093_ FILLER_0_18_107/a_2276_472# 0.001996f
C3459 FILLER_0_5_72/a_1020_375# _029_ 0.010208f
C3460 FILLER_0_5_117/a_124_375# _153_ 0.079379f
C3461 FILLER_0_22_177/a_1468_375# vss 0.028064f
C3462 FILLER_0_22_177/a_36_472# vdd 0.111906f
C3463 _016_ _131_ 0.017461f
C3464 net48 net76 0.069349f
C3465 _099_ _195_/a_67_603# 0.065049f
C3466 _114_ net14 0.127764f
C3467 FILLER_0_7_195/a_36_472# _072_ 0.008357f
C3468 _390_/a_36_68# _038_ 0.019355f
C3469 _143_ _141_ 0.192528f
C3470 net81 FILLER_0_9_270/a_36_472# 0.084422f
C3471 mask\[2\] FILLER_0_16_154/a_572_375# 0.026605f
C3472 net63 mask\[2\] 0.553545f
C3473 _401_/a_36_68# _179_ 0.007074f
C3474 FILLER_0_4_107/a_1468_375# _160_ 0.028099f
C3475 _443_/a_2665_112# _066_ 0.001654f
C3476 _412_/a_2248_156# cal_itt\[1\] 0.005868f
C3477 FILLER_0_4_213/a_124_375# vss 0.006145f
C3478 FILLER_0_4_213/a_572_375# vdd 0.026692f
C3479 net25 _213_/a_67_603# 0.027452f
C3480 net18 FILLER_0_17_282/a_36_472# 0.036965f
C3481 _070_ FILLER_0_5_164/a_572_375# 0.001083f
C3482 _024_ _023_ 0.005966f
C3483 FILLER_0_22_86/a_124_375# _098_ 0.011864f
C3484 _140_ _146_ 0.135012f
C3485 _418_/a_36_151# _007_ 0.007397f
C3486 _077_ _042_ 0.045685f
C3487 FILLER_0_17_72/a_1020_375# _131_ 0.005847f
C3488 fanout62/a_36_160# net79 0.011515f
C3489 _061_ _247_/a_36_160# 0.009993f
C3490 _136_ _451_/a_2225_156# 0.01289f
C3491 _065_ _235_/a_67_603# 0.004135f
C3492 _367_/a_36_68# vdd 0.010246f
C3493 net27 _015_ 0.103416f
C3494 _449_/a_796_472# vss 0.00143f
C3495 net32 _108_ 0.035815f
C3496 FILLER_0_21_286/a_36_472# net77 0.001557f
C3497 result[6] _421_/a_796_472# 0.004697f
C3498 net70 FILLER_0_14_123/a_36_472# 0.009456f
C3499 _103_ net77 0.004691f
C3500 net73 FILLER_0_17_133/a_124_375# 0.022541f
C3501 net32 net19 0.65591f
C3502 net4 cal_itt\[1\] 0.048147f
C3503 _057_ _074_ 0.013823f
C3504 FILLER_0_9_142/a_124_375# _315_/a_36_68# 0.028077f
C3505 _096_ _306_/a_36_68# 0.016266f
C3506 _026_ _437_/a_796_472# 0.008884f
C3507 _149_ _437_/a_1204_472# 0.024276f
C3508 _111_ _098_ 0.014998f
C3509 cal_count\[2\] _183_ 0.034303f
C3510 fanout49/a_36_160# FILLER_0_3_78/a_484_472# 0.003699f
C3511 _078_ _081_ 0.445443f
C3512 trim_val\[0\] vdd 0.056059f
C3513 _451_/a_1353_112# _040_ 0.005265f
C3514 state\[0\] _072_ 0.030642f
C3515 FILLER_0_5_109/a_124_375# FILLER_0_4_107/a_484_472# 0.001684f
C3516 _104_ output18/a_224_472# 0.08426f
C3517 _122_ FILLER_0_6_231/a_484_472# 0.017477f
C3518 _123_ FILLER_0_6_231/a_124_375# 0.001259f
C3519 _114_ _428_/a_36_151# 0.008132f
C3520 result[4] FILLER_0_17_282/a_124_375# 0.018106f
C3521 _176_ net14 0.031922f
C3522 _069_ mask\[2\] 0.032781f
C3523 FILLER_0_14_263/a_36_472# net30 0.003972f
C3524 net7 _446_/a_2248_156# 0.001166f
C3525 _057_ _076_ 0.041986f
C3526 FILLER_0_16_73/a_36_472# FILLER_0_17_72/a_124_375# 0.001723f
C3527 FILLER_0_7_72/a_1468_375# _376_/a_36_160# 0.02985f
C3528 net64 _282_/a_36_160# 0.014431f
C3529 output38/a_224_472# _445_/a_36_151# 0.199812f
C3530 FILLER_0_7_233/a_124_375# FILLER_0_6_231/a_484_472# 0.001684f
C3531 ctln[3] FILLER_0_0_266/a_124_375# 0.002726f
C3532 net41 _446_/a_448_472# 0.040165f
C3533 sample result[0] 0.081581f
C3534 _176_ fanout55/a_36_160# 0.070942f
C3535 output18/a_224_472# vss 0.086897f
C3536 net60 _109_ 0.021502f
C3537 _449_/a_36_151# _174_ 0.002252f
C3538 _196_/a_36_160# FILLER_0_14_263/a_124_375# 0.005732f
C3539 net16 _164_ 0.015161f
C3540 _425_/a_36_151# _317_/a_36_113# 0.002361f
C3541 _137_ FILLER_0_15_180/a_572_375# 0.028083f
C3542 _072_ _247_/a_36_160# 0.005008f
C3543 net18 FILLER_0_9_270/a_572_375# 0.005977f
C3544 _445_/a_2248_156# vdd 0.018573f
C3545 _091_ _092_ 0.028594f
C3546 _372_/a_2590_472# _059_ 0.002974f
C3547 FILLER_0_21_28/a_2724_472# vdd 0.001342f
C3548 net55 net17 0.056153f
C3549 _436_/a_1308_423# vdd 0.005258f
C3550 trimb[1] FILLER_0_19_28/a_36_472# 0.01233f
C3551 FILLER_0_3_221/a_572_375# vss 0.003292f
C3552 _423_/a_1204_472# _012_ 0.003181f
C3553 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_572_375# 0.007947f
C3554 net36 _438_/a_796_472# 0.016855f
C3555 _000_ vss 0.205593f
C3556 ctln[3] ctln[2] 0.012289f
C3557 net16 _404_/a_36_472# 0.001126f
C3558 _428_/a_2248_156# _427_/a_36_151# 0.035837f
C3559 FILLER_0_5_117/a_36_472# _360_/a_36_160# 0.003913f
C3560 _439_/a_448_472# vss 0.036535f
C3561 _439_/a_1308_423# vdd 0.002368f
C3562 _114_ FILLER_0_11_109/a_36_472# 0.023029f
C3563 _126_ FILLER_0_13_100/a_124_375# 0.00134f
C3564 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_124_375# 0.012222f
C3565 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1468_375# 0.001597f
C3566 FILLER_0_8_239/a_36_472# _123_ 0.011767f
C3567 mask\[0\] _095_ 0.006711f
C3568 FILLER_0_21_28/a_2812_375# _424_/a_36_151# 0.059049f
C3569 _427_/a_2665_112# net23 0.032729f
C3570 _095_ FILLER_0_13_100/a_36_472# 0.003036f
C3571 mask\[4\] net22 0.075713f
C3572 _132_ FILLER_0_19_125/a_124_375# 0.009167f
C3573 net63 FILLER_0_15_212/a_572_375# 0.001597f
C3574 net70 _136_ 0.032219f
C3575 _050_ _025_ 0.033887f
C3576 _119_ vdd 0.38257f
C3577 fanout62/a_36_160# FILLER_0_13_290/a_124_375# 0.001138f
C3578 mask\[7\] _147_ 0.295801f
C3579 trim[0] trim[1] 0.001567f
C3580 FILLER_0_10_37/a_124_375# FILLER_0_10_28/a_124_375# 0.003228f
C3581 FILLER_0_7_162/a_36_472# net57 0.015199f
C3582 FILLER_0_12_136/a_572_375# cal_count\[3\] 0.005006f
C3583 ctlp[1] fanout77/a_36_113# 0.012793f
C3584 _190_/a_36_160# net47 0.001489f
C3585 ctln[2] net5 0.001249f
C3586 net58 _425_/a_448_472# 0.002474f
C3587 net50 FILLER_0_6_90/a_124_375# 0.041764f
C3588 FILLER_0_12_2/a_124_375# vdd 0.0247f
C3589 FILLER_0_0_266/a_36_472# vss 0.003738f
C3590 _115_ net74 0.033145f
C3591 _375_/a_36_68# calibrate 0.048799f
C3592 FILLER_0_10_214/a_36_472# net22 0.001634f
C3593 output25/a_224_472# vdd 0.03413f
C3594 _112_ _425_/a_1204_472# 0.001132f
C3595 FILLER_0_6_239/a_36_472# net37 0.004187f
C3596 net56 FILLER_0_19_142/a_124_375# 0.003154f
C3597 FILLER_0_16_57/a_484_472# _176_ 0.013507f
C3598 FILLER_0_9_28/a_2364_375# _220_/a_67_603# 0.002082f
C3599 net3 _095_ 0.002383f
C3600 mask\[3\] _289_/a_36_472# 0.02347f
C3601 net53 _451_/a_2225_156# 0.011677f
C3602 FILLER_0_18_2/a_1380_472# _452_/a_448_472# 0.059367f
C3603 _141_ _341_/a_49_472# 0.006222f
C3604 _106_ mask\[1\] 0.005728f
C3605 FILLER_0_4_152/a_124_375# trim_mask\[4\] 0.01182f
C3606 _326_/a_36_160# vdd 0.066545f
C3607 net80 _147_ 0.022618f
C3608 net58 _082_ 0.004276f
C3609 net67 net6 0.345681f
C3610 _430_/a_2248_156# mask\[3\] 0.004211f
C3611 net15 FILLER_0_5_72/a_124_375# 0.006403f
C3612 net58 net82 0.022761f
C3613 FILLER_0_4_152/a_124_375# net47 0.009228f
C3614 net75 cal_itt\[0\] 0.032053f
C3615 _176_ FILLER_0_11_109/a_36_472# 0.002951f
C3616 _208_/a_36_160# vdd 0.014709f
C3617 net62 FILLER_0_15_228/a_124_375# 0.001408f
C3618 _065_ vdd 0.646511f
C3619 FILLER_0_21_150/a_36_472# _146_ 0.00236f
C3620 net55 _216_/a_67_603# 0.071821f
C3621 _370_/a_692_472# _152_ 0.005908f
C3622 _370_/a_1152_472# _081_ 0.001901f
C3623 net57 cal_count\[3\] 0.02848f
C3624 FILLER_0_21_125/a_484_472# net54 0.022347f
C3625 _359_/a_36_488# _062_ 0.005596f
C3626 net69 FILLER_0_3_78/a_124_375# 0.004201f
C3627 _087_ FILLER_0_3_172/a_1916_375# 0.001223f
C3628 fanout70/a_36_113# net70 0.073707f
C3629 mask\[4\] _433_/a_2665_112# 0.005353f
C3630 fanout61/a_36_113# net78 0.009579f
C3631 _343_/a_665_69# mask\[3\] 0.001405f
C3632 _126_ _055_ 0.01647f
C3633 _111_ net55 0.002855f
C3634 _013_ net72 0.006579f
C3635 FILLER_0_13_65/a_124_375# _095_ 0.002035f
C3636 fanout67/a_36_160# trim_val\[0\] 0.003096f
C3637 _414_/a_1000_472# _089_ 0.001754f
C3638 net63 FILLER_0_15_205/a_124_375# 0.001597f
C3639 result[0] FILLER_0_9_282/a_572_375# 0.042859f
C3640 net50 FILLER_0_4_91/a_484_472# 0.008749f
C3641 net82 _082_ 0.286003f
C3642 _127_ _120_ 0.198577f
C3643 net62 _417_/a_1204_472# 0.001941f
C3644 net32 _419_/a_448_472# 0.011757f
C3645 _413_/a_1308_423# net59 0.018948f
C3646 _053_ _312_/a_672_472# 0.001065f
C3647 _151_ vss 0.050544f
C3648 output48/a_224_472# output37/a_224_472# 0.005147f
C3649 FILLER_0_6_47/a_36_472# vss 0.002433f
C3650 FILLER_0_6_47/a_484_472# vdd 0.005065f
C3651 FILLER_0_9_282/a_124_375# vdd 0.01273f
C3652 net15 FILLER_0_15_72/a_36_472# 0.007185f
C3653 net82 fanout57/a_36_113# 0.017696f
C3654 mask\[4\] FILLER_0_20_177/a_484_472# 0.001215f
C3655 fanout58/a_36_160# vss 0.039959f
C3656 mask\[8\] FILLER_0_22_107/a_572_375# 0.030641f
C3657 net35 FILLER_0_22_107/a_124_375# 0.010439f
C3658 output24/a_224_472# vdd 0.08781f
C3659 net16 _217_/a_36_160# 0.00629f
C3660 FILLER_0_16_255/a_36_472# _006_ 0.006621f
C3661 _432_/a_2560_156# _091_ 0.001542f
C3662 FILLER_0_11_135/a_36_472# _120_ 0.012562f
C3663 FILLER_0_16_73/a_36_472# _175_ 0.006803f
C3664 FILLER_0_16_73/a_484_472# vss 0.007212f
C3665 _115_ _449_/a_2665_112# 0.00947f
C3666 cal_count\[2\] _402_/a_718_527# 0.004645f
C3667 _089_ _088_ 0.009863f
C3668 mask\[4\] vdd 0.794539f
C3669 mask\[0\] FILLER_0_12_236/a_36_472# 0.002801f
C3670 _402_/a_1296_93# _179_ 0.001692f
C3671 net70 net53 1.170795f
C3672 _322_/a_124_24# _118_ 0.04952f
C3673 FILLER_0_13_212/a_1020_375# vdd -0.014642f
C3674 FILLER_0_13_212/a_572_375# vss 0.007991f
C3675 _003_ net76 0.080782f
C3676 _429_/a_2665_112# FILLER_0_15_228/a_124_375# 0.001077f
C3677 output34/a_224_472# _106_ 0.01606f
C3678 net38 net49 0.117427f
C3679 FILLER_0_12_136/a_1020_375# _114_ 0.006974f
C3680 _069_ FILLER_0_15_205/a_124_375# 0.002728f
C3681 _395_/a_244_68# _070_ 0.001481f
C3682 FILLER_0_21_142/a_36_472# net35 0.003079f
C3683 net52 _158_ 0.001338f
C3684 FILLER_0_11_101/a_36_472# _120_ 0.007656f
C3685 FILLER_0_10_214/a_36_472# vdd 0.026621f
C3686 FILLER_0_10_214/a_124_375# vss 0.013034f
C3687 _421_/a_1204_472# vdd 0.002198f
C3688 result[9] FILLER_0_24_274/a_932_472# 0.001826f
C3689 _446_/a_1308_423# net17 0.033125f
C3690 fanout63/a_36_160# net36 0.004435f
C3691 net79 _101_ 0.014383f
C3692 _023_ mask\[6\] 0.077441f
C3693 FILLER_0_8_37/a_484_472# _054_ 0.022621f
C3694 result[8] FILLER_0_24_274/a_484_472# 0.005458f
C3695 FILLER_0_19_187/a_124_375# vdd 0.030349f
C3696 FILLER_0_7_162/a_124_375# net57 0.033245f
C3697 _404_/a_36_472# _041_ 0.003068f
C3698 _413_/a_36_151# FILLER_0_3_172/a_1828_472# 0.001723f
C3699 vss FILLER_0_21_60/a_572_375# 0.021222f
C3700 vdd FILLER_0_21_60/a_36_472# 0.08419f
C3701 net26 FILLER_0_23_44/a_484_472# 0.003796f
C3702 FILLER_0_9_223/a_124_375# _128_ 0.004252f
C3703 _105_ _297_/a_36_472# 0.03208f
C3704 _052_ mask\[9\] 0.007224f
C3705 FILLER_0_2_111/a_572_375# vdd 0.012666f
C3706 _429_/a_448_472# net22 0.054866f
C3707 _429_/a_36_151# _018_ 0.118135f
C3708 _093_ FILLER_0_17_104/a_36_472# 0.014431f
C3709 net41 _444_/a_448_472# 0.031876f
C3710 _315_/a_244_497# _059_ 0.00101f
C3711 fanout82/a_36_113# vdd 0.083174f
C3712 FILLER_0_1_98/a_124_375# trim_mask\[3\] 0.058544f
C3713 output47/a_224_472# _452_/a_2225_156# 0.012077f
C3714 _144_ _149_ 0.032178f
C3715 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_36_472# 0.001723f
C3716 net81 net5 0.006276f
C3717 _440_/a_448_472# vdd 0.007263f
C3718 _440_/a_36_151# vss 0.016458f
C3719 net76 net37 0.549565f
C3720 FILLER_0_5_128/a_36_472# _160_ 0.006214f
C3721 net29 _045_ 0.344478f
C3722 _098_ net21 0.133694f
C3723 _256_/a_36_68# vss 0.055568f
C3724 _430_/a_2560_156# _091_ 0.047345f
C3725 FILLER_0_8_37/a_484_472# vss 0.001267f
C3726 _415_/a_448_472# net27 0.05785f
C3727 net66 net49 0.657679f
C3728 FILLER_0_13_65/a_36_472# net72 0.00272f
C3729 _083_ net59 0.408831f
C3730 _132_ mask\[9\] 0.203851f
C3731 FILLER_0_21_28/a_3260_375# _012_ 0.016427f
C3732 net1 net8 0.00497f
C3733 FILLER_0_5_72/a_932_472# vss 0.003084f
C3734 FILLER_0_5_72/a_1380_472# vdd 0.001438f
C3735 net70 FILLER_0_14_107/a_124_375# 0.029975f
C3736 _205_/a_36_160# net21 0.020847f
C3737 _098_ FILLER_0_19_171/a_932_472# 0.003573f
C3738 FILLER_0_20_2/a_124_375# vdd 0.010886f
C3739 net81 FILLER_0_15_235/a_484_472# 0.0047f
C3740 result[5] net62 0.041722f
C3741 FILLER_0_5_54/a_932_472# _029_ 0.014976f
C3742 FILLER_0_5_54/a_1468_375# trim_mask\[1\] 0.010901f
C3743 FILLER_0_16_89/a_1468_375# net14 0.022582f
C3744 _057_ _090_ 0.112325f
C3745 FILLER_0_21_125/a_36_472# _022_ 0.002295f
C3746 _105_ result[8] 0.011678f
C3747 _360_/a_36_160# _163_ 0.008593f
C3748 ctlp[1] _419_/a_36_151# 0.015335f
C3749 _114_ _439_/a_2665_112# 0.011015f
C3750 _410_/a_36_68# cal_count\[0\] 0.007618f
C3751 FILLER_0_8_127/a_36_472# _062_ 0.01783f
C3752 fanout63/a_36_160# FILLER_0_15_228/a_36_472# 0.014197f
C3753 FILLER_0_3_204/a_36_472# FILLER_0_3_212/a_36_472# 0.002296f
C3754 fanout64/a_36_160# calibrate 0.001117f
C3755 net58 FILLER_0_9_270/a_484_472# 0.061043f
C3756 _451_/a_836_156# vdd 0.003786f
C3757 _430_/a_1000_472# net36 0.001836f
C3758 _232_/a_67_603# _167_ 0.014152f
C3759 _062_ FILLER_0_8_156/a_572_375# 0.002944f
C3760 _446_/a_2665_112# net40 0.027712f
C3761 _070_ FILLER_0_10_94/a_36_472# 0.001866f
C3762 _448_/a_36_151# net65 0.001983f
C3763 _426_/a_36_151# FILLER_0_8_247/a_932_472# 0.001723f
C3764 net57 _427_/a_2665_112# 0.016685f
C3765 FILLER_0_5_198/a_124_375# net37 0.009149f
C3766 _130_ vdd 0.046379f
C3767 vdd _034_ 0.424437f
C3768 net42 _039_ 0.001096f
C3769 mask\[5\] FILLER_0_19_171/a_124_375# 0.002206f
C3770 _443_/a_36_151# FILLER_0_2_127/a_36_472# 0.006095f
C3771 _162_ vss 0.08357f
C3772 _161_ vdd 0.262564f
C3773 _421_/a_2665_112# net19 0.01849f
C3774 _430_/a_36_151# FILLER_0_18_209/a_36_472# 0.002841f
C3775 _131_ FILLER_0_9_105/a_484_472# 0.004364f
C3776 net27 net62 0.008623f
C3777 FILLER_0_13_206/a_124_375# _043_ 0.014212f
C3778 _379_/a_36_472# net47 0.016584f
C3779 _053_ net59 0.145863f
C3780 output35/a_224_472# ctlp[2] 0.001465f
C3781 _282_/a_36_160# mask\[2\] 0.023533f
C3782 _095_ _402_/a_56_567# 0.010012f
C3783 _164_ FILLER_0_6_47/a_124_375# 0.069738f
C3784 state\[1\] _055_ 0.067603f
C3785 _129_ vdd 0.314544f
C3786 _131_ vss 0.549133f
C3787 _397_/a_36_472# _175_ 0.004667f
C3788 _070_ calibrate 0.675125f
C3789 _091_ FILLER_0_15_212/a_1380_472# 0.002787f
C3790 output9/a_224_472# _412_/a_1308_423# 0.001352f
C3791 _042_ _039_ 0.003075f
C3792 _165_ trim_mask\[1\] 0.002231f
C3793 output38/a_224_472# FILLER_0_3_2/a_36_472# 0.035046f
C3794 net16 _378_/a_224_472# 0.001007f
C3795 output33/a_224_472# net19 0.12997f
C3796 _431_/a_2248_156# FILLER_0_18_139/a_932_472# 0.001148f
C3797 FILLER_0_7_146/a_36_472# calibrate 0.060587f
C3798 _005_ _193_/a_36_160# 0.009892f
C3799 trim_mask\[2\] fanout49/a_36_160# 0.12844f
C3800 _363_/a_36_68# FILLER_0_7_104/a_572_375# 0.002308f
C3801 _372_/a_3662_472# _062_ 0.0012f
C3802 _418_/a_36_151# _417_/a_36_151# 0.005373f
C3803 net79 _094_ 0.301878f
C3804 _255_/a_224_552# _116_ 0.027303f
C3805 _070_ net21 0.03068f
C3806 _009_ _296_/a_224_472# 0.001278f
C3807 FILLER_0_20_87/a_36_472# _437_/a_36_151# 0.001723f
C3808 _052_ FILLER_0_21_28/a_1468_375# 0.001757f
C3809 result[8] output19/a_224_472# 0.001465f
C3810 FILLER_0_18_37/a_1020_375# vdd 0.020683f
C3811 _056_ net22 0.075673f
C3812 _432_/a_36_151# _333_/a_36_160# 0.032942f
C3813 _399_/a_224_472# vdd 0.001593f
C3814 mask\[3\] FILLER_0_17_161/a_124_375# 0.032905f
C3815 _447_/a_1308_423# net17 0.002531f
C3816 _030_ net14 0.079892f
C3817 _104_ net18 0.039321f
C3818 _429_/a_36_151# vss 0.026298f
C3819 _429_/a_448_472# vdd 0.008822f
C3820 _076_ _080_ 0.005433f
C3821 _294_/a_224_472# _106_ 0.001038f
C3822 _126_ state\[1\] 1.191746f
C3823 _411_/a_36_151# net8 0.012319f
C3824 net18 vss 1.110302f
C3825 _119_ _069_ 0.00226f
C3826 vdd result[3] 0.181788f
C3827 _030_ _164_ 0.036025f
C3828 net52 _066_ 0.022601f
C3829 _053_ _122_ 0.368823f
C3830 net75 FILLER_0_10_247/a_36_472# 0.001184f
C3831 fanout68/a_36_113# vss 0.006152f
C3832 net56 vss 0.367812f
C3833 ctln[5] _448_/a_448_472# 0.010887f
C3834 _255_/a_224_552# _118_ 0.002405f
C3835 output47/a_224_472# net44 0.077292f
C3836 FILLER_0_9_28/a_3172_472# FILLER_0_9_60/a_36_472# 0.013276f
C3837 _426_/a_2665_112# _055_ 0.00142f
C3838 _306_/a_36_68# _113_ 0.010109f
C3839 _437_/a_2560_156# net14 0.00349f
C3840 _096_ vdd 0.557569f
C3841 net80 _098_ 1.289178f
C3842 trim_mask\[1\] FILLER_0_6_79/a_124_375# 0.0042f
C3843 _053_ _169_ 0.014161f
C3844 _068_ net22 0.088209f
C3845 _310_/a_49_472# _090_ 0.059827f
C3846 net52 net23 0.093434f
C3847 _395_/a_1492_488# _121_ 0.002537f
C3848 vdd FILLER_0_22_107/a_124_375# 0.029828f
C3849 net20 FILLER_0_15_212/a_1468_375# 0.006824f
C3850 FILLER_0_13_80/a_36_472# vss 0.009445f
C3851 net58 calibrate 0.205792f
C3852 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_36_472# 0.002296f
C3853 result[4] vdd 0.205815f
C3854 sample fanout65/a_36_113# 0.050978f
C3855 _297_/a_36_472# mask\[6\] 0.02557f
C3856 net72 FILLER_0_21_28/a_572_375# 0.005742f
C3857 ctlp[0] net43 0.003786f
C3858 _431_/a_1204_472# net73 0.026905f
C3859 net78 net79 0.009641f
C3860 _054_ _220_/a_67_603# 0.004333f
C3861 mask\[4\] net63 0.043339f
C3862 _275_/a_224_472# _092_ 0.002138f
C3863 net55 _452_/a_2449_156# 0.015878f
C3864 _068_ _311_/a_2700_473# 0.001846f
C3865 _444_/a_1308_423# net17 0.028709f
C3866 FILLER_0_21_142/a_36_472# vdd 0.111749f
C3867 FILLER_0_18_177/a_3260_375# net21 0.005704f
C3868 ctln[1] vss 0.27233f
C3869 FILLER_0_5_117/a_36_472# FILLER_0_4_107/a_1020_375# 0.001684f
C3870 _394_/a_56_524# _174_ 0.015122f
C3871 _098_ mask\[1\] 1.476748f
C3872 FILLER_0_7_72/a_3172_472# _219_/a_36_160# 0.035111f
C3873 _425_/a_36_151# _122_ 0.063131f
C3874 _425_/a_448_472# calibrate 0.105581f
C3875 ctln[3] _411_/a_1000_472# 0.00283f
C3876 FILLER_0_8_24/a_572_375# net17 0.007101f
C3877 _424_/a_1000_472# _012_ 0.00675f
C3878 net62 FILLER_0_14_235/a_36_472# 0.00534f
C3879 output8/a_224_472# net58 0.018549f
C3880 mask\[5\] FILLER_0_20_177/a_1020_375# 0.013294f
C3881 _033_ _444_/a_1000_472# 0.00692f
C3882 _165_ _444_/a_2665_112# 0.044447f
C3883 FILLER_0_18_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001684f
C3884 _048_ vss 0.056146f
C3885 _232_/a_67_603# vdd 0.007565f
C3886 _417_/a_448_472# vss 0.005289f
C3887 _417_/a_1308_423# vdd 0.002263f
C3888 FILLER_0_4_123/a_36_472# vdd 0.091386f
C3889 fanout76/a_36_160# net18 0.003319f
C3890 FILLER_0_4_123/a_124_375# vss 0.009712f
C3891 net82 calibrate 0.002345f
C3892 FILLER_0_9_28/a_484_472# vdd 0.010868f
C3893 result[8] mask\[6\] 0.111221f
C3894 FILLER_0_19_47/a_484_472# vss 0.001338f
C3895 _220_/a_67_603# vss 0.001485f
C3896 net63 FILLER_0_19_187/a_124_375# 0.012282f
C3897 net18 _416_/a_2248_156# 0.002106f
C3898 trim_mask\[3\] net14 0.142743f
C3899 _421_/a_448_472# _419_/a_2665_112# 0.002393f
C3900 net27 net4 0.025834f
C3901 _016_ _427_/a_448_472# 0.016416f
C3902 _056_ vdd 0.423512f
C3903 net35 FILLER_0_22_86/a_1468_375# 0.010438f
C3904 mask\[8\] FILLER_0_22_86/a_36_472# 0.012471f
C3905 FILLER_0_5_72/a_124_375# net47 0.006974f
C3906 output35/a_224_472# net21 0.069263f
C3907 FILLER_0_7_59/a_36_472# vss 0.004006f
C3908 FILLER_0_7_59/a_484_472# vdd 0.00824f
C3909 FILLER_0_13_212/a_1468_375# _043_ 0.01418f
C3910 _132_ _022_ 0.001404f
C3911 FILLER_0_5_128/a_36_472# _133_ 0.001217f
C3912 _081_ _080_ 0.003905f
C3913 _453_/a_36_151# vdd 0.164654f
C3914 net20 net32 0.006161f
C3915 mask\[4\] _069_ 0.001182f
C3916 net35 FILLER_0_22_128/a_2276_472# 0.014483f
C3917 FILLER_0_15_116/a_36_472# _040_ 0.002896f
C3918 net82 net21 0.037271f
C3919 net22 _201_/a_67_603# 0.004491f
C3920 trim_mask\[2\] net17 0.084388f
C3921 _049_ _146_ 0.042698f
C3922 _164_ trim_mask\[3\] 0.016366f
C3923 FILLER_0_8_107/a_124_375# FILLER_0_9_105/a_484_472# 0.001684f
C3924 FILLER_0_12_2/a_572_375# net67 0.007509f
C3925 _432_/a_36_151# net80 0.035794f
C3926 _170_ vss 0.280383f
C3927 net68 FILLER_0_6_47/a_932_472# 0.014935f
C3928 FILLER_0_11_135/a_124_375# vdd 0.042201f
C3929 output8/a_224_472# net82 0.002936f
C3930 net35 _211_/a_36_160# 0.009886f
C3931 FILLER_0_8_107/a_124_375# vss 0.031335f
C3932 FILLER_0_10_214/a_36_472# _069_ 0.085701f
C3933 _098_ _437_/a_448_472# 0.050691f
C3934 _431_/a_36_151# FILLER_0_17_133/a_36_472# 0.001723f
C3935 FILLER_0_4_49/a_36_472# _167_ 0.063278f
C3936 _074_ vss 0.404343f
C3937 FILLER_0_11_101/a_572_375# FILLER_0_9_105/a_36_472# 0.0027f
C3938 net20 FILLER_0_12_220/a_484_472# 0.001758f
C3939 net55 FILLER_0_18_61/a_124_375# 0.040701f
C3940 _091_ FILLER_0_18_177/a_572_375# 0.004285f
C3941 _077_ _439_/a_1000_472# 0.030609f
C3942 _448_/a_448_472# net59 0.050956f
C3943 _286_/a_224_472# vdd 0.00154f
C3944 _238_/a_67_603# FILLER_0_2_93/a_36_472# 0.002778f
C3945 net3 _185_ 0.004236f
C3946 _106_ output18/a_224_472# 0.005393f
C3947 FILLER_0_11_101/a_572_375# vdd 0.023482f
C3948 FILLER_0_18_2/a_1828_472# vdd 0.001953f
C3949 _127_ _125_ 0.053419f
C3950 net20 _323_/a_36_113# 0.002161f
C3951 _021_ mask\[5\] 0.001088f
C3952 _068_ vdd 0.793549f
C3953 _076_ vss 1.132839f
C3954 _105_ _109_ 0.107328f
C3955 _291_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C3956 net15 cal_count\[1\] 0.089855f
C3957 FILLER_0_17_72/a_2724_472# _438_/a_36_151# 0.002529f
C3958 _052_ _424_/a_36_151# 0.010844f
C3959 cal_itt\[2\] _253_/a_672_68# 0.0016f
C3960 _432_/a_36_151# mask\[1\] 0.003001f
C3961 _429_/a_2665_112# FILLER_0_14_235/a_36_472# 0.007491f
C3962 FILLER_0_12_124/a_124_375# net74 0.049113f
C3963 FILLER_0_15_180/a_36_472# vss 0.00138f
C3964 FILLER_0_15_180/a_484_472# vdd 0.037927f
C3965 mask\[1\] FILLER_0_15_180/a_124_375# 0.004011f
C3966 FILLER_0_4_99/a_124_375# _160_ 0.005563f
C3967 _075_ _074_ 0.058521f
C3968 _238_/a_67_603# trim_mask\[2\] 0.003021f
C3969 _289_/a_36_472# _094_ 0.00922f
C3970 _116_ _120_ 0.005759f
C3971 trim_mask\[2\] FILLER_0_3_78/a_484_472# 0.008122f
C3972 output39/a_224_472# _033_ 0.045759f
C3973 FILLER_0_8_127/a_124_375# _077_ 0.005095f
C3974 output22/a_224_472# net22 0.032714f
C3975 net34 _435_/a_796_472# 0.002288f
C3976 FILLER_0_15_142/a_36_472# _136_ 0.003745f
C3977 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_36_472# 0.002296f
C3978 _086_ _077_ 0.058673f
C3979 fanout51/a_36_113# vdd 0.013496f
C3980 vdd FILLER_0_13_72/a_572_375# -0.001166f
C3981 vss FILLER_0_13_72/a_124_375# 0.043492f
C3982 _057_ _117_ 0.120323f
C3983 output36/a_224_472# _006_ 0.022685f
C3984 _412_/a_448_472# _001_ 0.01124f
C3985 output13/a_224_472# _387_/a_36_113# 0.020974f
C3986 FILLER_0_19_142/a_124_375# _145_ 0.009109f
C3987 _055_ _223_/a_36_160# 0.012271f
C3988 _420_/a_2560_156# _009_ 0.001487f
C3989 sample FILLER_0_9_290/a_124_375# 0.00195f
C3990 _086_ _267_/a_1120_472# 0.004245f
C3991 FILLER_0_20_169/a_124_375# vdd 0.03036f
C3992 FILLER_0_3_204/a_36_472# net22 0.036788f
C3993 en_co_clk vss 0.014954f
C3994 _056_ _373_/a_244_68# 0.00229f
C3995 cal_count\[3\] _453_/a_1000_472# 0.001123f
C3996 net19 _001_ 0.018424f
C3997 _181_ cal_count\[2\] 0.375819f
C3998 _069_ _161_ 0.017831f
C3999 _095_ _451_/a_1040_527# 0.002316f
C4000 _118_ _120_ 0.339442f
C4001 output35/a_224_472# mask\[7\] 0.004608f
C4002 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_484_472# 0.001963f
C4003 FILLER_0_17_72/a_1828_472# net36 0.028046f
C4004 _142_ FILLER_0_17_142/a_572_375# 0.012321f
C4005 _053_ FILLER_0_7_104/a_572_375# 0.005239f
C4006 FILLER_0_12_124/a_36_472# _428_/a_36_151# 0.001723f
C4007 _303_/a_36_472# mask\[9\] 0.013976f
C4008 _093_ _438_/a_2248_156# 0.004221f
C4009 net52 FILLER_0_3_142/a_36_472# 0.001122f
C4010 net69 vdd 1.102677f
C4011 vdd _201_/a_67_603# 0.031337f
C4012 mask\[9\] _438_/a_1204_472# 0.03521f
C4013 _030_ _153_ 0.026157f
C4014 FILLER_0_5_164/a_484_472# vss 0.003257f
C4015 _114_ _017_ 0.071595f
C4016 fanout78/a_36_113# _418_/a_36_151# 0.030244f
C4017 net52 _442_/a_1308_423# 0.017208f
C4018 FILLER_0_18_177/a_932_472# vdd 0.029926f
C4019 FILLER_0_18_177/a_484_472# vss -0.001894f
C4020 _005_ _416_/a_36_151# 0.018752f
C4021 _427_/a_2665_112# net36 0.009904f
C4022 _131_ _095_ 0.043211f
C4023 ctln[2] FILLER_0_0_266/a_124_375# 0.041898f
C4024 _115_ FILLER_0_10_107/a_124_375# 0.011098f
C4025 FILLER_0_9_28/a_1828_472# net51 0.001502f
C4026 net56 FILLER_0_16_154/a_1020_375# 0.002321f
C4027 _339_/a_36_160# FILLER_0_19_155/a_484_472# 0.00304f
C4028 _450_/a_2449_156# _039_ 0.013285f
C4029 net18 _419_/a_1000_472# 0.008295f
C4030 FILLER_0_19_28/a_124_375# _452_/a_36_151# 0.002709f
C4031 net16 FILLER_0_18_37/a_1380_472# 0.002932f
C4032 net57 net52 0.016136f
C4033 FILLER_0_24_130/a_124_375# ctlp[7] 0.002726f
C4034 output21/a_224_472# result[8] 0.149245f
C4035 net69 _441_/a_1204_472# 0.014374f
C4036 output20/a_224_472# _422_/a_36_151# 0.053592f
C4037 FILLER_0_17_104/a_1020_375# net14 0.002226f
C4038 _411_/a_2665_112# net19 0.00934f
C4039 _412_/a_36_151# net2 0.003823f
C4040 _114_ FILLER_0_10_107/a_36_472# 0.00263f
C4041 FILLER_0_21_125/a_484_472# _144_ 0.001616f
C4042 _216_/a_67_603# FILLER_0_18_61/a_124_375# 0.014522f
C4043 _425_/a_1000_472# vdd 0.019072f
C4044 result[7] _046_ 0.003397f
C4045 net73 FILLER_0_18_107/a_2724_472# 0.02814f
C4046 _069_ _429_/a_448_472# 0.035108f
C4047 net37 FILLER_0_6_231/a_36_472# 0.002982f
C4048 _152_ vdd 0.354509f
C4049 _081_ vss 0.733408f
C4050 net35 net71 0.042275f
C4051 mask\[7\] FILLER_0_22_128/a_932_472# 0.017448f
C4052 _053_ FILLER_0_7_72/a_1828_472# 0.013271f
C4053 _115_ FILLER_0_9_142/a_124_375# 0.010167f
C4054 _091_ _274_/a_3368_68# 0.001328f
C4055 _070_ _171_ 0.084342f
C4056 ctln[5] net12 0.41364f
C4057 net64 FILLER_0_9_270/a_36_472# 0.014971f
C4058 net53 _427_/a_1204_472# 0.004293f
C4059 FILLER_0_9_28/a_572_375# net16 0.042681f
C4060 _002_ FILLER_0_3_172/a_2724_472# 0.006713f
C4061 _067_ FILLER_0_12_20/a_36_472# 0.015608f
C4062 _448_/a_1204_472# net22 0.002283f
C4063 net15 FILLER_0_17_72/a_124_375# 0.006492f
C4064 _098_ FILLER_0_15_212/a_124_375# 0.008125f
C4065 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_484_472# 0.013277f
C4066 FILLER_0_18_76/a_484_472# _438_/a_36_151# 0.001723f
C4067 cal_itt\[2\] FILLER_0_3_221/a_1380_472# 0.015024f
C4068 net60 ctlp[1] 0.073021f
C4069 _099_ _098_ 0.018316f
C4070 net50 _439_/a_1000_472# 0.005154f
C4071 net52 _439_/a_2248_156# 0.00258f
C4072 _093_ mask\[8\] 0.004026f
C4073 _138_ vdd 0.090752f
C4074 net23 FILLER_0_8_156/a_36_472# 0.004939f
C4075 FILLER_0_4_49/a_36_472# vdd 0.090733f
C4076 FILLER_0_4_49/a_572_375# vss 0.008729f
C4077 _075_ _081_ 0.001195f
C4078 net54 _438_/a_2248_156# 0.014423f
C4079 net65 vss 0.471168f
C4080 FILLER_0_9_28/a_1916_375# _453_/a_36_151# 0.001543f
C4081 output22/a_224_472# vdd 0.111234f
C4082 trim[0] output40/a_224_472# 0.005306f
C4083 net38 net40 1.103743f
C4084 result[9] vdd 0.597071f
C4085 FILLER_0_15_142/a_36_472# net53 0.080484f
C4086 _307_/a_672_472# _126_ 0.00121f
C4087 _098_ FILLER_0_19_111/a_124_375# 0.001331f
C4088 net56 _095_ 0.004847f
C4089 ctlp[9] net26 0.02213f
C4090 net32 _009_ 0.003756f
C4091 _136_ _337_/a_665_69# 0.001794f
C4092 _015_ FILLER_0_8_247/a_932_472# 0.005458f
C4093 FILLER_0_9_28/a_36_472# FILLER_0_10_28/a_36_472# 0.05841f
C4094 _176_ FILLER_0_10_107/a_36_472# 0.009019f
C4095 _117_ _310_/a_49_472# 0.018229f
C4096 FILLER_0_3_204/a_36_472# vdd 0.092654f
C4097 FILLER_0_22_86/a_1468_375# vdd 0.035441f
C4098 net15 _120_ 0.028275f
C4099 net15 _038_ 0.078028f
C4100 net76 _037_ 0.010891f
C4101 FILLER_0_11_78/a_36_472# _120_ 0.014169f
C4102 _038_ FILLER_0_11_78/a_36_472# 0.001782f
C4103 _036_ fanout68/a_36_113# 0.007847f
C4104 FILLER_0_17_104/a_1380_472# FILLER_0_16_115/a_124_375# 0.001723f
C4105 FILLER_0_5_212/a_124_375# FILLER_0_3_212/a_36_472# 0.001512f
C4106 _095_ FILLER_0_13_80/a_36_472# 0.004187f
C4107 FILLER_0_22_128/a_2276_472# vdd 0.00565f
C4108 FILLER_0_22_128/a_1828_472# vss 0.009137f
C4109 FILLER_0_9_290/a_124_375# FILLER_0_9_282/a_572_375# 0.012001f
C4110 net81 FILLER_0_12_236/a_484_472# 0.001419f
C4111 result[8] _422_/a_1308_423# 0.001356f
C4112 ctlp[3] _422_/a_448_472# 0.001441f
C4113 _086_ _363_/a_692_472# 0.001353f
C4114 FILLER_0_8_138/a_36_472# _076_ 0.016628f
C4115 _077_ _313_/a_67_603# 0.007446f
C4116 net56 FILLER_0_18_139/a_484_472# 0.004375f
C4117 _412_/a_36_151# valid 0.009757f
C4118 fanout59/a_36_160# net59 0.021522f
C4119 _211_/a_36_160# vdd 0.030216f
C4120 FILLER_0_15_235/a_124_375# FILLER_0_14_235/a_124_375# 0.05841f
C4121 _094_ net19 0.06304f
C4122 FILLER_0_7_72/a_932_472# _053_ 0.01339f
C4123 _425_/a_2248_156# net19 0.010557f
C4124 _013_ vdd 0.372605f
C4125 _445_/a_1308_423# _034_ 0.002494f
C4126 _137_ _097_ 0.001654f
C4127 net66 net40 0.124825f
C4128 net17 output6/a_224_472# 0.047757f
C4129 net36 FILLER_0_18_76/a_572_375# 0.005153f
C4130 _185_ _402_/a_56_567# 0.107713f
C4131 net82 FILLER_0_3_172/a_484_472# 0.008052f
C4132 output45/a_224_472# vdd -0.026726f
C4133 FILLER_0_14_50/a_124_375# _179_ 0.021823f
C4134 net54 mask\[8\] 0.162104f
C4135 _067_ FILLER_0_12_28/a_36_472# 0.0127f
C4136 _067_ net40 0.040115f
C4137 FILLER_0_3_172/a_3260_375# net65 0.002696f
C4138 _322_/a_124_24# net74 0.05722f
C4139 net58 output48/a_224_472# 0.065357f
C4140 _091_ _136_ 0.075998f
C4141 FILLER_0_7_72/a_124_375# net52 0.029774f
C4142 ctlp[2] mask\[7\] 0.036719f
C4143 _132_ FILLER_0_11_109/a_124_375# 0.008627f
C4144 _069_ _056_ 0.035189f
C4145 FILLER_0_15_116/a_484_472# vss 0.003923f
C4146 _091_ net62 0.019946f
C4147 _443_/a_1308_423# vdd 0.00203f
C4148 _443_/a_448_472# vss 0.030448f
C4149 _120_ net51 1.716752f
C4150 fanout76/a_36_160# net65 0.018025f
C4151 FILLER_0_5_117/a_36_472# vss 0.001215f
C4152 ctlp[3] _108_ 0.009437f
C4153 net20 mask\[3\] 0.047107f
C4154 _415_/a_2248_156# output27/a_224_472# 0.001506f
C4155 output48/a_224_472# _425_/a_448_472# 0.001155f
C4156 _448_/a_1204_472# vdd 0.002228f
C4157 _272_/a_36_472# vdd 0.058326f
C4158 FILLER_0_16_107/a_484_472# vdd 0.02929f
C4159 net52 FILLER_0_6_47/a_2276_472# 0.003298f
C4160 net15 mask\[8\] 0.02403f
C4161 _020_ net70 0.014391f
C4162 calibrate net21 0.036773f
C4163 mask\[4\] _140_ 0.001697f
C4164 net12 net59 0.001028f
C4165 _090_ vss 0.267577f
C4166 _113_ vdd 0.774039f
C4167 _137_ mask\[2\] 0.440828f
C4168 _028_ FILLER_0_6_79/a_36_472# 0.016281f
C4169 _131_ _332_/a_36_472# 0.006825f
C4170 _425_/a_36_151# FILLER_0_8_247/a_572_375# 0.001597f
C4171 _392_/a_244_472# _067_ 0.001893f
C4172 FILLER_0_16_57/a_1020_375# net72 0.002937f
C4173 output48/a_224_472# _082_ 0.002393f
C4174 output37/a_224_472# net18 0.046654f
C4175 net15 FILLER_0_17_56/a_484_472# 0.001758f
C4176 FILLER_0_5_54/a_36_472# net47 0.00679f
C4177 _041_ FILLER_0_18_37/a_1380_472# 0.003776f
C4178 net68 _453_/a_448_472# 0.01245f
C4179 fanout59/a_36_160# net64 0.006298f
C4180 net57 _428_/a_1308_423# 0.018725f
C4181 FILLER_0_3_54/a_124_375# net40 0.005766f
C4182 output48/a_224_472# net82 0.048965f
C4183 _086_ _375_/a_960_497# 0.001454f
C4184 FILLER_0_7_72/a_3172_472# _058_ 0.001085f
C4185 net78 _108_ 0.056528f
C4186 _433_/a_2560_156# _145_ 0.007651f
C4187 FILLER_0_17_56/a_124_375# _041_ 0.001489f
C4188 net74 _372_/a_786_69# 0.00149f
C4189 FILLER_0_16_89/a_1020_375# _136_ 0.019549f
C4190 _413_/a_2665_112# net82 0.004306f
C4191 net78 net19 0.507249f
C4192 _069_ _068_ 0.003779f
C4193 ctln[2] net81 0.003762f
C4194 _414_/a_36_151# net21 0.007791f
C4195 FILLER_0_17_72/a_3260_375# vdd 0.007427f
C4196 _134_ FILLER_0_10_107/a_124_375# 0.009573f
C4197 FILLER_0_12_20/a_484_472# net47 0.020293f
C4198 _136_ FILLER_0_17_142/a_124_375# 0.001315f
C4199 cal_itt\[3\] _087_ 0.002881f
C4200 FILLER_0_8_263/a_36_472# net19 0.047387f
C4201 net3 net17 0.045911f
C4202 result[5] _419_/a_36_151# 0.006539f
C4203 output45/a_224_472# output17/a_224_472# 0.071473f
C4204 FILLER_0_16_89/a_36_472# _451_/a_2449_156# 0.001571f
C4205 FILLER_0_4_107/a_1380_472# vdd 0.007022f
C4206 vdd FILLER_0_6_37/a_124_375# 0.041381f
C4207 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001597f
C4208 net15 _175_ 0.052586f
C4209 _132_ FILLER_0_17_104/a_124_375# 0.001918f
C4210 result[6] FILLER_0_21_286/a_36_472# 0.015369f
C4211 _427_/a_448_472# vss 0.040679f
C4212 _427_/a_1308_423# vdd 0.002814f
C4213 trim_mask\[4\] _370_/a_848_380# 0.027744f
C4214 net72 FILLER_0_15_59/a_36_472# 0.049812f
C4215 output7/a_224_472# vss 0.00746f
C4216 net52 FILLER_0_2_111/a_484_472# 0.061249f
C4217 _029_ vss 0.11129f
C4218 _308_/a_848_380# _219_/a_36_160# 0.001045f
C4219 _043_ FILLER_0_13_72/a_36_472# 0.017766f
C4220 net41 _402_/a_728_93# 0.032823f
C4221 _091_ _429_/a_2665_112# 0.002597f
C4222 ctlp[2] _422_/a_2248_156# 0.001328f
C4223 cal_count\[3\] _405_/a_67_603# 0.011131f
C4224 FILLER_0_13_65/a_36_472# vdd 0.005885f
C4225 _370_/a_848_380# net47 0.004223f
C4226 FILLER_0_2_101/a_124_375# _154_ 0.003932f
C4227 FILLER_0_19_55/a_36_472# net36 0.001068f
C4228 _093_ FILLER_0_17_133/a_36_472# 0.010432f
C4229 trim_mask\[2\] FILLER_0_2_93/a_36_472# 0.281054f
C4230 FILLER_0_21_142/a_36_472# FILLER_0_21_133/a_36_472# 0.001963f
C4231 net63 FILLER_0_18_177/a_932_472# 0.063742f
C4232 _449_/a_36_151# _453_/a_36_151# 0.007757f
C4233 net52 _440_/a_1204_472# 0.003916f
C4234 net60 _421_/a_2560_156# 0.001951f
C4235 vss _145_ 0.399701f
C4236 FILLER_0_7_72/a_1468_375# net52 0.003576f
C4237 net5 net59 0.923076f
C4238 _414_/a_448_472# net21 0.040301f
C4239 _452_/a_448_472# _041_ 0.007f
C4240 _086_ cal_itt\[3\] 0.046874f
C4241 _178_ _408_/a_56_524# 0.014421f
C4242 net71 vdd 0.775031f
C4243 net49 _440_/a_1204_472# 0.006692f
C4244 output39/a_224_472# _444_/a_36_151# 0.062717f
C4245 FILLER_0_9_28/a_2812_375# vdd 0.016637f
C4246 net38 FILLER_0_15_2/a_484_472# 0.003391f
C4247 _235_/a_67_603# _064_ 0.003796f
C4248 en_co_clk _095_ 0.003753f
C4249 _350_/a_49_472# mask\[6\] 0.033488f
C4250 _415_/a_2248_156# _416_/a_36_151# 0.001495f
C4251 _447_/a_1204_472# vdd 0.001085f
C4252 FILLER_0_16_89/a_36_472# net36 0.010907f
C4253 _091_ FILLER_0_19_171/a_124_375# 0.028992f
C4254 net57 FILLER_0_8_156/a_36_472# 0.001544f
C4255 _114_ cal_count\[3\] 0.081644f
C4256 result[4] net77 0.003336f
C4257 net23 FILLER_0_22_128/a_2364_375# 0.018463f
C4258 _132_ FILLER_0_19_134/a_124_375# 0.00141f
C4259 FILLER_0_17_64/a_36_472# net36 0.00195f
C4260 _137_ FILLER_0_16_154/a_484_472# 0.00631f
C4261 _183_ _180_ 0.002621f
C4262 FILLER_0_19_125/a_36_472# _145_ 0.004858f
C4263 _314_/a_224_472# vss 0.001399f
C4264 net54 _433_/a_2248_156# 0.04755f
C4265 _093_ FILLER_0_18_107/a_124_375# 0.008393f
C4266 _447_/a_2665_112# _168_ 0.001107f
C4267 FILLER_0_5_72/a_36_472# _440_/a_36_151# 0.001723f
C4268 _164_ FILLER_0_6_47/a_3172_472# 0.001058f
C4269 FILLER_0_0_198/a_36_472# vss 0.00344f
C4270 _077_ FILLER_0_9_72/a_124_375# 0.008103f
C4271 _155_ vss 0.13648f
C4272 fanout60/a_36_160# net79 0.069956f
C4273 output22/a_224_472# net63 0.017997f
C4274 net15 _453_/a_2560_156# 0.049334f
C4275 _035_ _164_ 0.056332f
C4276 mask\[7\] net21 0.050718f
C4277 _308_/a_1084_68# net14 0.002892f
C4278 _091_ net4 0.125608f
C4279 FILLER_0_14_81/a_36_472# _394_/a_1936_472# 0.010394f
C4280 net74 _370_/a_848_380# 0.004546f
C4281 _365_/a_244_472# _156_ 0.003847f
C4282 _141_ _339_/a_36_160# 0.011118f
C4283 _077_ _061_ 0.031458f
C4284 _444_/a_1000_472# _054_ 0.002998f
C4285 _053_ FILLER_0_4_213/a_572_375# 0.003451f
C4286 trim[4] trim[1] 0.001879f
C4287 _077_ _453_/a_1308_423# 0.071515f
C4288 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_36_472# 0.001963f
C4289 _077_ _311_/a_66_473# 0.002605f
C4290 FILLER_0_8_24/a_484_472# _054_ 0.009315f
C4291 net64 net5 0.098088f
C4292 output8/a_224_472# _411_/a_448_472# 0.010723f
C4293 _449_/a_36_151# FILLER_0_13_72/a_572_375# 0.035849f
C4294 FILLER_0_7_72/a_1380_472# _053_ 0.01339f
C4295 _059_ FILLER_0_5_136/a_36_472# 0.001755f
C4296 cal_count\[1\] FILLER_0_15_59/a_484_472# 0.006408f
C4297 _132_ net57 0.029479f
C4298 net80 net21 0.016911f
C4299 net65 FILLER_0_2_177/a_36_472# 0.016652f
C4300 _125_ _118_ 0.239695f
C4301 net16 cal_count\[3\] 0.082821f
C4302 _354_/a_49_472# _098_ 0.009677f
C4303 _029_ FILLER_0_5_88/a_124_375# 0.006771f
C4304 _103_ _418_/a_36_151# 0.032388f
C4305 net80 _333_/a_36_160# 0.001594f
C4306 _176_ cal_count\[3\] 0.067683f
C4307 result[7] _103_ 0.298427f
C4308 _025_ _436_/a_2248_156# 0.001054f
C4309 _076_ _385_/a_36_68# 0.006512f
C4310 ctlp[1] FILLER_0_23_290/a_124_375# 0.053745f
C4311 _078_ net37 0.459092f
C4312 FILLER_0_7_72/a_2276_472# FILLER_0_6_90/a_124_375# 0.001684f
C4313 net33 _434_/a_448_472# 0.003049f
C4314 net64 FILLER_0_15_235/a_484_472# 0.005893f
C4315 _102_ net36 0.003446f
C4316 trim_mask\[2\] FILLER_0_4_91/a_124_375# 0.003591f
C4317 _444_/a_1204_472# vdd 0.001086f
C4318 state\[0\] FILLER_0_12_220/a_1380_472# 0.003733f
C4319 _411_/a_36_151# _073_ 0.00135f
C4320 FILLER_0_7_233/a_36_472# vss 0.005354f
C4321 FILLER_0_0_232/a_36_472# vdd 0.050082f
C4322 FILLER_0_0_232/a_124_375# vss 0.019863f
C4323 net31 output31/a_224_472# 0.002146f
C4324 _053_ trim_val\[0\] 0.446477f
C4325 _088_ _269_/a_36_472# 0.004438f
C4326 net78 _419_/a_448_472# 0.0122f
C4327 net54 FILLER_0_18_107/a_124_375# 0.001636f
C4328 _219_/a_36_160# net14 0.048037f
C4329 _136_ net14 0.417108f
C4330 net11 vss 0.057193f
C4331 _453_/a_2560_156# net51 0.013556f
C4332 mask\[1\] net21 0.023956f
C4333 FILLER_0_4_144/a_572_375# net23 0.019114f
C4334 _440_/a_2665_112# _164_ 0.067034f
C4335 _077_ _072_ 0.178678f
C4336 FILLER_0_4_144/a_36_472# trim_mask\[4\] 0.017557f
C4337 _375_/a_36_68# _162_ 0.011065f
C4338 _375_/a_1612_497# _161_ 0.003325f
C4339 _163_ vss 0.638066f
C4340 net38 _452_/a_1040_527# 0.002024f
C4341 FILLER_0_4_49/a_484_472# net68 0.027016f
C4342 FILLER_0_20_2/a_124_375# net43 0.001563f
C4343 _291_/a_36_160# _092_ 0.03297f
C4344 _010_ _420_/a_2665_112# 0.029378f
C4345 _431_/a_448_472# vdd 0.001932f
C4346 _438_/a_1000_472# net14 0.003275f
C4347 FILLER_0_4_144/a_36_472# net47 0.008498f
C4348 output35/a_224_472# FILLER_0_22_177/a_1468_375# 0.018187f
C4349 FILLER_0_4_185/a_124_375# net22 0.004776f
C4350 _130_ FILLER_0_11_124/a_124_375# 0.001943f
C4351 _273_/a_36_68# vdd 0.041825f
C4352 FILLER_0_21_28/a_572_375# vdd 0.013051f
C4353 _451_/a_1697_156# net14 0.001298f
C4354 output15/a_224_472# vss 0.067969f
C4355 FILLER_0_14_91/a_36_472# en_co_clk 0.007733f
C4356 FILLER_0_11_78/a_124_375# vss 0.006233f
C4357 FILLER_0_11_78/a_572_375# vdd -0.006646f
C4358 FILLER_0_15_72/a_484_472# _451_/a_3129_107# 0.005866f
C4359 net32 net33 0.467071f
C4360 fanout74/a_36_113# _371_/a_36_113# 0.01088f
C4361 FILLER_0_18_2/a_2276_472# vss 0.001865f
C4362 FILLER_0_0_96/a_36_472# trim_mask\[3\] 0.005343f
C4363 _144_ FILLER_0_22_128/a_2812_375# 0.001601f
C4364 _064_ vdd 0.874293f
C4365 net82 FILLER_0_4_213/a_124_375# 0.00123f
C4366 FILLER_0_6_239/a_36_472# _123_ 0.004433f
C4367 net67 FILLER_0_9_60/a_124_375# 0.003083f
C4368 FILLER_0_21_142/a_36_472# _140_ 0.009261f
C4369 FILLER_0_22_86/a_932_472# _149_ 0.001205f
C4370 FILLER_0_22_86/a_36_472# _026_ 0.001503f
C4371 _430_/a_448_472# net22 0.036303f
C4372 _253_/a_1732_68# cal_itt\[1\] 0.001829f
C4373 _131_ FILLER_0_11_124/a_36_472# 0.015445f
C4374 _086_ _325_/a_224_472# 0.003155f
C4375 _058_ _062_ 1.676625f
C4376 output39/a_224_472# _054_ 0.002121f
C4377 net39 _221_/a_36_160# 0.059979f
C4378 FILLER_0_4_107/a_124_375# net47 0.004586f
C4379 net15 _441_/a_1000_472# 0.025912f
C4380 output42/a_224_472# net40 0.003278f
C4381 _002_ _088_ 0.003969f
C4382 FILLER_0_6_90/a_124_375# vdd 0.020992f
C4383 _371_/a_36_113# FILLER_0_2_127/a_124_375# 0.002437f
C4384 net42 vdd 0.178782f
C4385 output29/a_224_472# _005_ 0.021351f
C4386 _418_/a_796_472# vss 0.00145f
C4387 _053_ _119_ 0.038651f
C4388 _093_ FILLER_0_17_161/a_36_472# 0.006224f
C4389 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_124_375# 0.012001f
C4390 FILLER_0_10_28/a_36_472# net51 0.00703f
C4391 _171_ FILLER_0_10_94/a_36_472# 0.001514f
C4392 _172_ FILLER_0_10_94/a_124_375# 0.003341f
C4393 FILLER_0_22_177/a_932_472# net33 0.014021f
C4394 _433_/a_1204_472# _022_ 0.005308f
C4395 _426_/a_2248_156# _076_ 0.015189f
C4396 _000_ net58 0.00389f
C4397 net52 FILLER_0_9_72/a_1020_375# 0.00799f
C4398 FILLER_0_21_286/a_484_472# vss 0.008522f
C4399 net80 mask\[7\] 0.020051f
C4400 FILLER_0_15_116/a_484_472# _095_ 0.001069f
C4401 FILLER_0_13_142/a_572_375# net23 0.009573f
C4402 FILLER_0_4_99/a_36_472# FILLER_0_4_107/a_36_472# 0.002296f
C4403 FILLER_0_19_187/a_484_472# _434_/a_2665_112# 0.001868f
C4404 _130_ _428_/a_2248_156# 0.006602f
C4405 FILLER_0_1_266/a_36_472# vdd 0.008551f
C4406 FILLER_0_1_266/a_572_375# vss 0.001919f
C4407 _042_ vdd 0.261947f
C4408 _069_ _113_ 0.027402f
C4409 _079_ _112_ 0.004464f
C4410 _117_ vss 0.048946f
C4411 _081_ _385_/a_36_68# 0.006303f
C4412 _331_/a_448_472# _134_ 0.001126f
C4413 FILLER_0_5_206/a_36_472# vss 0.003493f
C4414 _077_ FILLER_0_9_60/a_572_375# 0.018665f
C4415 fanout56/a_36_113# _097_ 0.062226f
C4416 net75 _426_/a_36_151# 0.070626f
C4417 _428_/a_2665_112# _131_ 0.006081f
C4418 output48/a_224_472# calibrate 0.003223f
C4419 _176_ FILLER_0_17_72/a_1828_472# 0.001028f
C4420 net53 net14 0.04525f
C4421 output37/a_224_472# net65 0.096416f
C4422 net82 FILLER_0_3_221/a_572_375# 0.005424f
C4423 FILLER_0_9_28/a_124_375# net17 0.009179f
C4424 _412_/a_36_151# cal_itt\[1\] 0.025078f
C4425 _075_ FILLER_0_5_206/a_36_472# 0.001503f
C4426 vdd FILLER_0_4_91/a_484_472# 0.007304f
C4427 input2/a_36_113# clk 0.021981f
C4428 FILLER_0_1_98/a_36_472# vss 0.002275f
C4429 FILLER_0_8_247/a_124_375# calibrate 0.008393f
C4430 FILLER_0_12_220/a_124_375# _090_ 0.001521f
C4431 ctlp[1] FILLER_0_24_274/a_484_472# 0.001875f
C4432 _000_ net82 0.032846f
C4433 output32/a_224_472# output31/a_224_472# 0.00289f
C4434 net1 net2 0.624657f
C4435 FILLER_0_5_212/a_124_375# vdd 0.024541f
C4436 FILLER_0_13_212/a_572_375# _070_ 0.003986f
C4437 FILLER_0_3_172/a_1828_472# net22 0.009883f
C4438 FILLER_0_8_37/a_572_375# _220_/a_67_603# 0.00744f
C4439 _021_ _091_ 0.016024f
C4440 FILLER_0_4_185/a_124_375# vdd 0.02924f
C4441 _028_ FILLER_0_8_107/a_36_472# 0.002173f
C4442 _422_/a_2248_156# mask\[7\] 0.015008f
C4443 net41 _160_ 0.006523f
C4444 _071_ _314_/a_224_472# 0.001359f
C4445 result[6] _420_/a_2248_156# 0.003418f
C4446 _414_/a_2248_156# FILLER_0_5_212/a_36_472# 0.035805f
C4447 net80 mask\[1\] 0.015535f
C4448 _116_ _043_ 0.002037f
C4449 _413_/a_2665_112# net21 0.002828f
C4450 net20 _014_ 0.008597f
C4451 FILLER_0_10_214/a_124_375# _070_ 0.017713f
C4452 output30/a_224_472# result[3] 0.019025f
C4453 output38/a_224_472# vdd -0.006652f
C4454 net74 _120_ 0.027885f
C4455 _093_ _150_ 0.406318f
C4456 _004_ _415_/a_448_472# 0.044374f
C4457 net74 _038_ 0.055774f
C4458 _427_/a_448_472# _095_ 0.063616f
C4459 net27 _426_/a_1308_423# 0.00384f
C4460 _053_ FILLER_0_6_47/a_484_472# 0.006301f
C4461 _093_ FILLER_0_17_72/a_3172_472# 0.012002f
C4462 FILLER_0_16_37/a_124_375# _179_ 0.005434f
C4463 mask\[0\] net21 0.050431f
C4464 _446_/a_36_151# trim[3] 0.00699f
C4465 net16 _408_/a_2215_68# 0.002096f
C4466 net31 _008_ 0.292444f
C4467 _430_/a_448_472# vdd 0.002959f
C4468 output8/a_224_472# _413_/a_2665_112# 0.010726f
C4469 _321_/a_170_472# _126_ 0.018831f
C4470 _408_/a_718_524# _043_ 0.003719f
C4471 _066_ _386_/a_848_380# 0.00416f
C4472 fanout52/a_36_160# trim_mask\[4\] 0.014356f
C4473 FILLER_0_5_198/a_484_472# net59 0.059394f
C4474 FILLER_0_9_223/a_124_375# _246_/a_36_68# 0.005308f
C4475 _431_/a_36_151# FILLER_0_18_107/a_3172_472# 0.00271f
C4476 FILLER_0_1_266/a_36_472# net9 0.041635f
C4477 FILLER_0_16_73/a_484_472# net55 0.004188f
C4478 FILLER_0_5_54/a_484_472# FILLER_0_6_47/a_1380_472# 0.026657f
C4479 FILLER_0_5_54/a_1468_375# FILLER_0_6_47/a_2276_472# 0.001597f
C4480 _428_/a_448_472# _017_ 0.056f
C4481 _428_/a_36_151# net53 0.001124f
C4482 fanout53/a_36_160# net56 0.196684f
C4483 FILLER_0_16_57/a_484_472# FILLER_0_17_56/a_572_375# 0.001723f
C4484 _369_/a_36_68# vdd 0.042534f
C4485 _044_ vdd 0.406979f
C4486 _192_/a_67_603# _044_ 0.002571f
C4487 _105_ ctlp[1] 0.158795f
C4488 _408_/a_56_524# _095_ 0.01643f
C4489 FILLER_0_20_169/a_124_375# _140_ 0.01799f
C4490 _177_ cal_count\[1\] 0.03631f
C4491 net76 _123_ 0.003431f
C4492 _104_ _422_/a_2560_156# 0.003223f
C4493 cal_itt\[2\] net75 0.143064f
C4494 _431_/a_2665_112# vdd 0.015335f
C4495 FILLER_0_2_177/a_484_472# net59 0.007829f
C4496 _256_/a_36_68# _070_ 0.019259f
C4497 FILLER_0_11_142/a_36_472# vss 0.008744f
C4498 FILLER_0_11_142/a_484_472# vdd 0.006641f
C4499 net45 vdd 0.087369f
C4500 _322_/a_1152_472# _129_ 0.002978f
C4501 net41 FILLER_0_18_37/a_124_375# 0.004639f
C4502 FILLER_0_18_107/a_3260_375# vdd 0.004983f
C4503 FILLER_0_18_107/a_2812_375# vss 0.002392f
C4504 _073_ net76 0.040554f
C4505 FILLER_0_4_144/a_36_472# FILLER_0_3_142/a_124_375# 0.001543f
C4506 state\[1\] _121_ 0.006184f
C4507 _434_/a_1308_423# mask\[6\] 0.022677f
C4508 net58 fanout58/a_36_160# 0.013794f
C4509 output31/a_224_472# FILLER_0_16_255/a_124_375# 0.001274f
C4510 FILLER_0_7_104/a_1468_375# vdd 0.026224f
C4511 _004_ net62 0.001201f
C4512 _173_ _120_ 0.004205f
C4513 net79 FILLER_0_12_220/a_1380_472# 0.010583f
C4514 FILLER_0_18_139/a_484_472# _145_ 0.002415f
C4515 net47 _386_/a_692_472# 0.003299f
C4516 FILLER_0_3_221/a_36_472# FILLER_0_3_212/a_36_472# 0.001963f
C4517 _239_/a_36_160# net41 0.006002f
C4518 FILLER_0_12_124/a_36_472# _017_ 0.004641f
C4519 result[6] _419_/a_2665_112# 0.001225f
C4520 output29/a_224_472# _416_/a_448_472# 0.008149f
C4521 _074_ _375_/a_36_68# 0.003157f
C4522 valid net1 0.00347f
C4523 mask\[4\] FILLER_0_18_177/a_2812_375# 0.013557f
C4524 trim_val\[4\] _386_/a_1084_68# 0.002659f
C4525 FILLER_0_5_109/a_484_472# FILLER_0_4_107/a_572_375# 0.001684f
C4526 net55 FILLER_0_21_60/a_572_375# 0.041903f
C4527 FILLER_0_15_142/a_572_375# net74 0.001652f
C4528 fanout78/a_36_113# _007_ 0.003126f
C4529 trim_val\[1\] FILLER_0_6_47/a_36_472# 0.00351f
C4530 FILLER_0_16_57/a_1468_375# _175_ 0.001654f
C4531 net52 _441_/a_36_151# 0.013755f
C4532 _308_/a_848_380# _058_ 0.031449f
C4533 FILLER_0_4_107/a_124_375# _154_ 0.00183f
C4534 mask\[3\] FILLER_0_18_177/a_1916_375# 0.003052f
C4535 _447_/a_1000_472# _036_ 0.002902f
C4536 trimb[1] output44/a_224_472# 0.046391f
C4537 net54 _150_ 0.001162f
C4538 FILLER_0_4_144/a_572_375# net57 0.001254f
C4539 FILLER_0_23_88/a_36_472# vss 0.003481f
C4540 _133_ _160_ 0.043549f
C4541 result[5] net60 0.16275f
C4542 net24 _050_ 0.049889f
C4543 net20 _094_ 0.677838f
C4544 _122_ FILLER_0_5_198/a_484_472# 0.002999f
C4545 _030_ _384_/a_224_472# 0.003019f
C4546 _417_/a_1308_423# output30/a_224_472# 0.001434f
C4547 _417_/a_36_151# net30 0.010021f
C4548 net47 _452_/a_836_156# 0.002075f
C4549 input5/a_36_113# rstn 0.019149f
C4550 _062_ _226_/a_860_68# 0.001842f
C4551 _072_ _375_/a_960_497# 0.001322f
C4552 _441_/a_448_472# _030_ 0.038429f
C4553 _441_/a_36_151# net49 0.010951f
C4554 FILLER_0_13_65/a_36_472# _449_/a_36_151# 0.001723f
C4555 _208_/a_36_160# _049_ 0.04568f
C4556 _431_/a_2248_156# _427_/a_36_151# 0.001081f
C4557 net64 _055_ 0.00384f
C4558 net15 _423_/a_2665_112# 0.061217f
C4559 _093_ FILLER_0_18_139/a_1468_375# 0.004939f
C4560 _328_/a_36_113# FILLER_0_11_101/a_484_472# 0.001826f
C4561 _437_/a_1000_472# vdd 0.001777f
C4562 _428_/a_36_151# FILLER_0_14_107/a_124_375# 0.001597f
C4563 cal_itt\[3\] _061_ 0.001311f
C4564 _449_/a_2665_112# _038_ 0.024406f
C4565 FILLER_0_18_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001684f
C4566 FILLER_0_3_172/a_1828_472# vdd 0.0083f
C4567 _131_ _070_ 0.161861f
C4568 result[7] _420_/a_2248_156# 0.034866f
C4569 FILLER_0_7_104/a_932_472# _058_ 0.002096f
C4570 _052_ net36 0.005689f
C4571 _144_ mask\[6\] 0.230129f
C4572 _144_ mask\[8\] 0.131592f
C4573 FILLER_0_19_171/a_36_472# _434_/a_36_151# 0.00271f
C4574 _052_ FILLER_0_18_37/a_932_472# 0.002749f
C4575 fanout75/a_36_113# _082_ 0.016843f
C4576 FILLER_0_12_50/a_36_472# _453_/a_36_151# 0.001748f
C4577 mask\[4\] _137_ 0.086066f
C4578 _114_ _267_/a_224_472# 0.001264f
C4579 _430_/a_796_472# mask\[2\] 0.006305f
C4580 state\[2\] net74 0.024462f
C4581 _346_/a_49_472# _145_ 0.001141f
C4582 mask\[2\] FILLER_0_15_235/a_484_472# 0.004683f
C4583 _053_ _161_ 0.001047f
C4584 vss net6 0.096009f
C4585 FILLER_0_9_28/a_1916_375# _042_ 0.002352f
C4586 _132_ net36 0.029615f
C4587 net45 output17/a_224_472# 0.01994f
C4588 FILLER_0_17_200/a_572_375# net21 0.011557f
C4589 fanout82/a_36_113# _425_/a_36_151# 0.030783f
C4590 _415_/a_2665_112# _416_/a_36_151# 0.001602f
C4591 FILLER_0_23_88/a_124_375# _437_/a_36_151# 0.002709f
C4592 FILLER_0_22_177/a_1380_472# mask\[6\] 0.006573f
C4593 net35 FILLER_0_22_177/a_932_472# 0.00643f
C4594 _098_ _048_ 0.092201f
C4595 mask\[9\] FILLER_0_18_76/a_484_472# 0.002672f
C4596 FILLER_0_9_28/a_1020_375# net16 0.012909f
C4597 ctlp[1] FILLER_0_23_282/a_124_375# 0.00324f
C4598 ctln[8] ctln[9] 0.003265f
C4599 net15 _043_ 0.042278f
C4600 result[9] _421_/a_448_472# 0.015264f
C4601 output32/a_224_472# _008_ 0.074809f
C4602 FILLER_0_14_181/a_124_375# vdd 0.040138f
C4603 _053_ _129_ 0.003479f
C4604 net57 FILLER_0_13_142/a_572_375# 0.011369f
C4605 _172_ vss 0.054608f
C4606 net34 FILLER_0_22_128/a_2364_375# 0.009656f
C4607 net55 _131_ 0.314732f
C4608 net54 _026_ 0.006401f
C4609 cal_itt\[3\] _072_ 2.019868f
C4610 _292_/a_36_160# _047_ 0.001291f
C4611 _205_/a_36_160# _048_ 0.040317f
C4612 net73 _438_/a_2665_112# 0.001708f
C4613 net48 vss 0.161385f
C4614 net75 FILLER_0_8_247/a_1380_472# 0.020589f
C4615 net20 net78 1.100401f
C4616 _140_ FILLER_0_22_128/a_2276_472# 0.002954f
C4617 _430_/a_36_151# net22 0.005321f
C4618 mask\[5\] _434_/a_2665_112# 0.003849f
C4619 _119_ FILLER_0_4_107/a_1468_375# 0.001695f
C4620 _188_ _067_ 0.001554f
C4621 _383_/a_36_472# vdd -0.002154f
C4622 result[7] _419_/a_2665_112# 0.002471f
C4623 _219_/a_36_160# _439_/a_2665_112# 0.002537f
C4624 FILLER_0_8_247/a_1468_375# vdd 0.011086f
C4625 _085_ _267_/a_672_472# 0.006682f
C4626 _116_ _267_/a_1568_472# 0.001147f
C4627 _421_/a_2665_112# net33 0.007127f
C4628 mask\[4\] _276_/a_36_160# 0.025336f
C4629 net81 _425_/a_1308_423# 0.004202f
C4630 net55 FILLER_0_18_37/a_572_375# 0.007169f
C4631 net72 FILLER_0_18_37/a_36_472# 0.043427f
C4632 mask\[0\] mask\[1\] 0.01742f
C4633 net76 FILLER_0_5_212/a_36_472# 0.00377f
C4634 net15 net68 0.205016f
C4635 _187_ _188_ 0.001453f
C4636 net47 _221_/a_36_160# 0.012197f
C4637 _093_ FILLER_0_18_209/a_484_472# 0.014737f
C4638 _415_/a_36_151# result[1] 0.012965f
C4639 _104_ _420_/a_2665_112# 0.053555f
C4640 _441_/a_1308_423# _164_ 0.001807f
C4641 state\[1\] FILLER_0_13_142/a_1380_472# 0.006475f
C4642 FILLER_0_17_200/a_36_472# FILLER_0_18_177/a_2724_472# 0.026657f
C4643 FILLER_0_3_221/a_124_375# net59 0.008996f
C4644 _058_ net14 0.40635f
C4645 net32 net22 0.042885f
C4646 FILLER_0_4_99/a_124_375# FILLER_0_4_91/a_572_375# 0.012001f
C4647 FILLER_0_10_78/a_484_472# FILLER_0_9_72/a_1020_375# 0.001543f
C4648 FILLER_0_10_28/a_36_472# net47 0.002783f
C4649 output33/a_224_472# net33 0.151281f
C4650 _013_ _424_/a_2665_112# 0.001222f
C4651 net38 _450_/a_36_151# 0.035458f
C4652 _420_/a_2560_156# vdd 0.001652f
C4653 _011_ _422_/a_36_151# 0.015698f
C4654 _420_/a_2665_112# vss 0.001749f
C4655 _086_ _395_/a_36_488# 0.00825f
C4656 FILLER_0_12_136/a_124_375# state\[2\] 0.001029f
C4657 FILLER_0_12_136/a_1020_375# net53 0.002709f
C4658 FILLER_0_7_72/a_1916_375# vss 0.001259f
C4659 FILLER_0_16_241/a_124_375# net36 0.004069f
C4660 _018_ FILLER_0_15_205/a_36_472# 0.00273f
C4661 _308_/a_848_380# _115_ 0.00763f
C4662 output26/a_224_472# FILLER_0_23_44/a_484_472# 0.0323f
C4663 _399_/a_224_472# _182_ 0.002729f
C4664 vss FILLER_0_16_115/a_36_472# 0.003243f
C4665 _098_ FILLER_0_15_180/a_36_472# 0.101593f
C4666 cal_count\[1\] _451_/a_2225_156# 0.006336f
C4667 _444_/a_2248_156# net67 0.028782f
C4668 result[1] net64 0.048458f
C4669 FILLER_0_4_197/a_124_375# net21 0.018398f
C4670 net52 _443_/a_2248_156# 0.045316f
C4671 FILLER_0_2_93/a_572_375# _367_/a_36_68# 0.001069f
C4672 mask\[9\] FILLER_0_20_107/a_36_472# 0.006047f
C4673 net31 _093_ 0.274432f
C4674 output14/a_224_472# _442_/a_36_151# 0.172111f
C4675 net58 net18 0.091503f
C4676 FILLER_0_16_57/a_1020_375# vdd 0.004428f
C4677 FILLER_0_16_57/a_572_375# vss 0.00372f
C4678 vdd _450_/a_2449_156# 0.003646f
C4679 FILLER_0_16_37/a_36_472# _402_/a_728_93# 0.0108f
C4680 _387_/a_36_113# _170_ 0.017801f
C4681 net35 _436_/a_1000_472# 0.009213f
C4682 FILLER_0_4_123/a_124_375# _070_ 0.001677f
C4683 net55 FILLER_0_13_80/a_36_472# 0.016536f
C4684 _062_ _134_ 0.024038f
C4685 _322_/a_1152_472# _068_ 0.001502f
C4686 _430_/a_448_472# net63 0.026599f
C4687 _265_/a_244_68# _001_ 0.008874f
C4688 _183_ vss 0.009822f
C4689 _374_/a_244_472# _076_ 0.001567f
C4690 FILLER_0_15_212/a_1020_375# vss 0.035883f
C4691 FILLER_0_15_212/a_1468_375# vdd 0.010445f
C4692 FILLER_0_15_212/a_124_375# mask\[1\] 0.007876f
C4693 ctln[6] vss 0.45431f
C4694 net68 net51 0.008885f
C4695 _099_ mask\[1\] 0.19135f
C4696 _063_ trim_mask\[1\] 0.127216f
C4697 _316_/a_1084_68# net37 0.001574f
C4698 FILLER_0_16_89/a_36_472# _176_ 0.012173f
C4699 FILLER_0_18_2/a_2724_472# vdd 0.004348f
C4700 net16 _233_/a_36_160# 0.01152f
C4701 trimb[1] vdd 0.225206f
C4702 FILLER_0_20_177/a_932_472# _434_/a_36_151# 0.001723f
C4703 ctln[4] ctln[3] 0.073214f
C4704 FILLER_0_16_154/a_1380_472# vdd 0.001901f
C4705 FILLER_0_16_154/a_932_472# vss 0.001652f
C4706 FILLER_0_4_177/a_124_375# _386_/a_848_380# 0.001277f
C4707 _065_ _447_/a_448_472# 0.049072f
C4708 FILLER_0_17_200/a_124_375# net22 0.003602f
C4709 net57 _386_/a_848_380# 0.041622f
C4710 net15 net67 0.109181f
C4711 net64 FILLER_0_12_236/a_484_472# 0.010321f
C4712 fanout68/a_36_113# net17 0.001252f
C4713 trim_mask\[1\] FILLER_0_6_47/a_1468_375# 0.007169f
C4714 _142_ net53 0.001961f
C4715 FILLER_0_19_111/a_484_472# vdd 0.009246f
C4716 trimb[1] FILLER_0_20_15/a_484_472# 0.001292f
C4717 net62 FILLER_0_15_282/a_124_375# 0.012711f
C4718 _434_/a_36_151# vss 0.006401f
C4719 _434_/a_448_472# vdd 0.020387f
C4720 _148_ _352_/a_49_472# 0.003082f
C4721 fanout80/a_36_113# vss 0.003526f
C4722 mask\[5\] FILLER_0_20_193/a_572_375# 0.036451f
C4723 _144_ _433_/a_2248_156# 0.021805f
C4724 FILLER_0_8_107/a_124_375# _070_ 0.003069f
C4725 trimb[2] trimb[3] 0.369908f
C4726 _074_ _070_ 0.102481f
C4727 _430_/a_36_151# vdd 0.112575f
C4728 _163_ _385_/a_36_68# 0.012699f
C4729 net76 net2 0.039533f
C4730 FILLER_0_15_59/a_572_375# vss 0.018573f
C4731 FILLER_0_15_59/a_36_472# vdd 0.031071f
C4732 ctln[2] net59 0.009218f
C4733 net15 FILLER_0_11_64/a_36_472# 0.020589f
C4734 _080_ net37 0.005467f
C4735 _053_ _220_/a_255_603# 0.001311f
C4736 _430_/a_448_472# _069_ 0.047845f
C4737 FILLER_0_19_47/a_484_472# net55 0.061087f
C4738 FILLER_0_11_101/a_124_375# _070_ 0.052406f
C4739 _270_/a_36_472# net21 0.001606f
C4740 _260_/a_36_68# FILLER_0_3_221/a_1380_472# 0.001652f
C4741 FILLER_0_12_136/a_1380_472# _127_ 0.001432f
C4742 output8/a_224_472# FILLER_0_3_221/a_572_375# 0.03228f
C4743 _070_ _076_ 0.198272f
C4744 mask\[7\] FILLER_0_22_177/a_1468_375# 0.001315f
C4745 ctln[1] net58 0.014147f
C4746 fanout69/a_36_113# vss 0.002239f
C4747 _028_ FILLER_0_7_72/a_572_375# 0.003837f
C4748 net35 FILLER_0_22_128/a_124_375# 0.010439f
C4749 trim_val\[4\] FILLER_0_3_172/a_36_472# 0.006208f
C4750 net76 FILLER_0_3_172/a_2276_472# 0.002531f
C4751 _053_ FILLER_0_7_59/a_484_472# 0.013665f
C4752 _162_ _312_/a_234_472# 0.003812f
C4753 FILLER_0_4_152/a_36_472# vss 0.009467f
C4754 FILLER_0_7_146/a_36_472# _076_ 0.001843f
C4755 FILLER_0_7_146/a_124_375# _068_ 0.033245f
C4756 output8/a_224_472# _000_ 0.182377f
C4757 net50 trim_mask\[1\] 0.502622f
C4758 FILLER_0_9_28/a_124_375# FILLER_0_8_24/a_572_375# 0.05841f
C4759 _432_/a_36_151# FILLER_0_15_180/a_36_472# 0.002018f
C4760 FILLER_0_22_128/a_2724_472# FILLER_0_21_150/a_124_375# 0.001543f
C4761 net75 _253_/a_1100_68# 0.001047f
C4762 output45/a_224_472# net43 0.024629f
C4763 _064_ _445_/a_1308_423# 0.01485f
C4764 net52 _176_ 0.004215f
C4765 FILLER_0_13_212/a_932_472# net79 0.006824f
C4766 FILLER_0_16_107/a_484_472# _451_/a_36_151# 0.027244f
C4767 net62 FILLER_0_13_212/a_1380_472# 0.059367f
C4768 net32 vdd 0.50705f
C4769 _140_ net71 0.005182f
C4770 _069_ FILLER_0_11_142/a_484_472# 0.005789f
C4771 _132_ FILLER_0_16_107/a_572_375# 0.007439f
C4772 net39 net67 0.049482f
C4773 mask\[5\] FILLER_0_18_177/a_1468_375# 0.002726f
C4774 net4 FILLER_0_3_221/a_1380_472# 0.003953f
C4775 FILLER_0_13_206/a_36_472# net22 0.053292f
C4776 net16 net49 0.055931f
C4777 ctlp[6] net54 0.00409f
C4778 net67 net51 0.010753f
C4779 ctlp[3] _009_ 0.018168f
C4780 FILLER_0_15_205/a_36_472# vss 0.003239f
C4781 FILLER_0_15_116/a_572_375# _131_ 0.051323f
C4782 _450_/a_448_472# clkc 0.003011f
C4783 _450_/a_1040_527# net6 0.019715f
C4784 _189_/a_67_603# _043_ 0.005635f
C4785 FILLER_0_12_124/a_36_472# cal_count\[3\] 0.004109f
C4786 _084_ _316_/a_124_24# 0.001501f
C4787 _372_/a_170_472# vdd 0.031606f
C4788 _181_ _180_ 0.216908f
C4789 ctlp[9] vss 0.013018f
C4790 output34/a_224_472# _099_ 0.001498f
C4791 net75 _015_ 0.025217f
C4792 FILLER_0_12_220/a_484_472# vdd 0.002383f
C4793 FILLER_0_12_220/a_36_472# vss 0.023702f
C4794 _053_ _068_ 0.066662f
C4795 FILLER_0_11_64/a_36_472# net51 0.009015f
C4796 net50 _447_/a_2665_112# 0.015374f
C4797 net10 vss 0.324553f
C4798 _115_ net14 0.037635f
C4799 _058_ FILLER_0_8_156/a_124_375# 0.006325f
C4800 _091_ FILLER_0_18_209/a_572_375# 0.001343f
C4801 ctln[1] net82 0.001141f
C4802 output35/a_224_472# _048_ 0.009509f
C4803 _087_ net22 0.028009f
C4804 net74 _125_ 0.071757f
C4805 FILLER_0_7_162/a_36_472# FILLER_0_8_156/a_572_375# 0.001543f
C4806 state\[0\] _128_ 0.228492f
C4807 _186_ _067_ 0.001907f
C4808 _074_ FILLER_0_5_164/a_572_375# 0.001307f
C4809 _323_/a_36_113# vdd 0.009958f
C4810 net78 _009_ 0.02395f
C4811 net39 _445_/a_448_472# 0.014537f
C4812 _093_ FILLER_0_18_107/a_3172_472# 0.008787f
C4813 FILLER_0_5_72/a_36_472# _029_ 0.007282f
C4814 FILLER_0_5_72/a_572_375# trim_mask\[1\] 0.010714f
C4815 FILLER_0_22_177/a_484_472# vss -0.001894f
C4816 FILLER_0_22_177/a_932_472# vdd 0.029547f
C4817 valid net76 0.285892f
C4818 _411_/a_2248_156# net19 0.001197f
C4819 net58 _074_ 0.004651f
C4820 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3260_375# 0.086905f
C4821 _426_/a_2665_112# net64 0.01548f
C4822 output34/a_224_472# _419_/a_2248_156# 0.022045f
C4823 _046_ net30 0.006105f
C4824 mask\[2\] FILLER_0_16_154/a_1468_375# 0.014254f
C4825 FILLER_0_4_107/a_484_472# _160_ 0.008194f
C4826 _079_ net1 0.099822f
C4827 _063_ _444_/a_2665_112# 0.001996f
C4828 _452_/a_36_151# net40 0.012138f
C4829 FILLER_0_4_213/a_484_472# vdd 0.007084f
C4830 FILLER_0_4_213/a_36_472# vss 0.003969f
C4831 _070_ FILLER_0_5_164/a_484_472# 0.003424f
C4832 _187_ _186_ 0.032149f
C4833 FILLER_0_17_200/a_124_375# vdd -0.010938f
C4834 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_36_472# 0.009654f
C4835 FILLER_0_5_109/a_484_472# vdd 0.007355f
C4836 _128_ _247_/a_36_160# 0.00163f
C4837 FILLER_0_17_72/a_1916_375# _131_ 0.006589f
C4838 _277_/a_36_160# _093_ 0.018101f
C4839 net55 FILLER_0_13_72/a_124_375# 0.00281f
C4840 _449_/a_2248_156# vdd -0.001225f
C4841 _449_/a_1204_472# vss 0.006048f
C4842 cal_count\[2\] net47 0.274891f
C4843 net26 _423_/a_36_151# 0.067024f
C4844 net53 FILLER_0_14_123/a_124_375# 0.003138f
C4845 result[6] _421_/a_1204_472# 0.005361f
C4846 _103_ _007_ 0.002514f
C4847 _086_ net22 0.00117f
C4848 _003_ vss 0.095366f
C4849 net82 _170_ 0.080348f
C4850 net28 _044_ 0.481924f
C4851 mask\[0\] _099_ 0.00418f
C4852 _411_/a_448_472# _000_ 0.073053f
C4853 fanout64/a_36_160# net65 0.214347f
C4854 _308_/a_848_380# _134_ 0.001299f
C4855 _149_ _437_/a_2665_112# 0.020763f
C4856 _026_ _437_/a_1204_472# 0.022954f
C4857 FILLER_0_1_266/a_124_375# FILLER_0_0_266/a_124_375# 0.05841f
C4858 _074_ _082_ 0.069835f
C4859 vss trim[3] 0.235724f
C4860 _070_ _081_ 0.00804f
C4861 _451_/a_836_156# _040_ 0.016371f
C4862 _074_ net82 0.123449f
C4863 _442_/a_36_151# vdd 0.102701f
C4864 FILLER_0_14_181/a_36_472# _043_ 0.008613f
C4865 net15 FILLER_0_6_47/a_1916_375# 0.029774f
C4866 _176_ FILLER_0_15_72/a_572_375# 0.005529f
C4867 net38 _445_/a_36_151# 0.112205f
C4868 net50 _444_/a_2665_112# 0.023342f
C4869 net25 _423_/a_2248_156# 0.005535f
C4870 _073_ FILLER_0_6_231/a_36_472# 0.001898f
C4871 _086_ _311_/a_2700_473# 0.00176f
C4872 net47 _450_/a_448_472# 0.012172f
C4873 _305_/a_36_159# vdd 0.017293f
C4874 net81 net59 0.074175f
C4875 fanout62/a_36_160# FILLER_0_11_282/a_36_472# 0.005262f
C4876 mask\[4\] FILLER_0_19_171/a_484_472# 0.004669f
C4877 FILLER_0_19_47/a_124_375# _013_ 0.023766f
C4878 net1 cal_itt\[1\] 0.229522f
C4879 _408_/a_56_524# _185_ 0.002484f
C4880 net73 vdd 0.44835f
C4881 FILLER_0_13_206/a_36_472# vdd 0.011681f
C4882 FILLER_0_19_155/a_572_375# vdd 0.01384f
C4883 FILLER_0_19_155/a_124_375# vss 0.00336f
C4884 FILLER_0_13_206/a_124_375# vss 0.051723f
C4885 sample vss 0.276162f
C4886 _137_ FILLER_0_15_180/a_484_472# 0.046411f
C4887 FILLER_0_7_104/a_932_472# _134_ 0.004249f
C4888 net37 vss 0.666835f
C4889 ctln[2] FILLER_0_1_266/a_124_375# 0.047145f
C4890 net18 FILLER_0_9_270/a_484_472# 0.004375f
C4891 _445_/a_2560_156# vdd 0.002586f
C4892 _445_/a_2665_112# vss 0.004455f
C4893 FILLER_0_21_28/a_3172_472# vss 0.001574f
C4894 _436_/a_1000_472# vdd 0.006522f
C4895 FILLER_0_3_221/a_36_472# vdd 0.018263f
C4896 FILLER_0_3_221/a_1468_375# vss 0.004085f
C4897 _105_ mask\[5\] 0.706158f
C4898 _423_/a_2665_112# _012_ 0.014394f
C4899 net73 FILLER_0_18_107/a_572_375# 0.008889f
C4900 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_484_472# 0.001963f
C4901 _413_/a_2560_156# net59 0.016463f
C4902 _303_/a_36_472# net36 0.006675f
C4903 net76 FILLER_0_5_172/a_124_375# 0.001526f
C4904 net36 _438_/a_1204_472# 0.012234f
C4905 _053_ _152_ 0.032961f
C4906 _256_/a_36_68# calibrate 0.02084f
C4907 _439_/a_796_472# vss 0.003859f
C4908 _149_ net14 0.102004f
C4909 net62 _429_/a_2248_156# 0.012262f
C4910 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_36_472# 0.086743f
C4911 FILLER_0_18_171/a_36_472# FILLER_0_18_177/a_36_472# 0.003468f
C4912 _087_ vdd 0.281159f
C4913 net20 _418_/a_2248_156# 0.003507f
C4914 _075_ net37 0.001054f
C4915 net15 _424_/a_2248_156# 0.00415f
C4916 _189_/a_67_603# FILLER_0_12_236/a_124_375# 0.00221f
C4917 _445_/a_36_151# net66 0.058093f
C4918 _415_/a_36_151# net81 0.046145f
C4919 mask\[3\] net22 0.036607f
C4920 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_36_472# 0.001963f
C4921 net79 _193_/a_36_160# 0.010228f
C4922 FILLER_0_13_212/a_36_472# net22 0.002402f
C4923 FILLER_0_14_99/a_36_472# vdd 0.095251f
C4924 FILLER_0_14_99/a_124_375# vss 0.017196f
C4925 FILLER_0_12_136/a_1468_375# cal_count\[3\] 0.004337f
C4926 _043_ net47 0.043824f
C4927 output31/a_224_472# FILLER_0_17_282/a_36_472# 0.008834f
C4928 net44 FILLER_0_12_2/a_124_375# 0.01836f
C4929 net50 FILLER_0_6_90/a_36_472# 0.049285f
C4930 FILLER_0_12_2/a_572_375# vss 0.017629f
C4931 FILLER_0_12_2/a_36_472# vdd 0.104425f
C4932 _122_ _160_ 0.004488f
C4933 net63 _434_/a_448_472# 0.008139f
C4934 _074_ _312_/a_234_472# 0.005755f
C4935 _162_ calibrate 0.228839f
C4936 net81 FILLER_0_10_256/a_36_472# 0.089055f
C4937 FILLER_0_16_57/a_1380_472# _176_ 0.01346f
C4938 FILLER_0_10_37/a_124_375# vdd 0.048346f
C4939 _077_ _067_ 0.090648f
C4940 _016_ _127_ 0.01898f
C4941 FILLER_0_8_127/a_124_375# vdd 0.019587f
C4942 result[7] _421_/a_1204_472# 0.014927f
C4943 _430_/a_36_151# net63 0.026607f
C4944 net81 net64 0.455159f
C4945 _448_/a_36_151# _037_ 0.012725f
C4946 _120_ FILLER_0_10_107/a_124_375# 0.001834f
C4947 _086_ vdd 1.212255f
C4948 net67 clkc 0.102244f
C4949 FILLER_0_22_128/a_124_375# vdd 0.013058f
C4950 _217_/a_36_160# FILLER_0_19_28/a_572_375# 0.058908f
C4951 _058_ _439_/a_2665_112# 0.001029f
C4952 net75 _084_ 0.045583f
C4953 output46/a_224_472# FILLER_0_21_28/a_124_375# 0.003337f
C4954 output34/a_224_472# output18/a_224_472# 0.002121f
C4955 _139_ vss 0.052996f
C4956 mask\[5\] output19/a_224_472# 0.092961f
C4957 _077_ _187_ 0.058967f
C4958 net58 net65 1.468105f
C4959 valid fanout65/a_36_113# 0.001646f
C4960 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1468_375# 0.086635f
C4961 net68 net47 0.063835f
C4962 _098_ _145_ 0.007514f
C4963 net69 FILLER_0_3_78/a_36_472# 0.002068f
C4964 FILLER_0_9_142/a_124_375# _120_ 0.04442f
C4965 net60 _418_/a_2665_112# 0.042307f
C4966 net69 FILLER_0_2_127/a_36_472# 0.019383f
C4967 _072_ _306_/a_36_68# 0.042843f
C4968 state\[1\] _097_ 0.004171f
C4969 _134_ net14 0.001303f
C4970 net41 _408_/a_728_93# 0.058816f
C4971 _081_ _082_ 0.008298f
C4972 net64 _223_/a_36_160# 0.007842f
C4973 _070_ _090_ 0.369847f
C4974 FILLER_0_0_130/a_124_375# net13 0.009149f
C4975 FILLER_0_4_197/a_1020_375# net22 0.040565f
C4976 _397_/a_36_472# FILLER_0_17_72/a_1020_375# 0.001781f
C4977 net62 _248_/a_36_68# 0.002178f
C4978 trim_val\[2\] _160_ 0.051804f
C4979 net54 FILLER_0_21_150/a_124_375# 0.007123f
C4980 ctlp[5] vss 0.032166f
C4981 _430_/a_36_151# _069_ 0.026308f
C4982 _065_ _441_/a_2665_112# 0.003318f
C4983 result[0] FILLER_0_9_282/a_484_472# 0.018647f
C4984 _132_ _114_ 0.08562f
C4985 net62 _417_/a_2665_112# 0.006083f
C4986 net47 _156_ 0.040298f
C4987 calibrate net18 0.014127f
C4988 net74 _043_ 0.65119f
C4989 FILLER_0_9_282/a_36_472# vdd 0.106034f
C4990 FILLER_0_9_282/a_572_375# vss 0.058599f
C4991 _137_ _138_ 0.045916f
C4992 FILLER_0_6_47/a_1380_472# vdd 0.002735f
C4993 _429_/a_36_151# net21 0.054289f
C4994 _013_ _182_ 0.001681f
C4995 net82 net65 0.630327f
C4996 _053_ _377_/a_36_472# 0.023504f
C4997 mask\[4\] FILLER_0_20_177/a_1380_472# 0.001215f
C4998 result[8] FILLER_0_24_290/a_124_375# 0.00562f
C4999 mask\[8\] FILLER_0_22_107/a_484_472# 0.024416f
C5000 net35 FILLER_0_22_107/a_36_472# 0.007196f
C5001 FILLER_0_10_78/a_484_472# _176_ 0.001731f
C5002 net56 fanout54/a_36_160# 0.044466f
C5003 net16 _052_ 0.022236f
C5004 _193_/a_36_160# FILLER_0_13_290/a_124_375# 0.005732f
C5005 fanout57/a_36_113# net65 0.035361f
C5006 net63 FILLER_0_22_177/a_932_472# 0.060639f
C5007 output36/a_224_472# result[9] 0.059164f
C5008 _322_/a_692_472# _118_ 0.002849f
C5009 mask\[3\] vdd 0.340612f
C5010 FILLER_0_13_212/a_1468_375# vss 0.062822f
C5011 FILLER_0_13_212/a_36_472# vdd 0.105926f
C5012 FILLER_0_9_223/a_124_375# net4 0.061757f
C5013 FILLER_0_4_185/a_36_472# net76 0.023698f
C5014 FILLER_0_12_136/a_36_472# _114_ 0.003953f
C5015 FILLER_0_17_200/a_124_375# net63 0.008905f
C5016 state\[0\] _274_/a_36_68# 0.001852f
C5017 ctlp[1] _420_/a_448_472# 0.038053f
C5018 net67 net47 0.126281f
C5019 _086_ _135_ 0.005637f
C5020 cal_count\[3\] FILLER_0_12_28/a_124_375# 0.013328f
C5021 _421_/a_2665_112# vdd 0.029293f
C5022 FILLER_0_20_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001543f
C5023 _446_/a_1000_472# net17 0.031119f
C5024 net19 cal_itt\[0\] 0.111163f
C5025 _072_ _395_/a_36_488# 0.024944f
C5026 net62 _005_ 0.097739f
C5027 result[8] FILLER_0_24_274/a_1380_472# 0.005458f
C5028 FILLER_0_19_187/a_572_375# vss 0.055266f
C5029 FILLER_0_19_187/a_36_472# vdd 0.09884f
C5030 _413_/a_36_151# FILLER_0_3_172/a_2724_472# 0.001723f
C5031 vss FILLER_0_21_60/a_484_472# 0.004134f
C5032 ctln[4] FILLER_0_1_212/a_124_375# 0.008197f
C5033 FILLER_0_9_28/a_2724_472# _077_ 0.006001f
C5034 mask\[5\] mask\[6\] 0.140269f
C5035 _094_ FILLER_0_17_282/a_124_375# 0.001151f
C5036 FILLER_0_2_111/a_1468_375# vdd 0.011806f
C5037 _429_/a_796_472# net22 0.020124f
C5038 _093_ FILLER_0_17_104/a_932_472# 0.014431f
C5039 net41 FILLER_0_16_37/a_36_472# 0.009425f
C5040 trim_mask\[2\] fanout68/a_36_113# 0.003509f
C5041 FILLER_0_4_91/a_572_375# _160_ 0.007391f
C5042 net15 _394_/a_728_93# 0.085551f
C5043 output33/a_224_472# vdd -0.031734f
C5044 net50 net66 0.016385f
C5045 net52 _030_ 0.035783f
C5046 FILLER_0_11_109/a_36_472# _134_ 0.007739f
C5047 _445_/a_448_472# net47 0.005429f
C5048 _149_ _148_ 0.001124f
C5049 _440_/a_1308_423# vss 0.028595f
C5050 _415_/a_1000_472# result[1] 0.005365f
C5051 _021_ _143_ 0.007778f
C5052 net66 _382_/a_224_472# 0.001902f
C5053 _379_/a_36_472# _164_ 0.026812f
C5054 net18 _418_/a_448_472# 0.026048f
C5055 _077_ net23 0.0245f
C5056 output26/a_224_472# ctlp[9] 0.034572f
C5057 _006_ net30 0.284414f
C5058 _030_ net49 0.046089f
C5059 _430_/a_2248_156# net36 0.001198f
C5060 clk net18 0.003519f
C5061 _313_/a_67_603# vdd -0.002183f
C5062 _132_ _124_ 0.005668f
C5063 _390_/a_36_68# vss 0.002334f
C5064 output25/a_224_472# _051_ 0.019651f
C5065 net82 _443_/a_448_472# 0.007335f
C5066 FILLER_0_4_197/a_1020_375# vdd 0.002455f
C5067 _115_ _439_/a_2665_112# 0.003617f
C5068 net34 _108_ 0.297364f
C5069 net44 FILLER_0_20_2/a_124_375# 0.001564f
C5070 net70 FILLER_0_14_107/a_1020_375# 0.011157f
C5071 FILLER_0_20_2/a_572_375# vss 0.001471f
C5072 FILLER_0_20_2/a_36_472# vdd 0.102471f
C5073 _079_ net76 2.404004f
C5074 fanout62/a_36_160# vdd 0.059299f
C5075 _103_ net30 0.013544f
C5076 output8/a_224_472# ctln[1] 0.020259f
C5077 FILLER_0_5_54/a_484_472# trim_mask\[1\] 0.013584f
C5078 FILLER_0_4_197/a_1380_472# _088_ 0.017451f
C5079 _057_ _060_ 0.033334f
C5080 net34 net19 0.039959f
C5081 _438_/a_36_151# vdd 0.111691f
C5082 _343_/a_665_69# _141_ 0.002451f
C5083 ctlp[1] _419_/a_1308_423# 0.00678f
C5084 net25 net24 0.031854f
C5085 _405_/a_67_603# net40 0.015326f
C5086 _132_ fanout71/a_36_113# 0.055078f
C5087 _451_/a_3129_107# vdd 0.008569f
C5088 _137_ _113_ 0.030279f
C5089 _062_ FILLER_0_8_156/a_484_472# 0.006123f
C5090 FILLER_0_5_198/a_36_472# net37 0.0114f
C5091 _369_/a_244_472# _160_ 0.00146f
C5092 mask\[5\] FILLER_0_19_171/a_1020_375# 0.007169f
C5093 result[4] _418_/a_36_151# 0.005556f
C5094 _074_ calibrate 0.046632f
C5095 net41 FILLER_0_23_44/a_36_472# 0.001116f
C5096 output7/a_224_472# net17 0.001164f
C5097 _370_/a_848_380# FILLER_0_5_136/a_124_375# 0.014613f
C5098 net4 _248_/a_36_68# 0.054512f
C5099 net50 FILLER_0_3_54/a_124_375# 0.00189f
C5100 _442_/a_2665_112# _157_ 0.001587f
C5101 FILLER_0_4_144/a_124_375# _059_ 0.031451f
C5102 _079_ FILLER_0_5_198/a_124_375# 0.013896f
C5103 _095_ _402_/a_718_527# 0.002109f
C5104 _033_ FILLER_0_6_37/a_36_472# 0.017695f
C5105 _236_/a_36_160# vdd 0.023428f
C5106 _164_ FILLER_0_6_47/a_1020_375# 0.004285f
C5107 _076_ calibrate 1.005804f
C5108 _069_ FILLER_0_13_206/a_36_472# 0.005793f
C5109 _430_/a_2665_112# mask\[3\] 0.002697f
C5110 _074_ net21 0.186175f
C5111 _447_/a_448_472# net69 0.001694f
C5112 net16 _165_ 0.021744f
C5113 _070_ FILLER_0_7_233/a_36_472# 0.07194f
C5114 ctln[1] clk 0.551557f
C5115 _073_ _078_ 0.098575f
C5116 _028_ FILLER_0_5_72/a_1020_375# 0.00123f
C5117 _154_ _156_ 0.019471f
C5118 _408_/a_56_524# net17 0.048018f
C5119 _177_ _150_ 0.002507f
C5120 net76 cal_itt\[1\] 0.027781f
C5121 _414_/a_36_151# _074_ 0.070632f
C5122 net45 net43 0.131763f
C5123 _418_/a_1308_423# _417_/a_36_151# 0.001518f
C5124 _417_/a_36_151# _006_ 0.015561f
C5125 FILLER_0_7_104/a_124_375# _131_ 0.001291f
C5126 _057_ _116_ 0.028033f
C5127 _076_ net21 0.031683f
C5128 _052_ FILLER_0_21_28/a_2364_375# 0.002388f
C5129 _093_ FILLER_0_18_177/a_2364_375# 0.001989f
C5130 _070_ _163_ 1.884485f
C5131 FILLER_0_18_37/a_1468_375# vss 0.054381f
C5132 FILLER_0_18_37/a_36_472# vdd 0.136723f
C5133 FILLER_0_9_28/a_932_472# net68 0.003603f
C5134 _061_ net22 0.123662f
C5135 net75 _316_/a_848_380# 0.044673f
C5136 _333_/a_36_160# FILLER_0_15_180/a_36_472# 0.016014f
C5137 net27 FILLER_0_11_282/a_124_375# 0.002857f
C5138 _429_/a_36_151# mask\[1\] 0.001021f
C5139 _429_/a_1308_423# vss 0.008906f
C5140 net52 trim_mask\[3\] 0.666362f
C5141 FILLER_0_16_73/a_36_472# vss 0.035175f
C5142 _317_/a_36_113# FILLER_0_7_233/a_124_375# 0.03227f
C5143 _331_/a_448_472# _120_ 0.001496f
C5144 cal_count\[3\] _136_ 0.00703f
C5145 net73 FILLER_0_18_139/a_36_472# 0.002491f
C5146 net8 vss 0.171128f
C5147 net79 _416_/a_36_151# 0.062626f
C5148 net62 _416_/a_448_472# 0.009111f
C5149 _044_ output30/a_224_472# 0.00717f
C5150 net49 trim_mask\[3\] 0.03723f
C5151 FILLER_0_5_72/a_1380_472# FILLER_0_5_88/a_36_472# 0.013277f
C5152 ctln[1] _411_/a_448_472# 0.039538f
C5153 FILLER_0_21_142/a_484_472# vss 0.034607f
C5154 _196_/a_36_160# mask\[1\] 0.003254f
C5155 FILLER_0_14_99/a_124_375# _095_ 0.012128f
C5156 ctln[5] _448_/a_796_472# 0.001484f
C5157 FILLER_0_3_2/a_36_472# net66 0.011419f
C5158 _414_/a_448_472# _074_ 0.008725f
C5159 _057_ _118_ 0.055726f
C5160 net38 _039_ 0.059899f
C5161 net16 net40 0.039189f
C5162 trimb[4] vdd 0.081023f
C5163 _147_ _434_/a_36_151# 0.001817f
C5164 result[8] FILLER_0_23_282/a_36_472# 0.001908f
C5165 _086_ _069_ 0.580351f
C5166 output41/a_224_472# trim[3] 0.042209f
C5167 FILLER_0_15_235/a_124_375# FILLER_0_15_228/a_124_375# 0.002868f
C5168 output21/a_224_472# mask\[5\] 0.009585f
C5169 net52 net13 0.018118f
C5170 _122_ FILLER_0_5_164/a_36_472# 0.002232f
C5171 _310_/a_49_472# _060_ 0.001122f
C5172 net81 mask\[2\] 0.002083f
C5173 vdd FILLER_0_22_107/a_36_472# 0.114332f
C5174 vss FILLER_0_22_107/a_572_375# 0.001944f
C5175 _423_/a_36_151# FILLER_0_23_60/a_36_472# 0.001723f
C5176 FILLER_0_19_55/a_124_375# _052_ 0.053626f
C5177 _181_ vss 0.003673f
C5178 _285_/a_36_472# vdd 0.073338f
C5179 output14/a_224_472# _031_ 0.001077f
C5180 _072_ net22 0.147672f
C5181 _431_/a_1000_472# vss 0.002491f
C5182 _178_ _181_ 0.188669f
C5183 _321_/a_170_472# _121_ 0.007364f
C5184 net60 _011_ 0.003094f
C5185 FILLER_0_10_37/a_36_472# net68 0.005405f
C5186 fanout49/a_36_160# FILLER_0_4_91/a_36_472# 0.001461f
C5187 net75 net4 0.031823f
C5188 net72 FILLER_0_21_28/a_1468_375# 0.001823f
C5189 net55 FILLER_0_11_78/a_124_375# 0.001597f
C5190 net16 FILLER_0_17_38/a_572_375# 0.018281f
C5191 FILLER_0_5_164/a_36_472# _169_ 0.00284f
C5192 FILLER_0_5_164/a_572_375# _163_ 0.046852f
C5193 FILLER_0_9_223/a_484_472# _076_ 0.001736f
C5194 FILLER_0_12_124/a_124_375# _428_/a_36_151# 0.058722f
C5195 _274_/a_36_68# net79 0.009814f
C5196 FILLER_0_18_2/a_2276_472# net55 0.006033f
C5197 input4/a_36_68# vdd 0.09828f
C5198 _444_/a_1000_472# net17 0.02064f
C5199 _068_ _311_/a_3740_473# 0.001409f
C5200 _070_ _117_ 0.080445f
C5201 mask\[3\] FILLER_0_16_154/a_572_375# 0.027873f
C5202 _142_ _020_ 0.010094f
C5203 net36 net19 0.031858f
C5204 FILLER_0_2_93/a_572_375# net69 0.015032f
C5205 net15 FILLER_0_5_54/a_932_472# 0.008904f
C5206 net63 mask\[3\] 0.37365f
C5207 _425_/a_796_472# calibrate 0.025807f
C5208 FILLER_0_8_24/a_484_472# net17 0.010321f
C5209 _140_ _434_/a_448_472# 0.00128f
C5210 _424_/a_2248_156# _012_ 0.009377f
C5211 _023_ vss 0.114191f
C5212 mask\[5\] FILLER_0_20_177/a_36_472# 0.017871f
C5213 _033_ _444_/a_2248_156# 0.011578f
C5214 _067_ _039_ 0.221585f
C5215 _053_ FILLER_0_6_90/a_124_375# 0.003061f
C5216 _417_/a_796_472# vss 0.001608f
C5217 result[9] result[6] 0.026511f
C5218 _024_ _435_/a_448_472# 0.039244f
C5219 FILLER_0_9_72/a_124_375# vdd -0.003896f
C5220 FILLER_0_20_98/a_36_472# vdd 0.095266f
C5221 FILLER_0_20_98/a_124_375# vss 0.013019f
C5222 _093_ _304_/a_224_472# 0.002907f
C5223 FILLER_0_10_214/a_36_472# _055_ 0.027657f
C5224 output37/a_224_472# sample 0.015298f
C5225 _081_ net21 0.030964f
C5226 net63 FILLER_0_19_187/a_36_472# 0.006753f
C5227 output34/a_224_472# net18 0.126175f
C5228 output37/a_224_472# net37 0.011407f
C5229 _255_/a_224_552# _062_ 0.009032f
C5230 _127_ vss 0.343764f
C5231 _016_ _427_/a_796_472# 0.001666f
C5232 _385_/a_36_68# net37 0.047762f
C5233 _061_ vdd 0.295557f
C5234 net35 FILLER_0_22_86/a_484_472# 0.008347f
C5235 mask\[8\] FILLER_0_22_86/a_932_472# 0.012284f
C5236 fanout66/a_36_113# vdd 0.049012f
C5237 FILLER_0_5_72/a_1020_375# net47 0.006974f
C5238 FILLER_0_21_28/a_124_375# net17 0.005751f
C5239 net65 calibrate 0.012434f
C5240 _187_ _039_ 0.228074f
C5241 FILLER_0_13_290/a_124_375# _416_/a_36_151# 0.026277f
C5242 FILLER_0_5_212/a_36_472# _078_ 0.002235f
C5243 FILLER_0_13_212/a_484_472# _043_ 0.011439f
C5244 _077_ net57 0.025864f
C5245 _414_/a_36_151# _081_ 0.016708f
C5246 _453_/a_1308_423# vdd 0.002896f
C5247 _453_/a_448_472# vss 0.00396f
C5248 _311_/a_66_473# vdd 0.106886f
C5249 net35 FILLER_0_22_128/a_3172_472# 0.014415f
C5250 net17 _452_/a_1697_156# 0.001184f
C5251 _414_/a_1308_423# net21 0.06986f
C5252 _015_ _426_/a_448_472# 0.035938f
C5253 FILLER_0_17_200/a_484_472# FILLER_0_18_177/a_3172_472# 0.026657f
C5254 FILLER_0_18_2/a_2276_472# net17 0.037088f
C5255 _053_ _042_ 0.00242f
C5256 mask\[2\] net30 0.089173f
C5257 mask\[3\] _069_ 0.025564f
C5258 net57 _267_/a_1120_472# 0.002885f
C5259 _069_ FILLER_0_13_212/a_36_472# 0.047013f
C5260 ctln[1] input2/a_36_113# 0.05197f
C5261 net82 _163_ 0.00269f
C5262 FILLER_0_12_2/a_484_472# net67 0.006435f
C5263 _141_ FILLER_0_17_161/a_124_375# 0.040332f
C5264 _397_/a_36_472# vss 0.003673f
C5265 _037_ vss 0.051886f
C5266 net68 FILLER_0_6_47/a_1828_472# 0.009096f
C5267 FILLER_0_11_135/a_36_472# vss 0.006739f
C5268 output31/a_224_472# vss -0.003316f
C5269 net65 net21 0.04444f
C5270 _001_ vdd 0.122898f
C5271 _131_ _179_ 0.034602f
C5272 net47 _380_/a_224_472# 0.001405f
C5273 _431_/a_448_472# _137_ 0.008493f
C5274 FILLER_0_18_2/a_3172_472# net41 0.00982f
C5275 FILLER_0_16_107/a_484_472# _040_ 0.003828f
C5276 _114_ FILLER_0_13_142/a_572_375# 0.00191f
C5277 net35 _050_ 0.28822f
C5278 net31 ctlp[1] 0.050993f
C5279 _189_/a_67_603# FILLER_0_13_228/a_124_375# 0.00744f
C5280 output43/a_224_472# trimb[2] 0.005445f
C5281 _098_ _437_/a_796_472# 0.0049f
C5282 ctln[5] net59 0.030363f
C5283 _412_/a_448_472# en 0.011052f
C5284 net20 FILLER_0_12_220/a_1380_472# 0.029747f
C5285 net54 FILLER_0_22_128/a_36_472# 0.020739f
C5286 output8/a_224_472# net65 0.084944f
C5287 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_36_472# 0.086635f
C5288 net32 _421_/a_448_472# 0.022214f
C5289 FILLER_0_17_72/a_1828_472# _136_ 0.004161f
C5290 _414_/a_1204_472# net21 0.007637f
C5291 net81 FILLER_0_15_212/a_572_375# 0.006974f
C5292 _077_ _439_/a_2248_156# 0.038814f
C5293 vdd _433_/a_36_151# 0.086874f
C5294 mask\[0\] _429_/a_36_151# 0.026729f
C5295 _448_/a_796_472# net59 0.004855f
C5296 ctln[5] FILLER_0_0_198/a_124_375# 0.002726f
C5297 _122_ _121_ 0.034975f
C5298 FILLER_0_21_133/a_124_375# vss 0.015693f
C5299 _101_ vdd 0.02756f
C5300 FILLER_0_11_101/a_36_472# vss 0.001641f
C5301 FILLER_0_11_101/a_484_472# vdd 0.009482f
C5302 FILLER_0_14_91/a_124_375# _177_ 0.00134f
C5303 _093_ FILLER_0_18_100/a_36_472# 0.077197f
C5304 FILLER_0_18_100/a_124_375# mask\[9\] 0.005751f
C5305 _414_/a_448_472# _081_ 0.024533f
C5306 state\[0\] _274_/a_1612_497# 0.001071f
C5307 _016_ _118_ 0.001549f
C5308 _052_ _424_/a_1308_423# 0.008633f
C5309 _238_/a_67_603# output15/a_224_472# 0.019027f
C5310 _053_ FILLER_0_5_212/a_124_375# 0.048501f
C5311 mask\[1\] FILLER_0_15_180/a_36_472# 0.001145f
C5312 _072_ vdd 0.715894f
C5313 net35 _214_/a_36_160# 0.0116f
C5314 output39/a_224_472# net17 0.041253f
C5315 FILLER_0_18_2/a_1020_375# net55 0.003942f
C5316 FILLER_0_4_107/a_572_375# _157_ 0.001032f
C5317 net76 FILLER_0_6_177/a_124_375# 0.00227f
C5318 _085_ _120_ 0.032964f
C5319 _161_ _055_ 0.078364f
C5320 _431_/a_36_151# vss 0.00849f
C5321 FILLER_0_19_195/a_124_375# vdd 0.03587f
C5322 _132_ FILLER_0_18_107/a_1380_472# 0.034976f
C5323 _411_/a_2665_112# vdd 0.026095f
C5324 _093_ FILLER_0_17_72/a_1020_375# 0.001994f
C5325 net39 _033_ 0.607942f
C5326 FILLER_0_16_73/a_124_375# _176_ 0.006386f
C5327 FILLER_0_16_107/a_36_472# net36 0.001245f
C5328 _412_/a_1000_472# vdd 0.002008f
C5329 _014_ vdd 0.035382f
C5330 _041_ net40 0.082688f
C5331 net34 _435_/a_1204_472# 0.004285f
C5332 trimb[1] net43 0.004299f
C5333 FILLER_0_7_195/a_124_375# vss 0.006314f
C5334 vss FILLER_0_13_72/a_36_472# 0.034188f
C5335 result[7] result[9] 1.21288f
C5336 net68 _440_/a_1000_472# 0.002604f
C5337 _176_ _451_/a_3081_151# 0.001255f
C5338 _345_/a_36_160# vss 0.003697f
C5339 output13/a_224_472# _170_ 0.024999f
C5340 net67 FILLER_0_6_47/a_1828_472# 0.001175f
C5341 net15 _304_/a_224_472# 0.001451f
C5342 _086_ _267_/a_1792_472# 0.002715f
C5343 _074_ FILLER_0_3_172/a_484_472# 0.001763f
C5344 FILLER_0_20_169/a_36_472# vss 0.005112f
C5345 _429_/a_36_151# FILLER_0_15_212/a_124_375# 0.059049f
C5346 _130_ _126_ 0.061836f
C5347 net26 _012_ 0.066032f
C5348 _181_ _184_ 0.022711f
C5349 _181_ _401_/a_36_68# 0.010647f
C5350 net57 _225_/a_36_160# 0.022745f
C5351 _075_ FILLER_0_7_195/a_124_375# 0.008178f
C5352 net27 result[0] 0.106157f
C5353 FILLER_0_17_38/a_572_375# _041_ 0.021754f
C5354 net81 FILLER_0_15_205/a_124_375# 0.015134f
C5355 FILLER_0_14_50/a_36_472# _174_ 0.015387f
C5356 _142_ FILLER_0_17_142/a_484_472# 0.01467f
C5357 FILLER_0_2_101/a_124_375# net14 0.0239f
C5358 FILLER_0_5_128/a_36_472# _152_ 0.013822f
C5359 _053_ FILLER_0_7_104/a_1468_375# 0.001492f
C5360 _031_ vdd 0.327674f
C5361 _090_ net21 0.038093f
C5362 mask\[9\] _438_/a_2665_112# 0.040085f
C5363 net72 _424_/a_36_151# 0.09381f
C5364 _064_ _446_/a_448_472# 0.01156f
C5365 _235_/a_67_603# _446_/a_2665_112# 0.017036f
C5366 _015_ FILLER_0_8_239/a_124_375# 0.007342f
C5367 _126_ _129_ 0.039006f
C5368 output23/a_224_472# _208_/a_36_160# 0.014541f
C5369 _093_ FILLER_0_19_142/a_124_375# 0.00346f
C5370 _413_/a_36_151# _088_ 0.001289f
C5371 FILLER_0_18_177/a_1380_472# vss -0.001894f
C5372 FILLER_0_18_177/a_1828_472# vdd 0.004845f
C5373 net52 _442_/a_1000_472# 0.016308f
C5374 _072_ _251_/a_1130_472# 0.004007f
C5375 _165_ FILLER_0_6_47/a_124_375# 0.014312f
C5376 net72 _067_ 0.055817f
C5377 _005_ _416_/a_1308_423# 0.020096f
C5378 _411_/a_448_472# net65 0.006279f
C5379 _115_ FILLER_0_10_107/a_36_472# 0.016715f
C5380 FILLER_0_14_81/a_124_375# _177_ 0.002725f
C5381 fanout53/a_36_160# FILLER_0_16_154/a_932_472# 0.001426f
C5382 _441_/a_36_151# _168_ 0.033578f
C5383 net20 FILLER_0_3_221/a_932_472# 0.054476f
C5384 output24/a_224_472# _436_/a_36_151# 0.053592f
C5385 _345_/a_36_160# FILLER_0_19_125/a_36_472# 0.006647f
C5386 net66 FILLER_0_5_54/a_484_472# 0.001863f
C5387 FILLER_0_9_60/a_124_375# vss 0.003217f
C5388 FILLER_0_9_60/a_572_375# vdd 0.031403f
C5389 _140_ FILLER_0_19_155/a_572_375# 0.040109f
C5390 _413_/a_796_472# net65 0.006888f
C5391 net18 _419_/a_2248_156# 0.014287f
C5392 _439_/a_1308_423# FILLER_0_6_47/a_3260_375# 0.001224f
C5393 ctlp[1] _421_/a_36_151# 0.010453f
C5394 net15 FILLER_0_23_60/a_36_472# 0.004561f
C5395 net61 fanout61/a_36_113# 0.023179f
C5396 _238_/a_67_603# FILLER_0_1_98/a_36_472# 0.02529f
C5397 net69 _441_/a_2665_112# 0.014995f
C5398 output20/a_224_472# _422_/a_1308_423# 0.005632f
C5399 FILLER_0_17_104/a_36_472# net14 0.012286f
C5400 net20 _088_ 0.001704f
C5401 _096_ _055_ 0.047639f
C5402 _057_ _228_/a_36_68# 0.002062f
C5403 _094_ vdd 0.717159f
C5404 FILLER_0_17_218/a_572_375# vdd 0.019414f
C5405 FILLER_0_17_218/a_124_375# vss 0.012673f
C5406 _100_ vss 0.020176f
C5407 _425_/a_2248_156# vdd 0.010067f
C5408 mask\[7\] FILLER_0_22_128/a_1828_472# 0.004503f
C5409 _069_ _429_/a_796_472# 0.003099f
C5410 net41 _450_/a_3129_107# 0.059083f
C5411 FILLER_0_11_101/a_124_375# _171_ 0.00105f
C5412 _432_/a_2665_112# vdd 0.009104f
C5413 _297_/a_36_472# vss 0.003601f
C5414 FILLER_0_17_72/a_932_472# _175_ 0.003281f
C5415 _070_ _172_ 0.237178f
C5416 FILLER_0_24_96/a_124_375# output25/a_224_472# 0.002633f
C5417 FILLER_0_0_198/a_124_375# net59 0.004565f
C5418 _170_ _241_/a_224_472# 0.001199f
C5419 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1380_472# 0.013276f
C5420 _104_ _008_ 0.135471f
C5421 net53 _427_/a_2665_112# 0.042564f
C5422 _360_/a_36_160# net47 0.011731f
C5423 trim_mask\[0\] vss 0.014228f
C5424 _103_ _046_ 0.010317f
C5425 fanout54/a_36_160# _145_ 0.009257f
C5426 net48 _070_ 0.264809f
C5427 _423_/a_36_151# FILLER_0_23_44/a_572_375# 0.059049f
C5428 _448_/a_2665_112# net22 0.010428f
C5429 net70 _043_ 0.045182f
C5430 _115_ FILLER_0_9_72/a_1468_375# 0.025664f
C5431 _098_ FILLER_0_15_212/a_1020_375# 0.00918f
C5432 _428_/a_1204_472# net74 0.009712f
C5433 net50 _439_/a_2248_156# 0.007461f
C5434 _008_ vss 0.355468f
C5435 _245_/a_672_472# net17 0.00121f
C5436 _367_/a_36_68# _160_ 0.013113f
C5437 FILLER_0_4_49/a_484_472# vss 0.002751f
C5438 FILLER_0_5_109/a_484_472# _363_/a_36_68# 0.001709f
C5439 _098_ FILLER_0_16_154/a_932_472# 0.001701f
C5440 _104_ result[8] 0.00201f
C5441 _432_/a_448_472# FILLER_0_19_171/a_572_375# 0.00184f
C5442 _431_/a_2665_112# _137_ 0.010924f
C5443 trim[0] net40 0.005988f
C5444 FILLER_0_9_28/a_1468_375# vdd 0.009854f
C5445 _319_/a_672_472# _125_ 0.002725f
C5446 net54 FILLER_0_19_142/a_124_375# 0.056556f
C5447 _096_ _126_ 0.258912f
C5448 _098_ _434_/a_36_151# 0.019342f
C5449 _098_ FILLER_0_19_111/a_36_472# 0.003915f
C5450 FILLER_0_19_47/a_572_375# _183_ 0.001186f
C5451 fanout80/a_36_113# _098_ 0.011559f
C5452 result[8] vss 0.235206f
C5453 ctlp[5] _147_ 0.001406f
C5454 ctlp[3] vdd 0.251098f
C5455 _308_/a_124_24# trim_mask\[0\] 0.018998f
C5456 _242_/a_36_160# _170_ 0.001933f
C5457 _117_ _310_/a_1133_69# 0.002654f
C5458 FILLER_0_22_86/a_36_472# vss 0.002319f
C5459 _122_ net59 0.041453f
C5460 _114_ _311_/a_1920_473# 0.005579f
C5461 en_co_clk _171_ 0.003472f
C5462 _140_ FILLER_0_22_128/a_124_375# 0.011452f
C5463 FILLER_0_19_125/a_124_375# vdd 0.032954f
C5464 FILLER_0_22_128/a_3172_472# vdd 0.003395f
C5465 FILLER_0_22_128/a_2724_472# vss 0.005195f
C5466 _108_ _295_/a_36_472# 0.014558f
C5467 _095_ _181_ 0.008117f
C5468 _299_/a_36_472# _109_ 0.030751f
C5469 FILLER_0_9_28/a_36_472# vss -0.001119f
C5470 result[8] _422_/a_1000_472# 0.001104f
C5471 net35 _435_/a_36_151# 0.038368f
C5472 _132_ _428_/a_448_472# 0.034825f
C5473 _056_ _055_ 0.155993f
C5474 _412_/a_1204_472# cal_itt\[1\] 0.001547f
C5475 net56 FILLER_0_18_139/a_1380_472# 0.048069f
C5476 ctln[6] _387_/a_36_113# 0.007687f
C5477 net64 net59 0.005832f
C5478 net68 _381_/a_36_472# 0.003421f
C5479 output38/a_224_472# _446_/a_448_472# 0.007649f
C5480 net78 vdd 0.265913f
C5481 _050_ vdd 0.484554f
C5482 FILLER_0_15_235/a_572_375# FILLER_0_14_235/a_572_375# 0.05841f
C5483 _442_/a_2248_156# net14 0.025334f
C5484 _431_/a_2560_156# FILLER_0_17_142/a_124_375# 0.001178f
C5485 _445_/a_1000_472# _034_ 0.007034f
C5486 _445_/a_2665_112# _166_ 0.002292f
C5487 net15 _447_/a_36_151# 0.001598f
C5488 FILLER_0_11_142/a_572_375# _121_ 0.003107f
C5489 _360_/a_36_160# net74 0.001912f
C5490 _030_ net40 0.002509f
C5491 net17 net6 0.063494f
C5492 _185_ _402_/a_718_527# 0.001973f
C5493 FILLER_0_24_96/a_124_375# output24/a_224_472# 0.00363f
C5494 net36 FILLER_0_18_76/a_484_472# 0.005765f
C5495 net82 FILLER_0_3_172/a_1380_472# 0.007879f
C5496 FILLER_0_5_54/a_36_472# _164_ 0.003923f
C5497 FILLER_0_8_263/a_124_375# vss 0.007944f
C5498 FILLER_0_8_263/a_36_472# vdd 0.092694f
C5499 _058_ _059_ 0.990213f
C5500 vdd FILLER_0_14_235/a_572_375# 0.006167f
C5501 vss FILLER_0_14_235/a_124_375# 0.002686f
C5502 en_co_clk FILLER_0_13_100/a_36_472# 0.001752f
C5503 FILLER_0_22_86/a_124_375# FILLER_0_23_88/a_36_472# 0.001684f
C5504 output42/a_224_472# _039_ 0.001254f
C5505 _132_ FILLER_0_12_124/a_36_472# 0.00101f
C5506 _101_ _283_/a_36_472# 0.002471f
C5507 _098_ FILLER_0_15_205/a_36_472# 0.010528f
C5508 FILLER_0_3_172/a_484_472# net65 0.003678f
C5509 _322_/a_692_472# net74 0.003192f
C5510 _446_/a_2665_112# vdd 0.044081f
C5511 result[8] _107_ 0.041984f
C5512 _210_/a_67_603# vss 0.038142f
C5513 FILLER_0_7_72/a_124_375# net50 0.009304f
C5514 _415_/a_36_151# FILLER_0_10_256/a_36_472# 0.004847f
C5515 _214_/a_36_160# vdd 0.010812f
C5516 _069_ _061_ 0.024151f
C5517 _161_ state\[1\] 0.002512f
C5518 net34 net20 0.003775f
C5519 _443_/a_796_472# vss 0.001654f
C5520 _430_/a_2665_112# FILLER_0_17_218/a_572_375# 0.002362f
C5521 _415_/a_36_151# net64 0.001735f
C5522 _112_ FILLER_0_8_247/a_932_472# 0.001185f
C5523 calibrate FILLER_0_7_233/a_36_472# 0.013262f
C5524 _068_ _055_ 0.443477f
C5525 _119_ _160_ 0.037232f
C5526 FILLER_0_12_136/a_932_472# net23 0.004375f
C5527 net20 FILLER_0_13_212/a_932_472# 0.003007f
C5528 net48 _425_/a_448_472# 0.013011f
C5529 _448_/a_2248_156# vss 0.003807f
C5530 _448_/a_2665_112# vdd 0.005876f
C5531 _122_ _227_/a_36_160# 0.005128f
C5532 output48/a_224_472# _081_ 0.007705f
C5533 net52 FILLER_0_6_47/a_3172_472# 0.047876f
C5534 _060_ vss 0.318005f
C5535 _126_ FILLER_0_11_135/a_124_375# 0.008245f
C5536 output18/a_224_472# net18 0.01698f
C5537 cal_itt\[3\] net57 0.001586f
C5538 net63 FILLER_0_19_195/a_124_375# 0.017284f
C5539 _414_/a_1000_472# cal_itt\[3\] 0.08528f
C5540 _122_ _169_ 0.014463f
C5541 calibrate _163_ 0.026892f
C5542 FILLER_0_16_57/a_572_375# net55 0.004559f
C5543 FILLER_0_16_57/a_36_472# net72 0.040135f
C5544 _017_ _134_ 0.017998f
C5545 _423_/a_36_151# vss 0.012999f
C5546 _423_/a_448_472# vdd 0.01351f
C5547 mask\[3\] _282_/a_36_160# 0.005823f
C5548 FILLER_0_14_181/a_124_375# _137_ 0.006021f
C5549 net48 _082_ 0.003853f
C5550 FILLER_0_5_54/a_932_472# net47 0.006386f
C5551 net68 _453_/a_796_472# 0.001516f
C5552 cal_count\[3\] _389_/a_36_148# 0.024777f
C5553 net57 _428_/a_1000_472# 0.024803f
C5554 net16 FILLER_0_18_53/a_36_472# 0.001532f
C5555 net55 _183_ 0.024948f
C5556 net21 net11 0.10869f
C5557 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_124_375# 0.004426f
C5558 _176_ FILLER_0_18_53/a_36_472# 0.001868f
C5559 FILLER_0_17_56/a_36_472# _041_ 0.004881f
C5560 _035_ net49 0.018245f
C5561 _073_ _080_ 0.455535f
C5562 _118_ _311_/a_3220_473# 0.001133f
C5563 fanout60/a_36_160# FILLER_0_17_282/a_124_375# 0.005489f
C5564 _343_/a_49_472# vss 0.002581f
C5565 FILLER_0_16_89/a_36_472# _136_ 0.00722f
C5566 _044_ FILLER_0_14_263/a_36_472# 0.002013f
C5567 _086_ _363_/a_36_68# 0.007567f
C5568 FILLER_0_18_100/a_36_472# FILLER_0_18_107/a_36_472# 0.002764f
C5569 output48/a_224_472# net65 0.015306f
C5570 _126_ _068_ 0.01065f
C5571 fanout62/a_36_160# FILLER_0_9_290/a_36_472# 0.001961f
C5572 fanout55/a_36_160# cal_count\[1\] 0.007256f
C5573 FILLER_0_14_81/a_36_472# _451_/a_3129_107# 0.001557f
C5574 FILLER_0_5_206/a_124_375# net59 0.008027f
C5575 _086_ FILLER_0_11_124/a_124_375# 0.016039f
C5576 FILLER_0_17_72/a_36_472# vss 0.036865f
C5577 _134_ FILLER_0_10_107/a_36_472# 0.006746f
C5578 _072_ _069_ 0.265737f
C5579 _181_ _402_/a_1296_93# 0.040412f
C5580 net22 _435_/a_36_151# 0.001559f
C5581 _413_/a_2665_112# net65 0.033675f
C5582 _414_/a_36_151# _163_ 0.001186f
C5583 net16 FILLER_0_10_28/a_124_375# 0.002225f
C5584 vss FILLER_0_6_37/a_36_472# 0.006755f
C5585 _132_ FILLER_0_17_104/a_1020_375# 0.009251f
C5586 _427_/a_796_472# vss 0.001131f
C5587 trim_mask\[4\] _370_/a_1152_472# 0.001449f
C5588 net17 _450_/a_2225_156# 0.033342f
C5589 net52 FILLER_0_2_111/a_1380_472# 0.050754f
C5590 trim_mask\[1\] vdd 0.241393f
C5591 output16/a_224_472# vdd 0.006151f
C5592 _436_/a_36_151# FILLER_0_22_107/a_124_375# 0.026916f
C5593 _105_ _292_/a_36_160# 0.027405f
C5594 _081_ _242_/a_36_160# 0.025059f
C5595 _033_ net47 0.056436f
C5596 net76 FILLER_0_3_172/a_124_375# 0.001186f
C5597 _444_/a_448_472# net42 0.002526f
C5598 _116_ vss 0.235141f
C5599 FILLER_0_12_220/a_36_472# _070_ 0.087648f
C5600 FILLER_0_7_146/a_124_375# _372_/a_170_472# 0.001188f
C5601 net63 FILLER_0_18_177/a_1828_472# 0.047684f
C5602 net52 _440_/a_2665_112# 0.005084f
C5603 FILLER_0_7_72/a_1468_375# net50 0.020186f
C5604 _321_/a_3662_472# vdd 0.001229f
C5605 FILLER_0_8_24/a_124_375# net42 0.032303f
C5606 _096_ state\[1\] 0.083332f
C5607 fanout74/a_36_113# trim_mask\[4\] 0.026261f
C5608 FILLER_0_19_55/a_124_375# FILLER_0_17_56/a_36_472# 0.001338f
C5609 _095_ FILLER_0_13_72/a_36_472# 0.00819f
C5610 FILLER_0_6_79/a_36_472# _164_ 0.008685f
C5611 _094_ _283_/a_36_472# 0.004373f
C5612 _452_/a_1040_527# _041_ 0.002066f
C5613 FILLER_0_8_107/a_36_472# _062_ 0.001832f
C5614 _046_ mask\[2\] 0.003147f
C5615 net41 _445_/a_2248_156# 0.065247f
C5616 net49 _440_/a_2665_112# 0.025303f
C5617 net39 _444_/a_36_151# 0.14155f
C5618 _157_ vdd 0.419501f
C5619 net63 FILLER_0_17_218/a_572_375# 0.006355f
C5620 ctln[1] FILLER_0_3_221/a_572_375# 0.001554f
C5621 _115_ cal_count\[3\] 0.004426f
C5622 _350_/a_665_69# mask\[6\] 0.001069f
C5623 _104_ _093_ 0.109158f
C5624 _239_/a_36_160# _065_ 0.032139f
C5625 _256_/a_1612_497# vss 0.004265f
C5626 _415_/a_2665_112# net62 0.003644f
C5627 _432_/a_2665_112# net63 0.067487f
C5628 _447_/a_2665_112# vdd 0.022038f
C5629 _447_/a_2248_156# vss 0.003961f
C5630 ctln[1] _000_ 0.223573f
C5631 FILLER_0_18_107/a_1468_375# net71 0.001292f
C5632 FILLER_0_16_73/a_572_375# _175_ 0.138524f
C5633 FILLER_0_16_89/a_932_472# net36 0.001709f
C5634 _373_/a_1060_68# _090_ 0.002234f
C5635 _091_ FILLER_0_19_171/a_1020_375# 0.005708f
C5636 _093_ vss 2.002012f
C5637 FILLER_0_16_57/a_484_472# cal_count\[1\] 0.001664f
C5638 _118_ vss 0.217218f
C5639 _117_ net21 0.016722f
C5640 mask\[9\] vdd 0.940144f
C5641 _053_ _372_/a_170_472# 0.05895f
C5642 ctln[3] FILLER_0_0_232/a_36_472# 0.015594f
C5643 net23 FILLER_0_22_128/a_3260_375# 0.012171f
C5644 FILLER_0_16_73/a_484_472# _131_ 0.007761f
C5645 _431_/a_796_472# net73 0.002306f
C5646 _137_ FILLER_0_16_154/a_1380_472# 0.005667f
C5647 net54 _433_/a_2560_156# 0.014333f
C5648 _093_ FILLER_0_18_107/a_1020_375# 0.006376f
C5649 FILLER_0_18_107/a_572_375# mask\[9\] 0.005368f
C5650 _077_ FILLER_0_9_72/a_1020_375# 0.008103f
C5651 net61 net79 0.159f
C5652 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_572_375# 0.086635f
C5653 sample fanout64/a_36_160# 0.007266f
C5654 _105_ _011_ 0.003998f
C5655 net81 fanout82/a_36_113# 0.061162f
C5656 net20 net36 0.03843f
C5657 _077_ _128_ 0.005311f
C5658 _008_ _419_/a_1000_472# 0.003267f
C5659 _104_ _109_ 0.029532f
C5660 ctln[1] FILLER_0_0_266/a_36_472# 0.011046f
C5661 FILLER_0_2_111/a_572_375# _160_ 0.001049f
C5662 _365_/a_36_68# _156_ 0.027744f
C5663 FILLER_0_16_89/a_36_472# net53 0.004701f
C5664 FILLER_0_17_218/a_572_375# _069_ 0.001464f
C5665 FILLER_0_7_59/a_484_472# _439_/a_36_151# 0.001061f
C5666 net7 output40/a_224_472# 0.006944f
C5667 _444_/a_2248_156# _054_ 0.002637f
C5668 FILLER_0_21_133/a_36_472# _433_/a_36_151# 0.001723f
C5669 net73 FILLER_0_17_104/a_1380_472# 0.003206f
C5670 _077_ _453_/a_1000_472# 0.033726f
C5671 _127_ _332_/a_36_472# 0.00288f
C5672 _440_/a_448_472# _160_ 0.004748f
C5673 _056_ state\[1\] 0.219625f
C5674 _109_ vss 0.023215f
C5675 net71 _437_/a_36_151# 0.055761f
C5676 result[9] _419_/a_1204_472# 0.019627f
C5677 _155_ FILLER_0_7_104/a_124_375# 0.007925f
C5678 output46/a_224_472# FILLER_0_20_2/a_572_375# 0.03228f
C5679 net31 mask\[5\] 0.017182f
C5680 _435_/a_36_151# vdd 0.059103f
C5681 _449_/a_36_151# FILLER_0_13_72/a_484_472# 0.001723f
C5682 fanout74/a_36_113# net74 0.007425f
C5683 _119_ _374_/a_36_68# 0.001756f
C5684 output44/a_224_472# net38 0.106923f
C5685 trimb[0] trimb[2] 0.00878f
C5686 _139_ _098_ 0.026578f
C5687 _103_ _418_/a_1308_423# 0.004778f
C5688 _065_ net41 0.001765f
C5689 _103_ _006_ 0.00205f
C5690 _000_ _074_ 0.003542f
C5691 _070_ net37 0.036662f
C5692 _126_ _138_ 0.003253f
C5693 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_124_375# 0.001597f
C5694 _443_/a_36_151# _032_ 0.0737f
C5695 _422_/a_1000_472# _109_ 0.003473f
C5696 _110_ mask\[8\] 0.05045f
C5697 _123_ vss 0.016878f
C5698 FILLER_0_21_142/a_572_375# _433_/a_2665_112# 0.001092f
C5699 FILLER_0_7_146/a_36_472# net37 0.00208f
C5700 net54 vss 0.715177f
C5701 trim_mask\[2\] FILLER_0_4_91/a_36_472# 0.003327f
C5702 FILLER_0_3_204/a_124_375# _413_/a_36_151# 0.035849f
C5703 _444_/a_2248_156# vss 0.001329f
C5704 _444_/a_2665_112# vdd 0.029351f
C5705 net34 _009_ 0.325819f
C5706 _073_ vss 0.216342f
C5707 _204_/a_67_603# _201_/a_67_603# 0.001129f
C5708 trim_val\[4\] _443_/a_36_151# 0.009986f
C5709 net25 FILLER_0_23_60/a_124_375# 0.004431f
C5710 net69 _367_/a_244_472# 0.001708f
C5711 _442_/a_2248_156# _153_ 0.0011f
C5712 net74 FILLER_0_2_127/a_124_375# 0.001389f
C5713 _079_ _078_ 0.03338f
C5714 net78 _419_/a_796_472# 0.00376f
C5715 _120_ net14 0.024442f
C5716 _160_ _034_ 0.00905f
C5717 net29 _417_/a_2665_112# 0.002977f
C5718 _412_/a_1308_423# net1 0.022273f
C5719 FILLER_0_4_144/a_484_472# net23 0.01239f
C5720 _415_/a_1204_472# net18 0.001828f
C5721 _147_ _023_ 0.004036f
C5722 net65 FILLER_0_1_212/a_36_472# 0.004414f
C5723 net20 FILLER_0_15_228/a_36_472# 0.020589f
C5724 _438_/a_2248_156# net14 0.045909f
C5725 _339_/a_36_160# FILLER_0_19_171/a_124_375# 0.006021f
C5726 _337_/a_257_69# vdd 0.002972f
C5727 _119_ _133_ 0.038875f
C5728 net52 _386_/a_124_24# 0.001051f
C5729 mask\[8\] _437_/a_2665_112# 0.007907f
C5730 _012_ FILLER_0_23_60/a_36_472# 0.001572f
C5731 _412_/a_796_472# net81 0.038712f
C5732 _129_ _160_ 0.001631f
C5733 FILLER_0_21_28/a_1468_375# vdd -0.008892f
C5734 _320_/a_36_472# _043_ 0.019162f
C5735 net15 vss 1.330044f
C5736 FILLER_0_11_78/a_36_472# vss 0.00471f
C5737 FILLER_0_11_78/a_484_472# vdd 0.001756f
C5738 ctlp[2] _420_/a_2665_112# 0.01544f
C5739 FILLER_0_21_142/a_572_375# vdd 0.002442f
C5740 net55 FILLER_0_21_28/a_3172_472# 0.06297f
C5741 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_572_375# 0.086635f
C5742 _265_/a_244_68# cal_itt\[0\] 0.003127f
C5743 _028_ _363_/a_244_472# 0.002693f
C5744 net82 FILLER_0_4_213/a_36_472# 0.003042f
C5745 _430_/a_2248_156# _092_ 0.003124f
C5746 net17 trim[3] 0.001664f
C5747 net66 _167_ 0.016569f
C5748 FILLER_0_22_86/a_932_472# _026_ 0.001587f
C5749 net28 _094_ 0.007842f
C5750 _055_ _113_ 0.153988f
C5751 net27 FILLER_0_12_236/a_124_375# 0.044776f
C5752 _125_ _062_ 0.061735f
C5753 FILLER_0_23_44/a_1380_472# vss 0.003905f
C5754 net39 _054_ 0.049797f
C5755 FILLER_0_4_107/a_1020_375# net47 0.011446f
C5756 net81 _429_/a_448_472# 0.018517f
C5757 _051_ net71 0.001617f
C5758 FILLER_0_5_164/a_572_375# net37 0.014025f
C5759 net58 sample 0.006906f
C5760 FILLER_0_18_209/a_124_375# _047_ 0.006317f
C5761 FILLER_0_6_90/a_36_472# vdd 0.00366f
C5762 FILLER_0_6_90/a_572_375# vss 0.006421f
C5763 net20 _128_ 0.041f
C5764 FILLER_0_2_171/a_124_375# net22 0.009924f
C5765 net58 net37 0.15273f
C5766 _159_ FILLER_0_2_127/a_124_375# 0.020951f
C5767 net29 _005_ 0.020239f
C5768 _418_/a_2248_156# vdd 0.00423f
C5769 _412_/a_2560_156# net1 0.005618f
C5770 fanout74/a_36_113# FILLER_0_3_142/a_124_375# 0.002073f
C5771 FILLER_0_9_28/a_1380_472# net51 0.002012f
C5772 _305_/a_36_159# _425_/a_36_151# 0.001404f
C5773 mask\[8\] net14 0.040566f
C5774 net52 FILLER_0_9_72/a_36_472# 0.014911f
C5775 _116_ _071_ 0.017991f
C5776 _122_ FILLER_0_5_181/a_36_472# 0.003016f
C5777 FILLER_0_13_142/a_1468_375# net23 0.011746f
C5778 _445_/a_2665_112# net17 0.006445f
C5779 FILLER_0_5_128/a_572_375# vss 0.057605f
C5780 ctlp[1] FILLER_0_24_290/a_124_375# 0.050488f
C5781 _036_ _446_/a_2248_156# 0.001763f
C5782 net39 vss 0.170972f
C5783 FILLER_0_1_266/a_484_472# vss 0.001113f
C5784 _445_/a_2665_112# trim_val\[1\] 0.015206f
C5785 net51 vss 0.21065f
C5786 _126_ _113_ 0.547055f
C5787 _425_/a_448_472# net37 0.002755f
C5788 FILLER_0_24_274/a_36_472# FILLER_0_23_274/a_36_472# 0.05841f
C5789 _016_ net74 0.568682f
C5790 _086_ _053_ 0.091538f
C5791 _077_ FILLER_0_9_60/a_484_472# 0.024249f
C5792 cal_count\[3\] _134_ 0.011364f
C5793 ctln[4] ctln[5] 0.031901f
C5794 net52 _453_/a_2248_156# 0.011419f
C5795 FILLER_0_11_109/a_36_472# _120_ 0.014554f
C5796 _258_/a_36_160# net76 0.015203f
C5797 net75 _426_/a_1308_423# 0.002552f
C5798 _402_/a_1948_68# cal_count\[1\] 0.037053f
C5799 cal_itt\[3\] FILLER_0_6_177/a_572_375# 0.00225f
C5800 _137_ FILLER_0_19_155/a_572_375# 0.030256f
C5801 net73 _137_ 0.047989f
C5802 net82 net37 0.037195f
C5803 net48 calibrate 0.482314f
C5804 _442_/a_36_151# FILLER_0_2_127/a_36_472# 0.012873f
C5805 net64 mask\[2\] 0.046428f
C5806 net82 FILLER_0_3_221/a_1468_375# 0.009095f
C5807 _140_ _433_/a_36_151# 0.020943f
C5808 _350_/a_49_472# vss 0.001319f
C5809 FILLER_0_8_247/a_1020_375# calibrate 0.008393f
C5810 vdd _022_ 0.082842f
C5811 trim_val\[4\] net59 0.062701f
C5812 FILLER_0_16_89/a_572_375# vdd 0.005006f
C5813 FILLER_0_1_204/a_124_375# vdd 0.047704f
C5814 ctlp[1] FILLER_0_24_274/a_1380_472# 0.008573f
C5815 _430_/a_1204_472# net22 0.028536f
C5816 _079_ _263_/a_224_472# 0.002505f
C5817 output26/a_224_472# _423_/a_36_151# 0.011936f
C5818 FILLER_0_3_172/a_2724_472# net22 0.012284f
C5819 FILLER_0_5_212/a_36_472# vss 0.00578f
C5820 FILLER_0_8_37/a_484_472# _220_/a_67_603# 0.005759f
C5821 _094_ net77 0.00405f
C5822 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_36_472# 0.086635f
C5823 _422_/a_2560_156# mask\[7\] 0.010664f
C5824 net41 _034_ 0.026084f
C5825 FILLER_0_12_20/a_572_375# net40 0.007477f
C5826 _000_ net65 0.093773f
C5827 net35 net25 0.129685f
C5828 _181_ _185_ 0.061846f
C5829 net35 net23 0.04007f
C5830 net30 result[3] 0.002746f
C5831 net58 _264_/a_224_472# 0.001803f
C5832 _093_ _027_ 0.047164f
C5833 net38 vdd 0.906502f
C5834 _106_ FILLER_0_17_218/a_124_375# 0.004655f
C5835 FILLER_0_15_290/a_124_375# net79 0.051113f
C5836 _427_/a_796_472# _095_ 0.007281f
C5837 net27 _426_/a_1000_472# 0.002971f
C5838 net62 FILLER_0_15_290/a_36_472# 0.009046f
C5839 _053_ FILLER_0_6_47/a_1380_472# 0.004472f
C5840 _232_/a_67_603# _160_ 0.001684f
C5841 net27 FILLER_0_9_290/a_124_375# 0.002657f
C5842 net16 _186_ 0.225785f
C5843 _228_/a_36_68# vss 0.031389f
C5844 FILLER_0_4_123/a_36_472# _160_ 0.050308f
C5845 FILLER_0_24_96/a_36_472# net14 0.002882f
C5846 net38 FILLER_0_20_15/a_484_472# 0.003376f
C5847 _092_ _293_/a_36_472# 0.004828f
C5848 net74 FILLER_0_13_142/a_36_472# 0.003568f
C5849 _428_/a_796_472# _017_ 0.025239f
C5850 FILLER_0_2_171/a_124_375# vdd 0.042659f
C5851 FILLER_0_5_54/a_932_472# FILLER_0_6_47/a_1828_472# 0.026657f
C5852 _158_ vdd 0.131365f
C5853 _008_ _106_ 0.034748f
C5854 _211_/a_36_160# _436_/a_36_151# 0.068534f
C5855 _013_ FILLER_0_21_28/a_1828_472# 0.003978f
C5856 _444_/a_36_151# net47 0.016691f
C5857 _016_ FILLER_0_12_136/a_124_375# 0.008914f
C5858 _256_/a_36_68# _076_ 0.079206f
C5859 _127_ FILLER_0_11_124/a_36_472# 0.001641f
C5860 net58 FILLER_0_9_282/a_572_375# 0.006142f
C5861 _390_/a_36_68# _070_ 0.047478f
C5862 net63 _435_/a_36_151# 0.017194f
C5863 _322_/a_1084_68# _129_ 0.00419f
C5864 result[4] net30 0.298966f
C5865 FILLER_0_8_107/a_36_472# net14 0.001596f
C5866 _307_/a_672_472# _096_ 0.001367f
C5867 FILLER_0_18_107/a_484_472# vdd 0.035309f
C5868 FILLER_0_18_107/a_36_472# vss 0.003245f
C5869 net31 _199_/a_36_160# 0.007888f
C5870 _434_/a_1000_472# mask\[6\] 0.021582f
C5871 _103_ mask\[2\] 0.002168f
C5872 net57 _306_/a_36_68# 0.042596f
C5873 net24 FILLER_0_22_86/a_1380_472# 0.003096f
C5874 _302_/a_224_472# vss 0.005149f
C5875 output29/a_224_472# net19 0.09445f
C5876 _132_ _136_ 0.034253f
C5877 FILLER_0_7_104/a_36_472# vss 0.002797f
C5878 FILLER_0_7_104/a_484_472# vdd 0.021325f
C5879 output32/a_224_472# result[5] 0.047325f
C5880 _424_/a_36_151# vdd 0.125156f
C5881 FILLER_0_18_2/a_3260_375# FILLER_0_19_28/a_484_472# 0.001684f
C5882 FILLER_0_18_139/a_1380_472# _145_ 0.002077f
C5883 net66 vdd 0.646189f
C5884 _426_/a_36_151# net19 0.04851f
C5885 mask\[4\] FILLER_0_18_171/a_36_472# 0.01222f
C5886 _119_ _121_ 0.007336f
C5887 _074_ _162_ 0.112872f
C5888 mask\[4\] FILLER_0_18_177/a_36_472# 0.018019f
C5889 ctln[1] net18 0.004646f
C5890 net55 FILLER_0_21_60/a_484_472# 0.098472f
C5891 _067_ vdd 0.853589f
C5892 net78 net77 0.252376f
C5893 _189_/a_67_603# vss 0.004088f
C5894 net50 _441_/a_36_151# 0.060777f
C5895 net52 _441_/a_1308_423# 0.059264f
C5896 FILLER_0_4_107/a_124_375# _153_ 0.073219f
C5897 FILLER_0_4_107/a_1020_375# _154_ 0.013746f
C5898 FILLER_0_12_28/a_124_375# net40 0.047331f
C5899 FILLER_0_19_47/a_36_472# FILLER_0_18_37/a_1020_375# 0.001684f
C5900 FILLER_0_18_2/a_2364_375# net40 0.002024f
C5901 _088_ FILLER_0_3_212/a_36_472# 0.005583f
C5902 FILLER_0_12_236/a_36_472# _060_ 0.014046f
C5903 FILLER_0_4_144/a_484_472# net57 0.003724f
C5904 _068_ _160_ 0.003424f
C5905 fanout60/a_36_160# vdd 0.090968f
C5906 ctln[4] net59 0.10527f
C5907 FILLER_0_21_142/a_484_472# _098_ 0.001158f
C5908 FILLER_0_8_107/a_124_375# _131_ 0.001624f
C5909 _162_ _076_ 0.008623f
C5910 _407_/a_36_472# _181_ 0.035594f
C5911 net2 vss 0.213737f
C5912 net18 _417_/a_448_472# 0.03772f
C5913 _030_ _168_ 0.015729f
C5914 _181_ cal_count\[0\] 0.001114f
C5915 _417_/a_36_151# result[3] 0.006379f
C5916 _417_/a_1308_423# net30 0.007538f
C5917 _072_ _375_/a_1612_497# 0.002646f
C5918 ctlp[1] _010_ 0.002794f
C5919 ctln[4] FILLER_0_0_198/a_124_375# 0.015879f
C5920 _441_/a_796_472# _030_ 0.024278f
C5921 _187_ vdd 0.194575f
C5922 _119_ _312_/a_672_472# 0.00145f
C5923 _028_ vss 0.410396f
C5924 _093_ FILLER_0_18_139/a_484_472# 0.008683f
C5925 _437_/a_2248_156# vdd 0.054674f
C5926 fanout75/a_36_113# _081_ 0.015843f
C5927 en_co_clk _390_/a_244_472# 0.001238f
C5928 net61 _422_/a_448_472# 0.006042f
C5929 fanout80/a_36_113# net21 0.021603f
C5930 FILLER_0_3_172/a_2724_472# vdd 0.006405f
C5931 _129_ _133_ 0.080636f
C5932 net32 result[6] 0.048987f
C5933 result[7] _420_/a_2560_156# 0.001179f
C5934 _127_ _428_/a_2665_112# 0.001162f
C5935 _077_ _114_ 0.047702f
C5936 FILLER_0_19_171/a_932_472# _434_/a_36_151# 0.00271f
C5937 FILLER_0_23_282/a_124_375# FILLER_0_23_274/a_124_375# 0.003732f
C5938 _273_/a_36_68# _055_ 0.081216f
C5939 state\[1\] _113_ 0.107642f
C5940 fanout61/a_36_113# net62 0.031315f
C5941 trimb[1] _452_/a_2225_156# 0.004072f
C5942 mask\[8\] _148_ 0.356546f
C5943 _012_ FILLER_0_23_44/a_572_375# 0.002827f
C5944 FILLER_0_4_213/a_572_375# net59 0.061684f
C5945 cal_count\[3\] FILLER_0_12_196/a_124_375# 0.007717f
C5946 FILLER_0_3_54/a_124_375# vdd 0.029897f
C5947 mask\[3\] _137_ 0.231419f
C5948 vdd rstn 0.160093f
C5949 _044_ _416_/a_2665_112# 0.01372f
C5950 result[4] _417_/a_36_151# 0.010571f
C5951 net57 _395_/a_36_488# 0.026081f
C5952 vss clkc 0.0311f
C5953 _035_ net40 0.068572f
C5954 FILLER_0_22_177/a_36_472# _146_ 0.002f
C5955 _098_ _023_ 0.004191f
C5956 _045_ vss 0.032891f
C5957 FILLER_0_22_177/a_124_375# _435_/a_36_151# 0.059049f
C5958 ctlp[1] FILLER_0_23_282/a_36_472# 0.003169f
C5959 FILLER_0_14_181/a_36_472# vss 0.002955f
C5960 net57 FILLER_0_13_142/a_1468_375# 0.011369f
C5961 _098_ FILLER_0_20_98/a_124_375# 0.012779f
C5962 FILLER_0_9_28/a_484_472# net41 0.042989f
C5963 net34 FILLER_0_22_128/a_3260_375# 0.006974f
C5964 net61 _108_ 0.030767f
C5965 net69 _160_ 0.077526f
C5966 FILLER_0_2_171/a_124_375# FILLER_0_2_165/a_124_375# 0.003598f
C5967 FILLER_0_15_205/a_36_472# net21 0.007503f
C5968 _412_/a_1308_423# net76 0.023786f
C5969 net34 net33 0.509436f
C5970 valid vss 0.308766f
C5971 _140_ FILLER_0_22_128/a_3172_472# 0.005458f
C5972 net61 net19 0.132027f
C5973 _322_/a_848_380# FILLER_0_9_142/a_36_472# 0.011591f
C5974 net23 _433_/a_2665_112# 0.015555f
C5975 FILLER_0_17_226/a_124_375# mask\[3\] 0.010642f
C5976 net20 _274_/a_36_68# 0.021022f
C5977 FILLER_0_18_107/a_124_375# net14 0.005202f
C5978 _077_ _176_ 0.00497f
C5979 net15 _095_ 0.056214f
C5980 _132_ net53 0.035348f
C5981 fanout76/a_36_160# net2 0.023033f
C5982 net64 FILLER_0_12_220/a_1468_375# 0.01836f
C5983 net71 _436_/a_36_151# 0.03535f
C5984 FILLER_0_8_247/a_36_472# vss 0.003706f
C5985 FILLER_0_8_247/a_484_472# vdd 0.005485f
C5986 FILLER_0_4_49/a_572_375# _440_/a_36_151# 0.073306f
C5987 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1468_375# 0.016748f
C5988 _096_ FILLER_0_15_180/a_572_375# 0.001972f
C5989 _050_ _140_ 0.001f
C5990 FILLER_0_24_96/a_36_472# ctlp[7] 0.001551f
C5991 _269_/a_36_472# _260_/a_36_68# 0.002875f
C5992 _426_/a_2248_156# _060_ 0.00106f
C5993 net55 FILLER_0_18_37/a_1468_375# 0.009059f
C5994 _066_ vdd 0.14893f
C5995 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_36_472# 0.086635f
C5996 net15 _036_ 0.036489f
C5997 _322_/a_848_380# _128_ 0.012288f
C5998 _168_ trim_mask\[3\] 0.007154f
C5999 net78 _421_/a_448_472# 0.025808f
C6000 net47 _054_ 0.171966f
C6001 FILLER_0_16_73/a_36_472# net55 0.002576f
C6002 FILLER_0_16_255/a_36_472# _094_ 0.005892f
C6003 _152_ _160_ 0.286108f
C6004 _091_ _043_ 0.041409f
C6005 _374_/a_36_68# _056_ 0.011052f
C6006 FILLER_0_21_133/a_124_375# _098_ 0.006462f
C6007 net81 _138_ 0.006815f
C6008 net38 _450_/a_1353_112# 0.02208f
C6009 result[7] net32 0.103491f
C6010 _011_ _422_/a_1308_423# 0.001997f
C6011 net47 _278_/a_36_160# 0.001838f
C6012 net4 _269_/a_36_472# 0.033296f
C6013 _086_ _395_/a_1492_488# 0.001769f
C6014 FILLER_0_12_136/a_1020_375# state\[2\] 0.001952f
C6015 net25 vdd 0.195306f
C6016 net23 vdd 1.576398f
C6017 _114_ _225_/a_36_160# 0.003628f
C6018 output26/a_224_472# FILLER_0_23_44/a_1380_472# 0.0323f
C6019 trim_mask\[4\] vss 0.641217f
C6020 FILLER_0_4_49/a_36_472# _160_ 0.00202f
C6021 FILLER_0_14_50/a_124_375# _181_ 0.00402f
C6022 FILLER_0_13_80/a_124_375# FILLER_0_13_72/a_572_375# 0.012001f
C6023 net47 vss 0.919407f
C6024 _444_/a_2560_156# net67 0.012781f
C6025 _178_ net47 0.09023f
C6026 net52 _443_/a_2560_156# 0.020855f
C6027 output6/a_224_472# net6 0.076605f
C6028 net58 net8 0.175026f
C6029 net80 _434_/a_36_151# 0.067037f
C6030 FILLER_0_16_57/a_1468_375# vss 0.062643f
C6031 FILLER_0_16_57/a_36_472# vdd 0.088011f
C6032 _315_/a_716_497# _120_ 0.001321f
C6033 _387_/a_36_113# _037_ 0.003577f
C6034 net35 _436_/a_2248_156# 0.014499f
C6035 net80 fanout80/a_36_113# 0.004615f
C6036 _132_ FILLER_0_14_107/a_124_375# 0.003315f
C6037 _112_ _316_/a_124_24# 0.032665f
C6038 _414_/a_36_151# _003_ 0.021191f
C6039 _115_ net52 0.022268f
C6040 _322_/a_1084_68# _068_ 0.001022f
C6041 _127_ _070_ 0.031272f
C6042 net15 _449_/a_448_472# 0.040076f
C6043 _012_ vss 0.454371f
C6044 FILLER_0_5_128/a_124_375# _360_/a_36_160# 0.005705f
C6045 sample calibrate 0.001861f
C6046 fanout54/a_36_160# FILLER_0_19_155/a_124_375# 0.005705f
C6047 FILLER_0_15_212/a_36_472# vss 0.002853f
C6048 FILLER_0_10_214/a_124_375# _090_ 0.072741f
C6049 FILLER_0_15_212/a_1020_375# mask\[1\] 0.017527f
C6050 _106_ _093_ 0.045972f
C6051 net72 _452_/a_36_151# 0.040035f
C6052 calibrate net37 0.101109f
C6053 FILLER_0_11_109/a_124_375# vdd 0.079069f
C6054 trimb[1] net44 0.089379f
C6055 net16 _063_ 0.038576f
C6056 fanout71/a_36_113# FILLER_0_20_107/a_36_472# 0.001645f
C6057 _195_/a_67_603# _045_ 0.004028f
C6058 _345_/a_36_160# _098_ 0.002041f
C6059 FILLER_0_5_172/a_124_375# vss 0.028247f
C6060 FILLER_0_5_172/a_36_472# vdd 0.092294f
C6061 FILLER_0_4_177/a_36_472# _386_/a_848_380# 0.007646f
C6062 _065_ _447_/a_796_472# 0.007495f
C6063 _110_ _423_/a_2665_112# 0.001668f
C6064 FILLER_0_20_169/a_36_472# _098_ 0.007354f
C6065 net79 FILLER_0_15_282/a_572_375# 0.01043f
C6066 trim_mask\[1\] FILLER_0_6_47/a_2364_375# 0.007169f
C6067 FILLER_0_9_223/a_36_472# vss 0.019592f
C6068 net62 FILLER_0_15_282/a_36_472# 0.013655f
C6069 _083_ _001_ 0.002625f
C6070 _067_ _450_/a_1353_112# 0.007106f
C6071 _025_ _352_/a_49_472# 0.003933f
C6072 _287_/a_36_472# _099_ 0.030964f
C6073 fanout80/a_36_113# mask\[1\] 0.020046f
C6074 net37 net21 0.03272f
C6075 _171_ _172_ 0.104216f
C6076 FILLER_0_15_142/a_124_375# vss 0.009207f
C6077 mask\[5\] FILLER_0_20_193/a_484_472# 0.02147f
C6078 _144_ _433_/a_2560_156# 0.01064f
C6079 _052_ FILLER_0_18_53/a_572_375# 0.001631f
C6080 _074_ _076_ 0.03553f
C6081 _000_ FILLER_0_0_232/a_124_375# 0.001391f
C6082 _411_/a_2248_156# vdd 0.006283f
C6083 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_124_375# 0.012222f
C6084 FILLER_0_15_59/a_484_472# vss 0.007866f
C6085 ctlp[8] net35 0.001859f
C6086 FILLER_0_4_197/a_932_472# net76 0.003693f
C6087 _414_/a_448_472# _003_ 0.023209f
C6088 _254_/a_448_472# _074_ 0.002163f
C6089 net10 _411_/a_448_472# 0.010544f
C6090 output48/a_224_472# net48 0.001786f
C6091 output9/a_224_472# _412_/a_448_472# 0.001025f
C6092 _119_ _122_ 0.155432f
C6093 FILLER_0_11_101/a_36_472# _070_ 0.033113f
C6094 _141_ FILLER_0_22_128/a_3260_375# 0.003544f
C6095 net65 net18 0.879399f
C6096 output8/a_224_472# FILLER_0_3_221/a_1468_375# 0.032044f
C6097 _133_ _068_ 0.002552f
C6098 output43/a_224_472# net40 0.014984f
C6099 trim_val\[4\] FILLER_0_3_172/a_932_472# 0.001407f
C6100 net75 _265_/a_916_472# 0.001686f
C6101 net35 FILLER_0_22_128/a_1020_375# 0.010202f
C6102 result[9] net30 0.231442f
C6103 net74 vss 0.589483f
C6104 _207_/a_67_603# mask\[6\] 0.072291f
C6105 _376_/a_36_160# FILLER_0_6_79/a_36_472# 0.003913f
C6106 output9/a_224_472# net19 0.070689f
C6107 _079_ _080_ 0.022852f
C6108 net50 net16 0.015448f
C6109 net75 _253_/a_1732_68# 0.001047f
C6110 _064_ _445_/a_1000_472# 0.015908f
C6111 _119_ _227_/a_36_160# 0.01123f
C6112 FILLER_0_4_177/a_124_375# net22 0.006125f
C6113 net57 net22 0.003595f
C6114 _397_/a_36_472# net55 0.039732f
C6115 _414_/a_1000_472# net22 0.001649f
C6116 _174_ FILLER_0_15_59/a_124_375# 0.00622f
C6117 _253_/a_36_68# vss 0.002481f
C6118 net61 _419_/a_448_472# 0.024246f
C6119 state\[0\] net4 0.13193f
C6120 mask\[5\] FILLER_0_18_177/a_2364_375# 0.002726f
C6121 _411_/a_2665_112# output10/a_224_472# 0.008469f
C6122 net80 FILLER_0_22_177/a_484_472# 0.005297f
C6123 FILLER_0_17_104/a_124_375# vdd 0.030663f
C6124 _430_/a_1204_472# net63 0.013728f
C6125 output13/a_224_472# ctln[6] 0.080817f
C6126 _144_ vss 0.411237f
C6127 FILLER_0_5_88/a_124_375# net47 0.005083f
C6128 FILLER_0_15_116/a_484_472# _131_ 0.042796f
C6129 mask\[1\] FILLER_0_15_205/a_36_472# 0.006921f
C6130 _155_ _151_ 0.10611f
C6131 _450_/a_1040_527# clkc 0.001412f
C6132 _415_/a_448_472# net79 0.001602f
C6133 output28/a_224_472# output29/a_224_472# 0.00289f
C6134 _440_/a_36_151# _029_ 0.00874f
C6135 mask\[9\] _140_ 0.00126f
C6136 trim_mask\[4\] FILLER_0_2_165/a_36_472# 0.265591f
C6137 FILLER_0_12_220/a_932_472# vss 0.003677f
C6138 FILLER_0_12_220/a_1380_472# vdd 0.002025f
C6139 _058_ FILLER_0_8_156/a_36_472# 0.011885f
C6140 _091_ FILLER_0_18_209/a_484_472# 0.001212f
C6141 output42/a_224_472# vdd 0.04917f
C6142 _139_ net21 0.004991f
C6143 FILLER_0_11_109/a_124_375# _135_ 0.009057f
C6144 _173_ vss 0.063821f
C6145 _088_ net22 0.17798f
C6146 _053_ _072_ 0.001774f
C6147 _202_/a_36_160# _047_ 0.02265f
C6148 _328_/a_36_113# _114_ 0.058671f
C6149 _074_ FILLER_0_5_164/a_484_472# 0.003556f
C6150 net39 _445_/a_796_472# 0.002296f
C6151 FILLER_0_5_72/a_932_472# _029_ 0.007801f
C6152 FILLER_0_5_72/a_1468_375# trim_mask\[1\] 0.017105f
C6153 FILLER_0_22_177/a_1380_472# vss 0.001502f
C6154 ctln[1] net65 0.073241f
C6155 _159_ vss 0.102545f
C6156 mask\[9\] _424_/a_2665_112# 0.015491f
C6157 mask\[2\] FILLER_0_16_154/a_484_472# 0.028444f
C6158 FILLER_0_4_107/a_1380_472# _160_ 0.020979f
C6159 net34 net35 2.497277f
C6160 FILLER_0_18_171/a_124_375# FILLER_0_19_171/a_124_375# 0.05841f
C6161 _452_/a_1353_112# net40 0.003745f
C6162 net73 _334_/a_36_160# 0.003275f
C6163 net79 _136_ 0.00111f
C6164 net52 FILLER_0_0_130/a_36_472# 0.002743f
C6165 FILLER_0_4_49/a_124_375# _232_/a_67_603# 0.002082f
C6166 FILLER_0_24_130/a_36_472# net54 0.06125f
C6167 _430_/a_1204_472# _069_ 0.001629f
C6168 FILLER_0_6_37/a_124_375# _160_ 0.04948f
C6169 FILLER_0_19_125/a_36_472# _144_ 0.153815f
C6170 _130_ _427_/a_36_151# 0.001056f
C6171 _418_/a_1000_472# _007_ 0.001051f
C6172 _057_ _311_/a_254_473# 0.002364f
C6173 FILLER_0_22_86/a_36_472# _098_ 0.182093f
C6174 FILLER_0_17_72/a_2812_375# _131_ 0.006589f
C6175 net75 _412_/a_36_151# 0.060039f
C6176 trim[4] net40 0.017911f
C6177 net62 net79 1.615103f
C6178 result[4] fanout78/a_36_113# 0.001531f
C6179 _150_ net14 0.001303f
C6180 FILLER_0_7_72/a_2276_472# _439_/a_2248_156# 0.013656f
C6181 net55 FILLER_0_13_72/a_36_472# 0.002172f
C6182 net31 _091_ 0.001465f
C6183 vdd FILLER_0_19_134/a_124_375# 0.027957f
C6184 _065_ trim_val\[2\] 0.002278f
C6185 _154_ vss 0.200253f
C6186 FILLER_0_17_72/a_3172_472# net14 0.046864f
C6187 FILLER_0_12_136/a_124_375# vss 0.004063f
C6188 FILLER_0_12_136/a_572_375# vdd 0.016972f
C6189 fanout73/a_36_113# vdd 0.048166f
C6190 _449_/a_2665_112# vss 0.007395f
C6191 _074_ _081_ 0.070546f
C6192 _130_ _321_/a_170_472# 0.001018f
C6193 result[6] _421_/a_2665_112# 0.034452f
C6194 FILLER_0_20_87/a_36_472# net71 0.003995f
C6195 _327_/a_36_472# _127_ 0.002934f
C6196 FILLER_0_4_185/a_36_472# vss 0.002627f
C6197 net64 FILLER_0_9_282/a_124_375# 0.046477f
C6198 output44/a_224_472# FILLER_0_18_2/a_572_375# 0.001296f
C6199 mask\[0\] FILLER_0_15_212/a_1020_375# 0.001158f
C6200 _151_ _163_ 0.501188f
C6201 FILLER_0_10_78/a_124_375# _176_ 0.002785f
C6202 FILLER_0_3_142/a_36_472# vdd 0.10948f
C6203 FILLER_0_3_142/a_124_375# vss 0.008128f
C6204 _142_ FILLER_0_17_133/a_36_472# 0.069383f
C6205 _414_/a_2665_112# _077_ 0.001675f
C6206 FILLER_0_5_54/a_124_375# vdd 0.007387f
C6207 _076_ _081_ 0.010091f
C6208 _133_ _152_ 0.124374f
C6209 _414_/a_1308_423# _074_ 0.005458f
C6210 _451_/a_3129_107# _040_ 0.004116f
C6211 _442_/a_1308_423# vdd 0.00782f
C6212 _442_/a_448_472# vss 0.001428f
C6213 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_36_472# 0.009654f
C6214 FILLER_0_18_177/a_124_375# FILLER_0_20_177/a_36_472# 0.0027f
C6215 _346_/a_257_69# _141_ 0.002092f
C6216 _183_ _179_ 0.017086f
C6217 _043_ net14 0.037706f
C6218 _104_ ctlp[1] 0.076863f
C6219 net75 _112_ 0.041092f
C6220 _321_/a_170_472# _129_ 0.024601f
C6221 _070_ trim_mask\[0\] 0.006144f
C6222 _307_/a_672_472# _113_ 0.006607f
C6223 output33/a_224_472# result[6] 0.035032f
C6224 trim[0] _445_/a_36_151# 0.008302f
C6225 net38 _445_/a_1308_423# 0.006454f
C6226 net15 FILLER_0_6_47/a_2812_375# 0.002944f
C6227 fanout55/a_36_160# _043_ 0.019538f
C6228 _098_ FILLER_0_14_235/a_124_375# 0.001228f
C6229 _176_ FILLER_0_15_72/a_484_472# 0.00753f
C6230 _074_ net65 0.002666f
C6231 fanout80/a_36_113# mask\[0\] 0.002212f
C6232 _126_ FILLER_0_14_181/a_124_375# 0.004632f
C6233 FILLER_0_4_177/a_124_375# vdd 0.021637f
C6234 _449_/a_36_151# _067_ 0.031377f
C6235 ctlp[1] vss 0.32843f
C6236 net68 FILLER_0_3_54/a_36_472# 0.049455f
C6237 net57 vdd 1.260693f
C6238 _414_/a_1000_472# vdd 0.002568f
C6239 mask\[4\] FILLER_0_19_171/a_1380_472# 0.002581f
C6240 FILLER_0_19_47/a_36_472# _013_ 0.03573f
C6241 FILLER_0_14_181/a_36_472# _095_ 0.071989f
C6242 FILLER_0_19_155/a_484_472# vdd 0.003341f
C6243 FILLER_0_19_155/a_36_472# vss 0.004125f
C6244 _425_/a_36_151# _014_ 0.12681f
C6245 _414_/a_1204_472# _074_ 0.003142f
C6246 fanout82/a_36_113# _122_ 0.007118f
C6247 _105_ _291_/a_36_160# 0.002075f
C6248 ctln[2] FILLER_0_1_266/a_36_472# 0.052489f
C6249 _436_/a_2248_156# vdd 0.011151f
C6250 FILLER_0_3_221/a_484_472# vss 0.005602f
C6251 FILLER_0_3_221/a_932_472# vdd 0.005654f
C6252 FILLER_0_11_124/a_36_472# _118_ 0.002798f
C6253 _341_/a_257_69# _137_ 0.004351f
C6254 net73 FILLER_0_18_107/a_1468_375# 0.024898f
C6255 FILLER_0_21_142/a_572_375# _140_ 0.018708f
C6256 FILLER_0_8_138/a_124_375# _059_ 0.007966f
C6257 _026_ net14 0.010792f
C6258 _439_/a_1204_472# vss 0.006567f
C6259 net62 _429_/a_2560_156# 0.002164f
C6260 _088_ vdd 0.140259f
C6261 _079_ vss 0.124667f
C6262 FILLER_0_22_128/a_484_472# _433_/a_36_151# 0.001653f
C6263 FILLER_0_21_125/a_36_472# _149_ 0.008849f
C6264 net20 _274_/a_1612_497# 0.002057f
C6265 _427_/a_3041_156# net23 0.001305f
C6266 _428_/a_36_151# _043_ 0.027757f
C6267 net68 _164_ 0.189377f
C6268 net34 net22 0.031404f
C6269 net63 FILLER_0_15_212/a_484_472# 0.059367f
C6270 net19 FILLER_0_23_274/a_36_472# 0.075097f
C6271 net56 _145_ 0.009307f
C6272 _068_ _121_ 0.008802f
C6273 net62 FILLER_0_13_290/a_124_375# 0.032026f
C6274 net80 _139_ 0.178583f
C6275 net14 _156_ 0.184287f
C6276 _081_ FILLER_0_5_164/a_484_472# 0.001105f
C6277 FILLER_0_12_136/a_484_472# cal_count\[3\] 0.007275f
C6278 _069_ net23 0.418375f
C6279 _350_/a_49_472# _147_ 0.016114f
C6280 ctlp[5] mask\[7\] 0.131468f
C6281 net44 FILLER_0_12_2/a_36_472# 0.011079f
C6282 _443_/a_448_472# _170_ 0.056211f
C6283 FILLER_0_12_2/a_484_472# vss 0.001748f
C6284 _177_ vss 0.074896f
C6285 net53 FILLER_0_13_142/a_572_375# 0.001597f
C6286 _003_ FILLER_0_5_181/a_124_375# 0.009929f
C6287 net16 _039_ 0.031852f
C6288 ctlp[8] vdd 0.115254f
C6289 FILLER_0_10_37/a_36_472# vss 0.003659f
C6290 FILLER_0_24_274/a_124_375# vss 0.002674f
C6291 _448_/a_1308_423# _037_ 0.034533f
C6292 FILLER_0_10_78/a_484_472# _115_ 0.005678f
C6293 _141_ net35 0.003655f
C6294 _095_ net47 0.508892f
C6295 output32/a_224_472# _418_/a_2665_112# 0.011048f
C6296 net15 FILLER_0_5_72/a_36_472# 0.006713f
C6297 _348_/a_257_69# mask\[6\] 0.00159f
C6298 FILLER_0_22_128/a_572_375# vss 0.00243f
C6299 FILLER_0_22_128/a_1020_375# vdd 0.002503f
C6300 _217_/a_36_160# FILLER_0_19_28/a_484_472# 0.006053f
C6301 _052_ FILLER_0_19_28/a_572_375# 0.011078f
C6302 _428_/a_2665_112# _118_ 0.001007f
C6303 _301_/a_36_472# net35 0.051887f
C6304 _019_ vss 0.10954f
C6305 _139_ mask\[1\] 0.017315f
C6306 FILLER_0_20_15/a_1020_375# net40 0.005742f
C6307 _162_ _163_ 0.011497f
C6308 net20 _092_ 0.001458f
C6309 _441_/a_36_151# FILLER_0_3_78/a_124_375# 0.035849f
C6310 cal_itt\[1\] vss 0.327626f
C6311 cal_itt\[0\] vdd 0.438996f
C6312 _359_/a_636_68# _062_ 0.001578f
C6313 _088_ FILLER_0_3_172/a_2812_375# 0.002239f
C6314 _031_ FILLER_0_2_127/a_36_472# 0.016207f
C6315 net79 net4 0.386068f
C6316 FILLER_0_5_181/a_124_375# net37 0.005396f
C6317 FILLER_0_21_206/a_36_472# _434_/a_2665_112# 0.00243f
C6318 _414_/a_1308_423# _081_ 0.003429f
C6319 _070_ _060_ 0.822179f
C6320 _140_ _022_ 0.001997f
C6321 _431_/a_36_151# FILLER_0_15_116/a_572_375# 0.001543f
C6322 net67 _164_ 0.030648f
C6323 _421_/a_2248_156# mask\[7\] 0.016229f
C6324 FILLER_0_7_72/a_124_375# vdd 0.01526f
C6325 _064_ _160_ 0.006705f
C6326 net57 FILLER_0_2_165/a_124_375# 0.007153f
C6327 output36/a_224_472# _094_ 0.001477f
C6328 net29 _102_ 0.056837f
C6329 FILLER_0_15_142/a_124_375# _095_ 0.003935f
C6330 FILLER_0_5_128/a_484_472# _160_ 0.003335f
C6331 _273_/a_36_68# _223_/a_36_160# 0.002786f
C6332 _093_ _098_ 0.556613f
C6333 valid output37/a_224_472# 0.039402f
C6334 _420_/a_36_151# FILLER_0_23_274/a_36_472# 0.001723f
C6335 FILLER_0_9_282/a_484_472# vss 0.00561f
C6336 FILLER_0_6_47/a_2276_472# vdd 0.002735f
C6337 FILLER_0_6_47/a_1828_472# vss 0.003457f
C6338 _256_/a_244_497# vss 0.001274f
C6339 output48/a_224_472# net37 0.095886f
C6340 FILLER_0_20_31/a_124_375# net40 0.011967f
C6341 FILLER_0_9_28/a_36_472# net17 0.012954f
C6342 result[8] output35/a_224_472# 0.016867f
C6343 net31 _292_/a_36_160# 0.010041f
C6344 net58 FILLER_0_8_263/a_124_375# 0.001876f
C6345 FILLER_0_17_226/a_124_375# FILLER_0_17_218/a_572_375# 0.012001f
C6346 _321_/a_170_472# FILLER_0_11_135/a_124_375# 0.001153f
C6347 net34 vdd 1.161282f
C6348 _021_ FILLER_0_18_171/a_124_375# 0.004621f
C6349 net74 _095_ 0.04188f
C6350 cal_count\[2\] _402_/a_1948_68# 0.010022f
C6351 FILLER_0_7_104/a_1020_375# _151_ 0.002336f
C6352 mask\[0\] FILLER_0_13_206/a_124_375# 0.005989f
C6353 _142_ FILLER_0_17_161/a_36_472# 0.00657f
C6354 FILLER_0_13_212/a_484_472# vss 0.002397f
C6355 _443_/a_36_151# net69 0.069715f
C6356 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_36_472# 0.086635f
C6357 net26 FILLER_0_21_28/a_1916_375# 0.008721f
C6358 output8/a_224_472# net8 0.034396f
C6359 FILLER_0_24_63/a_124_375# output25/a_224_472# 0.007304f
C6360 net55 _423_/a_36_151# 0.001124f
C6361 net20 cal_itt\[2\] 0.715447f
C6362 FILLER_0_12_136/a_932_472# _114_ 0.003953f
C6363 ctlp[1] _420_/a_796_472# 0.001468f
C6364 FILLER_0_4_197/a_484_472# net76 0.003719f
C6365 _056_ net59 0.001756f
C6366 _116_ _070_ 0.166494f
C6367 result[5] _010_ 0.00244f
C6368 FILLER_0_16_37/a_124_375# _181_ 0.001198f
C6369 _446_/a_2248_156# net17 0.008375f
C6370 net9 cal_itt\[0\] 0.110446f
C6371 _072_ _395_/a_1492_488# 0.003088f
C6372 _136_ FILLER_0_17_133/a_124_375# 0.001315f
C6373 _239_/a_36_160# _064_ 0.001292f
C6374 vss FILLER_0_5_148/a_124_375# 0.018465f
C6375 vdd FILLER_0_5_148/a_572_375# -0.009701f
C6376 output27/a_224_472# FILLER_0_9_270/a_124_375# 0.001274f
C6377 FILLER_0_19_187/a_484_472# vss 0.004504f
C6378 net36 net22 0.034258f
C6379 net20 net61 0.014444f
C6380 FILLER_0_4_177/a_572_375# net76 0.009573f
C6381 net55 FILLER_0_17_72/a_36_472# 0.020422f
C6382 _381_/a_244_68# _167_ 0.001153f
C6383 FILLER_0_12_20/a_124_375# _450_/a_448_472# 0.001597f
C6384 FILLER_0_16_89/a_124_375# _451_/a_448_472# 0.001597f
C6385 FILLER_0_2_111/a_484_472# vdd 0.005951f
C6386 net54 _098_ 0.116416f
C6387 _429_/a_1204_472# net22 0.001899f
C6388 _028_ FILLER_0_6_47/a_2812_375# 0.023189f
C6389 FILLER_0_4_91/a_484_472# _160_ 0.009925f
C6390 _258_/a_36_160# _078_ 0.006096f
C6391 net50 _030_ 0.073046f
C6392 _242_/a_36_160# net37 0.02401f
C6393 net47 _385_/a_36_68# 0.011168f
C6394 _443_/a_36_151# _152_ 0.002345f
C6395 FILLER_0_5_109/a_36_472# vdd 0.042799f
C6396 ctln[1] FILLER_0_0_232/a_124_375# 0.012033f
C6397 _440_/a_1000_472# vss 0.031704f
C6398 FILLER_0_14_99/a_124_375# FILLER_0_13_100/a_36_472# 0.001597f
C6399 FILLER_0_7_72/a_1468_375# vdd 0.001135f
C6400 net18 _418_/a_796_472# 0.003044f
C6401 _070_ _118_ 0.302298f
C6402 _340_/a_36_160# vdd 0.006001f
C6403 _053_ trim_mask\[1\] 0.110786f
C6404 _423_/a_36_151# net17 0.002865f
C6405 _432_/a_36_151# _093_ 0.018324f
C6406 _006_ result[3] 0.016909f
C6407 _049_ FILLER_0_22_128/a_3172_472# 0.01125f
C6408 _068_ net59 0.001388f
C6409 _392_/a_36_68# cal_count\[3\] 0.003072f
C6410 net16 net72 0.367221f
C6411 _132_ _149_ 0.087289f
C6412 net82 _443_/a_796_472# 0.00219f
C6413 _127_ calibrate 0.004656f
C6414 FILLER_0_21_28/a_1380_472# _012_ 0.004453f
C6415 net72 _176_ 0.059793f
C6416 FILLER_0_21_286/a_484_472# net18 0.001956f
C6417 _017_ FILLER_0_14_107/a_1020_375# 0.001363f
C6418 net44 FILLER_0_20_2/a_36_472# 0.037627f
C6419 _430_/a_448_472# net81 0.003775f
C6420 net70 FILLER_0_14_107/a_36_472# 0.054561f
C6421 fanout79/a_36_160# vss 0.002268f
C6422 FILLER_0_5_54/a_1380_472# trim_mask\[1\] 0.01205f
C6423 net60 _102_ 0.008212f
C6424 FILLER_0_16_89/a_1380_472# net14 0.049391f
C6425 FILLER_0_1_266/a_572_375# net18 0.080358f
C6426 net27 FILLER_0_9_270/a_572_375# 0.043797f
C6427 net32 _204_/a_67_603# 0.037639f
C6428 _142_ FILLER_0_16_154/a_124_375# 0.004001f
C6429 net41 FILLER_0_21_28/a_572_375# 0.054443f
C6430 ctlp[1] _419_/a_1000_472# 0.005263f
C6431 _438_/a_448_472# vss 0.00615f
C6432 FILLER_0_0_96/a_124_375# vdd 0.034959f
C6433 net15 _098_ 0.003965f
C6434 net52 FILLER_0_5_72/a_124_375# 0.029702f
C6435 _141_ _433_/a_2665_112# 0.013144f
C6436 _091_ _432_/a_1204_472# 0.00563f
C6437 FILLER_0_12_2/a_572_375# net3 0.001872f
C6438 _451_/a_2225_156# vss 0.003848f
C6439 _077_ _246_/a_36_68# 0.006077f
C6440 FILLER_0_7_72/a_3260_375# vdd 0.008342f
C6441 net41 _064_ 0.301777f
C6442 _369_/a_36_68# _160_ 0.015312f
C6443 mask\[5\] FILLER_0_19_171/a_36_472# 0.002923f
C6444 FILLER_0_5_72/a_124_375# net49 0.001158f
C6445 FILLER_0_3_204/a_124_375# net22 0.031438f
C6446 net38 net43 0.016358f
C6447 result[4] _006_ 0.271278f
C6448 _414_/a_2665_112# cal_itt\[3\] 0.02392f
C6449 FILLER_0_18_2/a_2812_375# _452_/a_36_151# 0.001597f
C6450 trim_val\[1\] FILLER_0_6_37/a_36_472# 0.011347f
C6451 FILLER_0_15_2/a_124_375# vdd 0.010829f
C6452 _093_ net55 0.182194f
C6453 _411_/a_448_472# net8 0.04545f
C6454 FILLER_0_17_56/a_124_375# FILLER_0_18_53/a_484_472# 0.001597f
C6455 _074_ FILLER_0_7_233/a_36_472# 0.001341f
C6456 net57 _069_ 0.026933f
C6457 output34/a_224_472# _421_/a_2248_156# 0.001144f
C6458 _415_/a_448_472# net19 0.03569f
C6459 _088_ FILLER_0_5_198/a_572_375# 0.001374f
C6460 _079_ FILLER_0_5_198/a_36_472# 0.012251f
C6461 FILLER_0_19_28/a_572_375# net40 0.00139f
C6462 FILLER_0_9_28/a_3260_375# net51 0.001597f
C6463 net68 FILLER_0_5_54/a_572_375# 0.040374f
C6464 FILLER_0_21_142/a_484_472# mask\[7\] 0.001603f
C6465 net15 FILLER_0_7_59/a_124_375# 0.004662f
C6466 _126_ FILLER_0_13_206/a_36_472# 0.026561f
C6467 _346_/a_49_472# _144_ 0.036821f
C6468 _068_ _122_ 0.096251f
C6469 net51 cal_count\[0\] 0.030963f
C6470 trim[0] FILLER_0_3_2/a_36_472# 0.017429f
C6471 FILLER_0_20_177/a_572_375# mask\[6\] 0.001158f
C6472 FILLER_0_6_177/a_124_375# vss 0.002362f
C6473 _073_ _070_ 0.001892f
C6474 FILLER_0_6_177/a_572_375# vdd 0.02743f
C6475 _074_ _163_ 0.446493f
C6476 net36 FILLER_0_15_235/a_572_375# 0.083299f
C6477 FILLER_0_8_127/a_36_472# _077_ 0.003023f
C6478 _132_ _020_ 0.037636f
C6479 _153_ _156_ 0.539362f
C6480 _070_ _330_/a_224_472# 0.001096f
C6481 _408_/a_718_524# net17 0.012884f
C6482 _141_ vdd 0.439746f
C6483 _077_ FILLER_0_8_156/a_572_375# 0.007238f
C6484 _068_ _227_/a_36_160# 0.053563f
C6485 _348_/a_49_472# vdd 0.038046f
C6486 _417_/a_1308_423# _006_ 0.022704f
C6487 FILLER_0_7_104/a_1020_375# _131_ 0.016404f
C6488 _132_ _134_ 0.029512f
C6489 _057_ _085_ 0.543871f
C6490 _301_/a_36_472# vdd 0.013061f
C6491 _438_/a_36_151# _437_/a_36_151# 0.002668f
C6492 _052_ FILLER_0_21_28/a_3260_375# 0.002388f
C6493 _093_ FILLER_0_18_177/a_3260_375# 0.002695f
C6494 _143_ FILLER_0_17_161/a_36_472# 0.00363f
C6495 ctln[1] FILLER_0_1_266/a_572_375# 0.004319f
C6496 net36 vdd 0.939735f
C6497 _128_ net22 0.03249f
C6498 result[8] ctlp[2] 0.068359f
C6499 _076_ _163_ 0.030003f
C6500 FILLER_0_18_37/a_932_472# vdd 0.01019f
C6501 _086_ _055_ 0.113385f
C6502 _429_/a_1000_472# vss 0.006901f
C6503 _091_ FILLER_0_13_228/a_124_375# 0.001657f
C6504 net50 trim_mask\[3\] 0.001654f
C6505 net39 FILLER_0_8_2/a_36_472# 0.010296f
C6506 net74 _332_/a_36_472# 0.003752f
C6507 FILLER_0_7_195/a_124_375# calibrate 0.00576f
C6508 _432_/a_36_151# _337_/a_49_472# 0.002462f
C6509 net62 net19 0.352148f
C6510 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2724_472# 0.026657f
C6511 cal_count\[3\] _120_ 4.687877f
C6512 cal_count\[3\] _038_ 0.682941f
C6513 FILLER_0_9_72/a_36_472# _453_/a_2665_112# 0.001167f
C6514 net79 _416_/a_1308_423# 0.030119f
C6515 _044_ net30 0.005104f
C6516 _059_ _120_ 0.0127f
C6517 _430_/a_1308_423# net36 0.003317f
C6518 _053_ _444_/a_2665_112# 0.001698f
C6519 _193_/a_36_160# vdd 0.092266f
C6520 FILLER_0_7_195/a_124_375# net21 0.007906f
C6521 _061_ _311_/a_3740_473# 0.006728f
C6522 net70 vss 0.175272f
C6523 ctln[5] _448_/a_1204_472# 0.005186f
C6524 net26 _424_/a_448_472# 0.063966f
C6525 net10 _000_ 0.001954f
C6526 trimb[4] net44 0.127019f
C6527 _390_/a_36_68# _171_ 0.001252f
C6528 _140_ net23 0.06742f
C6529 FILLER_0_5_128/a_484_472# _133_ 0.037369f
C6530 FILLER_0_8_127/a_124_375# _126_ 0.001799f
C6531 FILLER_0_10_247/a_124_375# vss 0.006235f
C6532 FILLER_0_10_247/a_36_472# vdd 0.111658f
C6533 _177_ _095_ 0.004392f
C6534 input4/a_36_68# net5 0.004765f
C6535 cal vdd 0.318671f
C6536 _414_/a_36_151# FILLER_0_7_195/a_124_375# 0.059049f
C6537 _114_ _306_/a_36_68# 0.032258f
C6538 _086_ _126_ 0.063495f
C6539 FILLER_0_9_105/a_484_472# FILLER_0_10_107/a_124_375# 0.001543f
C6540 _414_/a_796_472# _089_ 0.001426f
C6541 FILLER_0_21_206/a_124_375# net33 0.001579f
C6542 ctlp[6] ctlp[7] 0.002504f
C6543 FILLER_0_22_86/a_572_375# net71 0.002239f
C6544 vss FILLER_0_22_107/a_484_472# 0.003617f
C6545 net20 FILLER_0_15_212/a_1380_472# 0.001449f
C6546 net41 output38/a_224_472# 0.017358f
C6547 FILLER_0_5_72/a_1020_375# _164_ 0.018398f
C6548 net80 _023_ 0.261119f
C6549 FILLER_0_10_107/a_124_375# vss 0.003015f
C6550 FILLER_0_10_107/a_572_375# vdd 0.043678f
C6551 FILLER_0_15_228/a_124_375# vss 0.006435f
C6552 FILLER_0_15_228/a_36_472# vdd 0.084606f
C6553 FILLER_0_12_50/a_36_472# _067_ 0.011087f
C6554 FILLER_0_3_204/a_124_375# vdd 0.023302f
C6555 _431_/a_2248_156# net73 0.003228f
C6556 net58 _073_ 0.057725f
C6557 _452_/a_36_151# vdd 0.109842f
C6558 net15 net55 1.200864f
C6559 net55 FILLER_0_11_78/a_36_472# 0.059367f
C6560 net67 FILLER_0_12_20/a_124_375# 0.007044f
C6561 FILLER_0_6_239/a_36_472# _316_/a_124_24# 0.002228f
C6562 net34 net63 0.050865f
C6563 net16 FILLER_0_17_38/a_484_472# 0.032356f
C6564 net72 _041_ 0.467856f
C6565 FILLER_0_5_164/a_484_472# _163_ 0.029894f
C6566 FILLER_0_3_204/a_36_472# net59 0.001606f
C6567 en vdd 0.282941f
C6568 net61 _009_ 0.042703f
C6569 FILLER_0_2_93/a_484_472# net69 0.0127f
C6570 _425_/a_1204_472# calibrate 0.009749f
C6571 FILLER_0_9_142/a_36_472# vdd 0.107619f
C6572 FILLER_0_9_142/a_124_375# vss 0.006851f
C6573 _072_ _311_/a_3740_473# 0.005483f
C6574 _065_ trim_val\[3\] 1.235816f
C6575 _424_/a_2560_156# _012_ 0.002513f
C6576 _378_/a_224_472# net67 0.00211f
C6577 mask\[5\] FILLER_0_20_177/a_932_472# 0.016114f
C6578 net38 FILLER_0_15_10/a_36_472# 0.020589f
C6579 _053_ FILLER_0_6_90/a_36_472# 0.002495f
C6580 net75 net1 0.098901f
C6581 _144_ _147_ 0.057955f
C6582 FILLER_0_21_133/a_124_375# mask\[7\] 0.00145f
C6583 _417_/a_2248_156# vdd 0.004032f
C6584 net57 _385_/a_244_472# 0.001506f
C6585 net19 _316_/a_848_380# 0.00558f
C6586 _024_ _435_/a_796_472# 0.006511f
C6587 FILLER_0_9_72/a_572_375# vss 0.007993f
C6588 FILLER_0_9_72/a_1020_375# vdd -0.014642f
C6589 _096_ _097_ 0.038778f
C6590 _093_ _111_ 0.555171f
C6591 mask\[5\] vss 0.528441f
C6592 FILLER_0_21_133/a_36_472# _436_/a_2248_156# 0.001148f
C6593 FILLER_0_16_107/a_36_472# _136_ 0.011469f
C6594 _057_ _062_ 0.062063f
C6595 _128_ vdd 0.217501f
C6596 input1/a_36_113# vdd 0.099655f
C6597 _073_ _082_ 0.009987f
C6598 _421_/a_2248_156# _419_/a_2248_156# 0.001364f
C6599 _081_ _163_ 0.427672f
C6600 _085_ _310_/a_49_472# 0.001093f
C6601 _073_ net82 0.028504f
C6602 net35 FILLER_0_22_86/a_1380_472# 0.00813f
C6603 _430_/a_2665_112# net36 0.003477f
C6604 FILLER_0_5_72/a_36_472# net47 0.003953f
C6605 FILLER_0_21_28/a_1020_375# net17 0.001134f
C6606 ctln[3] _411_/a_2665_112# 0.003037f
C6607 FILLER_0_24_63/a_36_472# _423_/a_2665_112# 0.001873f
C6608 _114_ _395_/a_36_488# 0.005314f
C6609 FILLER_0_13_212/a_1380_472# _043_ 0.014431f
C6610 _127_ FILLER_0_11_142/a_124_375# 0.00205f
C6611 cal_count\[2\] FILLER_0_15_2/a_572_375# 0.015401f
C6612 _015_ _426_/a_796_472# 0.007696f
C6613 state\[2\] cal_count\[3\] 0.005312f
C6614 net52 FILLER_0_2_101/a_124_375# 0.007787f
C6615 output9/a_224_472# fanout81/a_36_160# 0.012218f
C6616 net55 net51 0.007067f
C6617 _341_/a_49_472# FILLER_0_17_161/a_36_472# 0.079018f
C6618 _000_ FILLER_0_3_221/a_1468_375# 0.054354f
C6619 FILLER_0_18_177/a_2724_472# net22 0.004297f
C6620 net47 _166_ 0.034342f
C6621 result[6] net78 0.027123f
C6622 _337_/a_257_69# _137_ 0.001822f
C6623 _114_ FILLER_0_13_142/a_1468_375# 0.001931f
C6624 _098_ _437_/a_1204_472# 0.005729f
C6625 net65 _163_ 0.013462f
C6626 FILLER_0_4_152/a_124_375# FILLER_0_4_144/a_572_375# 0.012001f
C6627 mask\[8\] _213_/a_67_603# 0.039626f
C6628 net54 FILLER_0_22_128/a_932_472# 0.014735f
C6629 result[8] net21 0.166555f
C6630 FILLER_0_17_72/a_2724_472# _136_ 0.03065f
C6631 FILLER_0_14_91/a_484_472# FILLER_0_14_99/a_36_472# 0.013276f
C6632 _131_ FILLER_0_16_115/a_36_472# 0.008241f
C6633 net81 FILLER_0_15_212/a_1468_375# 0.006906f
C6634 _077_ _439_/a_2560_156# 0.012523f
C6635 vss _433_/a_448_472# 0.005349f
C6636 mask\[0\] _429_/a_1308_423# 0.019225f
C6637 _106_ ctlp[1] 0.002631f
C6638 mask\[5\] _107_ 0.01249f
C6639 _027_ _438_/a_448_472# 0.053901f
C6640 net4 net19 0.050898f
C6641 FILLER_0_3_172/a_572_375# net22 0.013048f
C6642 net20 _015_ 0.005917f
C6643 FILLER_0_20_98/a_36_472# _437_/a_36_151# 0.001723f
C6644 _094_ _418_/a_36_151# 0.041823f
C6645 _143_ FILLER_0_18_139/a_1468_375# 0.001097f
C6646 _394_/a_1336_472# FILLER_0_15_72/a_124_375# 0.016876f
C6647 _052_ _424_/a_1000_472# 0.007574f
C6648 FILLER_0_16_57/a_572_375# _131_ 0.015859f
C6649 _185_ net47 0.185634f
C6650 net34 FILLER_0_22_177/a_124_375# 0.006974f
C6651 FILLER_0_18_2/a_1468_375# _452_/a_448_472# 0.001597f
C6652 FILLER_0_5_117/a_124_375# vdd 0.035079f
C6653 net39 net17 0.099429f
C6654 FILLER_0_8_263/a_124_375# calibrate 0.006928f
C6655 FILLER_0_11_142/a_36_472# _076_ 0.003047f
C6656 _395_/a_1044_488# _085_ 0.00391f
C6657 _395_/a_36_488# _176_ 0.010116f
C6658 FILLER_0_7_72/a_2812_375# trim_mask\[0\] 0.005302f
C6659 net17 net51 0.026974f
C6660 _415_/a_2248_156# FILLER_0_11_282/a_124_375# 0.001221f
C6661 net80 FILLER_0_20_169/a_36_472# 0.024142f
C6662 net72 FILLER_0_17_64/a_124_375# 0.002236f
C6663 FILLER_0_16_107/a_572_375# vdd 0.019922f
C6664 net23 FILLER_0_21_150/a_36_472# 0.016375f
C6665 _131_ _183_ 0.227229f
C6666 _430_/a_36_151# net81 0.017255f
C6667 FILLER_0_19_195/a_36_472# vss 0.005146f
C6668 _132_ FILLER_0_18_107/a_2276_472# 0.006713f
C6669 FILLER_0_7_104/a_1468_375# _133_ 0.003206f
C6670 _093_ FILLER_0_17_72/a_1916_375# 0.017467f
C6671 trim[1] _033_ 0.015549f
C6672 _008_ _418_/a_448_472# 0.052899f
C6673 _411_/a_36_151# net75 0.033786f
C6674 net15 _216_/a_67_603# 0.060076f
C6675 output27/a_224_472# vdd 0.070751f
C6676 FILLER_0_20_177/a_124_375# vdd 0.001964f
C6677 fanout52/a_36_160# _443_/a_2665_112# 0.007884f
C6678 _256_/a_3368_68# net22 0.001285f
C6679 fanout72/a_36_113# _043_ 0.017862f
C6680 net34 _435_/a_2665_112# 0.009214f
C6681 FILLER_0_14_181/a_36_472# _098_ 0.004669f
C6682 FILLER_0_5_206/a_36_472# _081_ 0.014328f
C6683 result[9] _006_ 0.05748f
C6684 result[5] vss 0.307366f
C6685 output16/a_224_472# _447_/a_448_472# 0.003175f
C6686 output13/a_224_472# _037_ 0.019694f
C6687 trim_val\[0\] FILLER_0_6_47/a_484_472# 0.001215f
C6688 net15 _111_ 0.049514f
C6689 _365_/a_36_68# vss 0.029516f
C6690 _086_ state\[1\] 0.043298f
C6691 _429_/a_36_151# FILLER_0_15_212/a_1020_375# 0.035849f
C6692 _326_/a_36_160# _119_ 0.003944f
C6693 FILLER_0_20_15/a_124_375# vdd 0.006513f
C6694 result[9] _103_ 0.034463f
C6695 net65 FILLER_0_1_266/a_572_375# 0.002969f
C6696 mask\[7\] _297_/a_36_472# 0.003196f
C6697 _095_ _451_/a_2225_156# 0.001102f
C6698 net63 net36 0.010544f
C6699 FILLER_0_18_2/a_36_472# cal_count\[2\] 0.001929f
C6700 _181_ _179_ 0.011848f
C6701 _155_ _029_ 0.174512f
C6702 cal_count\[2\] _452_/a_448_472# 0.003314f
C6703 _062_ _310_/a_49_472# 0.020509f
C6704 ctlp[2] _109_ 0.059999f
C6705 FILLER_0_17_38/a_484_472# _041_ 0.009607f
C6706 FILLER_0_5_117/a_36_472# _163_ 0.007418f
C6707 net74 FILLER_0_11_124/a_36_472# 0.020589f
C6708 _441_/a_36_151# vdd 0.098562f
C6709 _413_/a_1000_472# net82 0.002029f
C6710 _104_ output20/a_224_472# 0.019295f
C6711 _053_ FILLER_0_7_104/a_484_472# 0.005353f
C6712 net69 _369_/a_244_472# 0.002456f
C6713 _060_ net21 0.074356f
C6714 net27 vss 0.534444f
C6715 net78 _418_/a_36_151# 0.003648f
C6716 _058_ FILLER_0_9_105/a_124_375# 0.014234f
C6717 output33/a_224_472# _204_/a_67_603# 0.00401f
C6718 output20/a_224_472# vss -0.004787f
C6719 result[7] net78 0.019651f
C6720 net75 FILLER_0_6_239/a_36_472# 0.009325f
C6721 FILLER_0_18_177/a_2724_472# vdd 0.002749f
C6722 net52 _442_/a_2248_156# 0.022954f
C6723 _035_ _445_/a_36_151# 0.002276f
C6724 _005_ _416_/a_1000_472# 0.027013f
C6725 FILLER_0_2_101/a_36_472# trim_mask\[3\] 0.013363f
C6726 net56 FILLER_0_16_154/a_932_472# 0.001401f
C6727 _441_/a_1308_423# _168_ 0.044302f
C6728 valid fanout64/a_36_160# 0.001811f
C6729 output24/a_224_472# _436_/a_1308_423# 0.005632f
C6730 FILLER_0_9_60/a_484_472# vdd 0.005181f
C6731 FILLER_0_9_60/a_36_472# vss 0.001327f
C6732 _140_ FILLER_0_19_155/a_484_472# 0.004155f
C6733 output10/a_224_472# rstn 0.001656f
C6734 net18 _419_/a_2560_156# 0.008155f
C6735 result[8] mask\[7\] 0.110637f
C6736 fanout75/a_36_113# net37 0.010418f
C6737 ctlp[1] _421_/a_1308_423# 0.002417f
C6738 FILLER_0_21_206/a_36_472# mask\[6\] 0.015735f
C6739 vdd _295_/a_36_472# 0.0083f
C6740 _429_/a_2248_156# _043_ 0.001001f
C6741 FILLER_0_17_104/a_932_472# net14 0.002113f
C6742 _069_ net36 0.032818f
C6743 FILLER_0_19_125/a_124_375# _334_/a_36_160# 0.001633f
C6744 FILLER_0_3_172/a_572_375# vdd 0.007121f
C6745 _100_ mask\[1\] 0.002229f
C6746 FILLER_0_17_218/a_484_472# vdd 0.004777f
C6747 FILLER_0_17_218/a_36_472# vss 0.006061f
C6748 net48 _074_ 1.192591f
C6749 _425_/a_2560_156# vdd 0.001827f
C6750 _425_/a_2665_112# vss 0.002983f
C6751 mask\[7\] FILLER_0_22_128/a_2724_472# 0.001055f
C6752 _069_ _429_/a_1204_472# 0.025254f
C6753 _443_/a_2248_156# net22 0.001984f
C6754 mask\[2\] FILLER_0_15_180/a_484_472# 0.00848f
C6755 FILLER_0_20_31/a_124_375# FILLER_0_20_15/a_1468_375# 0.012001f
C6756 _116_ calibrate 0.018482f
C6757 _431_/a_1204_472# _136_ 0.007382f
C6758 net63 FILLER_0_15_228/a_36_472# 0.001669f
C6759 FILLER_0_14_181/a_36_472# FILLER_0_15_180/a_124_375# 0.001723f
C6760 state\[2\] _427_/a_2665_112# 0.007007f
C6761 _415_/a_2560_156# result[1] 0.002282f
C6762 _012_ _098_ 0.002778f
C6763 _013_ FILLER_0_18_61/a_36_472# 0.01628f
C6764 net48 _076_ 0.077031f
C6765 _423_/a_36_151# FILLER_0_23_44/a_1468_375# 0.059049f
C6766 fanout62/a_36_160# result[1] 0.036633f
C6767 net62 output28/a_224_472# 0.206137f
C6768 FILLER_0_5_72/a_124_375# FILLER_0_5_54/a_1468_375# 0.005439f
C6769 _017_ _043_ 0.02569f
C6770 FILLER_0_5_109/a_484_472# _160_ 0.001598f
C6771 net26 _217_/a_36_160# 0.021067f
C6772 _098_ FILLER_0_15_212/a_36_472# 0.011079f
C6773 _428_/a_2665_112# net74 0.048822f
C6774 net58 net2 0.070564f
C6775 net50 _439_/a_2560_156# 0.006321f
C6776 _323_/a_36_113# _223_/a_36_160# 0.238626f
C6777 _429_/a_36_151# FILLER_0_15_205/a_36_472# 0.001723f
C6778 vdd _416_/a_36_151# 0.142481f
C6779 _029_ _163_ 0.007545f
C6780 _116_ net21 0.036746f
C6781 _422_/a_36_151# _108_ 0.062205f
C6782 net32 net30 0.004658f
C6783 result[2] FILLER_0_15_282/a_124_375# 0.001114f
C6784 trim[0] trim[2] 0.002289f
C6785 net16 _167_ 0.001124f
C6786 _114_ FILLER_0_9_72/a_1380_472# 0.001043f
C6787 _422_/a_36_151# net19 0.033614f
C6788 _261_/a_36_160# vss 0.05095f
C6789 net70 _095_ 0.222423f
C6790 _098_ _434_/a_1308_423# 0.007057f
C6791 _104_ _199_/a_36_160# 0.095519f
C6792 _210_/a_67_603# mask\[7\] 0.039004f
C6793 FILLER_0_9_223/a_484_472# _060_ 0.001529f
C6794 _093_ fanout54/a_36_160# 0.003506f
C6795 _117_ _090_ 0.041465f
C6796 FILLER_0_22_86/a_1380_472# vdd 0.008224f
C6797 FILLER_0_22_86/a_932_472# vss -0.001553f
C6798 _114_ _311_/a_2700_473# 0.005178f
C6799 net16 _235_/a_67_603# 0.038585f
C6800 _199_/a_36_160# vss 0.004608f
C6801 en_co_clk _172_ 0.025699f
C6802 _132_ _428_/a_796_472# 0.001472f
C6803 _093_ net21 0.032584f
C6804 net2 _082_ 0.034094f
C6805 _258_/a_36_160# _080_ 0.261387f
C6806 _118_ net21 0.007371f
C6807 net82 net2 0.451147f
C6808 _077_ FILLER_0_10_78/a_1380_472# 0.001548f
C6809 _061_ _055_ 0.853642f
C6810 _077_ _219_/a_36_160# 0.01438f
C6811 ctln[6] _170_ 0.005146f
C6812 _036_ _381_/a_36_472# 0.023012f
C6813 FILLER_0_7_146/a_124_375# net23 0.00129f
C6814 _030_ FILLER_0_3_78/a_124_375# 0.010439f
C6815 _055_ _311_/a_66_473# 0.040326f
C6816 _070_ net47 0.071795f
C6817 _411_/a_796_472# vss 0.00159f
C6818 _069_ FILLER_0_9_142/a_36_472# 0.035528f
C6819 _320_/a_224_472# vdd 0.001757f
C6820 FILLER_0_0_198/a_36_472# net11 0.056269f
C6821 net52 FILLER_0_6_79/a_36_472# 0.012286f
C6822 net28 net36 0.002537f
C6823 net82 FILLER_0_3_172/a_2276_472# 0.007729f
C6824 FILLER_0_21_206/a_124_375# net22 0.05301f
C6825 _155_ _163_ 0.296236f
C6826 _405_/a_67_603# vdd 0.034681f
C6827 vdd FILLER_0_14_235/a_484_472# 0.010228f
C6828 vss FILLER_0_14_235/a_36_472# 0.001602f
C6829 FILLER_0_7_72/a_3172_472# vss 0.002425f
C6830 _144_ _098_ 1.252524f
C6831 _442_/a_2665_112# trim_mask\[3\] 0.019514f
C6832 FILLER_0_4_197/a_36_472# _088_ 0.067725f
C6833 net58 valid 0.149817f
C6834 _173_ cal_count\[0\] 0.517178f
C6835 _128_ _069_ 0.018491f
C6836 FILLER_0_12_136/a_124_375# _428_/a_2665_112# 0.029834f
C6837 calibrate _123_ 0.016296f
C6838 _115_ FILLER_0_9_105/a_124_375# 0.002316f
C6839 net61 net33 0.043271f
C6840 _443_/a_1204_472# vss 0.005425f
C6841 _443_/a_2248_156# vdd 0.010579f
C6842 FILLER_0_14_99/a_124_375# _451_/a_1040_527# 0.010005f
C6843 FILLER_0_22_86/a_484_472# _437_/a_36_151# 0.013806f
C6844 fanout54/a_36_160# net54 0.018583f
C6845 FILLER_0_5_164/a_124_375# _066_ 0.006762f
C6846 net75 net76 0.106326f
C6847 _009_ FILLER_0_23_274/a_36_472# 0.005531f
C6848 _053_ net23 0.031487f
C6849 ctln[1] net10 0.029592f
C6850 FILLER_0_16_89/a_124_375# FILLER_0_17_72/a_1916_375# 0.026339f
C6851 FILLER_0_9_223/a_36_472# _070_ 0.006158f
C6852 _343_/a_49_472# net80 0.001646f
C6853 FILLER_0_4_152/a_36_472# _170_ 0.005476f
C6854 FILLER_0_21_142/a_124_375# net35 0.00123f
C6855 _072_ _055_ 0.083351f
C6856 _446_/a_448_472# net66 0.017696f
C6857 net48 _081_ 0.137029f
C6858 net34 _140_ 0.033459f
C6859 _429_/a_36_151# FILLER_0_13_206/a_124_375# 0.001597f
C6860 net55 net47 0.049398f
C6861 output42/a_224_472# FILLER_0_8_2/a_124_375# 0.030009f
C6862 _449_/a_2248_156# FILLER_0_13_80/a_124_375# 0.001068f
C6863 _411_/a_2248_156# output10/a_224_472# 0.019736f
C6864 _033_ _164_ 0.007117f
C6865 FILLER_0_16_57/a_1468_375# net55 0.006307f
C6866 FILLER_0_16_57/a_932_472# net72 0.004262f
C6867 _425_/a_36_151# FILLER_0_8_247/a_484_472# 0.059367f
C6868 FILLER_0_9_28/a_3172_472# _077_ 0.011059f
C6869 _423_/a_1308_423# vss 0.001726f
C6870 _423_/a_796_472# vdd 0.001494f
C6871 _114_ vdd 1.30767f
C6872 _119_ _129_ 0.055585f
C6873 sample net18 0.103617f
C6874 _086_ _160_ 0.007038f
C6875 _032_ net69 0.347645f
C6876 cal_count\[3\] _389_/a_428_148# 0.001072f
C6877 valid net82 0.060784f
C6878 net57 _428_/a_2248_156# 0.022587f
C6879 mask\[0\] _100_ 0.005921f
C6880 net55 _012_ 0.060122f
C6881 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_36_472# 0.012267f
C6882 net74 _070_ 0.394108f
C6883 FILLER_0_16_89/a_932_472# _136_ 0.045229f
C6884 output8/a_224_472# _073_ 0.043098f
C6885 _126_ FILLER_0_11_101/a_484_472# 0.001488f
C6886 net56 FILLER_0_19_155/a_124_375# 0.006762f
C6887 mask\[4\] FILLER_0_19_187/a_124_375# 0.006236f
C6888 FILLER_0_15_72/a_572_375# cal_count\[1\] 0.135344f
C6889 _000_ net8 0.021422f
C6890 FILLER_0_17_72/a_1380_472# vdd 0.001762f
C6891 FILLER_0_17_72/a_932_472# vss 0.002754f
C6892 _072_ _126_ 0.012566f
C6893 _093_ FILLER_0_18_61/a_124_375# 0.031062f
C6894 _360_/a_36_160# _153_ 0.006561f
C6895 _214_/a_36_160# _437_/a_36_151# 0.001542f
C6896 FILLER_0_5_136/a_124_375# vss 0.053395f
C6897 FILLER_0_5_136/a_36_472# vdd 0.092379f
C6898 FILLER_0_4_107/a_484_472# _369_/a_36_68# 0.001049f
C6899 FILLER_0_12_20/a_572_375# _039_ 0.005679f
C6900 _105_ ctlp[4] 0.002221f
C6901 output45/a_224_472# ctlp[0] 0.007867f
C6902 FILLER_0_16_89/a_572_375# _040_ 0.004252f
C6903 net17 net47 2.009509f
C6904 FILLER_0_3_78/a_572_375# _164_ 0.055492f
C6905 _427_/a_2248_156# vdd -0.002315f
C6906 _427_/a_1204_472# vss 0.0041f
C6907 _032_ _152_ 0.001206f
C6908 trim_mask\[4\] _370_/a_1084_68# 0.005157f
C6909 trim_val\[1\] net47 0.34878f
C6910 _432_/a_448_472# vdd 0.035246f
C6911 FILLER_0_5_172/a_124_375# FILLER_0_5_164/a_572_375# 0.012001f
C6912 _372_/a_170_472# _133_ 0.031518f
C6913 cal_count\[3\] cal_count\[2\] 0.005307f
C6914 net16 vdd 2.255325f
C6915 _340_/a_36_160# _140_ 0.062613f
C6916 net20 net62 0.058892f
C6917 _085_ vss 0.132721f
C6918 _176_ vdd 0.874707f
C6919 net76 FILLER_0_3_172/a_1020_375# 0.007439f
C6920 FILLER_0_12_220/a_932_472# _070_ 0.001282f
C6921 ctlp[1] _098_ 0.0012f
C6922 net63 FILLER_0_18_177/a_2724_472# 0.001857f
C6923 net50 _440_/a_2665_112# 0.009767f
C6924 FILLER_0_5_212/a_124_375# net59 0.045135f
C6925 FILLER_0_21_206/a_124_375# vdd 0.038521f
C6926 _093_ net80 0.818824f
C6927 output13/a_224_472# _448_/a_2248_156# 0.009013f
C6928 FILLER_0_9_223/a_572_375# _128_ 0.006559f
C6929 net82 trim_mask\[4\] 0.21475f
C6930 FILLER_0_8_24/a_36_472# net42 0.010665f
C6931 net55 net74 0.048927f
C6932 _137_ net23 0.031218f
C6933 net15 trim_mask\[2\] 0.026132f
C6934 mask\[5\] _346_/a_49_472# 0.037629f
C6935 result[9] _420_/a_2248_156# 0.046636f
C6936 FILLER_0_15_142/a_36_472# vss 0.006166f
C6937 _100_ _099_ 0.03589f
C6938 net52 _120_ 0.023363f
C6939 net52 _038_ 0.001152f
C6940 net41 _445_/a_2560_156# 0.002221f
C6941 fanout57/a_36_113# trim_mask\[4\] 0.002404f
C6942 trim[1] _444_/a_36_151# 0.001391f
C6943 mask\[7\] _109_ 0.028117f
C6944 FILLER_0_18_107/a_2812_375# _145_ 0.030158f
C6945 net15 FILLER_0_23_44/a_1468_375# 0.001307f
C6946 trim_val\[0\] _453_/a_36_151# 0.001629f
C6947 net63 FILLER_0_17_218/a_484_472# 0.002672f
C6948 ctln[1] FILLER_0_3_221/a_1468_375# 0.001235f
C6949 _258_/a_36_160# vss 0.005039f
C6950 FILLER_0_13_65/a_36_472# _174_ 0.011724f
C6951 net46 FILLER_0_20_15/a_572_375# 0.029486f
C6952 _447_/a_2560_156# vss 0.00126f
C6953 _003_ _074_ 0.00476f
C6954 _077_ net4 0.656292f
C6955 _091_ FILLER_0_19_171/a_36_472# 0.029168f
C6956 FILLER_0_16_57/a_1380_472# cal_count\[1\] 0.001568f
C6957 _124_ vdd 0.040228f
C6958 _114_ _135_ 0.018715f
C6959 _008_ _099_ 0.006163f
C6960 _053_ _372_/a_2590_472# 0.001932f
C6961 FILLER_0_11_64/a_124_375# _453_/a_2248_156# 0.001901f
C6962 net54 mask\[7\] 0.262465f
C6963 mask\[0\] FILLER_0_14_235/a_124_375# 0.009674f
C6964 net23 _049_ 0.215528f
C6965 _089_ net76 0.017609f
C6966 FILLER_0_9_72/a_124_375# _439_/a_36_151# 0.059049f
C6967 FILLER_0_5_72/a_1020_375# _440_/a_2248_156# 0.001068f
C6968 _411_/a_448_472# _073_ 0.004279f
C6969 _077_ FILLER_0_9_72/a_36_472# 0.006408f
C6970 net19 _419_/a_36_151# 0.009613f
C6971 net60 net79 0.113281f
C6972 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_484_472# 0.013277f
C6973 FILLER_0_5_212/a_124_375# _122_ 0.001352f
C6974 FILLER_0_12_28/a_124_375# _039_ 0.004669f
C6975 _405_/a_255_603# cal_count\[2\] 0.001576f
C6976 FILLER_0_18_100/a_36_472# net14 0.046864f
C6977 _413_/a_1000_472# net21 0.041643f
C6978 fanout71/a_36_113# vdd 0.028178f
C6979 FILLER_0_2_111/a_1468_375# _160_ 0.001026f
C6980 net74 _370_/a_1084_68# 0.001301f
C6981 _141_ _140_ 0.131685f
C6982 _214_/a_36_160# _051_ 0.207388f
C6983 FILLER_0_16_89/a_932_472# net53 0.012534f
C6984 FILLER_0_18_2/a_1916_375# net55 0.008235f
C6985 _216_/a_67_603# _012_ 0.001014f
C6986 net20 _429_/a_2665_112# 0.062922f
C6987 net7 net40 0.025164f
C6988 _444_/a_2560_156# _054_ 0.003269f
C6989 net31 _291_/a_36_160# 0.005683f
C6990 _140_ _348_/a_49_472# 0.023816f
C6991 _077_ _453_/a_2248_156# 0.013877f
C6992 _077_ _311_/a_1660_473# 0.001653f
C6993 net15 FILLER_0_18_61/a_124_375# 0.001179f
C6994 _061_ state\[1\] 0.02716f
C6995 net71 _437_/a_1308_423# 0.023981f
C6996 _074_ net37 0.064705f
C6997 _435_/a_1308_423# vdd 0.012856f
C6998 output46/a_224_472# FILLER_0_20_2/a_484_472# 0.001699f
C6999 FILLER_0_16_57/a_1468_375# _111_ 0.001371f
C7000 net36 _282_/a_36_160# 0.002754f
C7001 net38 _444_/a_448_472# 0.031117f
C7002 _410_/a_36_68# net51 0.014342f
C7003 mask\[0\] _060_ 0.002039f
C7004 net82 net74 0.007059f
C7005 _119_ _056_ 0.008929f
C7006 _363_/a_36_68# FILLER_0_5_109/a_36_472# 0.001024f
C7007 _256_/a_2552_68# _072_ 0.001213f
C7008 FILLER_0_21_142/a_124_375# _433_/a_2665_112# 0.004834f
C7009 _019_ _098_ 0.010193f
C7010 trim_mask\[1\] FILLER_0_5_88/a_36_472# 0.038642f
C7011 _089_ FILLER_0_5_198/a_124_375# 0.001517f
C7012 net38 FILLER_0_8_24/a_124_375# 0.001013f
C7013 cal_count\[3\] _043_ 0.721078f
C7014 _103_ _418_/a_1000_472# 0.006239f
C7015 _449_/a_2665_112# net55 0.057694f
C7016 _076_ net37 0.072179f
C7017 FILLER_0_18_76/a_124_375# vdd 0.019258f
C7018 net80 _337_/a_49_472# 0.015686f
C7019 _134_ FILLER_0_9_105/a_124_375# 0.005919f
C7020 mask\[3\] net30 0.451388f
C7021 _253_/a_36_68# _082_ 0.013108f
C7022 _228_/a_36_68# net21 0.055313f
C7023 _327_/a_36_472# net74 0.009344f
C7024 _424_/a_2665_112# net36 0.028938f
C7025 net52 fanout52/a_36_160# 0.036543f
C7026 _253_/a_36_68# net82 0.016638f
C7027 _053_ FILLER_0_5_54/a_124_375# 0.001571f
C7028 _086_ _374_/a_36_68# 0.009872f
C7029 _062_ vss 0.58133f
C7030 net69 _367_/a_36_68# 0.008893f
C7031 net20 _260_/a_36_68# 0.033776f
C7032 _016_ _428_/a_36_151# 0.001824f
C7033 _088_ _083_ 0.007169f
C7034 _414_/a_2665_112# net22 0.004067f
C7035 FILLER_0_18_2/a_1916_375# net17 0.013121f
C7036 _415_/a_1308_423# net18 0.010051f
C7037 FILLER_0_18_2/a_3260_375# vss 0.026159f
C7038 _440_/a_3041_156# _164_ 0.001221f
C7039 _092_ net22 0.010937f
C7040 net38 _452_/a_2225_156# 0.034415f
C7041 _053_ net57 0.037224f
C7042 output34/a_224_472# _093_ 0.012298f
C7043 _414_/a_1000_472# _053_ 0.029433f
C7044 _438_/a_2560_156# net14 0.049389f
C7045 _119_ _068_ 0.040944f
C7046 output35/a_224_472# FILLER_0_22_177/a_1380_472# 0.002486f
C7047 _072_ state\[1\] 0.267762f
C7048 FILLER_0_21_142/a_124_375# vdd 0.020936f
C7049 _130_ _129_ 0.021732f
C7050 ctln[8] vss 0.351742f
C7051 FILLER_0_21_28/a_2364_375# vdd -0.011393f
C7052 net20 net4 0.650415f
C7053 net82 _159_ 0.001393f
C7054 net2 calibrate 0.003482f
C7055 _041_ vdd 0.19154f
C7056 ctlp[4] mask\[6\] 0.003054f
C7057 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_484_472# 0.013277f
C7058 _265_/a_244_68# _084_ 0.016463f
C7059 FILLER_0_8_127/a_124_375# _133_ 0.001928f
C7060 _274_/a_36_68# _069_ 0.02257f
C7061 net57 FILLER_0_5_164/a_124_375# 0.040872f
C7062 _148_ FILLER_0_22_128/a_36_472# 0.010386f
C7063 _086_ _133_ 0.035637f
C7064 net36 _451_/a_36_151# 0.02414f
C7065 _003_ _081_ 0.041822f
C7066 _053_ _439_/a_2248_156# 0.002486f
C7067 net27 FILLER_0_12_236/a_36_472# 0.005414f
C7068 net54 _437_/a_448_472# 0.004418f
C7069 FILLER_0_5_212/a_124_375# FILLER_0_5_206/a_124_375# 0.005439f
C7070 _267_/a_36_472# vdd 0.005477f
C7071 FILLER_0_4_107/a_36_472# net47 0.002982f
C7072 net81 _429_/a_796_472# 0.002847f
C7073 FILLER_0_5_164/a_484_472# net37 0.013857f
C7074 FILLER_0_16_255/a_36_472# net36 0.034335f
C7075 FILLER_0_18_209/a_36_472# _047_ 0.002672f
C7076 FILLER_0_6_90/a_484_472# vss 0.00243f
C7077 FILLER_0_9_28/a_1916_375# net16 0.001431f
C7078 mask\[7\] _350_/a_49_472# 0.035293f
C7079 result[2] _005_ 0.060821f
C7080 _418_/a_2665_112# vss 0.003519f
C7081 _418_/a_2560_156# vdd 0.001506f
C7082 output10/a_224_472# cal_itt\[0\] 0.008003f
C7083 net82 FILLER_0_3_142/a_124_375# 0.018696f
C7084 FILLER_0_3_172/a_2276_472# net21 0.003603f
C7085 net14 FILLER_0_10_94/a_124_375# 0.007086f
C7086 _091_ vss 0.56693f
C7087 _433_/a_1288_156# _022_ 0.001147f
C7088 _190_/a_36_160# _450_/a_36_151# 0.002486f
C7089 FILLER_0_16_73/a_572_375# vss 0.030752f
C7090 _131_ FILLER_0_18_37/a_1468_375# 0.001151f
C7091 net52 FILLER_0_9_72/a_932_472# 0.008749f
C7092 _085_ _071_ 0.127349f
C7093 net55 _177_ 0.327874f
C7094 net70 _451_/a_448_472# 0.043107f
C7095 FILLER_0_13_142/a_484_472# net23 0.006746f
C7096 trim[1] vss 0.085436f
C7097 output37/a_224_472# _425_/a_2665_112# 0.022027f
C7098 FILLER_0_19_55/a_124_375# vdd 0.035786f
C7099 FILLER_0_16_73/a_36_472# _131_ 0.008223f
C7100 _081_ net37 1.274337f
C7101 FILLER_0_9_60/a_572_375# _439_/a_36_151# 0.001107f
C7102 _077_ _058_ 3.018054f
C7103 _141_ FILLER_0_21_150/a_36_472# 0.002773f
C7104 _114_ _069_ 0.029875f
C7105 _432_/a_448_472# net63 0.002757f
C7106 net57 _137_ 0.006142f
C7107 _096_ _161_ 0.00104f
C7108 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_36_472# 0.001963f
C7109 net75 _426_/a_1000_472# 0.002727f
C7110 FILLER_0_11_64/a_36_472# cal_count\[3\] 0.0081f
C7111 output27/a_224_472# FILLER_0_9_290/a_36_472# 0.001711f
C7112 valid calibrate 0.002363f
C7113 fanout60/a_36_160# _418_/a_36_151# 0.029017f
C7114 output29/a_224_472# vdd 0.103437f
C7115 _414_/a_2665_112# vdd 0.006496f
C7116 _011_ _299_/a_36_472# 0.004407f
C7117 sample net65 0.148853f
C7118 net82 FILLER_0_3_221/a_484_472# 0.013492f
C7119 net48 FILLER_0_7_233/a_36_472# 0.01015f
C7120 _426_/a_36_151# vdd 0.086652f
C7121 _098_ _438_/a_448_472# 0.008962f
C7122 net2 clk 0.046099f
C7123 _077_ _251_/a_244_472# 0.002492f
C7124 net65 net37 0.008382f
C7125 _092_ vdd 0.140213f
C7126 FILLER_0_8_247/a_36_472# calibrate 0.008647f
C7127 FILLER_0_12_220/a_36_472# _090_ 0.023446f
C7128 FILLER_0_7_72/a_2812_375# _028_ 0.003873f
C7129 FILLER_0_16_89/a_1468_375# vdd 0.038266f
C7130 FILLER_0_1_204/a_36_472# vss 0.002247f
C7131 _079_ _082_ 0.709481f
C7132 output14/a_224_472# trim_mask\[3\] 0.001155f
C7133 net65 FILLER_0_3_221/a_1468_375# 0.001695f
C7134 fanout81/a_36_160# net4 0.002848f
C7135 _431_/a_1308_423# vdd 0.002397f
C7136 _427_/a_2665_112# _043_ 0.002612f
C7137 FILLER_0_7_72/a_124_375# _053_ 0.014569f
C7138 _094_ _007_ 0.170362f
C7139 _065_ net69 0.051511f
C7140 FILLER_0_12_20/a_484_472# FILLER_0_12_28/a_36_472# 0.013277f
C7141 _175_ FILLER_0_15_72/a_572_375# 0.04785f
C7142 FILLER_0_2_93/a_124_375# net14 0.007439f
C7143 FILLER_0_12_20/a_484_472# net40 0.003391f
C7144 _093_ _099_ 0.001725f
C7145 net72 FILLER_0_17_38/a_124_375# 0.041464f
C7146 FILLER_0_17_64/a_124_375# vdd 0.027957f
C7147 FILLER_0_17_142/a_572_375# vdd 0.012885f
C7148 FILLER_0_17_142/a_124_375# vss 0.008753f
C7149 net18 net8 0.072251f
C7150 net64 FILLER_0_8_247/a_1468_375# 0.002559f
C7151 _120_ FILLER_0_8_156/a_36_472# 0.005842f
C7152 FILLER_0_6_47/a_124_375# vdd 0.008011f
C7153 net58 cal_itt\[1\] 0.79493f
C7154 net38 net44 0.523774f
C7155 trim[0] vdd 0.125774f
C7156 _106_ FILLER_0_17_218/a_36_472# 0.002777f
C7157 _427_/a_1204_472# _095_ 0.006692f
C7158 _069_ _176_ 0.766885f
C7159 _288_/a_224_472# _102_ 0.002528f
C7160 net27 _426_/a_2248_156# 0.002303f
C7161 _093_ FILLER_0_19_111/a_124_375# 0.00186f
C7162 _053_ FILLER_0_6_47/a_2276_472# 0.004472f
C7163 _193_/a_36_160# output30/a_224_472# 0.018f
C7164 _446_/a_1000_472# trim[3] 0.001257f
C7165 FILLER_0_16_255/a_124_375# _417_/a_2665_112# 0.003856f
C7166 _308_/a_848_380# vss 0.043591f
C7167 FILLER_0_10_78/a_484_472# _120_ 0.004669f
C7168 FILLER_0_5_109/a_572_375# vss 0.055343f
C7169 _428_/a_1204_472# _017_ 0.005148f
C7170 FILLER_0_2_171/a_36_472# vss 0.002909f
C7171 FILLER_0_5_54/a_1380_472# FILLER_0_6_47/a_2276_472# 0.026657f
C7172 fanout66/a_36_113# _160_ 0.015681f
C7173 _161_ _056_ 0.065732f
C7174 _377_/a_36_472# trim_val\[0\] 0.135527f
C7175 net20 _422_/a_36_151# 0.083307f
C7176 _443_/a_36_151# _442_/a_36_151# 0.06169f
C7177 _050_ _436_/a_36_151# 0.037103f
C7178 FILLER_0_15_142/a_36_472# _095_ 0.001526f
C7179 FILLER_0_12_236/a_572_375# FILLER_0_14_235/a_484_472# 0.001026f
C7180 FILLER_0_8_138/a_36_472# _062_ 0.001109f
C7181 FILLER_0_16_37/a_124_375# net47 0.002638f
C7182 output47/a_224_472# trimb[4] 0.044883f
C7183 _444_/a_1308_423# net47 0.040252f
C7184 _016_ FILLER_0_12_136/a_1020_375# 0.001659f
C7185 FILLER_0_15_10/a_124_375# FILLER_0_15_2/a_572_375# 0.012001f
C7186 fanout50/a_36_160# vss 0.009871f
C7187 net81 _001_ 0.012492f
C7188 net51 output6/a_224_472# 0.006462f
C7189 _133_ _313_/a_67_603# 0.002974f
C7190 net58 FILLER_0_9_282/a_484_472# 0.091905f
C7191 _127_ _131_ 0.470047f
C7192 net63 _435_/a_1308_423# 0.003621f
C7193 net41 FILLER_0_18_37/a_36_472# 0.007459f
C7194 result[4] result[3] 0.089939f
C7195 FILLER_0_8_24/a_572_375# net47 0.0353f
C7196 FILLER_0_18_107/a_1380_472# vdd 0.009462f
C7197 _130_ FILLER_0_11_135/a_124_375# 0.001198f
C7198 FILLER_0_17_200/a_572_375# _093_ 0.002355f
C7199 cal_itt\[1\] _082_ 0.921465f
C7200 _434_/a_2248_156# mask\[6\] 0.022666f
C7201 _132_ _120_ 0.034714f
C7202 _110_ vss 0.131865f
C7203 output21/a_224_472# ctlp[4] 0.052556f
C7204 net29 net19 0.305661f
C7205 mask\[4\] _201_/a_67_603# 0.029139f
C7206 net82 cal_itt\[1\] 0.396149f
C7207 cal_itt\[2\] vdd 0.267121f
C7208 FILLER_0_7_104/a_1380_472# vdd 0.011752f
C7209 _424_/a_448_472# vss 0.002076f
C7210 _424_/a_1308_423# vdd 0.002386f
C7211 _413_/a_36_151# FILLER_0_3_172/a_1468_375# 0.001252f
C7212 _030_ vdd 0.244909f
C7213 result[2] _416_/a_448_472# 0.003015f
C7214 net65 _264_/a_224_472# 0.001866f
C7215 mask\[4\] FILLER_0_18_177/a_932_472# 0.016924f
C7216 ctln[1] net8 0.678616f
C7217 net44 _067_ 0.001203f
C7218 _150_ FILLER_0_18_76/a_572_375# 0.008337f
C7219 _106_ _199_/a_36_160# 0.003376f
C7220 mask\[3\] FILLER_0_18_171/a_36_472# 0.00262f
C7221 net78 _007_ 0.054904f
C7222 FILLER_0_16_57/a_1380_472# _175_ 0.002834f
C7223 _397_/a_36_472# _131_ 0.012338f
C7224 net50 _441_/a_1308_423# 0.032656f
C7225 net52 _441_/a_1000_472# 0.011506f
C7226 _129_ FILLER_0_11_135/a_124_375# 0.009882f
C7227 mask\[3\] FILLER_0_18_177/a_36_472# 0.005668f
C7228 FILLER_0_19_47/a_484_472# FILLER_0_18_37/a_1468_375# 0.001684f
C7229 net61 vdd 0.46584f
C7230 _161_ _068_ 0.026092f
C7231 output23/a_224_472# _050_ 0.014495f
C7232 net18 _417_/a_796_472# 0.006722f
C7233 _417_/a_1000_472# net30 0.004556f
C7234 net5 rstn 0.101356f
C7235 FILLER_0_7_72/a_1468_375# _053_ 0.014569f
C7236 _086_ _121_ 0.049499f
C7237 FILLER_0_21_28/a_2276_472# _423_/a_36_151# 0.013806f
C7238 _437_/a_2665_112# vss 0.002056f
C7239 _437_/a_2560_156# vdd 0.0026f
C7240 _093_ FILLER_0_18_139/a_1380_472# 0.007013f
C7241 _077_ _115_ 0.131611f
C7242 _428_/a_36_151# FILLER_0_14_107/a_36_472# 0.02628f
C7243 FILLER_0_3_172/a_36_472# FILLER_0_2_171/a_124_375# 0.001723f
C7244 net69 FILLER_0_2_111/a_572_375# 0.015789f
C7245 en_co_clk _390_/a_36_68# 0.086301f
C7246 _430_/a_2665_112# _092_ 0.004778f
C7247 FILLER_0_3_172/a_3172_472# vss 0.003689f
C7248 _412_/a_1000_472# net81 0.012828f
C7249 _129_ _068_ 0.104827f
C7250 output7/a_224_472# trim[3] 0.103375f
C7251 ctlp[1] ctlp[2] 0.002331f
C7252 net65 FILLER_0_9_282/a_572_375# 0.001388f
C7253 FILLER_0_13_65/a_124_375# net15 0.048002f
C7254 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_124_375# 0.009654f
C7255 _098_ FILLER_0_15_228/a_124_375# 0.080662f
C7256 FILLER_0_12_136/a_932_472# FILLER_0_13_142/a_124_375# 0.001684f
C7257 _367_/a_244_472# _157_ 0.002529f
C7258 mask\[8\] _025_ 0.036686f
C7259 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_124_375# 0.009654f
C7260 _028_ FILLER_0_7_104/a_124_375# 0.008248f
C7261 _012_ FILLER_0_23_44/a_1468_375# 0.002827f
C7262 _432_/a_2560_156# vdd 0.003219f
C7263 output31/a_224_472# net18 0.009938f
C7264 _431_/a_36_151# _131_ 0.03645f
C7265 FILLER_0_4_213/a_484_472# net59 0.048997f
C7266 _096_ _056_ 0.001946f
C7267 net55 _451_/a_2225_156# 0.031243f
C7268 FILLER_0_3_54/a_36_472# vss 0.002818f
C7269 trimb[3] vdd 0.283005f
C7270 _292_/a_36_160# vss 0.009517f
C7271 _053_ FILLER_0_7_72/a_3260_375# 0.071059f
C7272 _430_/a_448_472# mask\[2\] 0.045973f
C7273 net73 _427_/a_36_151# 0.006328f
C7274 _074_ net8 0.001023f
C7275 _132_ mask\[8\] 0.029292f
C7276 input2/a_36_113# net2 0.015844f
C7277 net45 ctlp[0] 0.001134f
C7278 FILLER_0_14_91/a_572_375# _176_ 0.002444f
C7279 _359_/a_36_488# vdd 0.083138f
C7280 _045_ mask\[1\] 0.024178f
C7281 FILLER_0_22_177/a_1020_375# _435_/a_36_151# 0.059049f
C7282 FILLER_0_19_155/a_124_375# _145_ 0.006057f
C7283 _372_/a_170_472# _122_ 0.018399f
C7284 ctln[4] FILLER_0_0_232/a_36_472# 0.012298f
C7285 result[9] _421_/a_1204_472# 0.014964f
C7286 FILLER_0_6_239/a_124_375# FILLER_0_8_239/a_36_472# 0.001512f
C7287 net57 FILLER_0_13_142/a_484_472# 0.011685f
C7288 vss net14 1.003274f
C7289 _406_/a_36_159# vdd 0.020825f
C7290 FILLER_0_14_181/a_36_472# mask\[1\] 0.006352f
C7291 FILLER_0_21_125/a_572_375# vdd -0.013698f
C7292 mask\[5\] _098_ 1.316993f
C7293 _031_ _160_ 0.004547f
C7294 FILLER_0_15_72/a_124_375# vdd 0.020511f
C7295 FILLER_0_2_171/a_36_472# FILLER_0_2_165/a_36_472# 0.003468f
C7296 fanout55/a_36_160# vss 0.005203f
C7297 net34 _049_ 0.048403f
C7298 net60 net19 0.102311f
C7299 _053_ FILLER_0_6_177/a_572_375# 0.01663f
C7300 FILLER_0_24_130/a_124_375# vdd 0.027763f
C7301 net43 FILLER_0_20_15/a_124_375# 0.005925f
C7302 _257_/a_36_472# _077_ 0.019883f
C7303 net10 FILLER_0_0_232/a_124_375# 0.022977f
C7304 mask\[5\] _205_/a_36_160# 0.003775f
C7305 trim_mask\[3\] vdd 0.233305f
C7306 _164_ vss 0.597051f
C7307 output42/a_224_472# FILLER_0_8_24/a_124_375# 0.001168f
C7308 net47 FILLER_0_4_91/a_124_375# 0.009482f
C7309 FILLER_0_8_247/a_1380_472# vdd 0.036604f
C7310 net10 net11 0.007522f
C7311 FILLER_0_4_49/a_484_472# _440_/a_36_151# 0.006095f
C7312 _104_ _011_ 0.021454f
C7313 _305_/a_36_159# net59 0.007898f
C7314 net81 _094_ 0.004737f
C7315 _323_/a_36_113# net64 0.06154f
C7316 net55 FILLER_0_18_37/a_484_472# 0.006153f
C7317 net81 _425_/a_2248_156# 0.058229f
C7318 _069_ _267_/a_36_472# 0.003607f
C7319 _431_/a_36_151# net56 0.001371f
C7320 FILLER_0_9_28/a_1020_375# net68 0.004803f
C7321 _308_/a_124_24# net14 0.005016f
C7322 _011_ vss 0.003987f
C7323 net72 FILLER_0_17_56/a_572_375# 0.004473f
C7324 _070_ FILLER_0_10_107/a_124_375# 0.009848f
C7325 _441_/a_2248_156# _164_ 0.040396f
C7326 _374_/a_36_68# _061_ 0.026111f
C7327 FILLER_0_3_221/a_36_472# net59 0.075858f
C7328 output31/a_224_472# _417_/a_448_472# 0.008149f
C7329 _428_/a_448_472# vdd 0.034564f
C7330 mask\[3\] _046_ 0.018595f
C7331 _428_/a_36_151# vss 0.00285f
C7332 _098_ _433_/a_448_472# 0.027678f
C7333 _092_ net63 0.008819f
C7334 net32 _006_ 0.0012f
C7335 _411_/a_2248_156# ctln[3] 0.001208f
C7336 net38 _450_/a_836_156# 0.0039f
C7337 _011_ _422_/a_1000_472# 0.005583f
C7338 FILLER_0_14_181/a_124_375# _097_ 0.001668f
C7339 output48/a_224_472# net2 0.06309f
C7340 trimb[3] output17/a_224_472# 0.047604f
C7341 net13 vdd 0.264116f
C7342 _020_ _431_/a_1204_472# 0.002176f
C7343 _129_ _152_ 0.041257f
C7344 _091_ _095_ 0.005006f
C7345 net1 _265_/a_468_472# 0.002612f
C7346 _086_ _321_/a_170_472# 0.046783f
C7347 output9/a_224_472# vdd 0.102412f
C7348 _189_/a_67_603# mask\[0\] 0.043158f
C7349 net32 _103_ 0.038496f
C7350 _410_/a_36_68# _173_ 0.009636f
C7351 output6/a_224_472# clkc 0.017846f
C7352 _422_/a_36_151# _009_ 0.015085f
C7353 FILLER_0_10_78/a_932_472# _176_ 0.0109f
C7354 ctln[7] _442_/a_36_151# 0.007057f
C7355 net80 _434_/a_1308_423# 0.006837f
C7356 FILLER_0_16_57/a_932_472# vdd 0.005518f
C7357 FILLER_0_16_57/a_484_472# vss 0.004107f
C7358 _170_ _037_ 0.05171f
C7359 net35 _436_/a_2560_156# 0.003198f
C7360 _132_ FILLER_0_14_107/a_1020_375# 0.029702f
C7361 _112_ _316_/a_692_472# 0.001614f
C7362 FILLER_0_12_124/a_36_472# vdd 0.040515f
C7363 _115_ net50 0.008628f
C7364 _127_ _076_ 0.137964f
C7365 net15 _449_/a_796_472# 0.006722f
C7366 cal_itt\[3\] _058_ 0.002207f
C7367 _091_ FILLER_0_12_220/a_124_375# 0.006907f
C7368 _056_ _068_ 0.127175f
C7369 _246_/a_36_68# vdd 0.047419f
C7370 fanout54/a_36_160# FILLER_0_19_155/a_36_472# 0.193804f
C7371 FILLER_0_15_212/a_1380_472# vdd 0.003213f
C7372 FILLER_0_15_212/a_932_472# vss 0.019114f
C7373 FILLER_0_15_212/a_36_472# mask\[1\] 0.006865f
C7374 FILLER_0_7_72/a_572_375# net52 0.022624f
C7375 FILLER_0_11_109/a_36_472# vss 0.003131f
C7376 _072_ _374_/a_36_68# 0.061028f
C7377 _141_ _137_ 0.40175f
C7378 _092_ _069_ 0.040267f
C7379 net20 _419_/a_36_151# 0.001225f
C7380 net54 _436_/a_448_472# 0.006129f
C7381 _094_ net30 0.188507f
C7382 _065_ _447_/a_1204_472# 0.017675f
C7383 net57 _386_/a_1084_68# 0.005716f
C7384 net79 FILLER_0_15_282/a_484_472# 0.006575f
C7385 _144_ mask\[7\] 0.111088f
C7386 net36 _137_ 0.048198f
C7387 trim_mask\[1\] FILLER_0_6_47/a_3260_375# 0.003764f
C7388 _434_/a_1204_472# vdd 0.005382f
C7389 FILLER_0_5_88/a_124_375# _164_ 0.006288f
C7390 _087_ _122_ 0.007241f
C7391 net81 FILLER_0_8_263/a_36_472# 0.007373f
C7392 _000_ _073_ 0.222349f
C7393 output36/a_224_472# net36 0.009109f
C7394 _163_ net37 0.079552f
C7395 net81 FILLER_0_14_235/a_572_375# 0.029643f
C7396 net17 _381_/a_36_472# 0.002796f
C7397 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_36_472# 0.086742f
C7398 FILLER_0_1_212/a_124_375# FILLER_0_1_204/a_124_375# 0.003732f
C7399 _008_ net18 0.113775f
C7400 _077_ _134_ 0.043815f
C7401 net57 fanout56/a_36_113# 0.079542f
C7402 _416_/a_36_151# output30/a_224_472# 0.012025f
C7403 output48/a_224_472# valid 0.046397f
C7404 FILLER_0_8_127/a_36_472# vdd 0.069117f
C7405 FILLER_0_2_171/a_36_472# FILLER_0_2_177/a_36_472# 0.003468f
C7406 FILLER_0_15_290/a_124_375# vdd 0.028723f
C7407 net65 net8 0.203388f
C7408 _446_/a_2665_112# _160_ 0.013745f
C7409 _079_ net21 0.065561f
C7410 vss FILLER_0_8_156/a_124_375# 0.001766f
C7411 vdd FILLER_0_8_156/a_572_375# 0.014611f
C7412 output8/a_224_472# FILLER_0_3_221/a_484_472# 0.001699f
C7413 _141_ _049_ 0.0035f
C7414 net35 FILLER_0_22_128/a_1916_375# 0.014552f
C7415 cal_count\[3\] FILLER_0_12_50/a_124_375# 0.060164f
C7416 _275_/a_224_472# vss 0.001498f
C7417 output24/a_224_472# net71 0.001495f
C7418 mask\[0\] FILLER_0_14_181/a_36_472# 0.001234f
C7419 FILLER_0_18_100/a_124_375# _136_ 0.002528f
C7420 _414_/a_36_151# _079_ 0.037562f
C7421 net68 FILLER_0_6_47/a_572_375# 0.007672f
C7422 _064_ _445_/a_2248_156# 0.013127f
C7423 _254_/a_244_472# _072_ 0.001552f
C7424 ctlp[7] vss 0.036681f
C7425 FILLER_0_4_123/a_36_472# net69 0.001015f
C7426 FILLER_0_4_177/a_36_472# net22 0.006506f
C7427 FILLER_0_7_195/a_124_375# _074_ 0.019559f
C7428 net15 _439_/a_448_472# 0.038829f
C7429 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_124_375# 0.001597f
C7430 _086_ _122_ 0.033097f
C7431 net60 _419_/a_448_472# 0.05959f
C7432 net61 _419_/a_796_472# 0.00438f
C7433 FILLER_0_17_104/a_1020_375# vdd 0.012531f
C7434 net47 output6/a_224_472# 0.070584f
C7435 _013_ FILLER_0_18_37/a_1020_375# 0.023067f
C7436 _161_ _113_ 0.201931f
C7437 FILLER_0_10_78/a_124_375# _115_ 0.001718f
C7438 output44/a_224_472# FILLER_0_18_2/a_2364_375# 0.032639f
C7439 net54 _354_/a_49_472# 0.002169f
C7440 _148_ vss 0.025751f
C7441 ctlp[1] FILLER_0_21_286/a_572_375# 0.026009f
C7442 _147_ _435_/a_448_472# 0.001008f
C7443 _450_/a_2225_156# net6 0.001143f
C7444 FILLER_0_16_73/a_124_375# FILLER_0_17_72/a_124_375# 0.026339f
C7445 _004_ vss 0.115789f
C7446 net28 output29/a_224_472# 0.028512f
C7447 _144_ FILLER_0_18_107/a_1916_375# 0.003148f
C7448 result[4] result[9] 0.101112f
C7449 net28 _426_/a_36_151# 0.004878f
C7450 _432_/a_2560_156# net63 0.00227f
C7451 output42/a_224_472# net44 0.079084f
C7452 _019_ net21 0.065941f
C7453 _327_/a_244_68# _130_ 0.00117f
C7454 FILLER_0_4_123/a_36_472# _152_ 0.003937f
C7455 net16 FILLER_0_8_37/a_124_375# 0.010358f
C7456 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_124_375# 0.003228f
C7457 net39 _445_/a_1204_472# 0.002681f
C7458 _317_/a_36_113# _014_ 0.037134f
C7459 _015_ vdd 0.27747f
C7460 FILLER_0_15_116/a_124_375# net36 0.003055f
C7461 FILLER_0_5_72/a_484_472# trim_mask\[1\] 0.012321f
C7462 mask\[5\] output35/a_224_472# 0.003461f
C7463 FILLER_0_5_206/a_36_472# net37 0.009858f
C7464 net68 net49 0.607379f
C7465 _430_/a_2665_112# FILLER_0_15_212/a_1380_472# 0.021761f
C7466 _093_ FILLER_0_21_60/a_572_375# 0.011177f
C7467 _426_/a_3041_156# net64 0.001046f
C7468 _452_/a_836_156# net40 0.023204f
C7469 mask\[2\] FILLER_0_16_154/a_1380_472# 0.017868f
C7470 trim_mask\[4\] _241_/a_224_472# 0.009431f
C7471 _233_/a_36_160# net67 0.001315f
C7472 net25 _051_ 0.090798f
C7473 net34 result[6] 0.072393f
C7474 output8/a_224_472# cal_itt\[1\] 0.003894f
C7475 fanout64/a_36_160# _425_/a_2665_112# 0.005704f
C7476 _256_/a_244_497# calibrate 0.002421f
C7477 _057_ _311_/a_1212_473# 0.004869f
C7478 _104_ FILLER_0_23_274/a_124_375# 0.002159f
C7479 FILLER_0_22_86/a_932_472# _098_ 0.001442f
C7480 output36/a_224_472# _417_/a_2248_156# 0.023576f
C7481 _176_ _451_/a_36_151# 0.003176f
C7482 FILLER_0_17_72/a_36_472# _131_ 0.002672f
C7483 trim_mask\[1\] _160_ 0.051511f
C7484 result[8] _048_ 0.006006f
C7485 _065_ _064_ 0.007356f
C7486 vss FILLER_0_19_134/a_36_472# 0.005204f
C7487 _369_/a_36_68# _367_/a_36_68# 0.038188f
C7488 _153_ vss 0.256017f
C7489 _430_/a_36_151# mask\[2\] 0.016265f
C7490 FILLER_0_12_136/a_1468_375# vdd 0.026145f
C7491 FILLER_0_15_116/a_572_375# net70 0.050592f
C7492 FILLER_0_12_136/a_1020_375# vss 0.018233f
C7493 _116_ _162_ 0.00156f
C7494 FILLER_0_23_274/a_36_472# vdd 0.010289f
C7495 FILLER_0_23_274/a_124_375# vss 0.017196f
C7496 _230_/a_244_68# _070_ 0.001641f
C7497 net26 _423_/a_1000_472# 0.001338f
C7498 net64 FILLER_0_9_282/a_36_472# 0.031302f
C7499 result[7] FILLER_0_24_274/a_572_375# 0.006125f
C7500 FILLER_0_5_54/a_572_375# vss 0.002617f
C7501 FILLER_0_5_54/a_1020_375# vdd -0.014642f
C7502 _091_ _106_ 0.001188f
C7503 FILLER_0_4_197/a_1020_375# net59 0.008989f
C7504 FILLER_0_17_72/a_1468_375# net36 0.047507f
C7505 _068_ _152_ 0.006744f
C7506 _451_/a_2449_156# _040_ 0.004434f
C7507 _157_ _160_ 0.010231f
C7508 _430_/a_2560_156# net63 0.009628f
C7509 _442_/a_1000_472# vdd 0.003088f
C7510 FILLER_0_18_177/a_572_375# FILLER_0_20_177/a_484_472# 0.0027f
C7511 _356_/a_36_472# _438_/a_36_151# 0.004432f
C7512 _114_ _428_/a_2248_156# 0.004516f
C7513 mask\[9\] FILLER_0_20_87/a_36_472# 0.00596f
C7514 _321_/a_2590_472# _129_ 0.005391f
C7515 _242_/a_36_160# net47 0.028264f
C7516 _096_ _113_ 0.650985f
C7517 _035_ _167_ 0.01574f
C7518 mask\[3\] net64 0.002654f
C7519 _178_ _402_/a_1948_68# 0.00815f
C7520 FILLER_0_4_177/a_572_375# vss 0.054783f
C7521 FILLER_0_4_177/a_36_472# vdd 0.114788f
C7522 net41 _446_/a_2665_112# 0.004501f
C7523 FILLER_0_18_177/a_572_375# vdd 0.031241f
C7524 FILLER_0_18_177/a_124_375# vss 0.00364f
C7525 _036_ FILLER_0_3_54/a_36_472# 0.002156f
C7526 _449_/a_1308_423# _067_ 0.021042f
C7527 net79 FILLER_0_11_282/a_124_375# 0.002239f
C7528 net62 FILLER_0_11_282/a_36_472# 0.00149f
C7529 FILLER_0_12_20/a_572_375# vdd 0.013384f
C7530 _004_ _416_/a_2248_156# 0.001078f
C7531 _162_ _118_ 0.005444f
C7532 _095_ net14 0.043065f
C7533 FILLER_0_16_73/a_484_472# net15 0.001946f
C7534 FILLER_0_21_142/a_124_375# _140_ 0.016087f
C7535 fanout55/a_36_160# _095_ 0.00409f
C7536 _142_ vss 0.121933f
C7537 _412_/a_2665_112# vdd 0.014403f
C7538 _436_/a_2665_112# vss 0.007905f
C7539 FILLER_0_3_221/a_1380_472# vss 0.002804f
C7540 FILLER_0_4_99/a_36_472# net47 0.003903f
C7541 net73 FILLER_0_18_107/a_2364_375# 0.015484f
C7542 _093_ _131_ 0.254316f
C7543 _131_ _118_ 0.001685f
C7544 mask\[7\] FILLER_0_22_128/a_572_375# 0.01909f
C7545 net72 FILLER_0_20_31/a_124_375# 0.011347f
C7546 net75 _263_/a_224_472# 0.004396f
C7547 _257_/a_36_472# cal_itt\[3\] 0.136487f
C7548 _273_/a_36_68# FILLER_0_10_214/a_36_472# 0.003036f
C7549 net74 FILLER_0_13_100/a_36_472# 0.003924f
C7550 net27 net58 0.190417f
C7551 ctln[3] cal_itt\[0\] 0.002081f
C7552 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1468_375# 0.086635f
C7553 _439_/a_2665_112# vss 0.003954f
C7554 FILLER_0_22_128/a_1380_472# _433_/a_36_151# 0.001973f
C7555 FILLER_0_19_171/a_1380_472# FILLER_0_19_187/a_36_472# 0.013277f
C7556 _002_ FILLER_0_3_172/a_2364_375# 0.016984f
C7557 _444_/a_2248_156# FILLER_0_8_37/a_484_472# 0.013656f
C7558 _379_/a_36_472# _063_ 0.071695f
C7559 net36 _040_ 0.429029f
C7560 FILLER_0_15_150/a_124_375# vdd 0.026143f
C7561 _428_/a_1308_423# _043_ 0.024052f
C7562 _036_ _164_ 0.011115f
C7563 FILLER_0_21_28/a_1828_472# _424_/a_36_151# 0.001723f
C7564 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3260_375# 0.001597f
C7565 _445_/a_448_472# net49 0.00122f
C7566 net15 FILLER_0_21_60/a_572_375# 0.03167f
C7567 _077_ FILLER_0_6_231/a_124_375# 0.009235f
C7568 _335_/a_49_472# vdd 0.085394f
C7569 _221_/a_36_160# net40 0.002952f
C7570 _412_/a_36_151# net19 0.03393f
C7571 net79 FILLER_0_13_290/a_36_472# 0.038324f
C7572 _115_ _322_/a_848_380# 0.011372f
C7573 _313_/a_67_603# _227_/a_36_160# 0.032438f
C7574 _307_/a_234_472# _085_ 0.001966f
C7575 FILLER_0_16_57/a_124_375# FILLER_0_15_59/a_36_472# 0.001543f
C7576 net80 _019_ 0.265857f
C7577 net69 _152_ 0.002532f
C7578 _415_/a_2560_156# net64 0.066438f
C7579 _126_ net23 0.030487f
C7580 FILLER_0_12_136/a_1380_472# cal_count\[3\] 0.00383f
C7581 _072_ _121_ 0.041039f
C7582 _428_/a_36_151# _095_ 0.006658f
C7583 net58 _425_/a_2665_112# 0.069807f
C7584 fanout62/a_36_160# net64 0.052109f
C7585 net15 _440_/a_36_151# 0.016061f
C7586 FILLER_0_10_28/a_36_472# net40 0.020589f
C7587 state\[2\] FILLER_0_13_142/a_572_375# 0.007511f
C7588 _056_ _113_ 0.052362f
C7589 net53 FILLER_0_13_142/a_1468_375# 0.002334f
C7590 net57 FILLER_0_3_172/a_36_472# 0.001007f
C7591 _190_/a_36_160# _039_ 0.003926f
C7592 FILLER_0_16_73/a_124_375# _175_ 0.005727f
C7593 _308_/a_124_24# _439_/a_2665_112# 0.002245f
C7594 mask\[3\] _103_ 0.055796f
C7595 FILLER_0_24_274/a_1020_375# vss 0.003553f
C7596 _119_ FILLER_0_7_104/a_1468_375# 0.022368f
C7597 _448_/a_2248_156# _170_ 0.00254f
C7598 _448_/a_1000_472# _037_ 0.03564f
C7599 FILLER_0_12_28/a_124_375# vdd 0.040988f
C7600 FILLER_0_18_2/a_2364_375# vdd 0.002983f
C7601 vss output40/a_224_472# 0.002459f
C7602 _375_/a_36_68# _062_ 0.012855f
C7603 net31 _102_ 0.060034f
C7604 _437_/a_2248_156# _436_/a_36_151# 0.001837f
C7605 FILLER_0_22_128/a_1468_375# vss 0.006619f
C7606 _052_ FILLER_0_19_28/a_484_472# 0.003325f
C7607 _093_ net56 0.040124f
C7608 net71 FILLER_0_22_107/a_124_375# 0.018295f
C7609 _408_/a_1936_472# cal_count\[0\] 0.001434f
C7610 _207_/a_67_603# vss 0.00837f
C7611 output34/a_224_472# ctlp[1] 0.00277f
C7612 _019_ mask\[1\] 0.007797f
C7613 _086_ FILLER_0_11_142/a_572_375# 0.011726f
C7614 mask\[5\] ctlp[2] 0.104304f
C7615 _028_ _439_/a_448_472# 0.017606f
C7616 FILLER_0_13_65/a_124_375# net74 0.020091f
C7617 _441_/a_36_151# FILLER_0_3_78/a_36_472# 0.001723f
C7618 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1380_472# 0.013276f
C7619 _084_ vdd 0.134578f
C7620 _077_ FILLER_0_8_239/a_36_472# 0.001289f
C7621 _131_ _330_/a_224_472# 0.001186f
C7622 _087_ FILLER_0_3_172/a_932_472# 0.001947f
C7623 _086_ FILLER_0_7_104/a_572_375# 0.003137f
C7624 _420_/a_36_151# FILLER_0_23_290/a_124_375# 0.026277f
C7625 net61 net77 0.986569f
C7626 net82 FILLER_0_3_172/a_124_375# 0.011418f
C7627 FILLER_0_15_282/a_124_375# vss 0.004893f
C7628 FILLER_0_15_282/a_572_375# vdd 0.002928f
C7629 _120_ FILLER_0_9_72/a_484_472# 0.001645f
C7630 FILLER_0_17_38/a_124_375# vdd 0.01443f
C7631 _064_ _034_ 1.397143f
C7632 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_572_375# 0.086635f
C7633 FILLER_0_3_172/a_124_375# fanout57/a_36_113# 0.006548f
C7634 FILLER_0_7_59/a_572_375# trim_mask\[1\] 0.001548f
C7635 _127_ _321_/a_2034_472# 0.003159f
C7636 net15 _131_ 0.037758f
C7637 _415_/a_2665_112# FILLER_0_9_290/a_124_375# 0.001597f
C7638 net32 _419_/a_2665_112# 0.027035f
C7639 _087_ FILLER_0_5_181/a_36_472# 0.154469f
C7640 _057_ cal_count\[3\] 0.416063f
C7641 fanout80/a_36_113# FILLER_0_15_205/a_36_472# 0.010419f
C7642 input4/a_36_68# net59 0.003625f
C7643 _120_ _453_/a_2665_112# 0.002925f
C7644 FILLER_0_14_123/a_36_472# vdd 0.088525f
C7645 FILLER_0_14_123/a_124_375# vss 0.004985f
C7646 FILLER_0_6_47/a_2724_472# vss 0.020876f
C7647 FILLER_0_6_47/a_3172_472# vdd 0.002089f
C7648 net48 net37 0.081653f
C7649 FILLER_0_18_2/a_572_375# net44 0.072627f
C7650 _035_ vdd 0.215473f
C7651 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_124_375# 0.026339f
C7652 net56 net54 0.018493f
C7653 _250_/a_36_68# cal_count\[3\] 0.004136f
C7654 _070_ FILLER_0_5_136/a_124_375# 0.001083f
C7655 net57 FILLER_0_13_100/a_124_375# 0.012636f
C7656 net72 FILLER_0_19_28/a_572_375# 0.010026f
C7657 _143_ vss 0.02001f
C7658 FILLER_0_0_266/a_124_375# rstn 0.073089f
C7659 net20 FILLER_0_6_231/a_124_375# 0.060499f
C7660 _402_/a_1948_68# _401_/a_36_68# 0.012664f
C7661 output48/a_224_472# _079_ 0.003556f
C7662 FILLER_0_12_2/a_572_375# net6 0.058881f
C7663 FILLER_0_22_177/a_36_472# _434_/a_448_472# 0.012285f
C7664 FILLER_0_4_144/a_124_375# vdd 0.005512f
C7665 fanout78/a_36_113# _094_ 0.01312f
C7666 fanout56/a_36_113# net36 0.021321f
C7667 FILLER_0_13_212/a_1380_472# vss 0.010223f
C7668 _002_ net76 0.213703f
C7669 _105_ _293_/a_36_472# 0.004667f
C7670 _443_/a_36_151# _031_ 0.014344f
C7671 _443_/a_1308_423# net69 0.004128f
C7672 _032_ _442_/a_36_151# 0.005632f
C7673 FILLER_0_10_256/a_124_375# FILLER_0_10_247/a_124_375# 0.002036f
C7674 net26 FILLER_0_21_28/a_2812_375# 0.001905f
C7675 _116_ _076_ 0.008283f
C7676 _085_ _070_ 0.058787f
C7677 net34 _422_/a_1204_472# 0.001029f
C7678 _086_ FILLER_0_5_181/a_36_472# 0.013437f
C7679 _132_ _043_ 0.038747f
C7680 _276_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C7681 _446_/a_2560_156# net17 0.00101f
C7682 _402_/a_56_567# net47 0.026503f
C7683 vss FILLER_0_5_148/a_36_472# 0.029152f
C7684 _415_/a_448_472# vdd 0.005273f
C7685 ctln[2] rstn 0.017812f
C7686 net20 net60 0.033919f
C7687 FILLER_0_4_177/a_484_472# net76 0.006746f
C7688 output44/a_224_472# _452_/a_1353_112# 0.001321f
C7689 net2 fanout58/a_36_160# 0.010424f
C7690 _028_ _151_ 0.020076f
C7691 net55 FILLER_0_17_72/a_932_472# 0.024922f
C7692 _001_ net59 0.001439f
C7693 _105_ _108_ 0.548284f
C7694 FILLER_0_12_20/a_36_472# _450_/a_448_472# 0.058631f
C7695 FILLER_0_2_111/a_932_472# vss -0.001894f
C7696 FILLER_0_2_111/a_1380_472# vdd 0.002688f
C7697 fanout69/a_36_113# _371_/a_36_113# 0.259508f
C7698 FILLER_0_9_142/a_124_375# calibrate 0.001505f
C7699 _256_/a_1612_497# _076_ 0.001111f
C7700 _105_ net19 0.049611f
C7701 ctln[1] _073_ 0.001457f
C7702 net20 FILLER_0_8_239/a_36_472# 0.004483f
C7703 _440_/a_2248_156# vss 0.010006f
C7704 _440_/a_2665_112# vdd -0.002297f
C7705 en fanout59/a_36_160# 0.242369f
C7706 net15 FILLER_0_13_80/a_36_472# 0.001122f
C7707 _029_ _365_/a_244_472# 0.001956f
C7708 net18 _418_/a_1204_472# 0.01349f
C7709 _076_ _118_ 0.06281f
C7710 FILLER_0_24_63/a_36_472# vss 0.008178f
C7711 _448_/a_448_472# FILLER_0_3_172/a_572_375# 0.00123f
C7712 _448_/a_36_151# FILLER_0_3_172/a_1020_375# 0.001512f
C7713 net62 FILLER_0_15_235/a_572_375# 0.001315f
C7714 trim_mask\[2\] _381_/a_36_472# 0.034251f
C7715 _428_/a_36_151# _332_/a_36_472# 0.004432f
C7716 net63 FILLER_0_18_177/a_572_375# 0.004407f
C7717 FILLER_0_16_107/a_572_375# _040_ 0.001244f
C7718 net57 FILLER_0_16_154/a_1468_375# 0.217874f
C7719 FILLER_0_22_86/a_1468_375# _211_/a_36_160# 0.010334f
C7720 _219_/a_36_160# vdd 0.013125f
C7721 ctlp[8] _051_ 0.010337f
C7722 _345_/a_36_160# _145_ 0.001141f
C7723 _136_ vdd 1.020301f
C7724 FILLER_0_18_2/a_36_472# _452_/a_3129_107# 0.035307f
C7725 state\[1\] net23 0.075055f
C7726 net82 _443_/a_1204_472# 0.004056f
C7727 FILLER_0_21_28/a_2276_472# _012_ 0.023696f
C7728 _065_ _383_/a_36_472# 0.02518f
C7729 net57 _055_ 0.008619f
C7730 FILLER_0_16_89/a_124_375# _131_ 0.017319f
C7731 output38/a_224_472# _034_ 0.039873f
C7732 net38 _160_ 0.00247f
C7733 net70 FILLER_0_14_107/a_932_472# 0.008396f
C7734 net53 FILLER_0_14_107/a_1468_375# 0.001642f
C7735 FILLER_0_4_107/a_484_472# _031_ 0.002521f
C7736 output20/a_224_472# ctlp[2] 0.085373f
C7737 FILLER_0_12_136/a_572_375# _126_ 0.01289f
C7738 _277_/a_36_160# _102_ 0.061995f
C7739 net62 vdd 1.53102f
C7740 FILLER_0_1_266/a_484_472# net18 0.010423f
C7741 FILLER_0_1_266/a_572_375# net8 0.016292f
C7742 net27 FILLER_0_9_270/a_484_472# 0.023461f
C7743 _438_/a_796_472# vss 0.001171f
C7744 FILLER_0_13_142/a_124_375# vdd 0.02675f
C7745 fanout72/a_36_113# vss 0.053396f
C7746 ctlp[1] _419_/a_2248_156# 0.028734f
C7747 FILLER_0_0_96/a_36_472# vss 0.00344f
C7748 net35 _352_/a_49_472# 0.02594f
C7749 mask\[8\] _352_/a_257_69# 0.003259f
C7750 net73 FILLER_0_19_111/a_572_375# 0.04458f
C7751 mask\[5\] net21 0.212814f
C7752 net52 FILLER_0_5_72/a_1020_375# 0.00799f
C7753 fanout78/a_36_113# net78 0.004202f
C7754 cal_count\[2\] net40 0.313209f
C7755 FILLER_0_9_28/a_124_375# net47 0.006757f
C7756 output23/a_224_472# net23 0.122379f
C7757 FILLER_0_24_274/a_484_472# _420_/a_36_151# 0.002841f
C7758 _412_/a_1000_472# net59 0.00147f
C7759 cal_count\[3\] _310_/a_49_472# 0.00277f
C7760 net16 _182_ 0.05291f
C7761 _158_ _160_ 0.018681f
C7762 mask\[5\] FILLER_0_19_171/a_932_472# 0.007596f
C7763 FILLER_0_9_28/a_2276_472# net68 0.023299f
C7764 _176_ _182_ 0.008217f
C7765 FILLER_0_5_72/a_1020_375# net49 0.002208f
C7766 _311_/a_254_473# net21 0.003733f
C7767 _074_ _123_ 0.157299f
C7768 _016_ cal_count\[3\] 0.004588f
C7769 FILLER_0_16_107/a_124_375# net36 0.001706f
C7770 output29/a_224_472# output30/a_224_472# 0.005147f
C7771 net44 FILLER_0_15_2/a_124_375# 0.017852f
C7772 output19/a_224_472# _108_ 0.005075f
C7773 FILLER_0_15_2/a_572_375# vss 0.055203f
C7774 FILLER_0_15_2/a_36_472# vdd 0.104741f
C7775 FILLER_0_17_56/a_36_472# FILLER_0_18_53/a_484_472# 0.026657f
C7776 net57 _126_ 0.021705f
C7777 FILLER_0_4_107/a_1380_472# _152_ 0.001297f
C7778 _074_ _073_ 0.040339f
C7779 net4 net22 0.036966f
C7780 FILLER_0_19_28/a_484_472# net40 0.020293f
C7781 mask\[3\] mask\[2\] 0.077703f
C7782 output19/a_224_472# net19 0.030721f
C7783 FILLER_0_17_200/a_484_472# net22 0.020589f
C7784 fanout70/a_36_113# vdd 0.015969f
C7785 _450_/a_448_472# net40 0.00222f
C7786 _095_ FILLER_0_12_20/a_124_375# 0.001588f
C7787 _430_/a_796_472# net36 0.00117f
C7788 net66 _160_ 0.097885f
C7789 FILLER_0_21_125/a_572_375# _140_ 0.01659f
C7790 FILLER_0_20_177/a_1468_375# mask\[6\] 0.001162f
C7791 FILLER_0_6_177/a_36_472# vss 0.001617f
C7792 _073_ _076_ 0.011358f
C7793 FILLER_0_6_177/a_484_472# vdd 0.007991f
C7794 _091_ _098_ 1.501073f
C7795 net36 FILLER_0_15_235/a_484_472# 0.019725f
C7796 _028_ FILLER_0_5_72/a_932_472# 0.003042f
C7797 _376_/a_36_160# vss 0.03081f
C7798 FILLER_0_9_223/a_124_375# vss 0.009569f
C7799 _070_ _062_ 0.06973f
C7800 _072_ FILLER_0_7_233/a_124_375# 0.002279f
C7801 _341_/a_49_472# vss 0.003485f
C7802 _077_ FILLER_0_8_156/a_484_472# 0.006446f
C7803 _417_/a_1000_472# _006_ 0.026299f
C7804 FILLER_0_7_104/a_36_472# _131_ 0.002019f
C7805 FILLER_0_7_104/a_1468_375# _129_ 0.001165f
C7806 FILLER_0_7_146/a_36_472# _062_ 0.011622f
C7807 FILLER_0_9_28/a_572_375# _054_ 0.002983f
C7808 output43/a_224_472# vdd -0.032713f
C7809 ctln[1] FILLER_0_1_266/a_484_472# 0.002068f
C7810 _086_ _268_/a_245_68# 0.001044f
C7811 _432_/a_448_472# _137_ 0.008956f
C7812 FILLER_0_24_96/a_124_375# net25 0.008342f
C7813 FILLER_0_18_37/a_1380_472# vss 0.002042f
C7814 _250_/a_36_68# _427_/a_2665_112# 0.002152f
C7815 FILLER_0_4_49/a_124_375# trim_mask\[1\] 0.006676f
C7816 _335_/a_257_69# _043_ 0.001043f
C7817 cal net5 0.039735f
C7818 net75 _316_/a_1084_68# 0.001531f
C7819 _014_ _122_ 0.001529f
C7820 _429_/a_2248_156# vss 0.040729f
C7821 _429_/a_2665_112# vdd 0.010552f
C7822 FILLER_0_17_56/a_124_375# vss 0.00143f
C7823 FILLER_0_17_56/a_572_375# vdd 0.003489f
C7824 _000_ _253_/a_36_68# 0.005121f
C7825 FILLER_0_13_212/a_484_472# mask\[0\] 0.001794f
C7826 _014_ FILLER_0_7_233/a_124_375# 0.00143f
C7827 net19 FILLER_0_23_282/a_124_375# 0.001668f
C7828 output47/a_224_472# net38 0.082174f
C7829 _188_ _120_ 0.046757f
C7830 _316_/a_124_24# vss 0.00516f
C7831 _316_/a_848_380# vdd 0.048727f
C7832 FILLER_0_19_195/a_36_472# net21 0.009159f
C7833 fanout80/a_36_113# _139_ 0.009968f
C7834 net79 _416_/a_1000_472# 0.024811f
C7835 net68 _165_ 0.002748f
C7836 _044_ result[3] 0.00251f
C7837 net53 vdd 0.78288f
C7838 _017_ vss 0.022624f
C7839 net26 _424_/a_796_472# 0.006496f
C7840 _186_ cal_count\[1\] 0.003341f
C7841 FILLER_0_7_195/a_124_375# _163_ 0.001308f
C7842 _453_/a_36_151# _042_ 0.035846f
C7843 _043_ net40 0.031043f
C7844 _390_/a_36_68# _172_ 0.033476f
C7845 FILLER_0_3_54/a_124_375# _160_ 0.004602f
C7846 FILLER_0_20_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001543f
C7847 FILLER_0_4_197/a_572_375# net22 0.016547f
C7848 en net5 0.892091f
C7849 _386_/a_124_24# vdd 0.014293f
C7850 mask\[5\] mask\[7\] 0.014384f
C7851 FILLER_0_8_138/a_124_375# _077_ 0.007238f
C7852 FILLER_0_18_2/a_3260_375# net55 0.004262f
C7853 _412_/a_2248_156# vdd 0.005671f
C7854 net27 calibrate 0.017426f
C7855 _260_/a_36_68# vdd 0.011119f
C7856 _119_ _372_/a_170_472# 0.003159f
C7857 _090_ _060_ 0.396493f
C7858 FILLER_0_19_171/a_124_375# vdd -0.009473f
C7859 FILLER_0_22_86/a_1468_375# net71 0.010224f
C7860 net41 net38 0.059214f
C7861 net15 FILLER_0_13_72/a_124_375# 0.006403f
C7862 _451_/a_448_472# net14 0.04399f
C7863 net36 _437_/a_36_151# 0.002694f
C7864 FILLER_0_18_2/a_3172_472# FILLER_0_18_37/a_36_472# 0.002765f
C7865 FILLER_0_18_2/a_36_472# vss 0.001872f
C7866 net27 FILLER_0_10_256/a_124_375# 0.006216f
C7867 FILLER_0_10_107/a_36_472# vss 0.003894f
C7868 FILLER_0_10_107/a_484_472# vdd 0.034172f
C7869 _069_ _315_/a_36_68# 0.002242f
C7870 net46 net40 0.254778f
C7871 mask\[1\] FILLER_0_15_228/a_124_375# 0.013558f
C7872 _091_ _070_ 0.162632f
C7873 FILLER_0_11_282/a_36_472# _416_/a_1308_423# 0.001295f
C7874 net2 net18 0.030437f
C7875 _108_ mask\[6\] 0.032481f
C7876 _452_/a_1353_112# vdd 0.008539f
C7877 trimb[3] net43 0.221036f
C7878 _091_ _432_/a_36_151# 0.054497f
C7879 _003_ net37 0.046745f
C7880 net67 FILLER_0_12_20/a_36_472# 0.054453f
C7881 mask\[5\] net80 0.036014f
C7882 _091_ FILLER_0_15_180/a_124_375# 0.001415f
C7883 _104_ fanout63/a_36_160# 0.007014f
C7884 _144_ _354_/a_49_472# 0.03742f
C7885 net68 net40 0.036106f
C7886 _320_/a_1792_472# net79 0.002091f
C7887 trim[4] vdd 0.198218f
C7888 net4 vdd 1.218939f
C7889 _211_/a_36_160# net71 0.035804f
C7890 FILLER_0_18_177/a_2276_472# net21 0.01016f
C7891 net60 _009_ 0.006086f
C7892 mask\[3\] FILLER_0_16_154/a_484_472# 0.002067f
C7893 output18/a_224_472# ctlp[1] 0.039734f
C7894 FILLER_0_17_200/a_484_472# vdd 0.008335f
C7895 fanout63/a_36_160# vss 0.008974f
C7896 _164_ _166_ 0.002368f
C7897 _425_/a_2665_112# calibrate 0.029064f
C7898 _104_ _291_/a_36_160# 0.006129f
C7899 _081_ _123_ 0.007811f
C7900 _248_/a_36_68# vss 0.027935f
C7901 FILLER_0_4_197/a_124_375# _079_ 0.004772f
C7902 _230_/a_244_68# net21 0.00165f
C7903 _067_ FILLER_0_13_80/a_124_375# 0.001857f
C7904 _274_/a_3368_68# _069_ 0.001414f
C7905 _165_ net67 0.045827f
C7906 FILLER_0_8_107/a_36_472# FILLER_0_9_105/a_124_375# 0.001684f
C7907 _012_ FILLER_0_21_60/a_572_375# 0.011991f
C7908 _440_/a_36_151# net47 0.013626f
C7909 _073_ _081_ 0.046537f
C7910 _291_/a_36_160# vss 0.012222f
C7911 result[5] _418_/a_448_472# 0.007308f
C7912 _417_/a_2665_112# vss 0.002571f
C7913 _417_/a_2560_156# vdd 0.001658f
C7914 FILLER_0_14_107/a_124_375# vdd 0.013327f
C7915 FILLER_0_24_130/a_36_472# ctlp[7] 0.012298f
C7916 FILLER_0_9_72/a_36_472# vdd 0.109576f
C7917 FILLER_0_9_72/a_1468_375# vss 0.013085f
C7918 _110_ _098_ 0.09704f
C7919 FILLER_0_10_78/a_36_472# FILLER_0_9_72/a_572_375# 0.001543f
C7920 _420_/a_36_151# FILLER_0_23_282/a_124_375# 0.059049f
C7921 net41 _424_/a_36_151# 0.00413f
C7922 _182_ _041_ 0.08834f
C7923 net41 net66 0.08664f
C7924 _421_/a_2665_112# _419_/a_2665_112# 0.002588f
C7925 _116_ _090_ 0.122467f
C7926 FILLER_0_5_72/a_932_472# net47 0.003953f
C7927 _095_ FILLER_0_14_123/a_124_375# 0.014486f
C7928 net41 _067_ 0.033696f
C7929 FILLER_0_16_73/a_572_375# net55 0.015207f
C7930 _453_/a_2248_156# vdd 0.010767f
C7931 _127_ FILLER_0_11_142/a_36_472# 0.004538f
C7932 _311_/a_1660_473# vdd 0.001435f
C7933 FILLER_0_22_128/a_3172_472# _146_ 0.008065f
C7934 cal_count\[2\] FILLER_0_15_2/a_484_472# 0.015036f
C7935 _015_ _426_/a_1204_472# 0.008883f
C7936 _073_ net65 0.775972f
C7937 net22 _047_ 0.132529f
C7938 net23 _160_ 0.030085f
C7939 net57 state\[1\] 0.154183f
C7940 ctln[1] net2 0.126801f
C7941 FILLER_0_10_78/a_1468_375# _114_ 0.01836f
C7942 _308_/a_124_24# FILLER_0_9_72/a_1468_375# 0.007188f
C7943 _187_ net41 0.002046f
C7944 net54 FILLER_0_22_86/a_1020_375# 0.001597f
C7945 _136_ FILLER_0_16_154/a_572_375# 0.003842f
C7946 _196_/a_36_160# _045_ 0.036714f
C7947 _162_ net47 0.004104f
C7948 _088_ FILLER_0_3_221/a_124_375# 0.002378f
C7949 _098_ _437_/a_2665_112# 0.003567f
C7950 net62 _283_/a_36_472# 0.002309f
C7951 valid net18 0.03851f
C7952 fanout60/a_36_160# _417_/a_36_151# 0.062739f
C7953 _352_/a_49_472# vdd 0.077542f
C7954 trimb[1] FILLER_0_20_2/a_124_375# 0.003431f
C7955 output40/a_224_472# output41/a_224_472# 0.292611f
C7956 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_36_472# 0.002765f
C7957 net67 net40 0.886781f
C7958 net54 FILLER_0_22_128/a_1828_472# 0.009504f
C7959 net35 _213_/a_255_603# 0.001597f
C7960 _301_/a_36_472# _051_ 0.001277f
C7961 _308_/a_848_380# _070_ 0.033275f
C7962 _430_/a_1000_472# vss 0.001626f
C7963 FILLER_0_4_197/a_572_375# vdd 0.002455f
C7964 _414_/a_2665_112# _053_ 0.032254f
C7965 _000_ _079_ 0.032884f
C7966 FILLER_0_5_128/a_484_472# _152_ 0.002283f
C7967 output27/a_224_472# net5 0.008663f
C7968 net81 FILLER_0_15_212/a_484_472# 0.00169f
C7969 _118_ _090_ 0.005469f
C7970 mask\[0\] _429_/a_1000_472# 0.020553f
C7971 _448_/a_2665_112# net59 0.005948f
C7972 _270_/a_36_472# _079_ 0.036715f
C7973 _077_ _255_/a_224_552# 0.025141f
C7974 _096_ FILLER_0_14_181/a_124_375# 0.002455f
C7975 _005_ vss 0.01812f
C7976 _005_ _192_/a_255_603# 0.001058f
C7977 _027_ _438_/a_796_472# 0.031292f
C7978 _150_ _438_/a_1204_472# 0.003696f
C7979 FILLER_0_3_172/a_1468_375# net22 0.012895f
C7980 net4 net9 0.008183f
C7981 FILLER_0_18_53/a_572_375# vdd 0.018416f
C7982 _094_ _418_/a_1308_423# 0.029276f
C7983 _394_/a_728_93# FILLER_0_15_72/a_572_375# 0.02852f
C7984 _094_ _006_ 0.090405f
C7985 _052_ _424_/a_2248_156# 0.005116f
C7986 _285_/a_36_472# mask\[2\] 0.002447f
C7987 FILLER_0_16_57/a_1468_375# _131_ 0.015859f
C7988 net34 FILLER_0_22_177/a_1020_375# 0.006974f
C7989 FILLER_0_18_107/a_2364_375# _433_/a_36_151# 0.002106f
C7990 _292_/a_36_160# _098_ 0.048643f
C7991 _412_/a_1308_423# net58 0.037719f
C7992 _412_/a_448_472# net1 0.035155f
C7993 _103_ _094_ 0.280781f
C7994 FILLER_0_4_107/a_484_472# _157_ 0.027364f
C7995 _151_ _154_ 0.108571f
C7996 net74 _390_/a_244_472# 0.001317f
C7997 _445_/a_448_472# net40 0.044285f
C7998 cal_itt\[2\] _083_ 0.10423f
C7999 FILLER_0_5_128/a_572_375# _081_ 0.023853f
C8000 _053_ FILLER_0_6_47/a_124_375# 0.002541f
C8001 output20/a_224_472# mask\[7\] 0.024731f
C8002 FILLER_0_21_28/a_484_472# net40 0.022617f
C8003 _292_/a_36_160# _205_/a_36_160# 0.105676f
C8004 _093_ FILLER_0_17_72/a_2812_375# 0.019521f
C8005 net70 FILLER_0_13_100/a_36_472# 0.00585f
C8006 _320_/a_36_472# net21 0.025762f
C8007 net79 _043_ 0.393702f
C8008 FILLER_0_10_78/a_1468_375# _176_ 0.013408f
C8009 FILLER_0_8_263/a_36_472# net64 0.00399f
C8010 net75 vss 0.662689f
C8011 net1 net19 0.024768f
C8012 FILLER_0_13_142/a_572_375# _043_ 0.009328f
C8013 FILLER_0_20_177/a_1020_375# vdd 0.005483f
C8014 _114_ FILLER_0_10_94/a_572_375# 0.008375f
C8015 net64 FILLER_0_14_235/a_572_375# 0.008689f
C8016 _098_ net14 0.061285f
C8017 mask\[8\] _423_/a_2248_156# 0.001648f
C8018 net62 _069_ 0.010033f
C8019 FILLER_0_21_125/a_124_375# _098_ 0.006462f
C8020 _176_ _040_ 0.272465f
C8021 net16 _447_/a_448_472# 0.063057f
C8022 _398_/a_36_113# vdd 0.030449f
C8023 FILLER_0_8_127/a_124_375# _119_ 0.013315f
C8024 fanout72/a_36_113# _095_ 0.001842f
C8025 _000_ cal_itt\[1\] 0.012692f
C8026 FILLER_0_24_63/a_36_472# output26/a_224_472# 0.023414f
C8027 FILLER_0_17_226/a_36_472# _104_ 0.013926f
C8028 _429_/a_36_151# FILLER_0_15_212/a_36_472# 0.001723f
C8029 _426_/a_36_151# _425_/a_36_151# 0.006252f
C8030 FILLER_0_20_15/a_1020_375# vdd 0.005198f
C8031 _086_ _119_ 0.419383f
C8032 net65 FILLER_0_1_266/a_484_472# 0.004635f
C8033 output21/a_224_472# _108_ 0.005356f
C8034 _422_/a_36_151# vdd 0.177717f
C8035 _384_/a_224_472# vss 0.004801f
C8036 FILLER_0_17_226/a_36_472# vss 0.007552f
C8037 cal_count\[2\] _452_/a_1040_527# 0.002003f
C8038 _432_/a_2248_156# net21 0.002329f
C8039 net20 FILLER_0_16_241/a_36_472# 0.001528f
C8040 FILLER_0_5_212/a_36_472# _081_ 0.01062f
C8041 _441_/a_1308_423# vdd 0.002837f
C8042 _441_/a_448_472# vss 0.025073f
C8043 _131_ net74 0.227843f
C8044 _412_/a_2560_156# net58 0.005111f
C8045 _233_/a_36_160# _033_ 0.017573f
C8046 vdd _047_ 0.175913f
C8047 net69 _369_/a_36_68# 0.008024f
C8048 _031_ _369_/a_244_472# 0.002741f
C8049 net55 _424_/a_448_472# 0.005273f
C8050 trim_val\[2\] _446_/a_2665_112# 0.012621f
C8051 net20 _413_/a_2248_156# 0.002515f
C8052 _288_/a_224_472# net19 0.002252f
C8053 FILLER_0_16_57/a_1380_472# _394_/a_728_93# 0.001627f
C8054 _413_/a_1000_472# net65 0.02866f
C8055 _058_ FILLER_0_9_105/a_36_472# 0.011426f
C8056 _326_/a_36_160# _086_ 0.063565f
C8057 FILLER_0_2_111/a_124_375# _154_ 0.004032f
C8058 _077_ _392_/a_36_68# 0.055912f
C8059 net52 _442_/a_2560_156# 0.008682f
C8060 FILLER_0_18_177/a_3172_472# vss 0.002639f
C8061 output36/a_224_472# output29/a_224_472# 0.007726f
C8062 mask\[4\] FILLER_0_19_155/a_572_375# 0.020261f
C8063 _005_ _416_/a_2248_156# 0.036714f
C8064 _176_ FILLER_0_10_94/a_572_375# 0.011743f
C8065 _431_/a_1308_423# _137_ 0.008805f
C8066 _441_/a_1000_472# _168_ 0.036305f
C8067 _058_ vdd 0.511536f
C8068 _356_/a_36_472# mask\[9\] 0.047632f
C8069 ctlp[1] _421_/a_1000_472# 0.007039f
C8070 FILLER_0_7_162/a_36_472# vss 0.006392f
C8071 _021_ vdd 0.022473f
C8072 FILLER_0_17_142/a_572_375# _137_ 0.006974f
C8073 FILLER_0_20_31/a_124_375# vdd 0.04619f
C8074 fanout77/a_36_113# vdd 0.032109f
C8075 FILLER_0_3_172/a_1468_375# vdd 0.045181f
C8076 _129_ _372_/a_170_472# 0.001985f
C8077 FILLER_0_15_290/a_124_375# output30/a_224_472# 0.02894f
C8078 _431_/a_1288_156# net73 0.001033f
C8079 _070_ net14 0.536953f
C8080 _079_ fanout75/a_36_113# 0.059598f
C8081 net16 _444_/a_448_472# 0.038803f
C8082 FILLER_0_4_123/a_124_375# trim_mask\[4\] 0.004312f
C8083 net54 _145_ 0.087336f
C8084 cal_count\[3\] _278_/a_36_160# 0.008398f
C8085 _147_ _207_/a_67_603# 0.001123f
C8086 _423_/a_36_151# FILLER_0_23_44/a_484_472# 0.001723f
C8087 net62 net28 0.05491f
C8088 net82 FILLER_0_2_171/a_36_472# 0.001777f
C8089 net26 _052_ 0.100927f
C8090 _115_ FILLER_0_9_72/a_1380_472# 0.007262f
C8091 _098_ FILLER_0_15_212/a_932_472# 0.011837f
C8092 FILLER_0_4_123/a_124_375# net47 0.011322f
C8093 vdd _416_/a_1308_423# 0.002623f
C8094 vss _416_/a_448_472# 0.004806f
C8095 FILLER_0_7_104/a_1468_375# _152_ 0.009263f
C8096 _422_/a_1308_423# _108_ 0.019345f
C8097 _412_/a_36_151# fanout81/a_36_160# 0.001725f
C8098 cal_count\[3\] vss 1.35143f
C8099 _033_ net49 0.003904f
C8100 _178_ cal_count\[3\] 0.002061f
C8101 FILLER_0_17_200/a_484_472# net63 0.003767f
C8102 net52 fanout74/a_36_113# 0.001514f
C8103 net34 output23/a_224_472# 0.021474f
C8104 FILLER_0_11_64/a_124_375# _120_ 0.004514f
C8105 _059_ vss 0.714648f
C8106 FILLER_0_19_47/a_484_472# _012_ 0.001667f
C8107 _092_ _276_/a_36_160# 0.06772f
C8108 _017_ _095_ 0.002789f
C8109 _098_ _434_/a_1000_472# 0.00725f
C8110 net15 _029_ 0.111797f
C8111 trim_mask\[4\] _170_ 0.09738f
C8112 net74 FILLER_0_13_80/a_36_472# 0.00679f
C8113 _295_/a_244_68# _107_ 0.00123f
C8114 FILLER_0_14_91/a_572_375# _136_ 0.049763f
C8115 _053_ _359_/a_36_488# 0.015831f
C8116 _131_ _154_ 0.019221f
C8117 net47 _170_ 0.010131f
C8118 _389_/a_36_148# vdd 0.039639f
C8119 _117_ _060_ 0.149558f
C8120 net79 FILLER_0_12_236/a_124_375# 0.010367f
C8121 _434_/a_36_151# _023_ 0.035162f
C8122 net10 net8 0.003331f
C8123 _089_ vss 0.018272f
C8124 FILLER_0_4_49/a_124_375# net66 0.017584f
C8125 fanout58/a_36_160# cal_itt\[1\] 0.010654f
C8126 output28/a_224_472# FILLER_0_11_282/a_124_375# 0.002977f
C8127 _074_ net47 0.012724f
C8128 net55 fanout55/a_36_160# 0.028425f
C8129 _132_ _428_/a_1204_472# 0.025555f
C8130 _128_ _055_ 1.887595f
C8131 ctlp[3] _422_/a_2665_112# 0.001024f
C8132 _077_ _120_ 0.205715f
C8133 trim_mask\[4\] _076_ 0.001824f
C8134 ctln[6] _037_ 0.031407f
C8135 FILLER_0_4_197/a_932_472# net82 0.001826f
C8136 output14/a_224_472# FILLER_0_0_130/a_36_472# 0.023414f
C8137 trim[0] _446_/a_448_472# 0.007307f
C8138 _030_ FILLER_0_3_78/a_36_472# 0.007376f
C8139 net49 FILLER_0_3_78/a_572_375# 0.066078f
C8140 _069_ net4 0.07542f
C8141 _055_ _311_/a_692_473# 0.003127f
C8142 FILLER_0_17_200/a_484_472# _069_ 0.001396f
C8143 _076_ net47 0.00115f
C8144 net2 net65 0.035908f
C8145 _009_ FILLER_0_23_290/a_124_375# 0.002666f
C8146 _320_/a_1120_472# vdd 0.001676f
C8147 trimb[2] vss 0.102375f
C8148 net50 FILLER_0_6_79/a_36_472# 0.001614f
C8149 _213_/a_67_603# vss 0.019344f
C8150 _431_/a_2248_156# net36 0.001441f
C8151 net82 FILLER_0_3_172/a_3172_472# 0.007677f
C8152 FILLER_0_4_185/a_124_375# _272_/a_36_472# 0.001781f
C8153 _119_ _313_/a_67_603# 0.015457f
C8154 _432_/a_2248_156# net80 0.059406f
C8155 _431_/a_36_151# FILLER_0_16_115/a_36_472# 0.004847f
C8156 output29/a_224_472# FILLER_0_14_263/a_36_472# 0.0323f
C8157 FILLER_0_4_123/a_124_375# net74 0.002449f
C8158 net20 _256_/a_1164_497# 0.001462f
C8159 _074_ FILLER_0_5_172/a_124_375# 0.068565f
C8160 FILLER_0_22_86/a_484_472# FILLER_0_23_88/a_124_375# 0.001684f
C8161 FILLER_0_3_172/a_2276_472# net65 0.001777f
C8162 output45/a_224_472# net45 0.019483f
C8163 _111_ _110_ 0.00195f
C8164 net55 _404_/a_36_472# 0.001746f
C8165 _070_ FILLER_0_11_109/a_36_472# 0.001091f
C8166 net62 net77 0.122747f
C8167 _128_ _126_ 0.008298f
C8168 _094_ mask\[2\] 0.089828f
C8169 _115_ FILLER_0_9_105/a_36_472# 0.004013f
C8170 net60 net33 0.008865f
C8171 _443_/a_2665_112# vss 0.007913f
C8172 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_572_375# 0.026339f
C8173 net27 mask\[0\] 0.067038f
C8174 FILLER_0_5_164/a_36_472# _066_ 0.00611f
C8175 FILLER_0_16_89/a_572_375# FILLER_0_17_72/a_2364_375# 0.026339f
C8176 _123_ FILLER_0_7_233/a_36_472# 0.002812f
C8177 _228_/a_36_68# _090_ 0.018462f
C8178 FILLER_0_12_220/a_124_375# _248_/a_36_68# 0.005308f
C8179 FILLER_0_9_223/a_36_472# _076_ 0.00146f
C8180 FILLER_0_7_162/a_124_375# vss 0.018732f
C8181 net17 _164_ 0.007595f
C8182 calibrate _062_ 2.032477f
C8183 _432_/a_2248_156# mask\[1\] 0.002293f
C8184 _115_ vdd 0.455713f
C8185 FILLER_0_19_28/a_572_375# vdd 0.034691f
C8186 _426_/a_36_151# FILLER_0_9_270/a_36_472# 0.008172f
C8187 _446_/a_796_472# net66 0.002296f
C8188 trim_val\[1\] _164_ 0.100504f
C8189 cal_count\[3\] _373_/a_438_68# 0.003743f
C8190 mask\[4\] mask\[3\] 1.118454f
C8191 ctlp[1] net18 0.088706f
C8192 _415_/a_2248_156# vss 0.00818f
C8193 trimb[0] vdd 0.10929f
C8194 FILLER_0_16_57/a_484_472# net55 0.001797f
C8195 _425_/a_448_472# FILLER_0_8_247/a_932_472# 0.012285f
C8196 FILLER_0_14_181/a_124_375# _138_ 0.001663f
C8197 _155_ FILLER_0_6_90/a_572_375# 0.001562f
C8198 _086_ _130_ 0.008816f
C8199 _062_ net21 0.025648f
C8200 net63 FILLER_0_20_177/a_1020_375# 0.005919f
C8201 _032_ _031_ 0.013851f
C8202 _070_ FILLER_0_8_156/a_124_375# 0.004329f
C8203 _086_ _161_ 0.077837f
C8204 net57 _428_/a_2560_156# 0.010877f
C8205 result[2] net79 0.077934f
C8206 output34/a_224_472# _199_/a_36_160# 0.003531f
C8207 _177_ _131_ 0.058938f
C8208 _118_ _117_ 0.032074f
C8209 net60 FILLER_0_17_282/a_124_375# 0.039003f
C8210 _214_/a_36_160# FILLER_0_23_88/a_124_375# 0.005398f
C8211 _238_/a_67_603# net14 0.004718f
C8212 _253_/a_36_68# _074_ 0.026327f
C8213 net56 FILLER_0_19_155/a_36_472# 0.00611f
C8214 mask\[4\] FILLER_0_19_187/a_36_472# 0.004669f
C8215 net81 cal_itt\[0\] 0.001048f
C8216 FILLER_0_15_72/a_484_472# cal_count\[1\] 0.013337f
C8217 FILLER_0_4_123/a_124_375# _159_ 0.023643f
C8218 valid net65 0.074257f
C8219 FILLER_0_14_91/a_572_375# net53 0.063988f
C8220 FILLER_0_8_127/a_124_375# _129_ 0.056784f
C8221 net36 state\[1\] 0.004105f
C8222 _440_/a_36_151# FILLER_0_6_47/a_1828_472# 0.001512f
C8223 FILLER_0_7_72/a_484_472# net52 0.049487f
C8224 _083_ _265_/a_224_472# 0.003404f
C8225 FILLER_0_17_72/a_1828_472# vss 0.001443f
C8226 FILLER_0_17_72/a_2276_472# vdd 0.001409f
C8227 _181_ _402_/a_718_527# 0.00461f
C8228 _086_ _129_ 0.051553f
C8229 _255_/a_224_552# cal_itt\[3\] 0.003266f
C8230 FILLER_0_22_86/a_124_375# net14 0.003962f
C8231 FILLER_0_9_223/a_572_375# net4 0.02077f
C8232 _419_/a_36_151# vdd -0.110366f
C8233 FILLER_0_12_20/a_484_472# _039_ 0.006288f
C8234 FILLER_0_16_89/a_1468_375# _040_ 0.004985f
C8235 _396_/a_224_472# net36 0.00114f
C8236 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2724_472# 0.026657f
C8237 FILLER_0_3_78/a_484_472# _164_ 0.05311f
C8238 FILLER_0_6_239/a_124_375# net76 0.001286f
C8239 _132_ FILLER_0_17_104/a_932_472# 0.006091f
C8240 trim_mask\[4\] _081_ 0.111668f
C8241 _427_/a_2665_112# vss 0.01229f
C8242 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_36_472# 0.026657f
C8243 net19 _420_/a_448_472# 0.05745f
C8244 FILLER_0_17_142/a_36_472# FILLER_0_19_142/a_124_375# 0.001512f
C8245 ctln[9] vdd 0.221231f
C8246 _372_/a_2034_472# _076_ 0.007461f
C8247 _372_/a_170_472# _068_ 0.037034f
C8248 net74 FILLER_0_13_72/a_124_375# 0.014594f
C8249 _081_ net47 1.302193f
C8250 _269_/a_36_472# _078_ 0.033601f
C8251 _257_/a_36_472# vdd -0.001779f
C8252 _190_/a_36_160# vdd 0.031799f
C8253 output15/a_224_472# net15 0.028578f
C8254 FILLER_0_1_204/a_124_375# net59 0.00999f
C8255 _412_/a_448_472# net76 0.026446f
C8256 net76 FILLER_0_3_172/a_1916_375# 0.019901f
C8257 _017_ _332_/a_36_472# 0.033837f
C8258 FILLER_0_21_206/a_36_472# vss 0.004971f
C8259 _321_/a_1194_69# vss 0.0011f
C8260 en_co_clk net74 0.039096f
C8261 net26 net40 0.001136f
C8262 result[9] _420_/a_2560_156# 0.002295f
C8263 net76 net19 0.02061f
C8264 FILLER_0_6_90/a_572_375# _163_ 0.007844f
C8265 net39 _444_/a_1000_472# 0.001323f
C8266 FILLER_0_4_152/a_124_375# vdd -0.001403f
C8267 FILLER_0_4_49/a_572_375# net47 0.00654f
C8268 mask\[5\] output18/a_224_472# 0.00133f
C8269 mask\[7\] _435_/a_448_472# 0.064472f
C8270 FILLER_0_8_138/a_36_472# _059_ 0.02252f
C8271 _412_/a_36_151# _265_/a_244_68# 0.072351f
C8272 _115_ _135_ 0.004345f
C8273 _394_/a_1336_472# cal_count\[1\] 0.018116f
C8274 _091_ net21 0.030022f
C8275 net55 _217_/a_36_160# 0.001311f
C8276 _091_ _333_/a_36_160# 0.031262f
C8277 cal_count\[3\] _071_ 0.214649f
C8278 net57 _374_/a_36_68# 0.001052f
C8279 net22 FILLER_0_18_209/a_572_375# 0.005202f
C8280 net25 FILLER_0_22_86/a_572_375# 0.002444f
C8281 _320_/a_36_472# mask\[0\] 0.001026f
C8282 cal_itt\[1\] net18 0.026586f
C8283 _069_ _047_ 0.001975f
C8284 FILLER_0_5_128/a_572_375# _163_ 0.007391f
C8285 _091_ FILLER_0_19_171/a_932_472# 0.002509f
C8286 _443_/a_2665_112# FILLER_0_2_165/a_36_472# 0.007491f
C8287 _149_ vdd 0.379674f
C8288 FILLER_0_2_171/a_124_375# net59 0.006603f
C8289 _053_ _372_/a_3662_472# 0.002006f
C8290 net23 FILLER_0_22_128/a_1380_472# 0.0019f
C8291 net80 _435_/a_448_472# 0.005274f
C8292 result[2] FILLER_0_13_290/a_124_375# 0.015011f
C8293 FILLER_0_18_139/a_124_375# vss 0.006869f
C8294 FILLER_0_18_139/a_572_375# vdd 0.004039f
C8295 mask\[0\] FILLER_0_14_235/a_36_472# 0.287093f
C8296 _408_/a_728_93# _067_ 0.006262f
C8297 FILLER_0_9_72/a_1020_375# _439_/a_36_151# 0.059049f
C8298 net78 _420_/a_2248_156# 0.001534f
C8299 _093_ FILLER_0_18_107/a_2812_375# 0.00626f
C8300 _036_ _384_/a_224_472# 0.001921f
C8301 FILLER_0_5_72/a_1468_375# _440_/a_2665_112# 0.001077f
C8302 _121_ net23 0.078786f
C8303 FILLER_0_15_282/a_572_375# output30/a_224_472# 0.029138f
C8304 _077_ FILLER_0_9_72/a_932_472# 0.006408f
C8305 net19 _419_/a_1308_423# 0.056469f
C8306 FILLER_0_0_130/a_36_472# vdd 0.050082f
C8307 FILLER_0_0_130/a_124_375# vss 0.018073f
C8308 FILLER_0_24_96/a_36_472# net24 0.028193f
C8309 FILLER_0_8_107/a_36_472# _077_ 0.007552f
C8310 ctln[2] cal 0.009784f
C8311 _233_/a_36_160# _444_/a_36_151# 0.032942f
C8312 net74 _081_ 0.093806f
C8313 _430_/a_36_151# _138_ 0.001123f
C8314 _187_ _408_/a_728_93# 0.002598f
C8315 FILLER_0_1_204/a_36_472# net21 0.076466f
C8316 _077_ _453_/a_2560_156# 0.001286f
C8317 _004_ net58 0.00116f
C8318 _106_ fanout63/a_36_160# 0.00715f
C8319 _105_ _009_ 0.01731f
C8320 net71 _437_/a_1000_472# 0.014459f
C8321 _155_ FILLER_0_7_104/a_36_472# 0.005042f
C8322 _435_/a_1000_472# vdd 0.032539f
C8323 _136_ _451_/a_36_151# 0.043941f
C8324 net38 _444_/a_796_472# 0.002641f
C8325 _119_ _061_ 0.132725f
C8326 state\[2\] _225_/a_36_160# 0.037565f
C8327 _291_/a_36_160# _106_ 0.054237f
C8328 FILLER_0_20_87/a_36_472# _438_/a_1308_423# 0.010224f
C8329 _089_ FILLER_0_5_198/a_36_472# 0.001314f
C8330 net38 FILLER_0_8_24/a_36_472# 0.015829f
C8331 _103_ _418_/a_2248_156# 0.012186f
C8332 _443_/a_36_151# net23 0.012359f
C8333 _449_/a_2665_112# en_co_clk 0.002966f
C8334 FILLER_0_18_76/a_36_472# vdd 0.014249f
C8335 FILLER_0_18_76/a_572_375# vss 0.007413f
C8336 ctln[2] en 0.001355f
C8337 _079_ _074_ 0.025058f
C8338 _134_ FILLER_0_9_105/a_36_472# 0.004375f
C8339 net33 _434_/a_2665_112# 0.001043f
C8340 _076_ FILLER_0_3_221/a_484_472# 0.001225f
C8341 FILLER_0_10_78/a_124_375# _120_ 0.006134f
C8342 _392_/a_36_68# _039_ 0.001522f
C8343 _372_/a_170_472# _152_ 0.037088f
C8344 _020_ vdd 0.194776f
C8345 FILLER_0_9_28/a_1020_375# _054_ 0.002273f
C8346 FILLER_0_10_37/a_124_375# _453_/a_36_151# 0.017882f
C8347 cal_count\[3\] _095_ 0.06065f
C8348 FILLER_0_5_117/a_36_472# net47 0.005919f
C8349 _086_ _056_ 0.043494f
C8350 _137_ FILLER_0_17_104/a_1020_375# 0.001676f
C8351 output39/a_224_472# net39 0.129913f
C8352 _134_ vdd 0.482157f
C8353 _028_ _155_ 0.049284f
C8354 _079_ _076_ 0.001575f
C8355 _016_ _428_/a_1308_423# 0.00107f
C8356 result[9] net32 0.001371f
C8357 result[6] net61 0.120359f
C8358 output11/a_224_472# _411_/a_36_151# 0.095813f
C8359 ctlp[2] _011_ 0.101324f
C8360 _448_/a_2665_112# trim_val\[4\] 0.004707f
C8361 FILLER_0_4_197/a_1380_472# net76 0.003767f
C8362 output38/a_224_472# _064_ 0.017666f
C8363 _159_ _081_ 0.003646f
C8364 FILLER_0_10_78/a_572_375# cal_count\[3\] 0.002314f
C8365 _339_/a_36_160# FILLER_0_19_171/a_36_472# 0.195478f
C8366 _337_/a_665_69# mask\[1\] 0.002125f
C8367 _086_ FILLER_0_11_135/a_124_375# 0.008238f
C8368 _444_/a_36_151# net49 0.007102f
C8369 _131_ _451_/a_2225_156# 0.008232f
C8370 net59 rstn 0.039664f
C8371 _128_ _426_/a_2665_112# 0.025626f
C8372 _442_/a_36_151# net69 0.048683f
C8373 _119_ _072_ 0.189217f
C8374 FILLER_0_18_209/a_124_375# vss 0.004598f
C8375 FILLER_0_18_209/a_572_375# vdd 0.021356f
C8376 FILLER_0_21_28/a_3260_375# vdd -0.001166f
C8377 _320_/a_1568_472# _043_ 0.00177f
C8378 net52 FILLER_0_2_93/a_124_375# 0.007787f
C8379 output19/a_224_472# _009_ 0.003174f
C8380 _126_ _320_/a_224_472# 0.003754f
C8381 FILLER_0_7_72/a_124_375# FILLER_0_7_59/a_572_375# 0.003228f
C8382 _091_ net80 0.23053f
C8383 net36 FILLER_0_20_87/a_36_472# 0.074773f
C8384 net57 FILLER_0_5_164/a_36_472# 0.032208f
C8385 _162_ FILLER_0_6_177/a_124_375# 0.031168f
C8386 _086_ _068_ 0.080666f
C8387 FILLER_0_2_93/a_572_375# _030_ 0.001718f
C8388 net36 _451_/a_1353_112# 0.01266f
C8389 _074_ cal_itt\[1\] 0.120296f
C8390 net81 net36 0.030215f
C8391 _427_/a_36_151# net23 0.006844f
C8392 FILLER_0_9_223/a_36_472# _090_ 0.001057f
C8393 _447_/a_1308_423# _164_ 0.001422f
C8394 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_36_472# 0.003468f
C8395 FILLER_0_4_107/a_932_472# net47 0.008252f
C8396 _414_/a_796_472# cal_itt\[3\] 0.019699f
C8397 _114_ _055_ 0.071738f
C8398 net81 _429_/a_1204_472# 0.005046f
C8399 net62 output30/a_224_472# 0.074425f
C8400 FILLER_0_4_197/a_932_472# net21 0.00663f
C8401 _186_ cal_count\[2\] 0.001605f
C8402 FILLER_0_20_107/a_124_375# vdd 0.04384f
C8403 _083_ _084_ 0.016693f
C8404 _029_ net47 2.210804f
C8405 FILLER_0_12_20/a_124_375# net17 0.002167f
C8406 _321_/a_170_472# net23 0.025371f
C8407 _449_/a_448_472# cal_count\[3\] 0.007511f
C8408 _028_ _163_ 0.199021f
C8409 result[1] _416_/a_36_151# 0.007739f
C8410 _009_ FILLER_0_23_282/a_124_375# 0.012402f
C8411 FILLER_0_3_172/a_3172_472# net21 0.037958f
C8412 net14 FILLER_0_10_94/a_36_472# 0.003391f
C8413 _091_ mask\[1\] 0.064614f
C8414 net72 cal_count\[1\] 0.13509f
C8415 _066_ net59 0.002935f
C8416 output43/a_224_472# net43 0.11662f
C8417 FILLER_0_18_107/a_124_375# FILLER_0_20_107/a_36_472# 0.00108f
C8418 _115_ _069_ 0.022355f
C8419 net53 _451_/a_36_151# 0.030715f
C8420 FILLER_0_13_142/a_1380_472# net23 0.026285f
C8421 net70 _451_/a_1040_527# 0.002679f
C8422 _120_ _039_ 0.148356f
C8423 _379_/a_36_472# vdd 0.004183f
C8424 FILLER_0_16_107/a_124_375# FILLER_0_16_89/a_1468_375# 0.005439f
C8425 _408_/a_56_524# net47 0.040511f
C8426 _425_/a_1204_472# net37 0.001403f
C8427 net81 FILLER_0_10_247/a_36_472# 0.015109f
C8428 _135_ _134_ 0.038135f
C8429 _077_ _125_ 0.017422f
C8430 _114_ _126_ 3.341247f
C8431 _093_ FILLER_0_16_115/a_36_472# 0.001526f
C8432 _165_ _033_ 0.022734f
C8433 FILLER_0_17_226/a_36_472# _106_ 0.050907f
C8434 FILLER_0_4_123/a_36_472# FILLER_0_2_111/a_1468_375# 0.00189f
C8435 net31 _293_/a_36_472# 0.005692f
C8436 net70 _131_ 0.57653f
C8437 _176_ _055_ 0.001694f
C8438 net20 _288_/a_224_472# 0.003019f
C8439 net48 _123_ 0.153061f
C8440 _119_ _319_/a_234_472# 0.004559f
C8441 net61 _418_/a_36_151# 0.042401f
C8442 net29 vdd 0.611195f
C8443 net81 FILLER_0_15_228/a_36_472# 0.003953f
C8444 _079_ _081_ 1.441057f
C8445 net29 _192_/a_67_603# 0.017997f
C8446 result[7] net61 0.021122f
C8447 net82 FILLER_0_3_221/a_1380_472# 0.008049f
C8448 _426_/a_1308_423# vdd 0.008509f
C8449 _077_ _251_/a_906_472# 0.001076f
C8450 FILLER_0_8_247/a_932_472# calibrate 0.008694f
C8451 _143_ _432_/a_36_151# 0.001486f
C8452 FILLER_0_16_89/a_36_472# vss 0.001289f
C8453 fanout77/a_36_113# net77 0.031558f
C8454 trim_mask\[2\] FILLER_0_3_54/a_36_472# 0.004063f
C8455 net81 en 0.071123f
C8456 _155_ net47 0.009532f
C8457 net71 FILLER_0_19_111/a_484_472# 0.004544f
C8458 _233_/a_36_160# vss 0.01649f
C8459 _175_ FILLER_0_15_72/a_484_472# 0.020589f
C8460 _427_/a_448_472# net74 0.051943f
C8461 FILLER_0_2_93/a_36_472# net14 0.005108f
C8462 net72 FILLER_0_17_38/a_36_472# 0.123542f
C8463 _122_ _066_ 0.001217f
C8464 FILLER_0_13_228/a_124_375# net79 0.008554f
C8465 FILLER_0_17_64/a_36_472# vss 0.006428f
C8466 FILLER_0_18_107/a_2364_375# _022_ 0.001902f
C8467 net20 FILLER_0_15_235/a_124_375# 0.001278f
C8468 FILLER_0_18_177/a_1380_472# _139_ 0.00195f
C8469 net23 _146_ 0.034955f
C8470 FILLER_0_17_142/a_36_472# vss 0.008239f
C8471 FILLER_0_17_142/a_484_472# vdd 0.004902f
C8472 mask\[4\] FILLER_0_19_195/a_124_375# 0.006236f
C8473 _431_/a_796_472# _136_ 0.009889f
C8474 net17 output40/a_224_472# 0.00187f
C8475 _335_/a_49_472# _137_ 0.03139f
C8476 _151_ _365_/a_36_68# 0.001944f
C8477 FILLER_0_6_47/a_1020_375# vdd 0.016637f
C8478 net57 _121_ 0.004182f
C8479 FILLER_0_14_107/a_124_375# _451_/a_36_151# 0.059049f
C8480 net31 net19 0.023019f
C8481 _072_ FILLER_0_10_214/a_36_472# 0.015199f
C8482 FILLER_0_18_107/a_3172_472# FILLER_0_17_133/a_124_375# 0.001543f
C8483 _427_/a_2665_112# _095_ 0.039612f
C8484 _126_ _176_ 0.057877f
C8485 net27 _426_/a_2560_156# 0.004199f
C8486 net20 _411_/a_36_151# 0.011179f
C8487 _053_ FILLER_0_6_47/a_3172_472# 0.001777f
C8488 mask\[9\] FILLER_0_19_111/a_572_375# 0.027695f
C8489 trim_mask\[2\] net14 0.060278f
C8490 FILLER_0_15_142/a_484_472# vdd 0.001097f
C8491 FILLER_0_5_117/a_36_472# _154_ 0.005034f
C8492 _186_ _043_ 0.045082f
C8493 _033_ net40 0.298492f
C8494 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1468_375# 0.086635f
C8495 _066_ _169_ 0.222791f
C8496 FILLER_0_3_142/a_36_472# _443_/a_36_151# 0.001723f
C8497 _122_ net23 0.276617f
C8498 vdd FILLER_0_12_196/a_124_375# 0.015159f
C8499 _274_/a_36_68# FILLER_0_12_236/a_484_472# 0.001237f
C8500 FILLER_0_10_78/a_124_375# FILLER_0_9_72/a_932_472# 0.001543f
C8501 _428_/a_2248_156# net53 0.001188f
C8502 _339_/a_36_160# vss 0.027338f
C8503 trim_mask\[2\] _164_ 1.859062f
C8504 _161_ _061_ 0.026347f
C8505 _144_ _145_ 0.671767f
C8506 _050_ _436_/a_1308_423# 0.022688f
C8507 _081_ cal_itt\[1\] 0.009747f
C8508 _444_/a_1000_472# net47 0.036015f
C8509 _161_ _311_/a_66_473# 0.021817f
C8510 _016_ FILLER_0_12_136/a_36_472# 0.016227f
C8511 FILLER_0_7_72/a_2812_375# net14 0.025092f
C8512 _227_/a_36_160# net23 0.055152f
C8513 vdd FILLER_0_6_231/a_124_375# 0.024542f
C8514 net52 vss 1.608047f
C8515 net74 _318_/a_224_472# 0.001513f
C8516 _000_ _411_/a_796_472# 0.044697f
C8517 net51 net6 0.142515f
C8518 _068_ _313_/a_67_603# 0.012208f
C8519 _415_/a_2665_112# vss 0.015461f
C8520 net63 _435_/a_1000_472# 0.002536f
C8521 net57 _443_/a_36_151# 0.003322f
C8522 FILLER_0_8_24/a_484_472# net47 0.042018f
C8523 net67 _450_/a_36_151# 0.067819f
C8524 FILLER_0_18_107/a_2276_472# vdd 0.004405f
C8525 net23 _169_ 0.00151f
C8526 _325_/a_224_472# _120_ 0.00233f
C8527 FILLER_0_4_197/a_1468_375# net22 0.009108f
C8528 _126_ _124_ 0.012466f
C8529 _434_/a_2560_156# mask\[6\] 0.010913f
C8530 trim_mask\[4\] _163_ 0.003686f
C8531 net35 _434_/a_2665_112# 0.024254f
C8532 FILLER_0_15_150/a_36_472# vdd 0.088307f
C8533 result[2] net19 0.065763f
C8534 _128_ _223_/a_36_160# 0.012824f
C8535 _102_ vss 0.068703f
C8536 _394_/a_1336_472# _175_ 0.002792f
C8537 _424_/a_1000_472# vdd 0.002952f
C8538 _413_/a_36_151# FILLER_0_3_172/a_2364_375# 0.059049f
C8539 _024_ net33 0.001047f
C8540 net49 vss 0.689397f
C8541 net47 _163_ 0.64626f
C8542 output29/a_224_472# _416_/a_2665_112# 0.011048f
C8543 net65 cal_itt\[1\] 0.049124f
C8544 mask\[4\] FILLER_0_18_177/a_1828_472# 0.014226f
C8545 _027_ FILLER_0_18_76/a_572_375# 0.08501f
C8546 _150_ FILLER_0_18_76/a_484_472# 0.003548f
C8547 _122_ FILLER_0_5_172/a_36_472# 0.003007f
C8548 net20 FILLER_0_6_239/a_36_472# 0.005138f
C8549 net50 _441_/a_1000_472# 0.02354f
C8550 net52 _441_/a_2248_156# 0.023959f
C8551 FILLER_0_4_107/a_36_472# _153_ 0.042459f
C8552 FILLER_0_4_107/a_932_472# _154_ 0.017867f
C8553 mask\[3\] FILLER_0_18_177/a_932_472# 0.005654f
C8554 _447_/a_2665_112# trim_val\[3\] 0.002721f
C8555 FILLER_0_23_290/a_124_375# FILLER_0_23_282/a_572_375# 0.012001f
C8556 FILLER_0_12_124/a_124_375# vdd -0.00168f
C8557 net54 FILLER_0_19_111/a_36_472# 0.003467f
C8558 net60 vdd 0.575502f
C8559 fanout73/a_36_113# _427_/a_36_151# 0.032681f
C8560 net18 _417_/a_1204_472# 0.01349f
C8561 FILLER_0_16_57/a_572_375# net15 0.013085f
C8562 _091_ mask\[0\] 0.04171f
C8563 _029_ _154_ 0.116532f
C8564 _417_/a_2248_156# net30 0.048831f
C8565 FILLER_0_18_2/a_2276_472# net47 0.001369f
C8566 _072_ _161_ 0.048567f
C8567 _441_/a_2248_156# net49 0.048164f
C8568 _415_/a_1204_472# net27 0.006198f
C8569 FILLER_0_5_117/a_124_375# _160_ 0.008534f
C8570 FILLER_0_21_206/a_124_375# _204_/a_67_603# 0.003591f
C8571 FILLER_0_21_125/a_124_375# mask\[7\] 0.00145f
C8572 FILLER_0_5_172/a_124_375# _163_ 0.006403f
C8573 FILLER_0_8_239/a_124_375# vss 0.017196f
C8574 FILLER_0_8_239/a_36_472# vdd 0.079402f
C8575 _074_ FILLER_0_6_177/a_124_375# 0.003608f
C8576 FILLER_0_5_72/a_124_375# vdd -0.005497f
C8577 _053_ _219_/a_36_160# 0.005244f
C8578 net15 _183_ 0.007353f
C8579 _031_ FILLER_0_2_111/a_572_375# 0.023633f
C8580 net69 FILLER_0_2_111/a_1468_375# 0.021524f
C8581 net14 FILLER_0_4_91/a_124_375# 0.009573f
C8582 _272_/a_36_472# _087_ 0.048282f
C8583 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_572_375# 0.086635f
C8584 net72 _038_ 0.013821f
C8585 net81 output27/a_224_472# 0.011872f
C8586 _050_ _208_/a_36_160# 0.001038f
C8587 _245_/a_234_472# _067_ 0.005071f
C8588 trim_val\[0\] trim_mask\[1\] 0.003033f
C8589 _174_ _067_ 0.002678f
C8590 ctlp[4] vss 0.102044f
C8591 FILLER_0_12_136/a_1380_472# FILLER_0_13_142/a_572_375# 0.001684f
C8592 net41 _452_/a_36_151# 0.036301f
C8593 _367_/a_36_68# _157_ 0.013352f
C8594 FILLER_0_9_223/a_124_375# _070_ 0.002989f
C8595 output25/a_224_472# _214_/a_36_160# 0.027335f
C8596 output46/a_224_472# FILLER_0_20_15/a_572_375# 0.00135f
C8597 _446_/a_36_151# net40 0.015376f
C8598 _028_ FILLER_0_7_104/a_1020_375# 0.004954f
C8599 _012_ FILLER_0_23_44/a_484_472# 0.001572f
C8600 _274_/a_244_497# net64 0.004085f
C8601 net16 _402_/a_728_93# 0.040925f
C8602 _114_ state\[1\] 0.087216f
C8603 _081_ FILLER_0_5_148/a_124_375# 0.021583f
C8604 _105_ net33 0.202272f
C8605 _421_/a_36_151# net19 0.016842f
C8606 _011_ mask\[7\] 0.043474f
C8607 _187_ _174_ 0.001321f
C8608 fanout63/a_36_160# _098_ 0.003627f
C8609 net15 FILLER_0_15_59/a_572_375# 0.033245f
C8610 net36 FILLER_0_15_180/a_572_375# 0.002531f
C8611 net74 _163_ 0.042013f
C8612 _116_ FILLER_0_13_206/a_124_375# 0.003926f
C8613 output32/a_224_472# net19 0.08441f
C8614 trim[4] FILLER_0_8_2/a_124_375# 0.028454f
C8615 _267_/a_36_472# _055_ 0.035376f
C8616 FILLER_0_14_91/a_484_472# _176_ 0.003624f
C8617 FILLER_0_19_155/a_36_472# _145_ 0.005521f
C8618 net51 _450_/a_2225_156# 0.009822f
C8619 _091_ FILLER_0_15_212/a_124_375# 0.025529f
C8620 _441_/a_36_151# _160_ 0.030777f
C8621 _086_ _113_ 0.072034f
C8622 net57 FILLER_0_13_142/a_1380_472# 0.011768f
C8623 _155_ _154_ 0.18488f
C8624 FILLER_0_21_125/a_36_472# vss 0.00143f
C8625 net34 FILLER_0_22_128/a_1380_472# 0.001011f
C8626 output21/a_224_472# _009_ 0.004164f
C8627 FILLER_0_21_125/a_484_472# vdd 0.002728f
C8628 mask\[4\] FILLER_0_22_128/a_3172_472# 0.001484f
C8629 FILLER_0_15_72/a_572_375# vss 0.007579f
C8630 FILLER_0_15_72/a_36_472# vdd 0.108844f
C8631 _004_ FILLER_0_10_256/a_124_375# 0.006989f
C8632 FILLER_0_17_200/a_36_472# vss 0.001182f
C8633 net73 net71 0.033964f
C8634 FILLER_0_10_78/a_932_472# _115_ 0.013773f
C8635 _053_ FILLER_0_6_177/a_484_472# 0.015994f
C8636 FILLER_0_4_197/a_1468_375# vdd 0.019672f
C8637 FILLER_0_20_193/a_572_375# net35 0.002196f
C8638 output24/a_224_472# _050_ 0.061723f
C8639 _419_/a_36_151# net77 0.163616f
C8640 ctlp[4] _107_ 0.080312f
C8641 _427_/a_2248_156# state\[1\] 0.001849f
C8642 mask\[5\] _048_ 0.062788f
C8643 net52 FILLER_0_2_165/a_36_472# 0.002601f
C8644 net64 FILLER_0_12_220/a_1380_472# 0.011079f
C8645 net47 FILLER_0_4_91/a_36_472# 0.005186f
C8646 net46 FILLER_0_21_28/a_36_472# 0.051176f
C8647 FILLER_0_3_2/a_124_375# vdd 0.021963f
C8648 _176_ state\[1\] 0.001641f
C8649 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1380_472# 0.003468f
C8650 _093_ FILLER_0_19_155/a_124_375# 0.001864f
C8651 _269_/a_36_472# _080_ 0.003981f
C8652 _083_ _260_/a_36_68# 0.047191f
C8653 net81 _425_/a_2560_156# 0.022037f
C8654 net55 FILLER_0_18_37/a_1380_472# 0.007432f
C8655 output9/a_224_472# net5 0.005189f
C8656 _136_ _137_ 0.417639f
C8657 _035_ _446_/a_448_472# 0.018273f
C8658 FILLER_0_2_111/a_1380_472# FILLER_0_2_127/a_36_472# 0.013276f
C8659 _322_/a_1084_68# _128_ 0.002629f
C8660 net55 FILLER_0_17_56/a_124_375# 0.014472f
C8661 net72 FILLER_0_17_56/a_484_472# 0.003359f
C8662 _413_/a_36_151# net76 0.084453f
C8663 _070_ FILLER_0_10_107/a_36_472# 0.013252f
C8664 net78 _421_/a_1204_472# 0.006482f
C8665 result[5] net18 0.173673f
C8666 _396_/a_224_472# _176_ 0.008359f
C8667 output19/a_224_472# net33 0.126671f
C8668 _441_/a_2560_156# _164_ 0.049213f
C8669 _056_ _061_ 0.445098f
C8670 FILLER_0_18_171/a_36_472# _141_ 0.002037f
C8671 _414_/a_2248_156# cal_itt\[3\] 0.032294f
C8672 FILLER_0_7_72/a_2724_472# _219_/a_36_160# 0.001448f
C8673 _077_ net68 0.003823f
C8674 _056_ _311_/a_66_473# 0.026074f
C8675 _428_/a_796_472# vdd 0.003502f
C8676 _098_ _433_/a_796_472# 0.002825f
C8677 output36/a_224_472# net62 0.317201f
C8678 FILLER_0_16_255/a_124_375# net19 0.008033f
C8679 net4 _083_ 0.135165f
C8680 net20 net76 0.021613f
C8681 _437_/a_448_472# net14 0.090442f
C8682 _127_ FILLER_0_11_135/a_36_472# 0.044488f
C8683 _088_ net59 0.270902f
C8684 _076_ FILLER_0_9_142/a_124_375# 0.001774f
C8685 net1 _265_/a_244_68# 0.023821f
C8686 _070_ _248_/a_36_68# 0.007095f
C8687 _086_ _321_/a_2590_472# 0.001522f
C8688 _065_ output16/a_224_472# 0.049052f
C8689 _163_ _154_ 0.190662f
C8690 net27 net18 0.092379f
C8691 _444_/a_2665_112# trim_val\[0\] 0.007249f
C8692 FILLER_0_11_142/a_572_375# net23 0.010863f
C8693 _081_ FILLER_0_6_177/a_124_375# 0.005524f
C8694 _422_/a_1308_423# _009_ 0.008875f
C8695 net6 clkc 0.036083f
C8696 output14/a_224_472# _442_/a_2248_156# 0.001723f
C8697 net80 _434_/a_1000_472# 0.01421f
C8698 FILLER_0_16_57/a_1380_472# vss 0.011192f
C8699 FILLER_0_4_197/a_484_472# net21 0.046864f
C8700 net57 _122_ 0.034045f
C8701 _132_ FILLER_0_14_107/a_36_472# 0.002187f
C8702 cal_count\[3\] FILLER_0_11_124/a_36_472# 0.00702f
C8703 _131_ _331_/a_448_472# 0.007271f
C8704 net15 _449_/a_1204_472# 0.01349f
C8705 _091_ FILLER_0_12_220/a_1020_375# 0.001598f
C8706 FILLER_0_20_177/a_572_375# _098_ 0.015373f
C8707 _061_ _068_ 1.857322f
C8708 FILLER_0_15_212/a_932_472# mask\[1\] 0.014799f
C8709 net7 vdd 0.321735f
C8710 FILLER_0_7_72/a_572_375# net50 0.012932f
C8711 net55 _452_/a_448_472# 0.05323f
C8712 trim_mask\[2\] _153_ 0.007934f
C8713 _123_ net37 0.002942f
C8714 _068_ _311_/a_66_473# 0.071325f
C8715 _072_ _056_ 0.061377f
C8716 net20 _419_/a_1308_423# 0.022245f
C8717 _425_/a_36_151# _316_/a_848_380# 0.035903f
C8718 net25 FILLER_0_23_88/a_124_375# 0.010782f
C8719 net76 FILLER_0_1_192/a_124_375# 0.00275f
C8720 _425_/a_2665_112# net18 0.003301f
C8721 _053_ net4 0.013559f
C8722 _073_ net37 0.013152f
C8723 _065_ _447_/a_2665_112# 0.034757f
C8724 net57 _169_ 0.033365f
C8725 trim_mask\[1\] FILLER_0_6_47/a_484_472# 0.022211f
C8726 _073_ FILLER_0_3_221/a_1468_375# 0.006377f
C8727 _274_/a_36_68# net81 0.014689f
C8728 _434_/a_2665_112# vdd 0.030225f
C8729 FILLER_0_18_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001684f
C8730 _171_ net14 0.020479f
C8731 _043_ _225_/a_36_160# 0.007958f
C8732 _148_ mask\[7\] 0.010238f
C8733 net35 _024_ 0.001335f
C8734 _412_/a_2665_112# fanout59/a_36_160# 0.016426f
C8735 _028_ FILLER_0_7_72/a_1916_375# 0.003862f
C8736 _431_/a_448_472# net73 0.050964f
C8737 net20 _043_ 0.094689f
C8738 _077_ net67 0.073924f
C8739 net81 FILLER_0_14_235/a_484_472# 0.015266f
C8740 ctln[4] FILLER_0_1_204/a_124_375# 0.008283f
C8741 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_36_472# 0.002296f
C8742 _322_/a_124_24# vdd 0.01572f
C8743 result[7] FILLER_0_23_274/a_36_472# 0.014434f
C8744 _421_/a_36_151# _419_/a_448_472# 0.002098f
C8745 _043_ FILLER_0_12_196/a_36_472# 0.001526f
C8746 _290_/a_224_472# _094_ 0.003006f
C8747 _411_/a_1204_472# vss 0.001746f
C8748 _446_/a_2665_112# _034_ 0.002484f
C8749 _187_ _450_/a_3129_107# 0.00126f
C8750 FILLER_0_15_290/a_36_472# vss 0.010015f
C8751 FILLER_0_2_101/a_124_375# vdd 0.044073f
C8752 vss FILLER_0_8_156/a_36_472# 0.00168f
C8753 vdd FILLER_0_8_156/a_484_472# 0.007249f
C8754 output8/a_224_472# FILLER_0_3_221/a_1380_472# 0.001699f
C8755 _188_ FILLER_0_12_50/a_124_375# 0.00157f
C8756 net35 FILLER_0_22_128/a_2812_375# 0.010399f
C8757 net53 _137_ 0.008376f
C8758 net17 _452_/a_448_472# 0.043154f
C8759 _077_ FILLER_0_11_64/a_36_472# 0.076102f
C8760 output32/a_224_472# _419_/a_448_472# 0.010723f
C8761 _072_ _068_ 0.185471f
C8762 net33 mask\[6\] 0.881813f
C8763 _415_/a_448_472# FILLER_0_9_270/a_36_472# 0.012285f
C8764 FILLER_0_13_100/a_36_472# net14 0.046864f
C8765 net68 FILLER_0_6_47/a_1468_375# 0.022624f
C8766 _064_ _445_/a_2560_156# 0.005361f
C8767 FILLER_0_10_78/a_484_472# vss 0.005854f
C8768 fanout81/a_36_160# net76 0.001905f
C8769 net15 _439_/a_796_472# 0.001822f
C8770 _185_ _405_/a_255_603# 0.002565f
C8771 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_572_375# 0.001597f
C8772 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_36_472# 0.026657f
C8773 FILLER_0_18_100/a_124_375# _438_/a_2248_156# 0.001068f
C8774 _052_ vss 0.077815f
C8775 vss _202_/a_36_160# 0.010418f
C8776 net60 _419_/a_796_472# 0.003097f
C8777 net61 _419_/a_1204_472# 0.012025f
C8778 mask\[5\] FILLER_0_18_177/a_484_472# 0.001063f
C8779 fanout66/a_36_113# net69 0.001345f
C8780 net47 net6 0.23883f
C8781 FILLER_0_17_104/a_1468_375# vss 0.001786f
C8782 FILLER_0_17_104/a_36_472# vdd 0.095484f
C8783 _444_/a_36_151# net40 0.032012f
C8784 mask\[2\] net23 0.431197f
C8785 net62 FILLER_0_14_263/a_36_472# 0.019591f
C8786 _025_ vss 0.016676f
C8787 cal_count\[3\] cal_count\[0\] 0.098735f
C8788 ctlp[1] FILLER_0_21_286/a_484_472# 0.045536f
C8789 _322_/a_848_380# _125_ 0.013667f
C8790 net28 net29 0.178557f
C8791 _004_ mask\[1\] 0.052788f
C8792 _440_/a_1000_472# _029_ 0.004334f
C8793 _269_/a_36_472# vss 0.014227f
C8794 FILLER_0_18_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001597f
C8795 _140_ _149_ 0.0088f
C8796 _132_ vss 0.492496f
C8797 net55 FILLER_0_18_53/a_124_375# 0.011674f
C8798 net72 FILLER_0_18_53/a_484_472# 0.001067f
C8799 net52 _036_ 0.013473f
C8800 net50 net68 0.224698f
C8801 FILLER_0_10_78/a_572_375# net52 0.003311f
C8802 FILLER_0_8_138/a_124_375# vdd 0.024547f
C8803 net16 FILLER_0_8_37/a_36_472# 0.012905f
C8804 _267_/a_36_472# state\[1\] 0.001647f
C8805 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_36_472# 0.007947f
C8806 FILLER_0_23_290/a_124_375# vdd 0.030435f
C8807 net39 _445_/a_2665_112# 0.002831f
C8808 FILLER_0_15_116/a_36_472# net36 0.013546f
C8809 FILLER_0_5_72/a_1380_472# trim_mask\[1\] 0.01221f
C8810 mask\[2\] FILLER_0_15_212/a_484_472# 0.001641f
C8811 _139_ _337_/a_49_472# 0.024331f
C8812 trimb[0] net43 0.109028f
C8813 _428_/a_36_151# FILLER_0_13_100/a_36_472# 0.004032f
C8814 _036_ net49 0.005235f
C8815 _093_ FILLER_0_21_60/a_484_472# 0.001396f
C8816 _404_/a_36_472# _179_ 0.00141f
C8817 _431_/a_2248_156# FILLER_0_17_142/a_572_375# 0.006739f
C8818 net34 _146_ 0.004718f
C8819 _063_ net67 0.039144f
C8820 FILLER_0_4_99/a_36_472# net14 0.022408f
C8821 net50 _156_ 0.020099f
C8822 _050_ FILLER_0_22_107/a_124_375# 0.002634f
C8823 FILLER_0_20_193/a_572_375# vdd 0.029393f
C8824 FILLER_0_17_72/a_932_472# _131_ 0.002672f
C8825 FILLER_0_9_28/a_2276_472# vss -0.001894f
C8826 trim_val\[4\] _066_ 0.015621f
C8827 _088_ FILLER_0_5_206/a_124_375# 0.001374f
C8828 _079_ FILLER_0_5_206/a_36_472# 0.008243f
C8829 net16 _160_ 0.354736f
C8830 _420_/a_448_472# _009_ 0.061681f
C8831 FILLER_0_19_111/a_124_375# net14 0.001837f
C8832 _136_ _040_ 0.788826f
C8833 FILLER_0_12_136/a_484_472# vdd 0.005304f
C8834 FILLER_0_12_136/a_36_472# vss 0.003185f
C8835 mask\[7\] _436_/a_2665_112# 0.004274f
C8836 FILLER_0_15_116/a_484_472# net70 0.049569f
C8837 FILLER_0_15_116/a_124_375# net53 0.009286f
C8838 cal_itt\[3\] net76 0.017174f
C8839 _438_/a_36_151# net71 0.053065f
C8840 fanout61/a_36_113# vss 0.05514f
C8841 _421_/a_2248_156# _109_ 0.001349f
C8842 _132_ FILLER_0_19_125/a_36_472# 0.008568f
C8843 _412_/a_36_151# vdd 0.080326f
C8844 _002_ vss 0.08396f
C8845 result[7] FILLER_0_24_274/a_1468_375# 0.006125f
C8846 FILLER_0_5_212/a_36_472# net37 0.007858f
C8847 FILLER_0_7_195/a_36_472# vss 0.002568f
C8848 _032_ net23 0.019676f
C8849 net52 _449_/a_448_472# 0.001042f
C8850 _286_/a_224_472# _094_ 0.008468f
C8851 _008_ output31/a_224_472# 0.051074f
C8852 FILLER_0_5_54/a_36_472# vdd 0.006056f
C8853 FILLER_0_5_54/a_1468_375# vss 0.053407f
C8854 _412_/a_2665_112# net5 0.042084f
C8855 FILLER_0_17_72/a_2364_375# net36 0.005483f
C8856 FILLER_0_16_241/a_36_472# FILLER_0_15_235/a_572_375# 0.001543f
C8857 net75 net58 0.061787f
C8858 FILLER_0_7_104/a_124_375# _153_ 0.001205f
C8859 FILLER_0_7_104/a_1020_375# _154_ 0.005051f
C8860 FILLER_0_18_177/a_1020_375# FILLER_0_20_177/a_932_472# 0.0027f
C8861 _442_/a_2248_156# vdd 0.038702f
C8862 trim_val\[4\] net23 0.014503f
C8863 _213_/a_67_603# _098_ 0.018092f
C8864 FILLER_0_10_37/a_124_375# _042_ 0.002437f
C8865 net74 _172_ 0.006643f
C8866 _165_ _054_ 0.001337f
C8867 net38 _445_/a_2248_156# 0.029721f
C8868 net50 net67 0.518421f
C8869 FILLER_0_4_185/a_124_375# _087_ 0.120668f
C8870 FILLER_0_18_177/a_1468_375# vdd 0.024167f
C8871 FILLER_0_16_241/a_36_472# vdd 0.012388f
C8872 FILLER_0_16_241/a_124_375# vss 0.04897f
C8873 FILLER_0_4_177/a_484_472# vss 0.002399f
C8874 net47 _450_/a_2225_156# 0.057106f
C8875 _449_/a_1000_472# _067_ 0.021759f
C8876 _307_/a_672_472# _114_ 0.0018f
C8877 _128_ _121_ 0.051501f
C8878 FILLER_0_12_20/a_484_472# vdd 0.003108f
C8879 _112_ vdd 0.086153f
C8880 cal_itt\[3\] FILLER_0_5_198/a_124_375# 0.01268f
C8881 _450_/a_448_472# _039_ 0.047559f
C8882 _413_/a_2248_156# vdd -0.006767f
C8883 net75 _425_/a_448_472# 0.038993f
C8884 cal_count\[3\] _070_ 0.059233f
C8885 net16 FILLER_0_18_37/a_124_375# 0.017482f
C8886 _053_ _058_ 0.075418f
C8887 _095_ FILLER_0_15_72/a_572_375# 0.00352f
C8888 net23 FILLER_0_16_154/a_484_472# 0.001369f
C8889 _105_ net22 0.01308f
C8890 output12/a_224_472# net76 0.00803f
C8891 net69 _031_ 0.450281f
C8892 _431_/a_2665_112# net73 0.001495f
C8893 _070_ _059_ 0.041498f
C8894 state\[0\] vss 0.126943f
C8895 _239_/a_36_160# net16 0.003137f
C8896 _370_/a_848_380# vdd -0.001256f
C8897 _370_/a_124_24# vss 0.005764f
C8898 result[6] net62 0.005382f
C8899 mask\[7\] FILLER_0_22_128/a_1468_375# 0.0178f
C8900 net17 FILLER_0_20_15/a_572_375# 0.018398f
C8901 net73 FILLER_0_18_107/a_3260_375# 0.001629f
C8902 _163_ FILLER_0_5_148/a_124_375# 0.001706f
C8903 _165_ vss 0.048027f
C8904 FILLER_0_7_146/a_36_472# _059_ 0.073041f
C8905 net75 _082_ 0.417366f
C8906 net75 net82 0.214597f
C8907 fanout53/a_36_160# _427_/a_2665_112# 0.00285f
C8908 _002_ FILLER_0_3_172/a_3260_375# 0.001683f
C8909 _255_/a_224_552# vdd 0.082462f
C8910 output21/a_224_472# net33 0.001166f
C8911 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1380_472# 0.026657f
C8912 net31 net20 0.238809f
C8913 _428_/a_1000_472# _043_ 0.020031f
C8914 FILLER_0_14_50/a_124_375# cal_count\[3\] 0.002524f
C8915 FILLER_0_21_28/a_2724_472# _424_/a_36_151# 0.001723f
C8916 cal_itt\[2\] FILLER_0_3_221/a_124_375# 0.006217f
C8917 net15 FILLER_0_21_60/a_484_472# 0.001552f
C8918 _077_ FILLER_0_6_231/a_36_472# 0.075292f
C8919 _054_ net40 0.072879f
C8920 _247_/a_36_160# vss 0.009308f
C8921 _412_/a_36_151# net9 0.005212f
C8922 _246_/a_36_68# _055_ 0.028938f
C8923 _356_/a_36_472# net36 0.004539f
C8924 FILLER_0_16_57/a_572_375# FILLER_0_15_59/a_484_472# 0.001543f
C8925 fanout69/a_36_113# trim_mask\[4\] 0.027938f
C8926 _024_ vdd 0.091532f
C8927 _176_ _394_/a_718_524# 0.00141f
C8928 FILLER_0_4_152/a_36_472# trim_mask\[4\] 0.011746f
C8929 ctln[7] FILLER_0_0_96/a_124_375# 0.025944f
C8930 net55 cal_count\[3\] 0.005157f
C8931 net57 _097_ 0.100409f
C8932 cal_count\[1\] vdd 0.516859f
C8933 _428_/a_1308_423# _095_ 0.001504f
C8934 _443_/a_1204_472# _170_ 0.002808f
C8935 net15 _440_/a_1308_423# 0.015192f
C8936 net2 net37 0.05083f
C8937 _061_ _113_ 0.012561f
C8938 state\[2\] FILLER_0_13_142/a_1468_375# 0.018691f
C8939 net53 FILLER_0_13_142/a_484_472# 0.059444f
C8940 FILLER_0_4_152/a_36_472# net47 0.007541f
C8941 net63 _434_/a_2665_112# 0.120476f
C8942 _091_ FILLER_0_13_212/a_572_375# 0.022882f
C8943 _043_ _039_ 0.001161f
C8944 net53 _040_ 0.035628f
C8945 FILLER_0_24_274/a_484_472# vdd 0.004641f
C8946 FILLER_0_24_274/a_36_472# vss 0.001013f
C8947 _367_/a_692_472# net14 0.00423f
C8948 _448_/a_2248_156# _037_ 0.027079f
C8949 _091_ FILLER_0_10_214/a_124_375# 0.006331f
C8950 FILLER_0_12_28/a_36_472# vss 0.003004f
C8951 _141_ _146_ 0.020044f
C8952 _162_ _062_ 0.033583f
C8953 _449_/a_2665_112# _172_ 0.003296f
C8954 vss net40 0.898805f
C8955 FILLER_0_2_93/a_484_472# FILLER_0_0_96/a_124_375# 0.001338f
C8956 FILLER_0_12_124/a_36_472# _126_ 0.056268f
C8957 _178_ net40 0.029542f
C8958 _348_/a_49_472# _146_ 0.001552f
C8959 FILLER_0_22_128/a_2812_375# vdd 0.003766f
C8960 FILLER_0_22_128/a_2364_375# vss 0.017496f
C8961 fanout56/a_36_113# _136_ 0.002316f
C8962 net71 FILLER_0_22_107/a_36_472# 0.034505f
C8963 net35 mask\[6\] 0.041818f
C8964 FILLER_0_9_28/a_1828_472# vdd 0.006263f
C8965 mask\[8\] net35 2.631701f
C8966 _292_/a_36_160# output18/a_224_472# 0.009736f
C8967 net41 net16 2.918931f
C8968 _086_ FILLER_0_11_142/a_484_472# 0.008338f
C8969 FILLER_0_4_177/a_572_375# FILLER_0_5_181/a_124_375# 0.05841f
C8970 _028_ _439_/a_796_472# 0.013039f
C8971 FILLER_0_20_15/a_932_472# net40 0.002705f
C8972 FILLER_0_18_171/a_124_375# vss 0.048769f
C8973 FILLER_0_6_79/a_124_375# vss 0.007008f
C8974 FILLER_0_6_79/a_36_472# vdd 0.087807f
C8975 _131_ _062_ 0.120189f
C8976 cal net59 0.297816f
C8977 _087_ FILLER_0_3_172/a_1828_472# 0.027954f
C8978 _086_ FILLER_0_7_104/a_1468_375# 0.065371f
C8979 net60 net77 0.046792f
C8980 _021_ _137_ 0.002807f
C8981 _232_/a_67_603# trim_mask\[1\] 0.022808f
C8982 cal_count\[3\] net17 0.068527f
C8983 net57 mask\[2\] 0.022012f
C8984 net82 FILLER_0_3_172/a_1020_375# 0.010679f
C8985 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_36_472# 0.002765f
C8986 _095_ _281_/a_672_472# 0.00134f
C8987 net16 FILLER_0_19_47/a_36_472# 0.009509f
C8988 _104_ _198_/a_67_603# 0.007168f
C8989 FILLER_0_15_282/a_36_472# vss 0.004616f
C8990 _120_ FILLER_0_9_72/a_1380_472# 0.001723f
C8991 FILLER_0_17_38/a_572_375# vss 0.007503f
C8992 FILLER_0_17_38/a_36_472# vdd 0.01637f
C8993 trim_mask\[4\] _371_/a_36_113# 0.007529f
C8994 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_484_472# 0.013276f
C8995 _143_ net80 0.023487f
C8996 _178_ FILLER_0_17_38/a_572_375# 0.031538f
C8997 net79 _018_ 0.069992f
C8998 _065_ net66 0.003956f
C8999 FILLER_0_3_172/a_124_375# net65 0.021073f
C9000 net65 _425_/a_2665_112# 0.00628f
C9001 mask\[5\] _145_ 0.012075f
C9002 FILLER_0_3_204/a_124_375# net59 0.007104f
C9003 _105_ vdd 0.565719f
C9004 result[9] _094_ 0.03984f
C9005 _392_/a_36_68# vdd 0.036386f
C9006 net72 cal_count\[2\] 0.073818f
C9007 vdd FILLER_0_3_212/a_124_375# 0.025095f
C9008 FILLER_0_6_177/a_124_375# _163_ 0.025831f
C9009 net62 _418_/a_36_151# 0.029844f
C9010 _198_/a_67_603# vss 0.003647f
C9011 _081_ _261_/a_36_160# 0.049069f
C9012 _144_ _434_/a_36_151# 0.004055f
C9013 _316_/a_124_24# calibrate 0.016936f
C9014 net64 net36 0.037523f
C9015 fanout69/a_36_113# net74 0.034782f
C9016 valid sample 0.103192f
C9017 en net59 0.490893f
C9018 FILLER_0_14_107/a_124_375# _040_ 0.001861f
C9019 _236_/a_36_160# _064_ 0.039922f
C9020 valid net37 0.051518f
C9021 _073_ net8 0.206839f
C9022 FILLER_0_9_28/a_2724_472# trim_val\[0\] 0.001183f
C9023 _256_/a_716_497# _128_ 0.001035f
C9024 FILLER_0_21_142/a_484_472# net54 0.038728f
C9025 _413_/a_36_151# FILLER_0_1_192/a_36_472# 0.046516f
C9026 net52 FILLER_0_6_47/a_2812_375# 0.018463f
C9027 net72 FILLER_0_19_28/a_484_472# 0.004312f
C9028 net55 FILLER_0_19_28/a_124_375# 0.002644f
C9029 FILLER_0_7_104/a_932_472# _151_ 0.002092f
C9030 net20 FILLER_0_6_231/a_36_472# 0.045553f
C9031 _136_ _334_/a_36_160# 0.005574f
C9032 _402_/a_1948_68# _179_ 0.005403f
C9033 net48 _079_ 0.012855f
C9034 FILLER_0_12_2/a_484_472# net6 0.005586f
C9035 trimb[2] net17 0.007637f
C9036 _127_ _118_ 0.141388f
C9037 FILLER_0_4_144/a_36_472# vdd 0.004289f
C9038 FILLER_0_4_144/a_572_375# vss 0.072463f
C9039 _443_/a_1000_472# net69 0.008276f
C9040 FILLER_0_10_256/a_36_472# FILLER_0_10_247/a_36_472# 0.001963f
C9041 FILLER_0_16_73/a_36_472# net15 0.005297f
C9042 FILLER_0_24_96/a_36_472# net35 0.002526f
C9043 FILLER_0_24_63/a_124_375# ctlp[8] 0.005758f
C9044 net54 FILLER_0_22_107/a_572_375# 0.002239f
C9045 net20 output32/a_224_472# 0.050019f
C9046 _426_/a_2248_156# FILLER_0_8_239/a_124_375# 0.001068f
C9047 net63 FILLER_0_20_193/a_572_375# 0.015818f
C9048 _433_/a_448_472# _145_ 0.045046f
C9049 FILLER_0_10_247/a_36_472# net64 0.059367f
C9050 net34 _422_/a_2665_112# 0.006103f
C9051 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_124_375# 0.004426f
C9052 FILLER_0_16_73/a_572_375# _131_ 0.011479f
C9053 net67 _039_ 0.302826f
C9054 FILLER_0_4_99/a_36_472# _153_ 0.066147f
C9055 FILLER_0_16_107/a_124_375# _136_ 0.00661f
C9056 _412_/a_2248_156# fanout59/a_36_160# 0.007753f
C9057 _093_ _397_/a_36_472# 0.001509f
C9058 net22 mask\[6\] 0.612004f
C9059 net71 _433_/a_36_151# 0.014126f
C9060 FILLER_0_17_72/a_124_375# vdd 0.0132f
C9061 _430_/a_36_151# FILLER_0_17_200/a_124_375# 0.059049f
C9062 FILLER_0_11_135/a_36_472# _118_ 0.002496f
C9063 FILLER_0_18_2/a_484_472# vdd 0.003495f
C9064 output19/a_224_472# vdd 0.063651f
C9065 net20 _277_/a_36_160# 0.015569f
C9066 net81 _426_/a_36_151# 0.060652f
C9067 FILLER_0_2_101/a_36_472# _156_ 0.001487f
C9068 net57 trim_val\[4\] 0.295336f
C9069 net55 FILLER_0_17_72/a_1828_472# 0.001217f
C9070 net29 FILLER_0_16_255/a_36_472# 0.086886f
C9071 FILLER_0_24_130/a_124_375# output23/a_224_472# 0.006051f
C9072 net36 _006_ 0.001331f
C9073 _132_ _095_ 0.042874f
C9074 FILLER_0_4_107/a_124_375# vdd 0.036972f
C9075 FILLER_0_16_89/a_36_472# _451_/a_448_472# 0.011974f
C9076 ctln[6] _442_/a_448_472# 0.003039f
C9077 FILLER_0_2_111/a_572_375# _158_ 0.031641f
C9078 fanout69/a_36_113# _159_ 0.005623f
C9079 net74 _371_/a_36_113# 0.027966f
C9080 _415_/a_2248_156# net58 0.001869f
C9081 _077_ FILLER_0_12_50/a_124_375# 0.008485f
C9082 result[9] net78 0.015761f
C9083 net16 FILLER_0_14_50/a_36_472# 0.001377f
C9084 FILLER_0_19_28/a_124_375# net17 0.007234f
C9085 _413_/a_448_472# net76 0.029504f
C9086 net47 net37 0.057409f
C9087 _445_/a_2665_112# net47 0.041188f
C9088 _440_/a_2560_156# vss 0.002793f
C9089 _091_ _429_/a_36_151# 0.006557f
C9090 en net64 0.01789f
C9091 _029_ _365_/a_36_68# 0.013994f
C9092 net54 FILLER_0_20_98/a_124_375# 0.001639f
C9093 net63 FILLER_0_18_177/a_1468_375# 0.020059f
C9094 _257_/a_36_472# _053_ 0.00507f
C9095 net57 FILLER_0_16_154/a_484_472# 0.001532f
C9096 _120_ vdd 0.750809f
C9097 _038_ vdd 0.043998f
C9098 net60 _421_/a_448_472# 0.052759f
C9099 net72 _043_ 0.05655f
C9100 FILLER_0_21_28/a_3172_472# _012_ 0.018785f
C9101 _128_ _122_ 0.019207f
C9102 _017_ FILLER_0_14_107/a_932_472# 0.001941f
C9103 FILLER_0_16_89/a_1020_375# _131_ 0.015706f
C9104 net38 _034_ 0.025823f
C9105 FILLER_0_16_73/a_124_375# vss 0.026383f
C9106 net79 vss 0.770834f
C9107 _119_ net23 0.0245f
C9108 FILLER_0_12_136/a_1468_375# _126_ 0.012732f
C9109 _414_/a_796_472# vdd 0.001497f
C9110 FILLER_0_23_282/a_124_375# vdd -0.003896f
C9111 _303_/a_36_472# vss 0.011549f
C9112 _431_/a_36_151# _093_ 0.004862f
C9113 FILLER_0_1_266/a_484_472# net8 0.016327f
C9114 _438_/a_2248_156# vdd 0.024595f
C9115 FILLER_0_13_142/a_1020_375# vdd 0.018221f
C9116 ctlp[1] _419_/a_2560_156# 0.002551f
C9117 _431_/a_796_472# _020_ 0.012284f
C9118 FILLER_0_13_142/a_572_375# vss 0.04084f
C9119 net66 _440_/a_448_472# 0.023934f
C9120 FILLER_0_5_172/a_124_375# net37 0.014083f
C9121 net73 FILLER_0_19_111/a_484_472# 0.007404f
C9122 net52 FILLER_0_5_72/a_36_472# 0.014911f
C9123 _184_ net40 0.122833f
C9124 _128_ net64 0.291788f
C9125 net41 _041_ 0.076779f
C9126 output25/a_224_472# net25 0.179738f
C9127 _211_/a_36_160# _050_ 0.010927f
C9128 _010_ _108_ 0.002048f
C9129 _151_ net14 0.009212f
C9130 FILLER_0_18_107/a_124_375# _438_/a_2665_112# 0.029834f
C9131 _010_ net19 0.408364f
C9132 net19 FILLER_0_14_263/a_124_375# 0.032085f
C9133 net44 FILLER_0_15_2/a_36_472# 0.007808f
C9134 output29/a_224_472# net30 0.044542f
C9135 FILLER_0_15_2/a_484_472# vss 0.003267f
C9136 _371_/a_36_113# _159_ 0.021612f
C9137 _081_ FILLER_0_5_136/a_124_375# 0.025819f
C9138 net23 _208_/a_36_160# 0.112626f
C9139 net69 _157_ 0.112249f
C9140 _164_ FILLER_0_6_47/a_36_472# 0.047981f
C9141 _074_ _062_ 0.005012f
C9142 net68 FILLER_0_5_54/a_484_472# 0.047601f
C9143 FILLER_0_21_133/a_124_375# net54 0.013027f
C9144 FILLER_0_11_282/a_124_375# vdd 0.026044f
C9145 net15 _453_/a_448_472# 0.040851f
C9146 net63 _024_ 0.001348f
C9147 _030_ _160_ 0.063581f
C9148 net66 _034_ 0.139638f
C9149 net49 _166_ 0.007445f
C9150 _155_ _365_/a_36_68# 0.053708f
C9151 FILLER_0_21_125/a_484_472# _140_ 0.013936f
C9152 FILLER_0_15_142/a_572_375# vdd -0.013698f
C9153 _447_/a_2665_112# net69 0.002067f
C9154 _430_/a_1000_472# net21 0.053061f
C9155 output9/a_224_472# ctln[2] 0.080206f
C9156 _076_ _062_ 0.978627f
C9157 mask\[6\] vdd 0.573103f
C9158 _417_/a_2248_156# _006_ 0.039121f
C9159 FILLER_0_7_104/a_932_472# _131_ 0.011713f
C9160 mask\[8\] vdd 0.423606f
C9161 output35/a_224_472# FILLER_0_21_206/a_36_472# 0.0323f
C9162 _114_ _121_ 0.002513f
C9163 _320_/a_36_472# _090_ 0.001941f
C9164 net56 FILLER_0_17_142/a_124_375# 0.004803f
C9165 _253_/a_36_68# FILLER_0_3_221/a_1468_375# 0.014131f
C9166 net75 calibrate 0.101912f
C9167 _429_/a_2560_156# vss 0.005255f
C9168 FILLER_0_17_56/a_36_472# vss 0.00167f
C9169 FILLER_0_17_56/a_484_472# vdd 0.002789f
C9170 _412_/a_2560_156# net18 0.015371f
C9171 FILLER_0_13_212/a_1380_472# mask\[0\] 0.002361f
C9172 fanout52/a_36_160# vdd 0.026513f
C9173 _412_/a_2248_156# net5 0.048919f
C9174 _258_/a_36_160# _081_ 0.00776f
C9175 _135_ _120_ 0.017522f
C9176 net75 FILLER_0_10_256/a_124_375# 0.027258f
C9177 fanout80/a_36_113# _019_ 0.003644f
C9178 net79 _416_/a_2248_156# 0.026136f
C9179 _093_ FILLER_0_17_218/a_124_375# 0.003338f
C9180 FILLER_0_5_128/a_124_375# _163_ 0.009765f
C9181 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_572_375# 0.086635f
C9182 net55 FILLER_0_18_76/a_572_375# 0.002278f
C9183 output27/a_224_472# net64 0.04953f
C9184 net62 _416_/a_2665_112# 0.037195f
C9185 vdd FILLER_0_13_290/a_36_472# 0.027484f
C9186 vss FILLER_0_13_290/a_124_375# 0.031844f
C9187 cal_count\[3\] _408_/a_1336_472# 0.010351f
C9188 mask\[4\] net23 0.111873f
C9189 state\[2\] vdd 0.392508f
C9190 _077_ _078_ 0.069858f
C9191 net26 _424_/a_1204_472# 0.00194f
C9192 _186_ _180_ 0.003034f
C9193 _453_/a_1308_423# _042_ 0.001778f
C9194 _453_/a_448_472# net51 0.006397f
C9195 output8/a_224_472# net75 0.044765f
C9196 output21/a_224_472# net22 0.022576f
C9197 FILLER_0_20_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001543f
C9198 net4 net5 0.104296f
C9199 _440_/a_36_151# _164_ 0.003699f
C9200 output44/a_224_472# FILLER_0_20_15/a_36_472# 0.0323f
C9201 _386_/a_848_380# vss 0.012638f
C9202 FILLER_0_10_78/a_1468_375# _389_/a_36_148# 0.001699f
C9203 _008_ _093_ 0.252609f
C9204 _175_ vdd 0.147794f
C9205 _010_ _420_/a_36_151# 0.001838f
C9206 _421_/a_36_151# _009_ 0.00246f
C9207 _163_ _365_/a_36_68# 0.004035f
C9208 FILLER_0_19_171/a_1020_375# vdd 0.025918f
C9209 _132_ _332_/a_36_472# 0.055537f
C9210 _176_ _121_ 0.035608f
C9211 FILLER_0_22_86/a_484_472# net71 0.00583f
C9212 net15 FILLER_0_13_72/a_36_472# 0.006713f
C9213 result[6] fanout77/a_36_113# 0.001469f
C9214 _095_ net40 0.674445f
C9215 net36 _097_ 0.022089f
C9216 _451_/a_1040_527# net14 0.029964f
C9217 FILLER_0_5_72/a_932_472# _164_ 0.011079f
C9218 _088_ FILLER_0_4_213/a_572_375# 0.022684f
C9219 fanout60/a_36_160# result[3] 0.00188f
C9220 _452_/a_836_156# vdd 0.002533f
C9221 net55 FILLER_0_21_28/a_2812_375# 0.004005f
C9222 _091_ FILLER_0_15_180/a_36_472# 0.00375f
C9223 FILLER_0_23_290/a_124_375# net77 0.001783f
C9224 FILLER_0_7_162/a_36_472# calibrate 0.014431f
C9225 _024_ FILLER_0_22_177/a_124_375# 0.005166f
C9226 _144_ _354_/a_665_69# 0.001518f
C9227 _036_ net40 0.599505f
C9228 FILLER_0_24_96/a_36_472# vdd 0.094828f
C9229 trim_mask\[4\] FILLER_0_2_111/a_1020_375# 0.02806f
C9230 trim[4] net44 0.188184f
C9231 _050_ net71 0.033192f
C9232 FILLER_0_18_177/a_3172_472# net21 0.010321f
C9233 fanout63/a_36_160# mask\[1\] 0.009907f
C9234 net20 FILLER_0_13_228/a_124_375# 0.047331f
C9235 _256_/a_2960_68# _056_ 0.001168f
C9236 _131_ net14 0.037705f
C9237 _377_/a_36_472# trim_mask\[1\] 0.001763f
C9238 _003_ _079_ 0.035497f
C9239 net34 _419_/a_2665_112# 0.001468f
C9240 _012_ FILLER_0_21_60/a_484_472# 0.01517f
C9241 _440_/a_1308_423# net47 0.009738f
C9242 _141_ mask\[2\] 0.084094f
C9243 _306_/a_36_68# _043_ 0.001086f
C9244 output22/a_224_472# _435_/a_36_151# 0.12978f
C9245 result[5] _418_/a_796_472# 0.001983f
C9246 FILLER_0_14_107/a_1020_375# vdd 0.008956f
C9247 FILLER_0_9_72/a_932_472# vdd 0.00604f
C9248 FILLER_0_9_72/a_484_472# vss 0.008087f
C9249 _430_/a_36_151# mask\[3\] 0.005848f
C9250 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_124_375# 0.012222f
C9251 _420_/a_36_151# FILLER_0_23_282/a_36_472# 0.001723f
C9252 _414_/a_2248_156# net22 0.062122f
C9253 _013_ mask\[9\] 0.011224f
C9254 FILLER_0_8_107/a_36_472# vdd 0.117254f
C9255 result[4] fanout60/a_36_160# 0.027276f
C9256 net36 mask\[2\] 0.871463f
C9257 net15 FILLER_0_9_60/a_124_375# 0.003602f
C9258 net1 vdd 0.63891f
C9259 _085_ _090_ 0.001012f
C9260 _116_ _060_ 0.020653f
C9261 _010_ _419_/a_448_472# 0.003295f
C9262 _020_ _137_ 0.228674f
C9263 FILLER_0_10_78/a_1468_375# _115_ 0.032403f
C9264 _453_/a_2665_112# vss 0.037567f
C9265 _311_/a_2180_473# vdd 0.001974f
C9266 calibrate _059_ 0.506928f
C9267 _430_/a_2248_156# vss 0.030251f
C9268 _015_ _426_/a_2665_112# 0.018623f
C9269 FILLER_0_18_2/a_3172_472# _452_/a_36_151# 0.059367f
C9270 net64 _416_/a_36_151# 0.013586f
C9271 _232_/a_67_603# net66 0.001758f
C9272 FILLER_0_19_55/a_36_472# net55 0.062683f
C9273 FILLER_0_19_47/a_36_472# _424_/a_1308_423# 0.010224f
C9274 output9/a_224_472# net81 0.02825f
C9275 output44/a_224_472# FILLER_0_18_2/a_1468_375# 0.032639f
C9276 _131_ _404_/a_36_472# 0.031567f
C9277 _079_ net37 0.408392f
C9278 FILLER_0_18_2/a_1828_472# net38 0.006713f
C9279 _411_/a_448_472# net75 0.072712f
C9280 _000_ FILLER_0_3_221/a_1380_472# 0.025567f
C9281 _119_ net57 0.30462f
C9282 _426_/a_36_151# _317_/a_36_113# 0.001082f
C9283 _136_ FILLER_0_16_154/a_1468_375# 0.0028f
C9284 _428_/a_36_151# _131_ 0.00821f
C9285 net3 FILLER_0_15_2/a_572_375# 0.004377f
C9286 _443_/a_2248_156# net59 0.002471f
C9287 net52 _387_/a_36_113# 0.02405f
C9288 net20 _078_ 0.105266f
C9289 fanout49/a_36_160# net49 0.032999f
C9290 trimb[1] FILLER_0_20_2/a_36_472# 0.003628f
C9291 net40 output41/a_224_472# 0.081551f
C9292 _091_ FILLER_0_18_177/a_484_472# 0.004272f
C9293 _261_/a_36_160# _163_ 0.002002f
C9294 output21/a_224_472# vdd 0.028725f
C9295 net32 _421_/a_2665_112# 0.019532f
C9296 net81 FILLER_0_15_212/a_1380_472# 0.003953f
C9297 _118_ _060_ 0.002868f
C9298 vdd _433_/a_2248_156# 0.008127f
C9299 mask\[0\] _429_/a_2248_156# 0.016246f
C9300 _089_ net21 0.006605f
C9301 _077_ _057_ 0.584179f
C9302 FILLER_0_13_65/a_124_375# fanout72/a_36_113# 0.005467f
C9303 fanout77/a_36_113# _418_/a_36_151# 0.001082f
C9304 _005_ mask\[1\] 0.246517f
C9305 FILLER_0_3_172/a_2364_375# net22 0.013028f
C9306 _288_/a_224_472# vdd 0.002071f
C9307 FILLER_0_18_53/a_484_472# vdd 0.002358f
C9308 FILLER_0_18_53/a_36_472# vss 0.001471f
C9309 _094_ _418_/a_1000_472# 0.053462f
C9310 _143_ FILLER_0_18_139/a_1380_472# 0.002226f
C9311 FILLER_0_17_133/a_124_375# vss 0.015434f
C9312 FILLER_0_17_133/a_36_472# vdd 0.097394f
C9313 _057_ _267_/a_1120_472# 0.001833f
C9314 input5/a_36_113# vss 0.005833f
C9315 _052_ _424_/a_2560_156# 0.003401f
C9316 FILLER_0_16_57/a_484_472# _131_ 0.008223f
C9317 _414_/a_36_151# _089_ 0.039611f
C9318 net34 FILLER_0_22_177/a_36_472# 0.003953f
C9319 _221_/a_36_160# vdd 0.073414f
C9320 FILLER_0_9_60/a_124_375# net51 0.002346f
C9321 _343_/a_49_472# _093_ 0.001926f
C9322 _187_ _453_/a_36_151# 0.001829f
C9323 fanout55/a_36_160# FILLER_0_13_80/a_36_472# 0.003699f
C9324 output33/a_224_472# net32 0.018183f
C9325 net55 FILLER_0_17_64/a_36_472# 0.034504f
C9326 _410_/a_36_68# cal_count\[3\] 0.001096f
C9327 _151_ _153_ 0.027868f
C9328 _115_ FILLER_0_10_94/a_572_375# 0.00887f
C9329 net74 _390_/a_36_68# 0.008011f
C9330 net36 FILLER_0_16_115/a_124_375# 0.001706f
C9331 _321_/a_170_472# _176_ 0.059301f
C9332 _415_/a_1204_472# _004_ 0.002391f
C9333 _053_ FILLER_0_6_47/a_1020_375# 0.015621f
C9334 FILLER_0_7_104/a_1380_472# _133_ 0.004838f
C9335 _274_/a_36_68# net64 0.036017f
C9336 _292_/a_36_160# _048_ 0.008475f
C9337 _093_ FILLER_0_17_72/a_36_472# 0.001971f
C9338 FILLER_0_10_28/a_124_375# vss 0.013087f
C9339 FILLER_0_10_28/a_36_472# vdd 0.092132f
C9340 _069_ _120_ 0.030804f
C9341 net16 _408_/a_728_93# 0.107634f
C9342 _008_ _418_/a_1204_472# 0.002933f
C9343 _126_ _136_ 0.086459f
C9344 FILLER_0_15_235/a_124_375# vdd -0.006807f
C9345 result[0] vdd 0.193436f
C9346 FILLER_0_9_105/a_572_375# vdd 0.074717f
C9347 net54 _210_/a_67_603# 0.001108f
C9348 FILLER_0_13_142/a_1468_375# _043_ 0.009636f
C9349 FILLER_0_20_177/a_1468_375# vss 0.053913f
C9350 FILLER_0_20_177/a_36_472# vdd 0.114932f
C9351 _114_ FILLER_0_10_94/a_484_472# 0.011954f
C9352 FILLER_0_21_142/a_572_375# FILLER_0_22_128/a_2276_472# 0.001543f
C9353 FILLER_0_17_200/a_124_375# mask\[3\] 0.01841f
C9354 net64 FILLER_0_14_235/a_484_472# 0.012355f
C9355 net35 _423_/a_2665_112# 0.019085f
C9356 _086_ _087_ 0.015938f
C9357 FILLER_0_21_125/a_36_472# _098_ 0.002923f
C9358 result[9] _418_/a_2248_156# 0.043716f
C9359 _411_/a_36_151# vdd 0.077963f
C9360 cal_itt\[1\] FILLER_0_3_221/a_1468_375# 0.020427f
C9361 _398_/a_36_113# net44 0.011803f
C9362 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1468_375# 0.086742f
C9363 ctln[9] _447_/a_448_472# 0.003564f
C9364 net16 _447_/a_796_472# 0.003278f
C9365 FILLER_0_7_162/a_124_375# calibrate 0.014255f
C9366 net36 FILLER_0_15_212/a_572_375# 0.004606f
C9367 _414_/a_2248_156# vdd 0.00901f
C9368 _104_ _422_/a_448_472# 0.001955f
C9369 net70 FILLER_0_16_115/a_36_472# 0.003407f
C9370 _414_/a_448_472# _089_ 0.003905f
C9371 net63 mask\[6\] 0.146994f
C9372 _276_/a_36_160# FILLER_0_18_209/a_572_375# 0.004736f
C9373 _429_/a_36_151# FILLER_0_15_212/a_932_472# 0.001723f
C9374 state\[0\] _426_/a_2248_156# 0.001198f
C9375 _426_/a_36_151# _425_/a_1308_423# 0.001518f
C9376 _116_ _118_ 0.054068f
C9377 FILLER_0_20_15/a_1468_375# vss 0.055156f
C9378 FILLER_0_20_15/a_36_472# vdd 0.086947f
C9379 _233_/a_36_160# net17 0.003831f
C9380 output25/a_224_472# ctlp[8] 0.018544f
C9381 FILLER_0_18_107/a_124_375# vdd 0.030961f
C9382 _321_/a_3126_472# _118_ 0.002754f
C9383 net52 net55 0.016401f
C9384 _267_/a_36_472# _121_ 0.041237f
C9385 _422_/a_1308_423# vdd 0.004083f
C9386 _168_ vss 0.171346f
C9387 _062_ _090_ 0.010805f
C9388 _412_/a_1308_423# net65 0.024499f
C9389 net79 FILLER_0_12_220/a_124_375# 0.010895f
C9390 _441_/a_796_472# vss 0.001231f
C9391 net31 net33 0.002465f
C9392 result[6] _419_/a_36_151# 0.001968f
C9393 _063_ _033_ 0.250192f
C9394 _031_ _369_/a_36_68# 0.050502f
C9395 net69 _158_ 0.033459f
C9396 _067_ FILLER_0_13_72/a_572_375# 0.001874f
C9397 mask\[9\] net71 0.344312f
C9398 _064_ _446_/a_2665_112# 0.039211f
C9399 _415_/a_448_472# result[1] 0.005209f
C9400 FILLER_0_16_241/a_36_472# _282_/a_36_160# 0.006647f
C9401 _293_/a_36_472# vss 0.014842f
C9402 output36/a_224_472# net29 0.077505f
C9403 FILLER_0_14_81/a_36_472# cal_count\[1\] 0.034486f
C9404 mask\[4\] FILLER_0_19_155/a_484_472# 0.024522f
C9405 _132_ _451_/a_448_472# 0.001197f
C9406 _005_ _416_/a_2560_156# 0.004273f
C9407 FILLER_0_19_55/a_36_472# _216_/a_67_603# 0.00254f
C9408 _176_ FILLER_0_10_94/a_484_472# 0.009483f
C9409 FILLER_0_9_28/a_36_472# net51 0.002082f
C9410 _125_ vdd 0.218505f
C9411 _131_ FILLER_0_17_104/a_572_375# 0.003214f
C9412 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_36_472# 0.003468f
C9413 _057_ _225_/a_36_160# 0.026341f
C9414 FILLER_0_21_142/a_36_472# net23 0.001629f
C9415 FILLER_0_6_239/a_36_472# vdd 0.092399f
C9416 FILLER_0_6_239/a_124_375# vss 0.017355f
C9417 net81 _015_ 0.002818f
C9418 _415_/a_2665_112# net58 0.005219f
C9419 ctlp[1] _421_/a_2248_156# 0.012937f
C9420 _139_ _019_ 0.094494f
C9421 net69 net66 0.09789f
C9422 net15 _423_/a_36_151# 0.003422f
C9423 FILLER_0_17_142/a_484_472# _137_ 0.003953f
C9424 _104_ _108_ 0.02837f
C9425 FILLER_0_20_31/a_36_472# vss 0.004923f
C9426 _444_/a_2665_112# FILLER_0_6_37/a_124_375# 0.005477f
C9427 _449_/a_36_151# _038_ 0.019666f
C9428 FILLER_0_3_172/a_2364_375# vdd -0.010717f
C9429 _359_/a_36_488# _133_ 0.04287f
C9430 FILLER_0_5_54/a_572_375# _440_/a_36_151# 0.026916f
C9431 net63 FILLER_0_19_171/a_1020_375# 0.004794f
C9432 FILLER_0_11_101/a_124_375# net14 0.011983f
C9433 _104_ net19 0.159483f
C9434 _108_ vss 0.160825f
C9435 ctlp[3] _296_/a_224_472# 0.005335f
C9436 _431_/a_2248_156# _136_ 0.030673f
C9437 net16 FILLER_0_16_37/a_36_472# 0.015199f
C9438 FILLER_0_9_28/a_2724_472# _453_/a_36_151# 0.013806f
C9439 _163_ FILLER_0_5_136/a_124_375# 0.009765f
C9440 _251_/a_468_472# vss 0.001679f
C9441 _413_/a_448_472# FILLER_0_1_192/a_36_472# 0.001462f
C9442 net19 vss 1.140787f
C9443 net50 _033_ 0.003088f
C9444 net36 FILLER_0_15_205/a_124_375# 0.004337f
C9445 _232_/a_255_603# net47 0.001241f
C9446 _423_/a_36_151# FILLER_0_23_44/a_1380_472# 0.001723f
C9447 net76 net22 0.118787f
C9448 net49 net17 0.029142f
C9449 FILLER_0_9_28/a_2364_375# _077_ 0.00397f
C9450 net62 result[1] 0.061866f
C9451 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1468_375# 0.016748f
C9452 net15 FILLER_0_17_72/a_36_472# 0.006905f
C9453 _077_ FILLER_0_7_72/a_484_472# 0.001332f
C9454 vss _416_/a_796_472# 0.001468f
C9455 _422_/a_1000_472# _108_ 0.027806f
C9456 _188_ vss 0.032923f
C9457 _069_ state\[2\] 0.023375f
C9458 _281_/a_672_472# _098_ 0.002084f
C9459 net65 FILLER_0_2_171/a_36_472# 0.023858f
C9460 FILLER_0_21_206/a_36_472# net21 0.132984f
C9461 net52 net82 0.108202f
C9462 FILLER_0_10_78/a_36_472# cal_count\[3\] 0.266339f
C9463 _140_ _024_ 0.00287f
C9464 _091_ _090_ 0.117348f
C9465 _189_/a_67_603# _100_ 0.002818f
C9466 net4 _055_ 0.216844f
C9467 FILLER_0_11_142/a_124_375# cal_count\[3\] 0.010782f
C9468 FILLER_0_22_177/a_124_375# mask\[6\] 0.002672f
C9469 _098_ _434_/a_2248_156# 0.016991f
C9470 output44/a_224_472# net46 0.003211f
C9471 FILLER_0_18_107/a_2276_472# _137_ 0.001752f
C9472 net75 output48/a_224_472# 0.070114f
C9473 cal_itt\[3\] _078_ 0.024443f
C9474 FILLER_0_14_91/a_484_472# _136_ 0.038919f
C9475 _053_ _359_/a_1492_488# 0.001437f
C9476 _093_ net54 0.003211f
C9477 net79 FILLER_0_12_236/a_36_472# 0.009225f
C9478 _238_/a_67_603# net52 0.006325f
C9479 net69 FILLER_0_3_54/a_124_375# 0.004245f
C9480 net34 _208_/a_36_160# 0.002666f
C9481 net16 trim_val\[2\] 0.124462f
C9482 FILLER_0_4_49/a_36_472# net66 0.012791f
C9483 net75 FILLER_0_8_247/a_124_375# 0.002085f
C9484 _140_ FILLER_0_22_128/a_2812_375# 0.003154f
C9485 net52 FILLER_0_3_78/a_484_472# 0.003143f
C9486 _108_ _107_ 0.018045f
C9487 en_co_clk fanout55/a_36_160# 0.041263f
C9488 mask\[5\] _434_/a_36_151# 0.00104f
C9489 net35 _435_/a_2248_156# 0.001854f
C9490 result[7] _419_/a_36_151# 0.001036f
C9491 _068_ net23 0.432092f
C9492 net68 _167_ 0.001302f
C9493 FILLER_0_2_177/a_124_375# net22 0.001318f
C9494 net49 FILLER_0_3_78/a_484_472# 0.048729f
C9495 FILLER_0_17_161/a_124_375# vss 0.00824f
C9496 FILLER_0_17_161/a_36_472# vdd 0.006972f
C9497 _125_ _135_ 0.001926f
C9498 _043_ net22 0.041447f
C9499 _320_/a_1792_472# vdd 0.001113f
C9500 net15 _447_/a_2248_156# 0.01843f
C9501 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_124_375# 0.012001f
C9502 net26 net72 0.868238f
C9503 _093_ net15 0.145303f
C9504 _098_ _202_/a_36_160# 0.006831f
C9505 cal_count\[2\] vdd 0.932907f
C9506 _235_/a_67_603# net68 0.027525f
C9507 FILLER_0_3_172/a_3172_472# net65 0.001777f
C9508 _005_ _099_ 0.001603f
C9509 _127_ net74 0.0588f
C9510 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_124_375# 0.012001f
C9511 _013_ _424_/a_36_151# 0.012928f
C9512 _095_ FILLER_0_14_107/a_572_375# 0.01418f
C9513 net72 FILLER_0_12_50/a_124_375# 0.011077f
C9514 net19 _416_/a_2248_156# 0.024466f
C9515 _420_/a_448_472# vdd 0.010071f
C9516 _420_/a_36_151# vss 0.043027f
C9517 net4 FILLER_0_12_220/a_572_375# 0.019052f
C9518 input3/a_36_113# vdd 0.117445f
C9519 FILLER_0_5_109/a_572_375# FILLER_0_5_117/a_36_472# 0.086635f
C9520 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_484_472# 0.001723f
C9521 FILLER_0_19_47/a_572_375# _052_ 0.020156f
C9522 _132_ _098_ 0.038463f
C9523 _228_/a_36_68# _060_ 0.016962f
C9524 FILLER_0_16_89/a_1020_375# FILLER_0_17_72/a_2812_375# 0.026339f
C9525 FILLER_0_16_89/a_36_472# FILLER_0_17_72/a_1916_375# 0.001723f
C9526 FILLER_0_4_49/a_572_375# FILLER_0_3_54/a_36_472# 0.001597f
C9527 _431_/a_2248_156# net53 0.003335f
C9528 net61 fanout78/a_36_113# 0.056484f
C9529 net34 mask\[4\] 0.001774f
C9530 FILLER_0_19_28/a_484_472# vdd 0.010504f
C9531 net47 _365_/a_244_472# 0.001431f
C9532 output46/a_224_472# net40 0.002542f
C9533 _446_/a_1204_472# net66 0.001885f
C9534 net76 vdd 1.272072f
C9535 vss _450_/a_36_151# 0.02803f
C9536 vdd _450_/a_448_472# 0.011591f
C9537 FILLER_0_4_197/a_1380_472# vss 0.007979f
C9538 cal_count\[3\] _373_/a_1060_68# 0.00165f
C9539 FILLER_0_10_78/a_932_472# _120_ 0.003672f
C9540 FILLER_0_7_72/a_572_375# vdd 0.004039f
C9541 net20 _010_ 0.016197f
C9542 trimb[0] net44 0.00246f
C9543 trim_mask\[1\] FILLER_0_4_91/a_484_472# 0.002806f
C9544 _423_/a_2248_156# vss 0.010039f
C9545 _423_/a_2665_112# vdd 0.022696f
C9546 FILLER_0_16_57/a_1380_472# net55 0.002219f
C9547 _431_/a_1308_423# _427_/a_36_151# 0.001256f
C9548 _155_ FILLER_0_6_90/a_484_472# 0.005297f
C9549 FILLER_0_8_127/a_36_472# _133_ 0.004423f
C9550 net69 net23 0.064573f
C9551 cal_count\[3\] _171_ 0.00961f
C9552 _076_ FILLER_0_8_156/a_124_375# 0.0062f
C9553 _070_ FILLER_0_8_156/a_36_472# 0.001338f
C9554 FILLER_0_20_193/a_124_375# _098_ 0.009717f
C9555 _062_ _163_ 0.001206f
C9556 _343_/a_257_69# _093_ 0.001043f
C9557 FILLER_0_16_154/a_124_375# vdd 0.00439f
C9558 _253_/a_672_68# _074_ 0.001857f
C9559 _096_ net57 0.05086f
C9560 FILLER_0_14_91/a_484_472# net53 0.00544f
C9561 _150_ vdd 0.05295f
C9562 FILLER_0_4_49/a_572_375# _164_ 0.005532f
C9563 _440_/a_36_151# FILLER_0_6_47/a_2724_472# 0.001653f
C9564 FILLER_0_7_72/a_484_472# net50 0.059395f
C9565 _142_ net56 0.028797f
C9566 FILLER_0_17_72/a_3172_472# vdd 0.002712f
C9567 net22 _435_/a_2248_156# 0.003453f
C9568 _079_ net8 0.001928f
C9569 FILLER_0_5_198/a_124_375# vdd 0.010749f
C9570 _057_ cal_itt\[3\] 0.014849f
C9571 FILLER_0_22_86/a_1020_375# net14 0.047331f
C9572 FILLER_0_5_109/a_572_375# FILLER_0_4_107/a_932_472# 0.001684f
C9573 _419_/a_1308_423# vdd 0.007543f
C9574 FILLER_0_21_133/a_124_375# _144_ 0.001885f
C9575 _185_ net40 0.048742f
C9576 FILLER_0_16_89/a_484_472# _040_ 0.009871f
C9577 mask\[0\] cal_count\[3\] 0.002612f
C9578 _116_ _228_/a_36_68# 0.013091f
C9579 _152_ net23 0.001895f
C9580 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3172_472# 0.026657f
C9581 _414_/a_2665_112# net59 0.010265f
C9582 FILLER_0_2_177/a_124_375# vdd 0.019296f
C9583 FILLER_0_12_136/a_124_375# _127_ 0.004013f
C9584 FILLER_0_16_89/a_124_375# _093_ 0.004086f
C9585 _372_/a_358_69# _070_ 0.001293f
C9586 net74 FILLER_0_13_72/a_36_472# 0.007448f
C9587 net44 _190_/a_36_160# 0.015628f
C9588 _043_ vdd 0.827689f
C9589 output33/a_224_472# _421_/a_2665_112# 0.010726f
C9590 net53 state\[1\] 0.00554f
C9591 trim_val\[4\] FILLER_0_3_172/a_572_375# 0.001076f
C9592 output15/a_224_472# ctln[8] 0.079231f
C9593 _114_ _097_ 0.004412f
C9594 _072_ FILLER_0_12_220/a_484_472# 0.028355f
C9595 net4 FILLER_0_12_236/a_484_472# 0.014212f
C9596 net70 FILLER_0_14_99/a_124_375# 0.002922f
C9597 net62 FILLER_0_13_212/a_124_375# 0.001597f
C9598 _291_/a_36_160# output18/a_224_472# 0.001175f
C9599 FILLER_0_6_90/a_484_472# _163_ 0.011711f
C9600 _058_ _055_ 0.070216f
C9601 _186_ vss 0.0718f
C9602 output22/a_224_472# net23 0.008048f
C9603 _035_ _160_ 0.120469f
C9604 _178_ _186_ 0.020123f
C9605 _369_/a_36_68# _157_ 0.068266f
C9606 net46 vdd 0.255965f
C9607 net4 FILLER_0_3_221/a_124_375# 0.015788f
C9608 FILLER_0_4_49/a_484_472# net47 0.002964f
C9609 mask\[7\] _435_/a_796_472# 0.009587f
C9610 _394_/a_56_524# cal_count\[1\] 0.022487f
C9611 _345_/a_36_160# _144_ 0.00465f
C9612 net55 _052_ 0.095046f
C9613 _131_ FILLER_0_14_123/a_124_375# 0.016964f
C9614 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1468_375# 0.086635f
C9615 _059_ _242_/a_36_160# 0.001942f
C9616 _062_ _117_ 0.042699f
C9617 net16 _174_ 0.022224f
C9618 net68 vdd 1.026897f
C9619 net22 FILLER_0_18_209/a_484_472# 0.005297f
C9620 _415_/a_36_151# _426_/a_36_151# 0.002121f
C9621 cal_itt\[1\] net8 0.040042f
C9622 _176_ _174_ 0.00677f
C9623 _026_ vdd 0.15542f
C9624 _414_/a_2665_112# _122_ 0.007441f
C9625 _020_ _334_/a_36_160# 0.028435f
C9626 net4 state\[1\] 0.010195f
C9627 net23 FILLER_0_22_128/a_2276_472# 0.011079f
C9628 FILLER_0_3_2/a_36_472# _446_/a_36_151# 0.004032f
C9629 FILLER_0_18_139/a_1020_375# vss 0.032606f
C9630 FILLER_0_17_200/a_572_375# FILLER_0_18_177/a_3172_472# 0.001597f
C9631 FILLER_0_18_139/a_1468_375# vdd 0.015542f
C9632 _426_/a_448_472# calibrate 0.002745f
C9633 _432_/a_2665_112# _430_/a_36_151# 0.030053f
C9634 _415_/a_448_472# net81 0.004045f
C9635 FILLER_0_9_72/a_36_472# _439_/a_36_151# 0.001723f
C9636 FILLER_0_15_282/a_124_375# net18 0.048284f
C9637 _093_ FILLER_0_18_107/a_36_472# 0.008683f
C9638 _036_ _168_ 0.01699f
C9639 FILLER_0_15_282/a_484_472# output30/a_224_472# 0.001711f
C9640 FILLER_0_7_72/a_1468_375# FILLER_0_5_72/a_1380_472# 0.00108f
C9641 net19 _419_/a_1000_472# 0.012949f
C9642 FILLER_0_9_28/a_36_472# net47 0.006712f
C9643 FILLER_0_10_256/a_36_472# _426_/a_36_151# 0.059238f
C9644 FILLER_0_12_28/a_36_472# cal_count\[0\] 0.001662f
C9645 _093_ _302_/a_224_472# 0.011376f
C9646 net15 net51 0.191328f
C9647 FILLER_0_18_177/a_3260_375# _202_/a_36_160# 0.001948f
C9648 mask\[4\] _141_ 0.948091f
C9649 vdd _156_ 0.178622f
C9650 _426_/a_36_151# net64 0.022056f
C9651 _063_ _444_/a_36_151# 0.030369f
C9652 cal_itt\[2\] net59 0.014956f
C9653 FILLER_0_14_81/a_36_472# _175_ 0.076977f
C9654 mask\[4\] _348_/a_49_472# 0.001241f
C9655 _392_/a_36_68# FILLER_0_12_50/a_36_472# 0.002811f
C9656 net31 net22 0.002533f
C9657 _439_/a_36_151# _453_/a_2248_156# 0.001082f
C9658 _140_ mask\[6\] 0.605898f
C9659 FILLER_0_1_204/a_36_472# net11 0.014707f
C9660 mask\[8\] _140_ 0.003375f
C9661 FILLER_0_7_72/a_1020_375# vss 0.004851f
C9662 net41 FILLER_0_12_28/a_124_375# 0.003909f
C9663 net71 _437_/a_2248_156# 0.025557f
C9664 _440_/a_2665_112# _160_ 0.008418f
C9665 net32 _094_ 0.027571f
C9666 net57 _068_ 0.029812f
C9667 _435_/a_2248_156# vdd 0.00571f
C9668 net73 _433_/a_36_151# 0.004541f
C9669 _112_ _083_ 0.003571f
C9670 _136_ _451_/a_1353_112# 0.058703f
C9671 net38 _444_/a_1204_472# 0.018432f
C9672 FILLER_0_17_72/a_2812_375# net14 0.018463f
C9673 net81 _136_ 0.021146f
C9674 _352_/a_49_472# _436_/a_36_151# 0.005127f
C9675 _074_ FILLER_0_3_221/a_1380_472# 0.001341f
C9676 _103_ _418_/a_2560_156# 0.002179f
C9677 fanout65/a_36_113# vdd 0.10473f
C9678 _443_/a_36_151# net13 0.001896f
C9679 _443_/a_1308_423# net23 0.034115f
C9680 FILLER_0_8_2/a_36_472# net40 0.002477f
C9681 output28/a_224_472# vss -0.0033f
C9682 net81 net62 0.245647f
C9683 FILLER_0_18_76/a_484_472# vss 0.005065f
C9684 FILLER_0_18_171/a_124_375# _098_ 0.032114f
C9685 ctln[2] net4 0.039098f
C9686 state\[0\] _070_ 0.009608f
C9687 _149_ _437_/a_36_151# 0.037766f
C9688 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_1020_375# 0.026339f
C9689 _392_/a_244_472# cal_count\[0\] 0.003287f
C9690 _070_ _370_/a_124_24# 0.00219f
C9691 _029_ net14 0.042032f
C9692 _326_/a_36_160# _128_ 0.02761f
C9693 net67 vdd 0.638702f
C9694 _053_ FILLER_0_5_54/a_36_472# 0.003309f
C9695 _426_/a_2665_112# net4 0.011288f
C9696 FILLER_0_11_124/a_124_375# _120_ 0.012164f
C9697 trim_val\[4\] _443_/a_2248_156# 0.050943f
C9698 output39/a_224_472# trim[1] 0.061797f
C9699 _086_ _061_ 0.152228f
C9700 net20 _080_ 0.093195f
C9701 net41 FILLER_0_17_38/a_124_375# 0.001109f
C9702 net54 FILLER_0_18_107/a_36_472# 0.002116f
C9703 _086_ _311_/a_66_473# 0.007295f
C9704 FILLER_0_5_109/a_572_375# _163_ 0.003096f
C9705 _126_ _389_/a_36_148# 0.007813f
C9706 _029_ _164_ 0.031781f
C9707 result[6] net60 0.094624f
C9708 output11/a_224_472# vss 0.083244f
C9709 FILLER_0_11_64/a_36_472# vdd 0.015144f
C9710 FILLER_0_11_64/a_124_375# vss 0.021069f
C9711 _070_ _247_/a_36_160# 0.0169f
C9712 FILLER_0_12_236/a_124_375# vdd 0.005169f
C9713 _010_ _009_ 0.030637f
C9714 output13/a_224_472# FILLER_0_0_130/a_124_375# 0.00363f
C9715 net38 _064_ 0.02996f
C9716 _335_/a_49_472# FILLER_0_15_180/a_572_375# 0.001126f
C9717 FILLER_0_14_91/a_124_375# vdd -0.010114f
C9718 FILLER_0_15_282/a_572_375# _417_/a_36_151# 0.001597f
C9719 FILLER_0_7_104/a_1020_375# _062_ 0.003073f
C9720 output12/a_224_472# _448_/a_36_151# 0.069748f
C9721 _442_/a_36_151# _031_ 0.013852f
C9722 _445_/a_36_151# vss 0.009726f
C9723 _445_/a_448_472# vdd 0.007946f
C9724 _000_ net75 0.096899f
C9725 FILLER_0_18_209/a_36_472# vss 0.005442f
C9726 FILLER_0_18_209/a_484_472# vdd 0.00367f
C9727 FILLER_0_21_28/a_484_472# vdd 0.011209f
C9728 _432_/a_2665_112# FILLER_0_17_200/a_124_375# 0.006271f
C9729 net50 FILLER_0_2_93/a_124_375# 0.007132f
C9730 net52 FILLER_0_2_93/a_36_472# 0.009026f
C9731 _035_ net41 0.048883f
C9732 FILLER_0_5_117/a_124_375# _119_ 0.002747f
C9733 _077_ FILLER_0_9_105/a_484_472# 0.002951f
C9734 _423_/a_36_151# _012_ 0.021631f
C9735 _052_ _216_/a_67_603# 0.006658f
C9736 output15/a_224_472# fanout50/a_36_160# 0.003531f
C9737 net38 net42 0.012245f
C9738 net32 net78 0.055231f
C9739 _161_ FILLER_0_6_177/a_572_375# 0.004064f
C9740 _162_ FILLER_0_6_177/a_36_472# 0.001723f
C9741 _077_ vss 1.071923f
C9742 FILLER_0_2_93/a_36_472# net49 0.001451f
C9743 FILLER_0_8_239/a_124_375# calibrate 0.008393f
C9744 net36 _451_/a_836_156# 0.007104f
C9745 _427_/a_1308_423# net23 0.004863f
C9746 net52 trim_mask\[2\] 0.036196f
C9747 net76 FILLER_0_5_198/a_572_375# 0.006974f
C9748 net68 fanout67/a_36_160# 0.02648f
C9749 FILLER_0_12_50/a_36_472# _120_ 0.005447f
C9750 _086_ _072_ 0.220767f
C9751 FILLER_0_13_212/a_572_375# _248_/a_36_68# 0.030745f
C9752 comp vdd 0.108153f
C9753 net27 net37 0.003648f
C9754 net81 _429_/a_2665_112# 0.012675f
C9755 net47 FILLER_0_6_37/a_36_472# 0.001161f
C9756 net62 net30 0.339141f
C9757 _155_ net14 0.10433f
C9758 _068_ _315_/a_244_497# 0.004768f
C9759 _186_ _184_ 0.047995f
C9760 FILLER_0_20_107/a_36_472# vss 0.004557f
C9761 net31 vdd 0.542738f
C9762 _002_ net82 0.034599f
C9763 FILLER_0_18_171/a_124_375# _432_/a_36_151# 0.001597f
C9764 trim_mask\[2\] net49 0.041781f
C9765 _064_ net66 0.304028f
C9766 net76 FILLER_0_2_177/a_572_375# 0.053951f
C9767 _075_ _077_ 0.004518f
C9768 output28/a_224_472# _416_/a_2248_156# 0.023576f
C9769 result[1] _416_/a_1308_423# 0.002597f
C9770 _009_ FILLER_0_23_282/a_36_472# 0.005974f
C9771 net24 vss 0.172755f
C9772 _112_ _425_/a_36_151# 0.032941f
C9773 net16 _450_/a_3129_107# 0.064714f
C9774 net72 _180_ 0.040135f
C9775 FILLER_0_12_136/a_36_472# _327_/a_36_472# 0.096379f
C9776 FILLER_0_16_57/a_124_375# _176_ 0.015872f
C9777 _131_ FILLER_0_18_37/a_1380_472# 0.035078f
C9778 _077_ _308_/a_124_24# 0.018118f
C9779 ctlp[4] net21 0.04068f
C9780 net53 _451_/a_1353_112# 0.028324f
C9781 _412_/a_448_472# output37/a_224_472# 0.001155f
C9782 _131_ FILLER_0_17_56/a_124_375# 0.001609f
C9783 _028_ net15 0.223301f
C9784 _425_/a_2665_112# net37 0.008519f
C9785 _128_ FILLER_0_10_214/a_36_472# 0.00186f
C9786 ctlp[6] vdd 0.207209f
C9787 _432_/a_1308_423# net80 0.030835f
C9788 FILLER_0_18_2/a_3172_472# _041_ 0.001503f
C9789 mask\[5\] FILLER_0_19_187/a_572_375# 0.005529f
C9790 net55 net40 0.043962f
C9791 _008_ ctlp[1] 0.002566f
C9792 FILLER_0_9_28/a_1916_375# net68 0.050307f
C9793 output47/a_224_472# FILLER_0_15_2/a_36_472# 0.035046f
C9794 _132_ FILLER_0_15_116/a_572_375# 0.003964f
C9795 _182_ cal_count\[1\] 0.166348f
C9796 result[0] FILLER_0_9_290/a_36_472# 0.020103f
C9797 _017_ _131_ 0.005879f
C9798 FILLER_0_14_81/a_124_375# vdd 0.023163f
C9799 _140_ _352_/a_665_69# 0.001363f
C9800 net60 _418_/a_36_151# 0.016348f
C9801 _053_ FILLER_0_6_79/a_36_472# 0.001777f
C9802 result[2] vdd 0.18482f
C9803 result[7] net60 0.778099f
C9804 output9/a_224_472# net59 0.051763f
C9805 _426_/a_1000_472# vdd 0.007031f
C9806 result[8] ctlp[1] 0.049662f
C9807 _028_ FILLER_0_6_90/a_572_375# 0.015802f
C9808 _303_/a_36_472# _098_ 0.021192f
C9809 net82 _370_/a_124_24# 0.001011f
C9810 _140_ _433_/a_2248_156# 0.003337f
C9811 FILLER_0_9_290/a_124_375# vdd 0.028723f
C9812 FILLER_0_12_220/a_932_472# _060_ 0.002471f
C9813 output38/a_224_472# net38 0.018882f
C9814 fanout67/a_36_160# net67 0.017633f
C9815 _106_ _293_/a_36_472# 0.04279f
C9816 FILLER_0_16_89/a_1380_472# vdd 0.010554f
C9817 _176_ FILLER_0_15_59/a_124_375# 0.007169f
C9818 _093_ _012_ 0.141641f
C9819 _163_ net14 0.040169f
C9820 FILLER_0_17_200/a_36_472# net21 0.036768f
C9821 _341_/a_49_472# net56 0.018486f
C9822 _065_ _441_/a_36_151# 0.00701f
C9823 ctln[7] trim_mask\[3\] 0.059414f
C9824 net81 net4 0.003327f
C9825 _413_/a_36_151# vss 0.003285f
C9826 _063_ vss 0.157186f
C9827 output27/a_224_472# FILLER_0_9_282/a_124_375# 0.029138f
C9828 _427_/a_796_472# net74 0.020124f
C9829 net55 FILLER_0_17_38/a_572_375# 0.007646f
C9830 net62 _417_/a_36_151# 0.044051f
C9831 net80 _339_/a_36_160# 0.016897f
C9832 _009_ _299_/a_36_472# 0.006927f
C9833 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_124_375# 0.012552f
C9834 net20 FILLER_0_15_235/a_36_472# 0.002227f
C9835 net64 FILLER_0_8_247/a_1380_472# 0.001021f
C9836 net73 FILLER_0_19_125/a_124_375# 0.005414f
C9837 output15/a_224_472# net14 0.003312f
C9838 net20 _104_ 0.482229f
C9839 net17 FILLER_0_12_28/a_36_472# 0.012286f
C9840 _163_ _164_ 0.021311f
C9841 net17 net40 1.095167f
C9842 _225_/a_36_160# vss 0.003244f
C9843 FILLER_0_6_47/a_1916_375# vdd -0.014642f
C9844 FILLER_0_6_47/a_1468_375# vss 0.003462f
C9845 _187_ _042_ 0.009526f
C9846 _069_ _043_ 0.04044f
C9847 _028_ net51 0.002321f
C9848 net50 _054_ 0.131493f
C9849 _231_/a_244_68# _059_ 0.004384f
C9850 FILLER_0_13_290/a_36_472# output30/a_224_472# 0.0323f
C9851 _076_ FILLER_0_5_148/a_36_472# 0.011563f
C9852 mask\[9\] FILLER_0_19_111/a_484_472# 0.041744f
C9853 net75 fanout75/a_36_113# 0.035159f
C9854 net20 vss 1.402494f
C9855 _193_/a_36_160# result[3] 0.002218f
C9856 FILLER_0_5_117/a_36_472# _153_ 0.028773f
C9857 mask\[4\] _346_/a_665_69# 0.001125f
C9858 output15/a_224_472# _164_ 0.031363f
C9859 FILLER_0_3_204/a_36_472# _088_ 0.004381f
C9860 _089_ _270_/a_36_472# 0.00437f
C9861 vss FILLER_0_12_196/a_36_472# 0.003551f
C9862 net4 _223_/a_36_160# 0.020711f
C9863 _128_ _161_ 0.027657f
C9864 _428_/a_2560_156# net53 0.002265f
C9865 _369_/a_36_68# _158_ 0.042315f
C9866 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_572_375# 0.086635f
C9867 _050_ _436_/a_1000_472# 0.02064f
C9868 output38/a_224_472# net66 0.148811f
C9869 _186_ _095_ 0.042856f
C9870 net27 FILLER_0_9_282/a_572_375# 0.002809f
C9871 vdd FILLER_0_6_231/a_36_472# 0.014642f
C9872 vss FILLER_0_6_231/a_572_375# 0.057794f
C9873 _086_ _331_/a_244_472# 0.001991f
C9874 _421_/a_36_151# vdd -0.053849f
C9875 net50 vss 1.178736f
C9876 FILLER_0_10_78/a_1020_375# _176_ 0.020379f
C9877 net74 _118_ 0.060991f
C9878 result[9] FILLER_0_24_274/a_572_375# 0.003576f
C9879 _128_ _129_ 0.029628f
C9880 FILLER_0_10_78/a_36_472# net52 0.014225f
C9881 net63 _435_/a_2248_156# 0.045342f
C9882 net67 _450_/a_1353_112# 0.025358f
C9883 ctlp[4] mask\[7\] 0.080163f
C9884 FILLER_0_18_107/a_2724_472# vss 0.003148f
C9885 FILLER_0_18_107/a_3172_472# vdd 0.004296f
C9886 _136_ FILLER_0_15_180/a_572_375# 0.001571f
C9887 net79 _070_ 0.009715f
C9888 result[8] FILLER_0_24_274/a_124_375# 0.00726f
C9889 _424_/a_2248_156# vdd -0.005751f
C9890 output32/a_224_472# vdd 0.082664f
C9891 _413_/a_36_151# FILLER_0_3_172/a_3260_375# 0.059049f
C9892 FILLER_0_1_192/a_124_375# vss 0.049811f
C9893 FILLER_0_1_192/a_36_472# vdd 0.011806f
C9894 net26 FILLER_0_23_44/a_124_375# 0.007775f
C9895 _320_/a_1120_472# state\[1\] 0.001998f
C9896 _265_/a_224_472# net59 0.001052f
C9897 net57 _113_ 0.012056f
C9898 mask\[4\] FILLER_0_18_177/a_2724_472# 0.014625f
C9899 _027_ FILLER_0_18_76/a_484_472# 0.00705f
C9900 net52 _441_/a_2560_156# 0.004721f
C9901 net50 _441_/a_2248_156# 0.027849f
C9902 mask\[3\] FILLER_0_18_177/a_1828_472# 0.004274f
C9903 net15 net47 0.035839f
C9904 _277_/a_36_160# vdd 0.115507f
C9905 _308_/a_124_24# net50 0.02221f
C9906 FILLER_0_12_136/a_572_375# _427_/a_1308_423# 0.001238f
C9907 _029_ _153_ 0.023421f
C9908 FILLER_0_16_57/a_1468_375# net15 0.012909f
C9909 FILLER_0_8_138/a_36_472# _077_ 0.005953f
C9910 _417_/a_2560_156# net30 0.049334f
C9911 _415_/a_1308_423# net27 0.02437f
C9912 _049_ FILLER_0_22_128/a_2812_375# 0.001905f
C9913 _057_ _306_/a_36_68# 0.019072f
C9914 mask\[4\] FILLER_0_17_218/a_484_472# 0.001232f
C9915 _449_/a_36_151# _043_ 0.001572f
C9916 _340_/a_36_160# FILLER_0_20_169/a_124_375# 0.005494f
C9917 FILLER_0_21_125/a_36_472# mask\[7\] 0.00344f
C9918 net15 _012_ 0.043755f
C9919 _074_ FILLER_0_6_177/a_36_472# 0.045576f
C9920 FILLER_0_19_134/a_36_472# _145_ 0.080913f
C9921 _431_/a_2560_156# _137_ 0.002967f
C9922 FILLER_0_5_72/a_572_375# vss 0.006023f
C9923 FILLER_0_5_72/a_1020_375# vdd 0.009501f
C9924 net21 _434_/a_2248_156# 0.001467f
C9925 mask\[3\] _094_ 0.00554f
C9926 mask\[3\] FILLER_0_17_218/a_572_375# 0.015907f
C9927 _050_ FILLER_0_22_128/a_124_375# 0.002607f
C9928 FILLER_0_1_98/a_36_472# net14 0.023583f
C9929 net69 FILLER_0_2_111/a_484_472# 0.010567f
C9930 _031_ FILLER_0_2_111/a_1468_375# 0.013595f
C9931 net14 FILLER_0_4_91/a_36_472# 0.005793f
C9932 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_484_472# 0.013277f
C9933 _420_/a_448_472# net77 0.001276f
C9934 net61 _422_/a_2665_112# 0.023601f
C9935 _098_ FILLER_0_19_171/a_572_375# 0.001946f
C9936 FILLER_0_5_54/a_572_375# _029_ 0.00494f
C9937 _413_/a_1204_472# net82 0.00291f
C9938 calibrate FILLER_0_8_156/a_36_472# 0.001283f
C9939 _122_ FILLER_0_8_156/a_572_375# 0.002572f
C9940 _315_/a_36_68# _121_ 0.031617f
C9941 _432_/a_2665_112# mask\[3\] 0.011428f
C9942 _441_/a_36_151# _440_/a_448_472# 0.002538f
C9943 FILLER_0_16_73/a_124_375# net55 0.007695f
C9944 _414_/a_796_472# _053_ 0.008213f
C9945 net16 trim_val\[0\] 0.00463f
C9946 _035_ FILLER_0_4_49/a_124_375# 0.00215f
C9947 fanout81/a_36_160# vss 0.02458f
C9948 FILLER_0_9_223/a_124_375# _076_ 0.004399f
C9949 _028_ FILLER_0_7_104/a_36_472# 0.006408f
C9950 _446_/a_1308_423# net40 0.038281f
C9951 _426_/a_36_151# FILLER_0_8_247/a_572_375# 0.059049f
C9952 _012_ FILLER_0_23_44/a_1380_472# 0.001572f
C9953 output13/a_224_472# net52 0.018089f
C9954 vdd _380_/a_224_472# 0.001733f
C9955 _081_ FILLER_0_5_148/a_36_472# 0.020403f
C9956 FILLER_0_21_150/a_124_375# _433_/a_2665_112# 0.029834f
C9957 FILLER_0_16_255/a_124_375# vdd 0.029925f
C9958 _421_/a_1308_423# net19 0.055838f
C9959 result[4] _417_/a_2248_156# 0.001436f
C9960 _119_ _114_ 0.001581f
C9961 _074_ _316_/a_124_24# 0.018608f
C9962 net15 FILLER_0_15_59/a_484_472# 0.015199f
C9963 FILLER_0_5_128/a_572_375# net47 0.010055f
C9964 FILLER_0_10_78/a_124_375# vss 0.006775f
C9965 net36 FILLER_0_15_180/a_484_472# 0.00702f
C9966 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_124_375# 0.012001f
C9967 net39 net47 0.13057f
C9968 _144_ net54 0.095482f
C9969 _253_/a_36_68# _073_ 0.027664f
C9970 net47 net51 0.007412f
C9971 _328_/a_36_113# vss 0.044028f
C9972 result[6] FILLER_0_23_290/a_124_375# 0.001492f
C9973 _005_ net18 0.073455f
C9974 net16 _445_/a_2248_156# 0.003321f
C9975 net50 FILLER_0_5_88/a_124_375# 0.03181f
C9976 FILLER_0_22_177/a_932_472# _435_/a_36_151# 0.001723f
C9977 _372_/a_3662_472# _122_ 0.002653f
C9978 output34/a_224_472# _102_ 0.008577f
C9979 _091_ FILLER_0_15_212/a_1020_375# 0.00799f
C9980 _432_/a_2248_156# _139_ 0.002904f
C9981 net21 _202_/a_36_160# 0.09166f
C9982 net15 net74 0.05717f
C9983 _155_ _153_ 0.033366f
C9984 net34 FILLER_0_22_128/a_2276_472# 0.005532f
C9985 FILLER_0_15_72/a_484_472# vss 0.010761f
C9986 _069_ FILLER_0_18_209/a_484_472# 0.013944f
C9987 FILLER_0_15_150/a_124_375# _427_/a_36_151# 0.001822f
C9988 _127_ FILLER_0_9_142/a_124_375# 0.005447f
C9989 net43 FILLER_0_20_15/a_36_472# 0.002803f
C9990 FILLER_0_8_107/a_124_375# FILLER_0_10_107/a_36_472# 0.0027f
C9991 _258_/a_36_160# net37 0.006865f
C9992 FILLER_0_21_150/a_124_375# vdd 0.020581f
C9993 FILLER_0_3_2/a_36_472# vss 0.004076f
C9994 _093_ FILLER_0_19_155/a_36_472# 0.001737f
C9995 net73 mask\[9\] 0.383862f
C9996 _015_ net64 1.212892f
C9997 _431_/a_36_151# net70 0.031018f
C9998 net26 vdd 0.487733f
C9999 _035_ _446_/a_796_472# 0.013039f
C10000 _308_/a_692_472# _115_ 0.001485f
C10001 net55 FILLER_0_17_56/a_36_472# 0.019193f
C10002 cal_itt\[3\] vss 0.15522f
C10003 _133_ FILLER_0_10_107/a_484_472# 0.001798f
C10004 _128_ _056_ 0.026612f
C10005 FILLER_0_23_88/a_36_472# net14 0.003077f
C10006 _104_ _009_ 0.284256f
C10007 _412_/a_2665_112# net59 0.055415f
C10008 FILLER_0_12_50/a_124_375# vdd 0.039185f
C10009 fanout81/a_36_160# fanout76/a_36_160# 0.01081f
C10010 output7/a_224_472# output40/a_224_472# 0.038066f
C10011 _061_ _311_/a_66_473# 0.030169f
C10012 _428_/a_1204_472# vdd 0.001231f
C10013 _077_ FILLER_0_10_78/a_572_375# 0.001886f
C10014 _071_ _225_/a_36_160# 0.002808f
C10015 _098_ _433_/a_1204_472# 0.014374f
C10016 FILLER_0_5_128/a_572_375# net74 0.050735f
C10017 FILLER_0_7_195/a_36_472# calibrate 0.010951f
C10018 _009_ vss 0.105833f
C10019 valid net2 0.062523f
C10020 _432_/a_1204_472# vdd 0.004019f
C10021 output47/a_224_472# _398_/a_36_113# 0.001605f
C10022 trimb[3] ctlp[0] 0.384753f
C10023 _068_ FILLER_0_9_142/a_36_472# 0.009073f
C10024 _075_ cal_itt\[3\] 0.731221f
C10025 _086_ _321_/a_3662_472# 0.002598f
C10026 _394_/a_728_93# vdd 0.006211f
C10027 _394_/a_1336_472# vss 0.040135f
C10028 cal_count\[1\] _040_ 0.019478f
C10029 _065_ net16 0.068602f
C10030 _163_ _153_ 0.243815f
C10031 _449_/a_36_151# FILLER_0_11_64/a_36_472# 0.046516f
C10032 FILLER_0_24_274/a_932_472# FILLER_0_23_282/a_36_472# 0.05841f
C10033 _002_ net21 0.056631f
C10034 FILLER_0_11_142/a_484_472# net23 0.006988f
C10035 _081_ FILLER_0_6_177/a_36_472# 0.00483f
C10036 FILLER_0_7_195/a_36_472# net21 0.005469f
C10037 _422_/a_1000_472# _009_ 0.007191f
C10038 _408_/a_1336_472# net40 0.020063f
C10039 trimb[1] net38 0.161478f
C10040 vss _039_ 0.180364f
C10041 FILLER_0_14_81/a_36_472# _043_ 0.001714f
C10042 FILLER_0_8_247/a_124_375# FILLER_0_8_239/a_124_375# 0.003732f
C10043 _132_ FILLER_0_14_107/a_932_472# 0.014911f
C10044 _093_ _177_ 0.001194f
C10045 FILLER_0_19_47/a_572_375# FILLER_0_18_53/a_36_472# 0.001684f
C10046 output42/a_224_472# net42 0.117956f
C10047 _414_/a_36_151# FILLER_0_7_195/a_36_472# 0.001723f
C10048 _128_ _068_ 0.863174f
C10049 _131_ cal_count\[3\] 0.035391f
C10050 _091_ FILLER_0_12_220/a_36_472# 0.003655f
C10051 output12/a_224_472# vss 0.013728f
C10052 net1 _083_ 0.30074f
C10053 ctln[1] net75 0.159105f
C10054 FILLER_0_20_177/a_1468_375# _098_ 0.012889f
C10055 result[7] FILLER_0_23_290/a_124_375# 0.018455f
C10056 net62 fanout78/a_36_113# 0.014177f
C10057 net55 _452_/a_1040_527# 0.021721f
C10058 FILLER_0_5_164/a_572_375# _386_/a_848_380# 0.001121f
C10059 _052_ FILLER_0_18_61/a_124_375# 0.006877f
C10060 _068_ _311_/a_692_473# 0.002377f
C10061 _072_ _061_ 0.448032f
C10062 net20 _419_/a_1000_472# 0.022734f
C10063 state\[0\] calibrate 0.001061f
C10064 _081_ _316_/a_124_24# 0.011421f
C10065 _072_ _311_/a_66_473# 0.031716f
C10066 _427_/a_36_151# FILLER_0_14_123/a_36_472# 0.004032f
C10067 _302_/a_224_472# _012_ 0.002675f
C10068 _062_ net37 0.082701f
C10069 _173_ net51 0.016607f
C10070 trim_mask\[1\] FILLER_0_6_47/a_1380_472# 0.006166f
C10071 _009_ _107_ 0.027726f
C10072 FILLER_0_18_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001684f
C10073 _360_/a_36_160# vdd 0.006439f
C10074 _102_ _099_ 0.151018f
C10075 _144_ _350_/a_49_472# 0.033348f
C10076 FILLER_0_15_116/a_36_472# _136_ 0.003818f
C10077 FILLER_0_13_228/a_124_375# vdd -0.007362f
C10078 FILLER_0_10_247/a_124_375# _100_ 0.001804f
C10079 _079_ _073_ 0.234533f
C10080 _322_/a_848_380# vss 0.026127f
C10081 net18 _416_/a_448_472# 0.05521f
C10082 mask\[5\] FILLER_0_20_169/a_36_472# 0.016469f
C10083 FILLER_0_8_107/a_36_472# _053_ 0.013669f
C10084 _095_ _225_/a_36_160# 0.001084f
C10085 FILLER_0_15_10/a_124_375# vdd 0.021578f
C10086 FILLER_0_2_101/a_36_472# vss 0.004743f
C10087 fanout61/a_36_113# FILLER_0_21_286/a_572_375# 0.015816f
C10088 _430_/a_2560_156# mask\[2\] 0.010268f
C10089 _126_ FILLER_0_12_196/a_124_375# 0.001392f
C10090 net35 FILLER_0_22_128/a_36_472# 0.00784f
C10091 _102_ _419_/a_2248_156# 0.001679f
C10092 net17 _452_/a_1040_527# 0.034254f
C10093 _285_/a_36_472# _094_ 0.045394f
C10094 fanout79/a_36_160# _060_ 0.005814f
C10095 _247_/a_36_160# net21 0.002254f
C10096 net75 _074_ 1.343862f
C10097 _265_/a_244_68# vss 0.009604f
C10098 net41 FILLER_0_20_31/a_124_375# 0.049106f
C10099 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_484_472# 0.026657f
C10100 _281_/a_234_472# _097_ 0.004169f
C10101 FILLER_0_4_197/a_36_472# net76 0.003914f
C10102 net60 _419_/a_1204_472# 0.023544f
C10103 net61 _419_/a_2665_112# 0.022394f
C10104 mask\[5\] FILLER_0_18_177/a_1380_472# 0.001063f
C10105 _013_ net36 0.032392f
C10106 _444_/a_1308_423# net40 0.043396f
C10107 net47 clkc 0.002956f
C10108 net20 FILLER_0_12_220/a_124_375# 0.003161f
C10109 net54 FILLER_0_22_128/a_572_375# 0.048634f
C10110 FILLER_0_17_104/a_932_472# vdd 0.020019f
C10111 _070_ FILLER_0_9_105/a_124_375# 0.017687f
C10112 _013_ FILLER_0_18_37/a_932_472# 0.010651f
C10113 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_124_375# 0.003732f
C10114 FILLER_0_17_72/a_2364_375# _136_ 0.047331f
C10115 _130_ _114_ 0.002404f
C10116 FILLER_0_8_24/a_572_375# net40 0.038492f
C10117 _114_ _161_ 0.024297f
C10118 FILLER_0_1_98/a_36_472# _153_ 0.001463f
C10119 _078_ vdd 0.181583f
C10120 _105_ result[6] 0.001477f
C10121 FILLER_0_18_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001597f
C10122 _411_/a_36_151# output10/a_224_472# 0.001362f
C10123 _374_/a_36_68# _058_ 0.010442f
C10124 _073_ cal_itt\[1\] 0.058541f
C10125 net55 FILLER_0_18_53/a_36_472# 0.00953f
C10126 _413_/a_796_472# _002_ 0.009261f
C10127 net50 _036_ 0.002727f
C10128 _057_ net22 0.163773f
C10129 FILLER_0_12_124/a_124_375# _126_ 0.02249f
C10130 FILLER_0_23_290/a_36_472# vss 0.0074f
C10131 mask\[2\] FILLER_0_15_212/a_1380_472# 0.001225f
C10132 _132_ FILLER_0_18_107/a_1916_375# 0.019011f
C10133 FILLER_0_9_223/a_484_472# state\[0\] 0.007034f
C10134 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3172_472# 0.013277f
C10135 _096_ _320_/a_224_472# 0.001285f
C10136 FILLER_0_16_107/a_484_472# net36 0.003765f
C10137 trim_mask\[2\] net40 0.401672f
C10138 FILLER_0_20_177/a_124_375# FILLER_0_20_169/a_124_375# 0.003732f
C10139 _050_ FILLER_0_22_107/a_36_472# 0.001098f
C10140 FILLER_0_20_193/a_36_472# vss 0.001978f
C10141 FILLER_0_20_193/a_484_472# vdd 0.00749f
C10142 FILLER_0_7_162/a_36_472# _074_ 0.003809f
C10143 result[9] _417_/a_2248_156# 0.046399f
C10144 FILLER_0_17_72/a_1828_472# _131_ 0.004882f
C10145 _431_/a_2248_156# FILLER_0_15_142/a_484_472# 0.016128f
C10146 net16 _034_ 0.096088f
C10147 FILLER_0_19_111/a_36_472# net14 0.00143f
C10148 _420_/a_796_472# _009_ 0.012395f
C10149 net73 _022_ 0.003246f
C10150 output44/a_224_472# FILLER_0_18_2/a_124_375# 0.001168f
C10151 _133_ _058_ 0.092697f
C10152 FILLER_0_12_136/a_932_472# vss 0.008682f
C10153 FILLER_0_12_136/a_1380_472# vdd 0.006419f
C10154 net72 vss 0.472104f
C10155 FILLER_0_15_116/a_36_472# net53 0.005099f
C10156 net68 FILLER_0_8_37/a_124_375# 0.004818f
C10157 _178_ net72 0.007093f
C10158 mask\[5\] result[8] 0.003797f
C10159 _414_/a_2248_156# _053_ 0.013478f
C10160 result[7] FILLER_0_24_274/a_484_472# 0.006641f
C10161 _415_/a_2248_156# net18 0.057604f
C10162 _136_ _356_/a_36_472# 0.004667f
C10163 _101_ _094_ 0.304499f
C10164 FILLER_0_18_107/a_3260_375# FILLER_0_19_134/a_124_375# 0.026339f
C10165 FILLER_0_17_161/a_124_375# _098_ 0.002013f
C10166 FILLER_0_5_54/a_484_472# vss 0.001929f
C10167 FILLER_0_5_54/a_932_472# vdd 0.003166f
C10168 _413_/a_1204_472# net21 0.011236f
C10169 result[6] output19/a_224_472# 0.001526f
C10170 trim_mask\[4\] net47 0.264421f
C10171 _176_ _129_ 0.036112f
C10172 _404_/a_36_472# _183_ 0.002637f
C10173 FILLER_0_7_104/a_1020_375# _153_ 0.026997f
C10174 FILLER_0_18_177/a_1468_375# FILLER_0_20_177/a_1380_472# 0.0027f
C10175 _093_ _438_/a_448_472# 0.0106f
C10176 _442_/a_2665_112# vss 0.001727f
C10177 _442_/a_2560_156# vdd 0.006195f
C10178 _442_/a_36_151# _158_ 0.001257f
C10179 FILLER_0_10_37/a_36_472# net51 0.002346f
C10180 mask\[9\] _438_/a_36_151# 0.060632f
C10181 _030_ _367_/a_36_68# 0.015584f
C10182 net20 FILLER_0_12_236/a_36_472# 0.003143f
C10183 _149_ FILLER_0_20_87/a_36_472# 0.001938f
C10184 _091_ _139_ 0.05535f
C10185 _079_ FILLER_0_5_212/a_36_472# 0.005671f
C10186 net15 FILLER_0_6_47/a_1828_472# 0.014911f
C10187 FILLER_0_10_28/a_124_375# net17 0.00917f
C10188 FILLER_0_18_177/a_2364_375# vdd 0.020562f
C10189 _096_ _114_ 0.066848f
C10190 _449_/a_2248_156# _067_ 0.040648f
C10191 cal_itt\[3\] FILLER_0_5_198/a_36_472# 0.07099f
C10192 _450_/a_1040_527# _039_ 0.015478f
C10193 FILLER_0_11_101/a_124_375# cal_count\[3\] 0.00419f
C10194 _186_ _185_ 0.007962f
C10195 FILLER_0_17_133/a_36_472# _137_ 0.001963f
C10196 net75 _425_/a_796_472# 0.001146f
C10197 net16 FILLER_0_18_37/a_1020_375# 0.005406f
C10198 _095_ FILLER_0_15_72/a_484_472# 0.002306f
C10199 FILLER_0_15_282/a_572_375# _006_ 0.001054f
C10200 net75 _081_ 0.060976f
C10201 _399_/a_224_472# net16 0.003817f
C10202 net46 net43 0.215092f
C10203 net69 _441_/a_36_151# 0.035817f
C10204 FILLER_0_16_89/a_124_375# _177_ 0.008257f
C10205 _415_/a_448_472# net64 0.02484f
C10206 _076_ _059_ 1.03702f
C10207 _028_ _154_ 0.174927f
C10208 net41 FILLER_0_19_28/a_572_375# 0.040551f
C10209 net73 FILLER_0_18_107/a_484_472# 0.0052f
C10210 mask\[7\] FILLER_0_22_128/a_2364_375# 0.003632f
C10211 net17 FILLER_0_20_15/a_1468_375# 0.010099f
C10212 _163_ FILLER_0_5_148/a_36_472# 0.002454f
C10213 _033_ vdd 0.509957f
C10214 _129_ _124_ 0.010499f
C10215 cal_count\[2\] FILLER_0_15_10/a_36_472# 0.015502f
C10216 FILLER_0_15_116/a_124_375# FILLER_0_14_107/a_1020_375# 0.026339f
C10217 net36 net71 0.148833f
C10218 FILLER_0_19_125/a_124_375# _433_/a_36_151# 0.001597f
C10219 _415_/a_36_151# net62 0.00514f
C10220 FILLER_0_24_290/a_124_375# vdd 0.026739f
C10221 net53 _427_/a_36_151# 0.13192f
C10222 net56 _427_/a_2665_112# 0.012193f
C10223 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1380_472# 0.013276f
C10224 _057_ vdd 0.801978f
C10225 state\[1\] FILLER_0_12_196/a_124_375# 0.063785f
C10226 _248_/a_36_68# _090_ 0.041161f
C10227 _448_/a_36_151# net22 0.027581f
C10228 _053_ _251_/a_906_472# 0.001696f
C10229 _428_/a_2248_156# _043_ 0.011841f
C10230 net75 net65 0.135447f
C10231 trim_val\[3\] trim_mask\[3\] 0.48462f
C10232 fanout74/a_36_113# vdd 0.099021f
C10233 cal_itt\[2\] FILLER_0_3_221/a_1020_375# 0.010951f
C10234 net52 _439_/a_448_472# 0.042072f
C10235 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_124_375# 0.012222f
C10236 _008_ result[5] 0.165753f
C10237 _335_/a_257_69# mask\[1\] 0.001543f
C10238 _021_ FILLER_0_18_171/a_36_472# 0.103755f
C10239 FILLER_0_18_2/a_484_472# _452_/a_2225_156# 0.019521f
C10240 net27 _100_ 0.006783f
C10241 _250_/a_36_68# vdd 0.014409f
C10242 net74 trim_mask\[4\] 0.548293f
C10243 net20 _106_ 0.050151f
C10244 _176_ _394_/a_1936_472# 0.001255f
C10245 _128_ _113_ 0.002117f
C10246 en_co_clk cal_count\[3\] 0.001359f
C10247 _180_ vdd 0.176915f
C10248 _428_/a_1000_472# _095_ 0.001101f
C10249 _412_/a_448_472# net58 0.044616f
C10250 _432_/a_36_151# FILLER_0_17_161/a_124_375# 0.035117f
C10251 FILLER_0_18_171/a_124_375# net80 0.024341f
C10252 net79 net21 0.645949f
C10253 net74 net47 0.030815f
C10254 net62 net64 0.078454f
C10255 _443_/a_2665_112# _170_ 0.019855f
C10256 net15 _440_/a_1000_472# 0.056791f
C10257 state\[2\] FILLER_0_13_142/a_484_472# 0.004186f
C10258 net53 FILLER_0_13_142/a_1380_472# 0.041222f
C10259 _091_ FILLER_0_13_212/a_1468_375# 0.003576f
C10260 _015_ FILLER_0_8_247/a_572_375# 0.00706f
C10261 _421_/a_36_151# net77 0.028951f
C10262 FILLER_0_3_78/a_124_375# vss 0.004739f
C10263 FILLER_0_3_78/a_572_375# vdd 0.014442f
C10264 _114_ _056_ 0.034246f
C10265 FILLER_0_2_127/a_124_375# vdd 0.013496f
C10266 _394_/a_1336_472# _095_ 0.031869f
C10267 FILLER_0_24_274/a_932_472# vss 0.001001f
C10268 mask\[5\] _343_/a_49_472# 0.002228f
C10269 _119_ FILLER_0_7_104/a_1380_472# 0.002603f
C10270 net58 net19 0.044785f
C10271 _104_ net33 0.037008f
C10272 _448_/a_2560_156# _037_ 0.011661f
C10273 vss trim[2] 0.026644f
C10274 FILLER_0_7_162/a_36_472# _081_ 0.002493f
C10275 FILLER_0_22_128/a_36_472# vdd 0.004601f
C10276 FILLER_0_22_128/a_3260_375# vss 0.006346f
C10277 _093_ net70 0.001888f
C10278 _348_/a_665_69# _146_ 0.001153f
C10279 FILLER_0_7_162/a_124_375# _074_ 0.007213f
C10280 _175_ _040_ 0.00133f
C10281 output46/a_224_472# FILLER_0_21_28/a_36_472# 0.010684f
C10282 net33 vss 0.674927f
C10283 _372_/a_170_472# net23 0.025555f
C10284 output15/a_224_472# FILLER_0_0_96/a_36_472# 0.023414f
C10285 net20 _426_/a_2248_156# 0.007902f
C10286 net56 FILLER_0_18_139/a_124_375# 0.00281f
C10287 FILLER_0_12_20/a_124_375# net6 0.003726f
C10288 _326_/a_36_160# FILLER_0_7_104/a_1380_472# 0.002051f
C10289 _079_ FILLER_0_3_172/a_2276_472# 0.00261f
C10290 _425_/a_448_472# net19 0.034226f
C10291 net60 _007_ 0.025806f
C10292 mask\[4\] _092_ 0.072581f
C10293 _412_/a_448_472# _082_ 0.022743f
C10294 result[8] output20/a_224_472# 0.038114f
C10295 net76 _083_ 0.002446f
C10296 _412_/a_2248_156# net59 0.008792f
C10297 net82 FILLER_0_3_172/a_1916_375# 0.010202f
C10298 _412_/a_448_472# net82 0.030379f
C10299 _260_/a_36_68# net59 0.004346f
C10300 FILLER_0_15_142/a_124_375# net74 0.005931f
C10301 FILLER_0_13_228/a_36_472# _043_ 0.02119f
C10302 FILLER_0_9_28/a_484_472# net16 0.021584f
C10303 _114_ FILLER_0_11_101/a_572_375# 0.051108f
C10304 FILLER_0_17_38/a_484_472# vss 0.001229f
C10305 _235_/a_67_603# _447_/a_36_151# 0.038675f
C10306 _114_ _068_ 1.097353f
C10307 _256_/a_716_497# net4 0.001936f
C10308 trim_mask\[4\] _159_ 0.049552f
C10309 _065_ _030_ 0.001499f
C10310 FILLER_0_3_172/a_1020_375# net65 0.006035f
C10311 net19 _082_ 0.029316f
C10312 _127_ _085_ 0.00179f
C10313 _446_/a_36_151# vdd 0.06703f
C10314 net79 _418_/a_448_472# 0.034736f
C10315 net82 net19 1.14585f
C10316 vss FILLER_0_3_212/a_36_472# 0.00838f
C10317 FILLER_0_6_177/a_36_472# _163_ 0.025039f
C10318 _159_ net47 0.01358f
C10319 _449_/a_36_151# FILLER_0_12_50/a_124_375# 0.017882f
C10320 net62 _006_ 0.136418f
C10321 _376_/a_36_160# _163_ 0.006811f
C10322 net16 _453_/a_36_151# 0.001634f
C10323 _322_/a_124_24# _126_ 0.019609f
C10324 result[7] FILLER_0_23_282/a_124_375# 0.016009f
C10325 net72 _401_/a_36_68# 0.006818f
C10326 FILLER_0_17_282/a_124_375# vss 0.024404f
C10327 FILLER_0_17_282/a_36_472# vdd 0.107351f
C10328 _081_ _059_ 0.04053f
C10329 _316_/a_848_380# _122_ 0.002234f
C10330 _316_/a_692_472# calibrate 0.006232f
C10331 _161_ _267_/a_36_472# 0.043279f
C10332 net79 FILLER_0_21_286/a_572_375# 0.001476f
C10333 FILLER_0_18_2/a_124_375# vdd 0.008721f
C10334 net4 net59 0.102012f
C10335 FILLER_0_9_142/a_124_375# _118_ 0.06224f
C10336 _429_/a_2665_112# net64 0.013014f
C10337 _306_/a_36_68# vss 0.008326f
C10338 trim_mask\[4\] _154_ 0.014658f
C10339 net27 FILLER_0_8_263/a_124_375# 0.016669f
C10340 _431_/a_448_472# net36 0.010914f
C10341 _089_ _081_ 0.002206f
C10342 _449_/a_36_151# _394_/a_728_93# 0.002727f
C10343 net33 _107_ 0.001322f
C10344 net2 cal_itt\[1\] 0.284695f
C10345 net31 FILLER_0_16_255/a_36_472# 0.003056f
C10346 FILLER_0_15_150/a_124_375# mask\[2\] 0.002588f
C10347 net27 FILLER_0_14_235/a_124_375# 0.002299f
C10348 _448_/a_36_151# vdd 0.133302f
C10349 net47 _154_ 0.055128f
C10350 _310_/a_49_472# vdd 0.043164f
C10351 FILLER_0_23_60/a_36_472# vdd 0.090554f
C10352 FILLER_0_23_60/a_124_375# vss 0.004081f
C10353 mask\[9\] FILLER_0_20_98/a_36_472# 0.005917f
C10354 cal_count\[2\] _182_ 0.044348f
C10355 net55 FILLER_0_19_28/a_36_472# 0.001572f
C10356 FILLER_0_3_142/a_124_375# trim_mask\[4\] 0.002514f
C10357 _053_ net76 0.022571f
C10358 net20 _421_/a_1308_423# 0.012036f
C10359 FILLER_0_7_72/a_572_375# _053_ 0.014569f
C10360 _119_ _359_/a_36_488# 0.003263f
C10361 FILLER_0_18_100/a_124_375# vss 0.025563f
C10362 FILLER_0_18_100/a_36_472# vdd 0.012574f
C10363 _442_/a_36_151# net23 0.00157f
C10364 FILLER_0_4_144/a_484_472# vss 0.033414f
C10365 net78 _094_ 0.050187f
C10366 _016_ vdd 0.114288f
C10367 _379_/a_36_472# _160_ 0.023459f
C10368 FILLER_0_5_117/a_124_375# FILLER_0_4_107/a_1380_472# 0.001684f
C10369 FILLER_0_9_28/a_2364_375# vdd 0.004562f
C10370 net55 _423_/a_2248_156# 0.001188f
C10371 _176_ FILLER_0_11_101/a_572_375# 0.00389f
C10372 _008_ _199_/a_36_160# 0.002015f
C10373 FILLER_0_14_99/a_124_375# net14 0.04852f
C10374 net54 FILLER_0_22_107/a_484_472# 0.005897f
C10375 net63 FILLER_0_20_193/a_484_472# 0.015851f
C10376 FILLER_0_14_263/a_124_375# vdd 0.026205f
C10377 _010_ vdd 0.121474f
C10378 _386_/a_124_24# _169_ 0.02709f
C10379 net27 _060_ 0.045136f
C10380 FILLER_0_17_72/a_572_375# vss 0.008057f
C10381 FILLER_0_17_72/a_1020_375# vdd 0.002541f
C10382 FILLER_0_18_2/a_484_472# net44 0.047503f
C10383 net81 _426_/a_1308_423# 0.002332f
C10384 FILLER_0_17_161/a_36_472# _137_ 0.013985f
C10385 FILLER_0_4_177/a_36_472# trim_val\[4\] 0.001889f
C10386 net4 _122_ 0.03487f
C10387 FILLER_0_4_107/a_1020_375# vdd 0.025121f
C10388 FILLER_0_7_72/a_3172_472# trim_mask\[0\] 0.001438f
C10389 net74 _159_ 0.129233f
C10390 FILLER_0_9_270/a_572_375# vdd 0.02345f
C10391 FILLER_0_19_28/a_36_472# net17 0.009277f
C10392 net38 FILLER_0_20_2/a_36_472# 0.002204f
C10393 _230_/a_244_68# _060_ 0.002039f
C10394 net17 _450_/a_36_151# 0.006157f
C10395 FILLER_0_21_125/a_36_472# _354_/a_49_472# 0.063744f
C10396 FILLER_0_16_241/a_124_375# _099_ 0.040547f
C10397 net52 FILLER_0_2_111/a_124_375# 0.00483f
C10398 FILLER_0_4_197/a_572_375# net59 0.001512f
C10399 ctlp[2] _422_/a_448_472# 0.011383f
C10400 _091_ _429_/a_1308_423# 0.031247f
C10401 _063_ _166_ 0.025402f
C10402 net4 net64 0.060449f
C10403 output34/a_224_472# _198_/a_67_603# 0.00179f
C10404 net63 FILLER_0_18_177/a_2364_375# 0.009893f
C10405 net52 _440_/a_36_151# 0.01571f
C10406 net57 FILLER_0_16_154/a_1380_472# 0.041458f
C10407 net60 _421_/a_796_472# 0.002046f
C10408 net74 _154_ 0.002976f
C10409 valid cal_itt\[1\] 0.011576f
C10410 _449_/a_2665_112# net74 0.001185f
C10411 _401_/a_244_472# _180_ 0.001689f
C10412 _065_ trim_mask\[3\] 0.020092f
C10413 FILLER_0_16_89/a_36_472# _131_ 0.013616f
C10414 net53 FILLER_0_14_107/a_1380_472# 0.059367f
C10415 trim[0] _034_ 0.044322f
C10416 FILLER_0_9_28/a_3260_375# _077_ 0.01495f
C10417 net79 mask\[1\] 0.029512f
C10418 FILLER_0_12_136/a_484_472# _126_ 0.014541f
C10419 _077_ cal_count\[0\] 0.018501f
C10420 FILLER_0_23_282/a_36_472# vdd 0.106034f
C10421 FILLER_0_23_282/a_572_375# vss 0.058599f
C10422 _438_/a_2560_156# vdd 0.001166f
C10423 _438_/a_2665_112# vss 0.001389f
C10424 FILLER_0_13_142/a_36_472# vdd 0.104785f
C10425 FILLER_0_13_142/a_1468_375# vss 0.00614f
C10426 net66 _440_/a_796_472# 0.002718f
C10427 net49 _440_/a_36_151# 0.021133f
C10428 _127_ _062_ 0.020537f
C10429 _131_ FILLER_0_17_64/a_36_472# 0.002638f
C10430 net52 FILLER_0_5_72/a_932_472# 0.008749f
C10431 FILLER_0_4_197/a_1380_472# net82 0.003084f
C10432 FILLER_0_19_142/a_124_375# vdd 0.022448f
C10433 net72 _095_ 0.136566f
C10434 net1 fanout59/a_36_160# 0.002325f
C10435 FILLER_0_17_56/a_572_375# FILLER_0_18_61/a_36_472# 0.001597f
C10436 cal_count\[3\] _090_ 0.243462f
C10437 _447_/a_36_151# vdd 0.067176f
C10438 _048_ FILLER_0_18_209/a_124_375# 0.001615f
C10439 _087_ FILLER_0_5_172/a_36_472# 0.00443f
C10440 _053_ net68 0.239882f
C10441 _086_ net23 0.037804f
C10442 net29 net30 0.053996f
C10443 result[2] output30/a_224_472# 0.045862f
C10444 _273_/a_36_68# _128_ 0.005719f
C10445 ctlp[2] _108_ 0.034027f
C10446 _152_ FILLER_0_5_136/a_36_472# 0.049485f
C10447 _137_ FILLER_0_16_154/a_124_375# 0.007998f
C10448 _031_ _157_ 0.104339f
C10449 net54 _433_/a_448_472# 0.008777f
C10450 ctlp[2] net19 0.017506f
C10451 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_572_375# 0.001597f
C10452 _164_ FILLER_0_6_47/a_932_472# 0.004272f
C10453 FILLER_0_11_282/a_36_472# vss 0.007114f
C10454 FILLER_0_20_107/a_36_472# _098_ 0.011046f
C10455 FILLER_0_24_130/a_124_375# output24/a_224_472# 0.00515f
C10456 _411_/a_1204_472# _000_ 0.002575f
C10457 _136_ _097_ 0.002577f
C10458 FILLER_0_17_38/a_572_375# _179_ 0.002825f
C10459 _430_/a_448_472# net36 0.011598f
C10460 FILLER_0_14_81/a_36_472# _394_/a_728_93# 0.005826f
C10461 _018_ net22 0.141743f
C10462 _133_ _134_ 0.015205f
C10463 _186_ net17 0.001172f
C10464 vdd FILLER_0_10_94/a_124_375# 0.020076f
C10465 _417_/a_2560_156# _006_ 0.007804f
C10466 net35 vss 0.434438f
C10467 _299_/a_36_472# vdd 0.098451f
C10468 _140_ FILLER_0_21_150/a_124_375# 0.019084f
C10469 _057_ _069_ 0.053765f
C10470 _320_/a_224_472# _113_ 0.00871f
C10471 net56 FILLER_0_17_142/a_36_472# 0.003603f
C10472 FILLER_0_8_127/a_36_472# _119_ 0.053962f
C10473 _137_ _043_ 0.007284f
C10474 _119_ FILLER_0_8_156/a_572_375# 0.01739f
C10475 _431_/a_2665_112# net36 0.001523f
C10476 _363_/a_244_472# vdd 0.002075f
C10477 _449_/a_448_472# net72 0.01383f
C10478 _025_ _436_/a_448_472# 0.044246f
C10479 trimb[4] net38 0.124219f
C10480 net75 FILLER_0_0_232/a_124_375# 0.00217f
C10481 _079_ _253_/a_36_68# 0.002433f
C10482 _316_/a_1084_68# vdd 0.001166f
C10483 net79 _416_/a_2560_156# 0.013576f
C10484 _093_ FILLER_0_17_218/a_36_472# 0.006994f
C10485 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_484_472# 0.013276f
C10486 net55 FILLER_0_18_76/a_484_472# 0.003745f
C10487 _444_/a_36_151# vdd 0.071209f
C10488 FILLER_0_7_195/a_124_375# _062_ 0.001983f
C10489 FILLER_0_4_197/a_124_375# _002_ 0.001406f
C10490 output14/a_224_472# vss 0.012129f
C10491 cal_count\[3\] _408_/a_56_524# 0.001685f
C10492 output44/a_224_472# vss 0.014054f
C10493 output31/a_224_472# _418_/a_2665_112# 0.008243f
C10494 _136_ mask\[2\] 1.822289f
C10495 _053_ net67 0.672744f
C10496 _193_/a_36_160# _044_ 0.025719f
C10497 _415_/a_2665_112# net18 0.004988f
C10498 _077_ _070_ 0.29321f
C10499 output20/a_224_472# _109_ 0.003452f
C10500 _390_/a_36_68# net14 0.010844f
C10501 _198_/a_67_603# _099_ 0.0109f
C10502 _453_/a_1000_472# _042_ 0.004985f
C10503 _306_/a_36_68# _071_ 0.054312f
C10504 _058_ FILLER_0_10_94/a_484_472# 0.002096f
C10505 _311_/a_1212_473# _117_ 0.001673f
C10506 FILLER_0_20_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001543f
C10507 output44/a_224_472# FILLER_0_20_15/a_932_472# 0.0323f
C10508 _448_/a_448_472# net76 0.003937f
C10509 FILLER_0_2_93/a_124_375# vdd 0.008901f
C10510 vss _167_ 0.043544f
C10511 _080_ vdd 0.123811f
C10512 _118_ _331_/a_448_472# 0.001166f
C10513 FILLER_0_19_171/a_36_472# vdd 0.004762f
C10514 FILLER_0_19_171/a_1468_375# vss 0.054352f
C10515 FILLER_0_22_86/a_1380_472# net71 0.011277f
C10516 net73 fanout73/a_36_113# 0.02062f
C10517 mask\[8\] _437_/a_36_151# 0.005179f
C10518 FILLER_0_18_139/a_1468_375# _137_ 0.004111f
C10519 net16 _013_ 0.060401f
C10520 _114_ _113_ 0.201729f
C10521 trimb[1] FILLER_0_18_2/a_572_375# 0.010125f
C10522 net20 _098_ 0.087341f
C10523 _036_ FILLER_0_3_78/a_124_375# 0.00215f
C10524 _088_ FILLER_0_4_213/a_484_472# 0.018066f
C10525 cal_count\[3\] _314_/a_224_472# 0.002143f
C10526 net60 net30 0.001168f
C10527 _452_/a_3129_107# vdd 0.016611f
C10528 input5/a_36_113# clk 0.01086f
C10529 net72 FILLER_0_21_28/a_1380_472# 0.048287f
C10530 _058_ _122_ 0.040376f
C10531 _235_/a_67_603# vss 0.002019f
C10532 net47 FILLER_0_5_148/a_124_375# 0.008947f
C10533 net1 net5 0.266194f
C10534 mask\[0\] net79 0.243338f
C10535 _253_/a_36_68# cal_itt\[1\] 0.039692f
C10536 FILLER_0_6_177/a_484_472# FILLER_0_5_181/a_36_472# 0.05841f
C10537 _093_ _199_/a_36_160# 0.05226f
C10538 _359_/a_36_488# _129_ 0.002527f
C10539 FILLER_0_23_44/a_572_375# vdd -0.011314f
C10540 FILLER_0_10_214/a_36_472# _246_/a_36_68# 0.001844f
C10541 _058_ _227_/a_36_160# 0.008511f
C10542 trim_mask\[2\] _168_ 0.00704f
C10543 FILLER_0_7_59/a_124_375# FILLER_0_6_47/a_1468_375# 0.05841f
C10544 _132_ _354_/a_49_472# 0.034372f
C10545 net22 vss 1.28233f
C10546 _018_ vdd 0.048119f
C10547 _440_/a_1000_472# net47 0.011283f
C10548 _415_/a_36_151# _416_/a_1308_423# 0.00119f
C10549 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_572_375# 0.086635f
C10550 output22/a_224_472# _435_/a_1308_423# 0.005111f
C10551 net19 calibrate 0.043159f
C10552 FILLER_0_14_107/a_1468_375# vss 0.055167f
C10553 FILLER_0_14_107/a_36_472# vdd 0.114495f
C10554 FILLER_0_9_72/a_1380_472# vss 0.007254f
C10555 _136_ FILLER_0_16_115/a_124_375# 0.006372f
C10556 _448_/a_36_151# FILLER_0_2_177/a_572_375# 0.001597f
C10557 _414_/a_2665_112# _068_ 0.002324f
C10558 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_36_472# 0.086742f
C10559 FILLER_0_22_177/a_572_375# net33 0.013337f
C10560 _433_/a_36_151# _022_ 0.017789f
C10561 cal_itt\[3\] _375_/a_36_68# 0.005168f
C10562 result[4] net61 0.023257f
C10563 FILLER_0_10_256/a_124_375# net19 0.002884f
C10564 _395_/a_36_488# _071_ 0.00276f
C10565 FILLER_0_17_72/a_1468_375# _150_ 0.001076f
C10566 _010_ _419_/a_796_472# 0.001613f
C10567 _445_/a_36_151# net17 0.009838f
C10568 _091_ FILLER_0_20_169/a_36_472# 0.007537f
C10569 _437_/a_2665_112# FILLER_0_22_107/a_572_375# 0.001597f
C10570 FILLER_0_21_28/a_36_472# net17 0.00347f
C10571 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_124_375# 0.003732f
C10572 _306_/a_36_68# _095_ 0.001366f
C10573 FILLER_0_4_177/a_124_375# _087_ 0.002288f
C10574 _075_ net22 0.180274f
C10575 _069_ _310_/a_49_472# 0.023925f
C10576 FILLER_0_10_78/a_36_472# _453_/a_2665_112# 0.007491f
C10577 _430_/a_2248_156# mask\[1\] 0.001498f
C10578 net50 fanout49/a_36_160# 0.059373f
C10579 net34 net32 0.330134f
C10580 net50 FILLER_0_7_59/a_124_375# 0.002292f
C10581 _071_ FILLER_0_13_142/a_1468_375# 0.007453f
C10582 ctln[3] _411_/a_36_151# 0.004014f
C10583 _308_/a_124_24# FILLER_0_9_72/a_1380_472# 0.003595f
C10584 _402_/a_728_93# cal_count\[1\] 0.057043f
C10585 net54 FILLER_0_22_86/a_932_472# 0.047897f
C10586 net79 _099_ 0.010543f
C10587 _136_ FILLER_0_16_154/a_484_472# 0.007583f
C10588 net53 mask\[2\] 0.005907f
C10589 net3 FILLER_0_15_2/a_484_472# 0.002224f
C10590 _428_/a_1308_423# _131_ 0.037599f
C10591 net48 _316_/a_124_24# 0.068708f
C10592 fanout66/a_36_113# net66 0.032757f
C10593 net52 _170_ 0.378738f
C10594 net20 _070_ 0.075448f
C10595 net60 _417_/a_36_151# 0.007446f
C10596 _432_/a_2248_156# _093_ 0.012955f
C10597 trim[2] output41/a_224_472# 0.005452f
C10598 output40/a_224_472# trim[3] 0.122003f
C10599 mask\[8\] _051_ 0.003475f
C10600 _059_ _163_ 0.038651f
C10601 result[0] net5 0.001104f
C10602 _087_ _088_ 0.001219f
C10603 vss _433_/a_2665_112# 0.035903f
C10604 mask\[0\] _429_/a_2560_156# 0.010913f
C10605 net16 FILLER_0_6_37/a_124_375# 0.010358f
C10606 cal_count\[3\] FILLER_0_11_78/a_124_375# 0.019818f
C10607 _402_/a_56_567# net40 0.033835f
C10608 FILLER_0_3_172/a_3260_375# net22 0.015274f
C10609 _086_ FILLER_0_4_177/a_124_375# 0.024433f
C10610 _094_ _418_/a_2248_156# 0.028557f
C10611 FILLER_0_7_72/a_1916_375# _376_/a_36_160# 0.001925f
C10612 _086_ net57 0.126563f
C10613 _105_ _204_/a_67_603# 0.061486f
C10614 FILLER_0_9_28/a_932_472# FILLER_0_10_37/a_36_472# 0.026657f
C10615 _057_ _267_/a_1792_472# 0.003005f
C10616 _422_/a_448_472# mask\[7\] 0.048658f
C10617 result[6] _420_/a_448_472# 0.017262f
C10618 FILLER_0_16_57/a_1380_472# _131_ 0.008223f
C10619 net44 _221_/a_36_160# 0.013363f
C10620 net34 FILLER_0_22_177/a_932_472# 0.003953f
C10621 _054_ vdd 0.360345f
C10622 FILLER_0_9_60/a_36_472# net51 0.059421f
C10623 _091_ FILLER_0_17_218/a_124_375# 0.013726f
C10624 FILLER_0_6_177/a_124_375# net47 0.002925f
C10625 _116_ _085_ 0.049304f
C10626 fanout77/a_36_113# _103_ 0.006045f
C10627 _410_/a_36_68# _188_ 0.007731f
C10628 _115_ FILLER_0_10_94/a_484_472# 0.015061f
C10629 _415_/a_1308_423# _004_ 0.002098f
C10630 _321_/a_2590_472# _176_ 0.001932f
C10631 _069_ _395_/a_1044_488# 0.002244f
C10632 _445_/a_1204_472# net40 0.003916f
C10633 _053_ FILLER_0_6_47/a_1916_375# 0.008103f
C10634 _093_ FILLER_0_17_72/a_932_472# 0.004367f
C10635 _126_ _120_ 0.055349f
C10636 _126_ _038_ 0.031198f
C10637 _008_ _418_/a_2665_112# 0.010862f
C10638 FILLER_0_15_235/a_572_375# vss 0.002683f
C10639 FILLER_0_15_235/a_36_472# vdd 0.019127f
C10640 FILLER_0_9_28/a_1380_472# vdd 0.01306f
C10641 vdd _278_/a_36_160# 0.016488f
C10642 FILLER_0_9_105/a_36_472# vss 0.002744f
C10643 FILLER_0_9_105/a_484_472# vdd 0.03152f
C10644 FILLER_0_13_142/a_484_472# _043_ 0.011974f
C10645 _104_ vdd 0.662413f
C10646 FILLER_0_20_177/a_484_472# vss 0.001256f
C10647 FILLER_0_20_177/a_932_472# vdd 0.035019f
C10648 vdd vss 15.42941f
C10649 fanout66/a_36_113# FILLER_0_3_54/a_124_375# 0.002853f
C10650 FILLER_0_2_101/a_124_375# _160_ 0.001047f
C10651 _192_/a_67_603# vss 0.007021f
C10652 net16 _447_/a_1204_472# 0.00194f
C10653 output16/a_224_472# _447_/a_2665_112# 0.005471f
C10654 _178_ vdd 0.440802f
C10655 _408_/a_1336_472# _186_ 0.010089f
C10656 net36 FILLER_0_15_212/a_1468_375# 0.005276f
C10657 _115_ _122_ 0.004082f
C10658 FILLER_0_24_63/a_36_472# ctlp[9] 0.012298f
C10659 input2/a_36_113# input5/a_36_113# 0.01088f
C10660 _276_/a_36_160# FILLER_0_18_209/a_484_472# 0.003913f
C10661 _013_ _041_ 0.00271f
C10662 FILLER_0_17_56/a_124_375# _183_ 0.019253f
C10663 FILLER_0_2_165/a_36_472# net22 0.028367f
C10664 FILLER_0_20_98/a_124_375# net14 0.05242f
C10665 FILLER_0_20_15/a_932_472# vdd 0.002617f
C10666 _079_ cal_itt\[1\] 0.012324f
C10667 FILLER_0_9_28/a_124_375# net40 0.047331f
C10668 cal_count\[3\] _117_ 0.00114f
C10669 mask\[7\] _108_ 0.785154f
C10670 FILLER_0_18_107/a_1020_375# vdd -0.008765f
C10671 FILLER_0_8_127/a_36_472# _129_ 0.060819f
C10672 _076_ FILLER_0_8_239/a_124_375# 0.007237f
C10673 _422_/a_1000_472# vdd 0.005284f
C10674 _063_ trim_val\[1\] 0.038045f
C10675 _115_ _227_/a_36_160# 0.00124f
C10676 mask\[7\] net19 0.003605f
C10677 net7 _239_/a_36_160# 0.068281f
C10678 cal_count\[2\] _452_/a_2225_156# 0.003086f
C10679 _062_ _060_ 0.032472f
C10680 FILLER_0_18_139/a_124_375# _145_ 0.00346f
C10681 _075_ vdd 0.190898f
C10682 net79 FILLER_0_12_220/a_1020_375# 0.010818f
C10683 _441_/a_2248_156# vdd -0.003818f
C10684 _441_/a_1204_472# vss 0.011996f
C10685 FILLER_0_3_221/a_124_375# FILLER_0_3_212/a_124_375# 0.002036f
C10686 _232_/a_255_603# _164_ 0.001274f
C10687 _430_/a_1308_423# vss 0.003054f
C10688 _031_ _158_ 0.015116f
C10689 mask\[4\] FILLER_0_18_177/a_572_375# 0.015941f
C10690 trim_val\[4\] _386_/a_124_24# 0.001172f
C10691 _430_/a_36_151# net36 0.003701f
C10692 _308_/a_124_24# vdd 0.011014f
C10693 _447_/a_448_472# net68 0.012962f
C10694 output36/a_224_472# result[2] 0.002356f
C10695 _165_ FILLER_0_6_47/a_36_472# 0.077573f
C10696 _106_ net33 0.001049f
C10697 _413_/a_36_151# net82 0.00601f
C10698 FILLER_0_19_125/a_36_472# vdd 0.003414f
C10699 FILLER_0_8_239/a_36_472# _317_/a_36_113# 0.00191f
C10700 _308_/a_1152_472# trim_mask\[0\] 0.004076f
C10701 FILLER_0_19_47/a_124_375# net26 0.008432f
C10702 _039_ cal_count\[0\] 0.219667f
C10703 _131_ FILLER_0_17_104/a_1468_375# 0.006022f
C10704 ctlp[1] _421_/a_2560_156# 0.001062f
C10705 fanout71/a_36_113# net71 0.087994f
C10706 vdd _107_ 0.038236f
C10707 FILLER_0_21_28/a_1916_375# _423_/a_36_151# 0.001597f
C10708 net69 _030_ 0.49547f
C10709 net15 _423_/a_1308_423# 0.001999f
C10710 _226_/a_1044_68# net21 0.001903f
C10711 FILLER_0_19_55/a_124_375# _013_ 0.009611f
C10712 _328_/a_36_113# _070_ 0.016264f
C10713 _442_/a_1308_423# FILLER_0_2_111/a_1468_375# 0.001048f
C10714 _449_/a_1308_423# _038_ 0.021006f
C10715 FILLER_0_3_172/a_3260_375# vdd -0.013516f
C10716 _359_/a_1492_488# _133_ 0.003815f
C10717 _308_/a_848_380# trim_mask\[0\] 0.035693f
C10718 FILLER_0_5_54/a_1468_375# _440_/a_36_151# 0.059049f
C10719 net50 net17 0.010654f
C10720 FILLER_0_15_290/a_36_472# net18 0.002452f
C10721 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_36_472# 0.086635f
C10722 result[7] _420_/a_448_472# 0.003274f
C10723 FILLER_0_15_290/a_124_375# result[3] 0.020277f
C10724 net20 net82 0.026007f
C10725 FILLER_0_11_101/a_36_472# net14 0.04522f
C10726 _189_/a_67_603# net27 0.008028f
C10727 _257_/a_36_472# _122_ 0.007741f
C10728 _132_ _131_ 0.444097f
C10729 net50 trim_val\[1\] 0.002079f
C10730 FILLER_0_7_104/a_572_375# _058_ 0.006125f
C10731 _127_ _428_/a_36_151# 0.030717f
C10732 output42/a_224_472# _236_/a_36_160# 0.001892f
C10733 FILLER_0_19_125/a_124_375# _022_ 0.055527f
C10734 _052_ FILLER_0_18_37/a_572_375# 0.00706f
C10735 FILLER_0_18_2/a_2724_472# _452_/a_36_151# 0.011733f
C10736 _251_/a_1130_472# vss 0.001211f
C10737 _267_/a_36_472# _113_ 0.014178f
C10738 FILLER_0_10_28/a_124_375# output6/a_224_472# 0.002633f
C10739 net9 vss 0.086497f
C10740 _147_ net33 0.001686f
C10741 fanout76/a_36_160# vdd 0.108854f
C10742 net7 net41 0.243942f
C10743 net15 FILLER_0_17_72/a_932_472# 0.001122f
C10744 output17/a_224_472# vss 0.009426f
C10745 FILLER_0_18_76/a_124_375# net71 0.008427f
C10746 net70 net74 0.017928f
C10747 _274_/a_716_497# net20 0.001321f
C10748 vdd _416_/a_2248_156# 0.004325f
C10749 _044_ _416_/a_36_151# 0.032206f
C10750 _422_/a_2248_156# _108_ 0.019477f
C10751 _412_/a_36_151# net81 0.014094f
C10752 _135_ vss 0.097337f
C10753 _126_ state\[2\] 0.030985f
C10754 FILLER_0_5_88/a_124_375# vdd 0.020896f
C10755 _091_ _060_ 0.085764f
C10756 _422_/a_2248_156# net19 0.003451f
C10757 FILLER_0_10_214/a_124_375# _247_/a_36_160# 0.005732f
C10758 FILLER_0_11_142/a_36_472# cal_count\[3\] 0.008454f
C10759 FILLER_0_22_177/a_1020_375# mask\[6\] 0.002657f
C10760 _098_ _434_/a_2560_156# 0.003888f
C10761 net35 FILLER_0_22_177/a_572_375# 0.007797f
C10762 _195_/a_67_603# vdd 0.022493f
C10763 net80 FILLER_0_17_161/a_124_375# 0.021914f
C10764 _258_/a_36_160# _073_ 0.079254f
C10765 net75 net48 0.10167f
C10766 _010_ net77 0.009534f
C10767 _430_/a_2665_112# vss 0.031646f
C10768 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3260_375# 0.086635f
C10769 _021_ _097_ 0.002219f
C10770 FILLER_0_5_128/a_484_472# FILLER_0_5_136/a_36_472# 0.013276f
C10771 _176_ FILLER_0_11_78/a_572_375# 0.013887f
C10772 _238_/a_67_603# net50 0.002229f
C10773 _365_/a_244_472# net14 0.001257f
C10774 _056_ _246_/a_36_68# 0.017953f
C10775 fanout81/a_36_160# net58 0.013959f
C10776 _289_/a_36_472# _099_ 0.035055f
C10777 FILLER_0_2_165/a_124_375# vss 0.008386f
C10778 FILLER_0_2_165/a_36_472# vdd -0.003333f
C10779 net16 _064_ 0.121797f
C10780 FILLER_0_4_49/a_572_375# net49 0.004345f
C10781 net75 FILLER_0_8_247/a_1020_375# 0.009573f
C10782 fanout54/a_36_160# FILLER_0_18_139/a_1020_375# 0.031033f
C10783 _140_ FILLER_0_22_128/a_36_472# 0.050084f
C10784 _118_ _062_ 0.029651f
C10785 result[1] FILLER_0_11_282/a_124_375# 0.018322f
C10786 _411_/a_1204_472# ctln[1] 0.031348f
C10787 fanout67/a_36_160# vss 0.005344f
C10788 output34/a_224_472# _293_/a_36_472# 0.001888f
C10789 _431_/a_2248_156# FILLER_0_15_142/a_572_375# 0.001374f
C10790 result[7] _419_/a_1308_423# 0.015718f
C10791 FILLER_0_4_197/a_1020_375# _088_ 0.013641f
C10792 _148_ FILLER_0_22_107/a_572_375# 0.00652f
C10793 _036_ _167_ 0.003223f
C10794 trim_mask\[1\] FILLER_0_6_90/a_36_472# 0.001162f
C10795 _072_ net23 0.006278f
C10796 ctln[7] FILLER_0_0_130/a_36_472# 0.012298f
C10797 FILLER_0_2_177/a_36_472# net22 0.002517f
C10798 result[9] net61 0.014374f
C10799 FILLER_0_9_28/a_1916_375# _054_ 0.005889f
C10800 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_124_375# 0.012001f
C10801 net15 _447_/a_2560_156# 0.001586f
C10802 _323_/a_36_113# FILLER_0_10_247/a_36_472# 0.00136f
C10803 FILLER_0_14_107/a_484_472# _043_ 0.001641f
C10804 _069_ _018_ 0.002777f
C10805 net44 cal_count\[2\] 0.191151f
C10806 result[2] FILLER_0_14_263/a_36_472# 0.001134f
C10807 _184_ vdd 0.202732f
C10808 _235_/a_67_603# _036_ 0.043345f
C10809 net69 trim_mask\[3\] 0.017779f
C10810 _183_ FILLER_0_18_53/a_124_375# 0.001032f
C10811 _401_/a_36_68# vdd 0.003745f
C10812 FILLER_0_5_128/a_124_375# net47 0.011156f
C10813 _279_/a_652_68# vdd 0.001562f
C10814 fanout61/a_36_113# net18 0.001668f
C10815 _374_/a_36_68# FILLER_0_8_156/a_484_472# 0.002559f
C10816 _068_ _246_/a_36_68# 0.059106f
C10817 fanout81/a_36_160# net82 0.027351f
C10818 _420_/a_1308_423# vss 0.001461f
C10819 output34/a_224_472# net19 0.001308f
C10820 _013_ _424_/a_1308_423# 0.007751f
C10821 _095_ FILLER_0_14_107/a_1468_375# 0.010523f
C10822 net16 _042_ 0.012486f
C10823 _141_ FILLER_0_19_155/a_572_375# 0.033271f
C10824 _359_/a_36_488# _152_ 0.032195f
C10825 FILLER_0_8_138/a_36_472# vdd 0.008749f
C10826 net44 input3/a_36_113# 0.016865f
C10827 FILLER_0_19_47/a_484_472# _052_ 0.01589f
C10828 FILLER_0_4_49/a_484_472# FILLER_0_3_54/a_36_472# 0.026657f
C10829 FILLER_0_16_89/a_1468_375# FILLER_0_17_72/a_3260_375# 0.026339f
C10830 FILLER_0_16_89/a_484_472# FILLER_0_17_72/a_2364_375# 0.001723f
C10831 FILLER_0_12_220/a_36_472# _248_/a_36_68# 0.006596f
C10832 FILLER_0_7_72/a_3172_472# FILLER_0_7_104/a_36_472# 0.013276f
C10833 mask\[5\] _144_ 0.38642f
C10834 _177_ _451_/a_2225_156# 0.031347f
C10835 _444_/a_448_472# net67 0.046278f
C10836 net73 net36 0.073334f
C10837 net72 _394_/a_244_524# 0.001083f
C10838 net52 _443_/a_448_472# 0.050192f
C10839 net47 _365_/a_36_68# 0.020511f
C10840 valid _425_/a_2665_112# 0.001839f
C10841 FILLER_0_10_78/a_572_375# FILLER_0_9_72/a_1380_472# 0.001543f
C10842 trim_mask\[0\] net14 0.499565f
C10843 net44 _450_/a_448_472# 0.050752f
C10844 ctln[0] net7 0.001209f
C10845 _446_/a_2665_112# net66 0.00195f
C10846 vdd _450_/a_1040_527# 0.005529f
C10847 _071_ vdd 0.074299f
C10848 mask\[8\] _436_/a_36_151# 0.032521f
C10849 FILLER_0_16_241/a_36_472# net30 0.001025f
C10850 _189_/a_67_603# FILLER_0_14_235/a_36_472# 0.002778f
C10851 _091_ _093_ 0.035503f
C10852 _322_/a_848_380# _070_ 0.006182f
C10853 _423_/a_2560_156# vss 0.002241f
C10854 net4 FILLER_0_4_213/a_572_375# 0.001015f
C10855 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001597f
C10856 output48/a_224_472# net19 0.054227f
C10857 _077_ FILLER_0_10_94/a_36_472# 0.001114f
C10858 net69 net13 0.005834f
C10859 net34 _421_/a_2665_112# 0.001056f
C10860 net63 FILLER_0_20_177/a_932_472# 0.004375f
C10861 _104_ net63 0.005363f
C10862 cal_count\[3\] _172_ 0.03048f
C10863 _316_/a_124_24# net37 0.011141f
C10864 _076_ FILLER_0_8_156/a_36_472# 0.006989f
C10865 _068_ FILLER_0_8_156/a_572_375# 0.00185f
C10866 FILLER_0_20_193/a_36_472# _098_ 0.006652f
C10867 net20 ctlp[2] 0.254928f
C10868 FILLER_0_20_177/a_572_375# _434_/a_36_151# 0.059049f
C10869 FILLER_0_16_154/a_1020_375# vdd 0.004279f
C10870 FILLER_0_16_154/a_572_375# vss 0.003976f
C10871 net63 vss 0.566021f
C10872 _323_/a_36_113# _128_ 0.014377f
C10873 _028_ FILLER_0_7_72/a_3172_472# 0.001873f
C10874 _027_ vdd 0.146607f
C10875 FILLER_0_4_49/a_484_472# _164_ 0.003258f
C10876 _421_/a_448_472# _010_ 0.039422f
C10877 _181_ _402_/a_1948_68# 0.001223f
C10878 FILLER_0_15_142/a_484_472# _427_/a_36_151# 0.001723f
C10879 net22 _435_/a_2560_156# 0.002281f
C10880 FILLER_0_5_198/a_572_375# vss 0.055087f
C10881 FILLER_0_5_198/a_36_472# vdd 0.088893f
C10882 _077_ calibrate 0.055446f
C10883 net31 result[6] 0.002094f
C10884 net34 output33/a_224_472# 0.077682f
C10885 FILLER_0_22_86/a_36_472# net14 0.003007f
C10886 _415_/a_796_472# net27 0.004502f
C10887 _144_ _433_/a_448_472# 0.075144f
C10888 output11/a_224_472# output8/a_224_472# 0.003437f
C10889 FILLER_0_5_128/a_124_375# net74 0.013683f
C10890 _419_/a_1000_472# vdd 0.004107f
C10891 _119_ _324_/a_224_472# 0.00368f
C10892 output45/a_224_472# trimb[3] 0.076387f
C10893 FILLER_0_16_89/a_1380_472# _040_ 0.008446f
C10894 _086_ FILLER_0_6_177/a_572_375# 0.012909f
C10895 FILLER_0_2_177/a_572_375# vss 0.008507f
C10896 FILLER_0_2_177/a_36_472# vdd 0.110255f
C10897 net17 _039_ 0.079171f
C10898 FILLER_0_16_89/a_1020_375# _093_ 0.004133f
C10899 net19 _420_/a_1204_472# 0.001828f
C10900 _077_ net21 0.032627f
C10901 _076_ _269_/a_36_472# 0.001618f
C10902 _078_ _083_ 0.01015f
C10903 state\[2\] state\[1\] 0.229832f
C10904 net15 ctln[8] 0.205163f
C10905 result[8] _011_ 0.001294f
C10906 net52 _029_ 0.03261f
C10907 _432_/a_1204_472# _137_ 0.006554f
C10908 _069_ vss 0.323941f
C10909 _093_ FILLER_0_17_142/a_124_375# 0.009328f
C10910 _096_ _335_/a_49_472# 0.00151f
C10911 FILLER_0_13_212/a_572_375# net79 0.009626f
C10912 net62 FILLER_0_13_212/a_1020_375# 0.001597f
C10913 _095_ vdd 1.051346f
C10914 _035_ _034_ 1.26804f
C10915 net49 _029_ 0.004408f
C10916 _430_/a_36_151# FILLER_0_18_177/a_2724_472# 0.001512f
C10917 _158_ _157_ 0.001663f
C10918 net4 FILLER_0_3_221/a_1020_375# 0.006974f
C10919 mask\[7\] _435_/a_1204_472# 0.007888f
C10920 ctln[1] _411_/a_2560_156# 0.001413f
C10921 _394_/a_718_524# cal_count\[1\] 0.009499f
C10922 net10 net75 0.073869f
C10923 _450_/a_36_151# output6/a_224_472# 0.134892f
C10924 _261_/a_36_160# net47 0.010976f
C10925 _036_ vdd 0.364747f
C10926 net57 _061_ 0.127011f
C10927 _091_ _337_/a_49_472# 0.014992f
C10928 FILLER_0_10_78/a_572_375# vdd -0.014642f
C10929 FILLER_0_7_195/a_36_472# _074_ 0.008706f
C10930 _077_ _410_/a_36_68# 0.020334f
C10931 output26/a_224_472# vdd 0.047141f
C10932 FILLER_0_5_128/a_124_375# _159_ 0.003644f
C10933 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_124_375# 0.001597f
C10934 net57 _311_/a_66_473# 0.013777f
C10935 FILLER_0_12_220/a_124_375# vdd -0.008946f
C10936 _053_ _078_ 0.137388f
C10937 net23 FILLER_0_22_128/a_3172_472# 0.015058f
C10938 FILLER_0_18_139/a_484_472# vdd 0.003106f
C10939 FILLER_0_18_139/a_36_472# vss 0.007877f
C10940 FILLER_0_4_123/a_124_375# _370_/a_124_24# 0.007188f
C10941 FILLER_0_16_73/a_572_375# net15 0.002076f
C10942 _165_ _220_/a_67_603# 0.004199f
C10943 FILLER_0_9_72/a_932_472# _439_/a_36_151# 0.001723f
C10944 FILLER_0_7_72/a_2812_375# _077_ 0.002969f
C10945 FILLER_0_15_282/a_36_472# net18 0.036858f
C10946 _093_ FILLER_0_18_107/a_932_472# 0.008683f
C10947 fanout65/a_36_113# net5 0.027955f
C10948 _126_ _125_ 0.032402f
C10949 FILLER_0_22_177/a_124_375# vss 0.002674f
C10950 FILLER_0_22_177/a_572_375# vdd -0.003694f
C10951 FILLER_0_18_107/a_484_472# mask\[9\] 0.001955f
C10952 FILLER_0_15_282/a_572_375# result[3] 0.038939f
C10953 net19 _419_/a_2248_156# 0.012726f
C10954 _093_ _110_ 0.08348f
C10955 _086_ FILLER_0_10_107/a_572_375# 0.001179f
C10956 _390_/a_692_472# _136_ 0.004782f
C10957 _050_ net23 0.003752f
C10958 trim_val\[3\] _441_/a_1308_423# 0.001312f
C10959 _426_/a_1308_423# net64 0.021119f
C10960 FILLER_0_4_107/a_124_375# _160_ 0.005906f
C10961 _255_/a_224_552# _374_/a_36_68# 0.00191f
C10962 mask\[3\] _141_ 0.361692f
C10963 net32 _295_/a_36_472# 0.002637f
C10964 net31 result[7] 0.231528f
C10965 net71 _437_/a_2560_156# 0.037081f
C10966 _413_/a_36_151# net21 0.012223f
C10967 _081_ _265_/a_468_472# 0.005156f
C10968 _435_/a_2560_156# vdd 0.001372f
C10969 _435_/a_2665_112# vss 0.002665f
C10970 mask\[3\] net36 0.002974f
C10971 result[0] result[1] 0.06045f
C10972 net20 calibrate 0.044792f
C10973 _449_/a_448_472# vdd 0.007757f
C10974 _449_/a_36_151# vss 0.014774f
C10975 net57 _072_ 0.108982f
C10976 _154_ _365_/a_36_68# 0.02267f
C10977 result[6] _421_/a_36_151# 0.032036f
C10978 net25 _214_/a_36_160# 0.019894f
C10979 _265_/a_244_68# _082_ 0.031951f
C10980 _443_/a_1308_423# net13 0.004098f
C10981 _443_/a_1000_472# net23 0.034596f
C10982 net72 net55 0.233515f
C10983 net28 vss 0.185012f
C10984 net28 _192_/a_255_603# 0.003166f
C10985 FILLER_0_9_223/a_572_375# vss 0.00704f
C10986 _026_ _437_/a_36_151# 0.012193f
C10987 _149_ _437_/a_1308_423# 0.015677f
C10988 vdd output41/a_224_472# 0.003282f
C10989 net44 net67 0.08001f
C10990 _053_ FILLER_0_5_54/a_932_472# 0.001578f
C10991 _086_ _128_ 0.085571f
C10992 _122_ FILLER_0_6_231/a_124_375# 0.013183f
C10993 _346_/a_49_472# vdd -0.002208f
C10994 trim_val\[4\] _443_/a_2560_156# 0.049334f
C10995 _448_/a_2560_156# trim_mask\[4\] 0.001306f
C10996 net39 trim[1] 0.115976f
C10997 net21 FILLER_0_12_196/a_36_472# 0.001298f
C10998 FILLER_0_17_200/a_124_375# FILLER_0_18_177/a_2724_472# 0.001597f
C10999 FILLER_0_14_263/a_124_375# output30/a_224_472# 0.011584f
C11000 _164_ FILLER_0_6_37/a_36_472# 0.001049f
C11001 _431_/a_36_151# _142_ 0.030496f
C11002 _402_/a_1296_93# vdd 0.017239f
C11003 _016_ _428_/a_2248_156# 0.048889f
C11004 net41 FILLER_0_17_38/a_36_472# 0.001308f
C11005 net20 output8/a_224_472# 0.084627f
C11006 FILLER_0_16_73/a_124_375# _131_ 0.015859f
C11007 _083_ _263_/a_224_472# 0.003191f
C11008 _020_ FILLER_0_18_107/a_2364_375# 0.003755f
C11009 net29 _006_ 0.135646f
C11010 FILLER_0_21_133/a_36_472# vss 0.004298f
C11011 net75 net37 0.07785f
C11012 net50 FILLER_0_8_24/a_572_375# 0.001597f
C11013 mask\[4\] FILLER_0_19_171/a_124_375# 0.001988f
C11014 FILLER_0_12_236/a_36_472# vdd 0.086431f
C11015 FILLER_0_12_236/a_572_375# vss 0.025768f
C11016 trim[0] _064_ 0.014422f
C11017 output37/a_224_472# vdd 0.082206f
C11018 FILLER_0_14_91/a_36_472# vdd 0.08739f
C11019 FILLER_0_14_91/a_572_375# vss 0.054783f
C11020 FILLER_0_15_282/a_484_472# _417_/a_36_151# 0.059367f
C11021 FILLER_0_15_282/a_36_472# _417_/a_448_472# 0.011962f
C11022 fanout82/a_36_113# _316_/a_848_380# 0.001292f
C11023 net52 _163_ 0.00157f
C11024 _385_/a_36_68# vdd 0.01625f
C11025 _442_/a_1308_423# _031_ 0.003679f
C11026 FILLER_0_21_28/a_1380_472# vdd 0.007073f
C11027 net72 net17 0.004503f
C11028 net50 FILLER_0_2_93/a_36_472# 0.008147f
C11029 ctlp[2] _009_ 0.220631f
C11030 output47/a_224_472# FILLER_0_18_2/a_484_472# 0.00175f
C11031 _423_/a_1308_423# _012_ 0.01389f
C11032 FILLER_0_1_192/a_124_375# net21 0.067765f
C11033 FILLER_0_13_100/a_124_375# _043_ 0.010818f
C11034 net36 _438_/a_36_151# 0.076525f
C11035 _093_ net14 0.11038f
C11036 output15/a_224_472# net52 0.007862f
C11037 net15 fanout50/a_36_160# 0.029852f
C11038 _001_ cal_itt\[0\] 0.004843f
C11039 _429_/a_36_151# net79 0.02414f
C11040 net52 FILLER_0_11_78/a_124_375# 0.006273f
C11041 FILLER_0_10_78/a_1020_375# _389_/a_36_148# 0.001335f
C11042 mask\[4\] FILLER_0_17_200/a_484_472# 0.001701f
C11043 net62 _429_/a_448_472# 0.002713f
C11044 _161_ FILLER_0_6_177/a_484_472# 0.001723f
C11045 net36 _451_/a_3129_107# 0.013154f
C11046 _077_ FILLER_0_10_78/a_36_472# 0.002486f
C11047 net15 _110_ 0.016359f
C11048 net54 _437_/a_2665_112# 0.061157f
C11049 _427_/a_1000_472# net23 0.003046f
C11050 net47 FILLER_0_5_136/a_124_375# 0.010674f
C11051 FILLER_0_21_28/a_1468_375# _424_/a_36_151# 0.059049f
C11052 net79 net18 0.222939f
C11053 net50 trim_mask\[2\] 0.267074f
C11054 net76 FILLER_0_5_198/a_484_472# 0.00169f
C11055 comp net44 0.079931f
C11056 output15/a_224_472# net49 0.005626f
C11057 FILLER_0_5_117/a_124_375# _086_ 0.003725f
C11058 _332_/a_36_472# vdd 0.017097f
C11059 net62 result[3] 0.451989f
C11060 FILLER_0_4_197/a_1468_375# net59 0.050218f
C11061 FILLER_0_14_50/a_36_472# cal_count\[1\] 0.030015f
C11062 _068_ _315_/a_36_68# 0.003516f
C11063 net64 FILLER_0_8_239/a_36_472# 0.002666f
C11064 net77 vss 0.327705f
C11065 output44/a_224_472# output46/a_224_472# 0.005749f
C11066 _096_ _136_ 0.022182f
C11067 FILLER_0_9_223/a_484_472# net20 0.002601f
C11068 net76 FILLER_0_2_177/a_484_472# 0.012872f
C11069 result[1] _416_/a_1000_472# 0.001529f
C11070 net28 _416_/a_2248_156# 0.001082f
C11071 FILLER_0_10_247/a_124_375# fanout79/a_36_160# 0.010334f
C11072 _274_/a_36_68# FILLER_0_12_220/a_484_472# 0.001048f
C11073 result[9] FILLER_0_23_274/a_36_472# 0.0064f
C11074 _002_ net65 0.042811f
C11075 FILLER_0_7_72/a_2812_375# net50 0.006598f
C11076 FILLER_0_16_57/a_1020_375# _176_ 0.006334f
C11077 FILLER_0_7_162/a_36_472# net37 0.090785f
C11078 net53 _451_/a_836_156# 0.006521f
C11079 _324_/a_224_472# _129_ 0.009728f
C11080 _106_ vdd 0.232973f
C11081 _131_ FILLER_0_17_56/a_36_472# 0.001491f
C11082 _130_ net53 0.00399f
C11083 _411_/a_2665_112# cal_itt\[0\] 0.010667f
C11084 output32/a_224_472# _418_/a_36_151# 0.07368f
C11085 net28 _195_/a_67_603# 0.012984f
C11086 output32/a_224_472# result[7] 0.063135f
C11087 mask\[5\] FILLER_0_19_187/a_484_472# 0.007596f
C11088 _089_ _003_ 0.014763f
C11089 result[4] net62 0.050684f
C11090 net20 _411_/a_448_472# 0.002167f
C11091 _370_/a_124_24# _081_ 0.015048f
C11092 net54 net14 0.121719f
C11093 trimb[4] FILLER_0_15_2/a_124_375# 0.003305f
C11094 _413_/a_448_472# net82 0.004927f
C11095 FILLER_0_21_125/a_124_375# net54 0.008377f
C11096 FILLER_0_10_78/a_932_472# vss 0.002987f
C11097 _132_ FILLER_0_15_116/a_484_472# 0.010148f
C11098 _182_ _180_ 0.090106f
C11099 FILLER_0_14_81/a_36_472# vss 0.007047f
C11100 net60 _418_/a_1308_423# 0.016365f
C11101 _119_ _058_ 0.692466f
C11102 net60 _006_ 0.006254f
C11103 output39/a_224_472# net49 0.039256f
C11104 output29/a_224_472# _044_ 0.087528f
C11105 _115_ FILLER_0_10_78/a_1020_375# 0.064761f
C11106 _011_ _109_ 0.055905f
C11107 _426_/a_2248_156# vdd 0.003943f
C11108 _028_ FILLER_0_6_90/a_484_472# 0.01566f
C11109 _439_/a_2665_112# trim_mask\[0\] 0.020363f
C11110 _147_ vdd 0.09215f
C11111 _098_ _438_/a_2665_112# 0.004321f
C11112 FILLER_0_9_290/a_36_472# vss 0.011755f
C11113 _431_/a_36_151# FILLER_0_14_123/a_124_375# 0.002807f
C11114 output38/a_224_472# trim[0] 0.026911f
C11115 _176_ FILLER_0_15_59/a_36_472# 0.00622f
C11116 net60 _103_ 0.066266f
C11117 _059_ net37 0.011845f
C11118 output27/a_224_472# FILLER_0_9_282/a_36_472# 0.001711f
C11119 net79 _417_/a_448_472# 0.028398f
C11120 _427_/a_1204_472# net74 0.003057f
C11121 FILLER_0_1_98/a_36_472# net52 0.005688f
C11122 net50 FILLER_0_4_91/a_124_375# 0.022557f
C11123 net55 FILLER_0_17_38/a_484_472# 0.013624f
C11124 net62 _417_/a_1308_423# 0.006676f
C11125 _326_/a_36_160# _058_ 0.003897f
C11126 FILLER_0_24_130/a_36_472# vdd 0.050082f
C11127 cal_itt\[3\] calibrate 1.141592f
C11128 _089_ net37 0.0326f
C11129 FILLER_0_14_107/a_36_472# _451_/a_36_151# 0.001723f
C11130 _335_/a_49_472# _138_ 0.005957f
C11131 output11/a_224_472# _413_/a_2665_112# 0.001492f
C11132 FILLER_0_6_47/a_2812_375# vdd 0.002455f
C11133 FILLER_0_6_47/a_2364_375# vss 0.008275f
C11134 _126_ _043_ 0.128227f
C11135 net18 FILLER_0_13_290/a_124_375# 0.007717f
C11136 _431_/a_2665_112# FILLER_0_17_142/a_572_375# 0.001092f
C11137 _068_ FILLER_0_5_148/a_484_472# 0.016952f
C11138 ctln[6] FILLER_0_0_130/a_124_375# 0.026786f
C11139 net20 mask\[1\] 0.09671f
C11140 FILLER_0_15_142/a_36_472# net74 0.003166f
C11141 net15 _164_ 0.026132f
C11142 net81 net1 0.03613f
C11143 cal_itt\[3\] net21 0.175781f
C11144 net63 FILLER_0_22_177/a_572_375# 0.001597f
C11145 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1380_472# 0.013277f
C11146 _285_/a_36_472# net36 0.003032f
C11147 cal_count\[2\] _402_/a_728_93# 0.036871f
C11148 FILLER_0_4_99/a_124_375# _156_ 0.081915f
C11149 _140_ vss 0.53195f
C11150 _282_/a_36_160# vss 0.005221f
C11151 _104_ _421_/a_448_472# 0.001106f
C11152 _414_/a_36_151# cal_itt\[3\] 0.049033f
C11153 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_484_472# 0.013276f
C11154 FILLER_0_6_90/a_572_375# net14 0.031929f
C11155 _050_ _436_/a_2248_156# 0.023725f
C11156 output35/a_224_472# net33 0.170613f
C11157 fanout71/a_36_113# FILLER_0_19_111/a_484_472# 0.007864f
C11158 net38 net66 0.040578f
C11159 net27 FILLER_0_9_282/a_484_472# 0.006955f
C11160 _395_/a_36_488# _070_ 0.005165f
C11161 FILLER_0_9_28/a_2364_375# _053_ 0.029866f
C11162 net35 _098_ 0.017288f
C11163 vss FILLER_0_6_231/a_484_472# 0.005629f
C11164 _421_/a_448_472# vss -0.001027f
C11165 _421_/a_1308_423# vdd 0.021664f
C11166 net38 _067_ 0.062447f
C11167 net63 _435_/a_2560_156# 0.023868f
C11168 _053_ FILLER_0_7_72/a_484_472# 0.00887f
C11169 _133_ _120_ 0.003762f
C11170 net67 _450_/a_836_156# 0.008805f
C11171 FILLER_0_8_37/a_124_375# _054_ 0.014206f
C11172 _132_ _145_ 0.010994f
C11173 _136_ FILLER_0_15_180/a_484_472# 0.002128f
C11174 result[8] FILLER_0_24_274/a_1020_375# 0.00726f
C11175 mask\[4\] _047_ 0.080091f
C11176 _424_/a_2665_112# vss 0.013462f
C11177 net26 FILLER_0_23_44/a_1020_375# 0.001646f
C11178 _320_/a_1792_472# state\[1\] 0.001901f
C11179 _210_/a_67_603# _436_/a_2665_112# 0.007103f
C11180 net55 FILLER_0_17_72/a_572_375# 0.023585f
C11181 _093_ FILLER_0_17_104/a_572_375# 0.01418f
C11182 net50 _441_/a_2560_156# 0.008865f
C11183 FILLER_0_7_162/a_124_375# net37 0.011644f
C11184 FILLER_0_21_142/a_572_375# net23 0.007884f
C11185 _443_/a_36_151# _370_/a_848_380# 0.001568f
C11186 _287_/a_36_472# _102_ 0.028733f
C11187 _414_/a_448_472# cal_itt\[3\] 0.109704f
C11188 mask\[4\] _021_ 0.018108f
C11189 net29 mask\[2\] 0.122202f
C11190 net82 FILLER_0_3_212/a_36_472# 0.011542f
C11191 FILLER_0_16_57/a_484_472# net15 0.008573f
C11192 cal input4/a_36_68# 0.054357f
C11193 FILLER_0_8_37/a_572_375# vdd 0.013575f
C11194 FILLER_0_8_37/a_124_375# vss 0.00252f
C11195 _132_ _318_/a_224_472# 0.001097f
C11196 state\[0\] _090_ 0.003121f
C11197 _449_/a_2248_156# _176_ 0.013753f
C11198 FILLER_0_21_28/a_1916_375# _012_ 0.023886f
C11199 _273_/a_36_68# _246_/a_36_68# 0.001168f
C11200 FILLER_0_5_72/a_36_472# vdd 0.107678f
C11201 FILLER_0_5_72/a_1468_375# vss 0.057097f
C11202 mask\[3\] FILLER_0_17_218/a_484_472# 0.017442f
C11203 _031_ FILLER_0_2_111/a_484_472# 0.027347f
C11204 net69 FILLER_0_2_111/a_1380_472# 0.021896f
C11205 _050_ FILLER_0_22_128/a_1020_375# 0.002647f
C11206 net81 FILLER_0_15_235/a_124_375# 0.008139f
C11207 FILLER_0_5_54/a_124_375# trim_mask\[1\] 0.024065f
C11208 FILLER_0_5_54/a_1468_375# _029_ 0.008339f
C11209 FILLER_0_4_144/a_572_375# _081_ 0.002236f
C11210 FILLER_0_4_144/a_124_375# _152_ 0.007333f
C11211 output46/a_224_472# vdd 0.043652f
C11212 _122_ FILLER_0_8_156/a_484_472# 0.007378f
C11213 _057_ _310_/a_741_69# 0.001002f
C11214 net20 output34/a_224_472# 0.023142f
C11215 FILLER_0_20_87/a_124_375# vdd 0.008846f
C11216 _410_/a_36_68# _039_ 0.016062f
C11217 _127_ _017_ 0.005836f
C11218 _449_/a_36_151# _095_ 0.003412f
C11219 _413_/a_1204_472# net65 0.017514f
C11220 _119_ _115_ 0.06747f
C11221 _451_/a_36_151# vss 0.028073f
C11222 _451_/a_448_472# vdd 0.04463f
C11223 _446_/a_1000_472# net40 0.0368f
C11224 _028_ FILLER_0_7_104/a_932_472# 0.003084f
C11225 _247_/a_36_160# _090_ 0.010285f
C11226 _426_/a_36_151# FILLER_0_8_247/a_1468_375# 0.059049f
C11227 ctlp[7] net54 0.004355f
C11228 vdd _166_ 0.108744f
C11229 net74 _062_ 0.062376f
C11230 _375_/a_36_68# vdd 0.010344f
C11231 FILLER_0_16_255/a_36_472# vss 0.00184f
C11232 input4/a_36_68# en 0.064323f
C11233 _421_/a_1000_472# net19 0.03394f
C11234 _187_ _067_ 0.035532f
C11235 result[4] _417_/a_2560_156# 0.001076f
C11236 _093_ FILLER_0_19_134/a_36_472# 0.002415f
C11237 FILLER_0_18_53/a_124_375# FILLER_0_18_37/a_1468_375# 0.012222f
C11238 _363_/a_36_68# vss 0.043707f
C11239 output9/a_224_472# FILLER_0_1_266/a_36_472# 0.001007f
C11240 net45 trimb[3] 0.001109f
C11241 _326_/a_36_160# _115_ 0.051266f
C11242 FILLER_0_14_91/a_484_472# _043_ 0.00134f
C11243 FILLER_0_11_124/a_124_375# vss 0.017354f
C11244 FILLER_0_11_124/a_36_472# vdd 0.005222f
C11245 net54 _148_ 0.098648f
C11246 _267_/a_1568_472# _055_ 0.001681f
C11247 _098_ net22 0.157058f
C11248 _091_ FILLER_0_15_212/a_36_472# 0.007355f
C11249 _412_/a_36_151# net59 0.003938f
C11250 mask\[7\] _009_ 0.078131f
C11251 output36/a_224_472# FILLER_0_14_263/a_124_375# 0.029138f
C11252 _185_ vdd 0.325358f
C11253 net43 vss 0.132286f
C11254 net20 _413_/a_2665_112# 0.015855f
C11255 net66 FILLER_0_3_54/a_124_375# 0.038548f
C11256 net34 FILLER_0_22_128/a_3172_472# 0.003953f
C11257 net20 _298_/a_224_472# 0.001861f
C11258 _086_ _114_ 1.371271f
C11259 net22 _205_/a_36_160# 0.109939f
C11260 input1/a_36_113# input4/a_36_68# 0.015796f
C11261 FILLER_0_14_91/a_572_375# _095_ 0.011885f
C11262 _350_/a_257_69# net23 0.003052f
C11263 _261_/a_36_160# FILLER_0_5_148/a_124_375# 0.005705f
C11264 _056_ net4 0.002408f
C11265 net79 _284_/a_224_472# 0.009327f
C11266 net20 mask\[0\] 0.103301f
C11267 ctln[2] net76 0.001008f
C11268 _419_/a_1000_472# net77 0.001113f
C11269 FILLER_0_18_107/a_36_472# net14 0.005297f
C11270 net63 _106_ 0.034574f
C11271 net34 _050_ 0.004662f
C11272 _372_/a_358_69# _163_ 0.001427f
C11273 state\[1\] _043_ 0.1587f
C11274 FILLER_0_21_150/a_36_472# vss 0.012815f
C11275 _161_ _058_ 0.101968f
C11276 net75 net8 0.553872f
C11277 _112_ net59 0.002846f
C11278 _083_ _080_ 0.043927f
C11279 _136_ _138_ 0.186242f
C11280 _142_ _093_ 0.492191f
C11281 _413_/a_2248_156# net59 0.05485f
C11282 cal_count\[3\] _390_/a_36_68# 0.003074f
C11283 _363_/a_244_472# _053_ 0.001236f
C11284 _128_ _061_ 0.76584f
C11285 vss output30/a_224_472# 0.030732f
C11286 fanout62/a_36_160# _416_/a_36_151# 0.016215f
C11287 FILLER_0_18_2/a_1828_472# _452_/a_1353_112# 0.001313f
C11288 _258_/a_36_160# _079_ 0.026618f
C11289 _129_ _058_ 0.050726f
C11290 ctlp[2] net33 0.004972f
C11291 net34 _210_/a_255_603# 0.002153f
C11292 net54 FILLER_0_19_134/a_36_472# 0.061344f
C11293 FILLER_0_16_57/a_1020_375# FILLER_0_17_64/a_124_375# 0.026339f
C11294 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_124_375# 0.012001f
C11295 FILLER_0_10_37/a_124_375# net16 0.010358f
C11296 FILLER_0_12_50/a_36_472# vss 0.0027f
C11297 output31/a_224_472# _417_/a_2665_112# 0.011048f
C11298 FILLER_0_16_37/a_124_375# net72 0.013591f
C11299 output7/a_224_472# net40 0.009154f
C11300 _428_/a_2665_112# vdd 0.004735f
C11301 net73 fanout71/a_36_113# 0.004833f
C11302 FILLER_0_20_193/a_36_472# net21 0.001099f
C11303 _098_ _433_/a_2665_112# 0.01601f
C11304 fanout53/a_36_160# vdd 0.016868f
C11305 result[9] net62 0.339372f
C11306 output44/a_224_472# net55 0.011586f
C11307 _028_ net14 0.066292f
C11308 FILLER_0_7_72/a_572_375# FILLER_0_6_47/a_3260_375# 0.026339f
C11309 net4 _068_ 0.040977f
C11310 _086_ _176_ 0.837546f
C11311 _437_/a_1204_472# net14 0.004949f
C11312 FILLER_0_4_144/a_36_472# _443_/a_36_151# 0.00271f
C11313 _307_/a_234_472# vdd 0.001209f
C11314 _106_ _069_ 0.006716f
C11315 ctln[1] input5/a_36_113# 0.01908f
C11316 FILLER_0_5_109/a_572_375# net47 0.011047f
C11317 _394_/a_56_524# vss 0.003797f
C11318 _065_ ctln[9] 0.123393f
C11319 FILLER_0_24_274/a_1380_472# FILLER_0_23_282/a_484_472# 0.058411f
C11320 FILLER_0_7_72/a_1916_375# net52 0.001608f
C11321 _070_ net22 0.032551f
C11322 _430_/a_36_151# _092_ 0.002363f
C11323 FILLER_0_5_128/a_36_472# _360_/a_36_160# 0.195479f
C11324 _028_ _164_ 0.019799f
C11325 FILLER_0_9_28/a_3260_375# vdd 0.017581f
C11326 _422_/a_2248_156# _009_ 0.061786f
C11327 _408_/a_56_524# net40 0.001367f
C11328 _407_/a_36_472# vdd 0.095308f
C11329 net20 _099_ 0.011124f
C11330 ctln[7] _442_/a_2248_156# 0.006094f
C11331 _121_ _120_ 0.069685f
C11332 vdd cal_count\[0\] 0.491891f
C11333 _112_ _122_ 0.120159f
C11334 FILLER_0_8_2/a_124_375# _054_ 0.001055f
C11335 FILLER_0_8_107/a_36_472# _133_ 0.00589f
C11336 net36 _094_ 0.086414f
C11337 FILLER_0_11_124/a_36_472# _135_ 0.110114f
C11338 _098_ FILLER_0_15_235/a_572_375# 0.001343f
C11339 _091_ FILLER_0_12_220/a_932_472# 0.001638f
C11340 FILLER_0_18_2/a_932_472# vdd 0.002342f
C11341 FILLER_0_20_177/a_484_472# _098_ 0.009817f
C11342 FILLER_0_8_127/a_124_375# _124_ 0.022175f
C11343 net27 FILLER_0_10_247/a_124_375# 0.015466f
C11344 output35/a_224_472# net35 0.007217f
C11345 _143_ _343_/a_49_472# 0.00918f
C11346 _072_ _128_ 0.072191f
C11347 _068_ _311_/a_1660_473# 0.003542f
C11348 FILLER_0_14_81/a_36_472# _095_ 0.014706f
C11349 FILLER_0_18_177/a_1916_375# net21 0.004339f
C11350 net20 _294_/a_224_472# 0.008053f
C11351 _086_ _124_ 0.063099f
C11352 net60 _420_/a_2248_156# 0.035104f
C11353 net15 FILLER_0_5_54/a_572_375# 0.002259f
C11354 _098_ vdd 2.272938f
C11355 mask\[5\] FILLER_0_19_195/a_36_472# 0.007596f
C11356 _412_/a_448_472# net18 0.049704f
C11357 ctln[6] net52 0.1064f
C11358 net54 _436_/a_2665_112# 0.042428f
C11359 output44/a_224_472# net17 0.07836f
C11360 _110_ _012_ 0.046196f
C11361 _413_/a_448_472# net21 0.052657f
C11362 _424_/a_448_472# _012_ 0.007299f
C11363 trim_mask\[1\] FILLER_0_6_47/a_2276_472# 0.006166f
C11364 _073_ FILLER_0_3_221/a_1380_472# 0.045839f
C11365 _033_ _444_/a_448_472# 0.047424f
C11366 _118_ _315_/a_716_497# 0.001968f
C11367 _205_/a_36_160# vdd 0.016131f
C11368 FILLER_0_8_2/a_36_472# vdd 0.104141f
C11369 FILLER_0_8_2/a_124_375# vss 0.003001f
C11370 fanout51/a_36_113# FILLER_0_9_72/a_36_472# 0.001391f
C11371 _028_ FILLER_0_7_72/a_2364_375# 0.003884f
C11372 net19 net18 0.028285f
C11373 net67 _439_/a_36_151# 0.136402f
C11374 FILLER_0_13_228/a_36_472# vss 0.006491f
C11375 FILLER_0_18_2/a_2812_375# net55 0.007169f
C11376 FILLER_0_19_47/a_572_375# vdd 0.019566f
C11377 FILLER_0_19_47/a_124_375# vss 0.002211f
C11378 net18 _416_/a_796_472# 0.007144f
C11379 net19 _196_/a_36_160# 0.027835f
C11380 net35 FILLER_0_22_86/a_124_375# 0.01209f
C11381 mask\[8\] FILLER_0_22_86/a_572_375# 0.013048f
C11382 _432_/a_448_472# mask\[3\] 0.005831f
C11383 FILLER_0_16_107/a_484_472# _136_ 0.013449f
C11384 net44 FILLER_0_15_10/a_124_375# 0.009108f
C11385 FILLER_0_15_10/a_36_472# vss 0.002605f
C11386 fanout49/a_36_160# vdd 0.099887f
C11387 _141_ FILLER_0_22_128/a_3172_472# 0.01947f
C11388 output11/a_224_472# _000_ 0.006606f
C11389 FILLER_0_7_59/a_124_375# vdd -0.006113f
C11390 _178_ FILLER_0_15_10/a_36_472# 0.001356f
C11391 FILLER_0_13_212/a_124_375# _043_ 0.011912f
C11392 FILLER_0_22_128/a_2812_375# _146_ 0.001336f
C11393 net35 FILLER_0_22_128/a_932_472# 0.007806f
C11394 net17 _452_/a_1293_527# 0.001011f
C11395 _235_/a_67_603# net17 0.018056f
C11396 FILLER_0_5_164/a_572_375# net22 0.002238f
C11397 FILLER_0_7_72/a_572_375# FILLER_0_5_72/a_484_472# 0.001512f
C11398 fanout64/a_36_160# vdd 0.010802f
C11399 _383_/a_36_472# trim_mask\[3\] 0.003193f
C11400 _387_/a_36_113# vdd 0.041853f
C11401 net59 FILLER_0_3_212/a_124_375# 0.057221f
C11402 trimb[0] FILLER_0_20_2/a_124_375# 0.006864f
C11403 net20 FILLER_0_1_212/a_36_472# 0.013846f
C11404 FILLER_0_18_177/a_3260_375# net22 0.049279f
C11405 net81 net76 0.236554f
C11406 net17 FILLER_0_23_44/a_124_375# 0.007634f
C11407 net65 _386_/a_848_380# 0.00123f
C11408 fanout66/a_36_113# _441_/a_36_151# 0.032681f
C11409 net60 _419_/a_2665_112# 0.059916f
C11410 mask\[5\] FILLER_0_18_177/a_2276_472# 0.001063f
C11411 _444_/a_1000_472# net40 0.038229f
C11412 output42/a_224_472# net38 0.066219f
C11413 net20 FILLER_0_12_220/a_1020_375# 0.047331f
C11414 net54 FILLER_0_22_128/a_1468_375# 0.004731f
C11415 output45/a_224_472# output43/a_224_472# 0.246888f
C11416 FILLER_0_17_104/a_1380_472# vss 0.001141f
C11417 _070_ FILLER_0_9_105/a_36_472# 0.023853f
C11418 _326_/a_36_160# _134_ 0.003299f
C11419 _143_ _093_ 0.003295f
C11420 FILLER_0_18_2/a_2812_375# net17 0.012909f
C11421 _077_ _439_/a_448_472# 0.052962f
C11422 _013_ FILLER_0_17_56/a_572_375# 0.001047f
C11423 FILLER_0_8_24/a_484_472# net40 0.004383f
C11424 _039_ output6/a_224_472# 0.012051f
C11425 result[1] result[2] 0.072492f
C11426 FILLER_0_16_107/a_36_472# _131_ 0.008817f
C11427 _083_ vss 0.0284f
C11428 _070_ vdd 1.546772f
C11429 _115_ _129_ 0.021405f
C11430 FILLER_0_18_107/a_1020_375# FILLER_0_17_104/a_1380_472# 0.001597f
C11431 ctln[1] net19 0.001327f
C11432 _056_ _058_ 0.988919f
C11433 FILLER_0_17_72/a_1380_472# _438_/a_36_151# 0.001221f
C11434 output10/a_224_472# vss 0.014205f
C11435 _432_/a_36_151# vdd 0.173104f
C11436 net47 net14 0.033547f
C11437 FILLER_0_15_180/a_124_375# vdd 0.016985f
C11438 FILLER_0_7_146/a_36_472# vdd 0.072981f
C11439 FILLER_0_7_146/a_124_375# vss 0.050543f
C11440 FILLER_0_6_90/a_572_375# _439_/a_2665_112# 0.001646f
C11441 net33 net21 0.052426f
C11442 _009_ _298_/a_224_472# 0.002441f
C11443 output35/a_224_472# net22 0.028095f
C11444 FILLER_0_22_86/a_1380_472# FILLER_0_22_107/a_36_472# 0.001963f
C11445 _053_ _054_ 0.015389f
C11446 result[7] FILLER_0_24_290/a_124_375# 0.005026f
C11447 net56 FILLER_0_17_161/a_124_375# 0.001108f
C11448 net82 net22 1.960347f
C11449 _132_ FILLER_0_18_107/a_2812_375# 0.002706f
C11450 net47 _164_ 0.118311f
C11451 FILLER_0_21_28/a_124_375# net40 0.060428f
C11452 net32 net61 0.056005f
C11453 trim_mask\[2\] FILLER_0_3_78/a_124_375# 0.010185f
C11454 _321_/a_170_472# _120_ 0.040613f
C11455 FILLER_0_9_28/a_3260_375# fanout67/a_36_160# 0.001925f
C11456 net23 _066_ 0.031928f
C11457 _096_ _320_/a_1120_472# 0.004315f
C11458 _420_/a_36_151# net18 0.001426f
C11459 fanout57/a_36_113# net22 0.024465f
C11460 FILLER_0_14_50/a_124_375# vdd 0.026996f
C11461 net34 _435_/a_36_151# 0.011954f
C11462 output47/a_224_472# cal_count\[2\] 0.080405f
C11463 FILLER_0_6_239/a_124_375# _074_ 0.010359f
C11464 result[9] _417_/a_2560_156# 0.00263f
C11465 FILLER_0_17_72/a_2724_472# _131_ 0.004095f
C11466 _176_ _451_/a_3129_107# 0.021559f
C11467 FILLER_0_5_109/a_572_375# _154_ 0.014669f
C11468 _127_ cal_count\[3\] 0.306114f
C11469 _420_/a_1204_472# _009_ 0.009314f
C11470 _086_ _267_/a_36_472# 0.070088f
C11471 _053_ vss 0.85895f
C11472 _144_ _437_/a_2665_112# 0.001186f
C11473 _133_ _125_ 0.014858f
C11474 _068_ _058_ 0.092852f
C11475 net55 vdd 1.248648f
C11476 net68 FILLER_0_8_37/a_36_472# 0.001088f
C11477 _431_/a_1308_423# net73 0.039024f
C11478 _127_ _059_ 0.002878f
C11479 cal_count\[3\] _453_/a_448_472# 0.001494f
C11480 result[6] _010_ 0.056004f
C11481 output47/a_224_472# input3/a_36_113# 0.001371f
C11482 result[7] FILLER_0_24_274/a_1380_472# 0.006454f
C11483 _095_ _451_/a_36_151# 0.008311f
C11484 _005_ _100_ 0.004305f
C11485 _074_ _251_/a_468_472# 0.001217f
C11486 FILLER_0_12_136/a_932_472# FILLER_0_11_142/a_124_375# 0.001543f
C11487 _074_ net19 0.035973f
C11488 FILLER_0_5_54/a_1380_472# vss 0.007301f
C11489 FILLER_0_15_142/a_572_375# _427_/a_36_151# 0.059049f
C11490 FILLER_0_17_72/a_484_472# net36 0.001629f
C11491 cal_count\[3\] FILLER_0_11_135/a_36_472# 0.005101f
C11492 FILLER_0_7_104/a_932_472# _154_ 0.002023f
C11493 _346_/a_49_472# _140_ 0.003436f
C11494 _093_ _438_/a_796_472# 0.001924f
C11495 _075_ _053_ 0.634359f
C11496 output23/a_224_472# ctlp[6] 0.024575f
C11497 mask\[9\] _438_/a_1308_423# 0.044336f
C11498 FILLER_0_5_164/a_572_375# vdd 0.0042f
C11499 net74 net14 0.034568f
C11500 _026_ FILLER_0_20_87/a_36_472# 0.004568f
C11501 _091_ _019_ 0.031681f
C11502 net41 cal_count\[2\] 0.079279f
C11503 output39/a_224_472# net40 0.087367f
C11504 _182_ vss 0.068928f
C11505 net15 FILLER_0_6_47/a_2724_472# 0.006158f
C11506 net58 vdd 0.929215f
C11507 _178_ _182_ 0.067534f
C11508 net68 _160_ 0.072339f
C11509 fanout55/a_36_160# net74 0.016856f
C11510 FILLER_0_18_177/a_3260_375# vdd 0.003399f
C11511 _449_/a_2560_156# _067_ 0.007511f
C11512 net20 FILLER_0_3_221/a_572_375# 0.004331f
C11513 FILLER_0_7_59/a_124_375# fanout67/a_36_160# 0.001597f
C11514 net66 FILLER_0_5_54/a_124_375# 0.002093f
C11515 FILLER_0_11_101/a_36_472# cal_count\[3\] 0.005101f
C11516 net18 _419_/a_448_472# 0.037373f
C11517 net75 _425_/a_1204_472# 0.015778f
C11518 mask\[4\] FILLER_0_18_209/a_572_375# 0.032112f
C11519 net16 FILLER_0_18_37/a_36_472# 0.001132f
C11520 FILLER_0_15_282/a_484_472# _006_ 0.00444f
C11521 net17 vdd 2.139315f
C11522 net20 _000_ 0.159624f
C11523 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_124_375# 0.012221f
C11524 net69 _441_/a_1308_423# 0.016223f
C11525 _035_ _064_ 0.02225f
C11526 calibrate FILLER_0_9_270/a_124_375# 0.002292f
C11527 trim_val\[1\] vdd 0.173304f
C11528 FILLER_0_7_72/a_1020_375# FILLER_0_5_72/a_932_472# 0.001512f
C11529 FILLER_0_21_125/a_124_375# _144_ 0.009117f
C11530 _201_/a_67_603# _047_ 0.013357f
C11531 _028_ _153_ 0.008011f
C11532 _425_/a_36_151# vss 0.00158f
C11533 _425_/a_448_472# vdd 0.029071f
C11534 net41 FILLER_0_19_28/a_484_472# 0.047447f
C11535 net73 FILLER_0_18_107/a_1380_472# 0.039646f
C11536 mask\[7\] FILLER_0_22_128/a_3260_375# 0.00186f
C11537 net17 FILLER_0_20_15/a_484_472# 0.011079f
C11538 _412_/a_1308_423# cal_itt\[1\] 0.009991f
C11539 _156_ _160_ 0.299745f
C11540 FILLER_0_15_116/a_36_472# FILLER_0_14_107/a_1020_375# 0.001723f
C11541 FILLER_0_15_116/a_572_375# FILLER_0_14_107/a_1468_375# 0.026339f
C11542 mask\[7\] net33 0.02491f
C11543 FILLER_0_23_60/a_124_375# FILLER_0_23_44/a_1468_375# 0.012001f
C11544 FILLER_0_24_290/a_36_472# vss 0.007621f
C11545 output35/a_224_472# vdd 0.064053f
C11546 net53 _427_/a_1308_423# 0.007426f
C11547 _122_ _120_ 0.143427f
C11548 net57 _067_ 0.018966f
C11549 _248_/a_36_68# _060_ 0.004581f
C11550 net67 FILLER_0_8_37/a_36_472# 0.001479f
C11551 _448_/a_36_151# net12 0.133216f
C11552 _448_/a_1308_423# net22 0.045644f
C11553 _082_ vdd 0.191411f
C11554 _428_/a_2560_156# _043_ 0.009909f
C11555 net82 vdd 1.014512f
C11556 FILLER_0_18_76/a_124_375# _438_/a_36_151# 0.001252f
C11557 _428_/a_36_151# net74 0.020444f
C11558 cal_itt\[2\] FILLER_0_3_221/a_36_472# 0.003825f
C11559 net50 _439_/a_448_472# 0.020872f
C11560 net52 _439_/a_796_472# 0.003099f
C11561 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_36_472# 0.086742f
C11562 _445_/a_2665_112# net49 0.03968f
C11563 _137_ vss 0.343959f
C11564 mask\[9\] net36 1.116767f
C11565 _098_ FILLER_0_16_154/a_572_375# 0.001791f
C11566 net63 _098_ 0.055686f
C11567 fanout57/a_36_113# vdd 0.005473f
C11568 net27 _425_/a_2665_112# 0.001323f
C11569 net80 net33 0.037227f
C11570 output36/a_224_472# vss -0.002521f
C11571 _013_ FILLER_0_18_53/a_572_375# 0.015534f
C11572 _327_/a_36_472# vdd 0.00142f
C11573 _239_/a_36_160# net68 0.043367f
C11574 _238_/a_67_603# vdd 0.004498f
C11575 _443_/a_2665_112# _037_ 0.004052f
C11576 _043_ FILLER_0_13_80/a_124_375# 0.013485f
C11577 state\[2\] FILLER_0_13_142/a_1380_472# 0.019965f
C11578 net63 _434_/a_3041_156# 0.001449f
C11579 _431_/a_448_472# _136_ 0.064724f
C11580 _091_ FILLER_0_13_212/a_484_472# 0.04953f
C11581 FILLER_0_17_226/a_36_472# _008_ 0.001842f
C11582 _274_/a_36_68# _072_ 0.001647f
C11583 FILLER_0_3_78/a_36_472# vss 0.004461f
C11584 net67 _160_ 0.003659f
C11585 _114_ _061_ 0.123371f
C11586 result[7] _010_ 0.054533f
C11587 FILLER_0_2_127/a_36_472# vss 0.002567f
C11588 _394_/a_56_524# _095_ 0.10007f
C11589 FILLER_0_22_86/a_124_375# vdd 0.024158f
C11590 _104_ FILLER_0_17_226/a_124_375# 0.024833f
C11591 _152_ _058_ 0.00259f
C11592 _415_/a_36_151# FILLER_0_11_282/a_124_375# 0.001822f
C11593 net58 net9 0.018829f
C11594 _154_ net14 0.02512f
C11595 _114_ _311_/a_66_473# 0.081048f
C11596 FILLER_0_22_128/a_932_472# vdd 0.004405f
C11597 FILLER_0_22_128/a_484_472# vss 0.002338f
C11598 mask\[6\] _146_ 0.181681f
C11599 _216_/a_67_603# vdd 0.030831f
C11600 FILLER_0_17_226/a_124_375# vss 0.025007f
C11601 net41 _043_ 0.03188f
C11602 _412_/a_2560_156# cal_itt\[1\] 0.00454f
C11603 _077_ _256_/a_36_68# 0.027906f
C11604 _049_ vss 0.026036f
C11605 net15 fanout72/a_36_113# 0.010284f
C11606 net56 FILLER_0_18_139/a_1020_375# 0.018398f
C11607 _411_/a_1308_423# vss 0.0013f
C11608 net75 FILLER_0_8_263/a_124_375# 0.001386f
C11609 output27/a_224_472# FILLER_0_8_263/a_36_472# 0.002002f
C11610 FILLER_0_12_20/a_36_472# net6 0.007073f
C11611 _441_/a_2665_112# FILLER_0_3_78/a_572_375# 0.010688f
C11612 _063_ FILLER_0_6_47/a_36_472# 0.007244f
C11613 _116_ _248_/a_36_68# 0.007314f
C11614 _174_ cal_count\[1\] 0.081252f
C11615 output17/a_224_472# net17 0.09023f
C11616 _132_ FILLER_0_16_115/a_36_472# 0.015199f
C11617 _069_ _098_ 0.029447f
C11618 _088_ FILLER_0_3_172/a_2724_472# 0.005827f
C11619 _086_ FILLER_0_7_104/a_1380_472# 0.034829f
C11620 _111_ vdd 0.3227f
C11621 _115_ _068_ 0.889978f
C11622 FILLER_0_16_241/a_36_472# mask\[2\] 0.025337f
C11623 net64 FILLER_0_11_282/a_124_375# 0.023042f
C11624 net82 FILLER_0_3_172/a_2812_375# 0.010439f
C11625 _140_ _147_ 0.08953f
C11626 FILLER_0_7_72/a_36_472# vss 0.033878f
C11627 _276_/a_36_160# vss 0.02914f
C11628 _092_ mask\[3\] 0.040554f
C11629 net46 net41 0.061224f
C11630 _004_ _415_/a_796_472# 0.005395f
C11631 _114_ FILLER_0_11_101/a_484_472# 0.025975f
C11632 _431_/a_448_472# fanout70/a_36_113# 0.001157f
C11633 FILLER_0_3_172/a_1916_375# net65 0.003745f
C11634 net9 _082_ 0.001006f
C11635 _412_/a_448_472# net65 0.043862f
C11636 _446_/a_1308_423# vdd 0.002346f
C11637 _035_ output38/a_224_472# 0.091395f
C11638 FILLER_0_18_2/a_572_375# net38 0.007477f
C11639 net82 net9 0.004599f
C11640 _077_ _162_ 0.013298f
C11641 _114_ _072_ 0.078148f
C11642 net41 net68 0.009755f
C11643 output28/a_224_472# net18 0.015144f
C11644 result[7] FILLER_0_23_282/a_36_472# 0.014869f
C11645 net72 _179_ 0.083699f
C11646 net35 net21 0.001845f
C11647 _316_/a_124_24# _123_ 0.009391f
C11648 FILLER_0_18_2/a_124_375# net44 0.051228f
C11649 FILLER_0_15_116/a_572_375# vdd 0.017636f
C11650 net65 net19 0.044106f
C11651 net63 _432_/a_36_151# 0.001392f
C11652 _076_ _226_/a_1044_68# 0.0023f
C11653 FILLER_0_12_136/a_572_375# net23 0.00281f
C11654 net20 fanout75/a_36_113# 0.001027f
C11655 _105_ _422_/a_2665_112# 0.011125f
C11656 _077_ _131_ 0.03465f
C11657 _095_ FILLER_0_15_10/a_36_472# 0.00335f
C11658 net20 FILLER_0_13_212/a_572_375# 0.002085f
C11659 _291_/a_36_160# _093_ 0.017281f
C11660 net57 _066_ 0.069098f
C11661 net27 FILLER_0_14_235/a_36_472# 0.003401f
C11662 _448_/a_1308_423# vdd 0.006042f
C11663 net47 _153_ 0.755476f
C11664 FILLER_0_3_142/a_36_472# net23 0.043034f
C11665 net20 _421_/a_1000_472# 0.012469f
C11666 _182_ _401_/a_36_68# 0.088487f
C11667 _442_/a_36_151# net13 0.009343f
C11668 net15 FILLER_0_17_56/a_124_375# 0.001854f
C11669 FILLER_0_5_54/a_572_375# net47 0.009717f
C11670 FILLER_0_7_59/a_572_375# net68 0.005738f
C11671 net26 FILLER_0_21_28/a_1828_472# 0.010367f
C11672 net55 _423_/a_2560_156# 0.002265f
C11673 net1 net59 0.920133f
C11674 _176_ FILLER_0_11_101/a_484_472# 0.001777f
C11675 _257_/a_36_472# _068_ 0.002986f
C11676 FILLER_0_14_263/a_36_472# vss 0.003195f
C11677 fanout57/a_36_113# FILLER_0_2_165/a_124_375# 0.008057f
C11678 net40 net6 0.00772f
C11679 net57 net23 0.324262f
C11680 _431_/a_448_472# net53 0.002087f
C11681 _072_ _176_ 0.298077f
C11682 _069_ _070_ 0.257147f
C11683 _386_/a_692_472# _169_ 0.004014f
C11684 _386_/a_848_380# _163_ 0.026484f
C11685 FILLER_0_13_65/a_124_375# net72 0.002341f
C11686 _177_ fanout55/a_36_160# 0.002687f
C11687 FILLER_0_17_72/a_1916_375# vdd 0.002595f
C11688 FILLER_0_17_72/a_1468_375# vss 0.003461f
C11689 FILLER_0_18_2/a_1380_472# net38 0.029747f
C11690 FILLER_0_12_20/a_124_375# net47 0.047331f
C11691 ctlp[2] vdd 0.617599f
C11692 _144_ _148_ 0.038002f
C11693 ctlp[5] ctlp[4] 0.001257f
C11694 FILLER_0_4_107/a_36_472# vdd 0.119007f
C11695 FILLER_0_4_107/a_1468_375# vss 0.055184f
C11696 FILLER_0_16_89/a_1380_472# _451_/a_1353_112# 0.010457f
C11697 FILLER_0_2_111/a_484_472# _158_ 0.003604f
C11698 _028_ FILLER_0_6_47/a_2724_472# 0.023218f
C11699 net41 net67 0.03408f
C11700 net20 _256_/a_36_68# 0.02797f
C11701 FILLER_0_9_270/a_36_472# vss 0.001642f
C11702 FILLER_0_9_270/a_484_472# vdd 0.006354f
C11703 calibrate net22 0.036525f
C11704 net52 FILLER_0_2_111/a_1020_375# 0.00245f
C11705 output19/a_224_472# _422_/a_2665_112# 0.024396f
C11706 _091_ _429_/a_1000_472# 0.029742f
C11707 _424_/a_2248_156# FILLER_0_21_60/a_124_375# 0.001068f
C11708 net31 net30 0.130396f
C11709 FILLER_0_2_101/a_124_375# _367_/a_36_68# 0.001176f
C11710 trim_mask\[2\] _167_ 0.027204f
C11711 net52 _440_/a_1308_423# 0.047012f
C11712 FILLER_0_21_133/a_36_472# _098_ 0.002964f
C11713 net61 _421_/a_2665_112# 0.001339f
C11714 net60 _421_/a_1204_472# 0.021679f
C11715 FILLER_0_4_197/a_1380_472# _081_ 0.001345f
C11716 output11/a_224_472# ctln[1] 0.004299f
C11717 FILLER_0_16_89/a_932_472# _131_ 0.008223f
C11718 FILLER_0_10_78/a_1468_375# vss 0.054053f
C11719 net22 net21 1.937266f
C11720 net50 FILLER_0_8_37/a_484_472# 0.003311f
C11721 FILLER_0_12_136/a_1380_472# _126_ 0.014722f
C11722 fanout71/a_36_113# _433_/a_36_151# 0.138322f
C11723 FILLER_0_18_2/a_2276_472# _452_/a_1040_527# 0.008652f
C11724 _431_/a_2665_112# _136_ 0.035394f
C11725 FILLER_0_11_142/a_572_375# _120_ 0.009014f
C11726 _273_/a_36_68# net4 0.06843f
C11727 _408_/a_1336_472# vdd 0.040992f
C11728 FILLER_0_23_282/a_484_472# vss 0.005378f
C11729 net41 _445_/a_448_472# 0.002211f
C11730 net62 _044_ 0.101165f
C11731 net41 FILLER_0_21_28/a_484_472# 0.060027f
C11732 FILLER_0_13_142/a_484_472# vss 0.024835f
C11733 net49 _440_/a_1308_423# 0.022006f
C11734 net35 mask\[7\] 0.954332f
C11735 _235_/a_67_603# trim_mask\[2\] 0.022726f
C11736 FILLER_0_7_59/a_572_375# net67 0.007538f
C11737 _412_/a_1204_472# net81 0.003435f
C11738 _414_/a_36_151# net22 0.014398f
C11739 FILLER_0_19_142/a_36_472# vss 0.011026f
C11740 ctlp[8] net25 0.055914f
C11741 FILLER_0_17_56/a_484_472# FILLER_0_18_61/a_36_472# 0.026657f
C11742 _040_ vss 0.216709f
C11743 _323_/a_36_113# _015_ 0.003795f
C11744 output33/a_224_472# net61 0.04987f
C11745 cal_count\[3\] _060_ 0.007037f
C11746 _447_/a_1308_423# vdd 0.004739f
C11747 net63 output35/a_224_472# 0.148302f
C11748 FILLER_0_16_89/a_572_375# net36 0.003629f
C11749 _174_ _120_ 0.002521f
C11750 net80 net35 0.028982f
C11751 result[2] net30 0.019568f
C11752 _057_ _055_ 0.290639f
C11753 FILLER_0_10_78/a_1468_375# _308_/a_124_24# 0.001565f
C11754 _137_ FILLER_0_16_154/a_1020_375# 0.010692f
C11755 _414_/a_2248_156# net59 0.004437f
C11756 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_484_472# 0.026657f
C11757 FILLER_0_5_72/a_572_375# _440_/a_36_151# 0.035849f
C11758 trim[4] net42 0.016428f
C11759 _321_/a_170_472# _125_ 0.008492f
C11760 _450_/a_2225_156# net40 0.04513f
C11761 FILLER_0_17_226/a_36_472# _093_ 0.004282f
C11762 _447_/a_2665_112# _441_/a_36_151# 0.028591f
C11763 _104_ result[6] 0.096535f
C11764 _414_/a_448_472# net22 0.047364f
C11765 FILLER_0_11_101/a_572_375# _134_ 0.0024f
C11766 net20 _429_/a_36_151# 0.002103f
C11767 vss FILLER_0_10_94/a_572_375# 0.013232f
C11768 vdd FILLER_0_10_94/a_36_472# 0.086035f
C11769 _444_/a_448_472# _054_ 0.017318f
C11770 net82 FILLER_0_2_177/a_572_375# 0.003837f
C11771 result[6] vss 0.310169f
C11772 trimb[1] FILLER_0_18_2/a_2364_375# 0.001523f
C11773 _093_ FILLER_0_18_177/a_3172_472# 0.003708f
C11774 ctln[4] _413_/a_2248_156# 0.001253f
C11775 FILLER_0_8_24/a_124_375# _054_ 0.008177f
C11776 _261_/a_36_160# FILLER_0_5_136/a_124_375# 0.003477f
C11777 _119_ _322_/a_124_24# 0.020461f
C11778 net20 net18 0.025322f
C11779 _057_ _126_ 0.022413f
C11780 cal_count\[1\] FILLER_0_15_59/a_124_375# 0.010034f
C11781 net7 _065_ 0.0295f
C11782 net75 _123_ 0.173358f
C11783 mask\[5\] _091_ 0.048311f
C11784 _154_ _153_ 0.719561f
C11785 _119_ FILLER_0_8_156/a_484_472# 0.00979f
C11786 _116_ cal_count\[3\] 0.384121f
C11787 _449_/a_796_472# net72 0.00138f
C11788 _449_/a_36_151# net55 0.003388f
C11789 output45/a_224_472# trimb[0] 0.003753f
C11790 _025_ _436_/a_796_472# 0.026852f
C11791 FILLER_0_9_28/a_1468_375# net16 0.005202f
C11792 net75 _073_ 0.34505f
C11793 _077_ FILLER_0_8_107/a_124_375# 0.010439f
C11794 _077_ _074_ 0.148596f
C11795 calibrate vdd 0.857987f
C11796 fanout54/a_36_160# vdd 0.008482f
C11797 _078_ FILLER_0_3_221/a_124_375# 0.002694f
C11798 _126_ _250_/a_36_68# 0.022134f
C11799 net64 FILLER_0_15_235/a_124_375# 0.025203f
C11800 result[0] net64 0.09782f
C11801 FILLER_0_16_37/a_124_375# vdd 0.038329f
C11802 _444_/a_1308_423# vdd 0.005677f
C11803 _326_/a_36_160# _322_/a_124_24# 0.004397f
C11804 _289_/a_244_68# _103_ 0.001153f
C11805 _414_/a_2248_156# _122_ 0.002838f
C11806 cal_count\[3\] _408_/a_718_524# 0.005968f
C11807 FILLER_0_10_256/a_124_375# vdd 0.041848f
C11808 FILLER_0_8_24/a_572_375# vdd 0.011353f
C11809 net34 net23 0.058486f
C11810 result[8] FILLER_0_21_206/a_36_472# 0.001292f
C11811 ctln[5] net76 0.001707f
C11812 _077_ _076_ 1.895143f
C11813 _096_ FILLER_0_12_196/a_124_375# 0.002309f
C11814 fanout59/a_36_160# vss 0.010949f
C11815 mask\[7\] net22 0.275179f
C11816 _411_/a_2248_156# cal_itt\[0\] 0.006897f
C11817 net21 vdd 1.653552f
C11818 _431_/a_2665_112# net53 0.004057f
C11819 net38 _452_/a_36_151# 0.010095f
C11820 _333_/a_36_160# vdd 0.107883f
C11821 net50 fanout68/a_36_113# 0.020067f
C11822 output32/a_224_472# net30 0.001139f
C11823 FILLER_0_4_49/a_124_375# net68 0.008422f
C11824 _028_ _376_/a_36_160# 0.026437f
C11825 _371_/a_36_113# _370_/a_124_24# 0.008354f
C11826 output46/a_224_472# net43 0.10562f
C11827 _072_ _267_/a_36_472# 0.024239f
C11828 _438_/a_448_472# net14 0.020612f
C11829 FILLER_0_2_93/a_572_375# vss 0.055237f
C11830 _414_/a_36_151# vdd 0.166006f
C11831 cal_count\[3\] _118_ 0.009058f
C11832 FILLER_0_19_171/a_484_472# vss 0.001913f
C11833 FILLER_0_19_171/a_932_472# vdd 0.011399f
C11834 output8/a_224_472# vdd 0.023187f
C11835 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_572_375# 0.086635f
C11836 mask\[8\] _437_/a_1308_423# 0.001928f
C11837 _288_/a_224_472# _006_ 0.001278f
C11838 net57 FILLER_0_3_142/a_36_472# 0.002298f
C11839 _053_ _385_/a_36_68# 0.018437f
C11840 _118_ _059_ 0.022651f
C11841 net23 FILLER_0_5_148/a_572_375# 0.039975f
C11842 FILLER_0_8_138/a_124_375# _119_ 0.006523f
C11843 _277_/a_36_160# net30 0.014059f
C11844 net20 ctln[1] 0.135151f
C11845 net44 _452_/a_3129_107# 0.067848f
C11846 net60 result[3] 0.001124f
C11847 _430_/a_1308_423# net21 0.008506f
C11848 fanout56/a_36_113# vss 0.03072f
C11849 _103_ _288_/a_224_472# 0.002992f
C11850 FILLER_0_21_28/a_124_375# FILLER_0_20_15/a_1468_375# 0.026339f
C11851 trim_mask\[2\] vdd 0.376424f
C11852 net47 FILLER_0_5_148/a_36_472# 0.004409f
C11853 FILLER_0_6_239/a_36_472# _122_ 0.01785f
C11854 _144_ _207_/a_67_603# 0.064623f
C11855 _024_ FILLER_0_22_177/a_36_472# 0.003242f
C11856 output35/a_224_472# _435_/a_2665_112# 0.008469f
C11857 FILLER_0_2_93/a_124_375# _441_/a_2665_112# 0.006271f
C11858 net16 _446_/a_2665_112# 0.045966f
C11859 _140_ _098_ 0.647503f
C11860 _282_/a_36_160# _098_ 0.00388f
C11861 _055_ _310_/a_49_472# 0.00384f
C11862 _410_/a_36_68# vdd 0.039824f
C11863 FILLER_0_23_44/a_1468_375# vdd -0.013698f
C11864 FILLER_0_16_89/a_36_472# _397_/a_36_472# 0.004546f
C11865 net15 _441_/a_448_472# 0.049213f
C11866 _104_ result[7] 0.475003f
C11867 FILLER_0_18_209/a_572_375# _201_/a_67_603# 0.008812f
C11868 _408_/a_728_93# cal_count\[2\] 0.001568f
C11869 FILLER_0_7_59/a_572_375# FILLER_0_6_47/a_1916_375# 0.05841f
C11870 net12 vss 0.043754f
C11871 mask\[1\] net22 0.029526f
C11872 _414_/a_448_472# vdd 0.013377f
C11873 _440_/a_2248_156# net47 0.017063f
C11874 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_484_472# 0.013276f
C11875 FILLER_0_7_72/a_2812_375# vdd 0.02125f
C11876 _418_/a_36_151# vss 0.041728f
C11877 FILLER_0_14_107/a_484_472# vss -0.001894f
C11878 FILLER_0_14_107/a_932_472# vdd 0.006908f
C11879 result[7] vss 0.49466f
C11880 _448_/a_448_472# FILLER_0_2_177/a_36_472# 0.001927f
C11881 _448_/a_36_151# FILLER_0_2_177/a_484_472# 0.059367f
C11882 FILLER_0_3_172/a_2812_375# net21 0.015743f
C11883 _433_/a_1308_423# _022_ 0.015376f
C11884 clk vdd 0.053789f
C11885 _056_ FILLER_0_12_196/a_124_375# 0.027077f
C11886 FILLER_0_22_177/a_1468_375# net33 0.017455f
C11887 cal_itt\[3\] _162_ 0.141474f
C11888 result[4] net60 0.244453f
C11889 _414_/a_2665_112# _072_ 0.025361f
C11890 FILLER_0_16_255/a_124_375# net30 0.001055f
C11891 FILLER_0_17_72/a_2364_375# _150_ 0.001083f
C11892 FILLER_0_15_116/a_124_375# _095_ 0.002659f
C11893 FILLER_0_21_286/a_124_375# vss 0.005049f
C11894 FILLER_0_21_286/a_572_375# vdd 0.03062f
C11895 _445_/a_1308_423# net17 0.002172f
C11896 _120_ _450_/a_3129_107# 0.001598f
C11897 _437_/a_2665_112# FILLER_0_22_107/a_484_472# 0.007376f
C11898 net50 _220_/a_67_603# 0.005566f
C11899 FILLER_0_9_223/a_484_472# vdd 0.004285f
C11900 FILLER_0_21_28/a_572_375# FILLER_0_20_31/a_124_375# 0.026339f
C11901 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_572_375# 0.086635f
C11902 net20 _074_ 0.038279f
C11903 net50 FILLER_0_7_59/a_36_472# 0.01018f
C11904 _016_ _126_ 0.051451f
C11905 ctln[3] vss 0.133697f
C11906 _402_/a_728_93# _180_ 0.008035f
C11907 FILLER_0_3_54/a_36_472# _381_/a_36_472# 0.010679f
C11908 _091_ net27 0.023019f
C11909 _143_ _144_ 0.001774f
C11910 FILLER_0_18_61/a_124_375# vdd 0.022663f
C11911 _136_ FILLER_0_16_154/a_1380_472# 0.006517f
C11912 net62 FILLER_0_15_212/a_1468_375# 0.001106f
C11913 _428_/a_1000_472# _131_ 0.035998f
C11914 output11/a_224_472# net65 0.001529f
C11915 _334_/a_36_160# vss 0.002713f
C11916 net52 _037_ 0.103749f
C11917 fanout66/a_36_113# _030_ 0.038252f
C11918 net20 _076_ 0.228128f
C11919 mask\[7\] vdd 1.098711f
C11920 net40 trim[3] 0.084824f
C11921 net70 net14 0.106631f
C11922 FILLER_0_14_81/a_36_472# net55 0.015878f
C11923 vdd FILLER_0_4_91/a_124_375# 0.019812f
C11924 FILLER_0_8_247/a_36_472# _316_/a_124_24# 0.001386f
C11925 _074_ FILLER_0_6_231/a_572_375# 0.009029f
C11926 net15 cal_count\[3\] 0.045013f
C11927 _413_/a_796_472# vdd 0.001569f
C11928 net76 net59 3.439686f
C11929 cal_count\[3\] FILLER_0_11_78/a_36_472# 0.031399f
C11930 ctlp[1] FILLER_0_24_274/a_1020_375# 0.004803f
C11931 _430_/a_36_151# _136_ 0.02044f
C11932 FILLER_0_3_172/a_484_472# net22 0.012284f
C11933 _086_ FILLER_0_4_177/a_36_472# 0.001464f
C11934 _427_/a_36_151# _043_ 0.002267f
C11935 _438_/a_2665_112# FILLER_0_19_111/a_124_375# 0.006271f
C11936 _094_ _418_/a_2560_156# 0.011088f
C11937 net16 trim_mask\[1\] 0.007065f
C11938 FILLER_0_16_107/a_124_375# vss 0.002683f
C11939 _057_ state\[1\] 0.284428f
C11940 net5 vss 0.326032f
C11941 _141_ net23 0.782974f
C11942 _422_/a_796_472# mask\[7\] 0.001755f
C11943 output16/a_224_472# net16 0.054603f
C11944 output13/a_224_472# net22 0.022308f
C11945 result[6] _420_/a_796_472# 0.002296f
C11946 net44 _054_ 0.003562f
C11947 _301_/a_36_472# net25 0.003165f
C11948 net80 vdd 1.045288f
C11949 _076_ FILLER_0_6_231/a_572_375# 0.001647f
C11950 net23 _348_/a_49_472# 0.0037f
C11951 output18/a_224_472# net33 0.135766f
C11952 _091_ FILLER_0_17_218/a_36_472# 0.066133f
C11953 FILLER_0_6_177/a_36_472# net47 0.011891f
C11954 FILLER_0_5_117/a_124_375# _158_ 0.001068f
C11955 _256_/a_2124_68# _070_ 0.002444f
C11956 net36 net23 0.028202f
C11957 FILLER_0_11_78/a_572_375# _389_/a_36_148# 0.021545f
C11958 _360_/a_36_160# _160_ 0.052885f
C11959 _321_/a_3662_472# _176_ 0.002006f
C11960 _150_ _356_/a_36_472# 0.007271f
C11961 _164_ _381_/a_36_472# 0.007224f
C11962 FILLER_0_16_37/a_36_472# cal_count\[2\] 0.008691f
C11963 _053_ FILLER_0_6_47/a_2812_375# 0.003818f
C11964 _250_/a_36_68# state\[1\] 0.103037f
C11965 _093_ FILLER_0_17_72/a_1828_472# 0.053526f
C11966 FILLER_0_5_181/a_124_375# net22 0.00205f
C11967 _408_/a_728_93# _043_ 0.029183f
C11968 _436_/a_2560_156# FILLER_0_22_128/a_124_375# 0.001178f
C11969 _436_/a_2665_112# FILLER_0_22_128/a_572_375# 0.001092f
C11970 FILLER_0_15_235/a_484_472# vss 0.003614f
C11971 FILLER_0_15_235/a_572_375# mask\[1\] 0.013718f
C11972 FILLER_0_13_142/a_1380_472# _043_ 0.011974f
C11973 FILLER_0_20_177/a_1380_472# vss 0.004504f
C11974 net38 FILLER_0_20_15/a_124_375# 0.012947f
C11975 mask\[5\] _292_/a_36_160# 0.007486f
C11976 FILLER_0_16_107/a_572_375# FILLER_0_18_107/a_484_472# 0.001512f
C11977 net58 FILLER_0_9_290/a_36_472# 0.005553f
C11978 fanout72/a_36_113# net74 0.02894f
C11979 FILLER_0_5_198/a_124_375# net59 0.00174f
C11980 _431_/a_36_151# FILLER_0_18_107/a_1828_472# 0.001221f
C11981 _428_/a_36_151# net70 0.040167f
C11982 net44 vss 0.477283f
C11983 cal_itt\[1\] FILLER_0_3_221/a_1380_472# 0.004939f
C11984 _192_/a_67_603# mask\[1\] 0.020097f
C11985 mask\[1\] vdd 0.741266f
C11986 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1380_472# 0.013276f
C11987 fanout52/a_36_160# trim_val\[4\] 0.019286f
C11988 FILLER_0_10_78/a_36_472# vdd 0.001865f
C11989 output29/a_224_472# _094_ 0.006731f
C11990 FILLER_0_20_169/a_36_472# _339_/a_36_160# 0.001448f
C11991 net36 FILLER_0_15_212/a_484_472# 0.007742f
C11992 net76 _122_ 0.028025f
C11993 FILLER_0_2_177/a_124_375# net59 0.005212f
C11994 FILLER_0_11_142/a_124_375# vdd 0.010672f
C11995 FILLER_0_17_56/a_36_472# _183_ 0.056523f
C11996 _429_/a_2665_112# FILLER_0_15_212/a_1468_375# 0.010688f
C11997 cal_count\[3\] net51 0.042416f
C11998 FILLER_0_20_15/a_1380_472# vss 0.003678f
C11999 _322_/a_124_24# _129_ 0.017754f
C12000 _092_ FILLER_0_17_218/a_572_375# 0.006125f
C12001 FILLER_0_18_107/a_1916_375# vdd 0.018831f
C12002 FILLER_0_10_78/a_1020_375# _120_ 0.003403f
C12003 _098_ FILLER_0_21_150/a_36_472# 0.002964f
C12004 FILLER_0_12_50/a_36_472# cal_count\[0\] 0.001857f
C12005 _004_ fanout79/a_36_160# 0.048599f
C12006 net24 FILLER_0_22_86/a_1020_375# 0.022658f
C12007 _422_/a_2248_156# vdd 0.005833f
C12008 FILLER_0_7_104/a_124_375# vdd 0.031505f
C12009 net41 net26 0.057852f
C12010 net79 FILLER_0_12_220/a_36_472# 0.005464f
C12011 _441_/a_2665_112# vss 0.005169f
C12012 _074_ _375_/a_960_497# 0.004175f
C12013 net55 _424_/a_2665_112# 0.056555f
C12014 _149_ net71 0.827628f
C12015 mask\[4\] FILLER_0_18_177/a_1468_375# 0.01587f
C12016 mask\[0\] net22 0.054097f
C12017 mask\[3\] FILLER_0_18_177/a_572_375# 0.002924f
C12018 _447_/a_796_472# net68 0.001593f
C12019 _447_/a_448_472# _036_ 0.015378f
C12020 FILLER_0_17_226/a_124_375# _106_ 0.061857f
C12021 result[9] net29 0.001272f
C12022 FILLER_0_21_28/a_124_375# FILLER_0_19_28/a_36_472# 0.001512f
C12023 FILLER_0_17_56/a_572_375# FILLER_0_15_59/a_36_472# 0.001188f
C12024 _115_ FILLER_0_11_78/a_572_375# 0.034089f
C12025 input2/a_36_113# vdd 0.096633f
C12026 _122_ FILLER_0_5_198/a_124_375# 0.001352f
C12027 FILLER_0_19_47/a_36_472# net26 0.050805f
C12028 net47 _452_/a_448_472# 0.005335f
C12029 net20 _081_ 0.024512f
C12030 _208_/a_36_160# FILLER_0_22_128/a_2812_375# 0.026361f
C12031 _131_ FILLER_0_17_104/a_484_472# 0.003483f
C12032 _086_ _315_/a_36_68# 0.003329f
C12033 net63 net21 0.278824f
C12034 _441_/a_36_151# net66 0.057618f
C12035 _413_/a_36_151# net65 0.033028f
C12036 FILLER_0_9_142/a_36_472# net23 0.001099f
C12037 net15 _423_/a_1000_472# 0.001786f
C12038 _437_/a_448_472# vdd 0.010432f
C12039 _437_/a_36_151# vss 0.006865f
C12040 _093_ FILLER_0_18_139/a_124_375# 0.008393f
C12041 output9/a_224_472# input4/a_36_68# 0.009732f
C12042 _411_/a_1204_472# net8 0.001768f
C12043 net31 _046_ 0.008368f
C12044 _449_/a_1000_472# _038_ 0.021492f
C12045 FILLER_0_3_172/a_36_472# vss 0.001848f
C12046 FILLER_0_3_172/a_484_472# vdd 0.007258f
C12047 _106_ _276_/a_36_160# 0.009097f
C12048 net63 FILLER_0_19_171/a_932_472# 0.00128f
C12049 FILLER_0_5_198/a_572_375# net21 0.023563f
C12050 FILLER_0_21_125/a_572_375# _433_/a_36_151# 0.059049f
C12051 FILLER_0_11_109/a_36_472# FILLER_0_10_107/a_124_375# 0.001684f
C12052 output13/a_224_472# vdd 0.045929f
C12053 net16 _444_/a_2665_112# 0.011295f
C12054 _144_ _348_/a_257_69# 0.001978f
C12055 fanout71/a_36_113# mask\[9\] 0.044939f
C12056 _052_ FILLER_0_18_37/a_1468_375# 0.001585f
C12057 FILLER_0_8_138/a_124_375# _129_ 0.006506f
C12058 FILLER_0_21_286/a_484_472# _420_/a_36_151# 0.027236f
C12059 net20 net65 0.335083f
C12060 FILLER_0_10_28/a_124_375# net6 0.007948f
C12061 cal_count\[3\] _228_/a_36_68# 0.01871f
C12062 _128_ net23 0.041791f
C12063 _147_ _049_ 0.001131f
C12064 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1380_472# 0.003468f
C12065 _017_ net74 0.041246f
C12066 net64 _043_ 0.004021f
C12067 output34/a_224_472# vdd 0.094191f
C12068 vdd _416_/a_2560_156# 0.00165f
C12069 vss _416_/a_2665_112# 0.002676f
C12070 _432_/a_2248_156# _091_ 0.007123f
C12071 _422_/a_2560_156# _108_ 0.008253f
C12072 FILLER_0_5_181/a_124_375# vdd 0.009553f
C12073 cal_itt\[3\] _074_ 0.584958f
C12074 vdd output6/a_224_472# 0.009312f
C12075 FILLER_0_5_88/a_36_472# vss 0.005793f
C12076 _069_ net21 0.032615f
C12077 FILLER_0_22_177/a_36_472# mask\[6\] 0.006882f
C12078 net35 FILLER_0_22_177/a_1468_375# 0.048182f
C12079 _093_ FILLER_0_18_76/a_572_375# 0.025143f
C12080 net73 _136_ 0.050578f
C12081 mask\[9\] FILLER_0_18_76/a_124_375# 0.004592f
C12082 _008_ _102_ 0.027578f
C12083 net75 valid 0.002077f
C12084 cal_itt\[3\] _076_ 0.002726f
C12085 net76 FILLER_0_5_206/a_124_375# 0.006974f
C12086 _176_ FILLER_0_11_78/a_484_472# 0.008724f
C12087 _171_ vdd 0.038202f
C12088 _430_/a_2665_112# mask\[1\] 0.004574f
C12089 FILLER_0_17_200/a_484_472# _430_/a_36_151# 0.001723f
C12090 FILLER_0_13_206/a_124_375# net79 0.009649f
C12091 net72 _131_ 0.186396f
C12092 _280_/a_224_472# _097_ 0.007508f
C12093 _365_/a_36_68# net14 0.017522f
C12094 FILLER_0_4_49/a_484_472# net49 0.006499f
C12095 output48/a_224_472# vdd 0.038342f
C12096 net75 FILLER_0_8_247/a_36_472# 0.002992f
C12097 net54 FILLER_0_18_139/a_124_375# 0.002807f
C12098 FILLER_0_7_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001723f
C12099 _004_ FILLER_0_10_247/a_124_375# 0.004573f
C12100 result[7] _419_/a_1000_472# 0.015362f
C12101 _413_/a_2665_112# vdd 0.02286f
C12102 _025_ FILLER_0_22_107/a_572_375# 0.090334f
C12103 _148_ FILLER_0_22_107/a_484_472# 0.004761f
C12104 fanout56/a_36_113# _095_ 0.004331f
C12105 fanout73/a_36_113# net36 0.01199f
C12106 result[9] net60 0.251903f
C12107 mask\[0\] vdd 0.181371f
C12108 FILLER_0_14_107/a_1380_472# _043_ 0.001641f
C12109 FILLER_0_13_100/a_36_472# vdd 0.021826f
C12110 FILLER_0_16_57/a_124_375# FILLER_0_18_53/a_484_472# 0.001512f
C12111 FILLER_0_13_100/a_124_375# vss 0.00513f
C12112 FILLER_0_14_50/a_36_472# FILLER_0_12_50/a_124_375# 0.0027f
C12113 _051_ vss 0.050185f
C12114 _093_ FILLER_0_18_209/a_124_375# 0.00333f
C12115 _119_ _120_ 0.036534f
C12116 FILLER_0_17_200/a_572_375# net22 0.047331f
C12117 _033_ _160_ 0.020281f
C12118 _136_ FILLER_0_14_99/a_36_472# 0.01535f
C12119 _105_ mask\[4\] 0.025209f
C12120 _126_ _018_ 0.001243f
C12121 ctlp[3] net61 0.007397f
C12122 net63 mask\[7\] 0.069252f
C12123 net73 fanout70/a_36_113# 0.21211f
C12124 trim_val\[2\] net68 0.010894f
C12125 _031_ trim_mask\[3\] 0.016747f
C12126 _183_ FILLER_0_18_53/a_36_472# 0.007412f
C12127 _179_ vdd 0.049022f
C12128 _061_ FILLER_0_8_156/a_572_375# 0.023346f
C12129 _255_/a_224_552# _161_ 0.025424f
C12130 _013_ _424_/a_1000_472# 0.037585f
C12131 _420_/a_1000_472# vss 0.002146f
C12132 FILLER_0_20_107/a_124_375# net71 0.03452f
C12133 _095_ FILLER_0_14_107/a_484_472# 0.014431f
C12134 net17 net43 0.144179f
C12135 _072_ _246_/a_36_68# 0.064797f
C12136 FILLER_0_9_223/a_572_375# calibrate 0.002082f
C12137 _435_/a_2665_112# net21 0.067461f
C12138 net4 FILLER_0_12_220/a_484_472# 0.022264f
C12139 _394_/a_1336_472# FILLER_0_13_72/a_124_375# 0.001597f
C12140 _141_ FILLER_0_19_155/a_484_472# 0.015625f
C12141 net3 vdd 0.118499f
C12142 net57 net36 0.087967f
C12143 FILLER_0_10_256/a_124_375# net28 0.034928f
C12144 FILLER_0_16_89/a_932_472# FILLER_0_17_72/a_2812_375# 0.001723f
C12145 _089_ FILLER_0_3_172/a_2276_472# 0.001522f
C12146 fanout65/a_36_113# net64 0.002858f
C12147 net63 net80 0.337396f
C12148 ctlp[4] result[8] 0.151286f
C12149 _242_/a_36_160# vdd 0.007995f
C12150 cal_itt\[3\] FILLER_0_5_164/a_484_472# 0.001518f
C12151 net61 net78 1.588656f
C12152 _360_/a_36_160# _133_ 0.001878f
C12153 _444_/a_796_472# net67 0.006859f
C12154 _113_ FILLER_0_12_196/a_124_375# 0.001597f
C12155 _323_/a_36_113# net4 0.005657f
C12156 _090_ FILLER_0_12_196/a_36_472# 0.002321f
C12157 net52 _443_/a_796_472# 0.004334f
C12158 FILLER_0_7_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001723f
C12159 _446_/a_2248_156# net49 0.006196f
C12160 net44 _450_/a_1040_527# 0.002267f
C12161 _099_ FILLER_0_15_235/a_572_375# 0.001327f
C12162 net67 FILLER_0_8_24/a_36_472# 0.001252f
C12163 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_36_472# 0.002296f
C12164 net35 _436_/a_448_472# 0.012374f
C12165 _174_ cal_count\[2\] 0.004821f
C12166 FILLER_0_3_78/a_572_375# _160_ 0.003506f
C12167 net48 _251_/a_468_472# 0.002731f
C12168 _322_/a_848_380# _076_ 0.006699f
C12169 net52 _448_/a_2248_156# 0.002555f
C12170 _233_/a_36_160# FILLER_0_6_37/a_36_472# 0.012692f
C12171 FILLER_0_15_212/a_124_375# vdd -0.004549f
C12172 _132_ _127_ 0.112364f
C12173 _431_/a_448_472# _020_ 0.05255f
C12174 _099_ vdd 0.326559f
C12175 output11/a_224_472# FILLER_0_0_232/a_124_375# 0.00515f
C12176 FILLER_0_4_107/a_572_375# _151_ 0.00162f
C12177 FILLER_0_20_177/a_1468_375# _434_/a_36_151# 0.001822f
C12178 FILLER_0_16_154/a_1468_375# vss 0.002071f
C12179 FILLER_0_16_154/a_36_472# vdd 0.00225f
C12180 FILLER_0_16_73/a_484_472# FILLER_0_17_72/a_572_375# 0.001723f
C12181 FILLER_0_4_99/a_36_472# vdd 0.094733f
C12182 FILLER_0_4_99/a_124_375# vss 0.017518f
C12183 _411_/a_2560_156# net8 0.013106f
C12184 FILLER_0_13_65/a_124_375# vdd 0.011301f
C12185 net63 mask\[1\] 0.120872f
C12186 net73 net53 0.094507f
C12187 output11/a_224_472# net11 0.003448f
C12188 cal_itt\[3\] _081_ 0.03503f
C12189 net64 FILLER_0_12_236/a_124_375# 0.043517f
C12190 output37/a_224_472# fanout59/a_36_160# 0.021845f
C12191 _055_ vss 0.365503f
C12192 trim_mask\[1\] FILLER_0_6_47/a_124_375# 0.005902f
C12193 _274_/a_2960_68# _070_ 0.001963f
C12194 FILLER_0_19_111/a_124_375# vdd 0.005128f
C12195 _421_/a_796_472# _010_ 0.037434f
C12196 FILLER_0_5_198/a_484_472# vss 0.001338f
C12197 FILLER_0_22_86/a_932_472# net14 0.020589f
C12198 _419_/a_2248_156# vdd 0.040646f
C12199 _144_ _433_/a_796_472# 0.008448f
C12200 _386_/a_848_380# net37 0.006086f
C12201 _414_/a_1308_423# cal_itt\[3\] 0.044184f
C12202 output25/a_224_472# mask\[8\] 0.015742f
C12203 FILLER_0_18_107/a_572_375# FILLER_0_19_111/a_124_375# 0.058411f
C12204 _086_ FILLER_0_6_177/a_484_472# 0.017841f
C12205 FILLER_0_4_197/a_124_375# net22 0.00145f
C12206 net19 _420_/a_2665_112# 0.012322f
C12207 FILLER_0_16_89/a_36_472# _093_ 0.001338f
C12208 FILLER_0_12_136/a_36_472# _127_ 0.023927f
C12209 _432_/a_1308_423# _093_ 0.016365f
C12210 _232_/a_67_603# FILLER_0_5_54/a_36_472# 0.025312f
C12211 mask\[7\] FILLER_0_22_177/a_124_375# 0.001315f
C12212 net76 FILLER_0_3_172/a_932_472# 0.005391f
C12213 fanout53/a_36_160# _137_ 0.001852f
C12214 _053_ FILLER_0_7_59/a_124_375# 0.015298f
C12215 net50 _029_ 0.025102f
C12216 mask\[8\] _354_/a_257_69# 0.003809f
C12217 FILLER_0_17_200/a_572_375# vdd 0.006861f
C12218 net75 _253_/a_36_68# 0.047906f
C12219 _079_ _260_/a_244_472# 0.00325f
C12220 _093_ FILLER_0_17_142/a_36_472# 0.011974f
C12221 _069_ mask\[1\] 0.029447f
C12222 _126_ vss 0.399848f
C12223 net53 FILLER_0_14_99/a_36_472# 0.004153f
C12224 _414_/a_1204_472# cal_itt\[3\] 0.052432f
C12225 FILLER_0_13_212/a_1468_375# net79 0.009597f
C12226 FILLER_0_24_130/a_124_375# _050_ 0.007643f
C12227 net62 FILLER_0_13_212/a_36_472# 0.015187f
C12228 FILLER_0_4_91/a_572_375# _156_ 0.004958f
C12229 _327_/a_36_472# _428_/a_2248_156# 0.001757f
C12230 _069_ FILLER_0_11_142/a_124_375# 0.030279f
C12231 FILLER_0_7_72/a_3172_472# net14 0.046751f
C12232 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_36_472# 0.026657f
C12233 net16 _424_/a_36_151# 0.002969f
C12234 FILLER_0_3_204/a_124_375# _088_ 0.00269f
C12235 net4 FILLER_0_3_221/a_36_472# 0.010517f
C12236 mask\[5\] FILLER_0_18_177/a_124_375# 0.002726f
C12237 _431_/a_36_151# _132_ 0.051016f
C12238 net16 net66 0.030521f
C12239 cal_count\[3\] net47 0.043032f
C12240 net80 FILLER_0_22_177/a_124_375# 0.013214f
C12241 mask\[7\] _435_/a_2665_112# 0.030393f
C12242 net69 FILLER_0_2_101/a_124_375# 0.015032f
C12243 net41 _033_ 0.033812f
C12244 _394_/a_1936_472# cal_count\[1\] 0.008364f
C12245 ctln[4] _411_/a_36_151# 0.0022f
C12246 net76 FILLER_0_5_181/a_36_472# 0.014784f
C12247 net18 net33 0.001671f
C12248 net57 _128_ 0.040656f
C12249 FILLER_0_1_212/a_124_375# vss 0.011796f
C12250 FILLER_0_1_212/a_36_472# vdd 0.10765f
C12251 net16 _067_ 0.039705f
C12252 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1380_472# 0.013277f
C12253 _450_/a_36_151# net6 0.035997f
C12254 _450_/a_1353_112# output6/a_224_472# 0.008732f
C12255 _059_ net47 0.00606f
C12256 _413_/a_1308_423# net82 0.003079f
C12257 _174_ _043_ 0.964645f
C12258 _176_ _067_ 0.046599f
C12259 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_572_375# 0.001597f
C12260 _412_/a_1204_472# net59 0.001824f
C12261 FILLER_0_12_220/a_1020_375# vdd -0.014642f
C12262 FILLER_0_12_220/a_572_375# vss 0.007775f
C12263 _053_ _070_ 2.345795f
C12264 _132_ _345_/a_36_160# 0.078243f
C12265 _426_/a_1204_472# calibrate 0.00182f
C12266 FILLER_0_18_139/a_932_472# vss 0.041568f
C12267 _137_ _098_ 0.07262f
C12268 FILLER_0_18_139/a_1380_472# vdd 0.005855f
C12269 _030_ _157_ 0.011014f
C12270 _270_/a_36_472# net22 0.002857f
C12271 _053_ FILLER_0_7_146/a_36_472# 0.001014f
C12272 _187_ net16 0.161791f
C12273 output39/a_224_472# _445_/a_36_151# 0.11862f
C12274 _093_ FILLER_0_18_107/a_1828_472# 0.001872f
C12275 FILLER_0_5_72/a_572_375# _029_ 0.010208f
C12276 FILLER_0_22_177/a_1468_375# vdd -0.007187f
C12277 FILLER_0_15_282/a_484_472# result[3] 0.026996f
C12278 net19 _419_/a_2560_156# 0.003213f
C12279 _093_ _102_ 0.008937f
C12280 _447_/a_2665_112# _030_ 0.001226f
C12281 FILLER_0_24_96/a_36_472# output25/a_224_472# 0.010475f
C12282 _426_/a_1000_472# net64 0.008796f
C12283 _004_ net27 0.080285f
C12284 FILLER_0_21_133/a_36_472# mask\[7\] 0.003404f
C12285 mask\[2\] FILLER_0_16_154/a_124_375# 0.087247f
C12286 FILLER_0_4_107/a_1020_375# _160_ 0.015684f
C12287 net18 FILLER_0_17_282/a_124_375# 0.048177f
C12288 _155_ net50 0.012085f
C12289 FILLER_0_4_213/a_124_375# vdd 0.009037f
C12290 _255_/a_224_552# _056_ 0.033615f
C12291 FILLER_0_17_282/a_36_472# net30 0.001189f
C12292 FILLER_0_1_192/a_36_472# net59 0.082738f
C12293 _136_ _438_/a_36_151# 0.030558f
C12294 net31 _006_ 0.307613f
C12295 FILLER_0_17_72/a_572_375# _131_ 0.006224f
C12296 _204_/a_67_603# vss 0.010366f
C12297 output10/a_224_472# net58 0.025878f
C12298 _081_ _265_/a_244_68# 0.03338f
C12299 fanout62/a_36_160# net62 0.02201f
C12300 net38 _444_/a_1288_156# 0.001147f
C12301 _449_/a_1308_423# vss 0.027539f
C12302 FILLER_0_21_286/a_572_375# net77 0.044323f
C12303 _153_ _365_/a_36_68# 0.056496f
C12304 net20 FILLER_0_7_233/a_36_472# 0.035074f
C12305 _130_ _120_ 0.014675f
C12306 net70 FILLER_0_14_123/a_124_375# 0.032077f
C12307 result[6] _421_/a_1308_423# 0.023269f
C12308 net31 _103_ 0.227588f
C12309 FILLER_0_4_197/a_124_375# vdd 0.011327f
C12310 output37/a_224_472# net5 0.072504f
C12311 net74 cal_count\[3\] 0.040777f
C12312 result[1] vss 0.311464f
C12313 _431_/a_2248_156# vss 0.041929f
C12314 mask\[0\] _283_/a_36_472# 0.004645f
C12315 net28 mask\[1\] 0.572459f
C12316 _443_/a_2665_112# trim_mask\[4\] 0.013708f
C12317 _026_ _437_/a_1308_423# 0.018479f
C12318 _149_ _437_/a_1000_472# 0.019115f
C12319 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_932_472# 0.001723f
C12320 net33 _048_ 0.017633f
C12321 net74 _059_ 0.004133f
C12322 _451_/a_448_472# _040_ 0.026819f
C12323 net15 FILLER_0_17_64/a_36_472# 0.015524f
C12324 _122_ FILLER_0_6_231/a_36_472# 0.015997f
C12325 _129_ _120_ 0.017802f
C12326 FILLER_0_7_162/a_124_375# net47 0.030995f
C12327 FILLER_0_14_263/a_124_375# net30 0.016642f
C12328 _255_/a_224_552# _068_ 0.002412f
C12329 _016_ _428_/a_2560_156# 0.003934f
C12330 _402_/a_56_567# vdd 0.014708f
C12331 _178_ _402_/a_728_93# 0.050963f
C12332 _114_ net23 0.029535f
C12333 net41 _446_/a_36_151# 0.143017f
C12334 _083_ _082_ 0.018442f
C12335 _141_ _340_/a_36_160# 0.00584f
C12336 output18/a_224_472# vdd -0.01545f
C12337 net82 _083_ 0.010347f
C12338 net55 _182_ 0.012838f
C12339 net50 FILLER_0_8_24/a_484_472# 0.059367f
C12340 mask\[4\] FILLER_0_19_171/a_1020_375# 0.006236f
C12341 _340_/a_36_160# _348_/a_49_472# 0.001528f
C12342 FILLER_0_12_236/a_484_472# vss 0.002739f
C12343 _432_/a_36_151# _137_ 0.051293f
C12344 _137_ FILLER_0_15_180/a_124_375# 0.003108f
C12345 FILLER_0_14_91/a_484_472# vss 0.003257f
C12346 FILLER_0_7_104/a_932_472# _062_ 0.001184f
C12347 net50 _163_ 0.068547f
C12348 _442_/a_1000_472# _031_ 0.004174f
C12349 FILLER_0_21_28/a_2276_472# vdd 0.002733f
C12350 FILLER_0_21_28/a_1828_472# vss -0.001894f
C12351 _436_/a_448_472# vdd 0.038494f
C12352 FILLER_0_3_221/a_124_375# vss 0.034009f
C12353 net75 _079_ 0.071974f
C12354 _423_/a_1000_472# _012_ 0.013415f
C12355 _053_ trim_val\[1\] 0.00385f
C12356 FILLER_0_17_282/a_36_472# _417_/a_36_151# 0.001723f
C12357 FILLER_0_1_192/a_124_375# net11 0.003537f
C12358 trim_mask\[3\] _157_ 0.052956f
C12359 net36 _438_/a_1308_423# 0.012976f
C12360 _069_ mask\[0\] 0.040599f
C12361 output15/a_224_472# net50 0.00515f
C12362 ctln[8] fanout50/a_36_160# 0.004838f
C12363 _000_ vdd 0.215988f
C12364 net15 net52 0.166073f
C12365 net52 FILLER_0_11_78/a_36_472# 0.005678f
C12366 _439_/a_36_151# vss 0.032466f
C12367 _439_/a_448_472# vdd 0.006996f
C12368 _114_ FILLER_0_11_109/a_124_375# 0.009676f
C12369 _270_/a_36_472# vdd 0.09815f
C12370 _283_/a_36_472# _099_ 0.004667f
C12371 FILLER_0_17_200/a_36_472# _093_ 0.005101f
C12372 output39/a_224_472# _063_ 0.001019f
C12373 net39 _233_/a_36_160# 0.017979f
C12374 FILLER_0_8_239/a_124_375# _123_ 0.001286f
C12375 _071_ _055_ 0.002641f
C12376 net36 _451_/a_2449_156# 0.016229f
C12377 FILLER_0_17_200/a_484_472# mask\[3\] 0.014805f
C12378 _427_/a_2248_156# net23 0.033973f
C12379 FILLER_0_21_28/a_2364_375# _424_/a_36_151# 0.059049f
C12380 net63 FILLER_0_15_212/a_124_375# 0.001597f
C12381 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_124_375# 0.003228f
C12382 _095_ FILLER_0_13_100/a_124_375# 0.001989f
C12383 state\[1\] vss 0.294171f
C12384 net15 net49 0.057277f
C12385 FILLER_0_14_50/a_36_472# _180_ 0.153222f
C12386 FILLER_0_9_28/a_124_375# vdd -0.004893f
C12387 _176_ net23 0.036283f
C12388 mask\[5\] _143_ 0.032539f
C12389 _007_ vss 0.017377f
C12390 _321_/a_786_69# net23 0.001073f
C12391 _449_/a_2665_112# cal_count\[3\] 0.001422f
C12392 FILLER_0_12_136/a_124_375# cal_count\[3\] 0.005006f
C12393 _239_/a_36_160# _447_/a_36_151# 0.137659f
C12394 result[1] _416_/a_2248_156# 0.001888f
C12395 FILLER_0_0_266/a_124_375# vss 0.007654f
C12396 FILLER_0_0_266/a_36_472# vdd 0.05043f
C12397 _326_/a_36_160# FILLER_0_9_105/a_572_375# 0.005489f
C12398 output23/a_224_472# vss 0.075684f
C12399 _112_ _425_/a_1000_472# 0.001973f
C12400 FILLER_0_6_239/a_124_375# net37 0.001989f
C12401 FILLER_0_16_57/a_36_472# _176_ 0.075537f
C12402 result[7] _421_/a_1308_423# 0.022204f
C12403 net53 _451_/a_3129_107# 0.002806f
C12404 _126_ _071_ 0.090032f
C12405 _141_ _348_/a_49_472# 0.037821f
C12406 FILLER_0_4_197/a_36_472# net21 0.011079f
C12407 output32/a_224_472# _006_ 0.001009f
C12408 net75 cal_itt\[1\] 0.704169f
C12409 net62 _285_/a_36_472# 0.001288f
C12410 net18 FILLER_0_11_282/a_36_472# 0.048657f
C12411 _354_/a_49_472# vdd -0.001073f
C12412 _069_ FILLER_0_15_212/a_124_375# 0.039975f
C12413 net52 net51 0.091698f
C12414 _370_/a_692_472# _081_ 0.00129f
C12415 _370_/a_848_380# _152_ 0.031499f
C12416 trimb[4] FILLER_0_15_2/a_36_472# 0.006046f
C12417 net19 net37 0.030961f
C12418 FILLER_0_21_125/a_36_472# net54 0.016672f
C12419 output32/a_224_472# _103_ 0.090957f
C12420 ctln[2] vss 0.256543f
C12421 FILLER_0_17_200/a_572_375# net63 0.007512f
C12422 _140_ mask\[7\] 0.064343f
C12423 net60 _418_/a_1000_472# 0.007557f
C12424 _119_ _125_ 0.11554f
C12425 net29 _044_ 0.01495f
C12426 net39 net49 0.158007f
C12427 _062_ net14 0.003317f
C12428 mask\[4\] _433_/a_2248_156# 0.001082f
C12429 _413_/a_448_472# net65 0.044062f
C12430 _256_/a_36_68# net22 0.019035f
C12431 net24 FILLER_0_23_88/a_36_472# 0.006289f
C12432 net82 _425_/a_36_151# 0.002959f
C12433 _426_/a_2665_112# vss 0.006288f
C12434 _277_/a_36_160# _103_ 0.032112f
C12435 _095_ _055_ 0.002933f
C12436 FILLER_0_10_78/a_124_375# FILLER_0_11_78/a_124_375# 0.05841f
C12437 FILLER_0_8_127/a_124_375# _058_ 0.007791f
C12438 result[0] FILLER_0_9_282/a_124_375# 0.00283f
C12439 net79 _417_/a_796_472# 0.001042f
C12440 FILLER_0_24_96/a_124_375# vss 0.017357f
C12441 net29 _287_/a_244_68# 0.001262f
C12442 net50 FILLER_0_4_91/a_36_472# 0.058499f
C12443 net62 _417_/a_1000_472# 0.005762f
C12444 net32 _419_/a_36_151# 0.006506f
C12445 net80 _140_ 0.188514f
C12446 _326_/a_36_160# _125_ 0.050008f
C12447 _086_ _058_ 0.054155f
C12448 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_36_472# 0.086904f
C12449 _151_ vdd 0.157764f
C12450 ctln[8] net14 0.001447f
C12451 net81 _018_ 0.081888f
C12452 output12/a_224_472# FILLER_0_0_198/a_36_472# 0.023414f
C12453 _120_ _453_/a_36_151# 0.001848f
C12454 FILLER_0_6_47/a_36_472# vdd 0.090192f
C12455 FILLER_0_6_47/a_3260_375# vss 0.061766f
C12456 net15 FILLER_0_15_72/a_572_375# 0.002741f
C12457 FILLER_0_4_197/a_1380_472# FILLER_0_4_213/a_36_472# 0.013277f
C12458 mask\[4\] FILLER_0_20_177/a_36_472# 0.001215f
C12459 FILLER_0_13_290/a_36_472# result[3] 0.001069f
C12460 fanout58/a_36_160# vdd 0.101571f
C12461 mask\[8\] FILLER_0_22_107/a_124_375# 0.015331f
C12462 trim[4] _236_/a_36_160# 0.004514f
C12463 FILLER_0_17_200/a_572_375# _069_ 0.011239f
C12464 FILLER_0_16_255/a_124_375# _006_ 0.02007f
C12465 FILLER_0_11_135/a_124_375# _120_ 0.017316f
C12466 FILLER_0_16_73/a_484_472# vdd 0.003462f
C12467 net63 FILLER_0_22_177/a_1468_375# 0.005028f
C12468 _105_ _201_/a_67_603# 0.003335f
C12469 cal_count\[2\] _402_/a_244_567# 0.004411f
C12470 _089_ _079_ 0.126206f
C12471 output22/a_224_472# _024_ 0.029795f
C12472 net36 FILLER_0_15_228/a_36_472# 0.008225f
C12473 _402_/a_728_93# _401_/a_36_68# 0.002178f
C12474 fanout75/a_36_113# vdd 0.028614f
C12475 cal_itt\[3\] _163_ 0.021146f
C12476 _077_ net48 0.142015f
C12477 net70 _017_ 0.015488f
C12478 FILLER_0_13_212/a_572_375# vdd 0.001551f
C12479 FILLER_0_13_212/a_124_375# vss 0.007116f
C12480 _429_/a_2248_156# FILLER_0_15_228/a_124_375# 0.030666f
C12481 FILLER_0_6_90/a_484_472# net14 0.014785f
C12482 _050_ _436_/a_2560_156# 0.01099f
C12483 _131_ FILLER_0_14_107/a_1468_375# 0.051201f
C12484 trim[0] net66 0.376153f
C12485 FILLER_0_12_136/a_572_375# _114_ 0.006974f
C12486 FILLER_0_11_101/a_572_375# _120_ 0.006382f
C12487 FILLER_0_12_220/a_1468_375# _043_ 0.002509f
C12488 _421_/a_1000_472# vdd 0.006281f
C12489 FILLER_0_20_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001543f
C12490 FILLER_0_10_214/a_124_375# vdd 0.018944f
C12491 _446_/a_448_472# net17 0.026011f
C12492 result[9] FILLER_0_24_274/a_484_472# 0.003507f
C12493 _068_ _120_ 0.447243f
C12494 net57 _443_/a_2248_156# 0.001117f
C12495 FILLER_0_1_98/a_124_375# net14 0.049552f
C12496 FILLER_0_8_37/a_36_472# _054_ 0.015053f
C12497 FILLER_0_13_65/a_124_375# _449_/a_36_151# 0.059049f
C12498 net62 _101_ 0.023932f
C12499 _412_/a_796_472# net1 0.002922f
C12500 _415_/a_1204_472# vdd 0.00108f
C12501 result[8] FILLER_0_24_274/a_36_472# 0.005458f
C12502 _394_/a_1936_472# _175_ 0.017848f
C12503 vdd FILLER_0_21_60/a_572_375# 0.022291f
C12504 vss FILLER_0_21_60/a_124_375# 0.003723f
C12505 net26 FILLER_0_23_44/a_36_472# 0.013977f
C12506 net55 FILLER_0_17_72/a_1468_375# 0.014449f
C12507 _422_/a_36_151# _421_/a_2665_112# 0.001725f
C12508 _431_/a_2665_112# FILLER_0_15_150/a_36_472# 0.035266f
C12509 fanout53/a_36_160# fanout56/a_36_113# 0.001636f
C12510 FILLER_0_2_111/a_124_375# vdd 0.024756f
C12511 _429_/a_36_151# net22 0.020582f
C12512 _093_ FILLER_0_17_104/a_1468_375# 0.010965f
C12513 net41 _444_/a_36_151# 0.013142f
C12514 output47/a_224_472# _452_/a_3129_107# 0.018181f
C12515 output12/a_224_472# net11 0.009336f
C12516 _413_/a_1308_423# net21 0.065716f
C12517 _114_ net57 0.22998f
C12518 _440_/a_36_151# vdd 0.117768f
C12519 net34 _295_/a_36_472# 0.032003f
C12520 FILLER_0_9_28/a_36_472# net40 0.020589f
C12521 _008_ _198_/a_67_603# 0.012332f
C12522 FILLER_0_16_57/a_1380_472# net15 0.017841f
C12523 fanout51/a_36_113# _120_ 0.014349f
C12524 cal en 0.482495f
C12525 FILLER_0_8_37/a_484_472# vdd 0.009603f
C12526 _021_ mask\[3\] 0.036781f
C12527 _132_ _093_ 0.105039f
C12528 net66 _030_ 0.087608f
C12529 _078_ net59 0.168928f
C12530 state\[0\] _060_ 0.047136f
C12531 _267_/a_36_472# net23 0.001178f
C12532 fanout74/a_36_113# _443_/a_36_151# 0.032681f
C12533 FILLER_0_21_28/a_2812_375# _012_ 0.016736f
C12534 FILLER_0_5_72/a_484_472# vss 0.003738f
C12535 FILLER_0_5_72/a_932_472# vdd 0.002735f
C12536 FILLER_0_7_72/a_2364_375# FILLER_0_6_90/a_484_472# 0.001684f
C12537 _031_ FILLER_0_2_111/a_1380_472# 0.01562f
C12538 net81 FILLER_0_15_235/a_36_472# 0.001855f
C12539 _098_ FILLER_0_19_171/a_484_472# 0.010731f
C12540 trimb[3] net38 0.002836f
C12541 FILLER_0_5_54/a_1020_375# trim_mask\[1\] 0.010745f
C12542 output46/a_224_472# net44 0.003804f
C12543 FILLER_0_18_2/a_932_472# _452_/a_2225_156# 0.001256f
C12544 FILLER_0_4_144/a_484_472# _081_ 0.001145f
C12545 FILLER_0_4_144/a_36_472# _152_ 0.008211f
C12546 FILLER_0_21_125/a_572_375# _022_ 0.006025f
C12547 FILLER_0_16_89/a_1020_375# net14 0.029702f
C12548 _028_ net52 0.150861f
C12549 FILLER_0_20_87/a_36_472# vss 0.006244f
C12550 state\[1\] _071_ 0.196063f
C12551 fanout63/a_36_160# FILLER_0_15_228/a_124_375# 0.001177f
C12552 net7 _064_ 0.001538f
C12553 _451_/a_1040_527# vdd 0.004038f
C12554 net81 vss 0.766885f
C12555 fanout56/a_36_113# _098_ 0.019463f
C12556 _446_/a_2248_156# net40 0.037373f
C12557 _062_ FILLER_0_8_156/a_124_375# 0.008116f
C12558 _247_/a_36_160# _060_ 0.055366f
C12559 _426_/a_36_151# FILLER_0_8_247/a_484_472# 0.001723f
C12560 _070_ FILLER_0_10_94/a_572_375# 0.009837f
C12561 net57 _427_/a_2248_156# 0.002706f
C12562 cal input1/a_36_113# 0.025739f
C12563 vss _160_ 1.119894f
C12564 _443_/a_36_151# FILLER_0_2_127/a_124_375# 0.073306f
C12565 net55 _040_ 0.107198f
C12566 _162_ vdd 0.073371f
C12567 fanout60/a_36_160# net61 0.001167f
C12568 input4/a_36_68# net4 0.004679f
C12569 _421_/a_2248_156# net19 0.016721f
C12570 FILLER_0_12_2/a_572_375# _450_/a_36_151# 0.001597f
C12571 net57 _176_ 0.192223f
C12572 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1468_375# 0.086742f
C12573 _415_/a_1308_423# net19 0.001498f
C12574 _308_/a_848_380# net14 0.021982f
C12575 _413_/a_2560_156# vss 0.001097f
C12576 _086_ _115_ 0.4112f
C12577 net54 _025_ 0.00573f
C12578 net20 net48 0.035427f
C12579 _058_ _313_/a_67_603# 0.010094f
C12580 output25/a_224_472# _423_/a_2665_112# 0.001396f
C12581 _131_ vdd 1.344823f
C12582 FILLER_0_16_107/a_572_375# net36 0.001706f
C12583 _091_ FILLER_0_15_212/a_932_472# 0.008749f
C12584 _078_ _122_ 0.185069f
C12585 _083_ calibrate 0.001446f
C12586 net68 trim_val\[0\] 0.052045f
C12587 _223_/a_36_160# vss 0.007187f
C12588 FILLER_0_7_146/a_124_375# calibrate 0.014163f
C12589 _423_/a_36_151# net40 0.004045f
C12590 _132_ net54 0.016007f
C12591 FILLER_0_19_55/a_36_472# _012_ 0.001667f
C12592 _346_/a_665_69# _141_ 0.002048f
C12593 net56 _433_/a_2665_112# 0.003434f
C12594 net22 _048_ 0.268142f
C12595 input1/a_36_113# en 0.036849f
C12596 _367_/a_36_68# _156_ 0.096366f
C12597 FILLER_0_14_91/a_484_472# _095_ 0.011772f
C12598 _261_/a_36_160# FILLER_0_5_148/a_36_472# 0.195478f
C12599 _059_ FILLER_0_5_148/a_124_375# 0.007657f
C12600 _128_ FILLER_0_9_142/a_36_472# 0.005101f
C12601 _432_/a_2665_112# _136_ 0.002691f
C12602 net79 _100_ 0.170973f
C12603 net31 _419_/a_2665_112# 0.004446f
C12604 net62 _094_ 0.04063f
C12605 FILLER_0_20_87/a_124_375# _437_/a_36_151# 0.059049f
C12606 net15 _052_ 0.001074f
C12607 _130_ _125_ 0.002745f
C12608 _372_/a_1194_69# _163_ 0.001328f
C12609 FILLER_0_20_169/a_124_375# mask\[6\] 0.001178f
C12610 FILLER_0_18_37/a_124_375# vss 0.002958f
C12611 FILLER_0_18_37/a_572_375# vdd 0.02259f
C12612 FILLER_0_0_130/a_36_472# _442_/a_36_151# 0.001723f
C12613 _429_/a_36_151# vdd 0.076815f
C12614 fanout50/a_36_160# _164_ 0.08721f
C12615 output11/a_224_472# net10 0.095679f
C12616 _104_ net30 0.001375f
C12617 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_124_375# 0.012222f
C12618 _233_/a_36_160# net47 0.054273f
C12619 _239_/a_36_160# vss 0.001596f
C12620 _126_ _332_/a_36_472# 0.009299f
C12621 FILLER_0_13_65/a_36_472# cal_count\[1\] 0.016393f
C12622 net20 _420_/a_2665_112# 0.030202f
C12623 net18 vdd 1.496006f
C12624 vss net30 0.17209f
C12625 _095_ state\[1\] 0.069906f
C12626 _129_ _125_ 0.069221f
C12627 _053_ calibrate 0.081635f
C12628 _275_/a_224_472# _091_ 0.003461f
C12629 net81 fanout76/a_36_160# 0.041089f
C12630 _196_/a_36_160# vdd 0.106963f
C12631 output7/a_224_472# trim[2] 0.008581f
C12632 fanout68/a_36_113# vdd 0.012621f
C12633 ctln[5] _448_/a_36_151# 0.009209f
C12634 net56 vdd 0.277166f
C12635 _430_/a_1308_423# _429_/a_36_151# 0.001722f
C12636 _074_ net22 0.079421f
C12637 output47/a_224_472# vss 0.002843f
C12638 _396_/a_224_472# _095_ 0.001351f
C12639 _437_/a_2665_112# net14 0.002936f
C12640 _053_ net21 0.036284f
C12641 _072_ net4 0.097916f
C12642 _394_/a_718_524# vss 0.002666f
C12643 output31/a_224_472# _289_/a_36_472# 0.00101f
C12644 _263_/a_224_472# net59 0.002558f
C12645 net41 _054_ 0.035503f
C12646 _076_ net22 0.03249f
C12647 net67 trim_val\[0\] 0.382079f
C12648 FILLER_0_7_72/a_1916_375# net50 0.059471f
C12649 net81 _195_/a_67_603# 0.002322f
C12650 net20 FILLER_0_15_212/a_1020_375# 0.001629f
C12651 net52 trim_mask\[4\] 0.034276f
C12652 FILLER_0_13_80/a_124_375# vss 0.042254f
C12653 FILLER_0_13_80/a_36_472# vdd 0.087291f
C12654 _422_/a_2560_156# _009_ 0.002551f
C12655 _053_ _414_/a_36_151# 0.035994f
C12656 _408_/a_718_524# net40 0.011463f
C12657 ctln[7] _442_/a_2560_156# 0.001742f
C12658 _254_/a_448_472# net22 0.009088f
C12659 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_124_375# 0.009654f
C12660 net52 net47 0.039912f
C12661 _131_ _135_ 0.068855f
C12662 FILLER_0_18_2/a_932_472# net44 0.012286f
C12663 _098_ FILLER_0_15_235/a_484_472# 0.004898f
C12664 FILLER_0_20_177/a_1380_472# _098_ 0.00679f
C12665 _099_ _282_/a_36_160# 0.005808f
C12666 net62 net78 0.001947f
C12667 _020_ net73 0.057454f
C12668 net55 _452_/a_2225_156# 0.022788f
C12669 net49 net47 0.53353f
C12670 _444_/a_448_472# net17 0.022222f
C12671 _068_ _311_/a_2180_473# 0.001454f
C12672 net41 vss 0.810444f
C12673 FILLER_0_18_177/a_2812_375# net21 0.048071f
C12674 net60 _420_/a_2560_156# 0.001358f
C12675 net15 FILLER_0_5_54/a_1468_375# 0.039975f
C12676 net41 _178_ 0.019945f
C12677 ctln[1] vdd 0.825166f
C12678 _394_/a_728_93# _174_ 0.012471f
C12679 _425_/a_36_151# calibrate 0.071513f
C12680 FILLER_0_3_54/a_36_472# _164_ 0.012512f
C12681 FILLER_0_8_24/a_124_375# net17 0.039695f
C12682 _065_ net68 0.194392f
C12683 trim_mask\[1\] FILLER_0_6_47/a_3172_472# 0.004605f
C12684 mask\[5\] FILLER_0_20_177/a_572_375# 0.013294f
C12685 net62 FILLER_0_14_235/a_572_375# 0.017549f
C12686 _411_/a_2560_156# _073_ 0.002649f
C12687 _033_ _444_/a_796_472# 0.0099f
C12688 _165_ _444_/a_2248_156# 0.006027f
C12689 _414_/a_2560_156# vss 0.001078f
C12690 net44 FILLER_0_8_2/a_36_472# 0.005851f
C12691 _245_/a_672_472# _039_ 0.001025f
C12692 _048_ vdd 0.270091f
C12693 _417_/a_36_151# vss 0.040392f
C12694 net19 net8 0.056454f
C12695 _414_/a_448_472# _053_ 0.065053f
C12696 FILLER_0_7_72/a_2812_375# _053_ 0.016329f
C12697 FILLER_0_4_123/a_124_375# vdd 0.027816f
C12698 FILLER_0_19_47/a_484_472# vdd 0.001133f
C12699 FILLER_0_19_47/a_36_472# vss 0.001559f
C12700 _220_/a_67_603# vdd 0.020078f
C12701 net18 _416_/a_1204_472# 0.027218f
C12702 _016_ _427_/a_36_151# 0.00483f
C12703 _374_/a_36_68# vss 0.047832f
C12704 mask\[8\] FILLER_0_22_86/a_1468_375# 0.015339f
C12705 net35 FILLER_0_22_86/a_1020_375# 0.010202f
C12706 FILLER_0_7_59/a_36_472# vdd 0.016778f
C12707 FILLER_0_7_59/a_572_375# vss 0.017487f
C12708 _075_ _414_/a_2560_156# 0.026328f
C12709 FILLER_0_13_212/a_1020_375# _043_ 0.01418f
C12710 _193_/a_36_160# _416_/a_36_151# 0.065269f
C12711 FILLER_0_5_128/a_36_472# _070_ 0.036f
C12712 _414_/a_2248_156# _056_ 0.001452f
C12713 net35 FILLER_0_22_128/a_1828_472# 0.016187f
C12714 net17 _452_/a_2225_156# 0.001943f
C12715 _093_ _198_/a_67_603# 0.004447f
C12716 net79 _060_ 0.019511f
C12717 net57 _267_/a_36_472# 0.032037f
C12718 _170_ vdd 0.18848f
C12719 net82 _386_/a_1084_68# 0.001068f
C12720 FILLER_0_12_2/a_124_375# net67 0.003339f
C12721 trimb[0] FILLER_0_20_2/a_36_472# 0.005458f
C12722 net68 FILLER_0_6_47/a_484_472# 0.005391f
C12723 _137_ _333_/a_36_160# 0.022811f
C12724 _077_ net37 0.003374f
C12725 FILLER_0_8_107/a_124_375# vdd 0.049132f
C12726 _098_ _437_/a_36_151# 0.092841f
C12727 _431_/a_36_151# FILLER_0_17_133/a_124_375# 0.059049f
C12728 FILLER_0_10_214/a_124_375# _069_ 0.014379f
C12729 _074_ vdd 1.221102f
C12730 _428_/a_36_151# net14 0.004485f
C12731 _091_ FILLER_0_18_177/a_124_375# 0.010316f
C12732 net20 net10 0.02842f
C12733 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_36_472# 0.009654f
C12734 _411_/a_1000_472# vss 0.002964f
C12735 FILLER_0_7_72/a_2364_375# net14 0.005919f
C12736 _077_ _439_/a_796_472# 0.007471f
C12737 _086_ _134_ 0.020487f
C12738 _013_ FILLER_0_17_56/a_484_472# 0.002659f
C12739 _448_/a_36_151# net59 0.062656f
C12740 _039_ net6 0.104745f
C12741 _413_/a_1000_472# _002_ 0.006249f
C12742 FILLER_0_11_101/a_124_375# vdd 0.024363f
C12743 _440_/a_2665_112# trim_mask\[1\] 0.007959f
C12744 _133_ vss 0.18326f
C12745 _076_ vdd 0.806117f
C12746 FILLER_0_18_100/a_36_472# _356_/a_36_472# 0.010679f
C12747 _081_ net22 0.103561f
C12748 mask\[4\] FILLER_0_18_139/a_1468_375# 0.023004f
C12749 _061_ _058_ 0.02828f
C12750 _144_ FILLER_0_18_107/a_1828_472# 0.001169f
C12751 _021_ _432_/a_796_472# 0.001666f
C12752 cal_itt\[2\] _253_/a_244_68# 0.001073f
C12753 FILLER_0_15_180/a_572_375# vss 0.010974f
C12754 FILLER_0_15_180/a_36_472# vdd 0.017678f
C12755 FILLER_0_9_28/a_1020_375# FILLER_0_10_37/a_36_472# 0.001597f
C12756 ctln[3] net58 0.00479f
C12757 _131_ _403_/a_224_472# 0.003274f
C12758 _414_/a_1308_423# net22 0.011978f
C12759 net32 net60 0.509175f
C12760 FILLER_0_1_98/a_36_472# _442_/a_2665_112# 0.002597f
C12761 ctln[0] vss 0.125714f
C12762 trim_mask\[2\] FILLER_0_3_78/a_36_472# 0.005209f
C12763 _116_ net79 0.081785f
C12764 _096_ _320_/a_1792_472# 0.001419f
C12765 output8/a_224_472# _411_/a_1308_423# 0.005111f
C12766 net65 net22 0.374917f
C12767 comp FILLER_0_12_2/a_124_375# 0.007468f
C12768 FILLER_0_14_50/a_36_472# vss 0.002954f
C12769 net34 _435_/a_1308_423# 0.008652f
C12770 _178_ FILLER_0_14_50/a_36_472# 0.001492f
C12771 vdd FILLER_0_13_72/a_124_375# -0.004549f
C12772 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_124_375# 0.009654f
C12773 net68 _440_/a_448_472# 0.02254f
C12774 _176_ _451_/a_2449_156# 0.038547f
C12775 FILLER_0_5_109/a_572_375# _153_ 0.03228f
C12776 net58 net5 0.387314f
C12777 _420_/a_2665_112# _009_ 0.001752f
C12778 _086_ _267_/a_672_472# 0.004515f
C12779 net55 net44 0.018961f
C12780 en_co_clk vdd 0.245319f
C12781 output31/a_224_472# net19 0.072666f
C12782 net23 net13 0.018808f
C12783 _072_ _058_ 0.029688f
C12784 _095_ _451_/a_1353_112# 0.00475f
C12785 _291_/a_36_160# _199_/a_36_160# 0.005575f
C12786 net52 _154_ 0.001512f
C12787 FILLER_0_12_136/a_1380_472# FILLER_0_11_142/a_572_375# 0.001543f
C12788 _136_ mask\[9\] 0.015204f
C12789 _074_ _251_/a_1130_472# 0.00237f
C12790 net75 net27 0.037524f
C12791 net73 FILLER_0_17_142/a_484_472# 0.001122f
C12792 _074_ net9 0.002862f
C12793 _063_ _445_/a_2665_112# 0.009759f
C12794 net63 _429_/a_36_151# 0.0144f
C12795 FILLER_0_17_72/a_1380_472# net36 0.021039f
C12796 result[6] ctlp[2] 0.001324f
C12797 _142_ FILLER_0_17_142/a_124_375# 0.011387f
C12798 _053_ FILLER_0_7_104/a_124_375# 0.012564f
C12799 _359_/a_1044_488# net74 0.005311f
C12800 _093_ _303_/a_36_472# 0.096502f
C12801 net52 FILLER_0_3_142/a_124_375# 0.002239f
C12802 _051_ _098_ 0.006332f
C12803 mask\[9\] _438_/a_1000_472# 0.056239f
C12804 FILLER_0_5_164/a_36_472# vss 0.001809f
C12805 FILLER_0_5_164/a_484_472# vdd 0.005235f
C12806 _251_/a_906_472# _068_ 0.001762f
C12807 fanout67/a_36_160# _220_/a_67_603# 0.005474f
C12808 net41 _184_ 0.065857f
C12809 net39 net40 0.279259f
C12810 FILLER_0_18_171/a_36_472# vss 0.0032f
C12811 net51 FILLER_0_12_28/a_36_472# 0.005661f
C12812 net20 net37 0.039674f
C12813 net52 _442_/a_448_472# 0.044149f
C12814 _036_ _160_ 0.034434f
C12815 net51 net40 0.060626f
C12816 _428_/a_36_151# FILLER_0_11_109/a_36_472# 0.001221f
C12817 FILLER_0_18_177/a_36_472# vss 0.002187f
C12818 FILLER_0_18_177/a_484_472# vdd 0.006177f
C12819 _427_/a_2248_156# net36 0.004462f
C12820 mask\[0\] FILLER_0_13_228/a_36_472# 0.002986f
C12821 net20 FILLER_0_3_221/a_1468_375# 0.007234f
C12822 FILLER_0_7_59/a_36_472# fanout67/a_36_160# 0.013068f
C12823 FILLER_0_9_28/a_1828_472# _042_ 0.001809f
C12824 net56 FILLER_0_16_154/a_572_375# 0.002321f
C12825 _450_/a_2225_156# _039_ 0.034731f
C12826 net18 _419_/a_796_472# 0.006586f
C12827 _439_/a_36_151# FILLER_0_6_47/a_2812_375# 0.001512f
C12828 mask\[4\] FILLER_0_18_209/a_484_472# 0.021522f
C12829 net16 FILLER_0_18_37/a_932_472# 0.008749f
C12830 net44 net17 0.046636f
C12831 _176_ net36 0.336675f
C12832 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_36_472# 0.086743f
C12833 net80 _137_ 0.260786f
C12834 net48 _265_/a_244_68# 0.00365f
C12835 FILLER_0_17_104/a_572_375# net14 0.004285f
C12836 net69 _441_/a_1000_472# 0.018209f
C12837 _429_/a_448_472# _043_ 0.003615f
C12838 calibrate FILLER_0_9_270/a_36_472# 0.00119f
C12839 FILLER_0_16_89/a_36_472# _177_ 0.048163f
C12840 FILLER_0_21_125/a_36_472# _144_ 0.008287f
C12841 _425_/a_796_472# vdd 0.002206f
C12842 net17 FILLER_0_20_15/a_1380_472# 0.012286f
C12843 FILLER_0_17_282/a_36_472# _418_/a_1308_423# 0.001295f
C12844 net73 FILLER_0_18_107/a_2276_472# 0.016723f
C12845 _081_ vdd 0.729534f
C12846 mask\[7\] FILLER_0_22_128/a_484_472# 0.010605f
C12847 FILLER_0_17_282/a_36_472# _006_ 0.002964f
C12848 _069_ _429_/a_36_151# 0.010076f
C12849 net37 FILLER_0_6_231/a_572_375# 0.001989f
C12850 mask\[8\] net71 0.424276f
C12851 FILLER_0_15_116/a_484_472# FILLER_0_14_107/a_1468_375# 0.001723f
C12852 mask\[7\] _049_ 0.234746f
C12853 FILLER_0_24_130/a_36_472# output23/a_224_472# 0.001994f
C12854 net53 _427_/a_1000_472# 0.008132f
C12855 net64 FILLER_0_9_270/a_572_375# 0.017924f
C12856 _247_/a_36_160# _228_/a_36_68# 0.001919f
C12857 _002_ FILLER_0_3_172/a_2276_472# 0.030358f
C12858 _067_ FILLER_0_12_20/a_572_375# 0.01186f
C12859 _448_/a_1000_472# net22 0.011389f
C12860 _414_/a_1308_423# vdd 0.004897f
C12861 FILLER_0_9_28/a_1916_375# _220_/a_67_603# 0.014522f
C12862 _050_ _352_/a_49_472# 0.005393f
C12863 _090_ net22 0.032492f
C12864 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3172_472# 0.026657f
C12865 _428_/a_1308_423# net74 0.0098f
C12866 cal_itt\[2\] FILLER_0_3_221/a_932_472# 0.016327f
C12867 net50 _439_/a_796_472# 0.002389f
C12868 net52 _439_/a_1204_472# 0.027632f
C12869 net3 FILLER_0_15_10/a_36_472# 0.002825f
C12870 _137_ mask\[1\] 0.782055f
C12871 net31 mask\[4\] 0.499009f
C12872 FILLER_0_4_49/a_572_375# vdd 0.005972f
C12873 _096_ _043_ 0.842762f
C12874 _098_ FILLER_0_16_154/a_1468_375# 0.009042f
C12875 net65 vdd 1.430654f
C12876 fanout54/a_36_160# FILLER_0_19_142/a_36_472# 0.002647f
C12877 _143_ _091_ 0.007204f
C12878 FILLER_0_18_2/a_2364_375# net38 0.001683f
C12879 cal_itt\[2\] _088_ 0.010847f
C12880 _307_/a_234_472# _126_ 0.00204f
C12881 _013_ FILLER_0_18_53/a_484_472# 0.012916f
C12882 output47/a_224_472# _095_ 0.012266f
C12883 _091_ FILLER_0_13_212/a_1380_472# 0.003507f
C12884 _136_ _337_/a_257_69# 0.002933f
C12885 _114_ _128_ 0.047516f
C12886 _015_ FILLER_0_8_247/a_484_472# 0.005458f
C12887 ctlp[6] output24/a_224_472# 0.004288f
C12888 _176_ FILLER_0_10_107/a_572_375# 0.012296f
C12889 FILLER_0_22_86/a_1020_375# vdd 0.008761f
C12890 _153_ net14 0.260217f
C12891 FILLER_0_11_78/a_572_375# _120_ 0.01683f
C12892 fanout77/a_36_113# _094_ 0.002244f
C12893 _095_ FILLER_0_13_80/a_124_375# 0.001989f
C12894 FILLER_0_22_128/a_1828_472# vdd 0.005724f
C12895 FILLER_0_22_128/a_1380_472# vss 0.007305f
C12896 FILLER_0_16_73/a_124_375# net15 0.005202f
C12897 _140_ _354_/a_49_472# 0.004731f
C12898 _186_ _181_ 0.018817f
C12899 result[8] _422_/a_448_472# 0.002989f
C12900 ctlp[3] _422_/a_36_151# 0.002627f
C12901 _411_/a_796_472# net75 0.006358f
C12902 _372_/a_3662_472# net23 0.002864f
C12903 _238_/a_67_603# _441_/a_2665_112# 0.015187f
C12904 net81 output37/a_224_472# 0.00641f
C12905 ctln[8] FILLER_0_0_96/a_36_472# 0.012298f
C12906 net56 FILLER_0_18_139/a_36_472# 0.002172f
C12907 _121_ vss 0.082882f
C12908 fanout78/a_36_113# vss 0.031944f
C12909 _174_ _180_ 0.102241f
C12910 _297_/a_36_472# _108_ 0.011437f
C12911 _445_/a_448_472# _034_ 0.03826f
C12912 _185_ _402_/a_728_93# 0.007151f
C12913 net36 FILLER_0_18_76/a_124_375# 0.001741f
C12914 net41 _095_ 0.641184f
C12915 net82 FILLER_0_3_172/a_36_472# 0.007612f
C12916 _080_ net59 0.038227f
C12917 _124_ FILLER_0_10_107/a_572_375# 0.002135f
C12918 _104_ _046_ 0.035267f
C12919 _067_ FILLER_0_12_28/a_124_375# 0.012779f
C12920 net78 _422_/a_36_151# 0.023285f
C12921 trim_mask\[2\] _447_/a_448_472# 0.002533f
C12922 trim_val\[2\] _447_/a_36_151# 0.022122f
C12923 FILLER_0_3_172/a_2812_375# net65 0.003745f
C12924 FILLER_0_3_172/a_36_472# fanout57/a_36_113# 0.19419f
C12925 _446_/a_1000_472# vdd 0.001598f
C12926 FILLER_0_4_197/a_36_472# _270_/a_36_472# 0.004546f
C12927 cal_itt\[2\] cal_itt\[0\] 0.011453f
C12928 _128_ _176_ 0.180252f
C12929 _391_/a_245_68# cal_count\[0\] 0.001201f
C12930 mask\[5\] FILLER_0_21_206/a_36_472# 0.019416f
C12931 _035_ net38 0.02987f
C12932 _003_ cal_itt\[3\] 0.054183f
C12933 _046_ vss 0.088886f
C12934 _008_ net19 0.027093f
C12935 _443_/a_448_472# vdd 0.007773f
C12936 _443_/a_36_151# vss 0.019802f
C12937 FILLER_0_22_86/a_124_375# _437_/a_36_151# 0.001597f
C12938 FILLER_0_15_116/a_484_472# vdd 0.006111f
C12939 net65 net9 0.061456f
C12940 _432_/a_36_151# FILLER_0_16_154/a_1468_375# 0.001107f
C12941 _414_/a_1288_156# cal_itt\[3\] 0.001354f
C12942 _120_ _042_ 0.031451f
C12943 ctln[5] vss 0.132862f
C12944 FILLER_0_12_136/a_1468_375# net23 0.021046f
C12945 _070_ _055_ 0.516713f
C12946 result[8] _108_ 0.007884f
C12947 net28 _196_/a_36_160# 0.060575f
C12948 FILLER_0_5_117/a_36_472# vdd 0.092171f
C12949 net20 FILLER_0_13_212/a_1468_375# 0.009573f
C12950 net68 _232_/a_67_603# 0.00184f
C12951 output48/a_224_472# _425_/a_36_151# 0.004037f
C12952 _439_/a_2665_112# net14 0.004943f
C12953 _448_/a_1000_472# vdd 0.004267f
C12954 net68 _220_/a_255_603# 0.001908f
C12955 _090_ vdd 0.751973f
C12956 _149_ FILLER_0_20_98/a_36_472# 0.067283f
C12957 _028_ FILLER_0_6_79/a_124_375# 0.015932f
C12958 _182_ _179_ 0.109377f
C12959 FILLER_0_16_57/a_572_375# net72 0.012909f
C12960 _425_/a_36_151# FILLER_0_8_247/a_124_375# 0.001597f
C12961 fanout77/a_36_113# net78 0.019286f
C12962 _128_ _124_ 0.111918f
C12963 FILLER_0_5_54/a_1468_375# net47 0.005049f
C12964 FILLER_0_7_59/a_484_472# net68 0.002785f
C12965 _261_/a_36_160# _059_ 0.004993f
C12966 net68 _453_/a_36_151# 0.039234f
C12967 net57 _428_/a_448_472# 0.032029f
C12968 _086_ _375_/a_692_497# 0.002565f
C12969 cal_itt\[3\] net37 0.03677f
C12970 net72 _183_ 0.093818f
C12971 _433_/a_2665_112# _145_ 0.018359f
C12972 FILLER_0_16_89/a_572_375# _136_ 0.069752f
C12973 _035_ net66 1.624557f
C12974 _098_ _204_/a_67_603# 0.00539f
C12975 net65 FILLER_0_2_165/a_124_375# 0.001177f
C12976 _242_/a_36_160# FILLER_0_5_164/a_124_375# 0.005705f
C12977 _132_ net74 0.031741f
C12978 _069_ _076_ 0.033276f
C12979 _274_/a_2552_68# vss 0.003123f
C12980 _126_ _070_ 0.089475f
C12981 _386_/a_1152_472# _163_ 0.004076f
C12982 _126_ FILLER_0_15_180/a_124_375# 0.001238f
C12983 FILLER_0_17_72/a_2812_375# vdd 0.005986f
C12984 FILLER_0_12_20/a_36_472# net47 0.020589f
C12985 FILLER_0_8_263/a_124_375# net19 0.039576f
C12986 _415_/a_2248_156# net27 0.022666f
C12987 mask\[0\] _137_ 0.009052f
C12988 net41 output41/a_224_472# 0.008587f
C12989 FILLER_0_4_107/a_932_472# vdd 0.00987f
C12990 FILLER_0_16_89/a_36_472# _451_/a_2225_156# 0.001329f
C12991 net34 net61 0.037731f
C12992 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_124_375# 0.001597f
C12993 result[6] FILLER_0_21_286/a_572_375# 0.015047f
C12994 trim_mask\[4\] _370_/a_124_24# 0.015021f
C12995 _132_ _144_ 0.185339f
C12996 _427_/a_36_151# vss 0.019281f
C12997 net72 FILLER_0_15_59/a_572_375# 0.00799f
C12998 output7/a_224_472# vdd 0.086699f
C12999 net52 FILLER_0_2_111/a_36_472# 0.0659f
C13000 _029_ vdd 0.223076f
C13001 _043_ FILLER_0_13_72/a_572_375# 0.013294f
C13002 net41 _402_/a_1296_93# 0.001707f
C13003 _091_ _429_/a_2248_156# 0.006148f
C13004 _370_/a_124_24# net47 0.017609f
C13005 net18 net77 0.378783f
C13006 _424_/a_2665_112# FILLER_0_21_60/a_572_375# 0.001077f
C13007 _093_ FILLER_0_17_133/a_124_375# 0.009649f
C13008 net63 FILLER_0_18_177/a_484_472# 0.061539f
C13009 FILLER_0_15_150/a_124_375# net23 0.03361f
C13010 trim_mask\[2\] FILLER_0_2_93/a_572_375# 0.002818f
C13011 net52 _440_/a_1000_472# 0.013793f
C13012 net60 _421_/a_2665_112# 0.044114f
C13013 vdd _145_ 0.082579f
C13014 _321_/a_170_472# vss 0.024882f
C13015 FILLER_0_14_50/a_36_472# _095_ 0.013704f
C13016 fanout74/a_36_113# _032_ 0.012909f
C13017 _452_/a_36_151# _041_ 0.013289f
C13018 _363_/a_36_68# _151_ 0.020916f
C13019 FILLER_0_11_142/a_484_472# _120_ 0.007893f
C13020 _408_/a_56_524# vdd 0.003158f
C13021 _408_/a_728_93# vss 0.001345f
C13022 _163_ net22 0.005017f
C13023 net49 _440_/a_1000_472# 0.020434f
C13024 FILLER_0_13_142/a_1380_472# vss 0.004953f
C13025 FILLER_0_7_59/a_484_472# net67 0.03109f
C13026 _235_/a_255_603# trim_val\[2\] 0.002471f
C13027 _078_ FILLER_0_4_213/a_572_375# 0.02957f
C13028 output33/a_224_472# net60 0.002526f
C13029 _447_/a_1000_472# vdd 0.003392f
C13030 state\[0\] FILLER_0_9_223/a_36_472# 0.002846f
C13031 _032_ FILLER_0_2_127/a_124_375# 0.002221f
C13032 net57 FILLER_0_8_156/a_572_375# 0.014948f
C13033 _318_/a_224_472# vdd 0.001873f
C13034 _136_ _067_ 0.051914f
C13035 _141_ FILLER_0_17_142/a_572_375# 0.029028f
C13036 _431_/a_1308_423# net36 0.002865f
C13037 _081_ FILLER_0_5_198/a_572_375# 0.001285f
C13038 FILLER_0_12_2/a_572_375# _039_ 0.005407f
C13039 FILLER_0_11_64/a_36_472# _453_/a_36_151# 0.001723f
C13040 result[2] result[3] 0.09741f
C13041 net23 FILLER_0_22_128/a_1916_375# 0.004205f
C13042 net59 vss 1.191297f
C13043 FILLER_0_5_109/a_124_375# _151_ 0.003377f
C13044 _189_/a_67_603# net79 0.008944f
C13045 _137_ FILLER_0_16_154/a_36_472# 0.005011f
C13046 output29/a_224_472# _193_/a_36_160# 0.006363f
C13047 net47 net40 0.635497f
C13048 FILLER_0_0_198/a_36_472# vdd 0.052226f
C13049 FILLER_0_0_198/a_124_375# vss 0.017602f
C13050 _315_/a_36_68# net23 0.030384f
C13051 FILLER_0_9_223/a_572_375# _076_ 0.034523f
C13052 _155_ vdd 0.193832f
C13053 net15 _453_/a_2665_112# 0.011775f
C13054 fanout60/a_36_160# net62 0.049222f
C13055 net68 net69 0.053856f
C13056 _008_ _419_/a_448_472# 0.01758f
C13057 output9/a_224_472# cal_itt\[0\] 0.008307f
C13058 net74 _370_/a_124_24# 0.083426f
C13059 _075_ net59 0.01129f
C13060 net20 _429_/a_1308_423# 0.001186f
C13061 vss FILLER_0_10_94/a_484_472# 0.001244f
C13062 _091_ _248_/a_36_68# 0.071763f
C13063 _444_/a_796_472# _054_ 0.001838f
C13064 _071_ _121_ 0.007734f
C13065 _077_ _453_/a_448_472# 0.057515f
C13066 output44/a_224_472# FILLER_0_18_2/a_1020_375# 0.032639f
C13067 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_124_375# 0.007947f
C13068 _418_/a_2665_112# _417_/a_2665_112# 0.00131f
C13069 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_36_472# 0.026657f
C13070 _146_ vss 0.078821f
C13071 result[9] _419_/a_1308_423# 0.012036f
C13072 net82 FILLER_0_2_177/a_484_472# 0.001777f
C13073 _293_/a_36_472# _093_ 0.004121f
C13074 FILLER_0_8_24/a_36_472# _054_ 0.007348f
C13075 _449_/a_36_151# FILLER_0_13_72/a_124_375# 0.059049f
C13076 cal_count\[1\] FILLER_0_15_59/a_36_472# 0.00544f
C13077 _180_ FILLER_0_15_59/a_124_375# 0.009926f
C13078 _138_ _043_ 0.005826f
C13079 ctln[0] output41/a_224_472# 0.001583f
C13080 _415_/a_36_151# vss 0.003124f
C13081 net65 FILLER_0_2_177/a_572_375# 0.017058f
C13082 FILLER_0_14_91/a_484_472# _070_ 0.001773f
C13083 _085_ cal_count\[3\] 0.653405f
C13084 _025_ _436_/a_1204_472# 0.01349f
C13085 net69 _156_ 0.008057f
C13086 _449_/a_1308_423# net55 0.001985f
C13087 _422_/a_448_472# _109_ 0.006344f
C13088 _430_/a_796_472# net21 0.015066f
C13089 FILLER_0_5_206/a_36_472# net22 0.049294f
C13090 _122_ vss 0.750387f
C13091 _090_ _279_/a_244_68# 0.001986f
C13092 net33 _434_/a_36_151# 0.002776f
C13093 _083_ FILLER_0_3_221/a_572_375# 0.001072f
C13094 net64 FILLER_0_15_235/a_36_472# 0.046292f
C13095 FILLER_0_16_37/a_36_472# vss 0.005874f
C13096 _444_/a_1000_472# vdd 0.004148f
C13097 state\[0\] FILLER_0_12_220/a_932_472# 0.001003f
C13098 FILLER_0_7_233/a_36_472# vdd 0.016804f
C13099 FILLER_0_7_233/a_124_375# vss 0.003952f
C13100 _178_ FILLER_0_16_37/a_36_472# 0.007425f
C13101 FILLER_0_4_185/a_36_472# _002_ 0.004231f
C13102 cal_count\[3\] _408_/a_1936_472# 0.007046f
C13103 _044_ FILLER_0_13_290/a_36_472# 0.001194f
C13104 ctln[7] vss 0.132613f
C13105 _411_/a_36_151# FILLER_0_0_232/a_36_472# 0.001723f
C13106 FILLER_0_0_232/a_124_375# vdd 0.012494f
C13107 _000_ _083_ 0.017601f
C13108 FILLER_0_10_256/a_36_472# vss 0.001792f
C13109 _327_/a_36_472# _126_ 0.011444f
C13110 FILLER_0_8_24/a_36_472# vss 0.001239f
C13111 FILLER_0_8_24/a_484_472# vdd 0.009032f
C13112 net78 _419_/a_36_151# 0.007437f
C13113 _227_/a_36_160# vss 0.010455f
C13114 net64 vss 0.636644f
C13115 _453_/a_2665_112# net51 0.046426f
C13116 net11 vdd 0.330644f
C13117 _411_/a_2248_156# _084_ 0.002258f
C13118 _166_ _160_ 0.492224f
C13119 FILLER_0_4_144/a_124_375# net23 0.011315f
C13120 fanout51/a_36_113# FILLER_0_11_64/a_36_472# 0.001396f
C13121 net35 FILLER_0_23_88/a_36_472# 0.00675f
C13122 _440_/a_2248_156# _164_ 0.054298f
C13123 FILLER_0_4_144/a_572_375# trim_mask\[4\] 0.014071f
C13124 _272_/a_36_472# net76 0.04597f
C13125 FILLER_0_10_78/a_1468_375# _171_ 0.034647f
C13126 _070_ state\[1\] 0.032046f
C13127 net38 _452_/a_1353_112# 0.005918f
C13128 _075_ _122_ 0.030339f
C13129 _169_ vss 0.037006f
C13130 _163_ vdd 0.418075f
C13131 FILLER_0_4_49/a_36_472# net68 0.00894f
C13132 _010_ _420_/a_2248_156# 0.047408f
C13133 _159_ _370_/a_124_24# 0.021983f
C13134 fanout61/a_36_113# ctlp[1] 0.019606f
C13135 FILLER_0_0_96/a_36_472# net14 0.009584f
C13136 FILLER_0_2_93/a_484_472# vss 0.003689f
C13137 FILLER_0_4_144/a_572_375# net47 0.011686f
C13138 FILLER_0_19_171/a_1380_472# vss 0.004488f
C13139 _430_/a_1000_472# _091_ 0.025041f
C13140 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_484_472# 0.013276f
C13141 net58 result[1] 0.004614f
C13142 trim[4] net38 0.095379f
C13143 mask\[8\] _437_/a_1000_472# 0.00112f
C13144 output15/a_224_472# vdd 0.025731f
C13145 FILLER_0_21_28/a_124_375# vdd 0.014155f
C13146 FILLER_0_11_78/a_124_375# vdd -0.011022f
C13147 net23 FILLER_0_5_148/a_484_472# 0.047258f
C13148 net44 _452_/a_2449_156# 0.0059f
C13149 output10/a_224_472# FILLER_0_0_266/a_36_472# 0.023414f
C13150 _109_ _108_ 0.001806f
C13151 net5 clk 0.042578f
C13152 FILLER_0_0_96/a_124_375# trim_mask\[3\] 0.006277f
C13153 FILLER_0_18_2/a_2276_472# vdd 0.004679f
C13154 trim_val\[2\] vss 0.027243f
C13155 FILLER_0_6_239/a_124_375# _123_ 0.044771f
C13156 output35/a_224_472# _204_/a_67_603# 0.012678f
C13157 net19 _109_ 0.005991f
C13158 FILLER_0_2_93/a_36_472# _441_/a_2665_112# 0.007491f
C13159 _253_/a_1528_68# cal_itt\[1\] 0.002251f
C13160 _131_ FILLER_0_11_124/a_124_375# 0.008946f
C13161 net15 _168_ 0.04897f
C13162 ctln[3] _411_/a_448_472# 0.00336f
C13163 FILLER_0_23_44/a_36_472# vss 0.002194f
C13164 FILLER_0_23_44/a_484_472# vdd 0.003276f
C13165 FILLER_0_2_165/a_36_472# net59 0.067972f
C13166 net15 _441_/a_796_472# 0.021664f
C13167 _305_/a_36_159# _112_ 0.001664f
C13168 FILLER_0_7_162/a_36_472# _062_ 0.016683f
C13169 FILLER_0_5_164/a_36_472# _385_/a_36_68# 0.001674f
C13170 _173_ FILLER_0_12_28/a_36_472# 0.001633f
C13171 _002_ _079_ 0.051048f
C13172 FILLER_0_18_209/a_484_472# _201_/a_67_603# 0.001605f
C13173 output45/a_224_472# net46 0.005906f
C13174 _408_/a_728_93# _184_ 0.001389f
C13175 _440_/a_2560_156# net47 0.003888f
C13176 net29 _101_ 0.007132f
C13177 _136_ net23 0.031512f
C13178 _105_ net32 2.08459f
C13179 _418_/a_1308_423# vss 0.001913f
C13180 FILLER_0_14_107/a_1380_472# vss 0.001338f
C13181 _006_ vss 0.111492f
C13182 _093_ FILLER_0_17_161/a_124_375# 0.002431f
C13183 mask\[5\] _339_/a_36_160# 0.007734f
C13184 FILLER_0_10_28/a_124_375# net51 0.00979f
C13185 trimb[1] FILLER_0_18_2/a_484_472# 0.009245f
C13186 FILLER_0_22_177/a_484_472# net33 0.013149f
C13187 _433_/a_1000_472# _022_ 0.05526f
C13188 _043_ _113_ 0.048005f
C13189 FILLER_0_15_116/a_36_472# _095_ 0.001098f
C13190 net52 FILLER_0_9_72/a_572_375# 0.022582f
C13191 FILLER_0_21_286/a_36_472# vss 0.004123f
C13192 FILLER_0_21_286/a_484_472# vdd 0.007903f
C13193 FILLER_0_13_142/a_124_375# net23 0.003962f
C13194 _103_ vss 0.098913f
C13195 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_36_472# 0.009654f
C13196 output39/a_224_472# vdd 0.022593f
C13197 net20 output31/a_224_472# 0.004424f
C13198 FILLER_0_1_266/a_572_375# vdd 0.030477f
C13199 _376_/a_36_160# _164_ 0.004503f
C13200 _069_ _090_ 1.067281f
C13201 _114_ _176_ 0.147182f
C13202 _117_ vdd 0.050188f
C13203 FILLER_0_16_73/a_124_375# FILLER_0_16_57/a_1468_375# 0.012222f
C13204 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_484_472# 0.013276f
C13205 FILLER_0_5_206/a_36_472# vdd 0.090007f
C13206 FILLER_0_5_206/a_124_375# vss 0.050652f
C13207 _077_ FILLER_0_9_60/a_124_375# 0.051389f
C13208 cal_count\[3\] _062_ 0.004405f
C13209 net31 _201_/a_67_603# 0.015773f
C13210 _377_/a_36_472# net68 0.001305f
C13211 _071_ FILLER_0_13_142/a_1380_472# 0.001617f
C13212 _059_ _062_ 0.161331f
C13213 _303_/a_36_472# _012_ 0.001735f
C13214 _402_/a_2172_497# cal_count\[1\] 0.008211f
C13215 FILLER_0_18_61/a_36_472# vss 0.00605f
C13216 _428_/a_2248_156# _131_ 0.005621f
C13217 FILLER_0_16_107/a_36_472# _093_ 0.001526f
C13218 trim[2] trim[3] 0.056575f
C13219 _017_ net14 0.014743f
C13220 _430_/a_2560_156# net36 0.00164f
C13221 net82 FILLER_0_3_221/a_124_375# 0.015932f
C13222 output47/a_224_472# _185_ 0.001177f
C13223 _075_ FILLER_0_5_206/a_124_375# 0.001024f
C13224 FILLER_0_1_98/a_36_472# vdd 0.009937f
C13225 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_36_472# 0.026657f
C13226 vss FILLER_0_4_91/a_572_375# 0.055113f
C13227 _077_ trim_mask\[0\] 0.090587f
C13228 _098_ FILLER_0_20_87/a_36_472# 0.016138f
C13229 _074_ FILLER_0_6_231/a_484_472# 0.004409f
C13230 vss _433_/a_3041_156# 0.001287f
C13231 fanout75/a_36_113# _083_ 0.002133f
C13232 FILLER_0_3_172/a_1380_472# net22 0.012284f
C13233 net81 _098_ 0.029506f
C13234 _438_/a_2665_112# FILLER_0_19_111/a_36_472# 0.007491f
C13235 net32 output19/a_224_472# 0.101682f
C13236 _422_/a_1204_472# mask\[7\] 0.025592f
C13237 output16/a_224_472# ctln[9] 0.08624f
C13238 output13/a_224_472# net12 0.002723f
C13239 result[6] _420_/a_1204_472# 0.002681f
C13240 FILLER_0_13_65/a_36_472# _043_ 0.013651f
C13241 net18 output30/a_224_472# 0.08667f
C13242 net57 _315_/a_36_68# 0.0036f
C13243 FILLER_0_11_78/a_484_472# _389_/a_36_148# 0.001043f
C13244 mask\[5\] ctlp[4] 0.001643f
C13245 ctln[2] net58 0.025352f
C13246 _053_ _151_ 0.538643f
C13247 _427_/a_36_151# _095_ 0.029048f
C13248 FILLER_0_16_37/a_36_472# _184_ 0.001522f
C13249 net27 _426_/a_448_472# 0.023676f
C13250 net38 _398_/a_36_113# 0.061273f
C13251 _093_ FILLER_0_17_72/a_2724_472# 0.02416f
C13252 FILLER_0_17_72/a_2276_472# mask\[9\] 0.006767f
C13253 FILLER_0_15_235/a_484_472# mask\[1\] 0.014415f
C13254 output34/a_224_472# result[7] 0.057094f
C13255 mask\[4\] FILLER_0_20_193/a_484_472# 0.001215f
C13256 FILLER_0_16_73/a_36_472# _394_/a_1336_472# 0.00108f
C13257 _066_ _386_/a_124_24# 0.059053f
C13258 net41 _185_ 0.029318f
C13259 net74 FILLER_0_13_142/a_572_375# 0.001412f
C13260 FILLER_0_5_198/a_36_472# net59 0.059378f
C13261 _431_/a_36_151# FILLER_0_18_107/a_2724_472# 0.00271f
C13262 _086_ _255_/a_224_552# 0.073601f
C13263 _428_/a_36_151# _017_ 0.021229f
C13264 fanout49/a_36_160# _160_ 0.009662f
C13265 _369_/a_692_472# vdd 0.003899f
C13266 _377_/a_36_472# net67 0.005639f
C13267 net29 _094_ 0.313846f
C13268 net36 FILLER_0_15_212/a_1380_472# 0.006416f
C13269 _408_/a_728_93# _095_ 0.040366f
C13270 net53 net23 0.501857f
C13271 _411_/a_1308_423# _000_ 0.004012f
C13272 _095_ FILLER_0_13_142/a_1380_472# 0.001782f
C13273 _104_ _422_/a_2665_112# 0.040586f
C13274 net2 input5/a_36_113# 0.007518f
C13275 input2/a_36_113# net5 0.001761f
C13276 FILLER_0_2_177/a_36_472# net59 0.007582f
C13277 FILLER_0_7_104/a_36_472# FILLER_0_9_105/a_124_375# 0.001188f
C13278 _176_ _124_ 0.036117f
C13279 FILLER_0_11_142/a_36_472# vdd 0.110248f
C13280 FILLER_0_11_142/a_572_375# vss 0.052505f
C13281 _188_ net51 0.044278f
C13282 _322_/a_692_472# _129_ 0.004891f
C13283 FILLER_0_7_162/a_124_375# _062_ 0.010242f
C13284 _092_ FILLER_0_17_218/a_484_472# 0.007838f
C13285 FILLER_0_18_107/a_2812_375# vdd 0.004212f
C13286 net23 _386_/a_124_24# 0.010805f
C13287 _434_/a_448_472# mask\[6\] 0.060756f
C13288 FILLER_0_20_193/a_36_472# FILLER_0_19_187/a_572_375# 0.001543f
C13289 trim_mask\[4\] _386_/a_848_380# 0.001657f
C13290 _422_/a_2665_112# vss 0.006352f
C13291 _287_/a_36_472# vdd 0.072871f
C13292 FILLER_0_7_104/a_1020_375# vdd 0.010571f
C13293 output9/a_224_472# cal 0.011495f
C13294 ctln[2] net82 0.005498f
C13295 FILLER_0_7_72/a_36_472# _439_/a_448_472# 0.008036f
C13296 _431_/a_2560_156# net73 0.001018f
C13297 FILLER_0_18_139/a_36_472# _145_ 0.002415f
C13298 FILLER_0_8_138/a_124_375# _313_/a_67_603# 0.00744f
C13299 net79 FILLER_0_12_220/a_932_472# 0.005532f
C13300 net47 _386_/a_848_380# 0.003045f
C13301 result[6] _419_/a_2248_156# 0.002634f
C13302 _074_ _375_/a_1612_497# 0.004567f
C13303 FILLER_0_9_28/a_2812_375# net68 0.012462f
C13304 output29/a_224_472# _416_/a_36_151# 0.07368f
C13305 FILLER_0_9_28/a_2364_375# trim_val\[0\] 0.006639f
C13306 _069_ _314_/a_224_472# 0.003461f
C13307 result[7] _298_/a_224_472# 0.007724f
C13308 _026_ net71 0.406369f
C13309 mask\[4\] FILLER_0_18_177/a_2364_375# 0.01602f
C13310 output14/a_224_472# ctln[6] 0.007421f
C13311 net55 FILLER_0_21_60/a_124_375# 0.015315f
C13312 _174_ vss 0.188373f
C13313 mask\[3\] FILLER_0_16_241/a_36_472# 0.00209f
C13314 FILLER_0_17_72/a_484_472# FILLER_0_18_76/a_36_472# 0.05841f
C13315 calibrate _055_ 0.006584f
C13316 _178_ _174_ 0.012157f
C13317 mask\[3\] FILLER_0_18_177/a_1468_375# 0.002924f
C13318 _447_/a_796_472# _036_ 0.006511f
C13319 result[9] result[2] 0.001669f
C13320 _070_ _160_ 0.065914f
C13321 FILLER_0_23_88/a_124_375# vss 0.014165f
C13322 FILLER_0_23_88/a_36_472# vdd 0.002576f
C13323 FILLER_0_21_28/a_572_375# FILLER_0_19_28/a_484_472# 0.001512f
C13324 _415_/a_2665_112# net27 0.030051f
C13325 _115_ FILLER_0_11_78/a_484_472# 0.003641f
C13326 _122_ FILLER_0_5_198/a_36_472# 0.00305f
C13327 net47 _452_/a_1040_527# 0.014695f
C13328 _062_ _226_/a_452_68# 0.001697f
C13329 _131_ FILLER_0_17_104/a_1380_472# 0.004125f
C13330 _072_ _375_/a_692_497# 0.001113f
C13331 _441_/a_36_151# _030_ 0.005324f
C13332 mask\[9\] _149_ 0.040342f
C13333 net15 _423_/a_2248_156# 0.048449f
C13334 _097_ vss 0.00839f
C13335 _053_ FILLER_0_8_37/a_484_472# 0.002095f
C13336 _055_ net21 0.025995f
C13337 _093_ FILLER_0_18_139/a_1020_375# 0.003529f
C13338 output9/a_224_472# en 0.011047f
C13339 net50 FILLER_0_9_60/a_124_375# 0.001715f
C13340 fanout73/a_36_113# _136_ 0.002661f
C13341 net67 FILLER_0_6_37/a_124_375# 0.002918f
C13342 _449_/a_2248_156# _038_ 0.016483f
C13343 FILLER_0_5_54/a_1380_472# _440_/a_36_151# 0.001723f
C13344 FILLER_0_3_172/a_1380_472# vdd 0.043045f
C13345 net32 mask\[6\] 0.003248f
C13346 FILLER_0_15_212/a_1380_472# FILLER_0_15_228/a_36_472# 0.013277f
C13347 FILLER_0_5_198/a_484_472# net21 0.051161f
C13348 net41 _407_/a_36_472# 0.003257f
C13349 FILLER_0_21_125/a_484_472# _433_/a_36_151# 0.001723f
C13350 FILLER_0_11_109/a_124_375# FILLER_0_10_107/a_484_472# 0.001684f
C13351 net41 cal_count\[0\] 0.001014f
C13352 net20 _008_ 0.153014f
C13353 FILLER_0_7_104/a_484_472# _058_ 0.006506f
C13354 _414_/a_36_151# _055_ 0.001987f
C13355 cal_itt\[0\] _084_ 0.061227f
C13356 _422_/a_2665_112# _107_ 0.005055f
C13357 _052_ FILLER_0_18_37/a_484_472# 0.003861f
C13358 _424_/a_36_151# FILLER_0_20_31/a_124_375# 0.012574f
C13359 _114_ _267_/a_36_472# 0.011923f
C13360 ctlp[0] vss 0.005302f
C13361 net50 trim_mask\[0\] 0.002835f
C13362 FILLER_0_5_181/a_36_472# vss 0.001068f
C13363 net20 result[8] 0.014571f
C13364 _053_ _162_ 0.00209f
C13365 net44 output6/a_224_472# 0.078248f
C13366 vdd net6 0.134918f
C13367 _104_ mask\[2\] 0.002737f
C13368 FILLER_0_24_63/a_124_375# vss 0.03143f
C13369 trimb[3] FILLER_0_20_15/a_124_375# 0.001391f
C13370 _126_ net21 0.024842f
C13371 ctln[6] net22 0.014307f
C13372 net57 _136_ 0.168299f
C13373 FILLER_0_22_177/a_932_472# mask\[6\] 0.006573f
C13374 ctlp[1] net79 0.002676f
C13375 mask\[2\] vss 0.536426f
C13376 net35 FILLER_0_22_177/a_484_472# 0.00632f
C13377 _093_ FILLER_0_18_76/a_484_472# 0.024853f
C13378 net60 _094_ 0.579872f
C13379 mask\[9\] FILLER_0_18_76/a_36_472# 0.002584f
C13380 _412_/a_448_472# net2 0.033994f
C13381 _053_ _131_ 0.086215f
C13382 _128_ _246_/a_36_68# 0.01024f
C13383 net57 FILLER_0_13_142/a_124_375# 0.011369f
C13384 fanout70/a_36_113# fanout73/a_36_113# 0.001578f
C13385 _172_ vdd 0.008764f
C13386 net34 FILLER_0_22_128/a_1916_375# 0.04185f
C13387 net16 _041_ 0.029736f
C13388 net81 net58 0.375649f
C13389 net48 vdd 0.35704f
C13390 net75 FILLER_0_8_247/a_932_472# 0.006746f
C13391 net54 FILLER_0_18_139/a_1020_375# 0.003589f
C13392 output32/a_224_472# result[9] 0.047198f
C13393 mask\[5\] _434_/a_2248_156# 0.003462f
C13394 net2 net19 0.031976f
C13395 _360_/a_36_160# FILLER_0_4_123/a_36_472# 0.001165f
C13396 result[7] _419_/a_2248_156# 0.001916f
C13397 _132_ net70 0.534228f
C13398 output12/a_224_472# _037_ 0.00827f
C13399 FILLER_0_8_247/a_1020_375# vdd -0.002559f
C13400 _085_ _267_/a_224_472# 0.002907f
C13401 _176_ _267_/a_36_472# 0.001681f
C13402 _025_ FILLER_0_22_107/a_484_472# 0.00892f
C13403 trim_val\[3\] FILLER_0_2_93/a_124_375# 0.001032f
C13404 FILLER_0_7_72/a_932_472# vss 0.002763f
C13405 FILLER_0_19_125/a_124_375# FILLER_0_18_107/a_2276_472# 0.001684f
C13406 FILLER_0_9_223/a_484_472# _055_ 0.026026f
C13407 net81 _425_/a_448_472# 0.056225f
C13408 net55 FILLER_0_18_37/a_124_375# 0.005899f
C13409 _131_ _182_ 0.113302f
C13410 FILLER_0_7_195/a_124_375# cal_itt\[3\] 0.034632f
C13411 trim_val\[1\] _160_ 0.024279f
C13412 net76 FILLER_0_5_212/a_124_375# 0.004635f
C13413 _322_/a_848_380# _127_ 0.018892f
C13414 _015_ FILLER_0_10_247/a_36_472# 0.007508f
C13415 _067_ _389_/a_36_148# 0.002789f
C13416 output37/a_224_472# net59 0.001014f
C13417 _093_ FILLER_0_18_209/a_36_472# 0.007068f
C13418 FILLER_0_4_185/a_124_375# net76 0.053929f
C13419 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_572_375# 0.086635f
C13420 _441_/a_448_472# _164_ 0.016938f
C13421 _104_ _420_/a_2248_156# 0.027923f
C13422 _064_ net68 0.059889f
C13423 trim_val\[2\] _036_ 0.279133f
C13424 _077_ _256_/a_1612_497# 0.002724f
C13425 net81 _082_ 0.001633f
C13426 _061_ FILLER_0_8_156/a_484_472# 0.00255f
C13427 _379_/a_36_472# trim_mask\[1\] 0.003592f
C13428 net81 net82 0.063498f
C13429 _057_ _161_ 1.09228f
C13430 _013_ _424_/a_2248_156# 0.001828f
C13431 _420_/a_2665_112# vdd 0.024431f
C13432 _420_/a_2248_156# vss -0.001f
C13433 _095_ FILLER_0_14_107/a_1380_472# 0.011439f
C13434 result[6] output18/a_224_472# 0.003068f
C13435 fanout73/a_36_113# net53 0.047141f
C13436 FILLER_0_7_72/a_1916_375# vdd 0.015888f
C13437 net4 FILLER_0_12_220/a_1380_472# 0.016375f
C13438 net44 net3 0.195171f
C13439 _394_/a_1336_472# FILLER_0_13_72/a_36_472# 0.008136f
C13440 _394_/a_728_93# FILLER_0_13_72/a_572_375# 0.001064f
C13441 FILLER_0_15_205/a_36_472# net22 0.037011f
C13442 _018_ FILLER_0_15_205/a_124_375# 0.002309f
C13443 output26/a_224_472# FILLER_0_23_44/a_36_472# 0.026108f
C13444 _032_ vss 0.02257f
C13445 _086_ _120_ 0.408014f
C13446 net20 _060_ 0.0426f
C13447 mask\[5\] _202_/a_36_160# 0.00164f
C13448 vdd FILLER_0_16_115/a_36_472# 0.093403f
C13449 vss FILLER_0_16_115/a_124_375# 0.006358f
C13450 ctln[1] output10/a_224_472# 0.083631f
C13451 output47/a_224_472# net55 0.160037f
C13452 _098_ FILLER_0_15_180/a_572_375# 0.01526f
C13453 output42/a_224_472# trim[4] 0.017153f
C13454 cal_count\[1\] _451_/a_3129_107# 0.028519f
C13455 FILLER_0_16_89/a_1380_472# FILLER_0_17_72/a_3260_375# 0.001723f
C13456 _069_ _117_ 0.041311f
C13457 net80 FILLER_0_16_154/a_1468_375# 0.013593f
C13458 _142_ _341_/a_49_472# 0.011026f
C13459 net60 net78 0.030634f
C13460 net52 _443_/a_1204_472# 0.005165f
C13461 _413_/a_2560_156# net82 0.00101f
C13462 mask\[9\] FILLER_0_20_107/a_124_375# 0.004716f
C13463 trim_val\[4\] vss 0.192567f
C13464 vdd _450_/a_2225_156# 0.020301f
C13465 _099_ FILLER_0_15_235/a_484_472# 0.002657f
C13466 FILLER_0_16_57/a_124_375# vss 0.001678f
C13467 FILLER_0_16_57/a_572_375# vdd 0.004039f
C13468 FILLER_0_16_37/a_36_472# _402_/a_1296_93# 0.001477f
C13469 mask\[8\] _436_/a_1000_472# 0.001091f
C13470 net35 _436_/a_796_472# 0.002146f
C13471 net55 FILLER_0_13_80/a_124_375# 0.069951f
C13472 _174_ _401_/a_36_68# 0.033989f
C13473 net72 _181_ 0.004503f
C13474 FILLER_0_3_78/a_484_472# _160_ 0.004988f
C13475 _105_ output33/a_224_472# 0.099107f
C13476 _265_/a_916_472# _001_ 0.001719f
C13477 _063_ FILLER_0_6_37/a_36_472# 0.014315f
C13478 valid net19 0.00646f
C13479 _183_ vdd 0.109252f
C13480 _239_/a_36_160# net17 0.014703f
C13481 FILLER_0_19_195/a_36_472# _434_/a_2248_156# 0.001731f
C13482 FILLER_0_15_212/a_572_375# vss 0.005835f
C13483 FILLER_0_15_212/a_1020_375# vdd -0.00211f
C13484 cal_count\[3\] net14 0.028995f
C13485 ctln[6] vdd 0.116327f
C13486 net68 _042_ 0.037716f
C13487 net57 net53 0.053565f
C13488 _122_ _385_/a_36_68# 0.003549f
C13489 _195_/a_67_603# mask\[2\] 0.003161f
C13490 FILLER_0_20_177/a_484_472# _434_/a_36_151# 0.001723f
C13491 FILLER_0_16_154/a_932_472# vdd 0.00549f
C13492 FILLER_0_16_154/a_484_472# vss 0.003464f
C13493 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_124_375# 0.003732f
C13494 FILLER_0_15_150/a_124_375# net36 0.005687f
C13495 _445_/a_2248_156# _444_/a_36_151# 0.001081f
C13496 output21/a_224_472# net32 0.017976f
C13497 net41 net55 0.033821f
C13498 _065_ _447_/a_36_151# 0.043351f
C13499 net57 _386_/a_124_24# 0.037058f
C13500 net64 FILLER_0_12_236/a_36_472# 0.052381f
C13501 output37/a_224_472# net64 0.110037f
C13502 _144_ _352_/a_257_69# 0.001662f
C13503 trim_mask\[1\] FILLER_0_6_47/a_1020_375# 0.007169f
C13504 _058_ net23 0.075446f
C13505 trimb[1] FILLER_0_20_15/a_36_472# 0.001292f
C13506 FILLER_0_4_144/a_572_375# FILLER_0_5_148/a_124_375# 0.05841f
C13507 _434_/a_36_151# vdd 0.104871f
C13508 FILLER_0_19_111/a_572_375# vss 0.003337f
C13509 FILLER_0_19_111/a_36_472# vdd 0.034386f
C13510 _431_/a_2665_112# FILLER_0_16_154/a_124_375# 0.006271f
C13511 output47/a_224_472# net17 0.081437f
C13512 fanout80/a_36_113# vdd 0.033884f
C13513 net38 _190_/a_36_160# 0.062343f
C13514 _064_ net67 0.006691f
C13515 _419_/a_2665_112# vss 0.004064f
C13516 _419_/a_2560_156# vdd 0.003021f
C13517 mask\[5\] FILLER_0_20_193/a_124_375# 0.015793f
C13518 _144_ _433_/a_1204_472# 0.009472f
C13519 _074_ _083_ 0.035769f
C13520 FILLER_0_15_59/a_572_375# vdd 0.03104f
C13521 FILLER_0_15_59/a_124_375# vss 0.003806f
C13522 _077_ _073_ 0.009611f
C13523 net15 FILLER_0_11_64/a_124_375# 0.047331f
C13524 FILLER_0_18_107/a_1020_375# FILLER_0_19_111/a_572_375# 0.05841f
C13525 _077_ _330_/a_224_472# 0.001921f
C13526 _053_ _220_/a_67_603# 0.065611f
C13527 _004_ _005_ 0.004158f
C13528 _116_ FILLER_0_12_196/a_36_472# 0.010951f
C13529 FILLER_0_16_89/a_932_472# _093_ 0.002018f
C13530 _080_ FILLER_0_3_221/a_1020_375# 0.001414f
C13531 FILLER_0_12_136/a_932_472# _127_ 0.002804f
C13532 output8/a_224_472# FILLER_0_3_221/a_124_375# 0.03228f
C13533 _070_ _133_ 0.436976f
C13534 FILLER_0_18_171/a_36_472# _098_ 0.020038f
C13535 _076_ _083_ 0.006023f
C13536 _068_ _078_ 0.002973f
C13537 net54 FILLER_0_20_107/a_36_472# 0.050184f
C13538 _096_ _057_ 0.001547f
C13539 output36/a_224_472# net18 0.010751f
C13540 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_1020_375# 0.026339f
C13541 FILLER_0_19_195/a_36_472# _202_/a_36_160# 0.002647f
C13542 fanout69/a_36_113# vdd 0.00378f
C13543 net76 FILLER_0_3_172/a_1828_472# 0.051851f
C13544 net56 _137_ 0.0313f
C13545 FILLER_0_4_152/a_36_472# vdd 0.087397f
C13546 _053_ FILLER_0_7_59/a_36_472# 0.073877f
C13547 net67 net42 0.101108f
C13548 FILLER_0_7_146/a_124_375# _076_ 0.00688f
C13549 FILLER_0_7_146/a_36_472# _133_ 0.009796f
C13550 state\[1\] net21 0.210202f
C13551 _415_/a_1308_423# FILLER_0_9_270/a_124_375# 0.001064f
C13552 _088_ _260_/a_36_68# 0.003476f
C13553 net75 _253_/a_672_68# 0.003771f
C13554 _064_ _445_/a_448_472# 0.080931f
C13555 output36/a_224_472# _196_/a_36_160# 0.001309f
C13556 FILLER_0_13_212/a_484_472# net79 0.00402f
C13557 output33/a_224_472# output19/a_224_472# 0.115114f
C13558 net41 net17 0.911377f
C13559 net62 FILLER_0_13_212/a_932_472# 0.059367f
C13560 FILLER_0_4_91/a_484_472# _156_ 0.009828f
C13561 _077_ net15 0.238832f
C13562 FILLER_0_16_73/a_484_472# _040_ 0.004877f
C13563 net41 trim_val\[1\] 0.001912f
C13564 _412_/a_2665_112# en 0.015256f
C13565 net20 _093_ 0.398457f
C13566 net4 FILLER_0_3_221/a_932_472# 0.002116f
C13567 _004_ net75 0.003999f
C13568 net80 FILLER_0_22_177/a_1020_375# 0.00258f
C13569 mask\[5\] FILLER_0_18_177/a_1020_375# 0.001604f
C13570 FILLER_0_13_206/a_124_375# net22 0.024537f
C13571 _031_ FILLER_0_2_101/a_124_375# 0.00179f
C13572 _053_ FILLER_0_8_107/a_124_375# 0.002386f
C13573 _415_/a_796_472# net19 0.001468f
C13574 _412_/a_36_151# _001_ 0.006762f
C13575 FILLER_0_15_205/a_124_375# vss 0.026372f
C13576 FILLER_0_15_205/a_36_472# vdd 0.010089f
C13577 _053_ _074_ 0.503728f
C13578 _161_ _310_/a_49_472# 0.022411f
C13579 _147_ _146_ 0.001164f
C13580 ctln[4] vss 0.244634f
C13581 net22 net37 0.03068f
C13582 _450_/a_1353_112# net6 0.054189f
C13583 _450_/a_36_151# clkc 0.033095f
C13584 _106_ net64 0.001587f
C13585 _305_/a_36_159# net1 0.013619f
C13586 _016_ _130_ 0.114514f
C13587 net45 net46 0.038161f
C13588 trim_val\[3\] vss 0.249446f
C13589 _013_ net26 0.174966f
C13590 _088_ net4 0.096522f
C13591 FILLER_0_10_78/a_1020_375# vss 0.002352f
C13592 ctlp[9] vdd 0.17413f
C13593 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_36_472# 0.026657f
C13594 _360_/a_36_160# _152_ 0.040508f
C13595 FILLER_0_12_220/a_36_472# vdd 0.027911f
C13596 FILLER_0_12_220/a_1468_375# vss 0.057853f
C13597 _053_ _076_ 0.108358f
C13598 FILLER_0_11_64/a_124_375# net51 0.027848f
C13599 _413_/a_1308_423# net65 0.022097f
C13600 net10 vdd 0.227004f
C13601 net50 _447_/a_2248_156# 0.007602f
C13602 _426_/a_2665_112# calibrate 0.004837f
C13603 cal_count\[3\] FILLER_0_11_109/a_36_472# 0.00702f
C13604 FILLER_0_17_72/a_2364_375# _451_/a_448_472# 0.001512f
C13605 net40 _381_/a_36_472# 0.020876f
C13606 output39/a_224_472# _445_/a_1308_423# 0.010408f
C13607 net39 _445_/a_36_151# 0.006056f
C13608 _174_ _095_ 0.977766f
C13609 FILLER_0_20_193/a_124_375# FILLER_0_19_195/a_36_472# 0.001543f
C13610 _093_ FILLER_0_18_107/a_2724_472# 0.00308f
C13611 trim_val\[4\] FILLER_0_2_165/a_36_472# 0.007765f
C13612 FILLER_0_5_72/a_1468_375# _029_ 0.007876f
C13613 FILLER_0_5_72/a_124_375# trim_mask\[1\] 0.010758f
C13614 _016_ _129_ 0.002216f
C13615 FILLER_0_22_177/a_36_472# vss 0.002984f
C13616 FILLER_0_22_177/a_484_472# vdd 0.006974f
C13617 _112_ _001_ 0.002527f
C13618 _099_ _195_/a_255_603# 0.002146f
C13619 trimb[1] FILLER_0_18_2/a_1468_375# 0.002041f
C13620 _313_/a_67_603# _120_ 0.005873f
C13621 trim_val\[3\] _441_/a_2248_156# 0.027464f
C13622 _371_/a_36_113# vdd 0.007666f
C13623 _369_/a_36_68# _156_ 0.001359f
C13624 _426_/a_2248_156# net64 0.01109f
C13625 mask\[2\] FILLER_0_16_154/a_1020_375# 0.020485f
C13626 FILLER_0_4_107/a_36_472# _160_ 0.009073f
C13627 FILLER_0_4_213/a_36_472# vdd 0.087733f
C13628 FILLER_0_4_213/a_572_375# vss 0.017689f
C13629 _057_ _056_ 0.167928f
C13630 trim_val\[0\] _054_ 0.010002f
C13631 _418_/a_448_472# _007_ 0.050316f
C13632 _095_ _097_ 0.030222f
C13633 _255_/a_224_552# _311_/a_66_473# 0.002588f
C13634 _077_ net51 0.76967f
C13635 fanout79/a_36_160# net79 0.011193f
C13636 FILLER_0_22_86/a_572_375# _098_ 0.001139f
C13637 FILLER_0_7_72/a_1380_472# vss 0.001117f
C13638 _432_/a_36_151# FILLER_0_18_171/a_36_472# 0.059367f
C13639 FILLER_0_17_72/a_1468_375# _131_ 0.006871f
C13640 net20 _123_ 0.034801f
C13641 _136_ _451_/a_2449_156# 0.004653f
C13642 _367_/a_36_68# vss 0.001589f
C13643 ctln[3] _000_ 0.008418f
C13644 _449_/a_1000_472# vss 0.029565f
C13645 mask\[7\] _436_/a_36_151# 0.030028f
C13646 FILLER_0_21_286/a_484_472# net77 0.02147f
C13647 result[5] fanout61/a_36_113# 0.001866f
C13648 result[6] _421_/a_1000_472# 0.024206f
C13649 net73 FILLER_0_17_133/a_36_472# 0.049294f
C13650 net20 _073_ 0.437482f
C13651 _003_ vdd 0.032367f
C13652 net4 cal_itt\[0\] 0.054266f
C13653 ctln[1] _411_/a_1308_423# 0.037098f
C13654 fanout58/a_36_160# fanout59/a_36_160# 0.001216f
C13655 _059_ FILLER_0_8_156/a_124_375# 0.00593f
C13656 _253_/a_36_68# net19 0.019615f
C13657 net33 _023_ 0.015172f
C13658 _149_ _437_/a_2248_156# 0.031905f
C13659 _026_ _437_/a_1000_472# 0.042316f
C13660 FILLER_0_17_38/a_124_375# _452_/a_36_151# 0.006111f
C13661 vdd trim[3] 0.147228f
C13662 FILLER_0_4_197/a_572_375# _088_ 0.013597f
C13663 _372_/a_1602_69# _152_ 0.00262f
C13664 _083_ _081_ 0.03934f
C13665 _115_ net23 0.018953f
C13666 _451_/a_1040_527# _040_ 0.007154f
C13667 trim_val\[0\] vss 0.11063f
C13668 FILLER_0_14_181/a_124_375# _043_ 0.008393f
C13669 result[4] FILLER_0_17_282/a_36_472# 0.017375f
C13670 _123_ FILLER_0_6_231/a_572_375# 0.00487f
C13671 trimb[1] cal_count\[2\] 0.003178f
C13672 _057_ _068_ 0.393271f
C13673 _402_/a_718_527# vdd 0.020893f
C13674 net15 FILLER_0_6_47/a_1468_375# 0.007439f
C13675 net50 _444_/a_2248_156# 0.005539f
C13676 ctln[3] FILLER_0_0_266/a_36_472# 0.012298f
C13677 net41 _446_/a_1308_423# 0.056251f
C13678 _086_ _311_/a_2180_473# 0.001744f
C13679 net47 _450_/a_36_151# 0.029201f
C13680 _126_ _171_ 0.01633f
C13681 _128_ _315_/a_36_68# 0.04902f
C13682 FILLER_0_5_128/a_124_375# _370_/a_124_24# 0.023285f
C13683 fanout62/a_36_160# FILLER_0_11_282/a_124_375# 0.058702f
C13684 mask\[4\] FILLER_0_19_171/a_36_472# 0.001776f
C13685 ctln[2] clk 0.004558f
C13686 _196_/a_36_160# FILLER_0_14_263/a_36_472# 0.004828f
C13687 output23/a_224_472# mask\[7\] 0.046766f
C13688 FILLER_0_19_155/a_124_375# vdd 0.019233f
C13689 FILLER_0_13_206/a_124_375# vdd 0.034528f
C13690 sample vdd 0.154389f
C13691 ctlp[5] net22 0.001542f
C13692 _137_ FILLER_0_15_180/a_36_472# 0.004437f
C13693 _131_ _040_ 0.211618f
C13694 _028_ FILLER_0_7_72/a_1020_375# 0.003837f
C13695 net37 vdd 0.544653f
C13696 FILLER_0_24_63/a_124_375# output26/a_224_472# 0.00515f
C13697 _136_ net36 1.151311f
C13698 _445_/a_2665_112# vdd 0.055628f
C13699 FILLER_0_21_28/a_2724_472# vss -0.001553f
C13700 _432_/a_1308_423# _091_ 0.008903f
C13701 FILLER_0_3_221/a_1020_375# vss 0.003948f
C13702 FILLER_0_3_221/a_1468_375# vdd 0.008815f
C13703 FILLER_0_12_124/a_36_472# _114_ 0.003953f
C13704 _436_/a_796_472# vdd 0.005009f
C13705 _423_/a_2248_156# _012_ 0.011646f
C13706 net73 FILLER_0_18_107/a_124_375# 0.003742f
C13707 FILLER_0_9_223/a_484_472# _426_/a_2665_112# 0.004209f
C13708 net62 net36 0.034265f
C13709 cal_itt\[3\] _116_ 0.001364f
C13710 _403_/a_224_472# _183_ 0.007508f
C13711 net36 _438_/a_1000_472# 0.072117f
C13712 _126_ mask\[0\] 0.067513f
C13713 ctln[8] net52 0.005231f
C13714 net15 net50 0.177988f
C13715 _363_/a_36_68# _155_ 0.013915f
C13716 _053_ _081_ 0.698311f
C13717 _428_/a_2665_112# _427_/a_36_151# 0.028591f
C13718 _439_/a_1308_423# vss 0.009355f
C13719 net39 _063_ 0.004732f
C13720 FILLER_0_10_78/a_36_472# _439_/a_36_151# 0.00271f
C13721 result[8] FILLER_0_23_290/a_36_472# 0.001414f
C13722 _427_/a_2560_156# net23 0.042069f
C13723 FILLER_0_21_28/a_3260_375# _424_/a_36_151# 0.035849f
C13724 net63 FILLER_0_15_212/a_1020_375# 0.001012f
C13725 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_36_472# 0.007947f
C13726 FILLER_0_4_152/a_124_375# _066_ 0.003354f
C13727 _414_/a_1308_423# _053_ 0.029387f
C13728 net57 _058_ 0.028536f
C13729 _119_ vss 0.22921f
C13730 _070_ _121_ 0.285424f
C13731 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_124_375# 0.007947f
C13732 _021_ net57 0.00736f
C13733 net62 _193_/a_36_160# 0.00227f
C13734 FILLER_0_14_99/a_124_375# vdd 0.040312f
C13735 net81 calibrate 0.047274f
C13736 FILLER_0_12_136/a_1020_375# cal_count\[3\] 0.002916f
C13737 output31/a_224_472# FILLER_0_17_282/a_124_375# 0.002977f
C13738 net50 FILLER_0_6_90/a_572_375# 0.010099f
C13739 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_572_375# 0.001597f
C13740 _056_ _310_/a_49_472# 0.003286f
C13741 FILLER_0_12_2/a_572_375# vdd 0.022401f
C13742 FILLER_0_12_2/a_124_375# vss 0.002871f
C13743 net63 _434_/a_36_151# 0.005153f
C13744 _091_ _339_/a_36_160# 0.031941f
C13745 _326_/a_36_160# FILLER_0_9_105/a_484_472# 0.002647f
C13746 FILLER_0_10_247/a_124_375# net79 0.00498f
C13747 output25/a_224_472# vss 0.080847f
C13748 net81 FILLER_0_10_256/a_124_375# 0.026113f
C13749 fanout70/a_36_113# net36 0.007807f
C13750 FILLER_0_16_57/a_932_472# _176_ 0.010635f
C13751 result[7] _421_/a_1000_472# 0.015328f
C13752 net53 _451_/a_2449_156# 0.015332f
C13753 fanout74/a_36_113# net69 0.006779f
C13754 FILLER_0_4_152/a_124_375# net23 0.039975f
C13755 _414_/a_1204_472# _053_ 0.003935f
C13756 _326_/a_36_160# vss 0.002357f
C13757 net81 net21 0.185411f
C13758 FILLER_0_1_98/a_124_375# net52 0.001167f
C13759 ctlp[1] net19 0.029153f
C13760 net7 output16/a_224_472# 0.001321f
C13761 _432_/a_1000_472# net80 0.033803f
C13762 FILLER_0_9_28/a_2364_375# _453_/a_36_151# 0.001597f
C13763 _175_ _451_/a_3129_107# 0.021546f
C13764 _408_/a_728_93# cal_count\[0\] 0.007633f
C13765 _208_/a_36_160# vss 0.012188f
C13766 _139_ vdd 0.085044f
C13767 net62 FILLER_0_15_228/a_36_472# 0.002128f
C13768 _065_ vss 0.230397f
C13769 net55 _216_/a_255_603# 0.001011f
C13770 _370_/a_1152_472# _152_ 0.001423f
C13771 _028_ _077_ 0.017713f
C13772 cal_count\[3\] FILLER_0_12_20/a_124_375# 0.008038f
C13773 FILLER_0_4_123/a_124_375# FILLER_0_4_107/a_1468_375# 0.012001f
C13774 net69 FILLER_0_3_78/a_572_375# 0.002984f
C13775 _363_/a_36_68# _163_ 0.005627f
C13776 _413_/a_2560_156# net21 0.002416f
C13777 net60 _418_/a_2248_156# 0.045472f
C13778 net69 FILLER_0_2_127/a_124_375# 0.08337f
C13779 result[2] _044_ 0.393081f
C13780 fanout58/a_36_160# net5 0.003758f
C13781 net41 _408_/a_1336_472# 0.063099f
C13782 result[6] net18 0.026875f
C13783 fanout74/a_36_113# _152_ 0.017267f
C13784 FILLER_0_4_49/a_124_375# trim_val\[1\] 0.024557f
C13785 trim_val\[2\] _166_ 0.014514f
C13786 trim_mask\[2\] _160_ 0.367302f
C13787 _127_ _395_/a_36_488# 0.00519f
C13788 ctlp[5] vdd 0.293399f
C13789 FILLER_0_8_127/a_124_375# _125_ 0.003105f
C13790 net63 FILLER_0_15_205/a_36_472# 0.047903f
C13791 net62 _417_/a_2248_156# 0.005537f
C13792 net32 _419_/a_1308_423# 0.00191f
C13793 _009_ _109_ 0.006736f
C13794 net53 net36 3.423337f
C13795 _086_ _125_ 0.490983f
C13796 FILLER_0_5_109/a_124_375# _163_ 0.002658f
C13797 _274_/a_2552_68# _070_ 0.001238f
C13798 FILLER_0_9_282/a_572_375# vdd 0.002928f
C13799 FILLER_0_9_282/a_124_375# vss 0.00451f
C13800 FILLER_0_6_47/a_932_472# vdd 0.003435f
C13801 net15 FILLER_0_15_72/a_484_472# 0.002925f
C13802 mask\[4\] _104_ 0.001621f
C13803 net35 FILLER_0_22_107/a_572_375# 0.010438f
C13804 mask\[8\] FILLER_0_22_107/a_36_472# 0.017159f
C13805 output24/a_224_472# vss 0.004078f
C13806 fanout59/a_36_160# net18 0.003981f
C13807 FILLER_0_2_101/a_124_375# _157_ 0.002818f
C13808 net63 FILLER_0_22_177/a_484_472# 0.059367f
C13809 mask\[4\] vss 0.426009f
C13810 _402_/a_728_93# _179_ 0.011717f
C13811 _431_/a_3041_156# vss 0.001312f
C13812 _322_/a_848_380# _118_ 0.047787f
C13813 net33 _297_/a_36_472# 0.00521f
C13814 FILLER_0_13_212/a_1468_375# vdd -0.013698f
C13815 FILLER_0_13_212/a_1020_375# vss 0.041631f
C13816 _412_/a_448_472# cal_itt\[1\] 0.043203f
C13817 net72 _423_/a_36_151# 0.024965f
C13818 FILLER_0_12_136/a_1468_375# _114_ 0.006974f
C13819 ctlp[1] _420_/a_36_151# 0.067975f
C13820 net34 _422_/a_36_151# 0.032272f
C13821 _098_ _146_ 0.004276f
C13822 FILLER_0_11_101/a_484_472# _120_ 0.011393f
C13823 _421_/a_2248_156# vdd 0.035239f
C13824 FILLER_0_20_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001543f
C13825 FILLER_0_10_214/a_36_472# vss 0.008006f
C13826 net19 cal_itt\[1\] 0.044717f
C13827 _415_/a_1308_423# vdd 0.004258f
C13828 _106_ mask\[2\] 0.039965f
C13829 net20 _189_/a_67_603# 0.011939f
C13830 net35 _023_ 0.008361f
C13831 fanout50/a_36_160# net52 0.037383f
C13832 result[8] FILLER_0_24_274/a_932_472# 0.005458f
C13833 FILLER_0_19_187/a_572_375# vdd 0.023383f
C13834 _413_/a_36_151# FILLER_0_3_172/a_2276_472# 0.001723f
C13835 vss FILLER_0_21_60/a_36_472# 0.001384f
C13836 vdd FILLER_0_21_60/a_484_472# 0.005181f
C13837 net26 FILLER_0_23_44/a_932_472# 0.001889f
C13838 mask\[0\] state\[1\] 0.064758f
C13839 _411_/a_1308_423# net65 0.004122f
C13840 _305_/a_36_159# net76 0.010842f
C13841 FILLER_0_9_223/a_484_472# _223_/a_36_160# 0.004695f
C13842 FILLER_0_16_107/a_572_375# _136_ 0.006445f
C13843 net56 fanout56/a_36_113# 0.015924f
C13844 _429_/a_1308_423# net22 0.001856f
C13845 FILLER_0_2_111/a_1020_375# vdd 0.007918f
C13846 net41 FILLER_0_16_37/a_124_375# 0.008195f
C13847 _429_/a_448_472# _018_ 0.035489f
C13848 fanout82/a_36_113# vss 0.023533f
C13849 _093_ FILLER_0_17_104/a_484_472# 0.014431f
C13850 net41 _444_/a_1308_423# 0.015841f
C13851 FILLER_0_4_91/a_124_375# _160_ 0.009765f
C13852 _173_ _186_ 0.002111f
C13853 net15 _394_/a_1336_472# 0.01144f
C13854 result[8] net33 0.474056f
C13855 fanout50/a_36_160# net49 0.030626f
C13856 FILLER_0_11_109/a_124_375# _134_ 0.027704f
C13857 _445_/a_36_151# net47 0.002364f
C13858 net41 FILLER_0_8_24/a_572_375# 0.003909f
C13859 _440_/a_1308_423# vdd 0.00218f
C13860 _440_/a_448_472# vss 0.032037f
C13861 net81 net80 0.006516f
C13862 net18 _418_/a_36_151# 0.017941f
C13863 net64 _098_ 0.281888f
C13864 _325_/a_224_472# _118_ 0.004845f
C13865 result[7] net18 0.098317f
C13866 cal net4 0.026084f
C13867 _390_/a_36_68# vdd 0.012472f
C13868 net82 _443_/a_36_151# 0.03565f
C13869 _115_ _439_/a_2248_156# 0.003553f
C13870 _412_/a_2248_156# en 0.022108f
C13871 FILLER_0_21_286/a_124_375# net18 0.015582f
C13872 net70 FILLER_0_14_107/a_572_375# 0.018214f
C13873 FILLER_0_5_72/a_1380_472# vss 0.004538f
C13874 result[5] net79 0.036275f
C13875 _087_ net76 0.529571f
C13876 FILLER_0_20_2/a_124_375# vss 0.002737f
C13877 FILLER_0_20_2/a_572_375# vdd 0.010844f
C13878 _098_ FILLER_0_19_171/a_1380_472# 0.001764f
C13879 FILLER_0_5_54/a_36_472# trim_mask\[1\] 0.101342f
C13880 FILLER_0_5_54/a_1380_472# _029_ 0.01027f
C13881 FILLER_0_8_138/a_36_472# _119_ 0.003894f
C13882 _057_ _113_ 0.339862f
C13883 FILLER_0_21_125/a_484_472# _022_ 0.004649f
C13884 FILLER_0_16_107/a_124_375# _131_ 0.016011f
C13885 _028_ _363_/a_692_472# 0.001416f
C13886 _028_ net50 0.087995f
C13887 ctlp[1] _419_/a_448_472# 0.020153f
C13888 net81 mask\[1\] 2.509493f
C13889 _446_/a_2560_156# net40 0.012204f
C13890 mask\[8\] _433_/a_36_151# 0.001402f
C13891 _448_/a_448_472# net65 0.001006f
C13892 _426_/a_36_151# FILLER_0_8_247/a_1380_472# 0.001723f
C13893 _070_ FILLER_0_10_94/a_484_472# 0.003573f
C13894 _130_ vss 0.090346f
C13895 _304_/a_224_472# _013_ 0.002769f
C13896 FILLER_0_5_198/a_572_375# net37 0.009149f
C13897 vss _034_ 0.008249f
C13898 mask\[5\] FILLER_0_19_171/a_572_375# 0.007169f
C13899 _161_ vss 0.134214f
C13900 fanout60/a_36_160# net60 0.019034f
C13901 en net4 0.125535f
C13902 _421_/a_2560_156# net19 0.006572f
C13903 _430_/a_36_151# FILLER_0_18_209/a_484_472# 0.001043f
C13904 FILLER_0_12_2/a_484_472# _450_/a_36_151# 0.059367f
C13905 fanout64/a_36_160# net64 0.043709f
C13906 net27 net79 0.059863f
C13907 _077_ FILLER_0_9_223/a_36_472# 0.005511f
C13908 _430_/a_2560_156# _092_ 0.001333f
C13909 _105_ net78 0.004705f
C13910 FILLER_0_13_206/a_36_472# _043_ 0.011439f
C13911 _442_/a_2248_156# _157_ 0.002731f
C13912 _033_ FILLER_0_6_37/a_124_375# 0.018812f
C13913 _164_ FILLER_0_6_47/a_572_375# 0.010099f
C13914 _129_ vss 0.141494f
C13915 _086_ net76 0.049988f
C13916 _069_ FILLER_0_13_206/a_124_375# 0.009695f
C13917 _133_ calibrate 0.0188f
C13918 _070_ _122_ 0.153373f
C13919 net51 _039_ 0.398642f
C13920 FILLER_0_16_255/a_36_472# _287_/a_36_472# 0.004546f
C13921 result[9] FILLER_0_14_263/a_124_375# 0.003706f
C13922 result[9] _010_ 0.121471f
C13923 _053_ _155_ 0.122798f
C13924 net5 net18 0.015361f
C13925 _447_/a_36_151# net69 0.001216f
C13926 net49 FILLER_0_3_54/a_36_472# 0.00186f
C13927 FILLER_0_4_152/a_124_375# net57 0.001947f
C13928 _070_ FILLER_0_7_233/a_124_375# 0.004917f
C13929 _115_ _315_/a_244_497# 0.00153f
C13930 _128_ net4 0.039671f
C13931 net1 input4/a_36_68# 0.056389f
C13932 _028_ FILLER_0_5_72/a_572_375# 0.00123f
C13933 _408_/a_728_93# net17 0.005494f
C13934 FILLER_0_15_150/a_124_375# _427_/a_2248_156# 0.001221f
C13935 output10/a_224_472# FILLER_0_0_232/a_124_375# 0.00363f
C13936 net52 net14 0.072003f
C13937 _059_ FILLER_0_5_148/a_36_472# 0.010977f
C13938 fanout81/a_36_160# net2 0.044793f
C13939 _070_ _227_/a_36_160# 0.00254f
C13940 _077_ net74 0.025882f
C13941 _072_ state\[2\] 0.002629f
C13942 _052_ FILLER_0_21_28/a_1916_375# 0.002388f
C13943 FILLER_0_7_72/a_3260_375# _058_ 0.00258f
C13944 _070_ _169_ 0.006335f
C13945 net58 net59 0.066534f
C13946 FILLER_0_18_37/a_1468_375# vdd 0.021186f
C13947 net75 _316_/a_124_24# 0.003078f
C13948 _317_/a_36_113# calibrate 0.011799f
C13949 mask\[3\] FILLER_0_17_161/a_36_472# 0.13873f
C13950 _429_/a_448_472# vss 0.035246f
C13951 net49 net14 0.00344f
C13952 net52 _164_ 0.313379f
C13953 net63 _139_ 0.003073f
C13954 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_36_472# 0.086742f
C13955 FILLER_0_16_73/a_36_472# vdd 0.08735f
C13956 _063_ net47 0.142088f
C13957 FILLER_0_14_99/a_36_472# _043_ 0.001242f
C13958 ctln[1] ctln[3] 0.926618f
C13959 net8 vdd 0.593788f
C13960 vss result[3] 0.28152f
C13961 _037_ net22 0.079675f
C13962 net62 _416_/a_36_151# 0.054002f
C13963 net45 net26 0.002978f
C13964 FILLER_0_15_142/a_484_472# net23 0.002884f
C13965 FILLER_0_16_57/a_932_472# FILLER_0_17_64/a_124_375# 0.001723f
C13966 net49 _164_ 0.428468f
C13967 FILLER_0_3_2/a_124_375# net66 0.027628f
C13968 FILLER_0_21_142/a_484_472# vdd 0.004917f
C13969 ctln[5] _448_/a_1308_423# 0.004061f
C13970 net31 net32 0.023293f
C13971 result[9] FILLER_0_23_282/a_36_472# 0.001324f
C13972 net16 FILLER_0_12_28/a_124_375# 0.002225f
C13973 _096_ vss 0.126096f
C13974 net1 _001_ 0.300335f
C13975 ctln[1] net5 0.050549f
C13976 _021_ _141_ 0.047816f
C13977 _394_/a_1936_472# vss 0.006085f
C13978 _082_ net59 0.004251f
C13979 FILLER_0_7_195/a_36_472# _062_ 0.0045f
C13980 net82 net59 0.102279f
C13981 _053_ _163_ 0.763235f
C13982 trim_mask\[1\] FILLER_0_6_79/a_36_472# 0.006265f
C13983 _122_ FILLER_0_5_164/a_572_375# 0.001352f
C13984 _310_/a_49_472# _113_ 0.020387f
C13985 _176_ _315_/a_36_68# 0.003811f
C13986 vss FILLER_0_22_107/a_124_375# 0.002881f
C13987 vdd FILLER_0_22_107/a_572_375# 0.005745f
C13988 _423_/a_36_151# FILLER_0_23_60/a_124_375# 0.005577f
C13989 _181_ vdd 0.209604f
C13990 FILLER_0_20_169/a_124_375# FILLER_0_19_171/a_36_472# 0.001543f
C13991 fanout57/a_36_113# net59 0.00178f
C13992 FILLER_0_15_150/a_36_472# net23 0.010444f
C13993 result[4] vss 0.306116f
C13994 net50 net47 0.040157f
C13995 FILLER_0_10_37/a_124_375# net68 0.012617f
C13996 net15 net72 0.157843f
C13997 net72 FILLER_0_21_28/a_1020_375# 0.040811f
C13998 net81 output48/a_224_472# 0.040059f
C13999 net47 _382_/a_224_472# 0.001795f
C14000 _114_ _308_/a_1084_68# 0.00178f
C14001 FILLER_0_9_28/a_484_472# _054_ 0.002831f
C14002 net16 FILLER_0_17_38/a_124_375# 0.046435f
C14003 net58 net64 0.590523f
C14004 _320_/a_36_472# net79 0.029189f
C14005 FILLER_0_5_164/a_124_375# _163_ 0.048663f
C14006 _068_ _311_/a_3220_473# 0.004371f
C14007 FILLER_0_21_142/a_36_472# vss 0.009084f
C14008 FILLER_0_2_93/a_124_375# net69 0.015032f
C14009 net15 FILLER_0_5_54/a_484_472# 0.002186f
C14010 _425_/a_448_472# _122_ 0.002863f
C14011 _425_/a_1308_423# calibrate 0.022697f
C14012 _065_ _036_ 0.031728f
C14013 FILLER_0_8_24/a_36_472# net17 0.045619f
C14014 _140_ _434_/a_36_151# 0.025956f
C14015 _424_/a_1204_472# _012_ 0.003572f
C14016 mask\[5\] FILLER_0_20_177/a_1468_375# 0.013222f
C14017 net81 mask\[0\] 0.320022f
C14018 net62 FILLER_0_14_235/a_484_472# 0.017862f
C14019 _033_ _444_/a_1204_472# 0.002294f
C14020 _023_ vdd 0.062542f
C14021 _412_/a_1000_472# net1 0.027748f
C14022 _174_ cal_count\[0\] 0.009645f
C14023 _024_ _435_/a_36_151# 0.10993f
C14024 _417_/a_1308_423# vss 0.002064f
C14025 net9 net8 0.027272f
C14026 _232_/a_67_603# vss 0.00988f
C14027 _306_/a_36_68# _116_ 0.00183f
C14028 FILLER_0_20_98/a_124_375# vdd 0.0135f
C14029 _035_ net16 0.034977f
C14030 FILLER_0_10_214/a_124_375# _055_ 0.001419f
C14031 FILLER_0_4_123/a_36_472# vss 0.004542f
C14032 net82 _122_ 0.001375f
C14033 result[8] net35 0.001362f
C14034 net63 FILLER_0_19_187/a_572_375# 0.049706f
C14035 _127_ vdd 0.155954f
C14036 output34/a_224_472# net30 0.002189f
C14037 _056_ vss 0.193804f
C14038 FILLER_0_5_72/a_572_375# net47 0.006974f
C14039 _385_/a_244_472# net37 0.001593f
C14040 net35 FILLER_0_22_86/a_36_472# 0.00797f
C14041 mask\[8\] FILLER_0_22_86/a_484_472# 0.012439f
C14042 FILLER_0_4_197/a_1020_375# net76 0.006026f
C14043 FILLER_0_5_212/a_124_375# _078_ 0.002018f
C14044 FILLER_0_7_59/a_484_472# vss 0.005804f
C14045 FILLER_0_17_226/a_36_472# _291_/a_36_160# 0.035111f
C14046 _453_/a_448_472# vdd 0.010005f
C14047 _453_/a_36_151# vss 0.007105f
C14048 FILLER_0_13_212/a_36_472# _043_ 0.011752f
C14049 _247_/a_36_160# _062_ 0.011327f
C14050 net35 FILLER_0_22_128/a_2724_472# 0.012359f
C14051 _015_ _426_/a_36_151# 0.01243f
C14052 FILLER_0_10_78/a_1380_472# _114_ 0.011079f
C14053 _114_ _136_ 0.003405f
C14054 trim_val\[2\] net17 0.019133f
C14055 _017_ cal_count\[3\] 0.003939f
C14056 net57 _267_/a_672_472# 0.004637f
C14057 _037_ vdd 0.158731f
C14058 FILLER_0_12_2/a_36_472# net67 0.013281f
C14059 _397_/a_36_472# vdd 0.094023f
C14060 net68 FILLER_0_6_47/a_1380_472# 0.049638f
C14061 FILLER_0_11_135/a_36_472# vdd 0.091206f
C14062 FILLER_0_11_135/a_124_375# vss 0.02843f
C14063 output31/a_224_472# vdd 0.083516f
C14064 _075_ _056_ 0.001957f
C14065 net17 FILLER_0_23_44/a_36_472# 0.071244f
C14066 _114_ FILLER_0_13_142/a_124_375# 0.00191f
C14067 mask\[8\] _050_ 0.001479f
C14068 _098_ _097_ 0.034041f
C14069 _064_ _033_ 0.001986f
C14070 _098_ _437_/a_1308_423# 0.005568f
C14071 _274_/a_716_497# net64 0.007904f
C14072 net60 _419_/a_3041_156# 0.001022f
C14073 net20 FILLER_0_12_220/a_932_472# 0.007397f
C14074 net55 FILLER_0_18_61/a_36_472# 0.022296f
C14075 _091_ FILLER_0_18_177/a_1020_375# 0.002226f
C14076 FILLER_0_9_60/a_484_472# FILLER_0_9_72/a_36_472# 0.002296f
C14077 FILLER_0_8_138/a_36_472# _129_ 0.055537f
C14078 net32 _421_/a_36_151# 0.008275f
C14079 net81 FILLER_0_15_212/a_124_375# 0.005049f
C14080 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_124_375# 0.012001f
C14081 _077_ _439_/a_1204_472# 0.016471f
C14082 net81 _099_ 0.140011f
C14083 _448_/a_1308_423# net59 0.014899f
C14084 _039_ clkc 0.003104f
C14085 FILLER_0_21_133/a_124_375# vdd 0.010519f
C14086 FILLER_0_11_101/a_572_375# vss 0.055325f
C14087 FILLER_0_11_101/a_36_472# vdd 0.093852f
C14088 _150_ _438_/a_36_151# 0.032532f
C14089 _068_ vss 0.547532f
C14090 _093_ FILLER_0_18_100/a_124_375# 0.011632f
C14091 FILLER_0_18_2/a_3260_375# net40 0.035372f
C14092 output32/a_224_472# net32 0.014826f
C14093 FILLER_0_18_107/a_36_472# FILLER_0_17_104/a_484_472# 0.026657f
C14094 FILLER_0_13_212/a_1020_375# FILLER_0_12_220/a_124_375# 0.05841f
C14095 _033_ net42 0.002707f
C14096 _052_ _424_/a_448_472# 0.017551f
C14097 FILLER_0_4_152/a_124_375# FILLER_0_5_148/a_572_375# 0.05841f
C14098 FILLER_0_15_180/a_484_472# vss 0.001207f
C14099 mask\[1\] FILLER_0_15_180/a_572_375# 0.011186f
C14100 FILLER_0_4_99/a_36_472# _160_ 0.006222f
C14101 state\[0\] _091_ 0.012343f
C14102 mask\[8\] _214_/a_36_160# 0.001264f
C14103 _432_/a_448_472# _136_ 0.001892f
C14104 _395_/a_36_488# _116_ 0.033784f
C14105 mask\[5\] _108_ 0.036539f
C14106 FILLER_0_4_107/a_124_375# _157_ 0.001427f
C14107 FILLER_0_10_78/a_1380_472# _176_ 0.009351f
C14108 _176_ _136_ 0.114837f
C14109 _431_/a_36_151# vdd 0.145005f
C14110 _132_ FILLER_0_18_107/a_932_472# 0.001369f
C14111 _093_ FILLER_0_17_72/a_572_375# 0.005609f
C14112 _018_ _138_ 0.008093f
C14113 _075_ _068_ 0.006297f
C14114 _098_ mask\[2\] 0.06158f
C14115 comp FILLER_0_12_2/a_36_472# 0.003875f
C14116 net34 _435_/a_1000_472# 0.007444f
C14117 FILLER_0_7_195/a_124_375# vdd 0.007788f
C14118 trimb[4] cal_count\[2\] 0.146942f
C14119 vdd FILLER_0_13_72/a_36_472# 0.108152f
C14120 vss FILLER_0_13_72/a_572_375# 0.061657f
C14121 fanout51/a_36_113# vss 0.0844f
C14122 net68 _440_/a_796_472# 0.021463f
C14123 _127_ _135_ 0.00622f
C14124 _345_/a_36_160# vdd 0.100094f
C14125 cal_itt\[3\] net47 0.00247f
C14126 result[8] net22 0.278936f
C14127 FILLER_0_19_142/a_36_472# _145_ 0.010377f
C14128 FILLER_0_18_171/a_36_472# net80 0.041571f
C14129 _086_ _267_/a_1568_472# 0.002143f
C14130 FILLER_0_20_169/a_124_375# vss 0.017635f
C14131 FILLER_0_20_169/a_36_472# vdd 0.010522f
C14132 _025_ _437_/a_2665_112# 0.001245f
C14133 _188_ _453_/a_796_472# 0.00103f
C14134 output47/a_224_472# net3 0.002186f
C14135 trimb[4] input3/a_36_113# 0.001221f
C14136 _443_/a_2248_156# _386_/a_124_24# 0.001257f
C14137 _432_/a_36_151# _097_ 0.003144f
C14138 mask\[4\] _346_/a_49_472# 0.079347f
C14139 _097_ FILLER_0_15_180/a_124_375# 0.007065f
C14140 _274_/a_36_68# net4 0.037848f
C14141 net20 ctlp[1] 0.024556f
C14142 FILLER_0_17_38/a_124_375# _041_ 0.009172f
C14143 _328_/a_36_113# net74 0.002214f
C14144 FILLER_0_17_72/a_2276_472# net36 0.004399f
C14145 _099_ net30 0.05959f
C14146 _142_ FILLER_0_17_142/a_36_472# 0.011216f
C14147 _053_ FILLER_0_7_104/a_1020_375# 0.002671f
C14148 FILLER_0_14_50/a_124_375# _174_ 0.033245f
C14149 _093_ _438_/a_2665_112# 0.003293f
C14150 net69 vss 0.34555f
C14151 _442_/a_2248_156# _158_ 0.001288f
C14152 vss _201_/a_67_603# 0.012925f
C14153 mask\[9\] _438_/a_2248_156# 0.036436f
C14154 _064_ _446_/a_36_151# 0.006723f
C14155 _114_ net53 0.001275f
C14156 _126_ _131_ 0.626666f
C14157 trim[1] net40 0.043114f
C14158 _413_/a_36_151# _079_ 0.0017f
C14159 _415_/a_1204_472# result[1] 0.004051f
C14160 net52 _442_/a_796_472# 0.004871f
C14161 _259_/a_455_68# _076_ 0.002372f
C14162 FILLER_0_18_177/a_1380_472# vdd 0.005692f
C14163 FILLER_0_18_177/a_932_472# vss -0.001894f
C14164 net47 _039_ 0.042757f
C14165 FILLER_0_18_171/a_124_375# _091_ 0.034351f
C14166 _005_ _416_/a_448_472# 0.04044f
C14167 ctln[2] FILLER_0_0_266/a_36_472# 0.049163f
C14168 _115_ FILLER_0_10_107/a_572_375# 0.040198f
C14169 fanout53/a_36_160# FILLER_0_16_154/a_484_472# 0.014774f
C14170 FILLER_0_9_60/a_124_375# vdd 0.005798f
C14171 _450_/a_1284_156# _039_ 0.001226f
C14172 _450_/a_3129_107# cal_count\[0\] 0.020971f
C14173 net15 FILLER_0_23_60/a_124_375# 0.038706f
C14174 FILLER_0_19_28/a_572_375# _452_/a_36_151# 0.0027f
C14175 net69 _441_/a_2248_156# 0.036635f
C14176 output20/a_224_472# _422_/a_448_472# 0.009204f
C14177 output21/a_224_472# ctlp[3] 0.021951f
C14178 net65 net5 0.004409f
C14179 net20 _079_ 0.177911f
C14180 FILLER_0_17_218/a_124_375# vdd 0.00593f
C14181 _100_ vdd 0.212037f
C14182 FILLER_0_18_2/a_3172_472# net55 0.00602f
C14183 _425_/a_1204_472# vdd 0.015969f
C14184 net73 FILLER_0_18_107/a_3172_472# 0.00533f
C14185 _152_ vss 0.140215f
C14186 mask\[7\] FILLER_0_22_128/a_1380_472# 0.015814f
C14187 _432_/a_36_151# mask\[2\] 0.031341f
C14188 _069_ _429_/a_1308_423# 0.027468f
C14189 net37 FILLER_0_6_231/a_484_472# 0.004323f
C14190 _115_ FILLER_0_9_142/a_36_472# 0.00336f
C14191 _297_/a_36_472# vdd 0.042391f
C14192 net53 _427_/a_2248_156# 0.038716f
C14193 trim_mask\[0\] vdd 0.154098f
C14194 net64 FILLER_0_9_270/a_484_472# 0.017924f
C14195 _002_ FILLER_0_3_172/a_3172_472# 0.002313f
C14196 output28/a_224_472# fanout79/a_36_160# 0.022393f
C14197 _067_ FILLER_0_12_20/a_484_472# 0.011046f
C14198 _147_ _208_/a_36_160# 0.006056f
C14199 result[5] net19 0.003542f
C14200 _423_/a_36_151# FILLER_0_23_44/a_124_375# 0.059049f
C14201 _394_/a_56_524# FILLER_0_15_59/a_572_375# 0.003413f
C14202 _448_/a_2248_156# net22 0.07925f
C14203 net15 FILLER_0_17_72/a_572_375# 0.003021f
C14204 _098_ FILLER_0_15_212/a_572_375# 0.009099f
C14205 _060_ net22 0.533421f
C14206 _428_/a_1000_472# net74 0.00735f
C14207 _176_ net53 0.083005f
C14208 fanout82/a_36_113# output37/a_224_472# 0.023409f
C14209 net52 _439_/a_2665_112# 0.00117f
C14210 _008_ vdd 0.284571f
C14211 _079_ FILLER_0_6_231/a_572_375# 0.002768f
C14212 _104_ result[9] 0.169685f
C14213 _093_ net35 0.00127f
C14214 _138_ vss 0.006962f
C14215 mask\[8\] mask\[9\] 0.078756f
C14216 FILLER_0_4_49/a_484_472# vdd 0.003356f
C14217 FILLER_0_4_49/a_36_472# vss 0.001931f
C14218 net54 _438_/a_2665_112# 0.032855f
C14219 _115_ _128_ 0.263909f
C14220 _256_/a_716_497# calibrate 0.001066f
C14221 net20 FILLER_0_24_274/a_124_375# 0.002751f
C14222 result[9] vss 0.348416f
C14223 mask\[4\] _106_ 0.091207f
C14224 output20/a_224_472# _108_ 0.022243f
C14225 result[8] vdd 0.590386f
C14226 net27 net19 0.036883f
C14227 net31 _421_/a_2665_112# 0.005428f
C14228 FILLER_0_18_2/a_3172_472# net17 0.002402f
C14229 _096_ _095_ 0.086147f
C14230 FILLER_0_3_204/a_36_472# vss 0.003572f
C14231 _176_ FILLER_0_10_107/a_484_472# 0.009571f
C14232 FILLER_0_22_86/a_36_472# vdd -0.001506f
C14233 FILLER_0_22_86/a_1468_375# vss 0.013146f
C14234 trim_val\[4\] _387_/a_36_113# 0.005339f
C14235 FILLER_0_11_78/a_484_472# _120_ 0.016839f
C14236 _038_ FILLER_0_11_78/a_484_472# 0.001782f
C14237 _114_ _311_/a_1660_473# 0.003304f
C14238 FILLER_0_22_128/a_2724_472# vdd 0.005923f
C14239 FILLER_0_22_128/a_2276_472# vss 0.02979f
C14240 FILLER_0_9_28/a_2364_375# _042_ 0.001216f
C14241 FILLER_0_9_28/a_36_472# vdd 0.086674f
C14242 _053_ net48 0.003159f
C14243 _132_ _428_/a_36_151# 0.013691f
C14244 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_572_375# 0.086635f
C14245 _236_/a_36_160# net67 0.009332f
C14246 net56 FILLER_0_18_139/a_932_472# 0.011079f
C14247 net31 output33/a_224_472# 0.005087f
C14248 net59 net21 0.157689f
C14249 output38/a_224_472# _446_/a_36_151# 0.117966f
C14250 ctlp[0] net17 0.006778f
C14251 _211_/a_36_160# vss 0.002041f
C14252 _013_ vss 0.163674f
C14253 _445_/a_796_472# _034_ 0.009261f
C14254 _116_ net22 0.122052f
C14255 FILLER_0_0_198/a_124_375# net21 0.004256f
C14256 output45/a_224_472# vss 0.00543f
C14257 net36 FILLER_0_18_76/a_36_472# 0.001728f
C14258 net82 FILLER_0_3_172/a_932_472# 0.007986f
C14259 FILLER_0_8_263/a_124_375# vdd 0.032664f
C14260 output8/a_224_472# net59 0.00398f
C14261 net54 net35 0.114666f
C14262 _124_ FILLER_0_10_107/a_484_472# 0.00438f
C14263 FILLER_0_24_130/a_36_472# output24/a_224_472# 0.023414f
C14264 en_co_clk FILLER_0_13_100/a_124_375# 0.002325f
C14265 vdd FILLER_0_14_235/a_124_375# -0.011193f
C14266 ctlp[5] _140_ 0.002123f
C14267 _020_ net36 0.001995f
C14268 _064_ _447_/a_36_151# 0.004185f
C14269 FILLER_0_3_172/a_36_472# net65 0.014671f
C14270 cal_itt\[2\] _084_ 0.061303f
C14271 _098_ FILLER_0_15_205/a_124_375# 0.009558f
C14272 _446_/a_2248_156# vdd 0.059236f
C14273 _322_/a_848_380# net74 0.00168f
C14274 net20 _256_/a_244_497# 0.005033f
C14275 _173_ _039_ 0.0326f
C14276 _035_ trim[0] 0.171633f
C14277 result[1] net18 0.056799f
C14278 _210_/a_67_603# vdd 0.028101f
C14279 _127_ _069_ 0.048146f
C14280 _415_/a_36_151# FILLER_0_10_256/a_124_375# 0.035117f
C14281 _091_ net79 0.052824f
C14282 calibrate _122_ 0.074949f
C14283 _132_ FILLER_0_11_109/a_36_472# 0.005748f
C14284 _116_ _311_/a_2700_473# 0.001555f
C14285 _443_/a_1308_423# vss 0.031091f
C14286 _412_/a_1000_472# net76 0.024114f
C14287 FILLER_0_14_99/a_124_375# _451_/a_36_151# 0.001441f
C14288 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3260_375# 0.086635f
C14289 FILLER_0_7_72/a_1916_375# _053_ 0.013335f
C14290 calibrate FILLER_0_7_233/a_124_375# 0.011958f
C14291 fanout67/a_36_160# FILLER_0_9_60/a_124_375# 0.02985f
C14292 _076_ _055_ 0.056585f
C14293 FILLER_0_12_136/a_484_472# net23 0.002172f
C14294 _119_ _375_/a_36_68# 0.007338f
C14295 _431_/a_2248_156# net56 0.013627f
C14296 _093_ net22 0.041918f
C14297 net20 FILLER_0_13_212/a_484_472# 0.001273f
C14298 net48 _425_/a_36_151# 0.020568f
C14299 _448_/a_2248_156# vdd 0.008296f
C14300 net52 FILLER_0_6_47/a_2724_472# 0.011079f
C14301 net64 calibrate 0.096329f
C14302 FILLER_0_16_107/a_484_472# vss 0.004223f
C14303 _444_/a_1308_423# FILLER_0_8_24/a_36_472# 0.009119f
C14304 net15 net35 0.01797f
C14305 _143_ _339_/a_36_160# 0.00507f
C14306 _122_ net21 0.026632f
C14307 _060_ vdd 0.349556f
C14308 _113_ vss 0.147905f
C14309 _165_ _164_ 0.351097f
C14310 calibrate _169_ 0.001883f
C14311 _392_/a_36_68# _067_ 0.020085f
C14312 _423_/a_36_151# vdd 0.088377f
C14313 fanout66/a_36_113# net68 0.01746f
C14314 FILLER_0_22_177/a_124_375# _023_ 0.001195f
C14315 FILLER_0_4_197/a_1468_375# _088_ 0.012367f
C14316 clk net59 0.052607f
C14317 FILLER_0_18_2/a_484_472# net38 0.003391f
C14318 FILLER_0_5_54/a_484_472# net47 0.006652f
C14319 net68 _453_/a_1308_423# 0.002195f
C14320 net57 _428_/a_796_472# 0.003017f
C14321 net72 _012_ 0.002382f
C14322 FILLER_0_3_54/a_36_472# net40 0.069702f
C14323 ctlp[1] _009_ 0.085933f
C14324 net62 output29/a_224_472# 0.138536f
C14325 _217_/a_36_160# _052_ 0.016695f
C14326 net74 _372_/a_1194_69# 0.002006f
C14327 FILLER_0_16_89/a_1468_375# _136_ 0.005791f
C14328 ctlp[7] _025_ 0.007483f
C14329 _343_/a_49_472# vdd 0.089707f
C14330 _242_/a_36_160# FILLER_0_5_164/a_36_472# 0.193804f
C14331 _044_ FILLER_0_14_263/a_124_375# 0.001047f
C14332 _126_ FILLER_0_11_101/a_124_375# 0.011403f
C14333 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_36_472# 0.012267f
C14334 _431_/a_1308_423# _136_ 0.027758f
C14335 fanout81/a_36_160# cal_itt\[1\] 0.069457f
C14336 _126_ _076_ 0.005517f
C14337 _187_ _392_/a_36_68# 0.058263f
C14338 FILLER_0_14_81/a_124_375# _451_/a_3129_107# 0.009542f
C14339 FILLER_0_17_72/a_3260_375# vss 0.052993f
C14340 FILLER_0_17_72/a_36_472# vdd 0.111688f
C14341 _134_ FILLER_0_10_107/a_572_375# 0.047331f
C14342 _048_ _204_/a_67_603# 0.004547f
C14343 _136_ FILLER_0_17_142/a_572_375# 0.001371f
C14344 cal_itt\[3\] _079_ 0.015743f
C14345 _064_ _444_/a_36_151# 0.001296f
C14346 result[5] _419_/a_448_472# 0.00232f
C14347 _148_ _025_ 0.007252f
C14348 FILLER_0_4_107/a_1380_472# vss 0.004455f
C14349 vss FILLER_0_6_37/a_124_375# 0.030885f
C14350 vdd FILLER_0_6_37/a_36_472# 0.138008f
C14351 _183_ _182_ 0.002134f
C14352 _370_/a_848_380# net23 0.001196f
C14353 result[6] FILLER_0_21_286/a_484_472# 0.011149f
C14354 _132_ FILLER_0_17_104/a_572_375# 0.003857f
C14355 _427_/a_1308_423# vss 0.030292f
C14356 net72 FILLER_0_15_59/a_484_472# 0.008749f
C14357 net17 _450_/a_3129_107# 0.004255f
C14358 net52 FILLER_0_2_111/a_932_472# 0.061249f
C14359 _043_ FILLER_0_13_72/a_484_472# 0.016114f
C14360 net41 _402_/a_56_567# 0.021641f
C14361 _132_ _148_ 0.002873f
C14362 _091_ _429_/a_2560_156# 0.001502f
C14363 _114_ _058_ 0.013316f
C14364 FILLER_0_13_65/a_36_472# vss 0.007545f
C14365 _370_/a_692_472# net47 0.001021f
C14366 net18 _007_ 0.060872f
C14367 ctln[5] output13/a_224_472# 0.023159f
C14368 _164_ net40 0.048933f
C14369 _413_/a_796_472# net59 0.006163f
C14370 _116_ vdd 0.399137f
C14371 net56 state\[1\] 0.007364f
C14372 _444_/a_36_151# net42 0.006866f
C14373 output34/a_224_472# _046_ 0.006059f
C14374 net63 FILLER_0_18_177/a_1380_472# 0.070445f
C14375 trim_mask\[2\] FILLER_0_2_93/a_484_472# 0.001424f
C14376 net52 _440_/a_2248_156# 0.028463f
C14377 net60 _421_/a_1288_156# 0.001147f
C14378 net10 output10/a_224_472# 0.012455f
C14379 net82 _032_ 0.014269f
C14380 net72 net74 0.035298f
C14381 net81 fanout58/a_36_160# 0.005575f
C14382 _095_ FILLER_0_13_72/a_572_375# 0.003559f
C14383 FILLER_0_6_79/a_124_375# _164_ 0.061565f
C14384 _100_ _283_/a_36_472# 0.033597f
C14385 _408_/a_718_524# vdd 0.002635f
C14386 _024_ net23 0.001994f
C14387 net71 vss 0.335256f
C14388 net49 _440_/a_2248_156# 0.025137f
C14389 net82 trim_val\[4\] 0.511271f
C14390 FILLER_0_7_59/a_124_375# trim_val\[0\] 0.002169f
C14391 net29 net36 0.370099f
C14392 trim_mask\[2\] trim_val\[2\] 0.21814f
C14393 ctln[1] FILLER_0_3_221/a_124_375# 0.001391f
C14394 net63 FILLER_0_17_218/a_124_375# 0.040329f
C14395 _431_/a_36_151# FILLER_0_18_139/a_36_472# 0.002529f
C14396 _078_ FILLER_0_4_213/a_484_472# 0.003702f
C14397 trim_val\[4\] fanout57/a_36_113# 0.078297f
C14398 _447_/a_2248_156# vdd 0.009094f
C14399 _303_/a_36_472# _110_ 0.001606f
C14400 FILLER_0_16_89/a_484_472# net36 0.003595f
C14401 ctln[2] net18 0.106494f
C14402 net57 FILLER_0_8_156/a_484_472# 0.008895f
C14403 _093_ vdd 1.439861f
C14404 _091_ FILLER_0_19_171/a_572_375# 0.013568f
C14405 FILLER_0_16_57/a_36_472# cal_count\[1\] 0.002116f
C14406 _067_ _120_ 0.031156f
C14407 _118_ vdd 0.292155f
C14408 _038_ _067_ 0.503045f
C14409 _141_ FILLER_0_17_142/a_484_472# 0.004527f
C14410 FILLER_0_12_2/a_484_472# _039_ 0.003082f
C14411 net80 _146_ 0.021227f
C14412 ctln[3] FILLER_0_0_232/a_124_375# 0.012394f
C14413 net23 FILLER_0_22_128/a_2812_375# 0.050811f
C14414 _021_ _432_/a_448_472# 0.032563f
C14415 _137_ FILLER_0_16_154/a_932_472# 0.004753f
C14416 net78 _420_/a_448_472# 0.001091f
C14417 net54 _433_/a_2665_112# 0.047439f
C14418 _093_ FILLER_0_18_107/a_572_375# 0.008393f
C14419 FILLER_0_5_72/a_484_472# _440_/a_36_151# 0.001723f
C14420 _077_ FILLER_0_9_72/a_572_375# 0.008103f
C14421 FILLER_0_18_107/a_124_375# mask\[9\] 0.006029f
C14422 FILLER_0_17_64/a_124_375# FILLER_0_17_56/a_572_375# 0.012001f
C14423 _274_/a_1612_497# net4 0.00807f
C14424 net61 net62 0.874859f
C14425 _114_ _389_/a_36_148# 0.009465f
C14426 _187_ _120_ 0.144679f
C14427 _036_ net69 0.353233f
C14428 _008_ _419_/a_796_472# 0.013039f
C14429 FILLER_0_15_142/a_484_472# net36 0.012033f
C14430 ctln[1] FILLER_0_0_266/a_124_375# 0.01186f
C14431 _365_/a_692_472# _156_ 0.001127f
C14432 net74 _370_/a_692_472# 0.005066f
C14433 net63 result[8] 0.013631f
C14434 FILLER_0_17_218/a_124_375# _069_ 0.003162f
C14435 _077_ _453_/a_796_472# 0.003409f
C14436 _440_/a_36_151# _160_ 0.002966f
C14437 _109_ vdd 0.059259f
C14438 result[9] _419_/a_1000_472# 0.012469f
C14439 output46/a_224_472# FILLER_0_20_2/a_124_375# 0.030009f
C14440 net52 _376_/a_36_160# 0.00267f
C14441 _256_/a_2552_68# _076_ 0.00144f
C14442 _449_/a_36_151# FILLER_0_13_72/a_36_472# 0.001723f
C14443 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_572_375# 0.001597f
C14444 net53 FILLER_0_17_142/a_572_375# 0.023771f
C14445 _180_ FILLER_0_15_59/a_36_472# 0.087308f
C14446 FILLER_0_5_128/a_36_472# _163_ 0.009857f
C14447 FILLER_0_8_37/a_484_472# _160_ 0.001767f
C14448 _432_/a_2560_156# _136_ 0.001178f
C14449 net65 FILLER_0_2_177/a_484_472# 0.01675f
C14450 _079_ _265_/a_244_68# 0.021777f
C14451 _029_ FILLER_0_5_88/a_36_472# 0.007596f
C14452 _103_ _418_/a_448_472# 0.002678f
C14453 _449_/a_1000_472# net55 0.001617f
C14454 ctlp[1] FILLER_0_23_290/a_36_472# 0.038596f
C14455 _422_/a_796_472# _109_ 0.002086f
C14456 _116_ _373_/a_244_68# 0.001213f
C14457 _053_ _003_ 0.021223f
C14458 FILLER_0_21_142/a_572_375# _433_/a_2248_156# 0.006739f
C14459 _123_ vdd 0.214703f
C14460 _113_ _279_/a_652_68# 0.001425f
C14461 _142_ _132_ 0.006253f
C14462 ctln[1] ctln[2] 0.047127f
C14463 FILLER_0_7_146/a_124_375# net37 0.005315f
C14464 net54 vdd 0.877573f
C14465 FILLER_0_15_150/a_36_472# net36 0.012318f
C14466 _000_ _411_/a_1000_472# 0.023042f
C14467 _444_/a_2248_156# vdd 0.041347f
C14468 _073_ vdd 0.258125f
C14469 _430_/a_2248_156# _091_ 0.053571f
C14470 FILLER_0_0_232/a_36_472# vss 0.007185f
C14471 FILLER_0_21_142/a_484_472# _140_ 0.011035f
C14472 _330_/a_224_472# vdd 0.001701f
C14473 _176_ _389_/a_36_148# 0.060256f
C14474 net78 _419_/a_1308_423# 0.018598f
C14475 output13/a_224_472# net59 0.007733f
C14476 _046_ _099_ 0.005245f
C14477 net64 mask\[1\] 0.038611f
C14478 _166_ _034_ 0.001936f
C14479 FILLER_0_4_144/a_36_472# net23 0.016933f
C14480 _440_/a_2560_156# _164_ 0.003934f
C14481 ctlp[2] _300_/a_224_472# 0.002954f
C14482 FILLER_0_4_144/a_484_472# trim_mask\[4\] 0.015778f
C14483 _375_/a_36_68# _161_ 0.028567f
C14484 net20 FILLER_0_15_228/a_124_375# 0.047331f
C14485 net65 FILLER_0_1_212/a_124_375# 0.005253f
C14486 net27 output28/a_224_472# 0.011692f
C14487 FILLER_0_20_2/a_572_375# net43 0.051705f
C14488 _010_ _420_/a_2560_156# 0.070902f
C14489 _431_/a_448_472# vss 0.005583f
C14490 _337_/a_49_472# vdd 0.028131f
C14491 FILLER_0_4_144/a_484_472# net47 0.008338f
C14492 FILLER_0_5_212/a_36_472# net22 0.0015f
C14493 _119_ _070_ 1.949038f
C14494 _115_ _114_ 0.148291f
C14495 trimb[1] FILLER_0_18_2/a_124_375# 0.01352f
C14496 FILLER_0_9_28/a_1468_375# net68 0.013121f
C14497 _130_ FILLER_0_11_124/a_36_472# 0.003572f
C14498 _273_/a_36_68# vss 0.095582f
C14499 mask\[8\] _437_/a_2248_156# 0.004415f
C14500 _012_ FILLER_0_23_60/a_124_375# 0.002827f
C14501 _238_/a_67_603# trim_val\[3\] 0.024283f
C14502 FILLER_0_21_28/a_1020_375# vdd 0.04353f
C14503 _131_ _160_ 0.003984f
C14504 net15 vdd 2.073988f
C14505 _053_ net37 0.080949f
C14506 FILLER_0_11_78/a_36_472# vdd -0.001328f
C14507 FILLER_0_11_78/a_572_375# vss 0.004808f
C14508 ctlp[2] _420_/a_2248_156# 0.001156f
C14509 net42 _054_ 0.006314f
C14510 net55 FILLER_0_21_28/a_2724_472# 0.049771f
C14511 _144_ FILLER_0_22_128/a_3260_375# 0.006444f
C14512 FILLER_0_15_290/a_124_375# FILLER_0_15_282/a_572_375# 0.012001f
C14513 _265_/a_244_68# cal_itt\[1\] 0.024108f
C14514 _064_ vss 0.228443f
C14515 mask\[4\] _098_ 0.041526f
C14516 net82 FILLER_0_4_213/a_572_375# 0.00123f
C14517 cal_itt\[2\] _260_/a_36_68# 0.004081f
C14518 net67 FILLER_0_9_60/a_572_375# 0.011073f
C14519 _144_ net33 0.042826f
C14520 _326_/a_36_160# _070_ 0.018037f
C14521 FILLER_0_19_55/a_36_472# FILLER_0_18_53/a_124_375# 0.001684f
C14522 _253_/a_1100_68# _084_ 0.001651f
C14523 _228_/a_36_68# net22 0.052558f
C14524 _116_ _279_/a_244_68# 0.001752f
C14525 _055_ _090_ 0.040233f
C14526 ctln[8] _168_ 0.001145f
C14527 FILLER_0_5_128/a_484_472# vss 0.004051f
C14528 output43/a_224_472# trimb[3] 0.070044f
C14529 FILLER_0_3_142/a_36_472# _370_/a_848_380# 0.001207f
C14530 FILLER_0_4_107/a_572_375# net47 0.006041f
C14531 net15 _441_/a_1204_472# 0.005939f
C14532 output48/a_224_472# net59 0.039277f
C14533 net81 _429_/a_36_151# 0.018551f
C14534 FILLER_0_5_164/a_124_375# net37 0.008158f
C14535 _140_ _023_ 0.079452f
C14536 FILLER_0_6_90/a_572_375# vdd 0.028324f
C14537 net42 vss 0.017902f
C14538 _413_/a_2665_112# net59 0.066623f
C14539 _418_/a_1000_472# vss 0.001193f
C14540 net81 net18 0.102876f
C14541 _120_ net23 0.147166f
C14542 FILLER_0_18_2/a_3260_375# FILLER_0_20_31/a_36_472# 0.001338f
C14543 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_36_472# 0.086635f
C14544 cal_itt\[2\] net4 0.333682f
C14545 _333_/a_36_160# _097_ 0.001332f
C14546 _115_ _176_ 1.300336f
C14547 _171_ FILLER_0_10_94/a_484_472# 0.001446f
C14548 FILLER_0_22_177/a_1380_472# net33 0.016037f
C14549 _073_ net9 0.005417f
C14550 result[8] _435_/a_2665_112# 0.001855f
C14551 _122_ FILLER_0_5_181/a_124_375# 0.001352f
C14552 net52 FILLER_0_9_72/a_1468_375# 0.003576f
C14553 _100_ FILLER_0_12_236/a_572_375# 0.015109f
C14554 FILLER_0_13_142/a_1020_375# net23 0.047331f
C14555 _445_/a_2248_156# net17 0.06175f
C14556 FILLER_0_5_128/a_572_375# vdd 0.008326f
C14557 net39 vdd 0.2282f
C14558 _130_ _428_/a_2665_112# 0.001241f
C14559 FILLER_0_1_266/a_484_472# vdd 0.003622f
C14560 _042_ vss 0.008272f
C14561 net51 vdd 0.692054f
C14562 _069_ _060_ 0.538161f
C14563 _126_ _090_ 0.003538f
C14564 _425_/a_36_151# net37 0.003145f
C14565 _040_ FILLER_0_16_115/a_36_472# 0.001876f
C14566 _077_ _319_/a_672_472# 0.001602f
C14567 _077_ FILLER_0_9_60/a_36_472# 0.038809f
C14568 FILLER_0_8_107/a_36_472# FILLER_0_7_104/a_484_472# 0.026657f
C14569 _095_ _113_ 0.004037f
C14570 FILLER_0_17_142/a_124_375# FILLER_0_17_133/a_124_375# 0.003228f
C14571 FILLER_0_11_109/a_124_375# _120_ 0.016902f
C14572 _378_/a_224_472# _165_ 0.00481f
C14573 net75 _426_/a_448_472# 0.041705f
C14574 _402_/a_2172_497# _180_ 0.001094f
C14575 _328_/a_36_113# net70 0.00292f
C14576 _137_ FILLER_0_19_155/a_124_375# 0.00129f
C14577 _428_/a_2560_156# _131_ 0.002853f
C14578 _442_/a_36_151# FILLER_0_2_127/a_124_375# 0.001597f
C14579 FILLER_0_5_88/a_36_472# _163_ 0.006541f
C14580 _413_/a_1000_472# vdd 0.002781f
C14581 mask\[2\] net21 0.033368f
C14582 _106_ _201_/a_67_603# 0.00327f
C14583 _115_ _124_ 0.045023f
C14584 net38 _221_/a_36_160# 0.029767f
C14585 net82 FILLER_0_3_221/a_1020_375# 0.010208f
C14586 _333_/a_36_160# mask\[2\] 0.022517f
C14587 _350_/a_49_472# vdd 0.026837f
C14588 vss FILLER_0_4_91/a_484_472# 0.003328f
C14589 FILLER_0_21_133/a_124_375# _140_ 0.018383f
C14590 FILLER_0_8_247/a_572_375# calibrate 0.008498f
C14591 FILLER_0_15_142/a_572_375# net23 0.006327f
C14592 FILLER_0_16_89/a_124_375# vdd 0.01011f
C14593 ctlp[1] FILLER_0_24_274/a_932_472# 0.003603f
C14594 mask\[9\] _423_/a_2665_112# 0.001735f
C14595 _027_ net71 0.057875f
C14596 FILLER_0_3_172/a_2276_472# net22 0.012151f
C14597 FILLER_0_5_212/a_36_472# vdd 0.107657f
C14598 FILLER_0_5_212/a_124_375# vss 0.006344f
C14599 output48/a_224_472# net64 0.002845f
C14600 net31 _094_ 0.203395f
C14601 FILLER_0_4_185/a_124_375# vss 0.024832f
C14602 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_124_375# 0.012001f
C14603 _422_/a_2665_112# mask\[7\] 0.028271f
C14604 FILLER_0_18_2/a_1020_375# net44 0.009108f
C14605 net16 ctln[9] 0.07797f
C14606 FILLER_0_17_56/a_36_472# _404_/a_36_472# 0.004546f
C14607 mask\[8\] net25 0.035648f
C14608 net23 mask\[6\] 0.025699f
C14609 FILLER_0_21_142/a_484_472# FILLER_0_21_150/a_36_472# 0.013277f
C14610 ctlp[1] net33 0.11288f
C14611 FILLER_0_10_214/a_36_472# _070_ 0.014734f
C14612 net63 _093_ 0.109689f
C14613 net18 net30 0.09055f
C14614 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_124_375# 0.005439f
C14615 _308_/a_848_380# FILLER_0_9_105/a_124_375# 0.005599f
C14616 net19 _418_/a_2665_112# 0.040822f
C14617 _427_/a_1308_423# _095_ 0.022677f
C14618 net27 _426_/a_796_472# 0.001678f
C14619 _069_ _116_ 0.390834f
C14620 _150_ mask\[9\] 0.162185f
C14621 _053_ FILLER_0_6_47/a_932_472# 0.011457f
C14622 net62 FILLER_0_15_290/a_124_375# 0.034614f
C14623 mask\[0\] net64 0.45093f
C14624 fanout75/a_36_113# _317_/a_36_113# 0.001442f
C14625 net20 result[5] 0.045364f
C14626 _346_/a_257_69# _144_ 0.001089f
C14627 _430_/a_448_472# vss 0.003371f
C14628 _028_ FILLER_0_7_72/a_2276_472# 0.001777f
C14629 FILLER_0_13_65/a_36_472# _095_ 0.003171f
C14630 _008_ net77 0.029049f
C14631 _065_ net17 0.035195f
C14632 fanout52/a_36_160# net23 0.009496f
C14633 _228_/a_36_68# vdd 0.036391f
C14634 FILLER_0_4_123/a_124_375# _160_ 0.038272f
C14635 _066_ _386_/a_692_472# 0.001958f
C14636 net38 FILLER_0_20_15/a_36_472# 0.070475f
C14637 _086_ _057_ 0.82902f
C14638 net35 _012_ 0.007543f
C14639 _428_/a_1308_423# _017_ 0.005962f
C14640 _428_/a_448_472# net53 0.001959f
C14641 net68 trim_mask\[1\] 0.054055f
C14642 _162_ _374_/a_36_68# 0.005729f
C14643 _369_/a_36_68# vss 0.002343f
C14644 output34/a_224_472# _103_ 0.027876f
C14645 _044_ vss 0.038421f
C14646 _122_ _242_/a_36_160# 0.005377f
C14647 FILLER_0_20_169/a_36_472# _140_ 0.023696f
C14648 state\[2\] net23 0.331644f
C14649 _431_/a_2665_112# vss 0.033886f
C14650 FILLER_0_7_104/a_484_472# FILLER_0_9_105/a_572_375# 0.001188f
C14651 FILLER_0_11_142/a_484_472# vss 0.033416f
C14652 net45 vss 0.028798f
C14653 net58 FILLER_0_9_282/a_124_375# 0.021949f
C14654 _086_ _250_/a_36_68# 0.001132f
C14655 FILLER_0_18_107/a_3260_375# vss 0.056926f
C14656 FILLER_0_18_107/a_36_472# vdd 0.116746f
C14657 _139_ _137_ 0.093639f
C14658 _093_ _069_ 0.008325f
C14659 _069_ _118_ 0.010986f
C14660 _434_/a_796_472# mask\[6\] 0.004416f
C14661 _004_ net79 0.27387f
C14662 net20 output20/a_224_472# 0.024692f
C14663 FILLER_0_7_104/a_36_472# vdd 0.096343f
C14664 FILLER_0_7_104/a_1468_375# vss 0.003442f
C14665 _242_/a_36_160# _169_ 0.051038f
C14666 trim_mask\[1\] _156_ 0.007519f
C14667 _114_ _134_ 0.015298f
C14668 fanout50/a_36_160# _168_ 0.033707f
C14669 net52 _384_/a_224_472# 0.001238f
C14670 mask\[4\] FILLER_0_18_177/a_3260_375# 0.013881f
C14671 net47 _167_ 0.003019f
C14672 net44 _245_/a_672_472# 0.001285f
C14673 net55 FILLER_0_21_60/a_36_472# 0.06794f
C14674 ctln[2] net65 0.113266f
C14675 _077_ FILLER_0_7_72/a_3172_472# 0.001923f
C14676 _238_/a_67_603# _065_ 0.005075f
C14677 _189_/a_67_603# vdd 0.01494f
C14678 net52 _441_/a_448_472# 0.04874f
C14679 FILLER_0_4_107/a_572_375# _154_ 0.052251f
C14680 FILLER_0_17_72/a_932_472# FILLER_0_18_76/a_484_472# 0.05841f
C14681 _088_ FILLER_0_3_212/a_124_375# 0.0042f
C14682 mask\[3\] FILLER_0_18_177/a_2364_375# 0.002935f
C14683 output40/a_224_472# net40 0.0374f
C14684 FILLER_0_12_236/a_572_375# _060_ 0.001597f
C14685 net64 _099_ 0.007017f
C14686 _076_ _160_ 0.006506f
C14687 _161_ _070_ 0.027757f
C14688 FILLER_0_1_212/a_36_472# net59 0.002567f
C14689 FILLER_0_24_96/a_36_472# net25 0.040228f
C14690 net2 vdd 0.434557f
C14691 net18 _417_/a_36_151# 0.020548f
C14692 _417_/a_448_472# net30 0.042386f
C14693 _062_ _226_/a_1044_68# 0.001944f
C14694 _072_ _375_/a_1388_497# 0.001138f
C14695 _441_/a_448_472# net49 0.001245f
C14696 mask\[9\] _026_ 0.002924f
C14697 _096_ _098_ 0.00638f
C14698 _157_ _156_ 0.005264f
C14699 _028_ vdd 0.626868f
C14700 net15 _423_/a_2560_156# 0.007083f
C14701 _093_ FILLER_0_18_139/a_36_472# 0.008761f
C14702 _097_ mask\[1\] 0.001232f
C14703 output9/a_224_472# net4 0.042449f
C14704 net50 FILLER_0_9_60/a_36_472# 0.001914f
C14705 _428_/a_36_151# FILLER_0_14_107/a_572_375# 0.001597f
C14706 FILLER_0_12_136/a_572_375# _120_ 0.001584f
C14707 _449_/a_2560_156# _038_ 0.010532f
C14708 ctlp[6] _050_ 0.100418f
C14709 net61 _422_/a_36_151# 0.003736f
C14710 net63 _337_/a_49_472# 0.001801f
C14711 FILLER_0_3_172/a_2276_472# vdd 0.00806f
C14712 _131_ _133_ 0.20118f
C14713 _129_ _070_ 0.056776f
C14714 result[7] _420_/a_2665_112# 0.039448f
C14715 trim_mask\[4\] net22 0.027368f
C14716 mask\[5\] _009_ 0.001095f
C14717 net67 trim_mask\[1\] 0.01761f
C14718 _076_ _223_/a_36_160# 0.001756f
C14719 net80 mask\[2\] 0.048734f
C14720 FILLER_0_19_171/a_484_472# _434_/a_36_151# 0.002841f
C14721 _144_ net35 0.036236f
C14722 fanout71/a_36_113# _149_ 0.001315f
C14723 state\[1\] _090_ 0.087906f
C14724 trimb[1] _452_/a_3129_107# 0.007229f
C14725 FILLER_0_18_2/a_1468_375# net38 0.016983f
C14726 _012_ FILLER_0_23_44/a_124_375# 0.002474f
C14727 net4 _246_/a_36_68# 0.003771f
C14728 _176_ _134_ 0.035146f
C14729 _114_ _267_/a_672_472# 0.001566f
C14730 FILLER_0_4_213/a_124_375# net59 0.039014f
C14731 output32/a_224_472# _094_ 0.005545f
C14732 net34 _024_ 0.009705f
C14733 _044_ _416_/a_2248_156# 0.005198f
C14734 FILLER_0_21_142/a_36_472# _098_ 0.002964f
C14735 net44 net6 0.005889f
C14736 vdd clkc 0.190259f
C14737 FILLER_0_9_28/a_1916_375# net51 0.001008f
C14738 FILLER_0_15_212/a_36_472# net22 0.003143f
C14739 net57 _120_ 0.012391f
C14740 net20 _199_/a_36_160# 0.05178f
C14741 _408_/a_728_93# _402_/a_56_567# 0.001359f
C14742 net52 cal_count\[3\] 0.348542f
C14743 net61 fanout77/a_36_113# 0.080943f
C14744 net35 FILLER_0_22_177/a_1380_472# 0.01447f
C14745 _045_ vdd 0.246567f
C14746 _277_/a_36_160# _094_ 0.007538f
C14747 mask\[2\] mask\[1\] 0.059794f
C14748 ctlp[1] FILLER_0_23_282/a_572_375# 0.009848f
C14749 FILLER_0_5_172/a_124_375# net22 0.002388f
C14750 _086_ _310_/a_49_472# 0.013039f
C14751 FILLER_0_4_197/a_124_375# net59 0.001026f
C14752 result[9] _421_/a_1308_423# 0.011854f
C14753 FILLER_0_14_181/a_36_472# vdd 0.027265f
C14754 FILLER_0_14_181/a_124_375# vss 0.009291f
C14755 net57 FILLER_0_13_142/a_1020_375# 0.009442f
C14756 output10/a_224_472# net8 0.010088f
C14757 net34 FILLER_0_22_128/a_2812_375# 0.005158f
C14758 _103_ _099_ 0.025799f
C14759 FILLER_0_15_205/a_124_375# net21 0.002912f
C14760 ctln[4] net21 0.009947f
C14761 fanout82/a_36_113# net82 0.003741f
C14762 FILLER_0_1_212/a_124_375# net11 0.029766f
C14763 valid vdd 0.148392f
C14764 _140_ FILLER_0_22_128/a_2724_472# 0.004196f
C14765 _322_/a_848_380# FILLER_0_9_142/a_124_375# 0.001721f
C14766 _124_ _134_ 0.002508f
C14767 net23 _433_/a_2248_156# 0.005588f
C14768 _430_/a_2248_156# FILLER_0_15_212/a_932_472# 0.035805f
C14769 net2 net9 0.001033f
C14770 FILLER_0_18_171/a_124_375# _143_ 0.005331f
C14771 _383_/a_36_472# vss 0.002794f
C14772 _132_ _017_ 0.155924f
C14773 net38 cal_count\[2\] 0.047195f
C14774 FILLER_0_8_247/a_1468_375# vss 0.054783f
C14775 FILLER_0_8_247/a_36_472# vdd 0.112197f
C14776 trim_val\[3\] FILLER_0_2_93/a_36_472# 0.015653f
C14777 net17 _034_ 0.020793f
C14778 _055_ _117_ 0.242156f
C14779 net55 FILLER_0_18_37/a_1020_375# 0.005661f
C14780 output44/a_224_472# FILLER_0_18_2/a_1916_375# 0.032639f
C14781 _136_ _335_/a_49_472# 0.039074f
C14782 trim_val\[1\] _034_ 0.001535f
C14783 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_124_375# 0.012001f
C14784 _322_/a_124_24# _128_ 0.02077f
C14785 _168_ _164_ 0.092012f
C14786 FILLER_0_10_78/a_572_375# FILLER_0_11_78/a_572_375# 0.05841f
C14787 net78 _421_/a_36_151# 0.001368f
C14788 _412_/a_796_472# net58 0.001182f
C14789 FILLER_0_16_255/a_124_375# _094_ 0.004398f
C14790 _081_ _160_ 0.00816f
C14791 _105_ net34 0.784678f
C14792 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_484_472# 0.013276f
C14793 _104_ _420_/a_2560_156# 0.002734f
C14794 _064_ _036_ 0.003286f
C14795 trim_mask\[2\] trim_val\[3\] 0.003342f
C14796 output32/a_224_472# net78 0.002901f
C14797 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_572_375# 0.086635f
C14798 ctln[1] _411_/a_1000_472# 0.040782f
C14799 net16 _379_/a_36_472# 0.01109f
C14800 _414_/a_2560_156# _074_ 0.001344f
C14801 net38 _450_/a_448_472# 0.031891f
C14802 _011_ _422_/a_448_472# 0.044695f
C14803 _000_ net59 0.004356f
C14804 FILLER_0_7_72/a_3172_472# net50 0.001428f
C14805 _086_ _395_/a_1044_488# 0.001091f
C14806 FILLER_0_12_136/a_572_375# state\[2\] 0.001955f
C14807 FILLER_0_16_241/a_36_472# net36 0.001988f
C14808 FILLER_0_12_136/a_1468_375# net53 0.002709f
C14809 _394_/a_728_93# FILLER_0_13_72/a_484_472# 0.018997f
C14810 net81 net65 0.083316f
C14811 output26/a_224_472# FILLER_0_23_44/a_932_472# 0.0323f
C14812 trim_mask\[4\] vdd 0.20602f
C14813 _098_ FILLER_0_15_180/a_484_472# 0.014511f
C14814 _444_/a_2665_112# net67 0.03521f
C14815 net47 vdd 2.422992f
C14816 FILLER_0_9_223/a_124_375# state\[0\] 0.002912f
C14817 _015_ net4 0.003985f
C14818 net52 _443_/a_2665_112# 0.05031f
C14819 _074_ _374_/a_36_68# 0.001447f
C14820 net57 fanout52/a_36_160# 0.122432f
C14821 _327_/a_36_472# _130_ 0.001474f
C14822 output14/a_224_472# _442_/a_448_472# 0.008149f
C14823 _315_/a_244_497# _120_ 0.006419f
C14824 FILLER_0_16_57/a_1468_375# vdd 0.020146f
C14825 FILLER_0_16_57/a_1020_375# vss 0.004487f
C14826 net35 _436_/a_1204_472# 0.005186f
C14827 _255_/a_224_552# FILLER_0_6_177/a_572_375# 0.001776f
C14828 FILLER_0_21_133/a_36_472# net54 0.02286f
C14829 _174_ _179_ 0.003183f
C14830 _413_/a_2560_156# net65 0.011101f
C14831 _415_/a_796_472# vdd 0.001842f
C14832 net15 _449_/a_36_151# 0.020788f
C14833 _012_ vdd 0.261844f
C14834 _374_/a_36_68# _076_ 0.026674f
C14835 _056_ _070_ 0.045548f
C14836 FILLER_0_15_212/a_572_375# mask\[1\] 0.012463f
C14837 FILLER_0_15_212/a_1468_375# vss 0.060206f
C14838 FILLER_0_15_212/a_36_472# vdd 0.105575f
C14839 net57 state\[2\] 1.25275f
C14840 FILLER_0_16_89/a_484_472# _176_ 0.004026f
C14841 trim_mask\[2\] _367_/a_36_68# 0.001302f
C14842 fanout71/a_36_113# FILLER_0_20_107/a_124_375# 0.002853f
C14843 trimb[1] vss 0.048527f
C14844 FILLER_0_16_154/a_1380_472# vss 0.003609f
C14845 FILLER_0_5_172/a_124_375# vdd 0.028449f
C14846 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_36_472# 0.009654f
C14847 _445_/a_2665_112# _444_/a_448_472# 0.001178f
C14848 net34 output19/a_224_472# 0.122464f
C14849 _065_ _447_/a_1308_423# 0.024822f
C14850 net57 _386_/a_692_472# 0.00409f
C14851 _011_ _108_ 0.036521f
C14852 FILLER_0_20_169/a_124_375# _098_ 0.019219f
C14853 net79 FILLER_0_15_282/a_124_375# 0.001058f
C14854 sample fanout59/a_36_160# 0.001854f
C14855 trim_mask\[1\] FILLER_0_6_47/a_1916_375# 0.007169f
C14856 FILLER_0_9_223/a_36_472# vdd 0.030289f
C14857 FILLER_0_19_111/a_484_472# vss 0.003811f
C14858 trimb[1] FILLER_0_20_15/a_932_472# 0.001069f
C14859 net62 FILLER_0_15_282/a_572_375# 0.007699f
C14860 _434_/a_1308_423# vdd 0.033494f
C14861 _067_ _450_/a_448_472# 0.003113f
C14862 _148_ _352_/a_257_69# 0.001417f
C14863 _181_ _182_ 0.02735f
C14864 net38 _043_ 0.117134f
C14865 _052_ FILLER_0_18_53/a_124_375# 0.001585f
C14866 FILLER_0_15_142/a_124_375# vdd -0.003809f
C14867 ctln[3] net10 0.873575f
C14868 _411_/a_1204_472# net75 0.008304f
C14869 FILLER_0_8_107/a_124_375# _133_ 0.048874f
C14870 mask\[5\] FILLER_0_20_193/a_36_472# 0.013533f
C14871 _144_ _433_/a_2665_112# 0.030413f
C14872 _430_/a_36_151# vss 0.011779f
C14873 net36 cal_count\[1\] 0.011481f
C14874 FILLER_0_15_59/a_484_472# vdd 0.010447f
C14875 FILLER_0_15_59/a_36_472# vss 0.00459f
C14876 ctlp[8] mask\[8\] 0.001554f
C14877 FILLER_0_4_185/a_36_472# net22 0.006506f
C14878 _254_/a_244_472# _074_ 0.002716f
C14879 _077_ _062_ 0.037598f
C14880 _098_ _201_/a_67_603# 0.005932f
C14881 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_124_375# 0.005439f
C14882 FILLER_0_12_124/a_124_375# _114_ 0.006974f
C14883 _119_ calibrate 0.062309f
C14884 FILLER_0_11_101/a_572_375# _070_ 0.011557f
C14885 _069_ _228_/a_36_68# 0.001676f
C14886 FILLER_0_15_150/a_124_375# net53 0.041074f
C14887 output8/a_224_472# FILLER_0_3_221/a_1020_375# 0.03228f
C14888 _133_ _076_ 0.11688f
C14889 _070_ _068_ 1.019801f
C14890 net35 FILLER_0_22_128/a_572_375# 0.010439f
C14891 trim_val\[4\] FILLER_0_3_172/a_484_472# 0.002633f
C14892 net74 vdd 1.451847f
C14893 FILLER_0_7_146/a_36_472# _068_ 0.012745f
C14894 _104_ net32 0.342568f
C14895 _376_/a_36_160# FILLER_0_6_79/a_124_375# 0.004736f
C14896 output13/a_224_472# trim_val\[4\] 0.001014f
C14897 _258_/a_36_160# net20 0.041584f
C14898 _074_ _317_/a_36_113# 0.003383f
C14899 _064_ _445_/a_796_472# 0.00673f
C14900 FILLER_0_13_212/a_1380_472# net79 0.006824f
C14901 FILLER_0_5_117/a_36_472# _160_ 0.005314f
C14902 FILLER_0_4_107/a_484_472# FILLER_0_2_111/a_124_375# 0.001404f
C14903 FILLER_0_7_72/a_1916_375# FILLER_0_5_88/a_36_472# 0.0027f
C14904 output42/a_224_472# _221_/a_36_160# 0.017421f
C14905 net32 vss 0.824307f
C14906 _126_ FILLER_0_11_142/a_36_472# 0.001428f
C14907 _253_/a_36_68# vdd 0.016219f
C14908 net61 _419_/a_36_151# 0.019141f
C14909 mask\[5\] FILLER_0_18_177/a_1916_375# 0.002014f
C14910 net80 FILLER_0_22_177/a_36_472# 0.018848f
C14911 net69 fanout49/a_36_160# 0.005942f
C14912 FILLER_0_5_109/a_36_472# FILLER_0_4_107/a_124_375# 0.001684f
C14913 _144_ vdd 0.40911f
C14914 _431_/a_1000_472# _137_ 0.010168f
C14915 fanout58/a_36_160# net59 0.048057f
C14916 mask\[1\] FILLER_0_15_205/a_124_375# 0.007883f
C14917 FILLER_0_9_28/a_572_375# net40 0.001406f
C14918 trimb[0] trimb[3] 0.549457f
C14919 _067_ _043_ 0.189767f
C14920 _411_/a_1308_423# net8 0.0176f
C14921 fanout78/a_36_113# net18 0.001419f
C14922 _372_/a_170_472# vss 0.027819f
C14923 _232_/a_67_603# trim_val\[1\] 0.009588f
C14924 _414_/a_2560_156# _081_ 0.008322f
C14925 FILLER_0_8_127/a_36_472# _058_ 0.003283f
C14926 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_484_472# 0.026657f
C14927 fanout75/a_36_113# net59 0.00817f
C14928 FILLER_0_12_220/a_484_472# vss 0.006724f
C14929 FILLER_0_12_220/a_932_472# vdd 0.003359f
C14930 trim_mask\[4\] FILLER_0_2_165/a_124_375# 0.011181f
C14931 FILLER_0_16_107/a_36_472# net14 0.004691f
C14932 FILLER_0_18_2/a_1828_472# net55 0.011802f
C14933 _058_ FILLER_0_8_156/a_572_375# 0.007692f
C14934 FILLER_0_17_133/a_36_472# FILLER_0_19_134/a_124_375# 0.001188f
C14935 _079_ net22 0.039221f
C14936 _173_ vdd 0.080629f
C14937 FILLER_0_17_72/a_1020_375# _451_/a_3129_107# 0.001202f
C14938 _187_ _043_ 0.011995f
C14939 net39 _445_/a_1308_423# 0.008252f
C14940 trim[1] _445_/a_36_151# 0.008362f
C14941 FILLER_0_20_193/a_484_472# FILLER_0_19_195/a_124_375# 0.001543f
C14942 _431_/a_2560_156# net36 0.001858f
C14943 FILLER_0_5_72/a_484_472# _029_ 0.004625f
C14944 FILLER_0_5_72/a_1020_375# trim_mask\[1\] 0.010728f
C14945 FILLER_0_22_177/a_932_472# vss -0.001894f
C14946 FILLER_0_22_177/a_1380_472# vdd 0.007188f
C14947 _099_ mask\[2\] 0.776725f
C14948 net68 net66 0.81104f
C14949 _093_ _424_/a_2665_112# 0.001854f
C14950 _159_ vdd 0.025131f
C14951 _020_ _431_/a_1308_423# 0.001997f
C14952 _426_/a_2560_156# net64 0.00801f
C14953 output34/a_224_472# _419_/a_2665_112# 0.010731f
C14954 FILLER_0_18_2/a_2364_375# _452_/a_1353_112# 0.001068f
C14955 net34 mask\[6\] 0.231853f
C14956 mask\[2\] FILLER_0_16_154/a_36_472# 0.312123f
C14957 _452_/a_448_472# net40 0.047031f
C14958 FILLER_0_4_107/a_932_472# _160_ 0.014254f
C14959 FILLER_0_4_213/a_484_472# vss 0.007857f
C14960 net52 FILLER_0_0_130/a_124_375# 0.004055f
C14961 _057_ _061_ 0.030546f
C14962 net32 _107_ 0.003155f
C14963 FILLER_0_14_99/a_36_472# FILLER_0_14_107/a_36_472# 0.002296f
C14964 _418_/a_796_472# _007_ 0.012286f
C14965 _057_ _311_/a_66_473# 0.042545f
C14966 FILLER_0_17_72/a_2364_375# _131_ 0.006037f
C14967 FILLER_0_5_109/a_484_472# vss 0.00212f
C14968 output38/a_224_472# output41/a_224_472# 0.00607f
C14969 trim_val\[4\] _241_/a_224_472# 0.003005f
C14970 _294_/a_224_472# mask\[2\] 0.001715f
C14971 net55 FILLER_0_13_72/a_572_375# 0.005919f
C14972 _065_ trim_mask\[2\] 0.002792f
C14973 fanout51/a_36_113# net55 0.010147f
C14974 net38 net67 1.762405f
C14975 FILLER_0_17_72/a_2724_472# net14 0.007133f
C14976 _136_ _451_/a_1697_156# 0.001053f
C14977 _154_ vdd 0.639978f
C14978 _449_/a_2248_156# vss 0.008071f
C14979 _449_/a_2665_112# vdd 0.012848f
C14980 FILLER_0_12_136/a_124_375# vdd 0.004378f
C14981 net26 _423_/a_448_472# 0.011612f
C14982 FILLER_0_20_87/a_124_375# net71 0.003629f
C14983 FILLER_0_18_2/a_1828_472# net17 0.008573f
C14984 net53 FILLER_0_14_123/a_36_472# 0.062713f
C14985 result[6] _421_/a_2248_156# 0.031832f
C14986 _092_ FILLER_0_18_209/a_572_375# 0.00609f
C14987 FILLER_0_4_185/a_36_472# vdd 0.122463f
C14988 net74 _135_ 0.002261f
C14989 FILLER_0_16_57/a_36_472# cal_count\[2\] 0.001952f
C14990 sample net5 0.359975f
C14991 mask\[0\] FILLER_0_15_212/a_572_375# 0.001158f
C14992 _443_/a_1456_156# net23 0.001009f
C14993 fanout75/a_36_113# _122_ 0.001035f
C14994 _131_ _427_/a_36_151# 0.0012f
C14995 FILLER_0_3_142/a_124_375# vdd 0.00167f
C14996 net4 _084_ 0.029194f
C14997 _142_ FILLER_0_17_133/a_124_375# 0.022066f
C14998 _059_ FILLER_0_8_156/a_36_472# 0.18373f
C14999 net54 _140_ 1.37516f
C15000 FILLER_0_18_177/a_1916_375# FILLER_0_19_195/a_36_472# 0.001684f
C15001 _149_ _437_/a_2560_156# 0.008064f
C15002 FILLER_0_17_38/a_36_472# _452_/a_36_151# 0.096503f
C15003 _070_ _152_ 0.114651f
C15004 _133_ _081_ 0.002847f
C15005 FILLER_0_10_78/a_484_472# cal_count\[3\] 0.001112f
C15006 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_124_375# 0.003732f
C15007 _442_/a_448_472# vdd 0.006758f
C15008 _442_/a_36_151# vss 0.021278f
C15009 _123_ FILLER_0_6_231/a_484_472# 0.001396f
C15010 mask\[4\] net21 0.049513f
C15011 mask\[5\] net33 0.251971f
C15012 output36/a_224_472# output31/a_224_472# 0.00289f
C15013 fanout70/a_36_113# _136_ 0.002788f
C15014 _004_ net19 0.112289f
C15015 _307_/a_234_472# _113_ 0.007518f
C15016 net38 _445_/a_448_472# 0.023336f
C15017 net15 FILLER_0_6_47/a_2364_375# 0.022624f
C15018 _176_ FILLER_0_15_72/a_36_472# 0.002101f
C15019 net50 _444_/a_2560_156# 0.001479f
C15020 _178_ _402_/a_2172_497# 0.003871f
C15021 net25 _423_/a_2665_112# 0.007096f
C15022 net41 _446_/a_1000_472# 0.01097f
C15023 net47 _450_/a_1353_112# 0.018879f
C15024 ctlp[1] vdd 0.942436f
C15025 net68 FILLER_0_3_54/a_124_375# 0.022559f
C15026 _126_ _172_ 0.017618f
C15027 _057_ _072_ 0.048392f
C15028 _305_/a_36_159# vss 0.003366f
C15029 _128_ _315_/a_1657_68# 0.0013f
C15030 mask\[4\] FILLER_0_19_171/a_932_472# 0.004669f
C15031 _340_/a_36_160# mask\[6\] 0.010151f
C15032 FILLER_0_19_47/a_572_375# _013_ 0.012993f
C15033 _411_/a_1000_472# net65 0.001916f
C15034 FILLER_0_14_181/a_124_375# _095_ 0.005538f
C15035 FILLER_0_19_155/a_572_375# vss 0.004538f
C15036 net73 vss 0.342554f
C15037 FILLER_0_13_206/a_36_472# vss 0.003985f
C15038 _411_/a_2560_156# net75 0.007047f
C15039 FILLER_0_9_28/a_932_472# vdd 0.04397f
C15040 net23 FILLER_0_16_154/a_124_375# 0.002689f
C15041 fanout82/a_36_113# calibrate 0.004982f
C15042 ctln[2] FILLER_0_1_266/a_572_375# 0.012126f
C15043 _132_ cal_count\[3\] 0.193553f
C15044 net67 _067_ 0.151887f
C15045 _072_ _250_/a_36_68# 0.007337f
C15046 FILLER_0_3_221/a_36_472# vss 0.046345f
C15047 FILLER_0_3_221/a_484_472# vdd 0.002974f
C15048 _401_/a_36_68# FILLER_0_15_59/a_36_472# 0.019798f
C15049 _436_/a_1204_472# vdd 0.003143f
C15050 FILLER_0_11_124/a_124_375# _118_ 0.030768f
C15051 _423_/a_2560_156# _012_ 0.004165f
C15052 net73 FILLER_0_18_107/a_1020_375# 0.04487f
C15053 _077_ _308_/a_848_380# 0.010515f
C15054 _431_/a_36_151# _137_ 0.011412f
C15055 mask\[7\] _208_/a_36_160# 0.105845f
C15056 ctln[8] net50 0.0032f
C15057 _098_ _113_ 0.001472f
C15058 _439_/a_1000_472# vss 0.032923f
C15059 FILLER_0_22_128/a_36_472# _433_/a_36_151# 0.001653f
C15060 net62 _429_/a_2665_112# 0.02887f
C15061 _087_ vss 0.09895f
C15062 _079_ vdd 0.476075f
C15063 ctln[4] _413_/a_2665_112# 0.001394f
C15064 net20 _418_/a_2665_112# 0.013517f
C15065 _053_ trim_mask\[0\] 0.007667f
C15066 net15 _424_/a_2665_112# 0.046592f
C15067 output29/a_224_472# net29 0.038602f
C15068 net63 FILLER_0_15_212/a_36_472# 0.059367f
C15069 _445_/a_448_472# net66 0.010949f
C15070 FILLER_0_8_24/a_484_472# FILLER_0_8_37/a_36_472# 0.001963f
C15071 net19 FILLER_0_23_274/a_124_375# 0.01233f
C15072 net20 _091_ 0.0557f
C15073 net23 _043_ 0.042095f
C15074 net53 _136_ 0.099584f
C15075 _076_ _121_ 0.013717f
C15076 FILLER_0_14_99/a_36_472# vss 0.003598f
C15077 FILLER_0_19_125/a_36_472# net73 0.004017f
C15078 _081_ FILLER_0_5_164/a_36_472# 0.001603f
C15079 net57 _280_/a_224_472# 0.001032f
C15080 FILLER_0_12_136/a_36_472# cal_count\[3\] 0.006102f
C15081 net50 FILLER_0_6_90/a_484_472# 0.012286f
C15082 net44 FILLER_0_12_2/a_572_375# 0.041552f
C15083 _443_/a_36_151# _170_ 0.014771f
C15084 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_1020_375# 0.001597f
C15085 FILLER_0_12_2/a_36_472# vss 0.003757f
C15086 net63 _434_/a_1308_423# 0.003686f
C15087 _177_ vdd 0.111636f
C15088 net53 FILLER_0_13_142/a_124_375# 0.001599f
C15089 mask\[0\] FILLER_0_12_220/a_1468_375# 0.001484f
C15090 _074_ _312_/a_672_472# 0.005399f
C15091 _161_ calibrate 0.044443f
C15092 FILLER_0_9_28/a_2724_472# net68 0.010755f
C15093 FILLER_0_10_37/a_124_375# vss 0.006228f
C15094 FILLER_0_10_37/a_36_472# vdd 0.141896f
C15095 FILLER_0_8_127/a_124_375# vss 0.019066f
C15096 net82 net69 0.005307f
C15097 FILLER_0_24_274/a_124_375# vdd 0.012632f
C15098 FILLER_0_15_142/a_572_375# net36 0.006382f
C15099 net18 net59 0.695067f
C15100 _448_/a_448_472# _037_ 0.044085f
C15101 _120_ FILLER_0_10_107/a_572_375# 0.002214f
C15102 _141_ mask\[6\] 0.009844f
C15103 _086_ vss 0.615299f
C15104 net28 _045_ 0.05144f
C15105 net7 net16 0.033509f
C15106 output32/a_224_472# _418_/a_2248_156# 0.024448f
C15107 output7/a_224_472# net41 0.003942f
C15108 FILLER_0_22_128/a_572_375# vdd 0.001473f
C15109 _348_/a_49_472# mask\[6\] 0.005525f
C15110 _129_ calibrate 0.04134f
C15111 _301_/a_36_472# mask\[8\] 0.016751f
C15112 _161_ net21 0.011799f
C15113 _019_ vdd 0.015401f
C15114 _002_ _089_ 0.002349f
C15115 _163_ _160_ 0.120564f
C15116 _236_/a_36_160# _444_/a_36_151# 0.034413f
C15117 _069_ FILLER_0_15_212/a_36_472# 0.046864f
C15118 cal_itt\[1\] vdd 0.410279f
C15119 net20 FILLER_0_1_204/a_36_472# 0.001278f
C15120 _259_/a_455_68# net37 0.0023f
C15121 _414_/a_36_151# _161_ 0.033054f
C15122 net69 FILLER_0_3_78/a_484_472# 0.002068f
C15123 _088_ FILLER_0_3_172/a_2364_375# 0.002377f
C15124 FILLER_0_9_142/a_36_472# _120_ 0.035902f
C15125 mask\[5\] _346_/a_257_69# 0.001764f
C15126 FILLER_0_18_139/a_1468_375# net23 0.04546f
C15127 fanout70/a_36_113# net53 0.031633f
C15128 net60 _418_/a_2560_156# 0.020147f
C15129 _031_ FILLER_0_2_127/a_124_375# 0.013811f
C15130 FILLER_0_21_206/a_124_375# _434_/a_2665_112# 0.002259f
C15131 _140_ _350_/a_49_472# 0.028997f
C15132 _013_ net55 0.239055f
C15133 FILLER_0_15_212/a_124_375# FILLER_0_15_205/a_124_375# 0.004426f
C15134 FILLER_0_0_130/a_36_472# net13 0.002757f
C15135 _070_ _113_ 0.01052f
C15136 net79 _248_/a_36_68# 0.018243f
C15137 net82 _152_ 0.001896f
C15138 _098_ net71 1.076897f
C15139 _397_/a_36_472# FILLER_0_17_72/a_1468_375# 0.001295f
C15140 _113_ FILLER_0_15_180/a_124_375# 0.001512f
C15141 net54 FILLER_0_21_150/a_36_472# 0.005439f
C15142 _415_/a_36_151# net18 0.015992f
C15143 mask\[4\] net80 0.034957f
C15144 _128_ _120_ 0.053476f
C15145 net62 _417_/a_2560_156# 0.003361f
C15146 _420_/a_36_151# FILLER_0_23_274/a_124_375# 0.059049f
C15147 FILLER_0_6_47/a_1828_472# vdd 0.002735f
C15148 FILLER_0_6_47/a_1380_472# vss 0.001431f
C15149 FILLER_0_9_282/a_36_472# vss 0.002224f
C15150 _429_/a_448_472# net21 0.014792f
C15151 ctln[1] net59 0.053978f
C15152 FILLER_0_7_72/a_2724_472# trim_mask\[0\] 0.006975f
C15153 result[8] FILLER_0_24_290/a_36_472# 0.004676f
C15154 cal_itt\[3\] _062_ 0.009718f
C15155 net35 FILLER_0_22_107/a_484_472# 0.008026f
C15156 net64 net18 1.557441f
C15157 _193_/a_36_160# FILLER_0_13_290/a_36_472# 0.004828f
C15158 _104_ mask\[3\] 0.078406f
C15159 _077_ net14 0.03359f
C15160 _233_/a_36_160# net49 0.035342f
C15161 net63 FILLER_0_22_177/a_1380_472# 0.062289f
C15162 FILLER_0_3_204/a_36_472# net82 0.008268f
C15163 _322_/a_1152_472# _118_ 0.001235f
C15164 _322_/a_124_24# _124_ 0.041337f
C15165 FILLER_0_22_177/a_124_375# _434_/a_1308_423# 0.001064f
C15166 mask\[3\] vss 0.664467f
C15167 FILLER_0_13_212/a_36_472# vss 0.005259f
C15168 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_124_375# 0.012001f
C15169 output45/a_224_472# net17 0.092967f
C15170 net26 FILLER_0_21_28/a_1468_375# 0.041169f
C15171 _131_ FILLER_0_14_107/a_1380_472# 0.01797f
C15172 FILLER_0_12_136/a_484_472# _114_ 0.003953f
C15173 ctlp[1] _420_/a_1308_423# 0.001418f
C15174 FILLER_0_20_107/a_36_472# net14 0.002543f
C15175 _421_/a_2665_112# vss 0.002792f
C15176 _421_/a_2560_156# vdd 0.001862f
C15177 _008_ FILLER_0_17_226/a_124_375# 0.006576f
C15178 cal_count\[3\] net40 0.080767f
C15179 _446_/a_1204_472# net17 0.003628f
C15180 _105_ _295_/a_36_472# 0.031356f
C15181 net9 cal_itt\[1\] 0.028339f
C15182 net24 net14 0.172253f
C15183 net79 _005_ 1.006306f
C15184 vdd FILLER_0_5_148/a_124_375# -0.011369f
C15185 fanout50/a_36_160# net50 0.052685f
C15186 FILLER_0_19_187/a_484_472# vdd 0.011023f
C15187 FILLER_0_19_187/a_36_472# vss 0.001951f
C15188 _104_ output33/a_224_472# 0.032929f
C15189 ctln[0] output7/a_224_472# 0.081823f
C15190 _170_ net59 0.002301f
C15191 _413_/a_36_151# FILLER_0_3_172/a_3172_472# 0.001723f
C15192 FILLER_0_4_177/a_124_375# net76 0.003962f
C15193 ctln[4] FILLER_0_1_212/a_36_472# 0.006408f
C15194 mask\[5\] net35 0.003646f
C15195 _429_/a_1000_472# net22 0.007429f
C15196 _429_/a_796_472# _018_ 0.002291f
C15197 FILLER_0_2_111/a_36_472# vdd 0.033758f
C15198 FILLER_0_2_111/a_1468_375# vss 0.055168f
C15199 _028_ FILLER_0_6_47/a_2364_375# 0.016593f
C15200 net41 _444_/a_1000_472# 0.002179f
C15201 _093_ FILLER_0_17_104/a_1380_472# 0.014431f
C15202 output33/a_224_472# vss 0.05089f
C15203 trimb[4] _452_/a_3129_107# 0.004943f
C15204 FILLER_0_4_91/a_36_472# _160_ 0.007864f
C15205 net15 _394_/a_56_524# 0.006099f
C15206 net52 net49 0.092082f
C15207 _074_ net59 0.030221f
C15208 _443_/a_36_151# _081_ 0.001923f
C15209 _440_/a_796_472# vss 0.001285f
C15210 net10 FILLER_0_1_212/a_124_375# 0.002314f
C15211 FILLER_0_7_72/a_2364_375# _077_ 0.002969f
C15212 net18 _418_/a_1308_423# 0.015651f
C15213 net18 _006_ 0.082256f
C15214 _076_ net59 0.005449f
C15215 _313_/a_67_603# vss 0.016047f
C15216 net82 _443_/a_1308_423# 0.006706f
C15217 FILLER_0_4_197/a_1020_375# vss 0.001981f
C15218 _449_/a_36_151# net74 0.032989f
C15219 _415_/a_2560_156# vss 0.001286f
C15220 _017_ FILLER_0_14_107/a_572_375# 0.003679f
C15221 FILLER_0_21_286/a_36_472# net18 0.18097f
C15222 net70 FILLER_0_14_107/a_1468_375# 0.007955f
C15223 _056_ calibrate 0.00931f
C15224 fanout79/a_36_160# vdd 0.099877f
C15225 _103_ net18 0.11279f
C15226 net44 FILLER_0_20_2/a_572_375# 0.002597f
C15227 _088_ net76 0.214494f
C15228 _050_ FILLER_0_22_128/a_36_472# 0.001098f
C15229 FILLER_0_20_2/a_484_472# vdd 0.001049f
C15230 FILLER_0_5_54/a_932_472# trim_mask\[1\] 0.016187f
C15231 fanout62/a_36_160# vss 0.01343f
C15232 _013_ _216_/a_67_603# 0.006454f
C15233 FILLER_0_16_89/a_932_472# net14 0.014714f
C15234 net27 FILLER_0_9_270/a_124_375# 0.079454f
C15235 _438_/a_448_472# vdd 0.009409f
C15236 _438_/a_36_151# vss 0.014203f
C15237 net41 FILLER_0_21_28/a_124_375# 0.003254f
C15238 ctlp[1] _419_/a_796_472# 0.001178f
C15239 _322_/a_848_380# _062_ 0.001872f
C15240 _255_/a_224_552# _114_ 0.005131f
C15241 _451_/a_2225_156# vdd 0.012404f
C15242 _451_/a_3129_107# vss 0.01f
C15243 mask\[4\] output34/a_224_472# 0.001777f
C15244 output19/a_224_472# _295_/a_36_472# 0.003896f
C15245 _056_ net21 0.484506f
C15246 FILLER_0_5_198/a_484_472# net37 0.009858f
C15247 _111_ _013_ 0.024203f
C15248 ctln[3] net8 0.003753f
C15249 cal net1 0.336092f
C15250 mask\[5\] FILLER_0_19_171/a_1468_375# 0.007169f
C15251 net61 net60 0.059237f
C15252 _063_ _164_ 0.326812f
C15253 result[4] _418_/a_448_472# 0.004918f
C15254 net57 _043_ 1.955053f
C15255 _074_ _122_ 0.300373f
C15256 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1380_472# 0.013276f
C15257 _414_/a_36_151# _056_ 0.00356f
C15258 ctlp[6] net23 0.006951f
C15259 trim_val\[1\] FILLER_0_6_37/a_124_375# 0.007292f
C15260 _370_/a_848_380# FILLER_0_5_136/a_36_472# 0.001177f
C15261 _343_/a_49_472# _137_ 0.001419f
C15262 _074_ FILLER_0_7_233/a_124_375# 0.003081f
C15263 _004_ output28/a_224_472# 0.024204f
C15264 _079_ FILLER_0_5_198/a_572_375# 0.011369f
C15265 _088_ FILLER_0_5_198/a_124_375# 0.001374f
C15266 FILLER_0_19_28/a_124_375# net40 0.047489f
C15267 _219_/a_36_160# _058_ 0.014194f
C15268 net68 FILLER_0_5_54/a_124_375# 0.018458f
C15269 _068_ calibrate 0.110297f
C15270 _076_ _122_ 0.097035f
C15271 _086_ _071_ 0.041029f
C15272 _126_ FILLER_0_13_206/a_124_375# 0.002746f
C15273 _042_ cal_count\[0\] 0.006265f
C15274 _033_ trim_mask\[1\] 0.001251f
C15275 net5 net8 0.001288f
C15276 trim[0] FILLER_0_3_2/a_124_375# 0.020708f
C15277 FILLER_0_20_177/a_124_375# mask\[6\] 0.001158f
C15278 _115_ _315_/a_36_68# 0.001683f
C15279 net36 FILLER_0_15_235/a_124_375# 0.007232f
C15280 net73 _095_ 0.003688f
C15281 _073_ _083_ 0.097365f
C15282 FILLER_0_6_177/a_124_375# vdd 0.017329f
C15283 _028_ FILLER_0_5_72/a_1468_375# 0.00123f
C15284 net1 en 0.068102f
C15285 net50 net14 0.192231f
C15286 _077_ FILLER_0_8_156/a_124_375# 0.00407f
C15287 output42/a_224_472# net67 0.05585f
C15288 result[9] ctlp[2] 0.105977f
C15289 _076_ _227_/a_36_160# 0.004997f
C15290 mask\[5\] net22 0.04021f
C15291 _417_/a_448_472# _006_ 0.068545f
C15292 FILLER_0_7_104/a_572_375# _131_ 0.003031f
C15293 _068_ net21 0.030836f
C15294 _093_ FILLER_0_18_177/a_2812_375# 0.001989f
C15295 _052_ FILLER_0_21_28/a_2812_375# 0.002388f
C15296 ctln[1] FILLER_0_1_266/a_124_375# 0.002958f
C15297 _410_/a_36_68# _453_/a_36_151# 0.002326f
C15298 _133_ _163_ 0.034905f
C15299 FILLER_0_18_37/a_484_472# vdd 0.008381f
C15300 FILLER_0_18_37/a_36_472# vss 0.003026f
C15301 net75 _316_/a_692_472# 0.00138f
C15302 net27 FILLER_0_11_282/a_36_472# 0.001526f
C15303 net50 _164_ 0.080818f
C15304 net63 _019_ 0.004471f
C15305 net39 FILLER_0_8_2/a_124_375# 0.008405f
C15306 _174_ _131_ 0.002314f
C15307 _372_/a_170_472# _385_/a_36_68# 0.009691f
C15308 _317_/a_36_113# FILLER_0_7_233/a_36_472# 0.003531f
C15309 _273_/a_36_68# _070_ 0.013247f
C15310 net16 cal_count\[1\] 0.007291f
C15311 _164_ _382_/a_224_472# 0.011658f
C15312 FILLER_0_9_72/a_36_472# _453_/a_2248_156# 0.013656f
C15313 net73 FILLER_0_18_139/a_484_472# 0.00131f
C15314 ctln[4] _000_ 0.002823f
C15315 input1/a_36_113# net1 0.003795f
C15316 net79 _416_/a_448_472# 0.078357f
C15317 _176_ cal_count\[1\] 0.297763f
C15318 _028_ _363_/a_36_68# 0.015609f
C15319 _037_ net12 0.007817f
C15320 net62 _416_/a_1308_423# 0.002665f
C15321 fanout82/a_36_113# output48/a_224_472# 0.009784f
C15322 _081_ net59 0.185504f
C15323 net70 vdd 0.858299f
C15324 FILLER_0_14_99/a_36_472# _095_ 0.011772f
C15325 ctln[5] _448_/a_1000_472# 0.007584f
C15326 ctlp[7] net24 0.078667f
C15327 net26 _424_/a_36_151# 0.062638f
C15328 trimb[4] vss 0.039934f
C15329 FILLER_0_10_247/a_124_375# vdd 0.040502f
C15330 FILLER_0_9_28/a_1828_472# net16 0.001946f
C15331 _287_/a_36_472# net30 0.005402f
C15332 _096_ mask\[1\] 0.010488f
C15333 result[8] FILLER_0_23_282/a_484_472# 0.001908f
C15334 _093_ _137_ 0.201779f
C15335 FILLER_0_9_105/a_124_375# FILLER_0_10_107/a_36_472# 0.001543f
C15336 vdd _381_/a_36_472# 0.014305f
C15337 FILLER_0_7_72/a_2364_375# net50 0.017301f
C15338 _122_ FILLER_0_5_164/a_484_472# 0.002997f
C15339 vdd FILLER_0_22_107/a_484_472# 0.035591f
C15340 vss FILLER_0_22_107/a_36_472# 0.001514f
C15341 FILLER_0_22_86/a_124_375# net71 0.002239f
C15342 _115_ _308_/a_1084_68# 0.001451f
C15343 FILLER_0_19_55/a_36_472# _052_ 0.019665f
C15344 net36 _280_/a_224_472# 0.001012f
C15345 net65 net59 0.790496f
C15346 FILLER_0_5_72/a_572_375# _164_ 0.005919f
C15347 FILLER_0_10_107/a_124_375# vdd 0.045066f
C15348 FILLER_0_12_50/a_124_375# _067_ 0.011869f
C15349 FILLER_0_16_255/a_36_472# _045_ 0.001653f
C15350 FILLER_0_15_228/a_124_375# vdd 0.013701f
C15351 _053_ net15 0.041871f
C15352 trim_mask\[0\] FILLER_0_10_94/a_572_375# 0.003359f
C15353 net55 FILLER_0_11_78/a_572_375# 0.002321f
C15354 FILLER_0_6_239/a_124_375# _316_/a_124_24# 0.003524f
C15355 net16 FILLER_0_17_38/a_36_472# 0.014381f
C15356 FILLER_0_5_164/a_36_472# _163_ 0.001777f
C15357 net16 _392_/a_36_68# 0.002191f
C15358 input4/a_36_68# vss 0.058179f
C15359 _444_/a_1204_472# net17 0.021952f
C15360 FILLER_0_2_93/a_36_472# net69 0.010977f
C15361 _111_ net71 0.002668f
C15362 mask\[3\] FILLER_0_16_154/a_1020_375# 0.001996f
C15363 net15 FILLER_0_5_54/a_1380_472# 0.047774f
C15364 _425_/a_796_472# _122_ 0.001701f
C15365 _425_/a_36_151# _123_ 0.006319f
C15366 _425_/a_1000_472# calibrate 0.027245f
C15367 FILLER_0_9_142/a_124_375# vdd 0.015952f
C15368 _328_/a_36_113# net14 0.002272f
C15369 FILLER_0_17_226/a_124_375# _093_ 0.001604f
C15370 _072_ _311_/a_3220_473# 0.001995f
C15371 _081_ _122_ 2.557248f
C15372 _152_ calibrate 0.020369f
C15373 _424_/a_2665_112# _012_ 0.01024f
C15374 mask\[5\] FILLER_0_20_177/a_484_472# 0.016114f
C15375 net38 FILLER_0_15_10/a_124_375# 0.047331f
C15376 _033_ _444_/a_2665_112# 0.004024f
C15377 _053_ FILLER_0_6_90/a_572_375# 0.073688f
C15378 _306_/a_36_68# _085_ 0.00755f
C15379 _024_ _435_/a_1308_423# 0.002661f
C15380 _417_/a_1000_472# vss 0.001822f
C15381 FILLER_0_8_138/a_36_472# _313_/a_67_603# 0.005759f
C15382 FILLER_0_9_72/a_124_375# vss 0.047932f
C15383 FILLER_0_9_72/a_572_375# vdd -0.014642f
C15384 FILLER_0_20_98/a_36_472# vss 0.00206f
C15385 trim_mask\[2\] net69 0.051795f
C15386 _304_/a_224_472# mask\[9\] 0.003125f
C15387 mask\[5\] vdd 0.79138f
C15388 net63 FILLER_0_19_187/a_484_472# 0.020823f
C15389 _121_ _314_/a_224_472# 0.00323f
C15390 _115_ FILLER_0_10_78/a_1380_472# 0.051132f
C15391 net18 _416_/a_1288_156# 0.001147f
C15392 _276_/a_36_160# _093_ 0.019339f
C15393 _115_ _219_/a_36_160# 0.001218f
C15394 _081_ _169_ 0.260462f
C15395 _061_ vss 0.046487f
C15396 FILLER_0_5_72/a_1468_375# net47 0.005049f
C15397 FILLER_0_21_28/a_572_375# net17 0.001455f
C15398 mask\[8\] FILLER_0_22_86/a_1380_472# 0.012151f
C15399 net35 FILLER_0_22_86/a_932_472# 0.007806f
C15400 fanout66/a_36_113# vss 0.014789f
C15401 FILLER_0_13_290/a_36_472# _416_/a_36_151# 0.001723f
C15402 _431_/a_36_151# _334_/a_36_160# 0.032942f
C15403 _453_/a_1308_423# vss 0.003012f
C15404 FILLER_0_13_212/a_932_472# _043_ 0.014431f
C15405 _311_/a_254_473# vdd 0.001207f
C15406 cal_count\[2\] FILLER_0_15_2/a_124_375# 0.033559f
C15407 _323_/a_36_113# _426_/a_2248_156# 0.001661f
C15408 _015_ _426_/a_1308_423# 0.029444f
C15409 _114_ _120_ 0.334426f
C15410 _064_ net17 0.108825f
C15411 _138_ net21 0.003242f
C15412 _141_ FILLER_0_17_161/a_36_472# 0.011708f
C15413 net65 net64 0.119915f
C15414 _001_ vss 0.004381f
C15415 _000_ FILLER_0_3_221/a_1020_375# 0.016709f
C15416 FILLER_0_1_98/a_124_375# _442_/a_2665_112# 0.003045f
C15417 _328_/a_36_113# _428_/a_36_151# 0.030244f
C15418 _114_ FILLER_0_13_142/a_1020_375# 0.001964f
C15419 _337_/a_49_472# _137_ 0.046633f
C15420 _189_/a_67_603# FILLER_0_13_228/a_36_472# 0.005759f
C15421 ctlp[1] net77 0.716304f
C15422 net56 mask\[2\] 0.090254f
C15423 _098_ _437_/a_1000_472# 0.007963f
C15424 FILLER_0_11_142/a_124_375# FILLER_0_11_135/a_124_375# 0.004426f
C15425 _144_ _140_ 0.415736f
C15426 FILLER_0_10_78/a_484_472# net52 0.004421f
C15427 net54 FILLER_0_22_128/a_484_472# 0.055436f
C15428 net32 _421_/a_1308_423# 0.005394f
C15429 FILLER_0_17_72/a_2276_472# _136_ 0.055635f
C15430 net17 net42 0.056318f
C15431 _131_ FILLER_0_16_115/a_124_375# 0.016715f
C15432 net81 FILLER_0_15_212/a_1020_375# 0.006974f
C15433 _077_ _439_/a_2665_112# 0.035688f
C15434 FILLER_0_3_204/a_36_472# net21 0.01535f
C15435 vdd _433_/a_448_472# 0.003821f
C15436 vss _433_/a_36_151# 0.00618f
C15437 mask\[0\] _429_/a_448_472# 0.061449f
C15438 _448_/a_1000_472# net59 0.007647f
C15439 ctln[5] FILLER_0_0_198/a_36_472# 0.012298f
C15440 _101_ vss 0.05721f
C15441 _251_/a_244_472# net4 0.005273f
C15442 FILLER_0_11_101/a_484_472# vss 0.003923f
C15443 FILLER_0_3_172/a_124_375# net22 0.01308f
C15444 _128_ _125_ 0.017316f
C15445 _027_ _438_/a_36_151# 0.010763f
C15446 _150_ _438_/a_1308_423# 0.001472f
C15447 FILLER_0_20_98/a_124_375# _437_/a_36_151# 0.059049f
C15448 FILLER_0_18_100/a_36_472# mask\[9\] 0.005719f
C15449 FILLER_0_13_212/a_1468_375# FILLER_0_12_220/a_572_375# 0.05841f
C15450 mask\[4\] FILLER_0_18_139/a_1380_472# 0.003851f
C15451 FILLER_0_18_107/a_484_472# FILLER_0_17_104/a_932_472# 0.026657f
C15452 _053_ FILLER_0_5_212/a_36_472# 0.007052f
C15453 _052_ _424_/a_796_472# 0.002115f
C15454 FILLER_0_16_57/a_124_375# _131_ 0.012982f
C15455 _072_ vss 0.439154f
C15456 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_572_375# 0.001597f
C15457 mask\[1\] FILLER_0_15_180/a_484_472# 0.003594f
C15458 _399_/a_224_472# _179_ 0.002288f
C15459 FILLER_0_11_142/a_572_375# _076_ 0.031784f
C15460 _395_/a_36_488# _085_ 0.020572f
C15461 net81 fanout80/a_36_113# 0.097873f
C15462 output27/a_224_472# result[0] 0.031252f
C15463 net16 _120_ 0.009918f
C15464 net80 FILLER_0_20_169/a_124_375# 0.054969f
C15465 net76 FILLER_0_6_177/a_572_375# 0.073022f
C15466 _176_ _120_ 0.169846f
C15467 _176_ _038_ 0.039948f
C15468 net23 FILLER_0_21_150/a_124_375# 0.045928f
C15469 net19 _417_/a_2665_112# 0.042961f
C15470 FILLER_0_5_109/a_124_375# net47 0.010784f
C15471 FILLER_0_5_128/a_124_375# vdd 0.008803f
C15472 FILLER_0_19_195/a_124_375# vss 0.020433f
C15473 FILLER_0_19_195/a_36_472# vdd 0.094409f
C15474 FILLER_0_7_104/a_1020_375# _133_ 0.008772f
C15475 _328_/a_36_113# FILLER_0_11_109/a_36_472# 0.0161f
C15476 _132_ FILLER_0_18_107/a_1828_472# 0.045833f
C15477 _413_/a_36_151# FILLER_0_4_197/a_484_472# 0.001512f
C15478 _093_ FILLER_0_17_72/a_1468_375# 0.005785f
C15479 _411_/a_2665_112# vss 0.00238f
C15480 _126_ _390_/a_36_68# 0.044675f
C15481 _011_ _009_ 0.035129f
C15482 _008_ _418_/a_36_151# 0.016984f
C15483 _096_ mask\[0\] 0.052773f
C15484 _014_ vss 0.034646f
C15485 _075_ _072_ 0.024301f
C15486 _085_ FILLER_0_13_142/a_1468_375# 0.001153f
C15487 net34 _435_/a_2248_156# 0.01519f
C15488 FILLER_0_5_206/a_124_375# _081_ 0.031751f
C15489 cal_count\[3\] FILLER_0_9_72/a_484_472# 0.004129f
C15490 FILLER_0_14_181/a_124_375# _098_ 0.005696f
C15491 trimb[0] output43/a_224_472# 0.043402f
C15492 vss FILLER_0_13_72/a_484_472# 0.008682f
C15493 FILLER_0_7_72/a_2724_472# FILLER_0_6_90/a_572_375# 0.001684f
C15494 FILLER_0_19_125/a_36_472# _433_/a_36_151# 0.059367f
C15495 result[5] vdd 0.142481f
C15496 output16/a_224_472# _447_/a_36_151# 0.200384f
C15497 _365_/a_36_68# vdd 0.004308f
C15498 fanout69/a_36_113# _160_ 0.005933f
C15499 result[7] result[8] 0.201281f
C15500 _343_/a_257_69# _137_ 0.003494f
C15501 _429_/a_36_151# FILLER_0_15_212/a_572_375# 0.059049f
C15502 net65 FILLER_0_1_266/a_124_375# 0.002654f
C15503 net27 FILLER_0_15_235/a_572_375# 0.001554f
C15504 ctln[5] net11 0.004569f
C15505 _150_ net36 0.108945f
C15506 FILLER_0_18_107/a_3172_472# FILLER_0_19_134/a_124_375# 0.001723f
C15507 _097_ FILLER_0_15_180/a_36_472# 0.005242f
C15508 cal_count\[2\] _452_/a_36_151# 0.006982f
C15509 FILLER_0_17_38/a_36_472# _041_ 0.003805f
C15510 net74 FILLER_0_11_124/a_124_375# 0.047331f
C15511 net81 FILLER_0_15_205/a_36_472# 0.081574f
C15512 FILLER_0_2_101/a_36_472# net14 0.051153f
C15513 _053_ FILLER_0_7_104/a_36_472# 0.01752f
C15514 _063_ _378_/a_224_472# 0.002323f
C15515 _031_ vss 0.18315f
C15516 mask\[9\] _438_/a_2560_156# 0.008709f
C15517 net72 _424_/a_448_472# 0.011745f
C15518 net27 vdd 0.88294f
C15519 output38/a_224_472# net17 0.04454f
C15520 _064_ _446_/a_1308_423# 0.001728f
C15521 net52 FILLER_0_5_54/a_1468_375# 0.003649f
C15522 _114_ state\[2\] 0.528838f
C15523 mask\[4\] output18/a_224_472# 0.017718f
C15524 _074_ FILLER_0_5_181/a_36_472# 0.002385f
C15525 _005_ net19 0.033451f
C15526 _015_ FILLER_0_8_239/a_36_472# 0.002627f
C15527 _093_ FILLER_0_19_142/a_36_472# 0.002415f
C15528 _415_/a_1308_423# result[1] 0.00761f
C15529 _320_/a_36_472# net22 0.005964f
C15530 output20/a_224_472# vdd 0.09529f
C15531 output22/a_224_472# mask\[7\] 0.05527f
C15532 net52 _442_/a_1204_472# 0.005558f
C15533 _384_/a_224_472# _168_ 0.003461f
C15534 net75 FILLER_0_6_239/a_124_375# 0.013962f
C15535 FILLER_0_18_177/a_1828_472# vss -0.001107f
C15536 FILLER_0_18_177/a_2276_472# vdd 0.005211f
C15537 _005_ _416_/a_796_472# 0.009162f
C15538 FILLER_0_2_101/a_124_375# trim_mask\[3\] 0.033692f
C15539 net38 _033_ 0.03598f
C15540 _115_ FILLER_0_10_107/a_484_472# 0.017642f
C15541 FILLER_0_14_81/a_36_472# _177_ 0.004294f
C15542 _441_/a_448_472# _168_ 0.033059f
C15543 net20 FILLER_0_3_221/a_1380_472# 0.008749f
C15544 FILLER_0_9_60/a_36_472# vdd 0.08419f
C15545 FILLER_0_9_60/a_572_375# vss 0.022532f
C15546 output24/a_224_472# _436_/a_448_472# 0.009204f
C15547 net66 FILLER_0_5_54/a_932_472# 0.001419f
C15548 _415_/a_1000_472# net18 0.006558f
C15549 FILLER_0_13_212/a_124_375# FILLER_0_13_206/a_124_375# 0.005439f
C15550 net18 _419_/a_2665_112# 0.0371f
C15551 FILLER_0_21_206/a_124_375# mask\[6\] 0.008881f
C15552 ctlp[1] _421_/a_448_472# 0.011026f
C15553 net80 _138_ 0.002053f
C15554 net69 _441_/a_2560_156# 0.002904f
C15555 mask\[0\] _056_ 0.001878f
C15556 FILLER_0_17_104/a_484_472# net14 0.004272f
C15557 _094_ vss 0.24519f
C15558 FILLER_0_17_218/a_572_375# vss 0.078608f
C15559 FILLER_0_17_218/a_36_472# vdd 0.084913f
C15560 FILLER_0_3_172/a_124_375# vdd 0.010886f
C15561 _028_ _053_ 0.891578f
C15562 _425_/a_2665_112# vdd 0.012933f
C15563 output22/a_224_472# net80 0.00955f
C15564 ctlp[5] output23/a_224_472# 0.005152f
C15565 FILLER_0_9_28/a_1468_375# _054_ 0.005381f
C15566 net75 net19 1.345314f
C15567 net45 net17 0.192181f
C15568 mask\[7\] FILLER_0_22_128/a_2276_472# 0.004398f
C15569 _069_ _429_/a_1000_472# 0.029501f
C15570 net41 _450_/a_2225_156# 0.024042f
C15571 _432_/a_2665_112# vss 0.002577f
C15572 _142_ FILLER_0_18_107/a_2724_472# 0.001549f
C15573 cal_itt\[2\] _413_/a_2248_156# 0.002527f
C15574 FILLER_0_14_181/a_124_375# FILLER_0_15_180/a_124_375# 0.026339f
C15575 net53 _427_/a_2560_156# 0.004594f
C15576 FILLER_0_22_128/a_36_472# _022_ 0.001541f
C15577 net28 fanout79/a_36_160# 0.036675f
C15578 trimb[1] FILLER_0_18_2/a_932_472# 0.011513f
C15579 _423_/a_36_151# FILLER_0_23_44/a_1020_375# 0.059049f
C15580 _350_/a_49_472# _049_ 0.025442f
C15581 _013_ FILLER_0_18_61/a_124_375# 0.016976f
C15582 _394_/a_56_524# FILLER_0_15_59/a_484_472# 0.001033f
C15583 _394_/a_718_524# FILLER_0_15_59/a_572_375# 0.001447f
C15584 _020_ _136_ 0.022753f
C15585 _448_/a_2560_156# net22 0.00766f
C15586 _233_/a_36_160# net40 0.001875f
C15587 _098_ FILLER_0_15_212/a_1468_375# 0.008327f
C15588 _429_/a_36_151# FILLER_0_15_205/a_124_375# 0.059049f
C15589 _428_/a_2248_156# net74 0.072805f
C15590 net50 _439_/a_2665_112# 0.007973f
C15591 _079_ FILLER_0_6_231/a_484_472# 0.008159f
C15592 net31 net34 0.080525f
C15593 _138_ mask\[1\] 0.085445f
C15594 _141_ FILLER_0_18_139/a_1468_375# 0.005239f
C15595 _331_/a_448_472# vdd 0.001343f
C15596 _098_ FILLER_0_16_154/a_1380_472# 0.00417f
C15597 _394_/a_56_524# net74 0.005616f
C15598 net54 FILLER_0_19_142/a_36_472# 0.07544f
C15599 _176_ _175_ 0.054439f
C15600 _104_ ctlp[3] 0.025066f
C15601 _363_/a_36_68# _154_ 0.149319f
C15602 _035_ _379_/a_36_472# 0.002226f
C15603 _261_/a_36_160# vdd 0.0109f
C15604 FILLER_0_11_101/a_36_472# FILLER_0_13_100/a_124_375# 0.001436f
C15605 _098_ _434_/a_448_472# 0.015893f
C15606 net48 _317_/a_36_113# 0.018494f
C15607 ctlp[3] vss 0.037106f
C15608 net2 _425_/a_36_151# 0.012359f
C15609 _105_ _092_ 0.006701f
C15610 _106_ mask\[3\] 0.249479f
C15611 _394_/a_2215_68# _095_ 0.001134f
C15612 FILLER_0_22_86/a_932_472# vdd 0.001826f
C15613 mask\[5\] net63 0.112147f
C15614 trim_val\[4\] _170_ 0.281942f
C15615 FILLER_0_4_152/a_124_375# _386_/a_124_24# 0.010472f
C15616 _114_ _311_/a_2180_473# 0.00515f
C15617 _199_/a_36_160# vdd 0.036579f
C15618 FILLER_0_19_125/a_124_375# vss 0.001974f
C15619 FILLER_0_22_128/a_3172_472# vss 0.006339f
C15620 _104_ net78 0.049954f
C15621 _132_ _428_/a_1308_423# 0.027389f
C15622 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_484_472# 0.013276f
C15623 net35 _435_/a_448_472# 0.007865f
C15624 FILLER_0_5_109/a_124_375# _154_ 0.058658f
C15625 _020_ fanout70/a_36_113# 0.001266f
C15626 FILLER_0_16_73/a_572_375# FILLER_0_17_72/a_572_375# 0.026339f
C15627 net81 net37 0.18149f
C15628 net59 net11 0.016998f
C15629 net78 vss 0.167812f
C15630 _053_ _257_/a_244_68# 0.001138f
C15631 _442_/a_2665_112# net14 0.011563f
C15632 _050_ vss 0.26237f
C15633 net37 _160_ 0.003563f
C15634 _320_/a_36_472# vdd 0.086964f
C15635 _445_/a_1204_472# _034_ 0.003057f
C15636 FILLER_0_0_198/a_124_375# net11 0.071885f
C15637 net15 _447_/a_448_472# 0.001766f
C15638 net49 net40 0.093233f
C15639 net52 FILLER_0_6_79/a_124_375# 0.010099f
C15640 net82 FILLER_0_3_172/a_1828_472# 0.004472f
C15641 FILLER_0_8_263/a_36_472# vss 0.001089f
C15642 FILLER_0_8_127/a_36_472# _322_/a_124_24# 0.00171f
C15643 _072_ _071_ 0.296543f
C15644 vss FILLER_0_14_235/a_572_375# 0.017196f
C15645 _442_/a_2248_156# trim_mask\[3\] 0.003039f
C15646 FILLER_0_7_72/a_3172_472# vdd 0.003913f
C15647 FILLER_0_3_172/a_932_472# net65 0.002604f
C15648 FILLER_0_4_197/a_36_472# _079_ 0.002448f
C15649 _446_/a_2560_156# vdd 0.003959f
C15650 _446_/a_2665_112# vss 0.001781f
C15651 ctln[1] ctln[4] 0.002283f
C15652 _028_ FILLER_0_7_72/a_2724_472# 0.001777f
C15653 FILLER_0_10_37/a_36_472# FILLER_0_8_37/a_124_375# 0.001512f
C15654 ctlp[3] _107_ 0.132316f
C15655 net72 _404_/a_36_472# 0.019911f
C15656 _210_/a_255_603# vss 0.001246f
C15657 _127_ _126_ 0.398279f
C15658 _094_ _195_/a_67_603# 0.043278f
C15659 _214_/a_36_160# vss 0.007045f
C15660 net58 FILLER_0_8_247/a_1468_375# 0.001669f
C15661 _443_/a_1000_472# vss 0.031435f
C15662 FILLER_0_22_86/a_36_472# _437_/a_36_151# 0.059367f
C15663 _009_ FILLER_0_23_274/a_124_375# 0.010723f
C15664 FILLER_0_12_136/a_1380_472# net23 0.011488f
C15665 _119_ _162_ 0.036701f
C15666 comp FILLER_0_15_2/a_124_375# 0.034135f
C15667 _432_/a_2248_156# vdd 0.02369f
C15668 net20 FILLER_0_13_212/a_1380_472# 0.006746f
C15669 cal_count\[3\] _188_ 0.048745f
C15670 _448_/a_2665_112# vss 0.009029f
C15671 _446_/a_36_151# net66 0.034846f
C15672 _053_ net47 0.011652f
C15673 result[7] _093_ 0.001096f
C15674 FILLER_0_17_72/a_124_375# FILLER_0_17_64/a_124_375# 0.003732f
C15675 _126_ FILLER_0_11_135/a_36_472# 0.002321f
C15676 mask\[1\] _113_ 0.032744f
C15677 net63 FILLER_0_19_195/a_36_472# 0.030832f
C15678 _122_ _163_ 0.156898f
C15679 _425_/a_36_151# FILLER_0_8_247/a_36_472# 0.02628f
C15680 _425_/a_1308_423# FILLER_0_8_247/a_1020_375# 0.001064f
C15681 FILLER_0_9_223/a_124_375# _077_ 0.008762f
C15682 _423_/a_1308_423# vdd 0.00335f
C15683 _423_/a_448_472# vss 0.002481f
C15684 FILLER_0_16_57/a_1020_375# net55 0.003303f
C15685 FILLER_0_16_57/a_484_472# net72 0.017841f
C15686 _119_ _131_ 0.073868f
C15687 fanout66/a_36_113# _036_ 0.014556f
C15688 FILLER_0_5_54/a_1380_472# net47 0.003924f
C15689 net68 _453_/a_1000_472# 0.001816f
C15690 output36/a_224_472# _045_ 0.041236f
C15691 net57 _428_/a_1204_472# 0.015233f
C15692 _105_ net61 0.020753f
C15693 _086_ _375_/a_36_68# 0.038443f
C15694 net81 _139_ 0.001762f
C15695 FILLER_0_7_72/a_36_472# _028_ 0.020625f
C15696 net62 net29 0.082455f
C15697 _118_ _311_/a_3740_473# 0.001244f
C15698 FILLER_0_16_89/a_484_472# _136_ 0.032722f
C15699 FILLER_0_7_195/a_124_375# _055_ 0.001597f
C15700 fanout60/a_36_160# FILLER_0_17_282/a_36_472# 0.002647f
C15701 net47 FILLER_0_5_164/a_124_375# 0.011983f
C15702 _126_ FILLER_0_11_101/a_36_472# 0.062336f
C15703 FILLER_0_18_2/a_2724_472# net55 0.007511f
C15704 FILLER_0_15_72/a_124_375# cal_count\[1\] 0.00816f
C15705 trimb[1] net55 0.017528f
C15706 trim_val\[4\] FILLER_0_5_164/a_484_472# 0.00172f
C15707 ctln[7] output15/a_224_472# 0.00838f
C15708 _169_ _163_ 0.013133f
C15709 FILLER_0_5_206/a_36_472# net59 0.060133f
C15710 _086_ FILLER_0_11_124/a_36_472# 0.010729f
C15711 _326_/a_36_160# _131_ 0.023688f
C15712 FILLER_0_17_72/a_484_472# vss 0.005334f
C15713 _181_ _402_/a_728_93# 0.064373f
C15714 _134_ FILLER_0_10_107/a_484_472# 0.020725f
C15715 net22 _435_/a_448_472# 0.001929f
C15716 _093_ _334_/a_36_160# 0.014676f
C15717 FILLER_0_5_136/a_124_375# vdd 0.035814f
C15718 net31 net36 0.00943f
C15719 mask\[0\] _138_ 0.22533f
C15720 FILLER_0_12_20/a_124_375# _039_ 0.004669f
C15721 _115_ _058_ 0.038308f
C15722 FILLER_0_16_89/a_124_375# _040_ 0.006315f
C15723 net41 trim[3] 0.005906f
C15724 FILLER_0_4_107/a_36_472# _369_/a_36_68# 0.001709f
C15725 FILLER_0_4_107/a_1020_375# _158_ 0.003535f
C15726 net27 _283_/a_36_472# 0.023243f
C15727 _132_ FILLER_0_17_104/a_1468_375# 0.051996f
C15728 FILLER_0_3_78/a_124_375# _164_ 0.023555f
C15729 _427_/a_1000_472# vss 0.012657f
C15730 net17 _450_/a_2449_156# 0.05017f
C15731 trim_mask\[1\] vss 0.449335f
C15732 net41 _402_/a_718_527# 0.019628f
C15733 _372_/a_170_472# _070_ 0.024545f
C15734 output16/a_224_472# vss 0.009875f
C15735 _436_/a_36_151# FILLER_0_22_107/a_572_375# 0.059049f
C15736 net76 FILLER_0_3_172/a_572_375# 0.003315f
C15737 _085_ vdd 0.227153f
C15738 FILLER_0_12_220/a_484_472# _070_ 0.004091f
C15739 FILLER_0_16_107/a_124_375# _093_ 0.003941f
C15740 net63 FILLER_0_18_177/a_2276_472# 0.012025f
C15741 net8 FILLER_0_0_266/a_124_375# 0.001181f
C15742 net52 _440_/a_2560_156# 0.004924f
C15743 fanout74/a_36_113# net23 0.005294f
C15744 _053_ net74 0.09773f
C15745 _155_ FILLER_0_4_91/a_572_375# 0.004038f
C15746 net73 _098_ 0.004745f
C15747 FILLER_0_18_2/a_2724_472# net17 0.017841f
C15748 trim_val\[0\] _220_/a_67_603# 0.005346f
C15749 _095_ FILLER_0_13_72/a_484_472# 0.027852f
C15750 trimb[1] net17 0.084269f
C15751 _452_/a_836_156# _041_ 0.001052f
C15752 FILLER_0_15_142/a_36_472# vdd 0.106034f
C15753 _408_/a_1936_472# vdd 0.022538f
C15754 _250_/a_36_68# net23 0.002628f
C15755 net41 _445_/a_2665_112# 0.056125f
C15756 net61 output19/a_224_472# 0.077658f
C15757 net49 _440_/a_2560_156# 0.011378f
C15758 net39 _444_/a_448_472# 0.002089f
C15759 _157_ vss 0.039512f
C15760 FILLER_0_7_59/a_36_472# trim_val\[0\] 0.003014f
C15761 ctln[1] FILLER_0_3_221/a_1020_375# 0.001554f
C15762 FILLER_0_5_206/a_36_472# _122_ 0.003017f
C15763 net63 FILLER_0_17_218/a_36_472# 0.003889f
C15764 FILLER_0_15_150/a_36_472# _136_ 0.002967f
C15765 _258_/a_36_160# vdd 0.00617f
C15766 net72 _217_/a_36_160# 0.068583f
C15767 trim_val\[4\] net65 0.015549f
C15768 _447_/a_2665_112# vss 0.012813f
C15769 FILLER_0_16_89/a_1380_472# net36 0.001657f
C15770 fanout77/a_36_113# _419_/a_36_151# 0.002361f
C15771 ctln[2] net8 0.057281f
C15772 _373_/a_1254_68# _090_ 0.001326f
C15773 _091_ FILLER_0_19_171/a_1468_375# 0.002731f
C15774 FILLER_0_16_57/a_932_472# cal_count\[1\] 0.002217f
C15775 mask\[9\] vss 0.649041f
C15776 _053_ _372_/a_2034_472# 0.00181f
C15777 _065_ fanout68/a_36_113# 0.005586f
C15778 _115_ _389_/a_36_148# 0.029505f
C15779 FILLER_0_10_37/a_124_375# cal_count\[0\] 0.016543f
C15780 _176_ _125_ 0.089769f
C15781 result[2] _193_/a_36_160# 0.040932f
C15782 _077_ FILLER_0_9_72/a_1468_375# 0.008273f
C15783 FILLER_0_18_107/a_1020_375# mask\[9\] 0.005758f
C15784 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_124_375# 0.026339f
C15785 _405_/a_67_603# cal_count\[2\] 0.021962f
C15786 net60 net62 0.002144f
C15787 net68 _441_/a_36_151# 0.031891f
C15788 FILLER_0_18_100/a_124_375# net14 0.04037f
C15789 state\[0\] _274_/a_1164_497# 0.002914f
C15790 FILLER_0_17_218/a_36_472# _069_ 0.001246f
C15791 net20 _429_/a_2248_156# 0.027661f
C15792 _444_/a_2665_112# _054_ 0.003576f
C15793 net18 FILLER_0_9_282/a_124_375# 0.024657f
C15794 _077_ _453_/a_1204_472# 0.011124f
C15795 _440_/a_1308_423# _160_ 0.002554f
C15796 net71 _437_/a_448_472# 0.060858f
C15797 _155_ FILLER_0_7_104/a_572_375# 0.002336f
C15798 output27/a_224_472# fanout65/a_36_113# 0.011564f
C15799 _435_/a_448_472# vdd 0.029967f
C15800 _091_ net22 0.031921f
C15801 net50 _376_/a_36_160# 0.018407f
C15802 net38 _444_/a_36_151# 0.009033f
C15803 _410_/a_36_68# _042_ 0.041079f
C15804 net75 output28/a_224_472# 0.00151f
C15805 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_484_472# 0.026657f
C15806 net53 FILLER_0_17_142/a_484_472# 0.001286f
C15807 mask\[0\] _113_ 0.01678f
C15808 ctln[0] trim[3] 0.216084f
C15809 trim_mask\[1\] FILLER_0_5_88/a_124_375# 0.072632f
C15810 _053_ _154_ 0.41707f
C15811 _125_ _124_ 0.085897f
C15812 net32 output35/a_224_472# 0.072991f
C15813 _449_/a_2248_156# net55 0.052445f
C15814 _443_/a_448_472# _032_ 0.036717f
C15815 _422_/a_1204_472# _109_ 0.001807f
C15816 _110_ net35 0.053239f
C15817 _093_ _437_/a_36_151# 0.056554f
C15818 FILLER_0_15_142/a_484_472# net53 0.044267f
C15819 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_36_472# 0.026657f
C15820 _083_ FILLER_0_3_221/a_484_472# 0.02695f
C15821 _430_/a_448_472# net21 0.03842f
C15822 trim_mask\[2\] FILLER_0_4_91/a_484_472# 0.0022f
C15823 _444_/a_2665_112# vss 0.002271f
C15824 _444_/a_2560_156# vdd 0.025035f
C15825 mask\[4\] net56 0.006006f
C15826 _424_/a_2248_156# net36 0.017101f
C15827 cal_count\[3\] _186_ 0.012453f
C15828 net25 FILLER_0_23_60/a_36_472# 0.005618f
C15829 trim_val\[4\] _443_/a_448_472# 0.038063f
C15830 _086_ _374_/a_244_472# 0.001496f
C15831 _062_ vdd 0.393862f
C15832 output11/a_224_472# net75 0.015211f
C15833 mask\[3\] fanout53/a_36_160# 0.001205f
C15834 net74 FILLER_0_2_127/a_36_472# 0.001261f
C15835 net20 _260_/a_244_472# 0.001593f
C15836 _079_ _083_ 0.872842f
C15837 _088_ _078_ 0.047558f
C15838 _119_ _074_ 0.153267f
C15839 net78 _419_/a_1000_472# 0.040603f
C15840 FILLER_0_18_2/a_3260_375# vdd 0.046682f
C15841 FILLER_0_9_28/a_572_375# net50 0.002807f
C15842 ctln[4] net65 0.020799f
C15843 net38 _452_/a_3129_107# 0.005269f
C15844 FILLER_0_20_2/a_484_472# net43 0.005543f
C15845 _438_/a_2665_112# net14 0.026903f
C15846 ctln[5] ctln[6] 0.017291f
C15847 _119_ _076_ 0.083673f
C15848 FILLER_0_15_150/a_36_472# net53 0.016925f
C15849 mask\[8\] _437_/a_2560_156# 0.001171f
C15850 _130_ _131_ 0.005955f
C15851 FILLER_0_21_28/a_1916_375# vdd -0.009753f
C15852 ctln[8] vdd 0.125219f
C15853 FILLER_0_11_78/a_484_472# vss 0.004063f
C15854 _432_/a_2248_156# net63 0.047337f
C15855 net20 fanout63/a_36_160# 0.084165f
C15856 FILLER_0_21_142/a_572_375# vss 0.097474f
C15857 FILLER_0_8_127/a_124_375# _070_ 0.003265f
C15858 net16 cal_count\[2\] 0.041089f
C15859 net82 FILLER_0_4_213/a_484_472# 0.002255f
C15860 _232_/a_67_603# FILLER_0_6_47/a_36_472# 0.010206f
C15861 net67 FILLER_0_9_60/a_484_472# 0.001345f
C15862 _144_ _049_ 0.100508f
C15863 _176_ cal_count\[2\] 0.005783f
C15864 FILLER_0_4_107/a_1468_375# trim_mask\[4\] 0.00157f
C15865 _086_ _070_ 0.123033f
C15866 FILLER_0_19_55/a_124_375# FILLER_0_18_53/a_484_472# 0.001684f
C15867 net20 _291_/a_36_160# 0.002375f
C15868 _055_ _060_ 0.181186f
C15869 net27 FILLER_0_12_236/a_572_375# 0.083731f
C15870 net54 _437_/a_36_151# 0.019307f
C15871 mask\[3\] _098_ 0.026156f
C15872 _053_ _079_ 0.007118f
C15873 _058_ _134_ 0.034211f
C15874 _131_ _129_ 0.017222f
C15875 FILLER_0_4_107/a_1468_375# net47 0.012534f
C15876 net48 net59 0.015963f
C15877 net81 _429_/a_1308_423# 0.008913f
C15878 FILLER_0_5_164/a_36_472# net37 0.008378f
C15879 net4 FILLER_0_6_231/a_124_375# 0.002212f
C15880 FILLER_0_2_171/a_36_472# net22 0.081357f
C15881 FILLER_0_6_90/a_36_472# vss 0.001409f
C15882 FILLER_0_6_90/a_484_472# vdd 0.003146f
C15883 _139_ FILLER_0_15_180/a_572_375# 0.022254f
C15884 _083_ cal_itt\[1\] 0.046464f
C15885 result[5] net77 0.142532f
C15886 _418_/a_2665_112# vdd 0.028061f
C15887 mask\[5\] _140_ 0.103728f
C15888 FILLER_0_18_177/a_3172_472# FILLER_0_18_209/a_36_472# 0.013276f
C15889 fanout74/a_36_113# FILLER_0_3_142/a_36_472# 0.016516f
C15890 _091_ vdd 1.011371f
C15891 FILLER_0_1_98/a_124_375# vdd 0.036865f
C15892 FILLER_0_16_73/a_572_375# vdd 0.005054f
C15893 FILLER_0_7_72/a_1828_472# _163_ 0.002095f
C15894 net35 net14 0.040959f
C15895 FILLER_0_17_72/a_1380_472# _150_ 0.014154f
C15896 net52 FILLER_0_9_72/a_484_472# 0.049391f
C15897 _100_ FILLER_0_12_236/a_484_472# 0.00195f
C15898 net70 _451_/a_36_151# 0.04524f
C15899 FILLER_0_13_142/a_36_472# net23 0.003007f
C15900 _445_/a_2560_156# net17 0.010829f
C15901 output37/a_224_472# _425_/a_2248_156# 0.00114f
C15902 net39 net44 0.0112f
C15903 ctlp[1] FILLER_0_24_290/a_36_472# 0.037615f
C15904 trim[1] vdd 0.089624f
C15905 _114_ _043_ 0.071339f
C15906 _057_ net57 0.873864f
C15907 _287_/a_36_472# _006_ 0.00121f
C15908 _425_/a_1308_423# net37 0.002601f
C15909 _408_/a_728_93# _450_/a_2225_156# 0.00128f
C15910 _141_ FILLER_0_21_150/a_124_375# 0.02192f
C15911 _412_/a_1308_423# vdd 0.003842f
C15912 net52 _453_/a_2665_112# 0.073881f
C15913 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_124_375# 0.007947f
C15914 _289_/a_36_472# _102_ 0.046918f
C15915 _430_/a_1308_423# _091_ 0.023198f
C15916 net75 _426_/a_796_472# 0.003146f
C15917 FILLER_0_11_64/a_124_375# cal_count\[3\] 0.002495f
C15918 _328_/a_36_113# _017_ 0.006485f
C15919 net57 _250_/a_36_68# 0.001141f
C15920 net4 FILLER_0_8_239/a_36_472# 0.008503f
C15921 output27/a_224_472# FILLER_0_9_290/a_124_375# 0.02894f
C15922 output14/a_224_472# net14 0.018674f
C15923 _116_ _055_ 0.72331f
C15924 _442_/a_448_472# FILLER_0_2_127/a_36_472# 0.008634f
C15925 net48 _122_ 0.110769f
C15926 FILLER_0_4_197/a_932_472# net22 0.0473f
C15927 _274_/a_2124_68# net4 0.00137f
C15928 net38 _054_ 0.640545f
C15929 net82 FILLER_0_3_221/a_36_472# 0.015923f
C15930 net48 FILLER_0_7_233/a_124_375# 0.013455f
C15931 net26 FILLER_0_18_37/a_932_472# 0.002613f
C15932 _098_ _438_/a_36_151# 0.009083f
C15933 _430_/a_448_472# net80 0.00896f
C15934 vss _022_ 0.067509f
C15935 FILLER_0_8_247/a_1468_375# calibrate 0.006404f
C15936 FILLER_0_12_220/a_572_375# _060_ 0.00145f
C15937 FILLER_0_16_89/a_1020_375# vdd 0.007416f
C15938 _443_/a_36_151# _371_/a_36_113# 0.001252f
C15939 FILLER_0_1_204/a_36_472# vdd 0.009339f
C15940 FILLER_0_1_204/a_124_375# vss 0.018397f
C15941 net65 FILLER_0_3_221/a_1020_375# 0.001641f
C15942 FILLER_0_3_172/a_3172_472# net22 0.010714f
C15943 valid fanout59/a_36_160# 0.029107f
C15944 _427_/a_2248_156# _043_ 0.001148f
C15945 _432_/a_36_151# mask\[3\] 0.002148f
C15946 _175_ FILLER_0_15_72/a_124_375# 0.009573f
C15947 net32 ctlp[2] 0.097138f
C15948 _256_/a_36_68# _056_ 0.008305f
C15949 net38 _278_/a_36_160# 0.010587f
C15950 net16 _043_ 0.049385f
C15951 _256_/a_1612_497# _055_ 0.001438f
C15952 _077_ cal_count\[3\] 0.176576f
C15953 _176_ _043_ 0.04106f
C15954 FILLER_0_17_142/a_124_375# vdd 0.020936f
C15955 ctln[6] net59 0.001267f
C15956 net20 net75 0.092951f
C15957 net18 result[3] 0.237732f
C15958 _120_ FILLER_0_8_156/a_572_375# 0.030218f
C15959 FILLER_0_11_78/a_572_375# _171_ 0.001028f
C15960 _308_/a_848_380# FILLER_0_9_105/a_36_472# 0.15783f
C15961 net38 vss 0.633752f
C15962 _106_ FILLER_0_17_218/a_572_375# 0.022684f
C15963 FILLER_0_16_107/a_124_375# FILLER_0_18_107/a_36_472# 0.001512f
C15964 FILLER_0_15_290/a_36_472# net79 0.04083f
C15965 _427_/a_1000_472# _095_ 0.021594f
C15966 _164_ _167_ 0.311625f
C15967 _077_ _059_ 0.020736f
C15968 _069_ _085_ 0.032519f
C15969 _027_ mask\[9\] 0.050723f
C15970 net38 _178_ 0.123812f
C15971 _118_ _055_ 0.042556f
C15972 _292_/a_36_160# net22 0.001864f
C15973 _053_ FILLER_0_6_47/a_1828_472# 0.006408f
C15974 net27 FILLER_0_9_290/a_36_472# 0.006729f
C15975 _321_/a_3126_472# _126_ 0.002939f
C15976 _321_/a_358_69# _069_ 0.001124f
C15977 FILLER_0_5_88/a_124_375# FILLER_0_6_90/a_36_472# 0.001543f
C15978 _308_/a_848_380# vdd 0.013895f
C15979 net42 output6/a_224_472# 0.009273f
C15980 net74 FILLER_0_13_142/a_484_472# 0.001771f
C15981 FILLER_0_5_109/a_572_375# vdd 0.024724f
C15982 _413_/a_1204_472# _002_ 0.003057f
C15983 net75 FILLER_0_6_231/a_572_375# 0.002577f
C15984 _428_/a_1000_472# _017_ 0.012268f
C15985 FILLER_0_2_171/a_124_375# vss 0.049142f
C15986 FILLER_0_2_171/a_36_472# vdd 0.029996f
C15987 _236_/a_36_160# FILLER_0_8_2/a_36_472# 0.01395f
C15988 _290_/a_224_472# net18 0.00868f
C15989 _162_ _056_ 0.018616f
C15990 FILLER_0_19_125/a_36_472# _022_ 0.013011f
C15991 _158_ vss 0.007784f
C15992 net16 net68 0.275467f
C15993 FILLER_0_16_241/a_124_375# _198_/a_67_603# 0.002082f
C15994 _408_/a_2215_68# _186_ 0.001205f
C15995 _444_/a_448_472# net47 0.030563f
C15996 _016_ fanout73/a_36_113# 0.001731f
C15997 _016_ FILLER_0_12_136/a_572_375# 0.00332f
C15998 net2 net5 0.47659f
C15999 fanout50/a_36_160# vdd 0.009536f
C16000 _256_/a_36_68# _068_ 0.029112f
C16001 net63 _435_/a_448_472# 0.009878f
C16002 result[4] net18 0.048179f
C16003 FILLER_0_8_24/a_124_375# net47 0.025599f
C16004 _070_ _313_/a_67_603# 0.004265f
C16005 net58 FILLER_0_9_282/a_36_472# 0.062389f
C16006 FILLER_0_18_107/a_932_472# vdd 0.009633f
C16007 _115_ _134_ 0.051655f
C16008 _430_/a_2665_112# _091_ 0.016404f
C16009 _126_ _118_ 0.215385f
C16010 _434_/a_36_151# _146_ 0.003818f
C16011 _434_/a_1204_472# mask\[6\] 0.006692f
C16012 _110_ vdd 0.041979f
C16013 FILLER_0_7_146/a_36_472# _313_/a_67_603# 0.002287f
C16014 FILLER_0_7_104/a_932_472# vdd 0.020291f
C16015 _424_/a_36_151# vss 0.030774f
C16016 _424_/a_448_472# vdd 0.014219f
C16017 cal_count\[2\] _041_ 0.02197f
C16018 net66 vss 0.265973f
C16019 _074_ _161_ 0.191658f
C16020 result[2] _416_/a_36_151# 0.010509f
C16021 mask\[4\] FILLER_0_18_177/a_484_472# 0.016924f
C16022 net52 _168_ 0.726039f
C16023 ctln[7] ctln[6] 0.00499f
C16024 trim_val\[4\] _163_ 0.03439f
C16025 _067_ vss 0.20904f
C16026 net50 _441_/a_448_472# 0.074088f
C16027 FILLER_0_4_107/a_1468_375# _154_ 0.005202f
C16028 FILLER_0_4_107/a_572_375# _153_ 0.010165f
C16029 FILLER_0_7_72/a_2276_472# net14 0.004375f
C16030 _308_/a_692_472# trim_mask\[0\] 0.004377f
C16031 FILLER_0_12_28/a_36_472# net40 0.020589f
C16032 output40/a_224_472# trim[2] 0.025041f
C16033 FILLER_0_12_236/a_484_472# _060_ 0.002678f
C16034 _016_ net57 0.028276f
C16035 fanout60/a_36_160# vss 0.035381f
C16036 _161_ _076_ 0.042123f
C16037 net49 _168_ 0.031157f
C16038 net18 _417_/a_1308_423# 0.015651f
C16039 FILLER_0_4_197/a_932_472# vdd 0.003395f
C16040 _417_/a_448_472# result[3] 0.003109f
C16041 _207_/a_67_603# FILLER_0_22_128/a_3260_375# 0.00744f
C16042 ctln[4] FILLER_0_0_198/a_36_472# 0.02582f
C16043 _187_ vss 0.080956f
C16044 _259_/a_271_68# net4 0.003663f
C16045 _207_/a_67_603# net33 0.005153f
C16046 FILLER_0_21_28/a_1828_472# _423_/a_36_151# 0.059367f
C16047 _437_/a_2665_112# vdd 0.050182f
C16048 net69 FILLER_0_2_111/a_124_375# 0.010762f
C16049 net61 _422_/a_1308_423# 0.002171f
C16050 net60 _422_/a_36_151# 0.008119f
C16051 FILLER_0_3_172/a_3172_472# vdd 0.003804f
C16052 _129_ _076_ 0.043637f
C16053 FILLER_0_4_144/a_124_375# _370_/a_848_380# 0.005599f
C16054 net41 _181_ 0.043679f
C16055 _430_/a_36_151# net21 0.019114f
C16056 FILLER_0_7_104/a_1380_472# _125_ 0.001279f
C16057 output23/a_224_472# _210_/a_67_603# 0.021084f
C16058 fanout61/a_36_113# net79 0.001865f
C16059 net16 net67 0.038448f
C16060 FILLER_0_5_117/a_36_472# _119_ 0.002628f
C16061 FILLER_0_19_171/a_1380_472# _434_/a_36_151# 0.00271f
C16062 state\[1\] _060_ 0.003973f
C16063 FILLER_0_12_136/a_572_375# FILLER_0_13_142/a_36_472# 0.001684f
C16064 fanout72/a_36_113# net72 0.02315f
C16065 trimb[1] _452_/a_2449_156# 0.001681f
C16066 net35 _148_ 0.114816f
C16067 FILLER_0_19_142/a_124_375# FILLER_0_19_134/a_124_375# 0.003732f
C16068 _431_/a_796_472# net70 0.001754f
C16069 _012_ FILLER_0_23_44/a_1020_375# 0.002827f
C16070 valid net5 0.044555f
C16071 FILLER_0_4_213/a_36_472# net59 0.044235f
C16072 cal_count\[3\] FILLER_0_12_196/a_36_472# 0.079338f
C16073 output31/a_224_472# net30 0.149277f
C16074 net55 _451_/a_3129_107# 0.098091f
C16075 FILLER_0_3_54/a_36_472# vdd 0.00827f
C16076 _292_/a_36_160# vdd 0.01694f
C16077 vss rstn 0.149553f
C16078 _069_ _062_ 0.029863f
C16079 result[4] _417_/a_448_472# 0.003485f
C16080 net57 _395_/a_1044_488# 0.002526f
C16081 net44 clkc 0.184915f
C16082 _415_/a_2560_156# net58 0.002325f
C16083 _102_ net19 0.011979f
C16084 _411_/a_1000_472# net8 0.007241f
C16085 FILLER_0_14_91/a_124_375# _176_ 0.019567f
C16086 FILLER_0_22_177/a_572_375# _435_/a_36_151# 0.059049f
C16087 ctlp[1] FILLER_0_23_282/a_484_472# 0.007608f
C16088 FILLER_0_24_130/a_36_472# _050_ 0.008605f
C16089 ctln[4] FILLER_0_0_232/a_124_375# 0.002726f
C16090 result[9] _421_/a_1000_472# 0.012144f
C16091 FILLER_0_14_181/a_124_375# mask\[1\] 0.044784f
C16092 net57 FILLER_0_13_142/a_36_472# 0.011199f
C16093 vdd net14 2.23064f
C16094 _098_ FILLER_0_20_98/a_36_472# 0.0127f
C16095 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3172_472# 0.013276f
C16096 FILLER_0_21_125/a_124_375# vdd -0.010326f
C16097 ctln[4] net11 0.194506f
C16098 fanout55/a_36_160# vdd 0.016488f
C16099 _091_ net63 0.767908f
C16100 net54 FILLER_0_18_139/a_932_472# 0.003365f
C16101 _432_/a_796_472# _098_ 0.038458f
C16102 _053_ FILLER_0_6_177/a_124_375# 0.009352f
C16103 output42/a_224_472# _444_/a_36_151# 0.002701f
C16104 _287_/a_36_472# mask\[2\] 0.00492f
C16105 FILLER_0_18_107/a_572_375# net14 0.00258f
C16106 FILLER_0_16_57/a_572_375# FILLER_0_18_61/a_36_472# 0.001512f
C16107 _177_ FILLER_0_17_72/a_1468_375# 0.026469f
C16108 _245_/a_234_472# net6 0.001301f
C16109 _164_ vdd 0.711488f
C16110 FILLER_0_5_109/a_124_375# _365_/a_36_68# 0.004633f
C16111 FILLER_0_8_247/a_484_472# vss -0.001894f
C16112 FILLER_0_8_247/a_932_472# vdd 0.008645f
C16113 net71 _436_/a_448_472# 0.005274f
C16114 _116_ state\[1\] 0.693219f
C16115 net81 _100_ 0.24831f
C16116 FILLER_0_4_197/a_1020_375# net82 0.00123f
C16117 FILLER_0_5_128/a_36_472# net47 0.008459f
C16118 ctlp[4] _108_ 0.002002f
C16119 net55 FILLER_0_18_37/a_36_472# 0.006084f
C16120 _066_ vss 0.08113f
C16121 output15/a_224_472# trim_val\[3\] 0.042209f
C16122 _011_ vdd 0.182751f
C16123 net72 FILLER_0_17_56/a_124_375# 0.018942f
C16124 sample net59 0.001181f
C16125 net78 _421_/a_1308_423# 0.015694f
C16126 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_572_375# 0.026339f
C16127 net37 net59 0.03883f
C16128 _404_/a_36_472# vdd 0.034854f
C16129 output31/a_224_472# _417_/a_36_151# 0.07368f
C16130 FILLER_0_17_200/a_124_375# net21 0.048656f
C16131 _428_/a_36_151# vdd 0.131612f
C16132 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_484_472# 0.013276f
C16133 _003_ _122_ 0.033778f
C16134 _098_ _433_/a_36_151# 0.023263f
C16135 _091_ _069_ 0.741596f
C16136 net38 _450_/a_1040_527# 0.027925f
C16137 _011_ _422_/a_796_472# 0.009261f
C16138 FILLER_0_7_72/a_2364_375# vdd 0.018287f
C16139 net25 vss 0.528437f
C16140 result[6] ctlp[1] 0.677825f
C16141 FILLER_0_12_136/a_1468_375# state\[2\] 0.035275f
C16142 net23 vss 1.922425f
C16143 _131_ _152_ 0.002949f
C16144 net1 _265_/a_224_472# 0.005504f
C16145 FILLER_0_4_49/a_484_472# _160_ 0.001336f
C16146 trimb[4] net55 0.01379f
C16147 FILLER_0_14_50/a_36_472# _181_ 0.001514f
C16148 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_572_375# 0.086635f
C16149 _177_ _040_ 0.061289f
C16150 _074_ _056_ 0.002397f
C16151 _341_/a_665_69# net23 0.001508f
C16152 FILLER_0_10_78/a_124_375# cal_count\[3\] 0.012197f
C16153 _149_ FILLER_0_20_107/a_124_375# 0.001244f
C16154 _315_/a_36_68# _120_ 0.00572f
C16155 net80 _434_/a_448_472# 0.113898f
C16156 FILLER_0_16_57/a_484_472# vdd 0.005894f
C16157 FILLER_0_16_57/a_36_472# vss 0.003789f
C16158 net35 _436_/a_2665_112# 0.012468f
C16159 FILLER_0_14_81/a_124_375# _176_ 0.001549f
C16160 _132_ FILLER_0_14_107/a_572_375# 0.007439f
C16161 _305_/a_36_159# calibrate 0.003505f
C16162 _112_ _316_/a_848_380# 0.022235f
C16163 FILLER_0_15_150/a_124_375# FILLER_0_15_142/a_572_375# 0.012001f
C16164 fanout68/a_36_113# net69 0.046009f
C16165 FILLER_0_5_117/a_124_375# _360_/a_36_160# 0.004736f
C16166 FILLER_0_11_109/a_124_375# FILLER_0_9_105/a_484_472# 0.0027f
C16167 _328_/a_36_113# cal_count\[3\] 0.006392f
C16168 net15 _449_/a_1308_423# 0.015651f
C16169 _354_/a_49_472# net71 0.010421f
C16170 _430_/a_36_151# net80 0.082603f
C16171 _056_ _076_ 0.938912f
C16172 _061_ _070_ 0.02813f
C16173 FILLER_0_15_212/a_932_472# vdd 0.001767f
C16174 FILLER_0_15_212/a_1468_375# mask\[1\] 0.045287f
C16175 FILLER_0_10_214/a_36_472# _090_ 0.011963f
C16176 net72 _452_/a_448_472# 0.001296f
C16177 FILLER_0_11_109/a_124_375# vss 0.006764f
C16178 FILLER_0_11_109/a_36_472# vdd 0.109453f
C16179 _359_/a_244_68# _059_ 0.002986f
C16180 _122_ net37 3.870625f
C16181 _072_ _374_/a_244_472# 0.001816f
C16182 _111_ _438_/a_36_151# 0.003619f
C16183 net32 mask\[7\] 0.01969f
C16184 FILLER_0_20_177/a_1468_375# _434_/a_2248_156# 0.001221f
C16185 FILLER_0_5_128/a_36_472# net74 0.01163f
C16186 FILLER_0_5_172/a_36_472# vss 0.003406f
C16187 FILLER_0_9_270/a_484_472# FILLER_0_9_282/a_36_472# 0.002296f
C16188 net54 _436_/a_36_151# 0.004179f
C16189 _427_/a_2665_112# _225_/a_36_160# 0.001394f
C16190 _065_ _447_/a_1000_472# 0.03162f
C16191 sample net64 0.209777f
C16192 FILLER_0_13_206/a_36_472# net21 0.00171f
C16193 net62 FILLER_0_15_282/a_484_472# 0.009524f
C16194 _434_/a_1000_472# vdd 0.032431f
C16195 _431_/a_2665_112# FILLER_0_16_154/a_36_472# 0.007491f
C16196 trimb[4] net17 0.004628f
C16197 _067_ _450_/a_1040_527# 0.007414f
C16198 _429_/a_36_151# _138_ 0.002064f
C16199 net81 FILLER_0_8_263/a_124_375# 0.026195f
C16200 _431_/a_2560_156# _136_ 0.013111f
C16201 _074_ _068_ 0.011897f
C16202 _169_ net37 0.03934f
C16203 net81 FILLER_0_14_235/a_124_375# 0.01391f
C16204 _174_ _183_ 0.008231f
C16205 _008_ net30 1.112351f
C16206 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_36_472# 0.016748f
C16207 _432_/a_1000_472# _093_ 0.007509f
C16208 _446_/a_2248_156# _160_ 0.002464f
C16209 FILLER_0_4_197/a_484_472# net22 0.007955f
C16210 FILLER_0_11_101/a_484_472# _070_ 0.017841f
C16211 net38 _095_ 0.032393f
C16212 _080_ FILLER_0_3_221/a_932_472# 0.003217f
C16213 output8/a_224_472# FILLER_0_3_221/a_36_472# 0.001699f
C16214 vdd FILLER_0_8_156/a_124_375# 0.005213f
C16215 _076_ _068_ 0.35956f
C16216 mask\[4\] _145_ 0.340415f
C16217 _013_ _131_ 0.001178f
C16218 result[9] net18 0.019413f
C16219 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001723f
C16220 net75 _265_/a_244_68# 0.046186f
C16221 net35 FILLER_0_22_128/a_1468_375# 0.015932f
C16222 _428_/a_36_151# _135_ 0.030608f
C16223 _072_ _070_ 2.141346f
C16224 net35 _207_/a_67_603# 0.005045f
C16225 _207_/a_255_603# mask\[6\] 0.003114f
C16226 _088_ _080_ 0.003418f
C16227 _414_/a_36_151# _087_ 0.010359f
C16228 net68 FILLER_0_6_47/a_124_375# 0.002491f
C16229 _064_ _445_/a_1204_472# 0.007445f
C16230 ctlp[7] vdd 0.481613f
C16231 output33/a_224_472# ctlp[2] 0.00175f
C16232 FILLER_0_4_177/a_572_375# net22 0.006125f
C16233 _089_ cal_itt\[3\] 0.049851f
C16234 net15 _439_/a_36_151# 0.068183f
C16235 _406_/a_36_159# cal_count\[2\] 0.028829f
C16236 FILLER_0_4_107/a_932_472# FILLER_0_2_111/a_572_375# 0.001512f
C16237 output42/a_224_472# _054_ 0.013225f
C16238 _397_/a_244_68# net55 0.001173f
C16239 _119_ _163_ 0.009297f
C16240 _086_ calibrate 0.041755f
C16241 _217_/a_36_160# vdd 0.092586f
C16242 result[7] ctlp[1] 0.07619f
C16243 net81 _060_ 0.019654f
C16244 _174_ FILLER_0_15_59/a_572_375# 0.007123f
C16245 net60 _419_/a_36_151# 0.016173f
C16246 net61 _419_/a_1308_423# 0.00793f
C16247 net80 FILLER_0_22_177/a_932_472# 0.002472f
C16248 FILLER_0_17_104/a_572_375# vdd 0.03661f
C16249 _013_ FILLER_0_18_37/a_572_375# 0.003828f
C16250 FILLER_0_5_88/a_36_472# net47 0.003953f
C16251 FILLER_0_3_172/a_36_472# FILLER_0_5_172/a_124_375# 0.0027f
C16252 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_124_375# 0.026339f
C16253 _161_ _090_ 0.207838f
C16254 _148_ vdd 0.01565f
C16255 ctlp[1] FILLER_0_21_286/a_124_375# 0.025059f
C16256 _147_ _435_/a_36_151# 0.003096f
C16257 cal_count\[3\] _039_ 0.004827f
C16258 _004_ vdd 0.448886f
C16259 _004_ _192_/a_67_603# 0.020219f
C16260 _440_/a_448_472# _029_ 0.043511f
C16261 _372_/a_2590_472# vss 0.00106f
C16262 net69 _170_ 0.006468f
C16263 FILLER_0_8_127/a_36_472# _125_ 0.003088f
C16264 FILLER_0_12_220/a_1380_472# vss 0.006172f
C16265 FILLER_0_16_107/a_484_472# _131_ 0.008223f
C16266 _058_ FILLER_0_8_156/a_484_472# 0.013955f
C16267 output42/a_224_472# vss 0.00418f
C16268 FILLER_0_11_109/a_36_472# _135_ 0.001891f
C16269 FILLER_0_17_72/a_3260_375# _451_/a_1040_527# 0.001117f
C16270 FILLER_0_4_123/a_124_375# _152_ 0.039668f
C16271 _086_ _414_/a_36_151# 0.002687f
C16272 _412_/a_2665_112# net1 0.063655f
C16273 _095_ _067_ 0.00784f
C16274 _060_ _223_/a_36_160# 0.002922f
C16275 net39 _445_/a_1000_472# 0.007782f
C16276 FILLER_0_5_72/a_36_472# trim_mask\[1\] 0.015775f
C16277 FILLER_0_5_72/a_1380_472# _029_ 0.007385f
C16278 _431_/a_2665_112# FILLER_0_18_139/a_1380_472# 0.001008f
C16279 FILLER_0_10_78/a_1380_472# _120_ 0.003228f
C16280 _136_ _038_ 0.061274f
C16281 _036_ net66 0.04474f
C16282 net68 _030_ 0.007737f
C16283 FILLER_0_5_206/a_124_375# net37 0.005485f
C16284 FILLER_0_20_193/a_124_375# FILLER_0_20_177/a_1468_375# 0.012222f
C16285 _008_ _417_/a_36_151# 0.001136f
C16286 _057_ _128_ 0.036548f
C16287 _452_/a_1040_527# net40 0.007832f
C16288 mask\[2\] FILLER_0_16_154/a_932_472# 0.021665f
C16289 net34 _299_/a_36_472# 0.003396f
C16290 FILLER_0_9_28/a_124_375# net42 0.007403f
C16291 mask\[5\] _137_ 0.002972f
C16292 FILLER_0_6_37/a_36_472# _160_ 0.008686f
C16293 _065_ output15/a_224_472# 0.037721f
C16294 _187_ _095_ 0.00765f
C16295 _439_/a_36_151# net51 0.00711f
C16296 _057_ _311_/a_692_473# 0.002083f
C16297 FILLER_0_22_86/a_484_472# _098_ 0.003294f
C16298 FILLER_0_17_72/a_3260_375# _131_ 0.004986f
C16299 trim_mask\[1\] _166_ 0.124855f
C16300 _415_/a_448_472# FILLER_0_11_282/a_124_375# 0.008952f
C16301 net16 _380_/a_224_472# 0.008718f
C16302 net67 FILLER_0_6_47/a_124_375# 0.005516f
C16303 FILLER_0_7_72/a_2276_472# _439_/a_2665_112# 0.001167f
C16304 net55 FILLER_0_13_72/a_484_472# 0.004375f
C16305 vss FILLER_0_19_134/a_124_375# 0.021427f
C16306 vdd FILLER_0_19_134/a_36_472# 0.092128f
C16307 _153_ vdd 0.672318f
C16308 fanout73/a_36_113# vss 0.01873f
C16309 _070_ _319_/a_234_472# 0.004015f
C16310 _449_/a_2560_156# vss 0.002544f
C16311 FILLER_0_12_136/a_1020_375# vdd 0.017472f
C16312 FILLER_0_12_136/a_572_375# vss 0.006091f
C16313 FILLER_0_15_116/a_124_375# net70 0.02416f
C16314 FILLER_0_23_274/a_124_375# vdd 0.014998f
C16315 _431_/a_2560_156# net53 0.002265f
C16316 _053_ _365_/a_36_68# 0.001572f
C16317 FILLER_0_7_72/a_1020_375# net52 0.00799f
C16318 result[6] _421_/a_2560_156# 0.006943f
C16319 net26 _423_/a_796_472# 0.001077f
C16320 _030_ _156_ 0.153053f
C16321 net64 FILLER_0_9_282/a_572_375# 0.002322f
C16322 _092_ FILLER_0_18_209/a_484_472# 0.006303f
C16323 result[7] FILLER_0_24_274/a_124_375# 0.006125f
C16324 _001_ _082_ 0.46787f
C16325 mask\[0\] FILLER_0_15_212/a_1468_375# 0.001182f
C16326 FILLER_0_3_142/a_36_472# vss 0.012379f
C16327 net82 _001_ 0.044461f
C16328 FILLER_0_8_138/a_124_375# _058_ 0.009863f
C16329 FILLER_0_4_197/a_484_472# vdd 0.002749f
C16330 _411_/a_2665_112# net58 0.018133f
C16331 FILLER_0_5_54/a_572_375# vdd 0.004086f
C16332 FILLER_0_17_72/a_1020_375# net36 0.001777f
C16333 _412_/a_1000_472# net58 0.030238f
C16334 output34/a_224_472# net32 0.027498f
C16335 _076_ _152_ 0.063574f
C16336 _068_ _081_ 0.006663f
C16337 _451_/a_2225_156# _040_ 0.015815f
C16338 _071_ net23 0.027895f
C16339 mask\[9\] FILLER_0_20_87/a_124_375# 0.004793f
C16340 mask\[5\] _049_ 0.008296f
C16341 _096_ _090_ 0.026104f
C16342 _402_/a_1948_68# vdd 0.001429f
C16343 output9/a_224_472# net76 0.002042f
C16344 mask\[3\] net21 0.100738f
C16345 _126_ FILLER_0_14_181/a_36_472# 0.008653f
C16346 net41 _446_/a_2248_156# 0.016492f
C16347 FILLER_0_18_177/a_124_375# vdd 0.033102f
C16348 _020_ FILLER_0_18_107/a_2276_472# 0.004069f
C16349 FILLER_0_4_177/a_572_375# vdd 0.001622f
C16350 FILLER_0_4_177/a_124_375# vss 0.002462f
C16351 _449_/a_448_472# _067_ 0.0432f
C16352 _036_ FILLER_0_3_54/a_124_375# 0.010221f
C16353 net57 vss 0.818311f
C16354 net4 FILLER_0_3_212/a_124_375# 0.001739f
C16355 _127_ _121_ 0.023125f
C16356 FILLER_0_12_20/a_124_375# vdd 0.017452f
C16357 FILLER_0_19_47/a_484_472# _013_ 0.009677f
C16358 net1 _084_ 0.008356f
C16359 net31 _092_ 0.04309f
C16360 FILLER_0_19_155/a_484_472# vss 0.004002f
C16361 FILLER_0_18_2/a_572_375# _452_/a_3129_107# 0.001073f
C16362 net66 output41/a_224_472# 0.015427f
C16363 _425_/a_448_472# _014_ 0.013561f
C16364 _256_/a_1164_497# net4 0.004729f
C16365 _214_/a_36_160# _098_ 0.001496f
C16366 mask\[2\] FILLER_0_15_205/a_36_472# 0.001204f
C16367 _142_ vdd 0.090938f
C16368 ctln[2] FILLER_0_1_266/a_484_472# 0.019076f
C16369 FILLER_0_24_63/a_124_375# ctlp[9] 0.002726f
C16370 FILLER_0_16_57/a_124_375# _183_ 0.005825f
C16371 net16 net26 0.273031f
C16372 FILLER_0_3_221/a_932_472# vss 0.002881f
C16373 FILLER_0_3_221/a_1380_472# vdd 0.003819f
C16374 FILLER_0_4_99/a_124_375# net47 0.001409f
C16375 _436_/a_2248_156# vss 0.002799f
C16376 _436_/a_2665_112# vdd 0.007946f
C16377 net73 FILLER_0_18_107/a_1916_375# 0.014643f
C16378 mask\[7\] FILLER_0_22_128/a_124_375# 0.01319f
C16379 _378_/a_224_472# vdd 0.002263f
C16380 _273_/a_36_68# FILLER_0_10_214/a_124_375# 0.003707f
C16381 net74 FILLER_0_13_100/a_124_375# 0.005049f
C16382 FILLER_0_9_28/a_1020_375# net50 0.001512f
C16383 state\[1\] _228_/a_36_68# 0.024977f
C16384 FILLER_0_14_123/a_124_375# FILLER_0_14_107/a_1468_375# 0.012001f
C16385 _439_/a_2248_156# vss 0.003954f
C16386 _439_/a_2665_112# vdd 0.015979f
C16387 calibrate _313_/a_67_603# 0.021436f
C16388 FILLER_0_22_128/a_932_472# _433_/a_36_151# 0.002841f
C16389 net41 _423_/a_36_151# 0.001134f
C16390 _289_/a_36_472# _198_/a_67_603# 0.027695f
C16391 _002_ FILLER_0_3_172/a_1916_375# 0.047331f
C16392 _088_ vss 0.326434f
C16393 _428_/a_448_472# _043_ 0.063478f
C16394 FILLER_0_21_28/a_1380_472# _424_/a_36_151# 0.001723f
C16395 output29/a_224_472# result[2] 0.058798f
C16396 net63 FILLER_0_15_212/a_932_472# 0.002269f
C16397 _077_ net52 0.047585f
C16398 FILLER_0_14_91/a_36_472# _067_ 0.004194f
C16399 net79 FILLER_0_13_290/a_124_375# 0.043673f
C16400 _115_ _322_/a_124_24# 0.019655f
C16401 net62 FILLER_0_13_290/a_36_472# 0.003157f
C16402 fanout69/a_36_113# _032_ 0.003681f
C16403 _176_ _394_/a_728_93# 0.002001f
C16404 net5 cal_itt\[1\] 0.057623f
C16405 FILLER_0_12_136/a_932_472# cal_count\[3\] 0.007247f
C16406 net72 cal_count\[3\] 0.059493f
C16407 net58 _425_/a_2248_156# 0.051603f
C16408 net44 FILLER_0_12_2/a_484_472# 0.046864f
C16409 _443_/a_1308_423# _170_ 0.043472f
C16410 FILLER_0_10_28/a_124_375# net40 0.047331f
C16411 _056_ _090_ 0.177189f
C16412 _003_ FILLER_0_5_181/a_36_472# 0.003545f
C16413 state\[2\] FILLER_0_13_142/a_124_375# 0.010494f
C16414 net63 _434_/a_1000_472# 0.002404f
C16415 _091_ _140_ 0.006511f
C16416 net53 FILLER_0_13_142/a_1020_375# 0.001597f
C16417 _430_/a_796_472# _019_ 0.006511f
C16418 ctln[5] _037_ 0.19244f
C16419 ctlp[8] vss 0.107975f
C16420 _095_ net23 0.053365f
C16421 _308_/a_124_24# _439_/a_2248_156# 0.01963f
C16422 FILLER_0_9_223/a_36_472# _055_ 0.014713f
C16423 _093_ net30 0.001859f
C16424 net70 _040_ 0.018254f
C16425 trim_mask\[3\] _156_ 0.002638f
C16426 net8 net59 0.062623f
C16427 _448_/a_2665_112# _387_/a_36_113# 0.010064f
C16428 _448_/a_796_472# _037_ 0.009263f
C16429 vdd output40/a_224_472# 0.079607f
C16430 net7 ctln[9] 0.005103f
C16431 FILLER_0_22_128/a_1020_375# vss 0.003747f
C16432 FILLER_0_22_128/a_1468_375# vdd 0.016807f
C16433 _233_/a_36_160# _063_ 0.002771f
C16434 _255_/a_224_552# _058_ 0.06267f
C16435 _408_/a_728_93# _181_ 0.018292f
C16436 _207_/a_67_603# vdd 0.034688f
C16437 _086_ FILLER_0_11_142/a_124_375# 0.009046f
C16438 _161_ _163_ 0.024512f
C16439 _028_ _439_/a_36_151# 0.009268f
C16440 FILLER_0_20_15/a_1468_375# net40 0.030032f
C16441 _081_ _152_ 0.172002f
C16442 _315_/a_244_497# vss 0.008724f
C16443 _077_ FILLER_0_8_239/a_124_375# 0.001772f
C16444 _275_/a_224_472# net63 0.002538f
C16445 cal_itt\[0\] vss 0.11965f
C16446 _088_ FILLER_0_3_172/a_3260_375# 0.002239f
C16447 _086_ FILLER_0_7_104/a_124_375# 0.001629f
C16448 net31 net61 0.053131f
C16449 net15 _160_ 0.046497f
C16450 FILLER_0_16_107/a_36_472# _132_ 0.001538f
C16451 FILLER_0_15_142/a_572_375# net53 0.021481f
C16452 FILLER_0_5_181/a_36_472# net37 0.010376f
C16453 FILLER_0_15_282/a_124_375# vdd 0.011964f
C16454 FILLER_0_7_72/a_124_375# vss 0.044754f
C16455 _431_/a_448_472# _131_ 0.006194f
C16456 _032_ _371_/a_36_113# 0.030245f
C16457 FILLER_0_17_200/a_572_375# _430_/a_36_151# 0.059049f
C16458 FILLER_0_16_37/a_124_375# FILLER_0_18_37/a_36_472# 0.001512f
C16459 fanout49/a_36_160# trim_mask\[1\] 0.00358f
C16460 net57 FILLER_0_2_165/a_36_472# 0.001562f
C16461 FILLER_0_7_59/a_124_375# trim_mask\[1\] 0.001548f
C16462 FILLER_0_8_107/a_36_472# _219_/a_36_160# 0.002767f
C16463 _053_ FILLER_0_7_72/a_3172_472# 0.032946f
C16464 FILLER_0_14_91/a_572_375# net14 0.005527f
C16465 _127_ _321_/a_170_472# 0.023836f
C16466 net32 _419_/a_2248_156# 0.034827f
C16467 mask\[3\] net80 0.02972f
C16468 _087_ FILLER_0_5_181/a_124_375# 0.068f
C16469 mask\[9\] _098_ 0.256513f
C16470 _141_ FILLER_0_19_171/a_36_472# 0.001292f
C16471 FILLER_0_6_47/a_2724_472# vdd 0.002467f
C16472 FILLER_0_6_47/a_2276_472# vss 0.004086f
C16473 FILLER_0_14_123/a_124_375# vdd 0.034436f
C16474 _126_ net74 1.001749f
C16475 net34 _104_ 0.293336f
C16476 _105_ _422_/a_36_151# 0.030571f
C16477 FILLER_0_20_31/a_36_472# net40 0.045181f
C16478 _275_/a_224_472# _069_ 0.004466f
C16479 FILLER_0_10_107/a_124_375# FILLER_0_10_94/a_572_375# 0.003228f
C16480 ctln[2] net2 0.004284f
C16481 net58 FILLER_0_8_263/a_36_472# 0.059769f
C16482 _063_ net49 0.002854f
C16483 fanout52/a_36_160# _386_/a_124_24# 0.004695f
C16484 net34 vss 0.481379f
C16485 _143_ vdd 0.074199f
C16486 mask\[0\] FILLER_0_13_206/a_36_472# 0.012766f
C16487 FILLER_0_12_2/a_36_472# output6/a_224_472# 0.00108f
C16488 _322_/a_1084_68# _118_ 0.002515f
C16489 net53 state\[2\] 0.001982f
C16490 FILLER_0_13_212/a_932_472# vss 0.022933f
C16491 output39/a_224_472# _034_ 0.002236f
C16492 _066_ _385_/a_36_68# 0.001405f
C16493 _346_/a_49_472# net23 0.022558f
C16494 _443_/a_448_472# net69 0.068491f
C16495 net55 _423_/a_448_472# 0.00206f
C16496 net26 FILLER_0_21_28/a_2364_375# 0.003691f
C16497 FILLER_0_15_142/a_484_472# FILLER_0_15_150/a_36_472# 0.013277f
C16498 FILLER_0_12_136/a_1380_472# _114_ 0.003953f
C16499 net20 _102_ 0.081029f
C16500 ctlp[1] _420_/a_1000_472# 0.001106f
C16501 FILLER_0_3_204/a_36_472# net65 0.001777f
C16502 _161_ _117_ 0.25528f
C16503 _086_ FILLER_0_5_181/a_124_375# 0.006872f
C16504 _276_/a_36_160# FILLER_0_17_218/a_36_472# 0.035111f
C16505 _431_/a_448_472# net56 0.001464f
C16506 _446_/a_2665_112# net17 0.00149f
C16507 _072_ _395_/a_244_68# 0.001406f
C16508 _446_/a_2665_112# trim_val\[1\] 0.001275f
C16509 _023_ _146_ 0.006636f
C16510 vdd FILLER_0_5_148/a_36_472# 0.001227f
C16511 vss FILLER_0_5_148/a_572_375# 0.042687f
C16512 net52 net50 0.702793f
C16513 output27/a_224_472# FILLER_0_9_270/a_572_375# 0.00135f
C16514 _037_ net59 0.799647f
C16515 FILLER_0_4_177/a_36_472# net76 0.003007f
C16516 output44/a_224_472# _452_/a_448_472# 0.004683f
C16517 net55 FILLER_0_17_72/a_484_472# 0.019636f
C16518 net57 _071_ 0.12089f
C16519 _139_ mask\[2\] 0.035793f
C16520 FILLER_0_16_89/a_572_375# _451_/a_448_472# 0.001597f
C16521 FILLER_0_2_111/a_932_472# vdd 0.003808f
C16522 FILLER_0_2_111/a_124_375# _369_/a_36_68# 0.001176f
C16523 FILLER_0_2_111/a_484_472# vss -0.001894f
C16524 _028_ FILLER_0_6_47/a_3260_375# 0.013006f
C16525 net41 _444_/a_2248_156# 0.028267f
C16526 net15 _394_/a_718_524# 0.027444f
C16527 net50 net49 0.238748f
C16528 net20 FILLER_0_8_239/a_124_375# 0.004302f
C16529 ctln[1] FILLER_0_0_232/a_36_472# 0.005158f
C16530 _440_/a_1204_472# vss 0.007007f
C16531 _440_/a_2248_156# vdd -0.003421f
C16532 FILLER_0_14_99/a_36_472# FILLER_0_13_100/a_36_472# 0.026657f
C16533 ctln[4] net10 0.1323f
C16534 trim_val\[4\] net37 0.003661f
C16535 net34 _107_ 0.017589f
C16536 output46/a_224_472# net38 0.003296f
C16537 FILLER_0_7_72/a_1468_375# vss 0.003253f
C16538 FILLER_0_18_2/a_1380_472# vss -0.001894f
C16539 FILLER_0_24_130/a_124_375# ctlp[6] 0.021926f
C16540 net18 _418_/a_1000_472# 0.050485f
C16541 FILLER_0_24_63/a_36_472# vdd 0.055524f
C16542 _340_/a_36_160# vss 0.029871f
C16543 _008_ _046_ 0.067769f
C16544 net63 FILLER_0_18_177/a_124_375# 0.001937f
C16545 net62 FILLER_0_15_235/a_124_375# 0.001315f
C16546 net57 FILLER_0_16_154/a_1020_375# 0.001902f
C16547 net82 _443_/a_1000_472# 0.008161f
C16548 FILLER_0_21_28/a_1828_472# _012_ 0.021162f
C16549 net70 FILLER_0_14_107/a_484_472# 0.010987f
C16550 net44 FILLER_0_20_2/a_484_472# 0.039736f
C16551 FILLER_0_12_136/a_124_375# _126_ 0.013041f
C16552 _050_ FILLER_0_22_128/a_932_472# 0.001098f
C16553 FILLER_0_1_266/a_124_375# net8 0.012703f
C16554 net27 FILLER_0_9_270/a_36_472# 0.041681f
C16555 FILLER_0_0_96/a_36_472# vdd 0.047982f
C16556 FILLER_0_0_96/a_124_375# vss 0.008342f
C16557 _306_/a_36_68# cal_count\[3\] 0.007663f
C16558 fanout72/a_36_113# vdd -0.002193f
C16559 net41 FILLER_0_21_28/a_1020_375# 0.010649f
C16560 ctlp[1] _419_/a_1204_472# 0.007338f
C16561 _432_/a_2248_156# _137_ 0.001775f
C16562 mask\[8\] _352_/a_49_472# 0.002573f
C16563 net73 FILLER_0_19_111/a_124_375# 0.005778f
C16564 fanout73/a_36_113# _095_ 0.003989f
C16565 net52 FILLER_0_5_72/a_572_375# 0.024148f
C16566 _057_ _114_ 0.30288f
C16567 FILLER_0_21_142/a_572_375# _098_ 0.006558f
C16568 FILLER_0_7_72/a_3260_375# vss 0.053035f
C16569 _061_ net21 0.049282f
C16570 FILLER_0_4_177/a_36_472# FILLER_0_2_177/a_124_375# 0.001512f
C16571 output34/a_224_472# mask\[3\] 0.002385f
C16572 mask\[5\] FILLER_0_19_171/a_484_472# 0.007647f
C16573 FILLER_0_5_72/a_572_375# net49 0.001158f
C16574 _311_/a_66_473# net21 0.02018f
C16575 _412_/a_2248_156# net1 0.044934f
C16576 _114_ _250_/a_36_68# 0.017773f
C16577 FILLER_0_15_2/a_572_375# vdd 0.017581f
C16578 FILLER_0_15_2/a_124_375# vss 0.002713f
C16579 output34/a_224_472# _421_/a_2665_112# 0.00151f
C16580 _004_ net28 0.082388f
C16581 _079_ FILLER_0_5_198/a_484_472# 0.008167f
C16582 FILLER_0_19_28/a_36_472# net40 0.020968f
C16583 trim_val\[1\] trim_mask\[1\] 0.519723f
C16584 _058_ _120_ 0.008566f
C16585 net68 FILLER_0_5_54/a_1020_375# 0.00648f
C16586 net15 FILLER_0_7_59/a_572_375# 0.033245f
C16587 FILLER_0_10_78/a_124_375# net52 0.008557f
C16588 _248_/a_36_68# net22 0.002193f
C16589 net57 _095_ 0.07431f
C16590 net66 _166_ 0.011066f
C16591 FILLER_0_21_125/a_124_375# _140_ 0.031374f
C16592 net16 _033_ 0.042852f
C16593 _072_ calibrate 0.539702f
C16594 fanout66/a_36_113# trim_mask\[2\] 0.015961f
C16595 net36 FILLER_0_15_235/a_36_472# 0.00664f
C16596 FILLER_0_6_177/a_36_472# vdd 0.109918f
C16597 FILLER_0_6_177/a_572_375# vss 0.008666f
C16598 _028_ FILLER_0_5_72/a_484_472# 0.003042f
C16599 _376_/a_36_160# vdd -0.006711f
C16600 FILLER_0_9_223/a_124_375# vdd 0.006153f
C16601 net1 net4 0.03357f
C16602 _141_ vss 0.308762f
C16603 _147_ net23 0.011375f
C16604 _341_/a_49_472# vdd 0.026636f
C16605 _077_ FILLER_0_8_156/a_36_472# 0.00563f
C16606 net41 net39 0.003649f
C16607 net81 net2 1.204674f
C16608 _057_ _176_ 0.001304f
C16609 _348_/a_49_472# vss 0.002301f
C16610 _417_/a_796_472# _006_ 0.014427f
C16611 result[5] result[6] 0.065361f
C16612 FILLER_0_7_104/a_1468_375# _131_ 0.029718f
C16613 FILLER_0_7_146/a_124_375# _062_ 0.028312f
C16614 _301_/a_36_472# vss 0.003975f
C16615 _438_/a_448_472# _437_/a_36_151# 0.00198f
C16616 net41 net51 0.031531f
C16617 ctln[1] FILLER_0_1_266/a_36_472# 0.002068f
C16618 net36 vss 1.788802f
C16619 _077_ _229_/a_224_472# 0.001293f
C16620 _068_ _163_ 0.04926f
C16621 _072_ net21 0.062333f
C16622 _335_/a_49_472# _043_ 0.00367f
C16623 ctlp[3] ctlp[2] 0.006764f
C16624 FILLER_0_18_37/a_1380_472# vdd 0.004422f
C16625 _141_ _341_/a_665_69# 0.001064f
C16626 _317_/a_36_113# _123_ 0.037893f
C16627 _014_ calibrate 0.403103f
C16628 _091_ FILLER_0_13_228/a_36_472# 0.001826f
C16629 _144_ _436_/a_36_151# 0.029716f
C16630 _429_/a_2248_156# vdd -0.006752f
C16631 _429_/a_1204_472# vss 0.002428f
C16632 _367_/a_244_472# _154_ 0.001775f
C16633 FILLER_0_17_56/a_124_375# vdd 0.008529f
C16634 net79 net19 0.03862f
C16635 _077_ FILLER_0_10_78/a_484_472# 0.002486f
C16636 FILLER_0_12_220/a_1380_472# FILLER_0_12_236/a_36_472# 0.013277f
C16637 FILLER_0_13_212/a_36_472# mask\[0\] 0.001366f
C16638 _273_/a_36_68# _076_ 0.001503f
C16639 _414_/a_36_151# _072_ 0.033026f
C16640 net16 _180_ 0.00101f
C16641 FILLER_0_19_195/a_124_375# net21 0.039225f
C16642 _316_/a_124_24# vdd 0.033047f
C16643 net79 _416_/a_796_472# 0.01137f
C16644 _176_ _180_ 0.030701f
C16645 net18 _044_ 0.174456f
C16646 net62 _416_/a_1000_472# 0.002399f
C16647 FILLER_0_9_28/a_572_375# vdd 0.023246f
C16648 _193_/a_36_160# vss 0.035228f
C16649 output31/a_224_472# _006_ 0.090006f
C16650 ctlp[2] net78 0.369805f
C16651 _056_ _117_ 0.065147f
C16652 _098_ _022_ 0.013131f
C16653 _017_ vdd 0.26981f
C16654 ctln[5] _448_/a_2248_156# 0.004396f
C16655 net26 _424_/a_1308_423# 0.001179f
C16656 _053_ _062_ 0.185944f
C16657 _120_ _389_/a_36_148# 0.022887f
C16658 _091_ _274_/a_2960_68# 0.001338f
C16659 _038_ _389_/a_36_148# 0.003749f
C16660 _430_/a_1000_472# net22 0.032221f
C16661 FILLER_0_10_247/a_36_472# vss 0.002828f
C16662 cal vss 0.424638f
C16663 _431_/a_2665_112# net56 0.048214f
C16664 output31/a_224_472# _103_ 0.006731f
C16665 FILLER_0_18_2/a_932_472# net38 0.020589f
C16666 trim[4] _221_/a_36_160# 0.002685f
C16667 FILLER_0_15_235/a_36_472# FILLER_0_15_228/a_36_472# 0.002765f
C16668 FILLER_0_9_105/a_572_375# FILLER_0_10_107/a_484_472# 0.001543f
C16669 _090_ _113_ 0.263235f
C16670 FILLER_0_21_206/a_36_472# net33 0.001447f
C16671 fanout51/a_36_113# FILLER_0_11_78/a_124_375# 0.005683f
C16672 _451_/a_36_151# net14 0.037503f
C16673 FILLER_0_18_2/a_36_472# vdd 0.104532f
C16674 _285_/a_36_472# mask\[1\] 0.036335f
C16675 FILLER_0_5_72/a_1468_375# _164_ 0.040819f
C16676 FILLER_0_10_107/a_36_472# vdd 0.117291f
C16677 FILLER_0_10_107/a_572_375# vss 0.017711f
C16678 FILLER_0_15_228/a_36_472# vss 0.006585f
C16679 FILLER_0_3_204/a_124_375# vss 0.017795f
C16680 FILLER_0_11_282/a_36_472# _416_/a_448_472# 0.011962f
C16681 _452_/a_36_151# vss 0.02741f
C16682 _452_/a_448_472# vdd 0.019824f
C16683 trim_mask\[0\] FILLER_0_10_94/a_484_472# 0.015575f
C16684 net81 valid 0.11798f
C16685 net55 FILLER_0_11_78/a_484_472# 0.038269f
C16686 _016_ _114_ 0.041462f
C16687 FILLER_0_5_128/a_572_375# _133_ 0.00134f
C16688 mask\[3\] _099_ 0.10534f
C16689 output35/a_224_472# _435_/a_36_151# 0.001362f
C16690 _320_/a_1568_472# net79 0.001157f
C16691 _432_/a_796_472# net80 0.007731f
C16692 FILLER_0_9_28/a_2276_472# _077_ 0.003256f
C16693 en vss 0.466499f
C16694 _068_ _117_ 0.011659f
C16695 FILLER_0_18_177/a_1828_472# net21 0.001887f
C16696 fanout63/a_36_160# vdd 0.020165f
C16697 _425_/a_2248_156# calibrate 0.022237f
C16698 FILLER_0_9_142/a_36_472# vss 0.004305f
C16699 _216_/a_67_603# mask\[9\] 0.003086f
C16700 _248_/a_36_68# vdd 0.038887f
C16701 mask\[5\] FILLER_0_20_177/a_1380_472# 0.016114f
C16702 _012_ FILLER_0_21_60/a_124_375# 0.016032f
C16703 _118_ _121_ 0.02882f
C16704 _067_ cal_count\[0\] 0.201595f
C16705 FILLER_0_14_123/a_36_472# _043_ 0.001782f
C16706 mask\[7\] _433_/a_36_151# 0.001832f
C16707 _294_/a_224_472# mask\[3\] 0.00233f
C16708 _174_ _181_ 0.079407f
C16709 result[5] _418_/a_36_151# 0.009705f
C16710 _291_/a_36_160# vdd 0.010802f
C16711 _053_ FILLER_0_6_90/a_484_472# 0.011443f
C16712 net57 _385_/a_36_68# 0.03315f
C16713 _024_ _435_/a_1000_472# 0.002902f
C16714 _417_/a_2665_112# vdd 0.03015f
C16715 FILLER_0_9_72/a_1020_375# vss 0.005622f
C16716 FILLER_0_9_72/a_1468_375# vdd 0.026475f
C16717 result[7] result[5] 0.016166f
C16718 net64 _100_ 0.001674f
C16719 _111_ mask\[9\] 0.127919f
C16720 net20 _274_/a_1164_497# 0.002879f
C16721 net36 _195_/a_67_603# 0.034361f
C16722 _432_/a_2665_112# net21 0.005773f
C16723 _115_ _120_ 0.076035f
C16724 _128_ vss 0.859962f
C16725 ctlp[4] _009_ 0.004522f
C16726 input1/a_36_113# vss 0.05331f
C16727 _421_/a_2665_112# _419_/a_2248_156# 0.001545f
C16728 _428_/a_36_151# _451_/a_36_151# 0.003608f
C16729 _152_ _163_ 0.05157f
C16730 FILLER_0_5_72/a_484_472# net47 0.00169f
C16731 _187_ cal_count\[0\] 0.645851f
C16732 _453_/a_1000_472# vss 0.001738f
C16733 _311_/a_1212_473# vdd 0.001387f
C16734 cal_count\[2\] FILLER_0_15_2/a_36_472# 0.037661f
C16735 FILLER_0_22_128/a_2724_472# _146_ 0.002471f
C16736 _015_ _426_/a_1000_472# 0.033582f
C16737 _093_ _046_ 0.061989f
C16738 _008_ net64 0.001427f
C16739 _017_ _135_ 0.094281f
C16740 FILLER_0_17_200/a_572_375# mask\[3\] 0.013879f
C16741 net52 FILLER_0_2_101/a_36_472# 0.00749f
C16742 FILLER_0_3_204/a_124_375# FILLER_0_3_172/a_3260_375# 0.012001f
C16743 trim_mask\[4\] _160_ 0.244284f
C16744 FILLER_0_7_72/a_1020_375# FILLER_0_6_79/a_124_375# 0.026339f
C16745 FILLER_0_18_177/a_3172_472# net22 0.037136f
C16746 net47 _160_ 0.2966f
C16747 _136_ FILLER_0_16_154/a_124_375# 0.00252f
C16748 _098_ _437_/a_2248_156# 0.008669f
C16749 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_124_375# 0.012267f
C16750 _150_ _136_ 0.039815f
C16751 _415_/a_796_472# net81 0.002008f
C16752 net54 FILLER_0_22_128/a_1380_472# 0.008765f
C16753 mask\[8\] _213_/a_255_603# 0.002776f
C16754 net35 _213_/a_67_603# 0.012955f
C16755 FILLER_0_5_128/a_484_472# _081_ 0.00169f
C16756 _140_ _148_ 0.011699f
C16757 net32 _421_/a_1000_472# 0.002275f
C16758 FILLER_0_17_72/a_3172_472# _136_ 0.002925f
C16759 net81 FILLER_0_15_212/a_36_472# 0.003945f
C16760 mask\[0\] _429_/a_796_472# 0.007281f
C16761 _448_/a_2248_156# net59 0.005684f
C16762 _270_/a_36_472# _087_ 0.02676f
C16763 vss _433_/a_1308_423# 0.002695f
C16764 FILLER_0_8_107/a_36_472# _058_ 0.015262f
C16765 _005_ _192_/a_67_603# 0.013886f
C16766 _101_ mask\[1\] 0.033941f
C16767 _005_ vdd 0.506158f
C16768 _150_ _438_/a_1000_472# 0.003452f
C16769 FILLER_0_3_172/a_1020_375# net22 0.013048f
C16770 _415_/a_36_151# FILLER_0_8_263/a_124_375# 0.001619f
C16771 FILLER_0_18_53/a_124_375# vdd 0.022f
C16772 _094_ _418_/a_448_472# 0.042782f
C16773 _057_ _267_/a_36_472# 0.038568f
C16774 FILLER_0_18_107/a_932_472# FILLER_0_17_104/a_1380_472# 0.026657f
C16775 _052_ _424_/a_1204_472# 0.002681f
C16776 FILLER_0_16_57/a_1020_375# _131_ 0.012481f
C16777 net34 FILLER_0_22_177/a_572_375# 0.006974f
C16778 FILLER_0_18_107/a_1916_375# _433_/a_36_151# 0.002709f
C16779 _180_ _041_ 0.00244f
C16780 FILLER_0_8_263/a_36_472# calibrate 0.006968f
C16781 FILLER_0_5_117/a_124_375# vss 0.001764f
C16782 _413_/a_36_151# _002_ 0.0076f
C16783 FILLER_0_16_107/a_572_375# vss 0.055104f
C16784 net72 FILLER_0_17_64/a_36_472# 0.001145f
C16785 _136_ _043_ 0.040107f
C16786 FILLER_0_4_107/a_36_472# _157_ 0.005289f
C16787 _028_ FILLER_0_7_59/a_572_375# 0.00133f
C16788 net76 FILLER_0_6_177/a_484_472# 0.016333f
C16789 _445_/a_36_151# net40 0.007227f
C16790 FILLER_0_21_28/a_36_472# net40 0.032105f
C16791 _132_ FILLER_0_18_107/a_2724_472# 0.002229f
C16792 _093_ FILLER_0_17_72/a_2364_375# 0.010888f
C16793 net70 FILLER_0_13_100/a_124_375# 0.017886f
C16794 _321_/a_1602_69# _120_ 0.00262f
C16795 _008_ _418_/a_1308_423# 0.027229f
C16796 _436_/a_448_472# FILLER_0_22_128/a_124_375# 0.006782f
C16797 net15 _216_/a_255_603# 0.002146f
C16798 _008_ _006_ 0.02963f
C16799 net38 net55 0.10956f
C16800 net62 _043_ 0.00426f
C16801 FILLER_0_8_263/a_124_375# net64 0.004793f
C16802 output27/a_224_472# vss 0.027374f
C16803 net75 vdd 1.265616f
C16804 FILLER_0_13_142/a_124_375# _043_ 0.009328f
C16805 FILLER_0_20_177/a_572_375# vdd -0.001627f
C16806 FILLER_0_20_177/a_124_375# vss 0.002674f
C16807 _114_ FILLER_0_10_94/a_124_375# 0.040691f
C16808 net34 _435_/a_2560_156# 0.002967f
C16809 net64 FILLER_0_14_235/a_124_375# 0.046554f
C16810 _070_ _067_ 0.001869f
C16811 _430_/a_2665_112# fanout63/a_36_160# 0.010365f
C16812 _091_ _137_ 0.486022f
C16813 _008_ _103_ 0.092504f
C16814 net16 _447_/a_36_151# 0.133348f
C16815 _141_ FILLER_0_16_154/a_1020_375# 0.003441f
C16816 _341_/a_49_472# FILLER_0_16_154/a_572_375# 0.001643f
C16817 net74 _160_ 0.165289f
C16818 fanout53/a_36_160# net23 0.007461f
C16819 _396_/a_224_472# _177_ 0.001254f
C16820 net80 FILLER_0_18_177/a_1828_472# 0.00195f
C16821 FILLER_0_10_78/a_932_472# _439_/a_2665_112# 0.001182f
C16822 FILLER_0_20_15/a_572_375# vdd 0.003301f
C16823 net65 FILLER_0_1_266/a_36_472# 0.003529f
C16824 output44/a_224_472# FILLER_0_19_28/a_124_375# 0.005166f
C16825 _095_ _451_/a_2449_156# 0.001843f
C16826 _028_ _133_ 0.007084f
C16827 _321_/a_170_472# _118_ 0.034852f
C16828 _027_ net36 0.185347f
C16829 FILLER_0_17_226/a_36_472# vdd 0.087587f
C16830 output47/a_224_472# net47 0.023797f
C16831 cal_count\[2\] _452_/a_1353_112# 0.002558f
C16832 net20 FILLER_0_16_241/a_124_375# 0.002327f
C16833 FILLER_0_17_104/a_124_375# _451_/a_448_472# 0.001718f
C16834 FILLER_0_17_104/a_572_375# _451_/a_36_151# 0.001619f
C16835 FILLER_0_5_212/a_124_375# _081_ 0.01149f
C16836 _441_/a_448_472# vdd 0.007984f
C16837 _441_/a_36_151# vss 0.015116f
C16838 _053_ FILLER_0_7_104/a_932_472# 0.002529f
C16839 _063_ _165_ 0.021839f
C16840 net64 _060_ 0.05104f
C16841 net55 _424_/a_36_151# 0.007344f
C16842 net38 net17 1.634286f
C16843 net48 _056_ 0.001581f
C16844 _432_/a_2665_112# net80 0.041304f
C16845 _058_ FILLER_0_9_105/a_572_375# 0.003832f
C16846 net52 _442_/a_2665_112# 0.031179f
C16847 FILLER_0_18_177/a_3172_472# vdd 0.002358f
C16848 net55 _067_ 0.053438f
C16849 mask\[4\] FILLER_0_19_155/a_124_375# 0.043876f
C16850 _033_ FILLER_0_6_47/a_124_375# 0.002521f
C16851 _176_ FILLER_0_10_94/a_124_375# 0.009888f
C16852 _005_ _416_/a_1204_472# 0.014873f
C16853 net20 state\[0\] 0.396139f
C16854 net53 FILLER_0_16_154/a_124_375# 0.003458f
C16855 FILLER_0_9_60/a_484_472# vss 0.005321f
C16856 _273_/a_36_68# _090_ 0.034955f
C16857 _093_ _356_/a_36_472# 0.009235f
C16858 net25 _098_ 0.001267f
C16859 _098_ net23 0.036637f
C16860 ctlp[3] mask\[7\] 0.103955f
C16861 ctlp[1] _421_/a_796_472# 0.001754f
C16862 FILLER_0_7_162/a_36_472# vdd 0.026981f
C16863 vss _295_/a_36_472# 0.009751f
C16864 FILLER_0_17_142/a_124_375# _137_ 0.006974f
C16865 _429_/a_2665_112# _043_ 0.007641f
C16866 net41 net47 0.19549f
C16867 FILLER_0_17_218/a_484_472# vss 0.035317f
C16868 _285_/a_36_472# _099_ 0.040922f
C16869 FILLER_0_3_172/a_1020_375# vdd 0.009809f
C16870 _131_ _372_/a_170_472# 0.002967f
C16871 _094_ mask\[1\] 0.49634f
C16872 net75 net9 0.006945f
C16873 _443_/a_2665_112# net22 0.00621f
C16874 _159_ _160_ 0.021804f
C16875 net76 net4 0.024291f
C16876 _132_ _328_/a_36_113# 0.006002f
C16877 output43/a_224_472# net46 0.0215f
C16878 _095_ net36 0.127549f
C16879 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1468_375# 0.086635f
C16880 net16 _444_/a_36_151# 0.010514f
C16881 FILLER_0_9_28/a_3172_472# net68 0.007929f
C16882 FILLER_0_12_220/a_932_472# _223_/a_36_160# 0.001323f
C16883 fanout72/a_36_113# _449_/a_36_151# 0.032681f
C16884 output33/a_224_472# output18/a_224_472# 0.111946f
C16885 net50 _165_ 0.056964f
C16886 output28/a_224_472# net79 0.04262f
C16887 net48 _068_ 0.054333f
C16888 _423_/a_36_151# FILLER_0_23_44/a_36_472# 0.001723f
C16889 net66 net17 0.023639f
C16890 net78 mask\[7\] 0.001437f
C16891 net82 FILLER_0_2_171/a_124_375# 0.003818f
C16892 _115_ FILLER_0_9_72/a_932_472# 0.001837f
C16893 _050_ mask\[7\] 0.128172f
C16894 _098_ FILLER_0_15_212/a_484_472# 0.00912f
C16895 net53 _043_ 0.053033f
C16896 _428_/a_2560_156# net74 0.002759f
C16897 FILLER_0_21_28/a_3172_472# FILLER_0_21_60/a_36_472# 0.013276f
C16898 vss _416_/a_36_151# 0.044403f
C16899 net32 net18 0.028135f
C16900 _134_ _120_ 0.047627f
C16901 _067_ net17 0.17227f
C16902 _422_/a_448_472# _108_ 0.03293f
C16903 _154_ _160_ 0.395185f
C16904 _086_ _151_ 0.002442f
C16905 mask\[8\] _149_ 0.0498f
C16906 fanout82/a_36_113# net37 0.046126f
C16907 cal_count\[3\] vdd 1.020669f
C16908 FILLER_0_7_72/a_2724_472# _308_/a_848_380# 0.001797f
C16909 net63 fanout63/a_36_160# 0.011149f
C16910 result[2] FILLER_0_15_282/a_572_375# 0.0011f
C16911 _114_ FILLER_0_14_107/a_36_472# 0.00191f
C16912 _058_ _125_ 0.016525f
C16913 _422_/a_448_472# net19 0.003382f
C16914 net20 FILLER_0_24_274/a_36_472# 0.009746f
C16915 _363_/a_36_68# _153_ 0.008003f
C16916 _003_ _161_ 0.004981f
C16917 net23 _387_/a_36_113# 0.031688f
C16918 _059_ vdd 0.161836f
C16919 FILLER_0_19_47/a_36_472# _012_ 0.001667f
C16920 _098_ _434_/a_796_472# 0.001383f
C16921 net34 _106_ 0.013009f
C16922 net74 FILLER_0_13_80/a_124_375# 0.012889f
C16923 FILLER_0_14_91/a_124_375# _136_ 0.013064f
C16924 _210_/a_255_603# mask\[7\] 0.001329f
C16925 _118_ _122_ 0.046796f
C16926 _117_ _113_ 0.09166f
C16927 _089_ vdd 0.087336f
C16928 trim_mask\[2\] trim_mask\[1\] 0.002186f
C16929 _053_ net14 0.713784f
C16930 trim_val\[4\] _037_ 0.258184f
C16931 _114_ _311_/a_3220_473# 0.003283f
C16932 net52 FILLER_0_3_78/a_124_375# 0.017889f
C16933 _073_ net59 0.028673f
C16934 _140_ _207_/a_67_603# 0.014923f
C16935 _118_ _227_/a_36_160# 0.017547f
C16936 _132_ _428_/a_1000_472# 0.027767f
C16937 ctlp[3] _422_/a_2248_156# 0.001888f
C16938 _070_ net23 0.047632f
C16939 FILLER_0_5_109/a_124_375# _153_ 0.040726f
C16940 net50 net40 0.005105f
C16941 FILLER_0_7_72/a_124_375# FILLER_0_6_47/a_2812_375# 0.026339f
C16942 _053_ _164_ 0.058788f
C16943 _095_ _452_/a_36_151# 0.002974f
C16944 FILLER_0_4_197/a_572_375# net76 0.006026f
C16945 output14/a_224_472# FILLER_0_0_130/a_124_375# 0.00515f
C16946 trim[0] _446_/a_36_151# 0.044586f
C16947 net38 _446_/a_1308_423# 0.010331f
C16948 net49 FILLER_0_3_78/a_124_375# 0.001597f
C16949 _030_ FILLER_0_3_78/a_572_375# 0.007667f
C16950 net34 _147_ 0.144404f
C16951 _412_/a_448_472# net19 0.001526f
C16952 trimb[2] vdd 0.084666f
C16953 _320_/a_672_472# vdd 0.008437f
C16954 _274_/a_36_68# vss 0.052669f
C16955 trim_mask\[2\] _157_ 0.002951f
C16956 _069_ _248_/a_36_68# 0.058746f
C16957 net20 _198_/a_67_603# 0.013603f
C16958 net50 FILLER_0_6_79/a_124_375# 0.004402f
C16959 _213_/a_67_603# vdd 0.014901f
C16960 net82 FILLER_0_3_172/a_2724_472# 0.007912f
C16961 FILLER_0_21_206/a_36_472# net22 0.012952f
C16962 output34/a_224_472# _094_ 0.002719f
C16963 _346_/a_49_472# _141_ 0.104653f
C16964 _431_/a_36_151# FILLER_0_16_115/a_124_375# 0.035117f
C16965 FILLER_0_4_123/a_36_472# fanout69/a_36_113# 0.007864f
C16966 _405_/a_67_603# vss 0.008564f
C16967 _405_/a_255_603# vdd 0.001044f
C16968 net73 _131_ 0.022043f
C16969 vss FILLER_0_14_235/a_484_472# 0.003246f
C16970 _398_/a_36_113# cal_count\[2\] 0.004895f
C16971 _178_ _405_/a_67_603# 0.02427f
C16972 _101_ _099_ 0.198807f
C16973 _430_/a_1000_472# net63 0.016386f
C16974 net32 _048_ 0.008647f
C16975 FILLER_0_7_195/a_36_472# cal_itt\[3\] 0.070665f
C16976 _070_ FILLER_0_11_109/a_124_375# 0.002358f
C16977 _122_ _123_ 0.242965f
C16978 _115_ FILLER_0_9_105/a_572_375# 0.003191f
C16979 _443_/a_2248_156# vss 0.008696f
C16980 _443_/a_2665_112# vdd 0.011824f
C16981 FILLER_0_22_86/a_484_472# _437_/a_448_472# 0.008036f
C16982 FILLER_0_7_72/a_2364_375# _053_ 0.015932f
C16983 _123_ FILLER_0_7_233/a_124_375# 0.007717f
C16984 _073_ _122_ 0.002157f
C16985 comp FILLER_0_15_2/a_36_472# 0.001941f
C16986 FILLER_0_7_162/a_124_375# vdd 0.011809f
C16987 FILLER_0_19_28/a_124_375# vdd 0.028695f
C16988 cal_count\[3\] _135_ 0.039115f
C16989 _446_/a_1308_423# net66 0.005976f
C16990 FILLER_0_16_73/a_572_375# _040_ 0.014453f
C16991 _143_ _140_ 0.00806f
C16992 _429_/a_36_151# FILLER_0_13_206/a_36_472# 0.059367f
C16993 cal_count\[3\] _373_/a_244_68# 0.002341f
C16994 _008_ mask\[2\] 0.003475f
C16995 _404_/a_36_472# _182_ 0.036415f
C16996 _449_/a_2665_112# FILLER_0_13_80/a_124_375# 0.010688f
C16997 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001597f
C16998 trim_mask\[1\] FILLER_0_4_91/a_124_375# 0.006803f
C16999 _415_/a_2248_156# vdd 0.009114f
C17000 _423_/a_1000_472# vdd 0.001833f
C17001 _114_ vss 0.365613f
C17002 FILLER_0_22_177/a_36_472# _023_ 0.007019f
C17003 ctlp[4] net33 0.001734f
C17004 net63 FILLER_0_20_177/a_572_375# 0.00281f
C17005 _093_ _103_ 0.124026f
C17006 net57 _428_/a_2665_112# 0.027291f
C17007 _105_ net60 0.042726f
C17008 _430_/a_1000_472# _069_ 0.00929f
C17009 _086_ _162_ 0.107276f
C17010 net81 _019_ 0.004079f
C17011 net57 fanout53/a_36_160# 0.009946f
C17012 net62 result[2] 0.311075f
C17013 net74 _133_ 0.696379f
C17014 FILLER_0_16_89/a_1380_472# _136_ 0.009079f
C17015 net47 FILLER_0_5_164/a_36_472# 0.046908f
C17016 mask\[4\] FILLER_0_19_187/a_572_375# 0.00553f
C17017 net81 cal_itt\[1\] 0.387207f
C17018 FILLER_0_4_99/a_124_375# _365_/a_36_68# 0.001918f
C17019 net16 _054_ 0.044357f
C17020 FILLER_0_15_72/a_36_472# cal_count\[1\] 0.006408f
C17021 FILLER_0_7_72/a_124_375# FILLER_0_5_72/a_36_472# 0.001512f
C17022 FILLER_0_14_91/a_124_375# net53 0.065572f
C17023 FILLER_0_20_193/a_572_375# _434_/a_2665_112# 0.002362f
C17024 FILLER_0_7_72/a_2724_472# net14 0.012436f
C17025 _440_/a_36_151# FILLER_0_6_47/a_1380_472# 0.001512f
C17026 _345_/a_36_160# FILLER_0_19_111/a_572_375# 0.132282f
C17027 FILLER_0_17_72/a_1828_472# vdd 0.001969f
C17028 FILLER_0_17_72/a_1380_472# vss 0.003698f
C17029 _086_ _131_ 0.886615f
C17030 _093_ FILLER_0_18_61/a_36_472# 0.004039f
C17031 FILLER_0_20_169/a_124_375# _434_/a_36_151# 0.026916f
C17032 trimb[2] output17/a_224_472# 0.008375f
C17033 net82 _066_ 0.029681f
C17034 FILLER_0_5_136/a_36_472# vss 0.007658f
C17035 FILLER_0_12_20/a_36_472# _039_ 0.007881f
C17036 _115_ _125_ 0.049021f
C17037 mask\[5\] _204_/a_67_603# 0.023791f
C17038 FILLER_0_16_89/a_1020_375# _040_ 0.004252f
C17039 ctln[6] net69 0.003695f
C17040 FILLER_0_9_28/a_1380_472# net16 0.005297f
C17041 _114_ _308_/a_124_24# 0.052818f
C17042 FILLER_0_17_226/a_36_472# net63 0.001822f
C17043 trim[4] net67 0.06366f
C17044 _413_/a_1000_472# net59 0.018099f
C17045 _132_ FILLER_0_17_104/a_484_472# 0.002737f
C17046 FILLER_0_3_78/a_36_472# _164_ 0.022063f
C17047 _427_/a_2248_156# vss 0.018484f
C17048 _427_/a_2665_112# vdd 0.033395f
C17049 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001597f
C17050 net19 _420_/a_36_151# 0.016882f
C17051 net20 net79 0.046876f
C17052 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_572_375# 0.086635f
C17053 _372_/a_2034_472# _133_ 0.001257f
C17054 _372_/a_170_472# _076_ 0.049892f
C17055 _436_/a_36_151# FILLER_0_22_107/a_484_472# 0.001723f
C17056 net16 vss 0.679042f
C17057 net16 _178_ 0.30147f
C17058 _398_/a_36_113# _043_ 0.005985f
C17059 net76 FILLER_0_3_172/a_1468_375# 0.039469f
C17060 _176_ vss 0.761803f
C17061 net57 _098_ 0.062604f
C17062 FILLER_0_5_212/a_36_472# net59 0.058827f
C17063 net82 net23 0.18994f
C17064 FILLER_0_21_206/a_36_472# vdd 0.00971f
C17065 FILLER_0_21_206/a_124_375# vss 0.05074f
C17066 output13/a_224_472# _448_/a_2665_112# 0.027303f
C17067 FILLER_0_5_128/a_484_472# _163_ 0.009861f
C17068 net4 FILLER_0_12_236/a_124_375# 0.001558f
C17069 output37/a_224_472# en 0.003788f
C17070 result[9] _420_/a_2665_112# 0.037019f
C17071 FILLER_0_6_90/a_124_375# _163_ 0.013948f
C17072 _094_ _099_ 0.193065f
C17073 FILLER_0_8_107/a_36_472# _134_ 0.005632f
C17074 _035_ _380_/a_224_472# 0.001921f
C17075 _411_/a_2248_156# net58 0.014884f
C17076 FILLER_0_18_107/a_3260_375# _145_ 0.00346f
C17077 FILLER_0_4_49/a_124_375# net47 0.006524f
C17078 mask\[7\] _435_/a_36_151# 0.037736f
C17079 net72 _052_ 0.138281f
C17080 fanout69/a_36_113# net69 0.040451f
C17081 net22 FILLER_0_18_209/a_124_375# 0.012909f
C17082 net25 FILLER_0_22_86/a_124_375# 0.004298f
C17083 net46 FILLER_0_20_15/a_1020_375# 0.0302f
C17084 _128_ FILLER_0_12_236/a_36_472# 0.001043f
C17085 _091_ FILLER_0_19_171/a_484_472# 0.013944f
C17086 _373_/a_1458_68# _113_ 0.001257f
C17087 _124_ vss 0.110847f
C17088 _443_/a_2665_112# FILLER_0_2_165/a_124_375# 0.006271f
C17089 _133_ _154_ 0.0133f
C17090 _053_ _372_/a_3126_472# 0.001056f
C17091 net80 _435_/a_36_151# 0.035259f
C17092 FILLER_0_18_139/a_124_375# vdd 0.023256f
C17093 mask\[0\] FILLER_0_14_235/a_572_375# 0.002003f
C17094 net28 _005_ 0.080653f
C17095 FILLER_0_9_72/a_572_375# _439_/a_36_151# 0.059049f
C17096 _091_ fanout56/a_36_113# 0.001254f
C17097 FILLER_0_5_72/a_1468_375# _440_/a_2248_156# 0.030666f
C17098 FILLER_0_5_72/a_1020_375# _440_/a_2665_112# 0.010688f
C17099 _077_ FILLER_0_9_72/a_484_472# 0.004472f
C17100 net19 _419_/a_448_472# 0.037199f
C17101 FILLER_0_15_282/a_124_375# output30/a_224_472# 0.029138f
C17102 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_36_472# 0.001723f
C17103 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_572_375# 0.026339f
C17104 FILLER_0_0_130/a_124_375# vdd 0.012493f
C17105 FILLER_0_5_212/a_36_472# _122_ 0.002272f
C17106 FILLER_0_12_28/a_36_472# _039_ 0.007926f
C17107 _405_/a_67_603# _184_ 0.010046f
C17108 _039_ net40 0.036781f
C17109 _036_ _441_/a_36_151# 0.005754f
C17110 fanout80/a_36_113# _138_ 0.002489f
C17111 fanout71/a_36_113# vss 0.007654f
C17112 _074_ _305_/a_36_159# 0.012602f
C17113 _064_ output39/a_224_472# 0.107406f
C17114 _187_ _408_/a_1336_472# 0.002191f
C17115 net20 _429_/a_2560_156# 0.002069f
C17116 _140_ _348_/a_257_69# 0.001089f
C17117 FILLER_0_1_204/a_124_375# net21 0.008041f
C17118 _077_ _453_/a_2665_112# 0.002824f
C17119 net18 FILLER_0_9_282/a_36_472# 0.041571f
C17120 net71 _437_/a_796_472# 0.006933f
C17121 net57 _070_ 0.202843f
C17122 _435_/a_796_472# vdd 0.003478f
C17123 net38 _444_/a_1308_423# 0.007915f
C17124 FILLER_0_15_142/a_572_375# FILLER_0_15_150/a_36_472# 0.086635f
C17125 _432_/a_36_151# net57 0.00484f
C17126 FILLER_0_17_72/a_124_375# FILLER_0_15_72/a_36_472# 0.001512f
C17127 FILLER_0_21_142/a_124_375# _433_/a_2560_156# 0.001178f
C17128 FILLER_0_20_87/a_36_472# _438_/a_448_472# 0.004782f
C17129 _053_ _153_ 0.015583f
C17130 _103_ _418_/a_1204_472# 0.00582f
C17131 net81 fanout79/a_36_160# 0.057526f
C17132 _013_ _183_ 0.00176f
C17133 net69 _371_/a_36_113# 0.016091f
C17134 net2 net59 0.334636f
C17135 _449_/a_2560_156# net55 0.004835f
C17136 _068_ net37 0.006392f
C17137 FILLER_0_18_76/a_124_375# vss 0.006877f
C17138 FILLER_0_18_76/a_572_375# vdd -0.009037f
C17139 _443_/a_36_151# trim_mask\[4\] 0.002625f
C17140 _087_ _074_ 0.004231f
C17141 _069_ cal_count\[3\] 0.012382f
C17142 _134_ FILLER_0_9_105/a_572_375# 0.02163f
C17143 _083_ FILLER_0_3_221/a_1380_472# 0.00181f
C17144 output42/a_224_472# net17 0.047757f
C17145 _099_ FILLER_0_14_235/a_572_375# 0.013281f
C17146 _069_ _059_ 0.002034f
C17147 _320_/a_36_472# _055_ 0.001393f
C17148 FILLER_0_16_107/a_484_472# FILLER_0_16_115/a_36_472# 0.013276f
C17149 mask\[3\] net56 0.002632f
C17150 _016_ _428_/a_448_472# 0.00347f
C17151 FILLER_0_10_78/a_932_472# FILLER_0_9_72/a_1468_375# 0.001543f
C17152 net78 _419_/a_2248_156# 0.001614f
C17153 output37/a_224_472# output27/a_224_472# 0.012653f
C17154 output14/a_224_472# net52 0.02346f
C17155 FILLER_0_6_90/a_36_472# FILLER_0_4_91/a_124_375# 0.001188f
C17156 _448_/a_2248_156# trim_val\[4\] 0.001534f
C17157 net38 _452_/a_2449_156# 0.058386f
C17158 net27 result[1] 0.187252f
C17159 net57 net55 0.001926f
C17160 _371_/a_36_113# _152_ 0.001083f
C17161 _131_ _451_/a_3129_107# 0.001608f
C17162 FILLER_0_21_142/a_124_375# vss 0.009345f
C17163 output33/a_224_472# net18 0.110644f
C17164 _128_ _426_/a_2248_156# 0.019019f
C17165 _114_ _071_ 0.040513f
C17166 FILLER_0_9_28/a_1020_375# vdd 0.033815f
C17167 FILLER_0_21_28/a_2812_375# vdd -0.014642f
C17168 FILLER_0_18_209/a_124_375# vdd 0.023676f
C17169 _040_ net14 0.069672f
C17170 _086_ _074_ 0.186795f
C17171 _320_/a_1120_472# _043_ 0.002242f
C17172 fanout58/a_36_160# input4/a_36_68# 0.059453f
C17173 _413_/a_448_472# _002_ 0.044695f
C17174 _093_ mask\[2\] 0.009354f
C17175 _077_ FILLER_0_9_105/a_124_375# 0.007189f
C17176 _016_ FILLER_0_12_124/a_36_472# 0.002661f
C17177 _041_ vss 0.012963f
C17178 _126_ _320_/a_36_472# 0.026216f
C17179 net16 _184_ 0.028159f
C17180 FILLER_0_21_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001723f
C17181 _402_/a_1948_68# _182_ 0.016049f
C17182 net36 FILLER_0_20_87/a_124_375# 0.005853f
C17183 cal_itt\[2\] _080_ 0.062471f
C17184 _189_/a_67_603# net64 0.064691f
C17185 net49 _167_ 0.031111f
C17186 _086_ _076_ 0.79237f
C17187 FILLER_0_2_93/a_124_375# _030_ 0.001641f
C17188 net36 _451_/a_448_472# 0.042223f
C17189 _176_ _401_/a_36_68# 0.004263f
C17190 trim_val\[1\] FILLER_0_5_54/a_124_375# 0.001814f
C17191 _053_ _439_/a_2665_112# 0.006037f
C17192 _415_/a_2560_156# net18 0.010318f
C17193 net27 FILLER_0_12_236/a_484_472# 0.042937f
C17194 _354_/a_49_472# _433_/a_36_151# 0.001715f
C17195 fanout63/a_36_160# _282_/a_36_160# 0.23939f
C17196 _125_ _134_ 0.00437f
C17197 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_124_375# 0.016748f
C17198 FILLER_0_4_107/a_484_472# net47 0.001975f
C17199 _267_/a_36_472# vss 0.001495f
C17200 _091_ _430_/a_796_472# 0.005465f
C17201 fanout62/a_36_160# net18 0.008106f
C17202 valid net59 0.577796f
C17203 net81 _429_/a_1000_472# 0.011018f
C17204 FILLER_0_18_209/a_484_472# _047_ 0.002188f
C17205 _139_ FILLER_0_15_180/a_484_472# 0.004763f
C17206 _095_ _405_/a_67_603# 0.012596f
C17207 output38/a_224_472# output39/a_224_472# 0.002978f
C17208 output28/a_224_472# net19 0.101711f
C17209 mask\[7\] _350_/a_257_69# 0.001135f
C17210 net74 _443_/a_36_151# 0.003682f
C17211 _052_ FILLER_0_17_38/a_484_472# 0.001368f
C17212 net15 _174_ 0.090215f
C17213 result[5] _007_ 0.0249f
C17214 _449_/a_36_151# cal_count\[3\] 0.018365f
C17215 trim_mask\[2\] net66 0.036211f
C17216 _427_/a_2248_156# _071_ 0.001131f
C17217 _430_/a_1204_472# net21 0.006991f
C17218 FILLER_0_13_212/a_1380_472# FILLER_0_13_228/a_36_472# 0.013277f
C17219 net82 FILLER_0_3_142/a_36_472# 0.0172f
C17220 FILLER_0_3_172/a_2724_472# net21 0.009426f
C17221 net14 FILLER_0_10_94/a_572_375# 0.047331f
C17222 net52 net22 0.017993f
C17223 net20 _430_/a_2248_156# 0.001893f
C17224 _305_/a_36_159# _081_ 0.039192f
C17225 _176_ _071_ 0.002542f
C17226 FILLER_0_17_72/a_1380_472# _027_ 0.00378f
C17227 FILLER_0_17_72/a_2276_472# _150_ 0.003968f
C17228 net70 _451_/a_1353_112# 0.00194f
C17229 net52 FILLER_0_9_72/a_1380_472# 0.003507f
C17230 FILLER_0_13_142/a_932_472# net23 0.020589f
C17231 fanout72/a_36_113# _394_/a_56_524# 0.002775f
C17232 FILLER_0_19_55/a_124_375# vss 0.001882f
C17233 FILLER_0_19_55/a_36_472# vdd 0.085984f
C17234 FILLER_0_21_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001723f
C17235 _425_/a_1000_472# net37 0.002879f
C17236 net81 FILLER_0_10_247/a_124_375# 0.044906f
C17237 net57 net82 0.91473f
C17238 net72 net40 0.001815f
C17239 net31 _047_ 0.029502f
C17240 _340_/a_36_160# _098_ 0.019601f
C17241 FILLER_0_13_80/a_36_472# _451_/a_3129_107# 0.001115f
C17242 _093_ FILLER_0_16_115/a_124_375# 0.003988f
C17243 net75 _426_/a_1204_472# 0.001592f
C17244 _114_ _095_ 0.001338f
C17245 net57 fanout57/a_36_113# 0.004316f
C17246 FILLER_0_15_142/a_124_375# _427_/a_36_151# 0.059049f
C17247 _187_ _410_/a_36_68# 0.038745f
C17248 _085_ _055_ 0.240451f
C17249 trim_mask\[4\] net59 0.012971f
C17250 net81 FILLER_0_15_228/a_124_375# 0.006974f
C17251 _414_/a_2665_112# vss 0.010021f
C17252 output29/a_224_472# vss 0.013148f
C17253 _087_ _081_ 0.002169f
C17254 _142_ _137_ 1.401722f
C17255 net82 FILLER_0_3_221/a_932_472# 0.004092f
C17256 _426_/a_36_151# vss 0.003014f
C17257 _426_/a_448_472# vdd 0.042167f
C17258 _098_ _438_/a_1308_423# 0.004124f
C17259 _092_ vss 0.346097f
C17260 FILLER_0_8_247/a_484_472# calibrate 0.009318f
C17261 _077_ _251_/a_468_472# 0.002497f
C17262 FILLER_0_12_220/a_1468_375# _060_ 0.001429f
C17263 FILLER_0_12_220/a_484_472# _090_ 0.006993f
C17264 _412_/a_2560_156# net5 0.007446f
C17265 _432_/a_1308_423# vdd 0.029938f
C17266 _337_/a_49_472# mask\[2\] 0.00188f
C17267 FILLER_0_16_89/a_1468_375# vss 0.048986f
C17268 FILLER_0_16_89/a_36_472# vdd 0.040085f
C17269 fanout66/a_36_113# _440_/a_36_151# 0.017895f
C17270 trim_mask\[2\] FILLER_0_3_54/a_124_375# 0.015198f
C17271 valid net64 0.022969f
C17272 _431_/a_1308_423# vss 0.003472f
C17273 _088_ net82 0.160444f
C17274 _233_/a_36_160# vdd 0.064615f
C17275 _427_/a_36_151# net74 0.04306f
C17276 FILLER_0_2_93/a_572_375# net14 0.044606f
C17277 _175_ FILLER_0_15_72/a_36_472# 0.006746f
C17278 net72 FILLER_0_17_38/a_572_375# 0.010272f
C17279 ctlp[4] net22 0.257841f
C17280 FILLER_0_17_64/a_124_375# vss 0.022351f
C17281 FILLER_0_17_64/a_36_472# vdd 0.094397f
C17282 fanout53/a_36_160# net36 0.028652f
C17283 _075_ _414_/a_2665_112# 0.050503f
C17284 _190_/a_36_160# _043_ 0.06415f
C17285 _077_ _188_ 0.1656f
C17286 FILLER_0_17_142/a_572_375# vss 0.049716f
C17287 FILLER_0_17_142/a_36_472# vdd 0.108843f
C17288 net58 cal_itt\[0\] 0.229955f
C17289 FILLER_0_6_47/a_572_375# vdd 0.003158f
C17290 _106_ FILLER_0_17_218/a_484_472# 0.012952f
C17291 trim[0] vss 0.132654f
C17292 FILLER_0_5_109/a_484_472# FILLER_0_5_117/a_36_472# 0.013276f
C17293 _321_/a_170_472# net74 0.020269f
C17294 _072_ FILLER_0_10_214/a_124_375# 0.033245f
C17295 _427_/a_2248_156# _095_ 0.022479f
C17296 _126_ _085_ 0.02154f
C17297 FILLER_0_2_93/a_124_375# trim_mask\[3\] 0.003033f
C17298 _093_ FILLER_0_19_111/a_572_375# 0.002743f
C17299 _053_ FILLER_0_6_47/a_2724_472# 0.001777f
C17300 mask\[9\] FILLER_0_19_111/a_124_375# 0.031474f
C17301 net16 _095_ 0.042842f
C17302 _086_ _081_ 0.033115f
C17303 FILLER_0_16_255/a_36_472# _417_/a_2665_112# 0.003221f
C17304 FILLER_0_24_290/a_124_375# FILLER_0_24_274/a_1468_375# 0.012001f
C17305 _176_ _095_ 0.064978f
C17306 output15/a_224_472# _383_/a_36_472# 0.001154f
C17307 net42 net6 0.166896f
C17308 FILLER_0_3_142/a_124_375# _443_/a_36_151# 0.059049f
C17309 calibrate net23 0.032259f
C17310 _130_ _127_ 0.195571f
C17311 clk rstn 0.541051f
C17312 fanout54/a_36_160# net23 0.05522f
C17313 net75 FILLER_0_6_231/a_484_472# 0.003485f
C17314 _339_/a_36_160# vdd 0.01226f
C17315 _272_/a_36_472# _003_ 0.001634f
C17316 _162_ _061_ 0.001665f
C17317 net16 _036_ 0.637538f
C17318 _122_ net47 0.030693f
C17319 _141_ _098_ 0.0697f
C17320 _050_ _436_/a_448_472# 0.064832f
C17321 _045_ _006_ 0.00216f
C17322 FILLER_0_16_37/a_36_472# net47 0.008304f
C17323 FILLER_0_10_78/a_572_375# _176_ 0.005927f
C17324 _098_ _348_/a_49_472# 0.011096f
C17325 _301_/a_36_472# _098_ 0.010091f
C17326 net52 vdd 1.32956f
C17327 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_572_375# 0.086635f
C17328 _415_/a_2665_112# vdd 0.017004f
C17329 net36 _098_ 3.387566f
C17330 _413_/a_2248_156# FILLER_0_3_212/a_124_375# 0.030666f
C17331 FILLER_0_8_24/a_36_472# net47 0.097212f
C17332 FILLER_0_10_78/a_124_375# _453_/a_2665_112# 0.006271f
C17333 _076_ _313_/a_67_603# 0.024219f
C17334 _127_ _129_ 0.716384f
C17335 FILLER_0_17_104/a_36_472# _438_/a_2248_156# 0.001731f
C17336 _139_ _138_ 0.00256f
C17337 FILLER_0_18_107/a_1828_472# vdd 0.004446f
C17338 cal_itt\[0\] _082_ 0.018597f
C17339 _256_/a_36_68# _072_ 0.027152f
C17340 _434_/a_2665_112# mask\[6\] 0.026286f
C17341 trim_mask\[4\] _169_ 0.042442f
C17342 net35 _434_/a_2248_156# 0.026885f
C17343 _010_ FILLER_0_23_274/a_36_472# 0.008718f
C17344 net82 cal_itt\[0\] 0.063072f
C17345 cal_itt\[2\] vss 0.249871f
C17346 FILLER_0_7_104/a_1380_472# vss 0.003236f
C17347 mask\[4\] _201_/a_255_603# 0.002111f
C17348 _102_ vdd 0.211559f
C17349 _285_/a_36_472# _196_/a_36_160# 0.004619f
C17350 _424_/a_796_472# vdd 0.001951f
C17351 FILLER_0_17_104/a_572_375# _040_ 0.001228f
C17352 _413_/a_36_151# FILLER_0_3_172/a_1916_375# 0.059049f
C17353 FILLER_0_8_138/a_124_375# _120_ 0.12254f
C17354 _030_ vss 0.117034f
C17355 net49 vdd 0.872948f
C17356 net47 _169_ 0.528536f
C17357 _320_/a_36_472# state\[1\] 0.013058f
C17358 output29/a_224_472# _416_/a_2248_156# 0.024448f
C17359 net50 _168_ 0.306226f
C17360 mask\[4\] FILLER_0_18_177/a_1380_472# 0.016924f
C17361 _104_ net61 1.149805f
C17362 _122_ FILLER_0_5_172/a_124_375# 0.001352f
C17363 _027_ FILLER_0_18_76/a_124_375# 0.001285f
C17364 net20 FILLER_0_6_239/a_124_375# 0.004897f
C17365 _173_ _408_/a_728_93# 0.022838f
C17366 net50 _441_/a_796_472# 0.010626f
C17367 FILLER_0_4_107/a_484_472# _154_ 0.040595f
C17368 _129_ FILLER_0_11_135/a_36_472# 0.078373f
C17369 mask\[3\] FILLER_0_18_177/a_484_472# 0.005654f
C17370 FILLER_0_19_47/a_124_375# FILLER_0_18_37/a_1380_472# 0.001684f
C17371 _429_/a_2248_156# FILLER_0_13_228/a_36_472# 0.035805f
C17372 _272_/a_36_472# net37 0.002669f
C17373 net61 vss 0.254538f
C17374 net18 _417_/a_1000_472# 0.056791f
C17375 FILLER_0_16_57/a_124_375# net15 0.001594f
C17376 _417_/a_1204_472# net30 0.001496f
C17377 _417_/a_796_472# result[3] 0.001206f
C17378 _062_ _055_ 0.29425f
C17379 _072_ _162_ 0.090175f
C17380 net20 _108_ 0.125627f
C17381 FILLER_0_18_2/a_1380_472# net55 0.007469f
C17382 output36/a_224_472# FILLER_0_15_282/a_124_375# 0.002977f
C17383 _441_/a_2248_156# _030_ 0.003495f
C17384 ctlp[5] output22/a_224_472# 0.024131f
C17385 _149_ _026_ 0.243704f
C17386 _207_/a_67_603# _049_ 0.003205f
C17387 FILLER_0_21_28/a_2276_472# _423_/a_448_472# 0.008036f
C17388 FILLER_0_8_239/a_124_375# vdd 0.035205f
C17389 _428_/a_36_151# FILLER_0_14_107/a_484_472# 0.059367f
C17390 net20 net19 0.384932f
C17391 net69 FILLER_0_2_111/a_1020_375# 0.018655f
C17392 _031_ FILLER_0_2_111/a_124_375# 0.05482f
C17393 FILLER_0_5_128/a_124_375# _160_ 0.001157f
C17394 FILLER_0_6_239/a_124_375# FILLER_0_6_231/a_572_375# 0.012001f
C17395 net61 _422_/a_1000_472# 0.001947f
C17396 FILLER_0_18_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001684f
C17397 net34 output35/a_224_472# 0.0731f
C17398 FILLER_0_4_144/a_36_472# _370_/a_848_380# 0.15783f
C17399 net38 output6/a_224_472# 0.060017f
C17400 ctlp[4] vdd 0.278868f
C17401 _144_ _146_ 0.333799f
C17402 _098_ FILLER_0_15_228/a_36_472# 0.022074f
C17403 FILLER_0_16_107/a_124_375# net14 0.004684f
C17404 _267_/a_36_472# _071_ 0.001682f
C17405 net67 _190_/a_36_160# 0.023989f
C17406 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_36_472# 0.002296f
C17407 FILLER_0_12_136/a_1020_375# FILLER_0_13_142/a_484_472# 0.001684f
C17408 _110_ _437_/a_36_151# 0.00125f
C17409 net35 _025_ 0.02169f
C17410 output46/a_224_472# FILLER_0_20_15/a_124_375# 0.029497f
C17411 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_36_472# 0.002296f
C17412 _143_ _137_ 0.009932f
C17413 _028_ FILLER_0_7_104/a_572_375# 0.003664f
C17414 FILLER_0_7_195/a_124_375# _161_ 0.005368f
C17415 net16 _402_/a_1296_93# 0.053493f
C17416 _432_/a_36_151# _141_ 0.008193f
C17417 trimb[3] vss 0.161605f
C17418 _114_ _332_/a_36_472# 0.021351f
C17419 net73 _427_/a_448_472# 0.00132f
C17420 net15 FILLER_0_15_59/a_124_375# 0.007439f
C17421 net36 FILLER_0_15_180/a_124_375# 0.004275f
C17422 _406_/a_36_159# _278_/a_36_160# 0.001331f
C17423 _086_ FILLER_0_5_117/a_36_472# 0.042352f
C17424 FILLER_0_18_2/a_1380_472# net17 0.003603f
C17425 FILLER_0_14_91/a_36_472# _176_ 0.076419f
C17426 _359_/a_36_488# vss 0.002427f
C17427 net73 _145_ 0.009144f
C17428 FILLER_0_22_177/a_1468_375# _435_/a_36_151# 0.059049f
C17429 net51 _450_/a_3129_107# 0.030082f
C17430 _086_ _090_ 0.065807f
C17431 net27 net81 1.118985f
C17432 FILLER_0_13_228/a_124_375# net4 0.002641f
C17433 _406_/a_36_159# vss 0.002509f
C17434 net57 FILLER_0_13_142/a_932_472# 0.01158f
C17435 _178_ _406_/a_36_159# 0.007052f
C17436 mask\[7\] net23 0.225177f
C17437 FILLER_0_21_125/a_36_472# vdd 0.007233f
C17438 FILLER_0_21_125/a_572_375# vss 0.054783f
C17439 FILLER_0_15_72/a_572_375# vdd 0.003801f
C17440 FILLER_0_15_72/a_124_375# vss 0.048711f
C17441 FILLER_0_17_200/a_36_472# vdd 0.001039f
C17442 _101_ _196_/a_36_160# 0.009836f
C17443 _091_ FILLER_0_16_154/a_1468_375# 0.003056f
C17444 _028_ FILLER_0_7_72/a_1828_472# 0.001777f
C17445 FILLER_0_20_193/a_572_375# mask\[6\] 0.001262f
C17446 _053_ FILLER_0_6_177/a_36_472# 0.00572f
C17447 FILLER_0_24_130/a_124_375# vss 0.018125f
C17448 net43 FILLER_0_20_15/a_572_375# 0.003924f
C17449 net10 FILLER_0_0_232/a_36_472# 0.016287f
C17450 _053_ _376_/a_36_160# 0.005109f
C17451 _091_ _055_ 0.003332f
C17452 result[4] output31/a_224_472# 0.049147f
C17453 _067_ output6/a_224_472# 0.001611f
C17454 trim_mask\[3\] vss 0.156544f
C17455 net52 FILLER_0_2_165/a_124_375# 0.002214f
C17456 FILLER_0_8_247/a_1380_472# vss 0.001338f
C17457 net47 FILLER_0_4_91/a_572_375# 0.008167f
C17458 comp _190_/a_36_160# 0.001891f
C17459 input2/a_36_113# rstn 0.002202f
C17460 _095_ _041_ 0.002104f
C17461 _085_ state\[1\] 0.182697f
C17462 _441_/a_2665_112# net14 0.00104f
C17463 net55 net36 0.273956f
C17464 _083_ _260_/a_244_472# 0.00134f
C17465 _412_/a_448_472# fanout81/a_36_160# 0.00998f
C17466 net81 _425_/a_2665_112# 0.010188f
C17467 net55 FILLER_0_18_37/a_932_472# 0.00769f
C17468 _035_ _446_/a_36_151# 0.012914f
C17469 net15 trim_val\[3\] 0.068273f
C17470 _430_/a_2560_156# vss 0.002924f
C17471 _067_ _171_ 0.007069f
C17472 net72 FILLER_0_17_56/a_36_472# 0.008058f
C17473 net78 _421_/a_1000_472# 0.022212f
C17474 _229_/a_224_472# net22 0.007346f
C17475 _070_ FILLER_0_10_107/a_572_375# 0.003959f
C17476 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_484_472# 0.001723f
C17477 net38 net3 0.103189f
C17478 _441_/a_2665_112# _164_ 0.021931f
C17479 FILLER_0_3_221/a_484_472# net59 0.001655f
C17480 _428_/a_1308_423# vdd 0.004352f
C17481 _098_ _433_/a_1308_423# 0.010653f
C17482 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_36_472# 0.007947f
C17483 net22 _202_/a_36_160# 0.052766f
C17484 net38 _450_/a_1293_527# 0.001307f
C17485 _011_ _422_/a_1204_472# 0.002176f
C17486 net4 _078_ 0.487587f
C17487 _437_/a_36_151# net14 0.014361f
C17488 net13 vss 0.071697f
C17489 _127_ FILLER_0_11_135/a_124_375# 0.040456f
C17490 _182_ FILLER_0_18_37/a_1380_472# 0.004074f
C17491 _079_ net59 0.102335f
C17492 net1 _265_/a_916_472# 0.002088f
C17493 FILLER_0_5_109/a_484_472# _163_ 0.005054f
C17494 ctlp[9] FILLER_0_23_44/a_932_472# 0.001195f
C17495 trimb[1] FILLER_0_18_2/a_1020_375# 0.01376f
C17496 _086_ _321_/a_2034_472# 0.001815f
C17497 output9/a_224_472# vss 0.007544f
C17498 FILLER_0_9_28/a_1828_472# _120_ 0.00108f
C17499 FILLER_0_11_142/a_124_375# net23 0.002992f
C17500 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_484_472# 0.013277f
C17501 _119_ _118_ 0.001596f
C17502 _074_ _061_ 0.007152f
C17503 _422_/a_448_472# _009_ 0.018984f
C17504 _105_ output19/a_224_472# 0.107668f
C17505 net80 _434_/a_796_472# 0.039593f
C17506 FILLER_0_16_57/a_932_472# vss 0.003388f
C17507 FILLER_0_16_57/a_1380_472# vdd 0.005673f
C17508 net57 calibrate 0.037299f
C17509 _132_ FILLER_0_14_107/a_1468_375# 0.019517f
C17510 _112_ _316_/a_1152_472# 0.001449f
C17511 ctln[1] _411_/a_2665_112# 0.004748f
C17512 _028_ FILLER_0_7_72/a_932_472# 0.001777f
C17513 FILLER_0_12_124/a_36_472# vss 0.001443f
C17514 cal_count\[3\] FILLER_0_11_124/a_124_375# 0.002147f
C17515 _127_ _068_ 0.052712f
C17516 _128_ _070_ 1.279188f
C17517 _131_ _331_/a_244_472# 0.002331f
C17518 net15 _449_/a_1000_472# 0.056791f
C17519 _091_ FILLER_0_12_220/a_572_375# 0.003075f
C17520 FILLER_0_20_177/a_124_375# _098_ 0.018701f
C17521 _061_ _076_ 0.024289f
C17522 FILLER_0_15_212/a_1380_472# vss 0.007595f
C17523 _246_/a_36_68# vss 0.024639f
C17524 mask\[4\] _343_/a_49_472# 0.036987f
C17525 FILLER_0_15_212/a_484_472# mask\[1\] 0.007258f
C17526 FILLER_0_10_214/a_36_472# _060_ 0.001378f
C17527 net55 _452_/a_36_151# 0.042427f
C17528 _076_ _311_/a_66_473# 0.003077f
C17529 _086_ _318_/a_224_472# 0.007024f
C17530 _341_/a_49_472# _137_ 0.059288f
C17531 net20 _419_/a_448_472# 0.025583f
C17532 _281_/a_672_472# vdd 0.001069f
C17533 cal net58 0.001209f
C17534 _094_ net18 0.468109f
C17535 _425_/a_36_151# _316_/a_124_24# 0.036238f
C17536 _414_/a_1000_472# net21 0.042244f
C17537 net54 _436_/a_1308_423# 0.002665f
C17538 _065_ _447_/a_2248_156# 0.038629f
C17539 _245_/a_234_472# net47 0.00188f
C17540 net34 ctlp[2] 0.953441f
C17541 net57 _333_/a_36_160# 0.008292f
C17542 _392_/a_36_68# _120_ 0.001738f
C17543 mask\[9\] _354_/a_49_472# 0.032687f
C17544 trim_mask\[1\] FILLER_0_6_47/a_36_472# 0.004319f
C17545 _073_ FILLER_0_3_221/a_1020_375# 0.002563f
C17546 _086_ _314_/a_224_472# 0.003715f
C17547 _434_/a_2248_156# vdd 0.019386f
C17548 FILLER_0_5_88/a_36_472# _164_ 0.011718f
C17549 _094_ _196_/a_36_160# 0.001668f
C17550 _079_ _122_ 0.003853f
C17551 cal_itt\[1\] net59 0.227495f
C17552 net81 FILLER_0_14_235/a_36_472# 0.002571f
C17553 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_124_375# 0.009654f
C17554 _002_ net22 0.038848f
C17555 _009_ _108_ 1.645945f
C17556 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_572_375# 0.026339f
C17557 _072_ _074_ 2.017168f
C17558 result[7] FILLER_0_23_274/a_124_375# 0.017938f
C17559 _421_/a_36_151# _419_/a_36_151# 0.561555f
C17560 FILLER_0_8_127/a_36_472# vss 0.004344f
C17561 _043_ FILLER_0_12_196/a_124_375# 0.003935f
C17562 output13/a_224_472# net23 0.00255f
C17563 output27/a_224_472# fanout64/a_36_160# 0.027335f
C17564 FILLER_0_15_290/a_36_472# vdd 0.092839f
C17565 FILLER_0_15_290/a_124_375# vss 0.032056f
C17566 net19 _009_ 0.055383f
C17567 _088_ net21 0.053843f
C17568 output8/a_224_472# FILLER_0_3_221/a_932_472# 0.001699f
C17569 vdd FILLER_0_8_156/a_36_472# 0.002891f
C17570 vss FILLER_0_8_156/a_572_375# 0.007969f
C17571 state\[1\] _062_ 0.001179f
C17572 net58 en 0.029072f
C17573 FILLER_0_13_65/a_124_375# _067_ 0.001283f
C17574 _077_ FILLER_0_11_64/a_124_375# 0.013507f
C17575 cal_count\[3\] FILLER_0_12_50/a_36_472# 0.063276f
C17576 net35 FILLER_0_22_128/a_2364_375# 0.012732f
C17577 net17 _452_/a_36_151# 0.041497f
C17578 _412_/a_36_151# net1 0.020184f
C17579 _087_ _163_ 0.004829f
C17580 output32/a_224_472# _419_/a_36_151# 0.129117f
C17581 _072_ _076_ 0.068172f
C17582 FILLER_0_18_100/a_36_472# _136_ 0.003419f
C17583 trimb[2] net43 0.011999f
C17584 _216_/a_67_603# net36 0.028132f
C17585 _074_ _014_ 0.001557f
C17586 FILLER_0_13_100/a_124_375# net14 0.041373f
C17587 net68 FILLER_0_6_47/a_1020_375# 0.029857f
C17588 _254_/a_448_472# _072_ 0.002611f
C17589 output9/a_224_472# fanout76/a_36_160# 0.016067f
C17590 _064_ _445_/a_2665_112# 0.004701f
C17591 FILLER_0_10_78/a_484_472# vdd 0.004673f
C17592 FILLER_0_4_177/a_484_472# net22 0.006506f
C17593 _185_ _405_/a_67_603# 0.060789f
C17594 FILLER_0_4_107/a_1380_472# FILLER_0_2_111/a_1020_375# 0.001512f
C17595 _052_ vdd 0.264744f
C17596 vdd _202_/a_36_160# 0.06338f
C17597 net61 _419_/a_1000_472# 0.017712f
C17598 net60 _419_/a_1308_423# 0.029697f
C17599 mask\[5\] FILLER_0_18_177/a_36_472# 0.001063f
C17600 _111_ net36 0.102444f
C17601 FILLER_0_17_104/a_1468_375# vdd 0.022331f
C17602 net75 _083_ 0.055491f
C17603 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_36_472# 0.001723f
C17604 _013_ FILLER_0_18_37/a_1468_375# 0.017213f
C17605 _175_ cal_count\[1\] 0.203153f
C17606 net62 FILLER_0_14_263/a_124_375# 0.037111f
C17607 _161_ _060_ 0.042838f
C17608 _008_ result[4] 0.134001f
C17609 FILLER_0_3_204/a_124_375# net82 0.014222f
C17610 _025_ vdd 0.259346f
C17611 net54 _354_/a_257_69# 0.001135f
C17612 mask\[4\] _093_ 0.469687f
C17613 ctlp[1] FILLER_0_21_286/a_36_472# 0.014043f
C17614 output44/a_224_472# net40 0.006489f
C17615 _188_ _039_ 0.002071f
C17616 _112_ net1 0.001653f
C17617 _322_/a_124_24# _125_ 0.01165f
C17618 _105_ mask\[6\] 0.029716f
C17619 net78 net18 1.351707f
C17620 net31 FILLER_0_18_209/a_572_375# 0.001813f
C17621 _440_/a_796_472# _029_ 0.009261f
C17622 _269_/a_36_472# vdd 0.03432f
C17623 _174_ net74 0.00916f
C17624 _144_ FILLER_0_18_107/a_2364_375# 0.002388f
C17625 net28 _426_/a_448_472# 0.00154f
C17626 _086_ _163_ 0.413768f
C17627 _132_ vdd 0.960634f
C17628 net40 _167_ 0.020177f
C17629 net16 FILLER_0_8_37/a_572_375# 0.004285f
C17630 _015_ vss 0.090048f
C17631 FILLER_0_15_116/a_572_375# net36 0.007321f
C17632 FILLER_0_2_111/a_124_375# _157_ 0.028285f
C17633 net39 _445_/a_2248_156# 0.003571f
C17634 FILLER_0_5_72/a_932_472# trim_mask\[1\] 0.014619f
C17635 mask\[2\] FILLER_0_15_212/a_36_472# 0.001181f
C17636 _428_/a_36_151# FILLER_0_13_100/a_124_375# 0.023595f
C17637 FILLER_0_4_197/a_1468_375# net76 0.007667f
C17638 _038_ _120_ 0.00117f
C17639 _036_ _030_ 0.430683f
C17640 _247_/a_36_160# net22 0.048614f
C17641 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1468_375# 0.086742f
C17642 _065_ net15 0.065255f
C17643 _235_/a_67_603# net40 0.001273f
C17644 FILLER_0_4_99/a_124_375# net14 0.003714f
C17645 FILLER_0_20_193/a_124_375# vdd 0.009092f
C17646 _242_/a_36_160# _066_ 0.044262f
C17647 _142_ _334_/a_36_160# 0.009001f
C17648 _057_ _311_/a_1660_473# 0.004637f
C17649 _104_ FILLER_0_23_274/a_36_472# 0.001642f
C17650 output36/a_224_472# _417_/a_2665_112# 0.008243f
C17651 _189_/a_67_603# FILLER_0_12_220/a_1468_375# 0.029786f
C17652 _176_ _451_/a_448_472# 0.007191f
C17653 FILLER_0_17_72/a_484_472# _131_ 0.002672f
C17654 _081_ _001_ 0.012101f
C17655 FILLER_0_9_28/a_2276_472# vdd 0.003276f
C17656 FILLER_0_17_200/a_36_472# net63 0.005648f
C17657 trim[0] output41/a_224_472# 0.018464f
C17658 net16 _166_ 0.146913f
C17659 _079_ FILLER_0_5_206/a_124_375# 0.009128f
C17660 _420_/a_36_151# _009_ 0.018171f
C17661 mask\[7\] _436_/a_2248_156# 0.003615f
C17662 output24/a_224_472# net54 0.177947f
C17663 FILLER_0_17_226/a_124_375# fanout63/a_36_160# 0.008215f
C17664 FILLER_0_15_116/a_36_472# net70 0.051129f
C17665 FILLER_0_12_136/a_1468_375# vss 0.043987f
C17666 _116_ _161_ 0.008003f
C17667 FILLER_0_23_274/a_36_472# vss 0.002346f
C17668 FILLER_0_7_72/a_1020_375# net50 0.014749f
C17669 fanout61/a_36_113# vdd 0.108255f
C17670 net80 net57 0.002913f
C17671 net26 _423_/a_1204_472# 0.001069f
C17672 _002_ vdd 0.152662f
C17673 net64 FILLER_0_9_282/a_484_472# 0.005717f
C17674 mask\[4\] net54 0.009909f
C17675 result[7] FILLER_0_24_274/a_1020_375# 0.006125f
C17676 FILLER_0_5_212/a_124_375# net37 0.005414f
C17677 FILLER_0_7_195/a_36_472# vdd 0.04565f
C17678 FILLER_0_18_2/a_2812_375# net40 0.018463f
C17679 _032_ trim_mask\[4\] 0.010578f
C17680 FILLER_0_8_138/a_124_375# _125_ 0.001589f
C17681 FILLER_0_5_54/a_1468_375# vdd 0.014683f
C17682 FILLER_0_5_54/a_1020_375# vss 0.003196f
C17683 net23 _242_/a_36_160# 0.007466f
C17684 FILLER_0_17_72/a_1916_375# net36 0.015395f
C17685 net58 output27/a_224_472# 0.121438f
C17686 output11/a_224_472# net20 0.036556f
C17687 FILLER_0_7_104/a_572_375# _154_ 0.020664f
C17688 _442_/a_1204_472# vdd 0.001128f
C17689 net16 _185_ 0.086347f
C17690 net34 net21 0.036237f
C17691 trim_val\[4\] trim_mask\[4\] 0.152123f
C17692 _114_ _428_/a_2665_112# 0.002329f
C17693 result[9] output31/a_224_472# 0.082001f
C17694 _016_ net53 0.180698f
C17695 FILLER_0_16_241/a_124_375# vdd 0.035603f
C17696 net41 _446_/a_2560_156# 0.005695f
C17697 trim_val\[4\] net47 0.003977f
C17698 _126_ net14 0.238336f
C17699 _086_ _117_ 0.010287f
C17700 net31 net29 0.009564f
C17701 FILLER_0_18_177/a_1020_375# vdd 0.040478f
C17702 FILLER_0_4_177/a_36_472# vss 0.001806f
C17703 FILLER_0_4_177/a_484_472# vdd 0.010663f
C17704 _449_/a_796_472# _067_ 0.004874f
C17705 net79 FILLER_0_11_282/a_36_472# 0.004358f
C17706 _130_ _118_ 0.053869f
C17707 FILLER_0_12_20/a_36_472# vdd 0.068477f
C17708 FILLER_0_12_20/a_572_375# vss 0.054934f
C17709 _004_ _416_/a_2665_112# 0.002631f
C17710 FILLER_0_21_142/a_36_472# _210_/a_67_603# 0.001547f
C17711 _291_/a_36_160# _276_/a_36_160# 0.239422f
C17712 _450_/a_36_151# _039_ 0.018559f
C17713 _161_ _118_ 0.023939f
C17714 _095_ _406_/a_36_159# 0.131137f
C17715 net75 _425_/a_36_151# 0.02868f
C17716 _095_ FILLER_0_15_72/a_124_375# 0.001474f
C17717 net23 FILLER_0_16_154/a_36_472# 0.035678f
C17718 FILLER_0_7_72/a_1380_472# _028_ 0.001777f
C17719 _132_ _135_ 0.345161f
C17720 FILLER_0_7_162/a_36_472# _053_ 0.004888f
C17721 net20 _077_ 0.094476f
C17722 _432_/a_1000_472# _091_ 0.026097f
C17723 _412_/a_2665_112# vss 0.011887f
C17724 output42/a_224_472# output6/a_224_472# 0.292612f
C17725 state\[0\] vdd 0.120171f
C17726 _411_/a_2560_156# vdd 0.001315f
C17727 net17 FILLER_0_20_15/a_124_375# 0.005919f
C17728 net73 FILLER_0_18_107/a_2812_375# 0.018753f
C17729 _370_/a_124_24# vdd 0.018613f
C17730 _129_ _118_ 0.213736f
C17731 _352_/a_49_472# FILLER_0_22_128/a_36_472# 0.063744f
C17732 mask\[7\] FILLER_0_22_128/a_1020_375# 0.035799f
C17733 net72 FILLER_0_20_31/a_36_472# 0.002751f
C17734 _165_ vdd 0.168803f
C17735 FILLER_0_7_146/a_124_375# _059_ 0.029514f
C17736 _092_ _106_ 0.140596f
C17737 net70 _427_/a_36_151# 0.029237f
C17738 _439_/a_2560_156# vss 0.001309f
C17739 fanout53/a_36_160# _427_/a_2248_156# 0.027388f
C17740 _002_ FILLER_0_3_172/a_2812_375# 0.006403f
C17741 _350_/a_49_472# _208_/a_36_160# 0.078981f
C17742 _444_/a_2665_112# FILLER_0_8_37/a_484_472# 0.001167f
C17743 _412_/a_1000_472# net65 0.00929f
C17744 FILLER_0_15_150/a_124_375# vss 0.01957f
C17745 _428_/a_796_472# _043_ 0.007935f
C17746 FILLER_0_21_28/a_2276_472# _424_/a_36_151# 0.001723f
C17747 net29 result[2] 0.001786f
C17748 _292_/a_36_160# _204_/a_67_603# 0.003478f
C17749 _077_ net50 0.312283f
C17750 _247_/a_36_160# vdd 0.060423f
C17751 _115_ _322_/a_692_472# 0.00171f
C17752 _126_ _428_/a_36_151# 0.032026f
C17753 _096_ _116_ 0.020685f
C17754 net74 _032_ 0.208799f
C17755 _428_/a_448_472# _095_ 0.008804f
C17756 net58 _425_/a_2560_156# 0.004835f
C17757 _274_/a_36_68# _070_ 0.032424f
C17758 _443_/a_1000_472# _170_ 0.012879f
C17759 _061_ _090_ 0.00832f
C17760 _056_ _060_ 0.085489f
C17761 state\[2\] FILLER_0_13_142/a_1020_375# 0.007311f
C17762 net32 _420_/a_2665_112# 0.002753f
C17763 net53 FILLER_0_13_142/a_36_472# 0.059367f
C17764 net15 _440_/a_448_472# 0.036624f
C17765 net16 _407_/a_36_472# 0.027354f
C17766 net63 _434_/a_2248_156# 0.063346f
C17767 _091_ FILLER_0_13_212/a_124_375# 0.025558f
C17768 _053_ _059_ 0.042128f
C17769 net16 cal_count\[0\] 0.152321f
C17770 _105_ output21/a_224_472# 0.034631f
C17771 result[7] _421_/a_1456_156# 0.001009f
C17772 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_124_375# 0.026339f
C17773 FILLER_0_24_274/a_36_472# vdd 0.107635f
C17774 FILLER_0_24_274/a_1468_375# vss 0.060201f
C17775 mask\[4\] _343_/a_257_69# 0.001786f
C17776 _448_/a_2665_112# _170_ 0.002715f
C17777 _448_/a_1204_472# _037_ 0.008883f
C17778 _062_ _160_ 0.001024f
C17779 FILLER_0_12_28/a_124_375# vss 0.013117f
C17780 FILLER_0_12_28/a_36_472# vdd 0.095598f
C17781 vdd net40 1.984115f
C17782 _437_/a_2665_112# _436_/a_36_151# 0.001466f
C17783 _411_/a_1308_423# net75 0.028281f
C17784 FILLER_0_22_128/a_1916_375# vss 0.018094f
C17785 FILLER_0_22_128/a_2364_375# vdd 0.015888f
C17786 net71 FILLER_0_22_107/a_572_375# 0.006403f
C17787 _430_/a_36_151# fanout80/a_36_113# 0.018169f
C17788 _057_ _058_ 0.098076f
C17789 _284_/a_224_472# _094_ 0.001731f
C17790 _432_/a_448_472# _098_ 0.032293f
C17791 net58 _416_/a_36_151# 0.001558f
C17792 _086_ FILLER_0_11_142/a_36_472# 0.006774f
C17793 FILLER_0_3_78/a_124_375# _168_ 0.009374f
C17794 _315_/a_36_68# vss 0.02467f
C17795 net34 mask\[7\] 0.901671f
C17796 _126_ FILLER_0_11_109/a_36_472# 0.00136f
C17797 FILLER_0_18_171/a_124_375# vdd 0.021417f
C17798 FILLER_0_6_79/a_124_375# vdd 0.015119f
C17799 result[5] fanout78/a_36_113# 0.018989f
C17800 _084_ vss 0.082779f
C17801 _098_ FILLER_0_21_206/a_124_375# 0.001882f
C17802 _420_/a_36_151# FILLER_0_23_290/a_36_472# 0.001723f
C17803 FILLER_0_18_139/a_1380_472# net23 0.013087f
C17804 _086_ FILLER_0_7_104/a_1020_375# 0.00757f
C17805 net31 net60 0.012623f
C17806 net82 FILLER_0_3_172/a_572_375# 0.010972f
C17807 FILLER_0_10_78/a_932_472# net52 0.00207f
C17808 _095_ _281_/a_234_472# 0.001467f
C17809 FILLER_0_21_206/a_124_375# _205_/a_36_160# 0.03126f
C17810 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_124_375# 0.012267f
C17811 _136_ _018_ 0.002892f
C17812 net63 _202_/a_36_160# 0.004414f
C17813 FILLER_0_15_282/a_572_375# vss 0.058168f
C17814 FILLER_0_15_282/a_36_472# vdd 0.10628f
C17815 _120_ FILLER_0_9_72/a_932_472# 0.001709f
C17816 FILLER_0_17_38/a_572_375# vdd 0.01525f
C17817 _072_ _090_ 0.091468f
C17818 _114_ _070_ 0.507391f
C17819 net79 net22 0.042486f
C17820 _032_ _159_ 0.053405f
C17821 net34 net80 0.041846f
C17822 net7 net68 0.032489f
C17823 fanout66/a_36_113# _029_ 0.001684f
C17824 net65 _425_/a_2248_156# 0.003451f
C17825 _173_ _450_/a_3129_107# 0.00264f
C17826 _198_/a_67_603# vdd 0.015843f
C17827 net48 _305_/a_36_159# 0.059079f
C17828 _274_/a_3368_68# vss 0.001714f
C17829 _116_ _056_ 0.30649f
C17830 _415_/a_2665_112# FILLER_0_9_290/a_36_472# 0.007376f
C17831 net32 _419_/a_2560_156# 0.029586f
C17832 FILLER_0_17_72/a_3172_472# FILLER_0_17_104/a_36_472# 0.013277f
C17833 _414_/a_36_151# FILLER_0_6_177/a_572_375# 0.073306f
C17834 net36 net21 0.034415f
C17835 _077_ FILLER_0_10_78/a_124_375# 0.001886f
C17836 output21/a_224_472# output19/a_224_472# 0.007877f
C17837 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_124_375# 0.004426f
C17838 FILLER_0_6_47/a_3172_472# vss 0.014726f
C17839 _413_/a_1204_472# vdd 0.001027f
C17840 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_36_472# 0.001723f
C17841 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_572_375# 0.007947f
C17842 _035_ vss 0.105648f
C17843 _091_ net81 0.03653f
C17844 _008_ result[9] 0.048497f
C17845 net52 FILLER_0_6_47/a_2364_375# 0.002577f
C17846 _053_ FILLER_0_7_162/a_124_375# 0.007494f
C17847 _070_ FILLER_0_5_136/a_36_472# 0.029293f
C17848 net57 FILLER_0_13_100/a_36_472# 0.077963f
C17849 FILLER_0_3_142/a_124_375# _032_ 0.001153f
C17850 FILLER_0_0_266/a_36_472# rstn 0.006108f
C17851 net20 FILLER_0_6_231/a_572_375# 0.01215f
C17852 fanout71/a_36_113# _098_ 0.012725f
C17853 _339_/a_36_160# _140_ 0.025058f
C17854 FILLER_0_12_136/a_1468_375# _071_ 0.002023f
C17855 FILLER_0_12_2/a_124_375# clkc 0.003601f
C17856 net33 _108_ 0.001901f
C17857 FILLER_0_4_144/a_124_375# vss 0.017638f
C17858 FILLER_0_4_144/a_572_375# vdd -0.013698f
C17859 _412_/a_36_151# net76 0.001169f
C17860 net39 _034_ 0.004367f
C17861 _443_/a_448_472# _031_ 0.001143f
C17862 _032_ _442_/a_448_472# 0.001977f
C17863 _443_/a_796_472# net69 0.020234f
C17864 _056_ _118_ 0.028015f
C17865 result[9] result[8] 0.242998f
C17866 net19 net33 0.254336f
C17867 net54 FILLER_0_22_107/a_124_375# 0.003502f
C17868 _412_/a_1308_423# net81 0.006961f
C17869 _405_/a_67_603# net17 0.014714f
C17870 net63 FILLER_0_20_193/a_124_375# 0.075841f
C17871 _433_/a_36_151# _145_ 0.004437f
C17872 _116_ _068_ 0.011673f
C17873 FILLER_0_10_247/a_124_375# net64 0.001597f
C17874 _176_ _070_ 0.467961f
C17875 net34 _422_/a_2248_156# 0.005617f
C17876 net80 _340_/a_36_160# 0.004225f
C17877 FILLER_0_4_99/a_124_375# _153_ 0.030839f
C17878 _091_ _223_/a_36_160# 0.001976f
C17879 _236_/a_36_160# output39/a_224_472# 0.042231f
C17880 vss FILLER_0_5_148/a_484_472# 0.009015f
C17881 _077_ cal_itt\[3\] 0.009816f
C17882 _098_ FILLER_0_18_76/a_124_375# 0.001831f
C17883 net29 FILLER_0_16_255/a_124_375# 0.085055f
C17884 FILLER_0_2_101/a_124_375# _156_ 0.022015f
C17885 _112_ net76 0.011948f
C17886 mask\[5\] _146_ 0.051687f
C17887 net55 FILLER_0_17_72/a_1380_472# 0.021108f
C17888 FILLER_0_12_20/a_484_472# _450_/a_448_472# 0.04564f
C17889 FILLER_0_21_142/a_36_472# net54 0.02217f
C17890 _422_/a_36_151# _010_ 0.006787f
C17891 _019_ mask\[2\] 0.155325f
C17892 ctln[6] _442_/a_36_151# 0.007031f
C17893 FILLER_0_2_111/a_1380_472# vss 0.001679f
C17894 _260_/a_36_68# _080_ 0.001888f
C17895 FILLER_0_3_204/a_124_375# net21 0.010054f
C17896 FILLER_0_9_142/a_124_375# _122_ 0.004711f
C17897 net15 _394_/a_1936_472# 0.001592f
C17898 _256_/a_1612_497# _068_ 0.002759f
C17899 _445_/a_2248_156# net47 0.028909f
C17900 FILLER_0_13_65/a_36_472# FILLER_0_13_72/a_36_472# 0.002765f
C17901 _440_/a_2665_112# vss 0.008703f
C17902 _029_ _365_/a_692_472# 0.001426f
C17903 FILLER_0_18_2/a_3260_375# net41 0.042057f
C17904 _068_ _118_ 1.374452f
C17905 _070_ _124_ 0.114614f
C17906 net63 FILLER_0_18_177/a_1020_375# 0.007516f
C17907 trim_val\[2\] _381_/a_36_472# 0.005253f
C17908 net16 net55 0.035875f
C17909 cal_count\[2\] cal_count\[1\] 0.067712f
C17910 FILLER_0_10_78/a_1380_472# vss 0.002096f
C17911 _219_/a_36_160# vss 0.00157f
C17912 net60 _421_/a_36_151# 0.224039f
C17913 _136_ vss 0.947188f
C17914 FILLER_0_21_28/a_2724_472# _012_ 0.020109f
C17915 net55 _176_ 0.300149f
C17916 _128_ calibrate 0.039365f
C17917 FILLER_0_16_89/a_572_375# _131_ 0.012481f
C17918 net4 _080_ 0.076128f
C17919 _017_ FILLER_0_14_107/a_484_472# 0.004583f
C17920 FILLER_0_16_73/a_124_375# vdd 0.008987f
C17921 net70 FILLER_0_14_107/a_1380_472# 0.003355f
C17922 net79 vdd 1.283563f
C17923 FILLER_0_12_136/a_1020_375# _126_ 0.012732f
C17924 net79 _192_/a_67_603# 0.017688f
C17925 _077_ _039_ 0.104126f
C17926 net62 vss 1.17087f
C17927 FILLER_0_1_266/a_36_472# net8 0.0138f
C17928 FILLER_0_21_142/a_124_375# _098_ 0.006558f
C17929 output32/a_224_472# net60 0.191561f
C17930 _303_/a_36_472# vdd 0.015964f
C17931 _386_/a_848_380# net22 0.00429f
C17932 _438_/a_1000_472# vss 0.001536f
C17933 net66 _440_/a_36_151# 0.041433f
C17934 FILLER_0_13_142/a_572_375# vdd 0.017472f
C17935 ctlp[1] _419_/a_2665_112# 0.009197f
C17936 _345_/a_36_160# net71 0.002396f
C17937 net73 FILLER_0_19_111/a_36_472# 0.001412f
C17938 FILLER_0_13_142/a_124_375# vss 0.009543f
C17939 _161_ _228_/a_36_68# 0.055774f
C17940 _374_/a_36_68# _062_ 0.004248f
C17941 output21/a_224_472# mask\[6\] 0.013037f
C17942 net34 output34/a_224_472# 0.031833f
C17943 _128_ net21 0.03068f
C17944 cal clk 0.033015f
C17945 FILLER_0_5_109/a_572_375# _160_ 0.004207f
C17946 fanout82/a_36_113# net2 0.008681f
C17947 FILLER_0_12_124/a_36_472# _332_/a_36_472# 0.004546f
C17948 _199_/a_36_160# _046_ 0.017122f
C17949 FILLER_0_4_177/a_484_472# FILLER_0_2_177/a_572_375# 0.001512f
C17950 mask\[5\] FILLER_0_19_171/a_1380_472# 0.007596f
C17951 _141_ net80 0.077957f
C17952 FILLER_0_5_72/a_1468_375# net49 0.001276f
C17953 _390_/a_244_472# _067_ 0.004031f
C17954 FILLER_0_10_78/a_1380_472# _308_/a_124_24# 0.037778f
C17955 net44 FILLER_0_15_2/a_572_375# 0.041552f
C17956 FILLER_0_15_2/a_36_472# vss 0.002136f
C17957 net80 net36 0.036729f
C17958 net16 net17 0.034209f
C17959 _004_ result[1] 0.005653f
C17960 _327_/a_36_472# _114_ 0.019746f
C17961 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_124_375# 0.012552f
C17962 _125_ _120_ 0.006198f
C17963 net68 FILLER_0_5_54/a_36_472# 0.012107f
C17964 net16 trim_val\[1\] 0.164715f
C17965 net15 FILLER_0_7_59/a_484_472# 0.015199f
C17966 net15 _453_/a_36_151# 0.009841f
C17967 FILLER_0_16_255/a_36_472# _102_ 0.004641f
C17968 FILLER_0_21_125/a_36_472# _140_ 0.101284f
C17969 _447_/a_2248_156# net69 0.001126f
C17970 en clk 0.067072f
C17971 _028_ FILLER_0_5_72/a_1380_472# 0.002164f
C17972 FILLER_0_9_28/a_3172_472# vss 0.001977f
C17973 _133_ _062_ 1.210949f
C17974 _072_ FILLER_0_7_233/a_36_472# 0.00241f
C17975 ctlp[7] _436_/a_36_151# 0.002655f
C17976 output43/a_224_472# vss -0.005182f
C17977 _417_/a_1204_472# _006_ 0.014354f
C17978 FILLER_0_7_104/a_484_472# _131_ 0.00432f
C17979 net36 mask\[1\] 0.28584f
C17980 output27/a_224_472# calibrate 0.010614f
C17981 _440_/a_2665_112# FILLER_0_5_88/a_124_375# 0.02132f
C17982 _429_/a_2665_112# vss 0.012165f
C17983 _367_/a_36_68# _154_ 0.028801f
C17984 FILLER_0_17_56/a_572_375# vss 0.05884f
C17985 FILLER_0_17_56/a_36_472# vdd 0.040007f
C17986 _442_/a_36_151# _371_/a_36_113# 0.001089f
C17987 _072_ _163_ 0.016226f
C17988 _148_ _436_/a_36_151# 0.032004f
C17989 _000_ _253_/a_244_68# 0.001243f
C17990 input1/a_36_113# clk 0.001121f
C17991 _014_ FILLER_0_7_233/a_36_472# 0.002089f
C17992 _119_ net74 0.02813f
C17993 _422_/a_36_151# _299_/a_36_472# 0.004432f
C17994 _069_ _247_/a_36_160# 0.046764f
C17995 FILLER_0_15_150/a_124_375# _095_ 0.003939f
C17996 cal_count\[1\] _043_ 0.002223f
C17997 _316_/a_692_472# vdd 0.001634f
C17998 net20 _009_ 0.026064f
C17999 net79 _416_/a_1204_472# 0.006493f
C18000 output46/a_224_472# trimb[3] 0.050924f
C18001 net55 FILLER_0_18_76/a_124_375# 0.001706f
C18002 FILLER_0_9_28/a_484_472# net51 0.001023f
C18003 FILLER_0_19_55/a_124_375# FILLER_0_19_47/a_572_375# 0.012001f
C18004 net62 _416_/a_2248_156# 0.043158f
C18005 FILLER_0_9_223/a_484_472# _128_ 0.005152f
C18006 vdd FILLER_0_13_290/a_124_375# 0.031436f
C18007 _424_/a_36_151# FILLER_0_18_37/a_572_375# 0.002807f
C18008 _430_/a_36_151# _139_ 0.012035f
C18009 _412_/a_796_472# net2 0.00566f
C18010 FILLER_0_3_172/a_124_375# net59 0.001045f
C18011 _413_/a_36_151# output12/a_224_472# 0.006251f
C18012 _061_ _117_ 0.046662f
C18013 net53 vss 0.426484f
C18014 net26 _424_/a_1000_472# 0.003207f
C18015 _453_/a_448_472# _042_ 0.053209f
C18016 _453_/a_36_151# net51 0.012537f
C18017 _415_/a_36_151# net27 0.019856f
C18018 net62 _195_/a_67_603# 0.002422f
C18019 FILLER_0_3_54/a_36_472# _160_ 0.00702f
C18020 _058_ FILLER_0_10_94/a_124_375# 0.001597f
C18021 _311_/a_66_473# _117_ 0.001055f
C18022 FILLER_0_20_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001543f
C18023 _070_ _267_/a_36_472# 0.002617f
C18024 _386_/a_124_24# vss 0.009702f
C18025 _386_/a_848_380# vdd 0.054849f
C18026 trim[4] _054_ 0.005511f
C18027 FILLER_0_19_125/a_124_375# _145_ 0.006777f
C18028 _260_/a_36_68# vss 0.030324f
C18029 _412_/a_2248_156# vss 0.005692f
C18030 _113_ _060_ 0.01991f
C18031 FILLER_0_19_171/a_572_375# vdd 0.022516f
C18032 FILLER_0_20_87/a_36_472# net14 0.001471f
C18033 _085_ _121_ 0.027373f
C18034 FILLER_0_22_86/a_36_472# net71 0.005766f
C18035 net15 FILLER_0_13_72/a_572_375# 0.003021f
C18036 net15 fanout51/a_36_113# 0.001562f
C18037 _423_/a_2248_156# FILLER_0_23_60/a_124_375# 0.001901f
C18038 fanout51/a_36_113# FILLER_0_11_78/a_36_472# 0.193759f
C18039 FILLER_0_18_2/a_36_472# net44 0.011079f
C18040 _451_/a_1353_112# net14 0.041814f
C18041 fanout68/a_36_113# net66 0.042828f
C18042 FILLER_0_5_72/a_484_472# _164_ 0.003769f
C18043 output42/a_224_472# FILLER_0_9_28/a_124_375# 0.003337f
C18044 FILLER_0_10_107/a_484_472# vss 0.00298f
C18045 _321_/a_358_69# _121_ 0.00135f
C18046 net27 FILLER_0_10_256/a_36_472# 0.008331f
C18047 fanout60/a_36_160# net18 0.004124f
C18048 mask\[1\] FILLER_0_15_228/a_36_472# 0.02055f
C18049 _088_ FILLER_0_4_213/a_124_375# 0.016013f
C18050 net14 _160_ 0.034023f
C18051 _452_/a_1040_527# vdd 0.004153f
C18052 net27 net64 1.364577f
C18053 _242_/a_36_160# FILLER_0_5_148/a_572_375# 0.00805f
C18054 _144_ _208_/a_36_160# 0.00717f
C18055 _143_ FILLER_0_16_154/a_1468_375# 0.002033f
C18056 net55 _041_ 0.972122f
C18057 trim[4] vss 0.033925f
C18058 net4 vss 0.774455f
C18059 FILLER_0_18_177/a_2724_472# net21 0.048803f
C18060 mask\[3\] FILLER_0_16_154/a_932_472# 0.002604f
C18061 FILLER_0_9_28/a_1828_472# net68 0.048468f
C18062 state\[0\] FILLER_0_9_223/a_572_375# 0.079258f
C18063 FILLER_0_17_200/a_484_472# vss 0.003134f
C18064 _164_ _160_ 1.863027f
C18065 _425_/a_2560_156# calibrate 0.010842f
C18066 _376_/a_36_160# FILLER_0_5_88/a_36_472# 0.001448f
C18067 net15 net69 0.034091f
C18068 _003_ _087_ 0.054908f
C18069 FILLER_0_4_197/a_124_375# _088_ 0.024641f
C18070 _406_/a_36_159# _185_ 0.001573f
C18071 _012_ FILLER_0_21_60/a_36_472# 0.017483f
C18072 _440_/a_448_472# net47 0.016997f
C18073 FILLER_0_24_96/a_124_375# ctlp[7] 0.004486f
C18074 output12/a_224_472# FILLER_0_1_192/a_124_375# 0.032639f
C18075 FILLER_0_14_107/a_572_375# vdd 0.021509f
C18076 FILLER_0_14_107/a_124_375# vss 0.002674f
C18077 _119_ _154_ 0.01697f
C18078 _305_/a_36_159# net37 0.015682f
C18079 FILLER_0_9_72/a_36_472# vss 0.0392f
C18080 FILLER_0_9_72/a_484_472# vdd 0.005654f
C18081 _056_ _228_/a_36_68# 0.043669f
C18082 _093_ _013_ 0.064462f
C18083 _420_/a_36_151# FILLER_0_23_282/a_572_375# 0.059049f
C18084 _389_/a_36_148# FILLER_0_10_94/a_124_375# 0.004673f
C18085 fanout61/a_36_113# net77 0.052643f
C18086 net18 rstn 0.015842f
C18087 _010_ _419_/a_36_151# 0.002099f
C18088 _116_ _113_ 0.179616f
C18089 result[5] _103_ 0.425479f
C18090 _412_/a_2665_112# output37/a_224_472# 0.002025f
C18091 _289_/a_36_472# vdd 0.006886f
C18092 _095_ FILLER_0_14_123/a_36_472# 0.014431f
C18093 FILLER_0_5_72/a_1380_472# net47 0.003924f
C18094 FILLER_0_19_187/a_36_472# _434_/a_36_151# 0.002398f
C18095 fanout51/a_36_113# net51 0.013081f
C18096 _453_/a_2248_156# vss 0.031525f
C18097 _453_/a_2665_112# vdd 0.005481f
C18098 _127_ FILLER_0_11_142/a_484_472# 0.001177f
C18099 fanout68/a_36_113# FILLER_0_3_54/a_124_375# 0.015816f
C18100 _311_/a_1920_473# vdd 0.007492f
C18101 ctln[3] net75 0.066513f
C18102 net17 _041_ 0.002779f
C18103 _015_ _426_/a_2248_156# 0.021465f
C18104 _430_/a_2248_156# vdd 0.008989f
C18105 input2/a_36_113# en 0.002108f
C18106 FILLER_0_19_55/a_124_375# net55 0.005311f
C18107 FILLER_0_19_47/a_36_472# _424_/a_448_472# 0.004782f
C18108 _256_/a_2960_68# _076_ 0.001292f
C18109 _087_ net37 0.23484f
C18110 _000_ FILLER_0_3_221/a_932_472# 0.008308f
C18111 net47 _034_ 0.052602f
C18112 net79 _283_/a_36_472# 0.010249f
C18113 net54 FILLER_0_22_86/a_1468_375# 0.001597f
C18114 mask\[4\] _144_ 0.268823f
C18115 _136_ FILLER_0_16_154/a_1020_375# 0.004387f
C18116 _098_ _437_/a_2560_156# 0.001174f
C18117 fanout49/a_36_160# _030_ 0.017759f
C18118 _091_ FILLER_0_18_171/a_36_472# 0.00395f
C18119 trimb[1] FILLER_0_20_2/a_572_375# 0.003431f
C18120 _091_ FILLER_0_18_177/a_36_472# 0.012695f
C18121 net32 _421_/a_2248_156# 0.038586f
C18122 net81 FILLER_0_15_212/a_932_472# 0.003953f
C18123 _118_ _113_ 0.005092f
C18124 vss _433_/a_1000_472# 0.002059f
C18125 mask\[0\] _429_/a_1204_472# 0.005396f
C18126 _448_/a_2560_156# net59 0.007516f
C18127 _096_ FILLER_0_14_181/a_36_472# 0.028078f
C18128 fanout69/a_36_113# FILLER_0_2_111/a_1468_375# 0.015816f
C18129 net80 FILLER_0_20_177/a_124_375# 0.001198f
C18130 _027_ _438_/a_1000_472# 0.010911f
C18131 _111_ FILLER_0_18_76/a_124_375# 0.002494f
C18132 input1/a_36_113# input2/a_36_113# 0.029417f
C18133 FILLER_0_3_172/a_1916_375# net22 0.00941f
C18134 FILLER_0_18_53/a_572_375# vss 0.057185f
C18135 FILLER_0_18_53/a_36_472# vdd 0.089087f
C18136 _029_ trim_mask\[1\] 1.002118f
C18137 _094_ _418_/a_796_472# 0.005889f
C18138 FILLER_0_17_133/a_124_375# vdd 0.010519f
C18139 input5/a_36_113# vdd 0.026855f
C18140 fanout76/a_36_160# net4 0.002206f
C18141 FILLER_0_8_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001597f
C18142 net54 _211_/a_36_160# 0.001244f
C18143 _132_ _140_ 0.019255f
C18144 _052_ _424_/a_2665_112# 0.003027f
C18145 FILLER_0_16_57/a_36_472# _131_ 0.00864f
C18146 _121_ _062_ 0.001616f
C18147 FILLER_0_12_124/a_36_472# FILLER_0_11_124/a_36_472# 0.05841f
C18148 net34 FILLER_0_22_177/a_1468_375# 0.006974f
C18149 ctln[1] rstn 0.62944f
C18150 _162_ FILLER_0_5_172/a_36_472# 0.001501f
C18151 fanout55/a_36_160# FILLER_0_13_80/a_124_375# 0.00805f
C18152 net55 FILLER_0_17_64/a_124_375# 0.020021f
C18153 _086_ net37 0.039329f
C18154 _115_ FILLER_0_10_94/a_124_375# 0.010311f
C18155 FILLER_0_15_142/a_36_472# _427_/a_36_151# 0.001723f
C18156 _445_/a_1308_423# net40 0.046345f
C18157 FILLER_0_5_128/a_572_375# _152_ 0.00813f
C18158 _053_ FILLER_0_6_47/a_572_375# 0.008213f
C18159 FILLER_0_7_104/a_932_472# _133_ 0.019721f
C18160 _131_ FILLER_0_11_109/a_124_375# 0.001048f
C18161 _017_ FILLER_0_13_100/a_124_375# 0.001274f
C18162 _093_ FILLER_0_17_72/a_3260_375# 0.011936f
C18163 FILLER_0_10_28/a_124_375# vdd 0.039012f
C18164 net16 _408_/a_1336_472# 0.022364f
C18165 _008_ _418_/a_1000_472# 0.01006f
C18166 net58 _426_/a_36_151# 0.002612f
C18167 FILLER_0_9_105/a_124_375# vdd 0.029831f
C18168 _398_/a_36_113# _278_/a_36_160# 0.001636f
C18169 FILLER_0_13_142/a_1020_375# _043_ 0.005672f
C18170 FILLER_0_20_177/a_1468_375# vdd 0.016422f
C18171 _114_ FILLER_0_10_94/a_36_472# 0.08191f
C18172 _069_ net79 0.045808f
C18173 net64 FILLER_0_14_235/a_36_472# 0.067888f
C18174 _136_ _095_ 0.043768f
C18175 net35 _423_/a_2248_156# 0.003899f
C18176 mask\[8\] _423_/a_2665_112# 0.004281f
C18177 FILLER_0_21_125/a_572_375# _098_ 0.006462f
C18178 net16 _447_/a_1308_423# 0.001178f
C18179 ctln[9] _447_/a_36_151# 0.010503f
C18180 output48/a_224_472# en 0.003074f
C18181 net15 _013_ 0.152142f
C18182 _398_/a_36_113# _178_ 0.004282f
C18183 _141_ FILLER_0_16_154/a_36_472# 0.00126f
C18184 net36 FILLER_0_15_212/a_124_375# 0.004391f
C18185 _130_ net74 0.001655f
C18186 net56 net23 0.930833f
C18187 net36 _099_ 0.325141f
C18188 _104_ _422_/a_36_151# 0.032235f
C18189 _035_ output41/a_224_472# 0.002168f
C18190 net70 FILLER_0_16_115/a_124_375# 0.025173f
C18191 FILLER_0_9_223/a_124_375# _055_ 0.014525f
C18192 net68 _120_ 0.001304f
C18193 _429_/a_36_151# FILLER_0_15_212/a_484_472# 0.001723f
C18194 FILLER_0_20_15/a_1468_375# vdd 0.009742f
C18195 output44/a_224_472# FILLER_0_19_28/a_36_472# 0.023414f
C18196 _053_ net52 0.042556f
C18197 FILLER_0_4_107/a_124_375# _156_ 0.00268f
C18198 _321_/a_2590_472# _118_ 0.002396f
C18199 _422_/a_36_151# vss 0.014056f
C18200 _422_/a_448_472# vdd 0.032865f
C18201 _168_ vdd 0.083621f
C18202 _155_ trim_mask\[1\] 0.006536f
C18203 FILLER_0_9_28/a_36_472# net42 0.038355f
C18204 _441_/a_1308_423# vss 0.016854f
C18205 _129_ net74 0.476969f
C18206 _093_ net71 0.133323f
C18207 _031_ _369_/a_692_472# 0.00359f
C18208 _067_ FILLER_0_13_72/a_124_375# 0.001782f
C18209 output23/a_224_472# FILLER_0_22_128/a_1468_375# 0.00242f
C18210 vss _047_ 0.070755f
C18211 net55 _424_/a_1308_423# 0.00168f
C18212 net34 output18/a_224_472# 0.17524f
C18213 _064_ _446_/a_2248_156# 0.04774f
C18214 net52 FILLER_0_5_54/a_1380_472# 0.00179f
C18215 trim_val\[1\] FILLER_0_6_47/a_124_375# 0.002577f
C18216 _004_ net81 0.993594f
C18217 _058_ FILLER_0_9_105/a_484_472# 0.00148f
C18218 _114_ net21 0.022033f
C18219 FILLER_0_16_241/a_124_375# _282_/a_36_160# 0.005398f
C18220 _293_/a_36_472# vdd 0.087136f
C18221 FILLER_0_14_81/a_124_375# cal_count\[1\] 0.070473f
C18222 _132_ _451_/a_36_151# 0.007777f
C18223 en_co_clk _067_ 0.272082f
C18224 _005_ _416_/a_2665_112# 0.014205f
C18225 mask\[4\] FILLER_0_19_155/a_36_472# 0.047448f
C18226 _258_/a_36_160# net59 0.003167f
C18227 _176_ FILLER_0_10_94/a_36_472# 0.009089f
C18228 FILLER_0_19_55/a_124_375# _216_/a_67_603# 0.003017f
C18229 FILLER_0_18_139/a_572_375# FILLER_0_19_142/a_124_375# 0.026339f
C18230 _432_/a_1308_423# _137_ 0.002078f
C18231 fanout70/a_36_113# _095_ 0.003087f
C18232 _441_/a_1204_472# _168_ 0.009437f
C18233 _273_/a_36_68# _060_ 0.010339f
C18234 _058_ vss 0.19427f
C18235 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_124_375# 0.016748f
C18236 _131_ FILLER_0_17_104/a_124_375# 0.006681f
C18237 FILLER_0_6_239/a_124_375# vdd 0.031271f
C18238 ctlp[1] _421_/a_1204_472# 0.003759f
C18239 _021_ vss 0.142648f
C18240 net48 _001_ 0.006122f
C18241 FILLER_0_17_142/a_36_472# _137_ 0.003953f
C18242 fanout77/a_36_113# vss 0.004099f
C18243 _105_ net31 0.054065f
C18244 FILLER_0_20_31/a_124_375# vss 0.049142f
C18245 FILLER_0_20_31/a_36_472# vdd 0.097195f
C18246 cal_itt\[2\] net58 0.003431f
C18247 _444_/a_2248_156# FILLER_0_6_37/a_124_375# 0.001101f
C18248 FILLER_0_3_172/a_1916_375# vdd -0.010166f
C18249 _412_/a_448_472# vdd 0.011f
C18250 _359_/a_36_488# _070_ 0.028563f
C18251 FILLER_0_15_290/a_36_472# output30/a_224_472# 0.001711f
C18252 _108_ vdd 0.298249f
C18253 net16 FILLER_0_16_37/a_124_375# 0.033245f
C18254 net16 _444_/a_1308_423# 0.002172f
C18255 _170_ _066_ 0.189122f
C18256 net75 _416_/a_2665_112# 0.001785f
C18257 FILLER_0_4_123/a_36_472# trim_mask\[4\] 0.003692f
C18258 net19 vdd 2.167778f
C18259 net28 net79 0.116857f
C18260 net16 FILLER_0_8_24/a_572_375# 0.002225f
C18261 net19 _192_/a_67_603# 0.003106f
C18262 _423_/a_36_151# FILLER_0_23_44/a_932_472# 0.001723f
C18263 FILLER_0_18_2/a_2812_375# FILLER_0_19_28/a_36_472# 0.001684f
C18264 _232_/a_67_603# net47 0.014888f
C18265 state\[2\] _043_ 0.028842f
C18266 _287_/a_36_472# _094_ 0.029751f
C18267 _098_ FILLER_0_15_212/a_1380_472# 0.009972f
C18268 FILLER_0_4_197/a_1380_472# net22 0.012286f
C18269 FILLER_0_4_123/a_36_472# net47 0.012399f
C18270 _072_ net48 0.037795f
C18271 vss _416_/a_1308_423# 0.001962f
C18272 FILLER_0_12_136/a_124_375# _130_ 0.010514f
C18273 _422_/a_796_472# _108_ 0.007356f
C18274 _141_ FILLER_0_18_139/a_1380_472# 0.016119f
C18275 trim_mask\[1\] _163_ 0.166315f
C18276 _153_ _160_ 0.304792f
C18277 mask\[8\] _026_ 0.001638f
C18278 _126_ _017_ 0.071134f
C18279 net54 net71 0.536043f
C18280 net65 FILLER_0_2_171/a_124_375# 0.023202f
C18281 _188_ vdd 0.022839f
C18282 _281_/a_234_472# _098_ 0.003724f
C18283 _175_ _043_ 0.001037f
C18284 FILLER_0_21_206/a_124_375# net21 0.035287f
C18285 FILLER_0_4_197/a_36_472# _002_ 0.006574f
C18286 _258_/a_36_160# _122_ 0.00102f
C18287 net76 net1 0.059026f
C18288 FILLER_0_11_64/a_36_472# _120_ 0.011673f
C18289 FILLER_0_11_64/a_36_472# _038_ 0.001822f
C18290 net13 _387_/a_36_113# 0.00189f
C18291 net23 _170_ 0.107532f
C18292 net53 _095_ 0.431214f
C18293 cal_itt\[2\] _082_ 0.032565f
C18294 _098_ _434_/a_1204_472# 0.006257f
C18295 _258_/a_36_160# FILLER_0_7_233/a_124_375# 0.001633f
C18296 cal_itt\[2\] net82 0.663246f
C18297 FILLER_0_13_65/a_36_472# net15 0.036527f
C18298 net48 _014_ 0.276733f
C18299 FILLER_0_14_91/a_36_472# _136_ 0.008573f
C18300 _053_ _359_/a_1044_488# 0.001474f
C18301 _389_/a_36_148# vss 0.001935f
C18302 net79 FILLER_0_12_236/a_572_375# 0.010684f
C18303 _434_/a_448_472# _023_ 0.03093f
C18304 ctln[1] _411_/a_2248_156# 0.013381f
C18305 FILLER_0_4_49/a_572_375# net66 0.074393f
C18306 net55 _406_/a_36_159# 0.001219f
C18307 net16 trim_mask\[2\] 0.002527f
C18308 _140_ FILLER_0_22_128/a_2364_375# 0.003037f
C18309 net52 FILLER_0_3_78/a_36_472# 0.034084f
C18310 output28/a_224_472# FILLER_0_11_282/a_36_472# 0.008834f
C18311 net52 FILLER_0_2_127/a_36_472# 0.001964f
C18312 _435_/a_2248_156# mask\[6\] 0.001778f
C18313 ctlp[3] _422_/a_2560_156# 0.001006f
C18314 _076_ net23 0.105196f
C18315 _430_/a_2248_156# net63 0.051057f
C18316 net49 FILLER_0_3_78/a_36_472# 0.059367f
C18317 _030_ FILLER_0_3_78/a_484_472# 0.007736f
C18318 FILLER_0_17_161/a_124_375# vdd 0.014253f
C18319 _431_/a_448_472# _093_ 0.002095f
C18320 _068_ net47 0.001491f
C18321 _055_ _311_/a_1212_473# 0.004259f
C18322 trimb[3] net17 0.005798f
C18323 _009_ FILLER_0_23_290/a_36_472# 0.002345f
C18324 net57 _131_ 0.030577f
C18325 _119_ _313_/a_255_603# 0.001151f
C18326 net41 _217_/a_36_160# 0.004517f
C18327 FILLER_0_4_123/a_36_472# net74 0.001578f
C18328 _074_ FILLER_0_5_172/a_36_472# 0.016713f
C18329 net19 net9 0.342451f
C18330 FILLER_0_3_172/a_2724_472# net65 0.001777f
C18331 FILLER_0_7_72/a_36_472# net52 0.014911f
C18332 _070_ _246_/a_36_68# 0.056186f
C18333 net79 net77 0.431572f
C18334 _095_ FILLER_0_14_107/a_124_375# 0.01418f
C18335 _420_/a_36_151# vdd 0.137919f
C18336 FILLER_0_20_107/a_36_472# _438_/a_2665_112# 0.035266f
C18337 _406_/a_36_159# net17 0.053547f
C18338 net58 FILLER_0_8_247/a_1380_472# 0.0597f
C18339 _115_ FILLER_0_9_105/a_484_472# 0.004075f
C18340 net4 FILLER_0_12_220/a_124_375# 0.016485f
C18341 _443_/a_2560_156# vss 0.002467f
C18342 FILLER_0_19_47/a_124_375# _052_ 0.019401f
C18343 _228_/a_36_68# _113_ 0.021898f
C18344 FILLER_0_9_223/a_36_472# _068_ 0.076678f
C18345 _430_/a_2248_156# _069_ 0.042876f
C18346 FILLER_0_16_107/a_36_472# vdd 0.110244f
C18347 _122_ _062_ 0.190871f
C18348 _115_ vss 0.372063f
C18349 FILLER_0_19_28/a_572_375# vss 0.002775f
C18350 FILLER_0_19_28/a_36_472# vdd 0.052986f
C18351 _446_/a_1000_472# net66 0.006158f
C18352 vdd _450_/a_36_151# 0.08588f
C18353 FILLER_0_4_197/a_1380_472# vdd 0.00581f
C18354 cal_count\[3\] _373_/a_632_68# 0.004529f
C18355 trim_mask\[1\] FILLER_0_4_91/a_36_472# 0.26171f
C18356 _423_/a_2248_156# vdd 0.013707f
C18357 trimb[0] vss 0.097724f
C18358 FILLER_0_16_57/a_932_472# net55 0.00179f
C18359 FILLER_0_14_181/a_36_472# _138_ 0.002748f
C18360 _062_ _227_/a_36_160# 0.015411f
C18361 FILLER_0_8_127/a_36_472# _070_ 0.005078f
C18362 net63 FILLER_0_20_177/a_1468_375# 0.018435f
C18363 trim_mask\[4\] net69 0.185121f
C18364 net57 net56 0.054294f
C18365 _022_ _145_ 0.199016f
C18366 _081_ _066_ 0.061358f
C18367 net60 FILLER_0_17_282/a_36_472# 0.009978f
C18368 _432_/a_448_472# net80 0.045963f
C18369 _002_ _413_/a_1308_423# 0.002178f
C18370 _214_/a_36_160# FILLER_0_23_88/a_36_472# 0.006647f
C18371 mask\[4\] FILLER_0_19_187/a_484_472# 0.004669f
C18372 FILLER_0_4_123/a_36_472# _159_ 0.004956f
C18373 FILLER_0_14_91/a_36_472# net53 0.005849f
C18374 output9/a_224_472# net58 0.050634f
C18375 _115_ _308_/a_124_24# 0.039354f
C18376 ctln[7] ctln[8] 0.004643f
C18377 FILLER_0_4_49/a_124_375# _164_ 0.017213f
C18378 _440_/a_36_151# FILLER_0_6_47/a_2276_472# 0.001512f
C18379 _345_/a_36_160# FILLER_0_19_111/a_484_472# 0.007907f
C18380 FILLER_0_8_138/a_36_472# _058_ 0.005325f
C18381 FILLER_0_17_72/a_2724_472# vdd 0.007064f
C18382 FILLER_0_17_72/a_2276_472# vss -0.001288f
C18383 _181_ _402_/a_2172_497# 0.001555f
C18384 _412_/a_1308_423# net59 0.00291f
C18385 FILLER_0_22_86/a_572_375# net14 0.009573f
C18386 _419_/a_36_151# vss -0.00139f
C18387 _419_/a_448_472# vdd 0.022174f
C18388 _238_/a_67_603# trim_mask\[3\] 0.028437f
C18389 net35 net24 0.01339f
C18390 _402_/a_56_567# _452_/a_36_151# 0.001915f
C18391 _412_/a_2248_156# output37/a_224_472# 0.001141f
C18392 net43 net40 0.018193f
C18393 FILLER_0_16_89/a_36_472# _040_ 0.015634f
C18394 ctln[6] _031_ 0.004486f
C18395 FILLER_0_4_107/a_932_472# _158_ 0.029116f
C18396 FILLER_0_4_123/a_36_472# _154_ 0.001043f
C18397 _081_ net23 0.081773f
C18398 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_36_472# 0.026657f
C18399 _132_ FILLER_0_17_104/a_1380_472# 0.02114f
C18400 FILLER_0_6_239/a_36_472# net76 0.011803f
C18401 _431_/a_1000_472# net73 0.035816f
C18402 _427_/a_2560_156# vss 0.003576f
C18403 trim_mask\[4\] _152_ 0.224909f
C18404 net19 _420_/a_1308_423# 0.010051f
C18405 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_484_472# 0.013276f
C18406 _016_ FILLER_0_12_124/a_124_375# 0.007335f
C18407 FILLER_0_13_142/a_1468_375# _225_/a_36_160# 0.027706f
C18408 FILLER_0_15_150/a_124_375# fanout53/a_36_160# 0.004079f
C18409 _372_/a_2590_472# _076_ 0.002268f
C18410 ctln[9] vss 0.167242f
C18411 _269_/a_36_472# _083_ 0.015096f
C18412 net74 FILLER_0_13_72/a_572_375# 0.012891f
C18413 _412_/a_796_472# cal_itt\[1\] 0.004226f
C18414 _152_ net47 0.242864f
C18415 _257_/a_36_472# vss 0.023401f
C18416 _413_/a_448_472# output12/a_224_472# 0.001495f
C18417 trim_val\[4\] FILLER_0_3_172/a_124_375# 0.002076f
C18418 FILLER_0_1_204/a_36_472# net59 0.067975f
C18419 net60 _010_ 0.108311f
C18420 _072_ FILLER_0_12_220/a_36_472# 0.01861f
C18421 FILLER_0_22_128/a_2364_375# FILLER_0_21_150/a_36_472# 0.001543f
C18422 _415_/a_1000_472# net27 0.017938f
C18423 net4 FILLER_0_12_236/a_36_472# 0.016315f
C18424 output9/a_224_472# net82 0.003636f
C18425 ctln[7] FILLER_0_1_98/a_124_375# 0.004533f
C18426 FILLER_0_6_90/a_36_472# _163_ 0.016147f
C18427 _186_ vdd 0.074983f
C18428 _035_ _166_ 0.034749f
C18429 net61 ctlp[2] 0.022612f
C18430 net66 _029_ 0.056971f
C18431 _369_/a_692_472# _157_ 0.0025f
C18432 FILLER_0_4_152/a_124_375# vss 0.019426f
C18433 FILLER_0_4_49/a_36_472# net47 0.002964f
C18434 _075_ _257_/a_36_472# 0.005709f
C18435 _091_ net64 0.079488f
C18436 mask\[7\] _435_/a_1308_423# 0.028235f
C18437 _394_/a_728_93# cal_count\[1\] 0.057049f
C18438 _411_/a_2665_112# net10 0.007912f
C18439 net74 net69 0.143604f
C18440 FILLER_0_8_263/a_124_375# FILLER_0_8_247/a_1468_375# 0.012001f
C18441 net22 FILLER_0_18_209/a_36_472# 0.018061f
C18442 _091_ FILLER_0_19_171/a_1380_472# 0.001044f
C18443 _149_ vss 0.005314f
C18444 FILLER_0_2_171/a_36_472# net59 0.066486f
C18445 net23 FILLER_0_22_128/a_1828_472# 0.003857f
C18446 FILLER_0_3_2/a_124_375# _446_/a_36_151# 0.023595f
C18447 _213_/a_67_603# _051_ 0.015959f
C18448 _426_/a_36_151# calibrate 0.004525f
C18449 FILLER_0_18_139/a_1020_375# vdd 0.001285f
C18450 FILLER_0_18_139/a_572_375# vss 0.009977f
C18451 mask\[0\] FILLER_0_14_235/a_484_472# 0.004688f
C18452 _335_/a_49_472# _098_ 0.001047f
C18453 result[1] _005_ 0.001478f
C18454 result[2] FILLER_0_13_290/a_36_472# 0.016496f
C18455 _077_ net22 0.049592f
C18456 net57 _170_ 0.057355f
C18457 _408_/a_56_524# _067_ 0.003678f
C18458 FILLER_0_14_181/a_36_472# _113_ 0.004214f
C18459 net78 _420_/a_2665_112# 0.039469f
C18460 FILLER_0_9_72/a_1468_375# _439_/a_36_151# 0.005577f
C18461 _093_ FILLER_0_18_107/a_3260_375# 0.008393f
C18462 FILLER_0_5_148/a_36_472# _160_ 0.001025f
C18463 _077_ FILLER_0_9_72/a_1380_472# 0.006408f
C18464 FILLER_0_15_282/a_36_472# output30/a_224_472# 0.001711f
C18465 FILLER_0_15_282/a_124_375# net30 0.00123f
C18466 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_484_472# 0.001723f
C18467 FILLER_0_12_28/a_124_375# cal_count\[0\] 0.001414f
C18468 FILLER_0_0_130/a_36_472# vss 0.00351f
C18469 FILLER_0_10_256/a_124_375# _426_/a_36_151# 0.001597f
C18470 FILLER_0_18_177/a_2812_375# _202_/a_36_160# 0.026361f
C18471 _308_/a_848_380# FILLER_0_10_94/a_484_472# 0.019491f
C18472 _114_ _171_ 0.203692f
C18473 cal_count\[3\] _055_ 0.039546f
C18474 net57 _074_ 0.026184f
C18475 _414_/a_1000_472# _074_ 0.00222f
C18476 FILLER_0_14_81/a_124_375# _175_ 0.005719f
C18477 _064_ net39 0.558387f
C18478 net74 _152_ 1.007413f
C18479 net67 _221_/a_36_160# 0.008581f
C18480 FILLER_0_1_204/a_124_375# net11 0.01048f
C18481 FILLER_0_7_72/a_1020_375# vdd 0.004039f
C18482 input3/a_36_113# cal_count\[2\] 0.00555f
C18483 net41 output40/a_224_472# 0.018977f
C18484 _155_ FILLER_0_7_104/a_484_472# 0.003068f
C18485 result[0] fanout65/a_36_113# 0.001816f
C18486 net57 _076_ 0.028356f
C18487 _435_/a_1204_472# vdd 0.013805f
C18488 net38 _444_/a_1000_472# 0.027886f
C18489 FILLER_0_7_72/a_2276_472# _077_ 0.00475f
C18490 _136_ _451_/a_448_472# 0.047841f
C18491 FILLER_0_9_28/a_2276_472# _053_ 0.002243f
C18492 net32 _297_/a_36_472# 0.001843f
C18493 FILLER_0_17_72/a_572_375# FILLER_0_15_72/a_484_472# 0.001512f
C18494 FILLER_0_13_212/a_36_472# _429_/a_1308_423# 0.009119f
C18495 _013_ _012_ 0.003113f
C18496 net38 FILLER_0_8_24/a_484_472# 0.001223f
C18497 _103_ _418_/a_2665_112# 0.0066f
C18498 net69 _159_ 0.010086f
C18499 _063_ _167_ 0.002201f
C18500 _443_/a_448_472# net23 0.038188f
C18501 FILLER_0_8_2/a_124_375# net40 0.002839f
C18502 output28/a_224_472# vdd 0.044767f
C18503 FILLER_0_18_76/a_36_472# vss 0.007456f
C18504 FILLER_0_4_197/a_932_472# net59 0.003599f
C18505 ctln[1] cal_itt\[0\] 0.003349f
C18506 _134_ FILLER_0_9_105/a_484_472# 0.011499f
C18507 _126_ cal_count\[3\] 0.418508f
C18508 _020_ vss 0.008954f
C18509 _372_/a_2034_472# _152_ 0.00171f
C18510 cal fanout58/a_36_160# 0.047586f
C18511 _086_ _127_ 0.042698f
C18512 FILLER_0_10_37/a_36_472# _453_/a_36_151# 0.003462f
C18513 _431_/a_36_151# net73 0.015086f
C18514 _099_ FILLER_0_14_235/a_484_472# 0.00281f
C18515 FILLER_0_4_107/a_36_472# trim_mask\[3\] 0.00152f
C18516 _134_ vss 0.088213f
C18517 _137_ FILLER_0_17_104/a_1468_375# 0.002679f
C18518 net7 _446_/a_36_151# 0.001237f
C18519 _176_ _171_ 0.049997f
C18520 net69 _154_ 0.05211f
C18521 FILLER_0_20_193/a_36_472# FILLER_0_18_177/a_1916_375# 0.0027f
C18522 net54 FILLER_0_18_107/a_3260_375# 0.001619f
C18523 _042_ net51 0.026776f
C18524 FILLER_0_6_90/a_484_472# FILLER_0_4_91/a_572_375# 0.00108f
C18525 FILLER_0_11_64/a_124_375# vdd 0.045435f
C18526 output11/a_224_472# vdd 0.01016f
C18527 net32 result[8] 0.024881f
C18528 FILLER_0_18_2/a_2276_472# net38 0.002313f
C18529 net57 en_co_clk 0.195533f
C18530 _159_ _152_ 0.035925f
C18531 _345_/a_36_160# net73 0.032139f
C18532 _121_ FILLER_0_8_156/a_124_375# 0.033427f
C18533 _086_ FILLER_0_11_135/a_36_472# 0.004074f
C18534 _132_ _137_ 0.023462f
C18535 _442_/a_448_472# net69 0.004308f
C18536 _445_/a_36_151# vdd 0.052935f
C18537 FILLER_0_21_28/a_3260_375# vss 0.054959f
C18538 FILLER_0_21_28/a_36_472# vdd 0.090954f
C18539 FILLER_0_18_209/a_572_375# vss 0.007545f
C18540 FILLER_0_18_209/a_36_472# vdd 0.089327f
C18541 fanout58/a_36_160# en 0.00568f
C18542 _320_/a_1792_472# _043_ 0.002235f
C18543 net52 FILLER_0_2_93/a_572_375# 0.007787f
C18544 output43/a_224_472# output46/a_224_472# 0.292611f
C18545 _077_ FILLER_0_9_105/a_36_472# 0.003177f
C18546 _126_ _320_/a_672_472# 0.003662f
C18547 _053_ _165_ 0.123461f
C18548 _356_/a_36_472# net14 0.001801f
C18549 cal_itt\[2\] output8/a_224_472# 0.05561f
C18550 net16 _179_ 0.007397f
C18551 _077_ vdd 1.61568f
C18552 FILLER_0_4_107/a_1380_472# trim_mask\[4\] 0.011766f
C18553 _074_ cal_itt\[0\] 0.076802f
C18554 net36 _451_/a_1040_527# 0.00974f
C18555 _427_/a_448_472# net23 0.014853f
C18556 FILLER_0_3_142/a_36_472# _081_ 0.001386f
C18557 net76 FILLER_0_5_198/a_124_375# 0.006974f
C18558 FILLER_0_12_50/a_124_375# _120_ 0.002753f
C18559 FILLER_0_4_107/a_1380_472# net47 0.008874f
C18560 net79 output30/a_224_472# 0.078502f
C18561 net81 _429_/a_2248_156# 0.017036f
C18562 fanout53/a_36_160# _136_ 0.001471f
C18563 _070_ _315_/a_36_68# 0.031892f
C18564 net38 output39/a_224_472# 0.036027f
C18565 mask\[4\] mask\[5\] 0.176881f
C18566 net28 net19 0.115252f
C18567 FILLER_0_20_107/a_124_375# vss 0.002749f
C18568 FILLER_0_20_107/a_36_472# vdd 0.117841f
C18569 FILLER_0_12_20/a_572_375# net17 0.041149f
C18570 net23 _145_ 0.035734f
C18571 trim_mask\[2\] _030_ 1.467465f
C18572 _412_/a_2665_112# net58 0.006815f
C18573 net76 FILLER_0_2_177/a_124_375# 0.00439f
C18574 ctln[0] output40/a_224_472# 0.017541f
C18575 _428_/a_2665_112# FILLER_0_13_142/a_124_375# 0.003325f
C18576 result[1] _416_/a_448_472# 0.008784f
C18577 _009_ FILLER_0_23_282/a_572_375# 0.016879f
C18578 net24 vdd 0.223761f
C18579 net14 FILLER_0_10_94/a_484_472# 0.020589f
C18580 _412_/a_1204_472# net1 0.019647f
C18581 _131_ net36 0.068899f
C18582 net57 _081_ 0.023513f
C18583 net53 _451_/a_448_472# 0.026909f
C18584 net70 _451_/a_836_156# 0.006451f
C18585 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_124_375# 0.026339f
C18586 _414_/a_1000_472# _081_ 0.006091f
C18587 _408_/a_244_524# net47 0.001066f
C18588 _425_/a_2248_156# net37 0.01491f
C18589 result[7] _102_ 0.010818f
C18590 mask\[5\] FILLER_0_19_187/a_124_375# 0.007169f
C18591 FILLER_0_18_2/a_2364_375# net55 0.005899f
C18592 _012_ net71 0.004946f
C18593 _136_ _098_ 0.049635f
C18594 _132_ FILLER_0_15_116/a_124_375# 0.047331f
C18595 FILLER_0_7_72/a_2276_472# net50 0.030391f
C18596 result[9] ctlp[1] 0.074012f
C18597 result[0] FILLER_0_9_290/a_124_375# 0.030628f
C18598 ctln[7] net14 0.197449f
C18599 FILLER_0_10_78/a_572_375# _115_ 0.004573f
C18600 net61 _418_/a_448_472# 0.001253f
C18601 _053_ FILLER_0_6_79/a_124_375# 0.003818f
C18602 _119_ _319_/a_672_472# 0.00488f
C18603 FILLER_0_18_2/a_1020_375# net38 0.047331f
C18604 net29 vss 0.259409f
C18605 output39/a_224_472# net66 0.009679f
C18606 _314_/a_224_472# net23 0.001238f
C18607 _426_/a_796_472# vdd 0.007178f
C18608 _028_ FILLER_0_6_90/a_124_375# 0.012573f
C18609 _098_ _438_/a_1000_472# 0.001492f
C18610 _255_/a_224_552# _057_ 0.024333f
C18611 FILLER_0_8_247/a_1380_472# calibrate 0.008605f
C18612 FILLER_0_12_220/a_484_472# _060_ 0.003379f
C18613 _141_ net56 0.012364f
C18614 FILLER_0_16_89/a_932_472# vdd 0.002218f
C18615 FILLER_0_16_89/a_484_472# vss -0.001894f
C18616 net7 _447_/a_36_151# 0.002494f
C18617 fanout49/a_36_160# _440_/a_2665_112# 0.00631f
C18618 _256_/a_36_68# _128_ 0.001702f
C18619 _413_/a_36_151# vdd 0.130213f
C18620 _063_ vdd 0.201806f
C18621 _427_/a_1308_423# net74 0.005627f
C18622 FILLER_0_2_93/a_484_472# net14 0.019214f
C18623 net72 FILLER_0_17_38/a_484_472# 0.00547f
C18624 net55 FILLER_0_17_38/a_124_375# 0.003236f
C18625 _091_ _097_ 0.036863f
C18626 _323_/a_36_113# _060_ 0.002584f
C18627 FILLER_0_13_228/a_36_472# net79 0.006824f
C18628 net36 _196_/a_36_160# 0.024527f
C18629 _131_ FILLER_0_10_107/a_572_375# 0.007252f
C18630 net56 net36 0.772486f
C18631 FILLER_0_13_65/a_36_472# net74 0.014937f
C18632 FILLER_0_17_142/a_484_472# vss 0.030872f
C18633 mask\[4\] FILLER_0_19_195/a_36_472# 0.004669f
C18634 net17 FILLER_0_12_28/a_124_375# 0.009108f
C18635 FILLER_0_18_2/a_2364_375# net17 0.048345f
C18636 FILLER_0_6_47/a_1468_375# vdd -0.014642f
C18637 _225_/a_36_160# vdd 0.058272f
C18638 FILLER_0_14_107/a_572_375# _451_/a_36_151# 0.02627f
C18639 net58 _084_ 0.141836f
C18640 cal_count\[3\] state\[1\] 0.236393f
C18641 _427_/a_2560_156# _095_ 0.009888f
C18642 FILLER_0_2_93/a_36_472# trim_mask\[3\] 0.003417f
C18643 _068_ FILLER_0_5_148/a_124_375# 0.003986f
C18644 _093_ FILLER_0_19_111/a_484_472# 0.001009f
C18645 net18 _193_/a_36_160# 0.114176f
C18646 mask\[9\] FILLER_0_19_111/a_36_472# 0.285112f
C18647 net20 vdd 2.14128f
C18648 FILLER_0_15_142/a_484_472# vss 0.029611f
C18649 net61 mask\[7\] 0.071542f
C18650 _066_ _163_ 0.006401f
C18651 _430_/a_36_151# _093_ 0.00184f
C18652 FILLER_0_17_38/a_572_375# _182_ 0.035561f
C18653 vdd FILLER_0_12_196/a_36_472# 0.019648f
C18654 vss FILLER_0_12_196/a_124_375# 0.042104f
C18655 cal net18 0.123815f
C18656 _432_/a_2665_112# _139_ 0.004089f
C18657 fanout53/a_36_160# net53 0.014917f
C18658 _428_/a_2665_112# net53 0.002379f
C18659 trim_val\[2\] _164_ 0.005847f
C18660 cal_count\[1\] _180_ 0.300952f
C18661 _050_ _436_/a_796_472# 0.007055f
C18662 FILLER_0_19_195/a_124_375# FILLER_0_19_187/a_572_375# 0.012001f
C18663 _081_ cal_itt\[0\] 0.036569f
C18664 _077_ fanout67/a_36_160# 0.017322f
C18665 FILLER_0_1_266/a_572_375# rstn 0.00328f
C18666 net27 FILLER_0_9_282/a_124_375# 0.003572f
C18667 _444_/a_1204_472# net47 0.007847f
C18668 _016_ FILLER_0_12_136/a_484_472# 0.001516f
C18669 vss FILLER_0_6_231/a_124_375# 0.00353f
C18670 vdd FILLER_0_6_231/a_572_375# 0.018694f
C18671 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_484_472# 0.013277f
C18672 net50 vdd 0.661261f
C18673 _091_ mask\[2\] 2.252217f
C18674 _415_/a_2248_156# result[1] 0.010922f
C18675 net38 _245_/a_672_472# 0.006341f
C18676 result[9] FILLER_0_24_274/a_124_375# 0.008195f
C18677 net57 _443_/a_448_472# 0.001956f
C18678 _068_ _313_/a_255_603# 0.001149f
C18679 net67 _450_/a_448_472# 0.068692f
C18680 _136_ _070_ 0.010577f
C18681 _019_ _138_ 0.003734f
C18682 _144_ net71 0.039862f
C18683 FILLER_0_18_107/a_2724_472# vdd 0.004677f
C18684 net23 _163_ 0.034799f
C18685 _084_ _082_ 0.044645f
C18686 _432_/a_36_151# _136_ 0.004543f
C18687 _382_/a_224_472# vdd 0.001663f
C18688 _136_ FILLER_0_15_180/a_124_375# 0.002442f
C18689 _429_/a_2665_112# _098_ 0.003225f
C18690 FILLER_0_15_150/a_36_472# vss 0.00975f
C18691 net82 _084_ 0.020793f
C18692 _394_/a_728_93# _175_ 0.010801f
C18693 _424_/a_1204_472# vdd 0.001573f
C18694 _413_/a_36_151# FILLER_0_3_172/a_2812_375# 0.059049f
C18695 FILLER_0_1_192/a_124_375# vdd 0.017212f
C18696 _143_ FILLER_0_18_171/a_36_472# 0.005167f
C18697 en net18 0.32189f
C18698 net65 cal_itt\[0\] 0.07564f
C18699 mask\[4\] FILLER_0_18_177/a_2276_472# 0.016876f
C18700 net81 _005_ 0.003646f
C18701 _104_ net60 0.063407f
C18702 net50 _441_/a_1204_472# 0.006986f
C18703 net52 _441_/a_2665_112# 0.004975f
C18704 _035_ net17 0.021052f
C18705 FILLER_0_4_107/a_484_472# _153_ 0.026082f
C18706 FILLER_0_4_107/a_1380_472# _154_ 0.005297f
C18707 FILLER_0_9_28/a_572_375# net41 0.025588f
C18708 mask\[3\] FILLER_0_18_177/a_1380_472# 0.005654f
C18709 comp cal_count\[2\] 0.015029f
C18710 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_572_375# 0.086635f
C18711 _132_ _040_ 0.023821f
C18712 cal_itt\[3\] net22 0.134309f
C18713 FILLER_0_12_124/a_124_375# vss 0.012672f
C18714 net60 vss 0.382678f
C18715 net54 FILLER_0_19_111/a_484_472# 0.00105f
C18716 net29 _195_/a_67_603# 0.048817f
C18717 _432_/a_2560_156# net80 0.01523f
C18718 net18 _417_/a_2248_156# 0.001601f
C18719 _417_/a_2665_112# net30 0.015638f
C18720 FILLER_0_16_57/a_1020_375# net15 0.048731f
C18721 net33 FILLER_0_22_128/a_3260_375# 0.001178f
C18722 output36/a_224_472# FILLER_0_15_282/a_36_472# 0.008834f
C18723 _064_ net47 0.110169f
C18724 _441_/a_2665_112# net49 0.062459f
C18725 ctln[1] cal 0.123834f
C18726 FILLER_0_21_206/a_36_472# _204_/a_67_603# 0.003123f
C18727 FILLER_0_5_172/a_36_472# _163_ 0.006934f
C18728 FILLER_0_8_239/a_36_472# vss 0.003115f
C18729 comp input3/a_36_113# 0.022213f
C18730 FILLER_0_19_134/a_124_375# _145_ 0.023167f
C18731 input1/a_36_113# net18 0.004922f
C18732 _074_ FILLER_0_6_177/a_572_375# 0.012642f
C18733 _428_/a_448_472# FILLER_0_14_107/a_932_472# 0.007f
C18734 FILLER_0_5_72/a_572_375# vdd -0.00211f
C18735 FILLER_0_5_72/a_124_375# vss 0.041166f
C18736 mask\[3\] FILLER_0_17_218/a_124_375# 0.016168f
C18737 net69 FILLER_0_2_111/a_36_472# 0.010759f
C18738 _031_ FILLER_0_2_111/a_1020_375# 0.016661f
C18739 net14 FILLER_0_4_91/a_572_375# 0.047331f
C18740 _272_/a_36_472# _079_ 0.0237f
C18741 FILLER_0_7_72/a_1916_375# FILLER_0_6_90/a_36_472# 0.001684f
C18742 net61 _422_/a_2248_156# 0.027973f
C18743 FILLER_0_18_177/a_1828_472# FILLER_0_19_187/a_572_375# 0.001684f
C18744 FILLER_0_5_128/a_484_472# net47 0.009309f
C18745 _420_/a_36_151# net77 0.023469f
C18746 _098_ FILLER_0_19_171/a_124_375# 0.040575f
C18747 net75 net81 0.420021f
C18748 net32 _109_ 0.038411f
C18749 _122_ FILLER_0_8_156/a_124_375# 0.032617f
C18750 _441_/a_36_151# _440_/a_36_151# 0.003983f
C18751 net38 net6 0.071232f
C18752 _267_/a_672_472# _071_ 0.00255f
C18753 net67 _043_ 0.003726f
C18754 FILLER_0_12_136/a_1468_375# FILLER_0_13_142/a_932_472# 0.001684f
C18755 net41 _452_/a_448_472# 0.052165f
C18756 fanout81/a_36_160# vdd 0.095319f
C18757 net42 net47 0.237866f
C18758 _273_/a_36_68# FILLER_0_9_223/a_36_472# 0.015795f
C18759 output46/a_224_472# FILLER_0_20_15/a_1020_375# 0.001274f
C18760 _446_/a_448_472# net40 0.05302f
C18761 _426_/a_36_151# FILLER_0_8_247/a_124_375# 0.059049f
C18762 _012_ FILLER_0_23_44/a_932_472# 0.001572f
C18763 FILLER_0_17_200/a_124_375# _093_ 0.00419f
C18764 _430_/a_36_151# _337_/a_49_472# 0.023882f
C18765 FILLER_0_16_107/a_572_375# _131_ 0.015859f
C18766 _227_/a_36_160# FILLER_0_8_156/a_124_375# 0.005398f
C18767 _008_ mask\[3\] 0.799138f
C18768 _375_/a_960_497# vdd 0.004471f
C18769 _081_ FILLER_0_5_148/a_572_375# 0.01425f
C18770 _421_/a_448_472# net19 0.058446f
C18771 output12/a_224_472# net22 0.002662f
C18772 _415_/a_36_151# _004_ 0.013592f
C18773 net20 _430_/a_2665_112# 0.005397f
C18774 net15 FILLER_0_15_59/a_36_472# 0.00464f
C18775 _324_/a_224_472# _070_ 0.00142f
C18776 FILLER_0_10_78/a_124_375# vdd -0.011193f
C18777 net36 FILLER_0_15_180/a_36_472# 0.007275f
C18778 _328_/a_36_113# vdd 0.136098f
C18779 _445_/a_2665_112# trim_mask\[1\] 0.00183f
C18780 trim[4] FILLER_0_8_2/a_36_472# 0.019134f
C18781 _384_/a_224_472# _160_ 0.00324f
C18782 FILLER_0_22_177/a_484_472# _435_/a_36_151# 0.001723f
C18783 _091_ FILLER_0_15_212/a_572_375# 0.022582f
C18784 net51 _450_/a_2449_156# 0.008215f
C18785 net68 net67 0.147318f
C18786 net34 FILLER_0_22_128/a_1828_472# 0.005158f
C18787 FILLER_0_21_125/a_484_472# vss 0.002399f
C18788 FILLER_0_15_72/a_484_472# vdd 0.002283f
C18789 FILLER_0_15_72/a_36_472# vss 0.038986f
C18790 _004_ FILLER_0_10_256/a_36_472# 0.00402f
C18791 ctln[1] input1/a_36_113# 0.004419f
C18792 FILLER_0_4_197/a_1468_375# vss 0.057762f
C18793 _004_ net64 0.001495f
C18794 _015_ calibrate 0.105287f
C18795 _427_/a_2665_112# state\[1\] 0.021573f
C18796 _419_/a_448_472# net77 0.007659f
C18797 _067_ net6 0.015232f
C18798 output34/a_224_472# net61 0.008309f
C18799 _411_/a_2665_112# net8 0.036782f
C18800 net46 FILLER_0_21_28/a_484_472# 0.001795f
C18801 net47 FILLER_0_4_91/a_484_472# 0.007531f
C18802 FILLER_0_5_128/a_484_472# net74 0.025425f
C18803 comp _043_ 0.003867f
C18804 FILLER_0_10_256/a_124_375# _015_ 0.001151f
C18805 FILLER_0_3_2/a_124_375# vss 0.007235f
C18806 FILLER_0_3_2/a_36_472# vdd 0.106665f
C18807 output27/a_224_472# net18 0.058296f
C18808 result[6] fanout61/a_36_113# 0.003917f
C18809 net73 _093_ 0.350073f
C18810 net50 fanout67/a_36_160# 0.007195f
C18811 _035_ _446_/a_1308_423# 0.002639f
C18812 ctln[8] trim_val\[3\] 0.007f
C18813 _067_ _172_ 0.010195f
C18814 net55 FILLER_0_17_56/a_572_375# 0.020564f
C18815 cal_itt\[3\] vdd 0.571239f
C18816 _070_ FILLER_0_10_107/a_484_472# 0.007421f
C18817 cal_itt\[2\] _413_/a_2665_112# 0.003007f
C18818 FILLER_0_23_88/a_124_375# net14 0.002894f
C18819 fanout81/a_36_160# net9 0.002274f
C18820 output28/a_224_472# net28 0.048681f
C18821 _056_ _311_/a_254_473# 0.005937f
C18822 _428_/a_1000_472# vdd 0.005345f
C18823 _098_ _433_/a_1000_472# 0.0184f
C18824 FILLER_0_16_255/a_36_472# net19 0.001273f
C18825 _009_ vdd 0.693198f
C18826 net4 _070_ 0.169392f
C18827 _086_ _116_ 1.316798f
C18828 FILLER_0_12_136/a_1380_472# state\[2\] 0.005779f
C18829 _437_/a_1308_423# net14 0.085815f
C18830 _068_ FILLER_0_9_142/a_124_375# 0.008226f
C18831 _076_ FILLER_0_9_142/a_36_472# 0.038562f
C18832 _411_/a_1204_472# ctln[3] 0.00185f
C18833 trim_mask\[4\] _369_/a_36_68# 0.00407f
C18834 _394_/a_1336_472# vdd 0.003226f
C18835 _086_ _321_/a_3126_472# 0.001522f
C18836 _290_/a_224_472# result[5] 0.001638f
C18837 output43/a_224_472# net17 0.083607f
C18838 FILLER_0_11_142/a_36_472# net23 0.002015f
C18839 _412_/a_1204_472# net76 0.020975f
C18840 _081_ FILLER_0_6_177/a_572_375# 0.007285f
C18841 _059_ _160_ 0.037235f
C18842 _422_/a_796_472# _009_ 0.001178f
C18843 output14/a_224_472# _442_/a_2665_112# 0.009771f
C18844 net80 _434_/a_1204_472# 0.003997f
C18845 vdd _039_ 0.219985f
C18846 FILLER_0_18_107/a_932_472# FILLER_0_16_115/a_124_375# 0.001512f
C18847 fanout68/a_36_113# _441_/a_36_151# 0.138322f
C18848 FILLER_0_1_98/a_124_375# trim_val\[3\] 0.001628f
C18849 result[4] result[5] 0.090472f
C18850 _132_ FILLER_0_14_107/a_484_472# 0.005391f
C18851 _112_ _316_/a_1084_68# 0.005773f
C18852 _328_/a_36_113# _135_ 0.005635f
C18853 net20 net63 0.045207f
C18854 _128_ _076_ 0.04562f
C18855 net15 _449_/a_2248_156# 0.001705f
C18856 output12/a_224_472# vdd 0.106635f
C18857 FILLER_0_20_177/a_1020_375# _098_ 0.013949f
C18858 FILLER_0_15_212/a_1380_472# mask\[1\] 0.041503f
C18859 net7 vss 0.117948f
C18860 net55 _452_/a_1353_112# 0.030679f
C18861 _413_/a_36_151# FILLER_0_2_177/a_572_375# 0.073306f
C18862 FILLER_0_5_164/a_124_375# _386_/a_848_380# 0.014613f
C18863 _068_ _311_/a_254_473# 0.002606f
C18864 _086_ _118_ 0.166544f
C18865 _077_ _449_/a_36_151# 0.002475f
C18866 net25 FILLER_0_23_88/a_36_472# 0.192699f
C18867 net76 FILLER_0_1_192/a_36_472# 0.003817f
C18868 _334_/a_36_160# FILLER_0_17_104/a_1468_375# 0.027706f
C18869 net54 _436_/a_1000_472# 0.002051f
C18870 _427_/a_36_151# FILLER_0_14_123/a_124_375# 0.023595f
C18871 _065_ _447_/a_2560_156# 0.012523f
C18872 FILLER_0_4_177/a_124_375# _163_ 0.004052f
C18873 net57 _163_ 0.759175f
C18874 _173_ _042_ 0.002294f
C18875 _412_/a_2248_156# net58 0.010702f
C18876 _424_/a_2665_112# _423_/a_2248_156# 0.001314f
C18877 trim_mask\[1\] FILLER_0_6_47/a_932_472# 0.007542f
C18878 _434_/a_2560_156# vdd 0.002922f
C18879 _434_/a_2665_112# vss 0.00127f
C18880 _067_ _450_/a_2225_156# 0.002584f
C18881 cal_itt\[3\] _251_/a_1130_472# 0.001099f
C18882 FILLER_0_15_116/a_572_375# _136_ 0.001706f
C18883 _132_ _334_/a_36_160# 0.026495f
C18884 net82 _316_/a_848_380# 0.087022f
C18885 ctln[4] FILLER_0_1_204/a_36_472# 0.006408f
C18886 FILLER_0_21_133/a_124_375# _433_/a_36_151# 0.059049f
C18887 fanout61/a_36_113# _418_/a_36_151# 0.001442f
C18888 _322_/a_124_24# vss 0.003731f
C18889 _322_/a_848_380# vdd 0.067623f
C18890 net18 _416_/a_36_151# 0.027435f
C18891 FILLER_0_4_99/a_36_472# _030_ 0.002699f
C18892 mask\[5\] FILLER_0_20_169/a_124_375# 0.011078f
C18893 FILLER_0_16_73/a_484_472# _176_ 0.010681f
C18894 _231_/a_652_68# _062_ 0.001555f
C18895 _057_ state\[2\] 0.054838f
C18896 _098_ _047_ 0.062495f
C18897 output13/a_224_472# net13 0.058196f
C18898 FILLER_0_2_101/a_124_375# vss 0.04897f
C18899 FILLER_0_2_101/a_36_472# vdd 0.099518f
C18900 vss FILLER_0_8_156/a_484_472# 0.004078f
C18901 net58 net4 0.858616f
C18902 FILLER_0_15_142/a_484_472# _095_ 0.001509f
C18903 _188_ FILLER_0_12_50/a_36_472# 0.006464f
C18904 net35 FILLER_0_22_128/a_3260_375# 0.012732f
C18905 net17 _452_/a_1353_112# 0.038603f
C18906 output32/a_224_472# _419_/a_1308_423# 0.005111f
C18907 _205_/a_36_160# _047_ 0.013528f
C18908 _207_/a_67_603# _146_ 0.026192f
C18909 _119_ _062_ 0.080398f
C18910 net55 _453_/a_2248_156# 0.001546f
C18911 net35 net33 1.594925f
C18912 _132_ FILLER_0_16_107/a_124_375# 0.003315f
C18913 _250_/a_36_68# state\[2\] 0.038165f
C18914 FILLER_0_16_107/a_36_472# _451_/a_36_151# 0.059367f
C18915 net68 FILLER_0_6_47/a_1916_375# 0.00799f
C18916 mask\[5\] _201_/a_67_603# 0.001222f
C18917 trimb[0] output46/a_224_472# 0.048191f
C18918 _265_/a_244_68# vdd 0.022571f
C18919 net15 _439_/a_1000_472# 0.001798f
C18920 _021_ _098_ 0.014179f
C18921 cal net65 0.023638f
C18922 FILLER_0_18_100/a_124_375# _438_/a_2665_112# 0.010688f
C18923 _411_/a_1000_472# net75 0.03227f
C18924 net60 _419_/a_1000_472# 0.028992f
C18925 net61 _419_/a_2248_156# 0.022159f
C18926 net54 FILLER_0_22_128/a_124_375# 0.032013f
C18927 FILLER_0_17_104/a_484_472# vdd 0.020339f
C18928 FILLER_0_17_104/a_36_472# vss 0.002744f
C18929 _444_/a_448_472# net40 0.055844f
C18930 FILLER_0_17_72/a_1916_375# _136_ 0.009573f
C18931 _326_/a_36_160# _062_ 0.007797f
C18932 fanout70/a_36_113# FILLER_0_15_116/a_572_375# 0.003553f
C18933 FILLER_0_8_24/a_124_375# net40 0.002431f
C18934 _450_/a_1697_156# net6 0.00236f
C18935 _345_/a_36_160# _433_/a_36_151# 0.015565f
C18936 _153_ FILLER_0_4_91/a_572_375# 0.001735f
C18937 mask\[3\] _093_ 2.443356f
C18938 FILLER_0_15_150/a_36_472# _095_ 0.001526f
C18939 FILLER_0_7_195/a_124_375# _072_ 0.012244f
C18940 ctlp[5] _435_/a_36_151# 0.003815f
C18941 FILLER_0_3_204/a_124_375# net65 0.003831f
C18942 net4 _082_ 0.004529f
C18943 _230_/a_244_68# _056_ 0.001844f
C18944 net82 net4 1.982825f
C18945 _300_/a_224_472# _011_ 0.007508f
C18946 fanout50/a_36_160# trim_val\[3\] 0.017252f
C18947 net55 FILLER_0_18_53/a_572_375# 0.015895f
C18948 net16 FILLER_0_8_37/a_484_472# 0.004272f
C18949 FILLER_0_8_138/a_124_375# vss 0.00629f
C18950 _267_/a_224_472# state\[1\] 0.001937f
C18951 net41 cal_count\[3\] 0.028902f
C18952 net75 _317_/a_36_113# 0.030797f
C18953 net65 en 0.001469f
C18954 _114_ _131_ 0.036548f
C18955 FILLER_0_23_290/a_36_472# vdd 0.089567f
C18956 FILLER_0_23_290/a_124_375# vss 0.033011f
C18957 FILLER_0_15_116/a_484_472# net36 0.009319f
C18958 net39 _445_/a_2560_156# 0.003401f
C18959 _132_ FILLER_0_18_107/a_1468_375# 0.089207f
C18960 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_124_375# 0.026339f
C18961 _096_ _320_/a_36_472# 0.052438f
C18962 _065_ ctln[8] 0.193903f
C18963 _092_ output18/a_224_472# 0.002205f
C18964 _050_ FILLER_0_22_107/a_572_375# 0.001825f
C18965 FILLER_0_20_193/a_572_375# vss 0.005887f
C18966 FILLER_0_20_193/a_36_472# vdd 0.091886f
C18967 output31/a_224_472# _094_ 0.004668f
C18968 FILLER_0_17_72/a_1380_472# _131_ 0.006873f
C18969 net20 FILLER_0_9_223/a_572_375# 0.03118f
C18970 _420_/a_1308_423# _009_ 0.014359f
C18971 _369_/a_36_68# _154_ 0.042308f
C18972 FILLER_0_12_136/a_932_472# vdd 0.005266f
C18973 FILLER_0_12_136/a_484_472# vss 0.007054f
C18974 _070_ _058_ 0.07307f
C18975 net72 vdd 1.425686f
C18976 FILLER_0_15_116/a_572_375# net53 0.012526f
C18977 _085_ _161_ 0.008926f
C18978 _438_/a_448_472# net71 0.044454f
C18979 _421_/a_2665_112# _109_ 0.002029f
C18980 _412_/a_36_151# vss 0.003515f
C18981 _077_ FILLER_0_10_78/a_932_472# 0.002503f
C18982 result[7] FILLER_0_24_274/a_36_472# 0.006454f
C18983 _118_ _313_/a_67_603# 0.001793f
C18984 FILLER_0_12_136/a_572_375# FILLER_0_11_142/a_36_472# 0.001543f
C18985 _101_ _100_ 0.012073f
C18986 _021_ _432_/a_36_151# 0.033849f
C18987 FILLER_0_5_109/a_36_472# _155_ 0.001872f
C18988 FILLER_0_16_107/a_484_472# net70 0.002732f
C18989 FILLER_0_5_54/a_36_472# vss 0.001756f
C18990 FILLER_0_5_54/a_484_472# vdd 0.003166f
C18991 net33 net22 0.066751f
C18992 net16 _131_ 0.001308f
C18993 FILLER_0_7_104/a_1468_375# _154_ 0.003683f
C18994 _176_ _131_ 1.798819f
C18995 _093_ _438_/a_36_151# 0.088469f
C18996 _442_/a_2665_112# vdd 0.056153f
C18997 _415_/a_2665_112# result[1] 0.010555f
C18998 FILLER_0_10_37/a_124_375# net51 0.006198f
C18999 _030_ _367_/a_692_472# 0.002082f
C19000 _149_ FILLER_0_20_87/a_124_375# 0.004191f
C19001 _079_ FILLER_0_5_212/a_124_375# 0.005363f
C19002 _016_ state\[2\] 0.002937f
C19003 net15 FILLER_0_6_47/a_1380_472# 0.00464f
C19004 FILLER_0_1_98/a_124_375# _065_ 0.001136f
C19005 FILLER_0_16_241/a_36_472# vss 0.004432f
C19006 FILLER_0_18_177/a_1916_375# vdd 0.021f
C19007 output10/a_224_472# net19 0.037774f
C19008 net47 _450_/a_2449_156# 0.004488f
C19009 _449_/a_1204_472# _067_ 0.014354f
C19010 _112_ vss 0.145781f
C19011 FILLER_0_12_20/a_484_472# vss 0.001783f
C19012 FILLER_0_5_128/a_124_375# _152_ 0.017496f
C19013 ctln[6] net23 0.003826f
C19014 _141_ _145_ 0.094128f
C19015 _450_/a_1353_112# _039_ 0.019843f
C19016 FILLER_0_10_78/a_1380_472# FILLER_0_10_94/a_36_472# 0.013277f
C19017 FILLER_0_17_133/a_124_375# _137_ 0.009198f
C19018 _413_/a_448_472# vdd 0.016117f
C19019 net75 _425_/a_1308_423# 0.034219f
C19020 _413_/a_2248_156# vss 0.004157f
C19021 net66 trim[3] 0.00567f
C19022 net16 FILLER_0_18_37/a_572_375# 0.03477f
C19023 FILLER_0_15_282/a_124_375# _006_ 0.002249f
C19024 _256_/a_3368_68# _076_ 0.001183f
C19025 _398_/a_36_113# net17 0.002702f
C19026 _035_ trim_mask\[2\] 0.004455f
C19027 FILLER_0_17_72/a_1916_375# net53 0.001657f
C19028 FILLER_0_16_57/a_36_472# _183_ 0.004107f
C19029 FILLER_0_18_2/a_2724_472# net47 0.001551f
C19030 _068_ _261_/a_36_160# 0.008557f
C19031 _133_ _059_ 0.039848f
C19032 _034_ 0 0.304805f
C19033 _160_ 0 1.542665f
C19034 _166_ 0 0.299751f
C19035 trim[3] 0 1.777626f
C19036 output41/a_224_472# 0 2.38465f
C19037 clkc 0 0.763769f
C19038 net6 0 1.112469f
C19039 output6/a_224_472# 0 2.38465f
C19040 FILLER_0_12_196/a_36_472# 0 0.417394f
C19041 FILLER_0_12_196/a_124_375# 0 0.246306f
C19042 result[3] 0 0.50376f
C19043 net30 0 1.81422f
C19044 output30/a_224_472# 0 2.38465f
C19045 _047_ 0 0.374694f
C19046 _201_/a_67_603# 0 0.345683f
C19047 _416_/a_2560_156# 0 0.016968f
C19048 _416_/a_2665_112# 0 0.62251f
C19049 _416_/a_2248_156# 0 0.371662f
C19050 _416_/a_1204_472# 0 0.012971f
C19051 _416_/a_1000_472# 0 0.291735f
C19052 _416_/a_796_472# 0 0.023206f
C19053 _416_/a_1308_423# 0 0.279043f
C19054 _416_/a_448_472# 0 0.684413f
C19055 _416_/a_36_151# 0 1.43589f
C19056 FILLER_0_13_290/a_36_472# 0 0.417394f
C19057 FILLER_0_13_290/a_124_375# 0 0.246306f
C19058 _278_/a_36_160# 0 0.696445f
C19059 _145_ 0 0.546455f
C19060 FILLER_0_13_72/a_484_472# 0 0.345058f
C19061 FILLER_0_13_72/a_36_472# 0 0.404746f
C19062 FILLER_0_13_72/a_572_375# 0 0.232991f
C19063 FILLER_0_13_72/a_124_375# 0 0.185089f
C19064 FILLER_0_14_235/a_484_472# 0 0.345058f
C19065 FILLER_0_14_235/a_36_472# 0 0.404746f
C19066 FILLER_0_14_235/a_572_375# 0 0.232991f
C19067 FILLER_0_14_235/a_124_375# 0 0.185089f
C19068 _156_ 0 0.593796f
C19069 _107_ 0 0.391583f
C19070 _295_/a_36_472# 0 0.031137f
C19071 _022_ 0 0.387773f
C19072 _433_/a_2560_156# 0 0.016968f
C19073 _433_/a_2665_112# 0 0.62251f
C19074 _433_/a_2248_156# 0 0.371662f
C19075 _433_/a_1204_472# 0 0.012971f
C19076 _433_/a_1000_472# 0 0.291735f
C19077 _433_/a_796_472# 0 0.023206f
C19078 _433_/a_1308_423# 0 0.279043f
C19079 _433_/a_448_472# 0 0.684413f
C19080 _433_/a_36_151# 0 1.43589f
C19081 FILLER_0_5_148/a_484_472# 0 0.345058f
C19082 FILLER_0_5_148/a_36_472# 0 0.404746f
C19083 FILLER_0_5_148/a_572_375# 0 0.232991f
C19084 FILLER_0_5_148/a_124_375# 0 0.185089f
C19085 _167_ 0 0.285904f
C19086 _381_/a_36_472# 0 0.031137f
C19087 trim[2] 0 0.79181f
C19088 net40 0 1.845219f
C19089 output40/a_224_472# 0 2.38465f
C19090 cal_count\[0\] 0 0.893784f
C19091 _039_ 0 0.412301f
C19092 _450_/a_2449_156# 0 0.049992f
C19093 _450_/a_2225_156# 0 0.434082f
C19094 _450_/a_3129_107# 0 0.58406f
C19095 _450_/a_836_156# 0 0.019766f
C19096 _450_/a_1040_527# 0 0.302082f
C19097 _450_/a_1353_112# 0 0.286513f
C19098 _450_/a_448_472# 0 1.21246f
C19099 _450_/a_36_151# 0 1.31409f
C19100 rstn 0 1.86494f
C19101 FILLER_0_8_156/a_484_472# 0 0.345058f
C19102 FILLER_0_8_156/a_36_472# 0 0.404746f
C19103 FILLER_0_8_156/a_572_375# 0 0.232991f
C19104 FILLER_0_8_156/a_124_375# 0 0.185089f
C19105 FILLER_0_6_37/a_36_472# 0 0.417394f
C19106 FILLER_0_6_37/a_124_375# 0 0.246306f
C19107 FILLER_0_21_60/a_484_472# 0 0.345058f
C19108 FILLER_0_21_60/a_36_472# 0 0.404746f
C19109 FILLER_0_21_60/a_572_375# 0 0.232991f
C19110 FILLER_0_21_60/a_124_375# 0 0.185089f
C19111 FILLER_0_22_107/a_484_472# 0 0.345058f
C19112 FILLER_0_22_107/a_36_472# 0 0.404746f
C19113 FILLER_0_22_107/a_572_375# 0 0.232991f
C19114 FILLER_0_22_107/a_124_375# 0 0.185089f
C19115 FILLER_0_16_115/a_36_472# 0 0.417394f
C19116 FILLER_0_16_115/a_124_375# 0 0.246306f
C19117 FILLER_0_19_134/a_36_472# 0 0.417394f
C19118 FILLER_0_19_134/a_124_375# 0 0.246306f
C19119 FILLER_0_3_212/a_36_472# 0 0.417394f
C19120 FILLER_0_3_212/a_124_375# 0 0.246306f
C19121 FILLER_0_10_94/a_484_472# 0 0.345058f
C19122 FILLER_0_10_94/a_36_472# 0 0.404746f
C19123 FILLER_0_10_94/a_572_375# 0 0.232991f
C19124 FILLER_0_10_94/a_124_375# 0 0.185089f
C19125 FILLER_0_4_91/a_484_472# 0 0.345058f
C19126 FILLER_0_4_91/a_36_472# 0 0.404746f
C19127 FILLER_0_4_91/a_572_375# 0 0.232991f
C19128 FILLER_0_4_91/a_124_375# 0 0.185089f
C19129 net14 0 1.508711f
C19130 _202_/a_36_160# 0 0.696445f
C19131 FILLER_0_6_231/a_484_472# 0 0.345058f
C19132 FILLER_0_6_231/a_36_472# 0 0.404746f
C19133 FILLER_0_6_231/a_572_375# 0 0.232991f
C19134 FILLER_0_6_231/a_124_375# 0 0.185089f
C19135 vss 0 65.60368f
C19136 vdd 0 1.086009p
C19137 _006_ 0 0.41456f
C19138 _417_/a_2560_156# 0 0.016968f
C19139 _417_/a_2665_112# 0 0.62251f
C19140 _417_/a_2248_156# 0 0.371662f
C19141 _417_/a_1204_472# 0 0.012971f
C19142 _417_/a_1000_472# 0 0.291735f
C19143 _417_/a_796_472# 0 0.023206f
C19144 _417_/a_1308_423# 0 0.279043f
C19145 _417_/a_448_472# 0 0.684413f
C19146 _417_/a_36_151# 0 1.43589f
C19147 _146_ 0 0.35443f
C19148 mask\[6\] 0 1.246962f
C19149 _348_/a_49_472# 0 0.054843f
C19150 _365_/a_36_68# 0 0.150048f
C19151 _023_ 0 0.345812f
C19152 _434_/a_2560_156# 0 0.016968f
C19153 _434_/a_2665_112# 0 0.62251f
C19154 _434_/a_2248_156# 0 0.371662f
C19155 _434_/a_1204_472# 0 0.012971f
C19156 _434_/a_1000_472# 0 0.291735f
C19157 _434_/a_796_472# 0 0.023206f
C19158 _434_/a_1308_423# 0 0.279043f
C19159 _434_/a_448_472# 0 0.684413f
C19160 _434_/a_36_151# 0 1.43589f
C19161 FILLER_0_5_136/a_36_472# 0 0.417394f
C19162 FILLER_0_5_136/a_124_375# 0 0.246306f
C19163 FILLER_0_18_209/a_484_472# 0 0.345058f
C19164 FILLER_0_18_209/a_36_472# 0 0.404746f
C19165 FILLER_0_18_209/a_572_375# 0 0.232991f
C19166 FILLER_0_18_209/a_124_375# 0 0.185089f
C19167 FILLER_0_12_28/a_36_472# 0 0.417394f
C19168 FILLER_0_12_28/a_124_375# 0 0.246306f
C19169 _040_ 0 0.355703f
C19170 _451_/a_2449_156# 0 0.049992f
C19171 _451_/a_2225_156# 0 0.434082f
C19172 _451_/a_3129_107# 0 0.58406f
C19173 _451_/a_836_156# 0 0.019766f
C19174 _451_/a_1040_527# 0 0.302082f
C19175 _451_/a_1353_112# 0 0.286513f
C19176 _451_/a_448_472# 0 1.21246f
C19177 _451_/a_36_151# 0 1.31409f
C19178 FILLER_0_6_47/a_3172_472# 0 0.345058f
C19179 FILLER_0_6_47/a_2724_472# 0 0.33241f
C19180 FILLER_0_6_47/a_2276_472# 0 0.33241f
C19181 FILLER_0_6_47/a_1828_472# 0 0.33241f
C19182 FILLER_0_6_47/a_1380_472# 0 0.33241f
C19183 FILLER_0_6_47/a_932_472# 0 0.33241f
C19184 FILLER_0_6_47/a_484_472# 0 0.33241f
C19185 FILLER_0_6_47/a_36_472# 0 0.404746f
C19186 FILLER_0_6_47/a_3260_375# 0 0.233093f
C19187 FILLER_0_6_47/a_2812_375# 0 0.17167f
C19188 FILLER_0_6_47/a_2364_375# 0 0.17167f
C19189 FILLER_0_6_47/a_1916_375# 0 0.17167f
C19190 FILLER_0_6_47/a_1468_375# 0 0.17167f
C19191 FILLER_0_6_47/a_1020_375# 0 0.17167f
C19192 FILLER_0_6_47/a_572_375# 0 0.17167f
C19193 FILLER_0_6_47/a_124_375# 0 0.185915f
C19194 FILLER_0_21_150/a_36_472# 0 0.417394f
C19195 FILLER_0_21_150/a_124_375# 0 0.246306f
C19196 FILLER_0_15_180/a_484_472# 0 0.345058f
C19197 FILLER_0_15_180/a_36_472# 0 0.404746f
C19198 FILLER_0_15_180/a_572_375# 0 0.232991f
C19199 FILLER_0_15_180/a_124_375# 0 0.185089f
C19200 FILLER_0_22_128/a_3172_472# 0 0.345058f
C19201 FILLER_0_22_128/a_2724_472# 0 0.33241f
C19202 FILLER_0_22_128/a_2276_472# 0 0.33241f
C19203 FILLER_0_22_128/a_1828_472# 0 0.33241f
C19204 FILLER_0_22_128/a_1380_472# 0 0.33241f
C19205 FILLER_0_22_128/a_932_472# 0 0.33241f
C19206 FILLER_0_22_128/a_484_472# 0 0.33241f
C19207 FILLER_0_22_128/a_36_472# 0 0.404746f
C19208 FILLER_0_22_128/a_3260_375# 0 0.233093f
C19209 FILLER_0_22_128/a_2812_375# 0 0.17167f
C19210 FILLER_0_22_128/a_2364_375# 0 0.17167f
C19211 FILLER_0_22_128/a_1916_375# 0 0.17167f
C19212 FILLER_0_22_128/a_1468_375# 0 0.17167f
C19213 FILLER_0_22_128/a_1020_375# 0 0.17167f
C19214 FILLER_0_22_128/a_572_375# 0 0.17167f
C19215 FILLER_0_22_128/a_124_375# 0 0.185915f
C19216 FILLER_0_19_111/a_484_472# 0 0.345058f
C19217 FILLER_0_19_111/a_36_472# 0 0.404746f
C19218 FILLER_0_19_111/a_572_375# 0 0.232991f
C19219 FILLER_0_19_111/a_124_375# 0 0.185089f
C19220 FILLER_0_19_155/a_484_472# 0 0.345058f
C19221 FILLER_0_19_155/a_36_472# 0 0.404746f
C19222 FILLER_0_19_155/a_572_375# 0 0.232991f
C19223 FILLER_0_19_155/a_124_375# 0 0.185089f
C19224 net11 0 1.328455f
C19225 net21 0 1.922829f
C19226 _007_ 0 0.309495f
C19227 net77 0 1.39077f
C19228 _418_/a_2560_156# 0 0.016968f
C19229 _418_/a_2665_112# 0 0.62251f
C19230 _418_/a_2248_156# 0 0.371662f
C19231 _418_/a_1204_472# 0 0.012971f
C19232 _418_/a_1000_472# 0 0.291735f
C19233 _418_/a_796_472# 0 0.023206f
C19234 _418_/a_1308_423# 0 0.279043f
C19235 _418_/a_448_472# 0 0.684413f
C19236 _418_/a_36_151# 0 1.43589f
C19237 _220_/a_67_603# 0 0.345683f
C19238 FILLER_0_9_282/a_484_472# 0 0.345058f
C19239 FILLER_0_9_282/a_36_472# 0 0.404746f
C19240 FILLER_0_9_282/a_572_375# 0 0.232991f
C19241 FILLER_0_9_282/a_124_375# 0 0.185089f
C19242 FILLER_0_18_37/a_1380_472# 0 0.345058f
C19243 FILLER_0_18_37/a_932_472# 0 0.33241f
C19244 FILLER_0_18_37/a_484_472# 0 0.33241f
C19245 FILLER_0_18_37/a_36_472# 0 0.404746f
C19246 FILLER_0_18_37/a_1468_375# 0 0.233029f
C19247 FILLER_0_18_37/a_1020_375# 0 0.171606f
C19248 FILLER_0_18_37/a_572_375# 0 0.171606f
C19249 FILLER_0_18_37/a_124_375# 0 0.185399f
C19250 FILLER_0_2_127/a_36_472# 0 0.417394f
C19251 FILLER_0_2_127/a_124_375# 0 0.246306f
C19252 _157_ 0 0.531763f
C19253 _435_/a_2560_156# 0 0.016968f
C19254 _435_/a_2665_112# 0 0.62251f
C19255 _435_/a_2248_156# 0 0.371662f
C19256 _435_/a_1204_472# 0 0.012971f
C19257 _435_/a_1000_472# 0 0.291735f
C19258 _435_/a_796_472# 0 0.023206f
C19259 _435_/a_1308_423# 0 0.279043f
C19260 _435_/a_448_472# 0 0.684413f
C19261 _435_/a_36_151# 0 1.43589f
C19262 _108_ 0 0.411979f
C19263 _297_/a_36_472# 0 0.031137f
C19264 trim_mask\[3\] 0 1.081535f
C19265 _164_ 0 1.3268f
C19266 _383_/a_36_472# 0 0.031137f
C19267 _041_ 0 0.299289f
C19268 _452_/a_2449_156# 0 0.049992f
C19269 _452_/a_2225_156# 0 0.434082f
C19270 _452_/a_3129_107# 0 0.58406f
C19271 _452_/a_836_156# 0 0.019766f
C19272 _452_/a_1040_527# 0 0.302082f
C19273 _452_/a_1353_112# 0 0.286513f
C19274 _452_/a_448_472# 0 1.21246f
C19275 _452_/a_36_151# 0 1.31409f
C19276 FILLER_0_6_79/a_36_472# 0 0.417394f
C19277 FILLER_0_6_79/a_124_375# 0 0.246306f
C19278 net59 0 5.044369f
C19279 FILLER_0_15_59/a_484_472# 0 0.345058f
C19280 FILLER_0_15_59/a_36_472# 0 0.404746f
C19281 FILLER_0_15_59/a_572_375# 0 0.232991f
C19282 FILLER_0_15_59/a_124_375# 0 0.185089f
C19283 FILLER_0_3_221/a_1380_472# 0 0.345058f
C19284 FILLER_0_3_221/a_932_472# 0 0.33241f
C19285 FILLER_0_3_221/a_484_472# 0 0.33241f
C19286 FILLER_0_3_221/a_36_472# 0 0.404746f
C19287 FILLER_0_3_221/a_1468_375# 0 0.233029f
C19288 FILLER_0_3_221/a_1020_375# 0 0.171606f
C19289 FILLER_0_3_221/a_572_375# 0 0.171606f
C19290 FILLER_0_3_221/a_124_375# 0 0.185399f
C19291 FILLER_0_19_187/a_484_472# 0 0.345058f
C19292 FILLER_0_19_187/a_36_472# 0 0.404746f
C19293 FILLER_0_19_187/a_572_375# 0 0.232991f
C19294 FILLER_0_19_187/a_124_375# 0 0.185089f
C19295 FILLER_0_20_15/a_1380_472# 0 0.345058f
C19296 FILLER_0_20_15/a_932_472# 0 0.33241f
C19297 FILLER_0_20_15/a_484_472# 0 0.33241f
C19298 FILLER_0_20_15/a_36_472# 0 0.404746f
C19299 FILLER_0_20_15/a_1468_375# 0 0.233029f
C19300 FILLER_0_20_15/a_1020_375# 0 0.171606f
C19301 FILLER_0_20_15/a_572_375# 0 0.171606f
C19302 FILLER_0_20_15/a_124_375# 0 0.185399f
C19303 _204_/a_67_603# 0 0.345683f
C19304 _419_/a_2560_156# 0 0.016968f
C19305 _419_/a_2665_112# 0 0.62251f
C19306 _419_/a_2248_156# 0 0.371662f
C19307 _419_/a_1204_472# 0 0.012971f
C19308 _419_/a_1000_472# 0 0.291735f
C19309 _419_/a_796_472# 0 0.023206f
C19310 _419_/a_1308_423# 0 0.279043f
C19311 _419_/a_448_472# 0 0.684413f
C19312 _419_/a_36_151# 0 1.43589f
C19313 _054_ 0 0.522819f
C19314 _221_/a_36_160# 0 0.386641f
C19315 FILLER_0_9_270/a_484_472# 0 0.345058f
C19316 FILLER_0_9_270/a_36_472# 0 0.404746f
C19317 FILLER_0_9_270/a_572_375# 0 0.232991f
C19318 FILLER_0_9_270/a_124_375# 0 0.185089f
C19319 FILLER_0_1_192/a_36_472# 0 0.417394f
C19320 FILLER_0_1_192/a_124_375# 0 0.246306f
C19321 FILLER_0_13_80/a_36_472# 0 0.417394f
C19322 FILLER_0_13_80/a_124_375# 0 0.246306f
C19323 _153_ 0 1.165862f
C19324 _154_ 0 1.167112f
C19325 _367_/a_36_68# 0 0.150048f
C19326 _436_/a_2560_156# 0 0.016968f
C19327 _436_/a_2665_112# 0 0.62251f
C19328 _436_/a_2248_156# 0 0.371662f
C19329 _436_/a_1204_472# 0 0.012971f
C19330 _436_/a_1000_472# 0 0.291735f
C19331 _436_/a_796_472# 0 0.023206f
C19332 _436_/a_1308_423# 0 0.279043f
C19333 _436_/a_448_472# 0 0.684413f
C19334 _436_/a_36_151# 0 1.43589f
C19335 FILLER_0_10_107/a_484_472# 0 0.345058f
C19336 FILLER_0_10_107/a_36_472# 0 0.404746f
C19337 FILLER_0_10_107/a_572_375# 0 0.232991f
C19338 FILLER_0_10_107/a_124_375# 0 0.185089f
C19339 _168_ 0 0.336537f
C19340 net51 0 2.105066f
C19341 _042_ 0 0.323587f
C19342 _453_/a_2560_156# 0 0.016968f
C19343 _453_/a_2665_112# 0 0.62251f
C19344 _453_/a_2248_156# 0 0.371662f
C19345 _453_/a_1204_472# 0 0.012971f
C19346 _453_/a_1000_472# 0 0.291735f
C19347 _453_/a_796_472# 0 0.023206f
C19348 _453_/a_1308_423# 0 0.279043f
C19349 _453_/a_448_472# 0 0.684413f
C19350 _453_/a_36_151# 0 1.43589f
C19351 FILLER_0_19_142/a_36_472# 0 0.417394f
C19352 FILLER_0_19_142/a_124_375# 0 0.246306f
C19353 _048_ 0 0.358805f
C19354 _205_/a_36_160# 0 0.696445f
C19355 net43 0 1.236377f
C19356 FILLER_0_3_78/a_484_472# 0 0.345058f
C19357 FILLER_0_3_78/a_36_472# 0 0.404746f
C19358 FILLER_0_3_78/a_572_375# 0 0.232991f
C19359 FILLER_0_3_78/a_124_375# 0 0.185089f
C19360 _437_/a_2560_156# 0 0.016968f
C19361 _437_/a_2665_112# 0 0.62251f
C19362 _437_/a_2248_156# 0 0.371662f
C19363 _437_/a_1204_472# 0 0.012971f
C19364 _437_/a_1000_472# 0 0.291735f
C19365 _437_/a_796_472# 0 0.023206f
C19366 _437_/a_1308_423# 0 0.279043f
C19367 _437_/a_448_472# 0 0.684413f
C19368 _437_/a_36_151# 0 1.43589f
C19369 _109_ 0 0.319326f
C19370 _299_/a_36_472# 0 0.031137f
C19371 net37 0 1.529713f
C19372 _385_/a_36_68# 0 0.112263f
C19373 FILLER_0_0_266/a_36_472# 0 0.417394f
C19374 FILLER_0_0_266/a_124_375# 0 0.246306f
C19375 net12 0 1.263595f
C19376 net22 0 2.108509f
C19377 FILLER_0_9_290/a_36_472# 0 0.417394f
C19378 FILLER_0_9_290/a_124_375# 0 0.246306f
C19379 _223_/a_36_160# 0 0.696445f
C19380 FILLER_0_14_263/a_36_472# 0 0.417394f
C19381 FILLER_0_14_263/a_124_375# 0 0.246306f
C19382 _158_ 0 0.309522f
C19383 _369_/a_36_68# 0 0.150048f
C19384 net71 0 1.420869f
C19385 _438_/a_2560_156# 0 0.016968f
C19386 _438_/a_2665_112# 0 0.62251f
C19387 _438_/a_2248_156# 0 0.371662f
C19388 _438_/a_1204_472# 0 0.012971f
C19389 _438_/a_1000_472# 0 0.291735f
C19390 _438_/a_796_472# 0 0.023206f
C19391 _438_/a_1308_423# 0 0.279043f
C19392 _438_/a_448_472# 0 0.684413f
C19393 _438_/a_36_151# 0 1.43589f
C19394 FILLER_0_23_274/a_36_472# 0 0.417394f
C19395 FILLER_0_23_274/a_124_375# 0 0.246306f
C19396 FILLER_0_17_282/a_36_472# 0 0.417394f
C19397 FILLER_0_17_282/a_124_375# 0 0.246306f
C19398 FILLER_0_5_198/a_484_472# 0 0.345058f
C19399 FILLER_0_5_198/a_36_472# 0 0.404746f
C19400 FILLER_0_5_198/a_572_375# 0 0.232991f
C19401 FILLER_0_5_198/a_124_375# 0 0.185089f
C19402 _163_ 0 1.03762f
C19403 _169_ 0 0.245383f
C19404 _386_/a_848_380# 0 0.40208f
C19405 _386_/a_124_24# 0 0.591898f
C19406 FILLER_0_20_2/a_484_472# 0 0.345058f
C19407 FILLER_0_20_2/a_36_472# 0 0.404746f
C19408 FILLER_0_20_2/a_572_375# 0 0.232991f
C19409 FILLER_0_20_2/a_124_375# 0 0.185089f
C19410 FILLER_0_16_154/a_1380_472# 0 0.345058f
C19411 FILLER_0_16_154/a_932_472# 0 0.33241f
C19412 FILLER_0_16_154/a_484_472# 0 0.33241f
C19413 FILLER_0_16_154/a_36_472# 0 0.404746f
C19414 FILLER_0_16_154/a_1468_375# 0 0.233029f
C19415 FILLER_0_16_154/a_1020_375# 0 0.171606f
C19416 FILLER_0_16_154/a_572_375# 0 0.171606f
C19417 FILLER_0_16_154/a_124_375# 0 0.185399f
C19418 FILLER_0_0_232/a_36_472# 0 0.417394f
C19419 FILLER_0_0_232/a_124_375# 0 0.246306f
C19420 FILLER_0_19_195/a_36_472# 0 0.417394f
C19421 FILLER_0_19_195/a_124_375# 0 0.246306f
C19422 _049_ 0 0.329957f
C19423 net33 0 1.934915f
C19424 _207_/a_67_603# 0 0.345683f
C19425 FILLER_0_3_54/a_36_472# 0 0.417394f
C19426 FILLER_0_3_54/a_124_375# 0 0.246306f
C19427 FILLER_0_2_101/a_36_472# 0 0.417394f
C19428 FILLER_0_2_101/a_124_375# 0 0.246306f
C19429 trim_mask\[0\] 0 0.605753f
C19430 _439_/a_2560_156# 0 0.016968f
C19431 _439_/a_2665_112# 0 0.62251f
C19432 _439_/a_2248_156# 0 0.371662f
C19433 _439_/a_1204_472# 0 0.012971f
C19434 _439_/a_1000_472# 0 0.291735f
C19435 _439_/a_796_472# 0 0.023206f
C19436 _439_/a_1308_423# 0 0.279043f
C19437 _439_/a_448_472# 0 0.684413f
C19438 _439_/a_36_151# 0 1.43589f
C19439 _066_ 0 0.333041f
C19440 FILLER_0_23_44/a_1380_472# 0 0.345058f
C19441 FILLER_0_23_44/a_932_472# 0 0.33241f
C19442 FILLER_0_23_44/a_484_472# 0 0.33241f
C19443 FILLER_0_23_44/a_36_472# 0 0.404746f
C19444 FILLER_0_23_44/a_1468_375# 0 0.233029f
C19445 FILLER_0_23_44/a_1020_375# 0 0.171606f
C19446 FILLER_0_23_44/a_572_375# 0 0.171606f
C19447 FILLER_0_23_44/a_124_375# 0 0.185399f
C19448 FILLER_0_23_88/a_36_472# 0 0.417394f
C19449 FILLER_0_23_88/a_124_375# 0 0.246306f
C19450 FILLER_0_5_164/a_484_472# 0 0.345058f
C19451 FILLER_0_5_164/a_36_472# 0 0.404746f
C19452 FILLER_0_5_164/a_572_375# 0 0.232991f
C19453 FILLER_0_5_164/a_124_375# 0 0.185089f
C19454 _060_ 0 2.485177f
C19455 _113_ 0 2.833205f
C19456 _090_ 0 2.629271f
C19457 _310_/a_49_472# 0 0.098072f
C19458 _037_ 0 0.467089f
C19459 _170_ 0 0.413995f
C19460 _387_/a_36_113# 0 0.418095f
C19461 _208_/a_36_160# 0 0.696445f
C19462 FILLER_0_18_76/a_484_472# 0 0.345058f
C19463 FILLER_0_18_76/a_36_472# 0 0.404746f
C19464 FILLER_0_18_76/a_572_375# 0 0.232991f
C19465 FILLER_0_18_76/a_124_375# 0 0.185089f
C19466 _225_/a_36_160# 0 0.386641f
C19467 FILLER_0_2_177/a_484_472# 0 0.345058f
C19468 FILLER_0_2_177/a_36_472# 0 0.404746f
C19469 FILLER_0_2_177/a_572_375# 0 0.232991f
C19470 FILLER_0_2_177/a_124_375# 0 0.185089f
C19471 FILLER_0_2_111/a_1380_472# 0 0.345058f
C19472 FILLER_0_2_111/a_932_472# 0 0.33241f
C19473 FILLER_0_2_111/a_484_472# 0 0.33241f
C19474 FILLER_0_2_111/a_36_472# 0 0.404746f
C19475 FILLER_0_2_111/a_1468_375# 0 0.233029f
C19476 FILLER_0_2_111/a_1020_375# 0 0.171606f
C19477 FILLER_0_2_111/a_572_375# 0 0.171606f
C19478 FILLER_0_2_111/a_124_375# 0 0.185399f
C19479 FILLER_0_15_228/a_36_472# 0 0.417394f
C19480 FILLER_0_15_228/a_124_375# 0 0.246306f
C19481 net47 0 2.314376f
C19482 _242_/a_36_160# 0 0.696445f
C19483 _117_ 0 1.266251f
C19484 _311_/a_66_473# 0 0.11665f
C19485 _043_ 0 0.487279f
C19486 _190_/a_36_160# 0 0.696445f
C19487 FILLER_0_9_105/a_484_472# 0 0.345058f
C19488 FILLER_0_9_105/a_36_472# 0 0.404746f
C19489 FILLER_0_9_105/a_572_375# 0 0.232991f
C19490 FILLER_0_9_105/a_124_375# 0 0.185089f
C19491 FILLER_0_13_100/a_36_472# 0 0.417394f
C19492 FILLER_0_13_100/a_124_375# 0 0.246306f
C19493 FILLER_0_22_177/a_1380_472# 0 0.345058f
C19494 FILLER_0_22_177/a_932_472# 0 0.33241f
C19495 FILLER_0_22_177/a_484_472# 0 0.33241f
C19496 FILLER_0_22_177/a_36_472# 0 0.404746f
C19497 FILLER_0_22_177/a_1468_375# 0 0.233029f
C19498 FILLER_0_22_177/a_1020_375# 0 0.171606f
C19499 FILLER_0_22_177/a_572_375# 0 0.171606f
C19500 FILLER_0_22_177/a_124_375# 0 0.185399f
C19501 FILLER_0_15_2/a_484_472# 0 0.345058f
C19502 FILLER_0_15_2/a_36_472# 0 0.404746f
C19503 FILLER_0_15_2/a_572_375# 0 0.232991f
C19504 FILLER_0_15_2/a_124_375# 0 0.185089f
C19505 FILLER_0_15_10/a_36_472# 0 0.417394f
C19506 FILLER_0_15_10/a_124_375# 0 0.246306f
C19507 FILLER_0_19_171/a_1380_472# 0 0.345058f
C19508 FILLER_0_19_171/a_932_472# 0 0.33241f
C19509 FILLER_0_19_171/a_484_472# 0 0.33241f
C19510 FILLER_0_19_171/a_36_472# 0 0.404746f
C19511 FILLER_0_19_171/a_1468_375# 0 0.233029f
C19512 FILLER_0_19_171/a_1020_375# 0 0.171606f
C19513 FILLER_0_19_171/a_572_375# 0 0.171606f
C19514 FILLER_0_19_171/a_124_375# 0 0.185399f
C19515 net13 0 1.176306f
C19516 net23 0 2.091399f
C19517 FILLER_0_20_87/a_36_472# 0 0.417394f
C19518 FILLER_0_20_87/a_124_375# 0 0.246306f
C19519 FILLER_0_20_98/a_36_472# 0 0.417394f
C19520 FILLER_0_20_98/a_124_375# 0 0.246306f
C19521 _055_ 0 1.782885f
C19522 FILLER_0_18_53/a_484_472# 0 0.345058f
C19523 FILLER_0_18_53/a_36_472# 0 0.404746f
C19524 FILLER_0_18_53/a_572_375# 0 0.232991f
C19525 FILLER_0_18_53/a_124_375# 0 0.185089f
C19526 FILLER_0_2_165/a_36_472# 0 0.417394f
C19527 FILLER_0_2_165/a_124_375# 0 0.246306f
C19528 FILLER_0_15_205/a_36_472# 0 0.417394f
C19529 FILLER_0_15_205/a_124_375# 0 0.246306f
C19530 FILLER_0_23_282/a_484_472# 0 0.345058f
C19531 FILLER_0_23_282/a_36_472# 0 0.404746f
C19532 FILLER_0_23_282/a_572_375# 0 0.232991f
C19533 FILLER_0_23_282/a_124_375# 0 0.185089f
C19534 net42 0 1.067446f
C19535 net17 0 2.210219f
C19536 _172_ 0 0.265782f
C19537 _171_ 0 0.300355f
C19538 _389_/a_36_148# 0 0.388358f
C19539 _080_ 0 0.328202f
C19540 _260_/a_36_68# 0 0.112263f
C19541 FILLER_0_0_96/a_36_472# 0 0.417394f
C19542 FILLER_0_0_96/a_124_375# 0 0.246306f
C19543 FILLER_0_9_72/a_1380_472# 0 0.345058f
C19544 FILLER_0_9_72/a_932_472# 0 0.33241f
C19545 FILLER_0_9_72/a_484_472# 0 0.33241f
C19546 FILLER_0_9_72/a_36_472# 0 0.404746f
C19547 FILLER_0_9_72/a_1468_375# 0 0.233029f
C19548 FILLER_0_9_72/a_1020_375# 0 0.171606f
C19549 FILLER_0_9_72/a_572_375# 0 0.171606f
C19550 FILLER_0_9_72/a_124_375# 0 0.185399f
C19551 FILLER_0_20_31/a_36_472# 0 0.417394f
C19552 FILLER_0_20_31/a_124_375# 0 0.246306f
C19553 _227_/a_36_160# 0 0.386641f
C19554 _120_ 0 1.533088f
C19555 _313_/a_67_603# 0 0.345683f
C19556 FILLER_0_5_172/a_36_472# 0 0.417394f
C19557 FILLER_0_5_172/a_124_375# 0 0.246306f
C19558 FILLER_0_12_20/a_484_472# 0 0.345058f
C19559 FILLER_0_12_20/a_36_472# 0 0.404746f
C19560 FILLER_0_12_20/a_572_375# 0 0.232991f
C19561 FILLER_0_12_20/a_124_375# 0 0.185089f
C19562 _134_ 0 0.365972f
C19563 _062_ 0 1.717773f
C19564 _059_ 0 1.686761f
C19565 _261_/a_36_160# 0 0.386641f
C19566 _044_ 0 0.388801f
C19567 mask\[1\] 0 1.295078f
C19568 _192_/a_67_603# 0 0.345683f
C19569 FILLER_0_13_142/a_1380_472# 0 0.345058f
C19570 FILLER_0_13_142/a_932_472# 0 0.33241f
C19571 FILLER_0_13_142/a_484_472# 0 0.33241f
C19572 FILLER_0_13_142/a_36_472# 0 0.404746f
C19573 FILLER_0_13_142/a_1468_375# 0 0.233029f
C19574 FILLER_0_13_142/a_1020_375# 0 0.171606f
C19575 FILLER_0_13_142/a_572_375# 0 0.171606f
C19576 FILLER_0_13_142/a_124_375# 0 0.185399f
C19577 FILLER_0_9_60/a_484_472# 0 0.345058f
C19578 FILLER_0_9_60/a_36_472# 0 0.404746f
C19579 FILLER_0_9_60/a_572_375# 0 0.232991f
C19580 FILLER_0_9_60/a_124_375# 0 0.185089f
C19581 FILLER_0_7_233/a_36_472# 0 0.417394f
C19582 FILLER_0_7_233/a_124_375# 0 0.246306f
C19583 _228_/a_36_68# 0 0.69549f
C19584 FILLER_0_21_206/a_36_472# 0 0.417394f
C19585 FILLER_0_21_206/a_124_375# 0 0.246306f
C19586 _067_ 0 0.851951f
C19587 _135_ 0 0.339478f
C19588 _193_/a_36_160# 0 0.696445f
C19589 _180_ 0 0.390598f
C19590 cal_count\[1\] 0 1.568289f
C19591 FILLER_0_4_213/a_484_472# 0 0.345058f
C19592 FILLER_0_4_213/a_36_472# 0 0.404746f
C19593 FILLER_0_4_213/a_572_375# 0 0.232991f
C19594 FILLER_0_4_213/a_124_375# 0 0.185089f
C19595 FILLER_0_11_282/a_36_472# 0 0.417394f
C19596 FILLER_0_11_282/a_124_375# 0 0.246306f
C19597 FILLER_0_18_61/a_36_472# 0 0.417394f
C19598 FILLER_0_18_61/a_124_375# 0 0.246306f
C19599 FILLER_0_15_235/a_484_472# 0 0.345058f
C19600 FILLER_0_15_235/a_36_472# 0 0.404746f
C19601 FILLER_0_15_235/a_572_375# 0 0.232991f
C19602 FILLER_0_15_235/a_124_375# 0 0.185089f
C19603 FILLER_0_23_290/a_36_472# 0 0.417394f
C19604 FILLER_0_23_290/a_124_375# 0 0.246306f
C19605 _121_ 0 0.532847f
C19606 _315_/a_36_68# 0 0.052951f
C19607 _246_/a_36_68# 0 0.69549f
C19608 FILLER_0_5_181/a_36_472# 0 0.417394f
C19609 FILLER_0_5_181/a_124_375# 0 0.246306f
C19610 _082_ 0 0.619901f
C19611 net8 0 1.163723f
C19612 net18 0 2.032159f
C19613 _332_/a_36_472# 0 0.031137f
C19614 _179_ 0 0.336984f
C19615 _401_/a_36_68# 0 0.112263f
C19616 FILLER_0_14_107/a_1380_472# 0 0.345058f
C19617 FILLER_0_14_107/a_932_472# 0 0.33241f
C19618 FILLER_0_14_107/a_484_472# 0 0.33241f
C19619 FILLER_0_14_107/a_36_472# 0 0.404746f
C19620 FILLER_0_14_107/a_1468_375# 0 0.233029f
C19621 FILLER_0_14_107/a_1020_375# 0 0.171606f
C19622 FILLER_0_14_107/a_572_375# 0 0.171606f
C19623 FILLER_0_14_107/a_124_375# 0 0.185399f
C19624 _097_ 0 0.592554f
C19625 FILLER_0_1_204/a_36_472# 0 0.417394f
C19626 FILLER_0_1_204/a_124_375# 0 0.246306f
C19627 FILLER_0_15_72/a_484_472# 0 0.345058f
C19628 FILLER_0_15_72/a_36_472# 0 0.404746f
C19629 FILLER_0_15_72/a_572_375# 0 0.232991f
C19630 FILLER_0_15_72/a_124_375# 0 0.185089f
C19631 FILLER_0_17_104/a_1380_472# 0 0.345058f
C19632 FILLER_0_17_104/a_932_472# 0 0.33241f
C19633 FILLER_0_17_104/a_484_472# 0 0.33241f
C19634 FILLER_0_17_104/a_36_472# 0 0.404746f
C19635 FILLER_0_17_104/a_1468_375# 0 0.233029f
C19636 FILLER_0_17_104/a_1020_375# 0 0.171606f
C19637 FILLER_0_17_104/a_572_375# 0 0.171606f
C19638 FILLER_0_17_104/a_124_375# 0 0.185399f
C19639 FILLER_0_8_37/a_484_472# 0 0.345058f
C19640 FILLER_0_8_37/a_36_472# 0 0.404746f
C19641 FILLER_0_8_37/a_572_375# 0 0.232991f
C19642 FILLER_0_8_37/a_124_375# 0 0.185089f
C19643 FILLER_0_15_212/a_1380_472# 0 0.345058f
C19644 FILLER_0_15_212/a_932_472# 0 0.33241f
C19645 FILLER_0_15_212/a_484_472# 0 0.33241f
C19646 FILLER_0_15_212/a_36_472# 0 0.404746f
C19647 FILLER_0_15_212/a_1468_375# 0 0.233029f
C19648 FILLER_0_15_212/a_1020_375# 0 0.171606f
C19649 FILLER_0_15_212/a_572_375# 0 0.171606f
C19650 FILLER_0_15_212/a_124_375# 0 0.185399f
C19651 FILLER_0_23_60/a_36_472# 0 0.417394f
C19652 FILLER_0_23_60/a_124_375# 0 0.246306f
C19653 _123_ 0 0.344874f
C19654 _122_ 0 0.600118f
C19655 calibrate 0 1.343796f
C19656 _316_/a_848_380# 0 0.40208f
C19657 _316_/a_124_24# 0 0.591898f
C19658 _247_/a_36_160# 0 0.696445f
C19659 FILLER_0_12_50/a_36_472# 0 0.417394f
C19660 FILLER_0_12_50/a_124_375# 0 0.246306f
C19661 _084_ 0 0.296163f
C19662 cal_itt\[0\] 0 1.831055f
C19663 cal_itt\[1\] 0 1.705665f
C19664 FILLER_0_11_109/a_36_472# 0 0.417394f
C19665 FILLER_0_11_109/a_124_375# 0 0.246306f
C19666 _182_ 0 0.34197f
C19667 _402_/a_1948_68# 0 0.022025f
C19668 _402_/a_718_527# 0 0.001795f
C19669 _402_/a_56_567# 0 0.424713f
C19670 _402_/a_728_93# 0 0.65929f
C19671 _402_/a_1296_93# 0 0.317801f
C19672 _045_ 0 0.349338f
C19673 mask\[2\] 0 1.335688f
C19674 _195_/a_67_603# 0 0.345683f
C19675 _333_/a_36_160# 0 0.386641f
C19676 _098_ 0 1.816151f
C19677 _147_ 0 0.322539f
C19678 _350_/a_49_472# 0 0.054843f
C19679 FILLER_0_12_236/a_484_472# 0 0.345058f
C19680 FILLER_0_12_236/a_36_472# 0 0.404746f
C19681 FILLER_0_12_236/a_572_375# 0 0.232991f
C19682 FILLER_0_12_236/a_124_375# 0 0.185089f
C19683 FILLER_0_2_171/a_36_472# 0 0.417394f
C19684 FILLER_0_2_171/a_124_375# 0 0.246306f
C19685 _014_ 0 0.363432f
C19686 _317_/a_36_113# 0 0.418095f
C19687 _248_/a_36_68# 0 0.69549f
C19688 FILLER_0_17_38/a_484_472# 0 0.345058f
C19689 FILLER_0_17_38/a_36_472# 0 0.404746f
C19690 FILLER_0_17_38/a_572_375# 0 0.232991f
C19691 FILLER_0_17_38/a_124_375# 0 0.185089f
C19692 _001_ 0 0.285216f
C19693 _265_/a_244_68# 0 0.138666f
C19694 _196_/a_36_160# 0 0.696445f
C19695 FILLER_0_6_90/a_484_472# 0 0.345058f
C19696 FILLER_0_6_90/a_36_472# 0 0.404746f
C19697 FILLER_0_6_90/a_572_375# 0 0.232991f
C19698 FILLER_0_6_90/a_124_375# 0 0.185089f
C19699 _183_ 0 0.356629f
C19700 _334_/a_36_160# 0 0.386641f
C19701 _282_/a_36_160# 0 0.386641f
C19702 _024_ 0 0.451815f
C19703 _009_ 0 0.397943f
C19704 _420_/a_2560_156# 0 0.016968f
C19705 _420_/a_2665_112# 0 0.62251f
C19706 _420_/a_2248_156# 0 0.371662f
C19707 _420_/a_1204_472# 0 0.012971f
C19708 _420_/a_1000_472# 0 0.291735f
C19709 _420_/a_796_472# 0 0.023206f
C19710 _420_/a_1308_423# 0 0.279043f
C19711 _420_/a_448_472# 0 0.684413f
C19712 _420_/a_36_151# 0 1.43589f
C19713 clk 0 1.162312f
C19714 FILLER_0_8_2/a_36_472# 0 0.417394f
C19715 FILLER_0_8_2/a_124_375# 0 0.246306f
C19716 FILLER_0_8_24/a_484_472# 0 0.345058f
C19717 FILLER_0_8_24/a_36_472# 0 0.404746f
C19718 FILLER_0_8_24/a_572_375# 0 0.232991f
C19719 FILLER_0_8_24/a_124_375# 0 0.185089f
C19720 _124_ 0 0.294081f
C19721 _118_ 0 1.378735f
C19722 _071_ 0 1.600488f
C19723 net9 0 1.13171f
C19724 net19 0 1.889339f
C19725 _138_ 0 0.33132f
C19726 _137_ 0 1.178616f
C19727 _335_/a_49_472# 0 0.054843f
C19728 _404_/a_36_472# 0 0.031137f
C19729 FILLER_0_20_107/a_36_472# 0 0.417394f
C19730 FILLER_0_20_107/a_124_375# 0 0.246306f
C19731 FILLER_0_9_142/a_36_472# 0 0.417394f
C19732 FILLER_0_9_142/a_124_375# 0 0.246306f
C19733 _099_ 0 1.152785f
C19734 _283_/a_36_472# 0 0.031137f
C19735 mask\[7\] 0 1.477838f
C19736 _352_/a_49_472# 0 0.054843f
C19737 _010_ 0 0.377779f
C19738 _421_/a_2560_156# 0 0.016968f
C19739 _421_/a_2665_112# 0 0.62251f
C19740 _421_/a_2248_156# 0 0.371662f
C19741 _421_/a_1204_472# 0 0.012971f
C19742 _421_/a_1000_472# 0 0.291735f
C19743 _421_/a_796_472# 0 0.023206f
C19744 _421_/a_1308_423# 0 0.279043f
C19745 _421_/a_448_472# 0 0.684413f
C19746 _421_/a_36_151# 0 1.43589f
C19747 FILLER_0_1_212/a_36_472# 0 0.417394f
C19748 FILLER_0_1_212/a_124_375# 0 0.246306f
C19749 FILLER_0_8_239/a_36_472# 0 0.417394f
C19750 FILLER_0_8_239/a_124_375# 0 0.246306f
C19751 _125_ 0 1.526603f
C19752 _058_ 0 1.483584f
C19753 FILLER_0_6_177/a_484_472# 0 0.345058f
C19754 FILLER_0_6_177/a_36_472# 0 0.404746f
C19755 FILLER_0_6_177/a_572_375# 0 0.232991f
C19756 FILLER_0_6_177/a_124_375# 0 0.185089f
C19757 state\[1\] 0 2.652405f
C19758 _267_/a_36_472# 0 0.137725f
C19759 _184_ 0 0.350066f
C19760 cal_count\[2\] 0 1.971854f
C19761 _405_/a_67_603# 0 0.345683f
C19762 _018_ 0 0.358633f
C19763 _046_ 0 0.361963f
C19764 _198_/a_67_603# 0 0.345683f
C19765 _094_ 0 1.263877f
C19766 _100_ 0 0.333135f
C19767 net36 0 2.262756f
C19768 FILLER_0_17_133/a_36_472# 0 0.417394f
C19769 FILLER_0_17_133/a_124_375# 0 0.246306f
C19770 _025_ 0 0.350324f
C19771 _148_ 0 0.325709f
C19772 _422_/a_2560_156# 0 0.016968f
C19773 _422_/a_2665_112# 0 0.62251f
C19774 _422_/a_2248_156# 0 0.371662f
C19775 _422_/a_1204_472# 0 0.012971f
C19776 _422_/a_1000_472# 0 0.291735f
C19777 _422_/a_796_472# 0 0.023206f
C19778 _422_/a_1308_423# 0 0.279043f
C19779 _422_/a_448_472# 0 0.684413f
C19780 _422_/a_36_151# 0 1.43589f
C19781 FILLER_0_1_266/a_484_472# 0 0.345058f
C19782 FILLER_0_1_266/a_36_472# 0 0.404746f
C19783 FILLER_0_1_266/a_572_375# 0 0.232991f
C19784 FILLER_0_1_266/a_124_375# 0 0.185089f
C19785 _152_ 0 0.918583f
C19786 _081_ 0 1.140656f
C19787 _370_/a_848_380# 0 0.40208f
C19788 _370_/a_124_24# 0 0.591898f
C19789 FILLER_0_24_274/a_1380_472# 0 0.345058f
C19790 FILLER_0_24_274/a_932_472# 0 0.33241f
C19791 FILLER_0_24_274/a_484_472# 0 0.33241f
C19792 FILLER_0_24_274/a_36_472# 0 0.404746f
C19793 FILLER_0_24_274/a_1468_375# 0 0.233029f
C19794 FILLER_0_24_274/a_1020_375# 0 0.171606f
C19795 FILLER_0_24_274/a_572_375# 0 0.171606f
C19796 FILLER_0_24_274/a_124_375# 0 0.185399f
C19797 _185_ 0 0.386917f
C19798 _406_/a_36_159# 0 0.374116f
C19799 _337_/a_49_472# 0 0.054843f
C19800 _199_/a_36_160# 0 0.696445f
C19801 _285_/a_36_472# 0 0.031137f
C19802 _354_/a_49_472# 0 0.054843f
C19803 _012_ 0 0.75195f
C19804 _423_/a_2560_156# 0 0.016968f
C19805 _423_/a_2665_112# 0 0.62251f
C19806 _423_/a_2248_156# 0 0.371662f
C19807 _423_/a_1204_472# 0 0.012971f
C19808 _423_/a_1000_472# 0 0.291735f
C19809 _423_/a_796_472# 0 0.023206f
C19810 _423_/a_1308_423# 0 0.279043f
C19811 _423_/a_448_472# 0 0.684413f
C19812 _423_/a_36_151# 0 1.43589f
C19813 FILLER_0_5_88/a_36_472# 0 0.417394f
C19814 FILLER_0_5_88/a_124_375# 0 0.246306f
C19815 trim_mask\[1\] 0 1.020743f
C19816 _029_ 0 0.308904f
C19817 _440_/a_2560_156# 0 0.016968f
C19818 _440_/a_2665_112# 0 0.62251f
C19819 _440_/a_2248_156# 0 0.371662f
C19820 _440_/a_1204_472# 0 0.012971f
C19821 _440_/a_1000_472# 0 0.291735f
C19822 _440_/a_796_472# 0 0.023206f
C19823 _440_/a_1308_423# 0 0.279043f
C19824 _440_/a_448_472# 0 0.684413f
C19825 _440_/a_36_151# 0 1.43589f
C19826 _159_ 0 0.351814f
C19827 _371_/a_36_113# 0 0.418095f
C19828 FILLER_0_17_56/a_484_472# 0 0.345058f
C19829 FILLER_0_17_56/a_36_472# 0 0.404746f
C19830 FILLER_0_17_56/a_572_375# 0 0.232991f
C19831 FILLER_0_17_56/a_124_375# 0 0.185089f
C19832 _083_ 0 0.527882f
C19833 _078_ 0 0.904554f
C19834 _269_/a_36_472# 0 0.031137f
C19835 _181_ 0 0.829168f
C19836 _407_/a_36_472# 0 0.031137f
C19837 _019_ 0 0.32907f
C19838 _139_ 0 0.346404f
C19839 FILLER_0_14_123/a_36_472# 0 0.417394f
C19840 FILLER_0_14_123/a_124_375# 0 0.246306f
C19841 _005_ 0 0.340993f
C19842 _101_ 0 0.280497f
C19843 _424_/a_2560_156# 0 0.016968f
C19844 _424_/a_2665_112# 0 0.62251f
C19845 _424_/a_2248_156# 0 0.371662f
C19846 _424_/a_1204_472# 0 0.012971f
C19847 _424_/a_1000_472# 0 0.291735f
C19848 _424_/a_796_472# 0 0.023206f
C19849 _424_/a_1308_423# 0 0.279043f
C19850 _424_/a_448_472# 0 0.684413f
C19851 _424_/a_36_151# 0 1.43589f
C19852 _026_ 0 0.320379f
C19853 _149_ 0 0.305496f
C19854 FILLER_0_5_54/a_1380_472# 0 0.345058f
C19855 FILLER_0_5_54/a_932_472# 0 0.33241f
C19856 FILLER_0_5_54/a_484_472# 0 0.33241f
C19857 FILLER_0_5_54/a_36_472# 0 0.404746f
C19858 FILLER_0_5_54/a_1468_375# 0 0.233029f
C19859 FILLER_0_5_54/a_1020_375# 0 0.171606f
C19860 FILLER_0_5_54/a_572_375# 0 0.171606f
C19861 FILLER_0_5_54/a_124_375# 0 0.185399f
C19862 FILLER_0_17_142/a_484_472# 0 0.345058f
C19863 FILLER_0_17_142/a_36_472# 0 0.404746f
C19864 FILLER_0_17_142/a_572_375# 0 0.232991f
C19865 FILLER_0_17_142/a_124_375# 0 0.185089f
C19866 _068_ 0 3.162692f
C19867 _076_ 0 3.812442f
C19868 _133_ 0 1.430901f
C19869 _070_ 0 3.115722f
C19870 _372_/a_170_472# 0 0.077257f
C19871 net49 0 5.140563f
C19872 _030_ 0 0.307083f
C19873 net66 0 1.472669f
C19874 _441_/a_2560_156# 0 0.016968f
C19875 _441_/a_2665_112# 0 0.62251f
C19876 _441_/a_2248_156# 0 0.371662f
C19877 _441_/a_1204_472# 0 0.012971f
C19878 _441_/a_1000_472# 0 0.291735f
C19879 _441_/a_796_472# 0 0.023206f
C19880 _441_/a_1308_423# 0 0.279043f
C19881 _441_/a_448_472# 0 0.684413f
C19882 _441_/a_36_151# 0 1.43589f
C19883 FILLER_0_5_206/a_36_472# 0 0.417394f
C19884 FILLER_0_5_206/a_124_375# 0 0.246306f
C19885 fanout49/a_36_160# 0 0.696445f
C19886 FILLER_0_8_247/a_1380_472# 0 0.345058f
C19887 FILLER_0_8_247/a_932_472# 0 0.33241f
C19888 FILLER_0_8_247/a_484_472# 0 0.33241f
C19889 FILLER_0_8_247/a_36_472# 0 0.404746f
C19890 FILLER_0_8_247/a_1468_375# 0 0.233029f
C19891 FILLER_0_8_247/a_1020_375# 0 0.171606f
C19892 FILLER_0_8_247/a_572_375# 0 0.171606f
C19893 FILLER_0_8_247/a_124_375# 0 0.185399f
C19894 FILLER_0_12_220/a_1380_472# 0 0.345058f
C19895 FILLER_0_12_220/a_932_472# 0 0.33241f
C19896 FILLER_0_12_220/a_484_472# 0 0.33241f
C19897 FILLER_0_12_220/a_36_472# 0 0.404746f
C19898 FILLER_0_12_220/a_1468_375# 0 0.233029f
C19899 FILLER_0_12_220/a_1020_375# 0 0.171606f
C19900 FILLER_0_12_220/a_572_375# 0 0.171606f
C19901 FILLER_0_12_220/a_124_375# 0 0.185399f
C19902 FILLER_0_21_286/a_484_472# 0 0.345058f
C19903 FILLER_0_21_286/a_36_472# 0 0.404746f
C19904 FILLER_0_21_286/a_572_375# 0 0.232991f
C19905 FILLER_0_21_286/a_124_375# 0 0.185089f
C19906 _140_ 0 1.276518f
C19907 _339_/a_36_160# 0 0.386641f
C19908 _095_ 0 2.689027f
C19909 _186_ 0 0.580923f
C19910 _408_/a_1936_472# 0 0.009918f
C19911 _408_/a_718_524# 0 0.005143f
C19912 _408_/a_56_524# 0 0.41096f
C19913 _408_/a_728_93# 0 0.654825f
C19914 _408_/a_1336_472# 0 0.316639f
C19915 FILLER_0_20_169/a_36_472# 0 0.417394f
C19916 FILLER_0_20_169/a_124_375# 0 0.246306f
C19917 _210_/a_67_603# 0 0.345683f
C19918 _425_/a_2560_156# 0 0.016968f
C19919 _425_/a_2665_112# 0 0.62251f
C19920 _425_/a_2248_156# 0 0.371662f
C19921 _425_/a_1204_472# 0 0.012971f
C19922 _425_/a_1000_472# 0 0.291735f
C19923 _425_/a_796_472# 0 0.023206f
C19924 _425_/a_1308_423# 0 0.279043f
C19925 _425_/a_448_472# 0 0.684413f
C19926 _425_/a_36_151# 0 1.43589f
C19927 net5 0 0.610761f
C19928 input5/a_36_113# 0 0.418095f
C19929 FILLER_0_11_78/a_484_472# 0 0.345058f
C19930 FILLER_0_11_78/a_36_472# 0 0.404746f
C19931 FILLER_0_11_78/a_572_375# 0 0.232991f
C19932 FILLER_0_11_78/a_124_375# 0 0.185089f
C19933 _102_ 0 0.335308f
C19934 _287_/a_36_472# 0 0.031137f
C19935 mask\[9\] 0 1.383606f
C19936 _356_/a_36_472# 0 0.031137f
C19937 _031_ 0 0.417351f
C19938 net69 0 1.020293f
C19939 _442_/a_2560_156# 0 0.016968f
C19940 _442_/a_2665_112# 0 0.62251f
C19941 _442_/a_2248_156# 0 0.371662f
C19942 _442_/a_1204_472# 0 0.012971f
C19943 _442_/a_1000_472# 0 0.291735f
C19944 _442_/a_796_472# 0 0.023206f
C19945 _442_/a_1308_423# 0 0.279043f
C19946 _442_/a_448_472# 0 0.684413f
C19947 _442_/a_36_151# 0 1.43589f
C19948 net64 0 2.598514f
C19949 fanout59/a_36_160# 0 0.696445f
C19950 FILLER_0_14_99/a_36_472# 0 0.417394f
C19951 FILLER_0_14_99/a_124_375# 0 0.246306f
C19952 _038_ 0 0.362839f
C19953 _136_ 0 1.345638f
C19954 _390_/a_36_68# 0 0.150048f
C19955 FILLER_0_15_282/a_484_472# 0 0.345058f
C19956 FILLER_0_15_282/a_36_472# 0 0.404746f
C19957 FILLER_0_15_282/a_572_375# 0 0.232991f
C19958 FILLER_0_15_282/a_124_375# 0 0.185089f
C19959 FILLER_0_11_124/a_36_472# 0 0.417394f
C19960 FILLER_0_11_124/a_124_375# 0 0.246306f
C19961 FILLER_0_11_135/a_36_472# 0 0.417394f
C19962 FILLER_0_11_135/a_124_375# 0 0.246306f
C19963 _188_ 0 0.349407f
C19964 cal_count\[3\] 0 1.862896f
C19965 _050_ 0 0.622354f
C19966 _211_/a_36_160# 0 0.386641f
C19967 net4 0 2.711508f
C19968 en 0 0.833743f
C19969 input4/a_36_68# 0 0.69549f
C19970 _426_/a_2560_156# 0 0.016968f
C19971 _426_/a_2665_112# 0 0.62251f
C19972 _426_/a_2248_156# 0 0.371662f
C19973 _426_/a_1204_472# 0 0.012971f
C19974 _426_/a_1000_472# 0 0.291735f
C19975 _426_/a_796_472# 0 0.023206f
C19976 _426_/a_1308_423# 0 0.279043f
C19977 _426_/a_448_472# 0 0.684413f
C19978 _426_/a_36_151# 0 1.43589f
C19979 _027_ 0 0.302949f
C19980 _150_ 0 0.320497f
C19981 FILLER_0_18_107/a_3172_472# 0 0.345058f
C19982 FILLER_0_18_107/a_2724_472# 0 0.33241f
C19983 FILLER_0_18_107/a_2276_472# 0 0.33241f
C19984 FILLER_0_18_107/a_1828_472# 0 0.33241f
C19985 FILLER_0_18_107/a_1380_472# 0 0.33241f
C19986 FILLER_0_18_107/a_932_472# 0 0.33241f
C19987 FILLER_0_18_107/a_484_472# 0 0.33241f
C19988 FILLER_0_18_107/a_36_472# 0 0.404746f
C19989 FILLER_0_18_107/a_3260_375# 0 0.233093f
C19990 FILLER_0_18_107/a_2812_375# 0 0.17167f
C19991 FILLER_0_18_107/a_2364_375# 0 0.17167f
C19992 FILLER_0_18_107/a_1916_375# 0 0.17167f
C19993 FILLER_0_18_107/a_1468_375# 0 0.17167f
C19994 FILLER_0_18_107/a_1020_375# 0 0.17167f
C19995 FILLER_0_18_107/a_572_375# 0 0.17167f
C19996 FILLER_0_18_107/a_124_375# 0 0.185915f
C19997 trim_mask\[4\] 0 0.987791f
C19998 _032_ 0 0.34876f
C19999 _443_/a_2560_156# 0 0.016968f
C20000 _443_/a_2665_112# 0 0.62251f
C20001 _443_/a_2248_156# 0 0.371662f
C20002 _443_/a_1204_472# 0 0.012971f
C20003 _443_/a_1000_472# 0 0.291735f
C20004 _443_/a_796_472# 0 0.023206f
C20005 _443_/a_1308_423# 0 0.279043f
C20006 _443_/a_448_472# 0 0.684413f
C20007 _443_/a_36_151# 0 1.43589f
C20008 _061_ 0 0.84986f
C20009 _056_ 0 2.393362f
C20010 _374_/a_36_68# 0 0.112263f
C20011 fanout58/a_36_160# 0 0.696445f
C20012 net74 0 1.237373f
C20013 fanout69/a_36_113# 0 0.418095f
C20014 _173_ 0 0.339446f
C20015 FILLER_0_3_142/a_36_472# 0 0.417394f
C20016 FILLER_0_3_142/a_124_375# 0 0.246306f
C20017 FILLER_0_17_64/a_36_472# 0 0.417394f
C20018 FILLER_0_17_64/a_124_375# 0 0.246306f
C20019 FILLER_0_11_101/a_484_472# 0 0.345058f
C20020 FILLER_0_11_101/a_36_472# 0 0.404746f
C20021 FILLER_0_11_101/a_572_375# 0 0.232991f
C20022 FILLER_0_11_101/a_124_375# 0 0.185089f
C20023 FILLER_0_22_86/a_1380_472# 0 0.345058f
C20024 FILLER_0_22_86/a_932_472# 0 0.33241f
C20025 FILLER_0_22_86/a_484_472# 0 0.33241f
C20026 FILLER_0_22_86/a_36_472# 0 0.404746f
C20027 FILLER_0_22_86/a_1468_375# 0 0.233029f
C20028 FILLER_0_22_86/a_1020_375# 0 0.171606f
C20029 FILLER_0_22_86/a_572_375# 0 0.171606f
C20030 FILLER_0_22_86/a_124_375# 0 0.185399f
C20031 net24 0 1.61895f
C20032 net3 0 0.740676f
C20033 input3/a_36_113# 0 0.418095f
C20034 _103_ 0 0.350464f
C20035 _289_/a_36_472# 0 0.031137f
C20036 _151_ 0 0.300777f
C20037 _427_/a_2560_156# 0 0.016968f
C20038 _427_/a_2665_112# 0 0.91969f
C20039 _427_/a_2248_156# 0 0.30886f
C20040 _427_/a_1204_472# 0 0.012971f
C20041 _427_/a_1000_472# 0 0.291735f
C20042 _427_/a_796_472# 0 0.023206f
C20043 _427_/a_1308_423# 0 0.279043f
C20044 _427_/a_448_472# 0 0.684413f
C20045 _427_/a_36_151# 0 1.43587f
C20046 FILLER_0_17_161/a_36_472# 0 0.417394f
C20047 FILLER_0_17_161/a_124_375# 0 0.246306f
C20048 FILLER_0_18_139/a_1380_472# 0 0.345058f
C20049 FILLER_0_18_139/a_932_472# 0 0.33241f
C20050 FILLER_0_18_139/a_484_472# 0 0.33241f
C20051 FILLER_0_18_139/a_36_472# 0 0.404746f
C20052 FILLER_0_18_139/a_1468_375# 0 0.233029f
C20053 FILLER_0_18_139/a_1020_375# 0 0.171606f
C20054 FILLER_0_18_139/a_572_375# 0 0.171606f
C20055 FILLER_0_18_139/a_124_375# 0 0.185399f
C20056 _161_ 0 0.592909f
C20057 _162_ 0 0.597238f
C20058 _375_/a_36_68# 0 0.048026f
C20059 trim_val\[0\] 0 0.742779f
C20060 net67 0 1.662327f
C20061 _444_/a_2560_156# 0 0.016968f
C20062 _444_/a_2665_112# 0 0.62251f
C20063 _444_/a_2248_156# 0 0.371662f
C20064 _444_/a_1204_472# 0 0.012971f
C20065 _444_/a_1000_472# 0 0.291735f
C20066 _444_/a_796_472# 0 0.023206f
C20067 _444_/a_1308_423# 0 0.279043f
C20068 _444_/a_448_472# 0 0.684413f
C20069 _444_/a_36_151# 0 1.43589f
C20070 net65 0 0.804072f
C20071 fanout57/a_36_113# 0 0.418095f
C20072 fanout68/a_36_113# 0 0.418095f
C20073 FILLER_0_12_2/a_484_472# 0 0.345058f
C20074 FILLER_0_12_2/a_36_472# 0 0.404746f
C20075 FILLER_0_12_2/a_572_375# 0 0.232991f
C20076 FILLER_0_12_2/a_124_375# 0 0.185089f
C20077 net79 0 1.584979f
C20078 fanout79/a_36_160# 0 0.386641f
C20079 _392_/a_36_68# 0 0.112263f
C20080 FILLER_0_13_228/a_36_472# 0 0.417394f
C20081 FILLER_0_13_228/a_124_375# 0 0.246306f
C20082 FILLER_0_13_206/a_36_472# 0 0.417394f
C20083 FILLER_0_13_206/a_124_375# 0 0.246306f
C20084 FILLER_0_20_177/a_1380_472# 0 0.345058f
C20085 FILLER_0_20_177/a_932_472# 0 0.33241f
C20086 FILLER_0_20_177/a_484_472# 0 0.33241f
C20087 FILLER_0_20_177/a_36_472# 0 0.404746f
C20088 FILLER_0_20_177/a_1468_375# 0 0.233029f
C20089 FILLER_0_20_177/a_1020_375# 0 0.171606f
C20090 FILLER_0_20_177/a_572_375# 0 0.171606f
C20091 FILLER_0_20_177/a_124_375# 0 0.185399f
C20092 _051_ 0 0.349381f
C20093 _213_/a_67_603# 0 0.345683f
C20094 net2 0 0.461658f
C20095 input2/a_36_113# 0 0.418095f
C20096 _129_ 0 0.926508f
C20097 _131_ 0 1.734297f
C20098 _359_/a_36_488# 0 0.101145f
C20099 FILLER_0_11_64/a_36_472# 0 0.417394f
C20100 FILLER_0_11_64/a_124_375# 0 0.246306f
C20101 state\[2\] 0 0.607433f
C20102 net53 0 4.483899f
C20103 _017_ 0 0.334329f
C20104 net70 0 1.238296f
C20105 _428_/a_2560_156# 0 0.016968f
C20106 _428_/a_2665_112# 0 0.62251f
C20107 _428_/a_2248_156# 0 0.371662f
C20108 _428_/a_1204_472# 0 0.012971f
C20109 _428_/a_1000_472# 0 0.291735f
C20110 _428_/a_796_472# 0 0.023206f
C20111 _428_/a_1308_423# 0 0.279043f
C20112 _428_/a_448_472# 0 0.684413f
C20113 _428_/a_36_151# 0 1.43589f
C20114 FILLER_0_5_72/a_1380_472# 0 0.345058f
C20115 FILLER_0_5_72/a_932_472# 0 0.33241f
C20116 FILLER_0_5_72/a_484_472# 0 0.33241f
C20117 FILLER_0_5_72/a_36_472# 0 0.404746f
C20118 FILLER_0_5_72/a_1468_375# 0 0.233029f
C20119 FILLER_0_5_72/a_1020_375# 0 0.171606f
C20120 FILLER_0_5_72/a_572_375# 0 0.171606f
C20121 FILLER_0_5_72/a_124_375# 0 0.185399f
C20122 _376_/a_36_160# 0 0.386641f
C20123 trim_val\[1\] 0 0.683578f
C20124 _445_/a_2560_156# 0 0.016968f
C20125 _445_/a_2665_112# 0 0.62251f
C20126 _445_/a_2248_156# 0 0.371662f
C20127 _445_/a_1204_472# 0 0.012971f
C20128 _445_/a_1000_472# 0 0.291735f
C20129 _445_/a_796_472# 0 0.023206f
C20130 _445_/a_1308_423# 0 0.279043f
C20131 _445_/a_448_472# 0 0.684413f
C20132 _445_/a_36_151# 0 1.43589f
C20133 fanout67/a_36_160# 0 0.386641f
C20134 fanout56/a_36_113# 0 0.418095f
C20135 net78 0 0.686263f
C20136 fanout78/a_36_113# 0 0.418095f
C20137 _174_ 0 0.979741f
C20138 FILLER_0_0_198/a_36_472# 0 0.417394f
C20139 FILLER_0_0_198/a_124_375# 0 0.246306f
C20140 FILLER_0_15_290/a_36_472# 0 0.417394f
C20141 FILLER_0_15_290/a_124_375# 0 0.246306f
C20142 FILLER_0_24_290/a_36_472# 0 0.417394f
C20143 FILLER_0_24_290/a_124_375# 0 0.246306f
C20144 FILLER_0_4_107/a_1380_472# 0 0.345058f
C20145 FILLER_0_4_107/a_932_472# 0 0.33241f
C20146 FILLER_0_4_107/a_484_472# 0 0.33241f
C20147 FILLER_0_4_107/a_36_472# 0 0.404746f
C20148 FILLER_0_4_107/a_1468_375# 0 0.233029f
C20149 FILLER_0_4_107/a_1020_375# 0 0.171606f
C20150 FILLER_0_4_107/a_572_375# 0 0.171606f
C20151 FILLER_0_4_107/a_124_375# 0 0.185399f
C20152 FILLER_0_7_104/a_1380_472# 0 0.345058f
C20153 FILLER_0_7_104/a_932_472# 0 0.33241f
C20154 FILLER_0_7_104/a_484_472# 0 0.33241f
C20155 FILLER_0_7_104/a_36_472# 0 0.404746f
C20156 FILLER_0_7_104/a_1468_375# 0 0.233029f
C20157 FILLER_0_7_104/a_1020_375# 0 0.171606f
C20158 FILLER_0_7_104/a_572_375# 0 0.171606f
C20159 FILLER_0_7_104/a_124_375# 0 0.185399f
C20160 _214_/a_36_160# 0 0.386641f
C20161 net1 0 0.364811f
C20162 input1/a_36_113# 0 0.418095f
C20163 _429_/a_2560_156# 0 0.016968f
C20164 _429_/a_2665_112# 0 0.62251f
C20165 _429_/a_2248_156# 0 0.371662f
C20166 _429_/a_1204_472# 0 0.012971f
C20167 _429_/a_1000_472# 0 0.291735f
C20168 _429_/a_796_472# 0 0.023206f
C20169 _429_/a_1308_423# 0 0.279043f
C20170 _429_/a_448_472# 0 0.684413f
C20171 _429_/a_36_151# 0 1.43589f
C20172 _011_ 0 0.278979f
C20173 _377_/a_36_472# 0 0.031137f
C20174 fanout66/a_36_113# 0 0.418095f
C20175 _035_ 0 0.327801f
C20176 _446_/a_2560_156# 0 0.016968f
C20177 _446_/a_2665_112# 0 0.62251f
C20178 _446_/a_2248_156# 0 0.371662f
C20179 _446_/a_1204_472# 0 0.012971f
C20180 _446_/a_1000_472# 0 0.291735f
C20181 _446_/a_796_472# 0 0.023206f
C20182 _446_/a_1308_423# 0 0.279043f
C20183 _446_/a_448_472# 0 0.684413f
C20184 _446_/a_36_151# 0 1.43589f
C20185 fanout77/a_36_113# 0 0.418095f
C20186 FILLER_0_5_212/a_36_472# 0 0.417394f
C20187 FILLER_0_5_212/a_124_375# 0 0.246306f
C20188 fanout55/a_36_160# 0 0.696445f
C20189 _175_ 0 0.344159f
C20190 _394_/a_1936_472# 0 0.009918f
C20191 _394_/a_718_524# 0 0.005143f
C20192 _394_/a_56_524# 0 0.41096f
C20193 _394_/a_728_93# 0 0.654825f
C20194 _394_/a_1336_472# 0 0.316639f
C20195 FILLER_0_3_172/a_3172_472# 0 0.345058f
C20196 FILLER_0_3_172/a_2724_472# 0 0.33241f
C20197 FILLER_0_3_172/a_2276_472# 0 0.33241f
C20198 FILLER_0_3_172/a_1828_472# 0 0.33241f
C20199 FILLER_0_3_172/a_1380_472# 0 0.33241f
C20200 FILLER_0_3_172/a_932_472# 0 0.33241f
C20201 FILLER_0_3_172/a_484_472# 0 0.33241f
C20202 FILLER_0_3_172/a_36_472# 0 0.404746f
C20203 FILLER_0_3_172/a_3260_375# 0 0.233093f
C20204 FILLER_0_3_172/a_2812_375# 0 0.17167f
C20205 FILLER_0_3_172/a_2364_375# 0 0.17167f
C20206 FILLER_0_3_172/a_1916_375# 0 0.17167f
C20207 FILLER_0_3_172/a_1468_375# 0 0.17167f
C20208 FILLER_0_3_172/a_1020_375# 0 0.17167f
C20209 FILLER_0_3_172/a_572_375# 0 0.17167f
C20210 FILLER_0_3_172/a_124_375# 0 0.185915f
C20211 FILLER_0_17_72/a_3172_472# 0 0.345058f
C20212 FILLER_0_17_72/a_2724_472# 0 0.33241f
C20213 FILLER_0_17_72/a_2276_472# 0 0.33241f
C20214 FILLER_0_17_72/a_1828_472# 0 0.33241f
C20215 FILLER_0_17_72/a_1380_472# 0 0.33241f
C20216 FILLER_0_17_72/a_932_472# 0 0.33241f
C20217 FILLER_0_17_72/a_484_472# 0 0.33241f
C20218 FILLER_0_17_72/a_36_472# 0 0.404746f
C20219 FILLER_0_17_72/a_3260_375# 0 0.233093f
C20220 FILLER_0_17_72/a_2812_375# 0 0.17167f
C20221 FILLER_0_17_72/a_2364_375# 0 0.17167f
C20222 FILLER_0_17_72/a_1916_375# 0 0.17167f
C20223 FILLER_0_17_72/a_1468_375# 0 0.17167f
C20224 FILLER_0_17_72/a_1020_375# 0 0.17167f
C20225 FILLER_0_17_72/a_572_375# 0 0.17167f
C20226 FILLER_0_17_72/a_124_375# 0 0.185915f
C20227 FILLER_0_2_93/a_484_472# 0 0.345058f
C20228 FILLER_0_2_93/a_36_472# 0 0.404746f
C20229 FILLER_0_2_93/a_572_375# 0 0.232991f
C20230 FILLER_0_2_93/a_124_375# 0 0.185089f
C20231 FILLER_0_11_142/a_484_472# 0 0.345058f
C20232 FILLER_0_11_142/a_36_472# 0 0.404746f
C20233 FILLER_0_11_142/a_572_375# 0 0.232991f
C20234 FILLER_0_11_142/a_124_375# 0 0.185089f
C20235 net25 0 1.803174f
C20236 _232_/a_67_603# 0 0.345683f
C20237 net35 0 1.844415f
C20238 mask\[8\] 0 1.276111f
C20239 _301_/a_36_472# 0 0.031137f
C20240 _033_ 0 0.323682f
C20241 _165_ 0 0.331995f
C20242 FILLER_0_3_2/a_36_472# 0 0.417394f
C20243 FILLER_0_3_2/a_124_375# 0 0.246306f
C20244 trim_val\[3\] 0 0.719615f
C20245 _036_ 0 0.369206f
C20246 net68 0 1.735004f
C20247 _447_/a_2560_156# 0 0.016968f
C20248 _447_/a_2665_112# 0 0.62251f
C20249 _447_/a_2248_156# 0 0.371662f
C20250 _447_/a_1204_472# 0 0.012971f
C20251 _447_/a_1000_472# 0 0.291735f
C20252 _447_/a_796_472# 0 0.023206f
C20253 _447_/a_1308_423# 0 0.279043f
C20254 _447_/a_448_472# 0 0.684413f
C20255 _447_/a_36_151# 0 1.43589f
C20256 FILLER_0_19_28/a_484_472# 0 0.345058f
C20257 FILLER_0_19_28/a_36_472# 0 0.404746f
C20258 FILLER_0_19_28/a_572_375# 0 0.232991f
C20259 FILLER_0_19_28/a_124_375# 0 0.185089f
C20260 fanout65/a_36_113# 0 0.418095f
C20261 fanout76/a_36_160# 0 0.386641f
C20262 net54 0 5.456963f
C20263 fanout54/a_36_160# 0 0.696445f
C20264 FILLER_0_4_49/a_484_472# 0 0.345058f
C20265 FILLER_0_4_49/a_36_472# 0 0.404746f
C20266 FILLER_0_4_49/a_572_375# 0 0.232991f
C20267 FILLER_0_4_49/a_124_375# 0 0.185089f
C20268 _176_ 0 0.804011f
C20269 _085_ 0 2.280803f
C20270 _116_ 0 1.959915f
C20271 _395_/a_36_488# 0 0.101145f
C20272 FILLER_0_14_50/a_36_472# 0 0.417394f
C20273 FILLER_0_14_50/a_124_375# 0 0.246306f
C20274 FILLER_0_8_263/a_36_472# 0 0.417394f
C20275 FILLER_0_8_263/a_124_375# 0 0.246306f
C20276 FILLER_0_0_130/a_36_472# 0 0.417394f
C20277 FILLER_0_0_130/a_124_375# 0 0.246306f
C20278 FILLER_0_16_255/a_36_472# 0 0.417394f
C20279 FILLER_0_16_255/a_124_375# 0 0.246306f
C20280 FILLER_0_7_59/a_484_472# 0 0.345058f
C20281 FILLER_0_7_59/a_36_472# 0 0.404746f
C20282 FILLER_0_7_59/a_572_375# 0 0.232991f
C20283 FILLER_0_7_59/a_124_375# 0 0.185089f
C20284 ctlp[2] 0 0.17528f
C20285 output19/a_224_472# 0 2.38465f
C20286 FILLER_0_7_146/a_36_472# 0 0.417394f
C20287 FILLER_0_7_146/a_124_375# 0 0.246306f
C20288 _216_/a_67_603# 0 0.345683f
C20289 FILLER_0_15_116/a_484_472# 0 0.345058f
C20290 FILLER_0_15_116/a_36_472# 0 0.404746f
C20291 FILLER_0_15_116/a_572_375# 0 0.232991f
C20292 FILLER_0_15_116/a_124_375# 0 0.185089f
C20293 _063_ 0 0.370155f
C20294 _233_/a_36_160# 0 0.386641f
C20295 FILLER_0_21_28/a_3172_472# 0 0.345058f
C20296 FILLER_0_21_28/a_2724_472# 0 0.33241f
C20297 FILLER_0_21_28/a_2276_472# 0 0.33241f
C20298 FILLER_0_21_28/a_1828_472# 0 0.33241f
C20299 FILLER_0_21_28/a_1380_472# 0 0.33241f
C20300 FILLER_0_21_28/a_932_472# 0 0.33241f
C20301 FILLER_0_21_28/a_484_472# 0 0.33241f
C20302 FILLER_0_21_28/a_36_472# 0 0.404746f
C20303 FILLER_0_21_28/a_3260_375# 0 0.233093f
C20304 FILLER_0_21_28/a_2812_375# 0 0.17167f
C20305 FILLER_0_21_28/a_2364_375# 0 0.17167f
C20306 FILLER_0_21_28/a_1916_375# 0 0.17167f
C20307 FILLER_0_21_28/a_1468_375# 0 0.17167f
C20308 FILLER_0_21_28/a_1020_375# 0 0.17167f
C20309 FILLER_0_21_28/a_572_375# 0 0.17167f
C20310 FILLER_0_21_28/a_124_375# 0 0.185915f
C20311 _110_ 0 0.323912f
C20312 _379_/a_36_472# 0 0.031137f
C20313 trim_val\[4\] 0 0.662409f
C20314 net76 0 1.454269f
C20315 _448_/a_2560_156# 0 0.016968f
C20316 _448_/a_2665_112# 0 0.62251f
C20317 _448_/a_2248_156# 0 0.371662f
C20318 _448_/a_1204_472# 0 0.012971f
C20319 _448_/a_1000_472# 0 0.291735f
C20320 _448_/a_796_472# 0 0.023206f
C20321 _448_/a_1308_423# 0 0.279043f
C20322 _448_/a_448_472# 0 0.684413f
C20323 _448_/a_36_151# 0 1.43589f
C20324 fanout64/a_36_160# 0 0.386641f
C20325 fanout75/a_36_113# 0 0.418095f
C20326 _250_/a_36_68# 0 0.69549f
C20327 net56 0 0.843396f
C20328 fanout53/a_36_160# 0 0.696445f
C20329 _177_ 0 0.358286f
C20330 result[2] 0 0.230851f
C20331 net29 0 1.802718f
C20332 output29/a_224_472# 0 2.38465f
C20333 ctlp[1] 0 0.17418f
C20334 output18/a_224_472# 0 2.38465f
C20335 FILLER_0_14_181/a_36_472# 0 0.417394f
C20336 FILLER_0_14_181/a_124_375# 0 0.246306f
C20337 _052_ 0 0.569133f
C20338 _217_/a_36_160# 0 0.386641f
C20339 net44 0 1.407054f
C20340 _303_/a_36_472# 0 0.031137f
C20341 en_co_clk 0 0.346872f
C20342 net55 0 5.119958f
C20343 net72 0 1.366255f
C20344 _449_/a_2560_156# 0 0.016968f
C20345 _449_/a_2665_112# 0 0.62251f
C20346 _449_/a_2248_156# 0 0.371662f
C20347 _449_/a_1204_472# 0 0.012971f
C20348 _449_/a_1000_472# 0 0.291735f
C20349 _449_/a_796_472# 0 0.023206f
C20350 _449_/a_1308_423# 0 0.279043f
C20351 _449_/a_448_472# 0 0.684413f
C20352 _449_/a_36_151# 0 1.43589f
C20353 fanout52/a_36_160# 0 0.696445f
C20354 net82 0 0.706042f
C20355 fanout74/a_36_113# 0 0.418095f
C20356 FILLER_0_10_28/a_36_472# 0 0.417394f
C20357 FILLER_0_10_28/a_124_375# 0 0.246306f
C20358 mask\[0\] 0 2.242948f
C20359 _320_/a_36_472# 0 0.137725f
C20360 fanout63/a_36_160# 0 0.696445f
C20361 FILLER_0_14_81/a_36_472# 0 0.417394f
C20362 FILLER_0_14_81/a_124_375# 0 0.246306f
C20363 _397_/a_36_472# 0 0.031137f
C20364 FILLER_0_13_212/a_1380_472# 0 0.345058f
C20365 FILLER_0_13_212/a_932_472# 0 0.33241f
C20366 FILLER_0_13_212/a_484_472# 0 0.33241f
C20367 FILLER_0_13_212/a_36_472# 0 0.404746f
C20368 FILLER_0_13_212/a_1468_375# 0 0.233029f
C20369 FILLER_0_13_212/a_1020_375# 0 0.171606f
C20370 FILLER_0_13_212/a_572_375# 0 0.171606f
C20371 FILLER_0_13_212/a_124_375# 0 0.185399f
C20372 trim[1] 0 0.793787f
C20373 net39 0 1.445128f
C20374 output39/a_224_472# 0 2.38465f
C20375 result[1] 0 0.229507f
C20376 net28 0 1.759728f
C20377 output28/a_224_472# 0 2.38465f
C20378 ctlp[0] 0 1.002286f
C20379 output17/a_224_472# 0 2.38465f
C20380 FILLER_0_16_37/a_36_472# 0 0.417394f
C20381 FILLER_0_16_37/a_124_375# 0 0.246306f
C20382 net26 0 1.671545f
C20383 _064_ 0 0.581481f
C20384 trim_val\[2\] 0 0.65354f
C20385 trim_mask\[2\] 0 0.92551f
C20386 _235_/a_67_603# 0 0.345683f
C20387 _013_ 0 0.48783f
C20388 _111_ 0 0.369652f
C20389 FILLER_0_18_177/a_3172_472# 0 0.345058f
C20390 FILLER_0_18_177/a_2724_472# 0 0.33241f
C20391 FILLER_0_18_177/a_2276_472# 0 0.33241f
C20392 FILLER_0_18_177/a_1828_472# 0 0.33241f
C20393 FILLER_0_18_177/a_1380_472# 0 0.33241f
C20394 FILLER_0_18_177/a_932_472# 0 0.33241f
C20395 FILLER_0_18_177/a_484_472# 0 0.33241f
C20396 FILLER_0_18_177/a_36_472# 0 0.404746f
C20397 FILLER_0_18_177/a_3260_375# 0 0.233093f
C20398 FILLER_0_18_177/a_2812_375# 0 0.17167f
C20399 FILLER_0_18_177/a_2364_375# 0 0.17167f
C20400 FILLER_0_18_177/a_1916_375# 0 0.17167f
C20401 FILLER_0_18_177/a_1468_375# 0 0.17167f
C20402 FILLER_0_18_177/a_1020_375# 0 0.17167f
C20403 FILLER_0_18_177/a_572_375# 0 0.17167f
C20404 FILLER_0_18_177/a_124_375# 0 0.185915f
C20405 FILLER_0_18_100/a_36_472# 0 0.417394f
C20406 FILLER_0_18_100/a_124_375# 0 0.246306f
C20407 _073_ 0 0.953711f
C20408 _126_ 0 2.036767f
C20409 _069_ 0 2.034557f
C20410 _321_/a_170_472# 0 0.077257f
C20411 fanout51/a_36_113# 0 0.418095f
C20412 net62 0 4.932099f
C20413 fanout62/a_36_160# 0 0.696445f
C20414 fanout73/a_36_113# 0 0.418095f
C20415 FILLER_0_19_47/a_484_472# 0 0.345058f
C20416 FILLER_0_19_47/a_36_472# 0 0.404746f
C20417 FILLER_0_19_47/a_572_375# 0 0.232991f
C20418 FILLER_0_19_47/a_124_375# 0 0.185089f
C20419 FILLER_0_14_91/a_484_472# 0 0.345058f
C20420 FILLER_0_14_91/a_36_472# 0 0.404746f
C20421 FILLER_0_14_91/a_572_375# 0 0.232991f
C20422 FILLER_0_14_91/a_124_375# 0 0.185089f
C20423 FILLER_0_10_214/a_36_472# 0 0.417394f
C20424 FILLER_0_10_214/a_124_375# 0 0.246306f
C20425 FILLER_0_10_247/a_36_472# 0 0.417394f
C20426 FILLER_0_10_247/a_124_375# 0 0.246306f
C20427 _178_ 0 1.252435f
C20428 _398_/a_36_113# 0 0.418095f
C20429 FILLER_0_16_241/a_36_472# 0 0.417394f
C20430 FILLER_0_16_241/a_124_375# 0 0.246306f
C20431 trim[0] 0 0.796081f
C20432 net38 0 1.529392f
C20433 output38/a_224_472# 0 2.38465f
C20434 ctln[9] 0 0.904836f
C20435 net16 0 1.295744f
C20436 output16/a_224_472# 0 2.38465f
C20437 result[0] 0 0.56622f
C20438 output27/a_224_472# 0 2.38465f
C20439 _219_/a_36_160# 0 0.386641f
C20440 FILLER_0_20_193/a_484_472# 0 0.345058f
C20441 FILLER_0_20_193/a_36_472# 0 0.404746f
C20442 FILLER_0_20_193/a_572_375# 0 0.232991f
C20443 FILLER_0_20_193/a_124_375# 0 0.185089f
C20444 _236_/a_36_160# 0 0.696445f
C20445 _112_ 0 0.308886f
C20446 _305_/a_36_159# 0 0.374116f
C20447 _074_ 0 1.813232f
C20448 _253_/a_36_68# 0 0.061249f
C20449 net50 0 4.486121f
C20450 net52 0 3.536016f
C20451 fanout50/a_36_160# 0 0.696445f
C20452 FILLER_0_10_37/a_36_472# 0 0.417394f
C20453 FILLER_0_10_37/a_124_375# 0 0.246306f
C20454 fanout72/a_36_113# 0 0.418095f
C20455 fanout61/a_36_113# 0 0.418095f
C20456 _128_ 0 0.447252f
C20457 _127_ 0 1.291729f
C20458 _322_/a_848_380# 0 0.40208f
C20459 _322_/a_124_24# 0 0.591898f
C20460 _088_ 0 0.457961f
C20461 _079_ 0 1.114894f
C20462 _087_ 0 0.601674f
C20463 _270_/a_36_472# 0 0.031137f
C20464 FILLER_0_4_123/a_36_472# 0 0.417394f
C20465 FILLER_0_4_123/a_124_375# 0 0.246306f
C20466 FILLER_0_17_218/a_484_472# 0 0.345058f
C20467 FILLER_0_17_218/a_36_472# 0 0.404746f
C20468 FILLER_0_17_218/a_572_375# 0 0.232991f
C20469 FILLER_0_17_218/a_124_375# 0 0.185089f
C20470 sample 0 0.508149f
C20471 output37/a_224_472# 0 2.38465f
C20472 valid 0 0.272072f
C20473 net48 0 1.219262f
C20474 output48/a_224_472# 0 2.38465f
C20475 ctln[8] 0 1.547984f
C20476 net15 0 1.440851f
C20477 output15/a_224_472# 0 2.38465f
C20478 ctlp[9] 0 0.73349f
C20479 output26/a_224_472# 0 2.38465f
C20480 FILLER_0_16_57/a_1380_472# 0 0.345058f
C20481 FILLER_0_16_57/a_932_472# 0 0.33241f
C20482 FILLER_0_16_57/a_484_472# 0 0.33241f
C20483 FILLER_0_16_57/a_36_472# 0 0.404746f
C20484 FILLER_0_16_57/a_1468_375# 0 0.233029f
C20485 FILLER_0_16_57/a_1020_375# 0 0.171606f
C20486 FILLER_0_16_57/a_572_375# 0 0.171606f
C20487 FILLER_0_16_57/a_124_375# 0 0.185399f
C20488 _306_/a_36_68# 0 0.69549f
C20489 _072_ 0 2.604301f
C20490 fanout82/a_36_113# 0 0.418095f
C20491 _015_ 0 0.406653f
C20492 _323_/a_36_113# 0 0.418095f
C20493 net60 0 5.024503f
C20494 net61 0 1.666523f
C20495 fanout60/a_36_160# 0 0.696445f
C20496 fanout71/a_36_113# 0 0.418095f
C20497 FILLER_0_6_239/a_36_472# 0 0.417394f
C20498 FILLER_0_6_239/a_124_375# 0 0.246306f
C20499 FILLER_0_4_99/a_36_472# 0 0.417394f
C20500 FILLER_0_4_99/a_124_375# 0 0.246306f
C20501 net57 0 1.383718f
C20502 FILLER_0_10_256/a_36_472# 0 0.417394f
C20503 FILLER_0_10_256/a_124_375# 0 0.246306f
C20504 cal_itt\[3\] 0 1.854962f
C20505 _340_/a_36_160# 0 0.386641f
C20506 FILLER_0_4_177/a_484_472# 0 0.345058f
C20507 FILLER_0_4_177/a_36_472# 0 0.404746f
C20508 FILLER_0_4_177/a_572_375# 0 0.232991f
C20509 FILLER_0_4_177/a_124_375# 0 0.185089f
C20510 FILLER_0_4_144/a_484_472# 0 0.345058f
C20511 FILLER_0_4_144/a_36_472# 0 0.404746f
C20512 FILLER_0_4_144/a_572_375# 0 0.232991f
C20513 FILLER_0_4_144/a_124_375# 0 0.185089f
C20514 ctln[7] 0 1.265946f
C20515 output14/a_224_472# 0 2.38465f
C20516 result[9] 0 0.8197f
C20517 output36/a_224_472# 0 2.38465f
C20518 trimb[4] 0 0.752332f
C20519 output47/a_224_472# 0 2.38465f
C20520 ctlp[8] 0 1.136333f
C20521 output25/a_224_472# 0 2.38465f
C20522 FILLER_0_12_136/a_1380_472# 0 0.345058f
C20523 FILLER_0_12_136/a_932_472# 0 0.33241f
C20524 FILLER_0_12_136/a_484_472# 0 0.33241f
C20525 FILLER_0_12_136/a_36_472# 0 0.404746f
C20526 FILLER_0_12_136/a_1468_375# 0 0.233029f
C20527 FILLER_0_12_136/a_1020_375# 0 0.171606f
C20528 FILLER_0_12_136/a_572_375# 0 0.171606f
C20529 FILLER_0_12_136/a_124_375# 0 0.185399f
C20530 FILLER_0_16_89/a_1380_472# 0 0.345058f
C20531 FILLER_0_16_89/a_932_472# 0 0.33241f
C20532 FILLER_0_16_89/a_484_472# 0 0.33241f
C20533 FILLER_0_16_89/a_36_472# 0 0.404746f
C20534 FILLER_0_16_89/a_1468_375# 0 0.233029f
C20535 FILLER_0_16_89/a_1020_375# 0 0.171606f
C20536 FILLER_0_16_89/a_572_375# 0 0.171606f
C20537 FILLER_0_16_89/a_124_375# 0 0.185399f
C20538 FILLER_0_21_125/a_484_472# 0 0.345058f
C20539 FILLER_0_21_125/a_36_472# 0 0.404746f
C20540 FILLER_0_21_125/a_572_375# 0 0.232991f
C20541 FILLER_0_21_125/a_124_375# 0 0.185089f
C20542 _238_/a_67_603# 0 0.345683f
C20543 _096_ 0 2.205532f
C20544 _093_ 0 1.893313f
C20545 FILLER_0_19_55/a_36_472# 0 0.417394f
C20546 FILLER_0_19_55/a_124_375# 0 0.246306f
C20547 net81 0 1.738987f
C20548 fanout81/a_36_160# 0 0.386641f
C20549 _057_ 0 1.600886f
C20550 _255_/a_224_552# 0 1.31114f
C20551 net73 0 1.058857f
C20552 fanout70/a_36_113# 0 0.418095f
C20553 _003_ 0 0.3064f
C20554 _089_ 0 0.36777f
C20555 _272_/a_36_472# 0 0.031137f
C20556 _187_ 0 0.311229f
C20557 _410_/a_36_68# 0 0.112263f
C20558 _141_ 0 1.249289f
C20559 mask\[3\] 0 1.26722f
C20560 _341_/a_49_472# 0 0.054843f
C20561 cal 0 0.793393f
C20562 FILLER_0_7_195/a_36_472# 0 0.417394f
C20563 FILLER_0_7_195/a_124_375# 0 0.246306f
C20564 FILLER_0_7_162/a_36_472# 0 0.417394f
C20565 FILLER_0_7_162/a_124_375# 0 0.246306f
C20566 ctln[6] 0 1.451644f
C20567 output13/a_224_472# 0 2.38465f
C20568 FILLER_0_18_2/a_3172_472# 0 0.345058f
C20569 FILLER_0_18_2/a_2724_472# 0 0.33241f
C20570 FILLER_0_18_2/a_2276_472# 0 0.33241f
C20571 FILLER_0_18_2/a_1828_472# 0 0.33241f
C20572 FILLER_0_18_2/a_1380_472# 0 0.33241f
C20573 FILLER_0_18_2/a_932_472# 0 0.33241f
C20574 FILLER_0_18_2/a_484_472# 0 0.33241f
C20575 FILLER_0_18_2/a_36_472# 0 0.404746f
C20576 FILLER_0_18_2/a_3260_375# 0 0.233093f
C20577 FILLER_0_18_2/a_2812_375# 0 0.17167f
C20578 FILLER_0_18_2/a_2364_375# 0 0.17167f
C20579 FILLER_0_18_2/a_1916_375# 0 0.17167f
C20580 FILLER_0_18_2/a_1468_375# 0 0.17167f
C20581 FILLER_0_18_2/a_1020_375# 0 0.17167f
C20582 FILLER_0_18_2/a_572_375# 0 0.17167f
C20583 FILLER_0_18_2/a_124_375# 0 0.185915f
C20584 trimb[3] 0 0.34698f
C20585 net46 0 1.13395f
C20586 output46/a_224_472# 0 2.38465f
C20587 result[8] 0 0.68837f
C20588 output35/a_224_472# 0 2.38465f
C20589 ctlp[7] 0 0.83567f
C20590 output24/a_224_472# 0 2.38465f
C20591 FILLER_0_8_107/a_36_472# 0 0.417394f
C20592 FILLER_0_8_107/a_124_375# 0 0.246306f
C20593 FILLER_0_12_124/a_36_472# 0 0.417394f
C20594 FILLER_0_12_124/a_124_375# 0 0.246306f
C20595 net41 0 1.746759f
C20596 _065_ 0 0.523724f
C20597 _239_/a_36_160# 0 0.696445f
C20598 FILLER_0_1_98/a_36_472# 0 0.417394f
C20599 FILLER_0_1_98/a_124_375# 0 0.246306f
C20600 _115_ 0 1.281516f
C20601 _114_ 0 2.293579f
C20602 _308_/a_848_380# 0 0.40208f
C20603 _308_/a_124_24# 0 0.591898f
C20604 _256_/a_36_68# 0 0.063181f
C20605 FILLER_0_10_78/a_1380_472# 0 0.345058f
C20606 FILLER_0_10_78/a_932_472# 0 0.33241f
C20607 FILLER_0_10_78/a_484_472# 0 0.33241f
C20608 FILLER_0_10_78/a_36_472# 0 0.404746f
C20609 FILLER_0_10_78/a_1468_375# 0 0.233029f
C20610 FILLER_0_10_78/a_1020_375# 0 0.171606f
C20611 FILLER_0_10_78/a_572_375# 0 0.171606f
C20612 FILLER_0_10_78/a_124_375# 0 0.185399f
C20613 _130_ 0 0.304085f
C20614 net80 0 1.375599f
C20615 fanout80/a_36_113# 0 0.418095f
C20616 net58 0 5.308423f
C20617 _000_ 0 0.382358f
C20618 net75 0 1.474299f
C20619 _411_/a_2560_156# 0 0.016968f
C20620 _411_/a_2665_112# 0 0.62251f
C20621 _411_/a_2248_156# 0 0.371662f
C20622 _411_/a_1204_472# 0 0.012971f
C20623 _411_/a_1000_472# 0 0.291735f
C20624 _411_/a_796_472# 0 0.023206f
C20625 _411_/a_1308_423# 0 0.279043f
C20626 _411_/a_448_472# 0 0.684413f
C20627 _411_/a_36_151# 0 1.43589f
C20628 state\[0\] 0 0.680109f
C20629 _273_/a_36_68# 0 0.69549f
C20630 _142_ 0 0.324372f
C20631 FILLER_0_9_223/a_484_472# 0 0.345058f
C20632 FILLER_0_9_223/a_36_472# 0 0.404746f
C20633 FILLER_0_9_223/a_572_375# 0 0.232991f
C20634 FILLER_0_9_223/a_124_375# 0 0.185089f
C20635 FILLER_0_4_197/a_1380_472# 0 0.345058f
C20636 FILLER_0_4_197/a_932_472# 0 0.33241f
C20637 FILLER_0_4_197/a_484_472# 0 0.33241f
C20638 FILLER_0_4_197/a_36_472# 0 0.404746f
C20639 FILLER_0_4_197/a_1468_375# 0 0.233029f
C20640 FILLER_0_4_197/a_1020_375# 0 0.171606f
C20641 FILLER_0_4_197/a_572_375# 0 0.171606f
C20642 FILLER_0_4_197/a_124_375# 0 0.185399f
C20643 FILLER_0_17_226/a_36_472# 0 0.417394f
C20644 FILLER_0_17_226/a_124_375# 0 0.246306f
C20645 FILLER_0_5_109/a_484_472# 0 0.345058f
C20646 FILLER_0_5_109/a_36_472# 0 0.404746f
C20647 FILLER_0_5_109/a_572_375# 0 0.232991f
C20648 FILLER_0_5_109/a_124_375# 0 0.185089f
C20649 ctln[5] 0 1.585113f
C20650 output12/a_224_472# 0 2.38465f
C20651 result[7] 0 0.24756f
C20652 net34 0 1.724665f
C20653 output34/a_224_472# 0 2.38465f
C20654 trimb[2] 0 0.839614f
C20655 net45 0 1.12041f
C20656 output45/a_224_472# 0 2.38465f
C20657 ctlp[6] 0 1.243017f
C20658 output23/a_224_472# 0 2.38465f
C20659 FILLER_0_15_142/a_484_472# 0 0.345058f
C20660 FILLER_0_15_142/a_36_472# 0 0.404746f
C20661 FILLER_0_15_142/a_572_375# 0 0.232991f
C20662 FILLER_0_15_142/a_124_375# 0 0.185089f
C20663 _077_ 0 1.645892f
C20664 _075_ 0 0.374516f
C20665 _257_/a_36_472# 0 0.031137f
C20666 _326_/a_36_160# 0 0.696445f
C20667 _412_/a_2560_156# 0 0.016968f
C20668 _412_/a_2665_112# 0 0.62251f
C20669 _412_/a_2248_156# 0 0.371662f
C20670 _412_/a_1204_472# 0 0.012971f
C20671 _412_/a_1000_472# 0 0.291735f
C20672 _412_/a_796_472# 0 0.023206f
C20673 _412_/a_1308_423# 0 0.279043f
C20674 _412_/a_448_472# 0 0.684413f
C20675 _412_/a_36_151# 0 1.43589f
C20676 _091_ 0 1.841339f
C20677 _274_/a_36_68# 0 0.063181f
C20678 _143_ 0 0.329289f
C20679 mask\[4\] 0 1.300438f
C20680 _343_/a_49_472# 0 0.054843f
C20681 FILLER_0_13_65/a_36_472# 0 0.417394f
C20682 FILLER_0_13_65/a_124_375# 0 0.246306f
C20683 _360_/a_36_160# 0 0.386641f
C20684 FILLER_0_4_185/a_36_472# 0 0.417394f
C20685 FILLER_0_4_185/a_124_375# 0 0.246306f
C20686 FILLER_0_4_152/a_36_472# 0 0.417394f
C20687 FILLER_0_4_152/a_124_375# 0 0.246306f
C20688 _291_/a_36_160# 0 0.386641f
C20689 ctln[2] 0 1.833091f
C20690 output9/a_224_472# 0 2.38465f
C20691 ctln[4] 0 1.461847f
C20692 output11/a_224_472# 0 2.38465f
C20693 trimb[1] 0 0.378532f
C20694 output44/a_224_472# 0 2.38465f
C20695 result[6] 0 0.19512f
C20696 output33/a_224_472# 0 2.38465f
C20697 ctlp[5] 0 1.282822f
C20698 output22/a_224_472# 0 2.38465f
C20699 FILLER_0_8_127/a_36_472# 0 0.417394f
C20700 FILLER_0_8_127/a_124_375# 0 0.246306f
C20701 FILLER_0_8_138/a_36_472# 0 0.417394f
C20702 FILLER_0_8_138/a_124_375# 0 0.246306f
C20703 FILLER_0_21_133/a_36_472# 0 0.417394f
C20704 FILLER_0_21_133/a_124_375# 0 0.246306f
C20705 FILLER_0_24_130/a_36_472# 0 0.417394f
C20706 FILLER_0_24_130/a_124_375# 0 0.246306f
C20707 FILLER_0_18_171/a_36_472# 0 0.417394f
C20708 FILLER_0_18_171/a_124_375# 0 0.246306f
C20709 _258_/a_36_160# 0 0.386641f
C20710 _016_ 0 0.314121f
C20711 _327_/a_36_472# 0 0.031137f
C20712 _189_/a_67_603# 0 0.345683f
C20713 FILLER_0_24_63/a_36_472# 0 0.417394f
C20714 FILLER_0_24_63/a_124_375# 0 0.246306f
C20715 FILLER_0_24_96/a_36_472# 0 0.417394f
C20716 FILLER_0_24_96/a_124_375# 0 0.246306f
C20717 cal_itt\[2\] 0 1.473514f
C20718 _002_ 0 0.289553f
C20719 _413_/a_2560_156# 0 0.016968f
C20720 _413_/a_2665_112# 0 0.62251f
C20721 _413_/a_2248_156# 0 0.371662f
C20722 _413_/a_1204_472# 0 0.012971f
C20723 _413_/a_1000_472# 0 0.291735f
C20724 _413_/a_796_472# 0 0.023206f
C20725 _413_/a_1308_423# 0 0.279043f
C20726 _413_/a_448_472# 0 0.684413f
C20727 _413_/a_36_151# 0 1.43589f
C20728 _092_ 0 0.680239f
C20729 FILLER_0_7_72/a_3172_472# 0 0.345058f
C20730 FILLER_0_7_72/a_2724_472# 0 0.33241f
C20731 FILLER_0_7_72/a_2276_472# 0 0.33241f
C20732 FILLER_0_7_72/a_1828_472# 0 0.33241f
C20733 FILLER_0_7_72/a_1380_472# 0 0.33241f
C20734 FILLER_0_7_72/a_932_472# 0 0.33241f
C20735 FILLER_0_7_72/a_484_472# 0 0.33241f
C20736 FILLER_0_7_72/a_36_472# 0 0.404746f
C20737 FILLER_0_7_72/a_3260_375# 0 0.233093f
C20738 FILLER_0_7_72/a_2812_375# 0 0.17167f
C20739 FILLER_0_7_72/a_2364_375# 0 0.17167f
C20740 FILLER_0_7_72/a_1916_375# 0 0.17167f
C20741 FILLER_0_7_72/a_1468_375# 0 0.17167f
C20742 FILLER_0_7_72/a_1020_375# 0 0.17167f
C20743 FILLER_0_7_72/a_572_375# 0 0.17167f
C20744 FILLER_0_7_72/a_124_375# 0 0.185915f
C20745 _086_ 0 2.45259f
C20746 _119_ 0 1.237181f
C20747 net63 0 5.362473f
C20748 _430_/a_2560_156# 0 0.016968f
C20749 _430_/a_2665_112# 0 0.62251f
C20750 _430_/a_2248_156# 0 0.371662f
C20751 _430_/a_1204_472# 0 0.012971f
C20752 _430_/a_1000_472# 0 0.291735f
C20753 _430_/a_796_472# 0 0.023206f
C20754 _430_/a_1308_423# 0 0.279043f
C20755 _430_/a_448_472# 0 0.684413f
C20756 _430_/a_36_151# 0 1.43589f
C20757 _292_/a_36_160# 0 0.386641f
C20758 comp 0 1.022965f
C20759 ctln[1] 0 1.11973f
C20760 output8/a_224_472# 0 2.38465f
C20761 ctln[3] 0 0.835391f
C20762 output10/a_224_472# 0 2.38465f
C20763 result[5] 0 0.206867f
C20764 net32 0 1.78884f
C20765 output32/a_224_472# 0 2.38465f
C20766 trimb[0] 0 0.847787f
C20767 output43/a_224_472# 0 2.38465f
C20768 ctlp[4] 0 0.37565f
C20769 output21/a_224_472# 0 2.38465f
C20770 _053_ 0 1.705161f
C20771 FILLER_0_16_107/a_484_472# 0 0.345058f
C20772 FILLER_0_16_107/a_36_472# 0 0.404746f
C20773 FILLER_0_16_107/a_572_375# 0 0.232991f
C20774 FILLER_0_16_107/a_124_375# 0 0.185089f
C20775 FILLER_0_3_204/a_36_472# 0 0.417394f
C20776 FILLER_0_3_204/a_124_375# 0 0.246306f
C20777 FILLER_0_9_28/a_3172_472# 0 0.345058f
C20778 FILLER_0_9_28/a_2724_472# 0 0.33241f
C20779 FILLER_0_9_28/a_2276_472# 0 0.33241f
C20780 FILLER_0_9_28/a_1828_472# 0 0.33241f
C20781 FILLER_0_9_28/a_1380_472# 0 0.33241f
C20782 FILLER_0_9_28/a_932_472# 0 0.33241f
C20783 FILLER_0_9_28/a_484_472# 0 0.33241f
C20784 FILLER_0_9_28/a_36_472# 0 0.404746f
C20785 FILLER_0_9_28/a_3260_375# 0 0.233093f
C20786 FILLER_0_9_28/a_2812_375# 0 0.17167f
C20787 FILLER_0_9_28/a_2364_375# 0 0.17167f
C20788 FILLER_0_9_28/a_1916_375# 0 0.17167f
C20789 FILLER_0_9_28/a_1468_375# 0 0.17167f
C20790 FILLER_0_9_28/a_1020_375# 0 0.17167f
C20791 FILLER_0_9_28/a_572_375# 0 0.17167f
C20792 FILLER_0_9_28/a_124_375# 0 0.185915f
C20793 _132_ 0 1.491425f
C20794 _328_/a_36_113# 0 0.418095f
C20795 _414_/a_2560_156# 0 0.016968f
C20796 _414_/a_2665_112# 0 0.62251f
C20797 _414_/a_2248_156# 0 0.371662f
C20798 _414_/a_1204_472# 0 0.012971f
C20799 _414_/a_1000_472# 0 0.291735f
C20800 _414_/a_796_472# 0 0.023206f
C20801 _414_/a_1308_423# 0 0.279043f
C20802 _414_/a_448_472# 0 0.684413f
C20803 _414_/a_36_151# 0 1.43589f
C20804 _276_/a_36_160# 0 0.386641f
C20805 _144_ 0 1.173846f
C20806 _345_/a_36_160# 0 0.386641f
C20807 _155_ 0 0.638535f
C20808 _020_ 0 0.316793f
C20809 _431_/a_2560_156# 0 0.016968f
C20810 _431_/a_2665_112# 0 0.62251f
C20811 _431_/a_2248_156# 0 0.371662f
C20812 _431_/a_1204_472# 0 0.012971f
C20813 _431_/a_1000_472# 0 0.291735f
C20814 _431_/a_796_472# 0 0.023206f
C20815 _431_/a_1308_423# 0 0.279043f
C20816 _431_/a_448_472# 0 0.684413f
C20817 _431_/a_36_151# 0 1.43589f
C20818 _105_ 0 1.21281f
C20819 _293_/a_36_472# 0 0.031137f
C20820 FILLER_0_5_128/a_484_472# 0 0.345058f
C20821 FILLER_0_5_128/a_36_472# 0 0.404746f
C20822 FILLER_0_5_128/a_572_375# 0 0.232991f
C20823 FILLER_0_5_128/a_124_375# 0 0.185089f
C20824 FILLER_0_5_117/a_36_472# 0 0.417394f
C20825 FILLER_0_5_117/a_124_375# 0 0.246306f
C20826 ctln[0] 0 1.423102f
C20827 net7 0 1.174913f
C20828 output7/a_224_472# 0 2.38465f
C20829 trim[4] 0 0.763069f
C20830 output42/a_224_472# 0 2.38465f
C20831 result[4] 0 0.038878f
C20832 net31 0 1.912935f
C20833 output31/a_224_472# 0 2.38465f
C20834 ctlp[3] 0 1.14968f
C20835 output20/a_224_472# 0 2.38465f
C20836 FILLER_0_16_73/a_484_472# 0 0.345058f
C20837 FILLER_0_16_73/a_36_472# 0 0.404746f
C20838 FILLER_0_16_73/a_572_375# 0 0.232991f
C20839 FILLER_0_16_73/a_124_375# 0 0.185089f
C20840 FILLER_0_21_142/a_484_472# 0 0.345058f
C20841 FILLER_0_21_142/a_36_472# 0 0.404746f
C20842 FILLER_0_21_142/a_572_375# 0 0.232991f
C20843 FILLER_0_21_142/a_124_375# 0 0.185089f
C20844 FILLER_0_15_150/a_36_472# 0 0.417394f
C20845 FILLER_0_15_150/a_124_375# 0 0.246306f
C20846 FILLER_0_19_125/a_36_472# 0 0.417394f
C20847 FILLER_0_19_125/a_124_375# 0 0.246306f
C20848 net10 0 1.480101f
C20849 net20 0 2.034189f
C20850 _277_/a_36_160# 0 0.386641f
C20851 net27 0 2.023744f
C20852 _004_ 0 0.390107f
C20853 _415_/a_2560_156# 0 0.016968f
C20854 _415_/a_2665_112# 0 0.62251f
C20855 _415_/a_2248_156# 0 0.371662f
C20856 _415_/a_1204_472# 0 0.012971f
C20857 _415_/a_1000_472# 0 0.291735f
C20858 _415_/a_796_472# 0 0.023206f
C20859 _415_/a_1308_423# 0 0.279043f
C20860 _415_/a_448_472# 0 0.684413f
C20861 _415_/a_36_151# 0 1.43589f
C20862 mask\[5\] 0 1.334568f
C20863 _346_/a_49_472# 0 0.054843f
C20864 _028_ 0 0.386029f
C20865 _363_/a_36_68# 0 0.150048f
C20866 _021_ 0 0.316776f
C20867 _432_/a_2560_156# 0 0.016968f
C20868 _432_/a_2665_112# 0 0.62251f
C20869 _432_/a_2248_156# 0 0.371662f
C20870 _432_/a_1204_472# 0 0.012971f
C20871 _432_/a_1000_472# 0 0.291735f
C20872 _432_/a_796_472# 0 0.023206f
C20873 _432_/a_1308_423# 0 0.279043f
C20874 _432_/a_448_472# 0 0.684413f
C20875 _432_/a_36_151# 0 1.43589f
C20876 _008_ 0 0.423631f
C20877 _104_ 0 1.435764f
C20878 _106_ 0 0.378703f
C20879 FILLER_0_17_200/a_484_472# 0 0.345058f
C20880 FILLER_0_17_200/a_36_472# 0 0.404746f
C20881 FILLER_0_17_200/a_572_375# 0 0.232991f
C20882 FILLER_0_17_200/a_124_375# 0 0.185089f
.ends

.subckt saradc vdd vss vinp vinn result[0] result[1] result[2] result[3] result[4]
+ result[5] result[6] result[7] result[8] result[9] valid cal en clk rstn
Xlatch_0 latch_0/tutyuu1 latch_0/tutyuu2 latch_0/Qn latch_0/Q latch_0/S latch_0/R
+ vdd vss latch
Xbuffer_0 buffer_0/middle buffer_0/out buffer_0/in vdd vss buffer_0/buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162#
+ buffer
Xdacp_0 vdd dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9 dacp_0/ctl10 vinp dacp_0/sample dacp_0/ctl2
+ dacp_0/ctl1 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/ndum dacp_0/ctl4 dacp_0/ctl6
+ dacp_0/bootstrapped_sw_p_0/enb dacp_0/out dacp_0/bootstrapped_sw_p_0/vbsl dacp_0/ctl3
+ dacp_0/bootstrapped_sw_p_0/vg dacp_0/bootstrapped_sw_p_0/vbsh dacp_0/carray_p_0/n8
+ dacp_0/carray_p_0/n9 dacp_0/ctl5 vdd vss dacp
Xcomparator_0 vdd dacp_0/out dacn_0/out sarlogic_0/trim[4] sarlogic_0/trim[1] sarlogic_0/trim[0]
+ sarlogic_0/trimb[4] sarlogic_0/trimb[1] sarlogic_0/trimb[0] sarlogic_0/trimb[2]
+ sarlogic_0/trimb[3] comparator_0/diff comparator_0/in comparator_0/trim_right_0/trim_switch_right_0/XM2_trim_right_0/D
+ comparator_0/trim_right_0/trim_switch_right_0/XM3_trim_right_0/D buffer_0/out comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D
+ latch_0/S latch_0/R comparator_0/trim_left_0/trim_switch_left_0/n4 comparator_0/trim_left_0/trim_switch_left_0/n3
+ comparator_0/trim_left_0/trim_switch_left_0/n2 comparator_0/ip sarlogic_0/trim[3]
+ sarlogic_0/trim[2] vss comparator
Xdacn_0 dacn_0/ctl1 dacn_0/ctl2 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5 dacn_0/ctl6 dacn_0/ctl7
+ dacn_0/ctl8 dacn_0/ctl9 dacn_0/ctl10 vinn dacn_0/bootstrapped_sw_n_0/vg dacn_0/bootstrapped_sw_n_0/enb
+ dacn_0/carray_n_0/n9 dacp_0/sample dacn_0/carray_n_0/n0 dacn_0/out dacn_0/carray_n_0/n8
+ vdd vdd dacn_0/bootstrapped_sw_n_0/vbsh vss dacn_0/bootstrapped_sw_n_0/vbsl dacn_0/carray_n_0/ndum
+ dacn
Xmim_cap_boss_0 vss vdd vss mim_cap_boss
Xsarlogic_0 dacn_0/ctl10 dacn_0/ctl1 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5 dacn_0/ctl6
+ dacn_0/ctl8 dacp_0/ctl10 dacp_0/ctl1 dacp_0/ctl2 dacp_0/ctl3 dacp_0/ctl4 dacp_0/ctl5
+ dacp_0/ctl6 dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9 clk buffer_0/in latch_0/Q en result[0]
+ result[1] result[2] result[3] result[4] result[5] result[6] result[7] result[8]
+ result[9] rstn dacp_0/sample sarlogic_0/trim[0] sarlogic_0/trim[1] sarlogic_0/trim[2]
+ sarlogic_0/trim[3] sarlogic_0/trim[4] sarlogic_0/trimb[0] sarlogic_0/trimb[1] sarlogic_0/trimb[2]
+ sarlogic_0/trimb[3] sarlogic_0/trimb[4] valid sarlogic_0/net10 sarlogic_0/output13/a_224_472#
+ sarlogic_0/output23/a_224_472# sarlogic_0/net59 sarlogic_0/net16 sarlogic_0/net27
+ sarlogic_0/output25/a_224_472# sarlogic_0/cal_itt\[1\] sarlogic_0/fanout65/a_36_113#
+ dacn_0/ctl2 dacn_0/ctl7 sarlogic_0/net15 dacn_0/ctl9 sarlogic_0/output10/a_224_472#
+ sarlogic_0/net26 sarlogic_0/net24 sarlogic_0/output11/a_224_472# sarlogic_0/output21/a_224_472#
+ sarlogic_0/net14 sarlogic_0/output12/a_224_472# sarlogic_0/output22/a_224_472# cal
+ sarlogic_0/net62 sarlogic_0/net20 vss vdd sarlogic
Xmim_cap_boss_1 vss vdd vss mim_cap_boss
C0 sarlogic_0/trim[1] vdd 0.113951f
C1 sarlogic_0/trim[4] sarlogic_0/trim[1] 2.925859f
C2 comparator_0/ip comparator_0/trim_right_0/trim_switch_right_0/XM2_trim_right_0/D 3.21246f
C3 sarlogic_0/net62 dacp_0/sample 0.160765f
C4 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n6 11.2161f
C5 dacp_0/sample sarlogic_0/fanout65/a_36_113# 0.001365f
C6 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n5 3.36878f
C7 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/n1 8.469265f
C8 latch_0/S latch_0/tutyuu1 0.005228f
C9 valid vdd 3.413481f
C10 dacn_0/ctl9 vdd 0.593962f
C11 dacp_0/carray_p_0/n9 dacp_0/out 0.846152p
C12 comparator_0/trim_right_0/trim_switch_right_0/XM3_trim_right_0/D vdd 0.248007f
C13 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/ndum 0.127951f
C14 dacp_0/ctl7 vdd 0.444612f
C15 dacp_0/sample sarlogic_0/cal_itt\[1\] 0.004307f
C16 dacp_0/bootstrapped_sw_p_0/vg vdd 0.026792f
C17 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n0 0.051666f
C18 dacp_0/ctl8 dacp_0/ctl7 2.592389f
C19 dacn_0/bootstrapped_sw_n_0/vg vdd 0.026792f
C20 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n4 2.84323f
C21 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D comparator_0/trim_right_0/trim_switch_right_0/XM0_trim_right_0/D 0.032158f
C22 dacp_0/carray_p_0/n8 vdd 0.031782f
C23 dacp_0/ctl9 dacp_0/ctl10 2.076966f
C24 dacn_0/carray_n_0/n3 dacn_0/carray_n_0/n1 0.137399f
C25 sarlogic_0/output22/a_224_472# vdd 0.006461f
C26 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n3 0.336612f
C27 dacn_0/bootstrapped_sw_n_0/vbsh dacn_0/out -0.061493f
C28 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n1 0.137399f
C29 m5_121216_n195240# vdd 1.18282f
C30 dacn_0/carray_n_0/n0 dacn_0/carray_n_0/n1 8.469265f
C31 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n0 0.025424f
C32 dacn_0/ctl8 vdd 0.393337f
C33 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n0 0.025424f
C34 dacn_0/out dacn_0/carray_n_0/n1 3.365905f
C35 dacn_0/carray_n_0/n8 vdd 0.031782f
C36 dacn_0/carray_n_0/n1 dacn_0/carray_n_0/n9 0.342393f
C37 comparator_0/ip vdd 0.39079f
C38 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n1 0.134826f
C39 dacn_0/carray_n_0/n6 dacn_0/out 0.105055p
C40 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/ndum 0.097254f
C41 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n9 14.716781f
C42 dacp_0/out dacp_0/carray_p_0/n8 0.420152p
C43 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n2 0.485242f
C44 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n6 0.614078f
C45 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n1 0.134705f
C46 result[7] result[8] 3.472163f
C47 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/ndum 0.097254f
C48 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n6 28.589401f
C49 dacn_0/ctl7 vdd 0.448862f
C50 dacp_0/ctl4 dacp_0/ctl3 3.636019f
C51 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/ndum 0.041162f
C52 sarlogic_0/trim[0] sarlogic_0/trim[1] 2.987179f
C53 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n1 0.134562f
C54 dacp_0/sample result[8] 0.161003f
C55 dacp_0/ctl9 vdd 0.673812f
C56 comparator_0/in buffer_0/out 0.016561f
C57 comparator_0/trim_left_0/trim_switch_left_0/n2 comparator_0/in 3.21246f
C58 dacp_0/ctl9 dacp_0/ctl8 2.331489f
C59 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n0 0.040502f
C60 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n5 7.39935f
C61 sarlogic_0/output12/a_224_472# vdd 0.006182f
C62 m5_n124784_86040# vdd 1.18282f
C63 sarlogic_0/trimb[4] vdd 0.165113f
C64 dacp_0/bootstrapped_sw_p_0/vbsl vinp 0.012179f
C65 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n3 0.336612f
C66 cal en 3.472141f
C67 sarlogic_0/net16 vdd 0.001182f
C68 sarlogic_0/trimb[1] sarlogic_0/trimb[4] 2.933839f
C69 cal vdd 3.379161f
C70 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/ndum 0.06073f
C71 vdd sarlogic_0/net14 0.005269f
C72 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n1 0.134826f
C73 dacp_0/sample valid 0.161748f
C74 dacn_0/ctl10 sarlogic_0/trim[3] 0.097876f
C75 comparator_0/ip comparator_0/trim_right_0/trim_switch_right_0/XM1_trim_right_0/D 1.60623f
C76 latch_0/R buffer_0/out 0.136735f
C77 sarlogic_0/net26 vdd 0.001136f
C78 dacp_0/out dacp_0/carray_p_0/n0 1.702719f
C79 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n3 25.8929f
C80 result[9] vdd 3.421719f
C81 comparator_0/trim_right_0/trim_switch_right_0/XM2_trim_right_0/D vdd 0.037004f
C82 m5_n124784_n195240# vdd 1.18282f
C83 dacp_0/ctl6 dacp_0/ctl5 3.114209f
C84 comparator_0/in vdd 0.39079f
C85 dacp_0/ctl1 vdd 0.85682f
C86 dacp_0/out dacp_0/carray_p_0/n1 3.365905f
C87 buffer_0/out vdd 0.039903f
C88 comparator_0/trim_left_0/trim_switch_left_0/n2 vdd 0.037004f
C89 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n5 5.60732f
C90 dacp_0/carray_p_0/n1 dacp_0/carray_p_0/ndum 8.161696f
C91 sarlogic_0/trimb[0] sarlogic_0/trimb[2] 3.097479f
C92 dacn_0/ctl10 vdd 0.357034f
C93 dacp_0/ctl6 vdd 0.474034f
C94 dacn_0/bootstrapped_sw_n_0/enb vdd 0.028031f
C95 vinn vdd 4.8626f
C96 dacp_0/ctl10 vdd 0.357034f
C97 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n2 0.996568f
C98 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n1 0.134562f
C99 sarlogic_0/trim[2] sarlogic_0/trim[3] 2.959509f
C100 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n4 0.614078f
C101 dacp_0/out dacp_0/carray_p_0/n3 13.201303f
C102 sarlogic_0/trim[3] vdd 0.565475f
C103 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/ndum 0.025424f
C104 buffer_0/buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vdd 0.011155f
C105 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n3 1.46111f
C106 latch_0/R vdd 0.172958f
C107 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n7 29.51607f
C108 dacn_0/ctl5 vdd 0.464997f
C109 comparator_0/in comparator_0/trim_left_0/trim_switch_left_0/n0 1.60623f
C110 result[5] vdd 3.379161f
C111 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n3 22.8406f
C112 dacp_0/ctl5 vdd 0.464997f
C113 comparator_0/ip comparator_0/trim_right_0/trim_switch_right_0/XM0_trim_right_0/D 1.60623f
C114 latch_0/Qn vdd 0.044756f
C115 en vdd 3.379161f
C116 dacn_0/ctl3 vdd 0.54157f
C117 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n0 0.097254f
C118 sarlogic_0/trim[2] vdd 0.142474f
C119 dacp_0/out dacp_0/carray_p_0/n6 0.105055p
C120 dacn_0/carray_n_0/n8 dacn_0/out 0.420152p
C121 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/ndum 0.025424f
C122 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n9 87.10265f
C123 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n0 0.099202f
C124 dacp_0/sample sarlogic_0/net27 0.004307f
C125 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n8 2.84323f
C126 sarlogic_0/trim[4] vdd 0.167468f
C127 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n0 0.025424f
C128 sarlogic_0/trimb[1] vdd 0.116601f
C129 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n5 5.60732f
C130 dacn_0/carray_n_0/n2 dacn_0/out 6.640605f
C131 dacp_0/ctl8 vdd 0.393337f
C132 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n9 0.996568f
C133 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n4 0.213096f
C134 comparator_0/trim_left_0/trim_switch_left_0/n1 comparator_0/in 1.60623f
C135 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n2 0.770114f
C136 dacp_0/sample cal 0.161292f
C137 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n5 0.207999f
C138 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n3 0.891504f
C139 buffer_0/buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# buffer_0/in 0.051091f
C140 comparator_0/in comparator_0/trim_left_0/trim_switch_left_0/n4 12.849839f
C141 dacp_0/bootstrapped_sw_p_0/enb vdd 0.028031f
C142 comparator_0/in comparator_0/trim_left_0/trim_switch_left_0/n3 6.42492f
C143 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n1 0.134705f
C144 comparator_0/trim_left_0/trim_switch_left_0/n2 comparator_0/trim_left_0/trim_switch_left_0/n4 0.128631f
C145 result[0] vdd 3.413481f
C146 dacp_0/out dacp_0/carray_p_0/n4 26.32268f
C147 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D comparator_0/trim_right_0/trim_switch_right_0/XM3_trim_right_0/D 0.241184f
C148 dacp_0/out vdd 1.294434f
C149 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n7 50.178104f
C150 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/ndum 0.025424f
C151 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n0 0.06073f
C152 dacp_0/ctl1 dacp_0/ctl2 4.157828f
C153 result[1] vdd 3.379161f
C154 dacp_0/sample result[9] 0.161326f
C155 dacn_0/carray_n_0/n7 dacn_0/out 0.210032p
C156 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n9 29.51607f
C157 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n7 1.70387f
C158 buffer_0/in vdd 0.334395f
C159 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n3 0.346757f
C160 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n5 3.36878f
C161 dacn_0/ctl1 vdd 0.862936f
C162 dacp_0/bootstrapped_sw_p_0/vbsh vdd 1.163764f
C163 result[2] vdd 3.379161f
C164 sarlogic_0/trimb[3] sarlogic_0/trimb[2] 2.951539f
C165 dacp_0/out dacp_0/carray_p_0/ndum 1.640173f
C166 result[1] result[0] 3.472163f
C167 latch_0/tutyuu1 vdd 0.004699f
C168 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/n2 0.099202f
C169 result[4] result[5] 3.472163f
C170 sarlogic_0/trim[2] sarlogic_0/trim[0] 3.097479f
C171 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n5 28.589401f
C172 comparator_0/trim_left_0/trim_switch_left_0/n4 vdd 0.063975f
C173 result[6] result[5] 3.472163f
C174 dacp_0/out dacp_0/bootstrapped_sw_p_0/vbsh -0.061493f
C175 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D comparator_0/ip 12.849839f
C176 sarlogic_0/trim[0] vdd 0.115811f
C177 comparator_0/trim_left_0/trim_switch_left_0/n3 vdd 0.248007f
C178 vdd result[3] 3.379161f
C179 dacp_0/sample result[5] 0.160929f
C180 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n0 0.06073f
C181 dacp_0/carray_p_0/n1 dacp_0/carray_p_0/n2 16.597801f
C182 result[4] vdd 3.379161f
C183 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n1 0.278221f
C184 result[2] result[1] 3.472163f
C185 dacp_0/ctl2 vdd 1.255808f
C186 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n6 11.2161f
C187 result[6] vdd 3.379161f
C188 dacp_0/sample en 0.18575f
C189 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n1 16.597801f
C190 result[7] vdd 3.379161f
C191 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n6 0.207877f
C192 comparator_0/trim_left_0/trim_switch_left_0/n1 comparator_0/trim_left_0/trim_switch_left_0/n0 0.032158f
C193 dacp_0/sample vdd 6.670178f
C194 vinn dacn_0/bootstrapped_sw_n_0/vbsl 0.01281f
C195 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n1 0.205173f
C196 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n2 22.8406f
C197 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n4 27.491999f
C198 dacp_0/sample dacn_0/carray_n_0/ndum 0.002948f
C199 sarlogic_0/net24 vdd 0.004775f
C200 comparator_0/trim_left_0/trim_switch_left_0/n4 comparator_0/trim_left_0/trim_switch_left_0/n0 0.032158f
C201 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n3 0.025424f
C202 dacp_0/ctl3 vdd 0.54157f
C203 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n8 87.10265f
C204 dacn_0/ctl5 dacn_0/ctl4 3.37511f
C205 en clk 3.472163f
C206 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n3 0.891504f
C207 dacn_0/ctl6 dacn_0/ctl7 2.853301f
C208 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n1 0.205173f
C209 clk vdd 3.37924f
C210 dacp_0/sample result[0] 0.161748f
C211 dacn_0/out vdd 1.294433f
C212 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n6 34.326103f
C213 dacn_0/carray_n_0/n9 vdd 0.037587f
C214 dacn_0/ctl3 dacn_0/ctl4 3.636021f
C215 result[2] result[3] 3.472163f
C216 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n2 0.207877f
C217 dacn_0/out dacn_0/carray_n_0/ndum 1.640173f
C218 dacp_0/out dacp_0/carray_p_0/n5 52.565495f
C219 vdd rstn 3.41356f
C220 dacp_0/sample dacp_0/carray_p_0/ndum 0.002948f
C221 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n9 0.127951f
C222 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/ndum 0.025424f
C223 dacn_0/ctl4 vdd 0.62371f
C224 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/ndum 0.025424f
C225 buffer_0/buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# buffer_0/middle 0.00331f
C226 dacp_0/sample result[1] 0.160984f
C227 comparator_0/trim_left_0/trim_switch_left_0/n1 comparator_0/trim_left_0/trim_switch_left_0/n4 0.032158f
C228 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/ndum 0.025424f
C229 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D comparator_0/trim_right_0/trim_switch_right_0/XM2_trim_right_0/D 0.128631f
C230 latch_0/R buffer_0/middle 0.009828f
C231 dacn_0/bootstrapped_sw_n_0/vbsl vdd 1.266964f
C232 result[2] dacp_0/sample 0.160984f
C233 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n6 34.326103f
C234 comparator_0/trim_left_0/trim_switch_left_0/n4 comparator_0/trim_left_0/trim_switch_left_0/n3 0.241184f
C235 dacp_0/sample sarlogic_0/net59 0.022016f
C236 sarlogic_0/net20 vdd 0.004671f
C237 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n2 0.213096f
C238 buffer_0/middle vdd 0.138765f
C239 dacn_0/ctl9 dacn_0/ctl8 2.33149f
C240 dacn_0/ctl2 dacn_0/ctl3 3.89692f
C241 result[4] result[3] 3.472163f
C242 comparator_0/trim_right_0/trim_switch_right_0/XM0_trim_right_0/D comparator_0/trim_right_0/trim_switch_right_0/XM1_trim_right_0/D 0.032158f
C243 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n0 0.184985f
C244 sarlogic_0/trimb[0] vdd 0.115811f
C245 dacn_0/ctl2 vdd 1.173819f
C246 comparator_0/trim_right_0/trim_switch_right_0/XM3_trim_right_0/D comparator_0/ip 6.42492f
C247 sarlogic_0/trimb[1] sarlogic_0/trimb[0] 2.995159f
C248 dacp_0/bootstrapped_sw_p_0/vbsl vdd 1.266964f
C249 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n4 1.70387f
C250 dacp_0/sample result[3] 0.160929f
C251 dacp_0/sample result[4] 0.160929f
C252 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n1 0.342393f
C253 result[6] result[7] 3.472163f
C254 sarlogic_0/output10/a_224_472# vdd 0.006335f
C255 result[9] result[8] 3.472163f
C256 dacp_0/out dacp_0/carray_p_0/n2 6.640605f
C257 dacp_0/sample result[6] 0.161003f
C258 vinp vdd 4.8626f
C259 dacp_0/sample result[7] 0.161003f
C260 dacp_0/carray_p_0/n2 dacp_0/carray_p_0/ndum 0.041162f
C261 dacn_0/bootstrapped_sw_n_0/vbsh vdd 1.163766f
C262 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D vdd 0.063975f
C263 dacp_0/ctl3 dacp_0/ctl2 3.896919f
C264 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n3 1.911225f
C265 buffer_0/in buffer_0/middle 0.005044f
C266 cal valid 3.472163f
C267 latch_0/R latch_0/S 0.235348f
C268 dacp_0/out dacp_0/bootstrapped_sw_p_0/vbsl -0.035593f
C269 dacp_0/out dacp_0/carray_p_0/n7 0.210032p
C270 latch_0/R latch_0/tutyuu2 0.004541f
C271 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/ndum 0.06073f
C272 dacn_0/ctl1 dacn_0/ctl2 4.157831f
C273 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n0 0.097254f
C274 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n1 8.161696f
C275 dacn_0/ctl6 dacn_0/ctl5 3.114201f
C276 latch_0/S latch_0/Qn 0.002019f
C277 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n8 0.770114f
C278 dacn_0/ctl7 dacn_0/ctl8 2.59239f
C279 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/ndum 0.025424f
C280 m5_121216_86040# vdd 1.18282f
C281 dacp_0/sample clk 0.171212f
C282 latch_0/S vdd 0.04502f
C283 dacn_0/carray_n_0/n0 dacn_0/carray_n_0/n3 0.051666f
C284 dacp_0/ctl5 dacp_0/ctl4 3.375109f
C285 dacn_0/out dacn_0/carray_n_0/n3 13.201303f
C286 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n6 14.716781f
C287 sarlogic_0/trimb[3] dacp_0/ctl10 0.087957f
C288 dacn_0/carray_n_0/n3 dacn_0/carray_n_0/n9 1.911225f
C289 dacp_0/sample rstn 0.161326f
C290 latch_0/tutyuu2 vdd 0.077568f
C291 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n3 25.8929f
C292 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n1 0.278221f
C293 dacn_0/ctl6 vdd 0.474034f
C294 dacp_0/ctl4 vdd 0.624893f
C295 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n3 0.346757f
C296 latch_0/R latch_0/Q 0.001863f
C297 dacn_0/ctl10 dacn_0/ctl9 2.076967f
C298 dacn_0/out dacn_0/carray_n_0/n0 1.702719f
C299 dacn_0/carray_n_0/n0 dacn_0/carray_n_0/n9 0.184985f
C300 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n8 50.178104f
C301 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n0 0.040502f
C302 sarlogic_0/trimb[2] vdd 0.139824f
C303 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D comparator_0/trim_right_0/trim_switch_right_0/XM1_trim_right_0/D 0.032158f
C304 result[8] vdd 3.530239f
C305 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n3 1.46111f
C306 dacn_0/out dacn_0/carray_n_0/n9 0.846152p
C307 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n0 0.025424f
C308 dacp_0/ctl7 dacp_0/ctl6 2.853299f
C309 dacn_0/carray_n_0/n4 dacn_0/out 26.32268f
C310 clk rstn 3.472163f
C311 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n7 0.485242f
C312 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n9 3.740571f
C313 latch_0/Q vdd 0.314864f
C314 dacn_0/carray_n_0/n5 dacn_0/out 52.565495f
C315 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n9 7.39935f
C316 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n4 3.740571f
C317 dacp_0/carray_p_0/n9 vdd 0.037587f
C318 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n5 27.491999f
C319 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n2 0.207999f
C320 dacn_0/out dacn_0/bootstrapped_sw_n_0/vbsl -0.035593f
C321 sarlogic_0/trimb[3] vdd 0.565475f
C322 m5_158680_n100000# vss 0.718816p $ **FLOATING
C323 m5_121216_n195240# vss 81.3617f $ **FLOATING
C324 m5_n124784_n195240# vss 81.3617f $ **FLOATING
C325 m5_121216_86040# vss 81.3617f $ **FLOATING
C326 m5_n124784_86040# vss 81.3617f $ **FLOATING
C327 m5_n161680_n100000# vss 0.718816p $ **FLOATING
C328 sarlogic_0/_034_ vss 0.304805f
C329 sarlogic_0/_160_ vss 1.542665f
C330 sarlogic_0/_166_ vss 0.299751f
C331 sarlogic_0/output41/a_224_472# vss 2.38465f
C332 sarlogic_0/net6 vss 1.112469f
C333 sarlogic_0/output6/a_224_472# vss 2.38465f
C334 sarlogic_0/FILLER_0_12_196/a_36_472# vss 0.417394f
C335 sarlogic_0/FILLER_0_12_196/a_124_375# vss 0.246306f
C336 result[3] vss 25.244722f
C337 sarlogic_0/net30 vss 1.81422f
C338 sarlogic_0/output30/a_224_472# vss 2.38465f
C339 sarlogic_0/_047_ vss 0.374694f
C340 sarlogic_0/_201_/a_67_603# vss 0.345683f
C341 sarlogic_0/_416_/a_2560_156# vss 0.016968f
C342 sarlogic_0/_416_/a_2665_112# vss 0.62251f
C343 sarlogic_0/_416_/a_2248_156# vss 0.371662f
C344 sarlogic_0/_416_/a_1204_472# vss 0.012971f
C345 sarlogic_0/_416_/a_1000_472# vss 0.291735f
C346 sarlogic_0/_416_/a_796_472# vss 0.023206f
C347 sarlogic_0/_416_/a_1308_423# vss 0.279043f
C348 sarlogic_0/_416_/a_448_472# vss 0.684413f
C349 sarlogic_0/_416_/a_36_151# vss 1.43589f
C350 sarlogic_0/FILLER_0_13_290/a_36_472# vss 0.417394f
C351 sarlogic_0/FILLER_0_13_290/a_124_375# vss 0.246306f
C352 sarlogic_0/_278_/a_36_160# vss 0.696445f
C353 sarlogic_0/_145_ vss 0.546455f
C354 sarlogic_0/FILLER_0_13_72/a_484_472# vss 0.345058f
C355 sarlogic_0/FILLER_0_13_72/a_36_472# vss 0.404746f
C356 sarlogic_0/FILLER_0_13_72/a_572_375# vss 0.232991f
C357 sarlogic_0/FILLER_0_13_72/a_124_375# vss 0.185089f
C358 sarlogic_0/FILLER_0_14_235/a_484_472# vss 0.345058f
C359 sarlogic_0/FILLER_0_14_235/a_36_472# vss 0.404746f
C360 sarlogic_0/FILLER_0_14_235/a_572_375# vss 0.232991f
C361 sarlogic_0/FILLER_0_14_235/a_124_375# vss 0.185089f
C362 sarlogic_0/_156_ vss 0.593796f
C363 sarlogic_0/_107_ vss 0.391583f
C364 sarlogic_0/_295_/a_36_472# vss 0.031137f
C365 sarlogic_0/_022_ vss 0.387773f
C366 sarlogic_0/_433_/a_2560_156# vss 0.016968f
C367 sarlogic_0/_433_/a_2665_112# vss 0.62251f
C368 sarlogic_0/_433_/a_2248_156# vss 0.371662f
C369 sarlogic_0/_433_/a_1204_472# vss 0.012971f
C370 sarlogic_0/_433_/a_1000_472# vss 0.291735f
C371 sarlogic_0/_433_/a_796_472# vss 0.023206f
C372 sarlogic_0/_433_/a_1308_423# vss 0.279043f
C373 sarlogic_0/_433_/a_448_472# vss 0.684413f
C374 sarlogic_0/_433_/a_36_151# vss 1.43589f
C375 sarlogic_0/FILLER_0_5_148/a_484_472# vss 0.345058f
C376 sarlogic_0/FILLER_0_5_148/a_36_472# vss 0.404746f
C377 sarlogic_0/FILLER_0_5_148/a_572_375# vss 0.232991f
C378 sarlogic_0/FILLER_0_5_148/a_124_375# vss 0.185089f
C379 sarlogic_0/_167_ vss 0.285904f
C380 sarlogic_0/_381_/a_36_472# vss 0.031137f
C381 sarlogic_0/net40 vss 1.845219f
C382 sarlogic_0/output40/a_224_472# vss 2.38465f
C383 sarlogic_0/cal_count\[0\] vss 0.893784f
C384 sarlogic_0/_039_ vss 0.412301f
C385 sarlogic_0/_450_/a_2449_156# vss 0.049992f
C386 sarlogic_0/_450_/a_2225_156# vss 0.434082f
C387 sarlogic_0/_450_/a_3129_107# vss 0.58406f
C388 sarlogic_0/_450_/a_836_156# vss 0.019766f
C389 sarlogic_0/_450_/a_1040_527# vss 0.302082f
C390 sarlogic_0/_450_/a_1353_112# vss 0.286513f
C391 sarlogic_0/_450_/a_448_472# vss 1.21246f
C392 sarlogic_0/_450_/a_36_151# vss 1.31409f
C393 rstn vss 31.165571f
C394 sarlogic_0/FILLER_0_8_156/a_484_472# vss 0.345058f
C395 sarlogic_0/FILLER_0_8_156/a_36_472# vss 0.404746f
C396 sarlogic_0/FILLER_0_8_156/a_572_375# vss 0.232991f
C397 sarlogic_0/FILLER_0_8_156/a_124_375# vss 0.185089f
C398 sarlogic_0/FILLER_0_6_37/a_36_472# vss 0.417394f
C399 sarlogic_0/FILLER_0_6_37/a_124_375# vss 0.246306f
C400 sarlogic_0/FILLER_0_21_60/a_484_472# vss 0.345058f
C401 sarlogic_0/FILLER_0_21_60/a_36_472# vss 0.404746f
C402 sarlogic_0/FILLER_0_21_60/a_572_375# vss 0.232991f
C403 sarlogic_0/FILLER_0_21_60/a_124_375# vss 0.185089f
C404 sarlogic_0/FILLER_0_22_107/a_484_472# vss 0.345058f
C405 sarlogic_0/FILLER_0_22_107/a_36_472# vss 0.404746f
C406 sarlogic_0/FILLER_0_22_107/a_572_375# vss 0.232991f
C407 sarlogic_0/FILLER_0_22_107/a_124_375# vss 0.185089f
C408 sarlogic_0/FILLER_0_16_115/a_36_472# vss 0.417394f
C409 sarlogic_0/FILLER_0_16_115/a_124_375# vss 0.246306f
C410 sarlogic_0/FILLER_0_19_134/a_36_472# vss 0.417394f
C411 sarlogic_0/FILLER_0_19_134/a_124_375# vss 0.246306f
C412 sarlogic_0/FILLER_0_3_212/a_36_472# vss 0.417394f
C413 sarlogic_0/FILLER_0_3_212/a_124_375# vss 0.246306f
C414 sarlogic_0/FILLER_0_10_94/a_484_472# vss 0.345058f
C415 sarlogic_0/FILLER_0_10_94/a_36_472# vss 0.404746f
C416 sarlogic_0/FILLER_0_10_94/a_572_375# vss 0.232991f
C417 sarlogic_0/FILLER_0_10_94/a_124_375# vss 0.185089f
C418 sarlogic_0/FILLER_0_4_91/a_484_472# vss 0.345058f
C419 sarlogic_0/FILLER_0_4_91/a_36_472# vss 0.404746f
C420 sarlogic_0/FILLER_0_4_91/a_572_375# vss 0.232991f
C421 sarlogic_0/FILLER_0_4_91/a_124_375# vss 0.185089f
C422 sarlogic_0/net14 vss 1.508711f
C423 sarlogic_0/_202_/a_36_160# vss 0.696445f
C424 sarlogic_0/FILLER_0_6_231/a_484_472# vss 0.345058f
C425 sarlogic_0/FILLER_0_6_231/a_36_472# vss 0.404746f
C426 sarlogic_0/FILLER_0_6_231/a_572_375# vss 0.232991f
C427 sarlogic_0/FILLER_0_6_231/a_124_375# vss 0.185089f
C428 vdd vss 16.715534p
C429 sarlogic_0/_006_ vss 0.41456f
C430 sarlogic_0/_417_/a_2560_156# vss 0.016968f
C431 sarlogic_0/_417_/a_2665_112# vss 0.62251f
C432 sarlogic_0/_417_/a_2248_156# vss 0.371662f
C433 sarlogic_0/_417_/a_1204_472# vss 0.012971f
C434 sarlogic_0/_417_/a_1000_472# vss 0.291735f
C435 sarlogic_0/_417_/a_796_472# vss 0.023206f
C436 sarlogic_0/_417_/a_1308_423# vss 0.279043f
C437 sarlogic_0/_417_/a_448_472# vss 0.684413f
C438 sarlogic_0/_417_/a_36_151# vss 1.43589f
C439 sarlogic_0/_146_ vss 0.35443f
C440 sarlogic_0/mask\[6\] vss 1.246962f
C441 sarlogic_0/_348_/a_49_472# vss 0.054843f
C442 sarlogic_0/_365_/a_36_68# vss 0.150048f
C443 sarlogic_0/_023_ vss 0.345812f
C444 sarlogic_0/_434_/a_2560_156# vss 0.016968f
C445 sarlogic_0/_434_/a_2665_112# vss 0.62251f
C446 sarlogic_0/_434_/a_2248_156# vss 0.371662f
C447 sarlogic_0/_434_/a_1204_472# vss 0.012971f
C448 sarlogic_0/_434_/a_1000_472# vss 0.291735f
C449 sarlogic_0/_434_/a_796_472# vss 0.023206f
C450 sarlogic_0/_434_/a_1308_423# vss 0.279043f
C451 sarlogic_0/_434_/a_448_472# vss 0.684413f
C452 sarlogic_0/_434_/a_36_151# vss 1.43589f
C453 sarlogic_0/FILLER_0_5_136/a_36_472# vss 0.417394f
C454 sarlogic_0/FILLER_0_5_136/a_124_375# vss 0.246306f
C455 sarlogic_0/FILLER_0_18_209/a_484_472# vss 0.345058f
C456 sarlogic_0/FILLER_0_18_209/a_36_472# vss 0.404746f
C457 sarlogic_0/FILLER_0_18_209/a_572_375# vss 0.232991f
C458 sarlogic_0/FILLER_0_18_209/a_124_375# vss 0.185089f
C459 sarlogic_0/FILLER_0_12_28/a_36_472# vss 0.417394f
C460 sarlogic_0/FILLER_0_12_28/a_124_375# vss 0.246306f
C461 sarlogic_0/_040_ vss 0.355703f
C462 sarlogic_0/_451_/a_2449_156# vss 0.049992f
C463 sarlogic_0/_451_/a_2225_156# vss 0.434082f
C464 sarlogic_0/_451_/a_3129_107# vss 0.58406f
C465 sarlogic_0/_451_/a_836_156# vss 0.019766f
C466 sarlogic_0/_451_/a_1040_527# vss 0.302082f
C467 sarlogic_0/_451_/a_1353_112# vss 0.286513f
C468 sarlogic_0/_451_/a_448_472# vss 1.21246f
C469 sarlogic_0/_451_/a_36_151# vss 1.31409f
C470 sarlogic_0/FILLER_0_6_47/a_3172_472# vss 0.345058f
C471 sarlogic_0/FILLER_0_6_47/a_2724_472# vss 0.33241f
C472 sarlogic_0/FILLER_0_6_47/a_2276_472# vss 0.33241f
C473 sarlogic_0/FILLER_0_6_47/a_1828_472# vss 0.33241f
C474 sarlogic_0/FILLER_0_6_47/a_1380_472# vss 0.33241f
C475 sarlogic_0/FILLER_0_6_47/a_932_472# vss 0.33241f
C476 sarlogic_0/FILLER_0_6_47/a_484_472# vss 0.33241f
C477 sarlogic_0/FILLER_0_6_47/a_36_472# vss 0.404746f
C478 sarlogic_0/FILLER_0_6_47/a_3260_375# vss 0.233093f
C479 sarlogic_0/FILLER_0_6_47/a_2812_375# vss 0.17167f
C480 sarlogic_0/FILLER_0_6_47/a_2364_375# vss 0.17167f
C481 sarlogic_0/FILLER_0_6_47/a_1916_375# vss 0.17167f
C482 sarlogic_0/FILLER_0_6_47/a_1468_375# vss 0.17167f
C483 sarlogic_0/FILLER_0_6_47/a_1020_375# vss 0.17167f
C484 sarlogic_0/FILLER_0_6_47/a_572_375# vss 0.17167f
C485 sarlogic_0/FILLER_0_6_47/a_124_375# vss 0.185915f
C486 sarlogic_0/FILLER_0_21_150/a_36_472# vss 0.417394f
C487 sarlogic_0/FILLER_0_21_150/a_124_375# vss 0.246306f
C488 sarlogic_0/FILLER_0_15_180/a_484_472# vss 0.345058f
C489 sarlogic_0/FILLER_0_15_180/a_36_472# vss 0.404746f
C490 sarlogic_0/FILLER_0_15_180/a_572_375# vss 0.232991f
C491 sarlogic_0/FILLER_0_15_180/a_124_375# vss 0.185089f
C492 sarlogic_0/FILLER_0_22_128/a_3172_472# vss 0.345058f
C493 sarlogic_0/FILLER_0_22_128/a_2724_472# vss 0.33241f
C494 sarlogic_0/FILLER_0_22_128/a_2276_472# vss 0.33241f
C495 sarlogic_0/FILLER_0_22_128/a_1828_472# vss 0.33241f
C496 sarlogic_0/FILLER_0_22_128/a_1380_472# vss 0.33241f
C497 sarlogic_0/FILLER_0_22_128/a_932_472# vss 0.33241f
C498 sarlogic_0/FILLER_0_22_128/a_484_472# vss 0.33241f
C499 sarlogic_0/FILLER_0_22_128/a_36_472# vss 0.404746f
C500 sarlogic_0/FILLER_0_22_128/a_3260_375# vss 0.233093f
C501 sarlogic_0/FILLER_0_22_128/a_2812_375# vss 0.17167f
C502 sarlogic_0/FILLER_0_22_128/a_2364_375# vss 0.17167f
C503 sarlogic_0/FILLER_0_22_128/a_1916_375# vss 0.17167f
C504 sarlogic_0/FILLER_0_22_128/a_1468_375# vss 0.17167f
C505 sarlogic_0/FILLER_0_22_128/a_1020_375# vss 0.17167f
C506 sarlogic_0/FILLER_0_22_128/a_572_375# vss 0.17167f
C507 sarlogic_0/FILLER_0_22_128/a_124_375# vss 0.185915f
C508 sarlogic_0/FILLER_0_19_111/a_484_472# vss 0.345058f
C509 sarlogic_0/FILLER_0_19_111/a_36_472# vss 0.404746f
C510 sarlogic_0/FILLER_0_19_111/a_572_375# vss 0.232991f
C511 sarlogic_0/FILLER_0_19_111/a_124_375# vss 0.185089f
C512 sarlogic_0/FILLER_0_19_155/a_484_472# vss 0.345058f
C513 sarlogic_0/FILLER_0_19_155/a_36_472# vss 0.404746f
C514 sarlogic_0/FILLER_0_19_155/a_572_375# vss 0.232991f
C515 sarlogic_0/FILLER_0_19_155/a_124_375# vss 0.185089f
C516 sarlogic_0/net11 vss 1.328455f
C517 sarlogic_0/net21 vss 1.922829f
C518 sarlogic_0/_007_ vss 0.309495f
C519 sarlogic_0/net77 vss 1.39077f
C520 sarlogic_0/_418_/a_2560_156# vss 0.016968f
C521 sarlogic_0/_418_/a_2665_112# vss 0.62251f
C522 sarlogic_0/_418_/a_2248_156# vss 0.371662f
C523 sarlogic_0/_418_/a_1204_472# vss 0.012971f
C524 sarlogic_0/_418_/a_1000_472# vss 0.291735f
C525 sarlogic_0/_418_/a_796_472# vss 0.023206f
C526 sarlogic_0/_418_/a_1308_423# vss 0.279043f
C527 sarlogic_0/_418_/a_448_472# vss 0.684413f
C528 sarlogic_0/_418_/a_36_151# vss 1.43589f
C529 sarlogic_0/_220_/a_67_603# vss 0.345683f
C530 sarlogic_0/FILLER_0_9_282/a_484_472# vss 0.345058f
C531 sarlogic_0/FILLER_0_9_282/a_36_472# vss 0.404746f
C532 sarlogic_0/FILLER_0_9_282/a_572_375# vss 0.232991f
C533 sarlogic_0/FILLER_0_9_282/a_124_375# vss 0.185089f
C534 sarlogic_0/FILLER_0_18_37/a_1380_472# vss 0.345058f
C535 sarlogic_0/FILLER_0_18_37/a_932_472# vss 0.33241f
C536 sarlogic_0/FILLER_0_18_37/a_484_472# vss 0.33241f
C537 sarlogic_0/FILLER_0_18_37/a_36_472# vss 0.404746f
C538 sarlogic_0/FILLER_0_18_37/a_1468_375# vss 0.233029f
C539 sarlogic_0/FILLER_0_18_37/a_1020_375# vss 0.171606f
C540 sarlogic_0/FILLER_0_18_37/a_572_375# vss 0.171606f
C541 sarlogic_0/FILLER_0_18_37/a_124_375# vss 0.185399f
C542 sarlogic_0/FILLER_0_2_127/a_36_472# vss 0.417394f
C543 sarlogic_0/FILLER_0_2_127/a_124_375# vss 0.246306f
C544 sarlogic_0/_157_ vss 0.531763f
C545 sarlogic_0/_435_/a_2560_156# vss 0.016968f
C546 sarlogic_0/_435_/a_2665_112# vss 0.62251f
C547 sarlogic_0/_435_/a_2248_156# vss 0.371662f
C548 sarlogic_0/_435_/a_1204_472# vss 0.012971f
C549 sarlogic_0/_435_/a_1000_472# vss 0.291735f
C550 sarlogic_0/_435_/a_796_472# vss 0.023206f
C551 sarlogic_0/_435_/a_1308_423# vss 0.279043f
C552 sarlogic_0/_435_/a_448_472# vss 0.684413f
C553 sarlogic_0/_435_/a_36_151# vss 1.43589f
C554 sarlogic_0/_108_ vss 0.411979f
C555 sarlogic_0/_297_/a_36_472# vss 0.031137f
C556 sarlogic_0/trim_mask\[3\] vss 1.081535f
C557 sarlogic_0/_164_ vss 1.3268f
C558 sarlogic_0/_383_/a_36_472# vss 0.031137f
C559 sarlogic_0/_041_ vss 0.299289f
C560 sarlogic_0/_452_/a_2449_156# vss 0.049992f
C561 sarlogic_0/_452_/a_2225_156# vss 0.434082f
C562 sarlogic_0/_452_/a_3129_107# vss 0.58406f
C563 sarlogic_0/_452_/a_836_156# vss 0.019766f
C564 sarlogic_0/_452_/a_1040_527# vss 0.302082f
C565 sarlogic_0/_452_/a_1353_112# vss 0.286513f
C566 sarlogic_0/_452_/a_448_472# vss 1.21246f
C567 sarlogic_0/_452_/a_36_151# vss 1.31409f
C568 sarlogic_0/FILLER_0_6_79/a_36_472# vss 0.417394f
C569 sarlogic_0/FILLER_0_6_79/a_124_375# vss 0.246306f
C570 sarlogic_0/net59 vss 5.044369f
C571 sarlogic_0/FILLER_0_15_59/a_484_472# vss 0.345058f
C572 sarlogic_0/FILLER_0_15_59/a_36_472# vss 0.404746f
C573 sarlogic_0/FILLER_0_15_59/a_572_375# vss 0.232991f
C574 sarlogic_0/FILLER_0_15_59/a_124_375# vss 0.185089f
C575 sarlogic_0/FILLER_0_3_221/a_1380_472# vss 0.345058f
C576 sarlogic_0/FILLER_0_3_221/a_932_472# vss 0.33241f
C577 sarlogic_0/FILLER_0_3_221/a_484_472# vss 0.33241f
C578 sarlogic_0/FILLER_0_3_221/a_36_472# vss 0.404746f
C579 sarlogic_0/FILLER_0_3_221/a_1468_375# vss 0.233029f
C580 sarlogic_0/FILLER_0_3_221/a_1020_375# vss 0.171606f
C581 sarlogic_0/FILLER_0_3_221/a_572_375# vss 0.171606f
C582 sarlogic_0/FILLER_0_3_221/a_124_375# vss 0.185399f
C583 sarlogic_0/FILLER_0_19_187/a_484_472# vss 0.345058f
C584 sarlogic_0/FILLER_0_19_187/a_36_472# vss 0.404746f
C585 sarlogic_0/FILLER_0_19_187/a_572_375# vss 0.232991f
C586 sarlogic_0/FILLER_0_19_187/a_124_375# vss 0.185089f
C587 sarlogic_0/FILLER_0_20_15/a_1380_472# vss 0.345058f
C588 sarlogic_0/FILLER_0_20_15/a_932_472# vss 0.33241f
C589 sarlogic_0/FILLER_0_20_15/a_484_472# vss 0.33241f
C590 sarlogic_0/FILLER_0_20_15/a_36_472# vss 0.404746f
C591 sarlogic_0/FILLER_0_20_15/a_1468_375# vss 0.233029f
C592 sarlogic_0/FILLER_0_20_15/a_1020_375# vss 0.171606f
C593 sarlogic_0/FILLER_0_20_15/a_572_375# vss 0.171606f
C594 sarlogic_0/FILLER_0_20_15/a_124_375# vss 0.185399f
C595 sarlogic_0/_204_/a_67_603# vss 0.345683f
C596 sarlogic_0/_419_/a_2560_156# vss 0.016968f
C597 sarlogic_0/_419_/a_2665_112# vss 0.62251f
C598 sarlogic_0/_419_/a_2248_156# vss 0.371662f
C599 sarlogic_0/_419_/a_1204_472# vss 0.012971f
C600 sarlogic_0/_419_/a_1000_472# vss 0.291735f
C601 sarlogic_0/_419_/a_796_472# vss 0.023206f
C602 sarlogic_0/_419_/a_1308_423# vss 0.279043f
C603 sarlogic_0/_419_/a_448_472# vss 0.684413f
C604 sarlogic_0/_419_/a_36_151# vss 1.43589f
C605 sarlogic_0/_054_ vss 0.522819f
C606 sarlogic_0/_221_/a_36_160# vss 0.386641f
C607 sarlogic_0/FILLER_0_9_270/a_484_472# vss 0.345058f
C608 sarlogic_0/FILLER_0_9_270/a_36_472# vss 0.404746f
C609 sarlogic_0/FILLER_0_9_270/a_572_375# vss 0.232991f
C610 sarlogic_0/FILLER_0_9_270/a_124_375# vss 0.185089f
C611 sarlogic_0/FILLER_0_1_192/a_36_472# vss 0.417394f
C612 sarlogic_0/FILLER_0_1_192/a_124_375# vss 0.246306f
C613 sarlogic_0/FILLER_0_13_80/a_36_472# vss 0.417394f
C614 sarlogic_0/FILLER_0_13_80/a_124_375# vss 0.246306f
C615 sarlogic_0/_153_ vss 1.165862f
C616 sarlogic_0/_154_ vss 1.167112f
C617 sarlogic_0/_367_/a_36_68# vss 0.150048f
C618 sarlogic_0/_436_/a_2560_156# vss 0.016968f
C619 sarlogic_0/_436_/a_2665_112# vss 0.62251f
C620 sarlogic_0/_436_/a_2248_156# vss 0.371662f
C621 sarlogic_0/_436_/a_1204_472# vss 0.012971f
C622 sarlogic_0/_436_/a_1000_472# vss 0.291735f
C623 sarlogic_0/_436_/a_796_472# vss 0.023206f
C624 sarlogic_0/_436_/a_1308_423# vss 0.279043f
C625 sarlogic_0/_436_/a_448_472# vss 0.684413f
C626 sarlogic_0/_436_/a_36_151# vss 1.43589f
C627 sarlogic_0/FILLER_0_10_107/a_484_472# vss 0.345058f
C628 sarlogic_0/FILLER_0_10_107/a_36_472# vss 0.404746f
C629 sarlogic_0/FILLER_0_10_107/a_572_375# vss 0.232991f
C630 sarlogic_0/FILLER_0_10_107/a_124_375# vss 0.185089f
C631 sarlogic_0/_168_ vss 0.336537f
C632 sarlogic_0/net51 vss 2.105066f
C633 sarlogic_0/_042_ vss 0.323587f
C634 sarlogic_0/_453_/a_2560_156# vss 0.016968f
C635 sarlogic_0/_453_/a_2665_112# vss 0.62251f
C636 sarlogic_0/_453_/a_2248_156# vss 0.371662f
C637 sarlogic_0/_453_/a_1204_472# vss 0.012971f
C638 sarlogic_0/_453_/a_1000_472# vss 0.291735f
C639 sarlogic_0/_453_/a_796_472# vss 0.023206f
C640 sarlogic_0/_453_/a_1308_423# vss 0.279043f
C641 sarlogic_0/_453_/a_448_472# vss 0.684413f
C642 sarlogic_0/_453_/a_36_151# vss 1.43589f
C643 sarlogic_0/FILLER_0_19_142/a_36_472# vss 0.417394f
C644 sarlogic_0/FILLER_0_19_142/a_124_375# vss 0.246306f
C645 sarlogic_0/_048_ vss 0.358805f
C646 sarlogic_0/_205_/a_36_160# vss 0.696445f
C647 sarlogic_0/net43 vss 1.236377f
C648 sarlogic_0/FILLER_0_3_78/a_484_472# vss 0.345058f
C649 sarlogic_0/FILLER_0_3_78/a_36_472# vss 0.404746f
C650 sarlogic_0/FILLER_0_3_78/a_572_375# vss 0.232991f
C651 sarlogic_0/FILLER_0_3_78/a_124_375# vss 0.185089f
C652 sarlogic_0/_437_/a_2560_156# vss 0.016968f
C653 sarlogic_0/_437_/a_2665_112# vss 0.62251f
C654 sarlogic_0/_437_/a_2248_156# vss 0.371662f
C655 sarlogic_0/_437_/a_1204_472# vss 0.012971f
C656 sarlogic_0/_437_/a_1000_472# vss 0.291735f
C657 sarlogic_0/_437_/a_796_472# vss 0.023206f
C658 sarlogic_0/_437_/a_1308_423# vss 0.279043f
C659 sarlogic_0/_437_/a_448_472# vss 0.684413f
C660 sarlogic_0/_437_/a_36_151# vss 1.43589f
C661 sarlogic_0/_109_ vss 0.319326f
C662 sarlogic_0/_299_/a_36_472# vss 0.031137f
C663 sarlogic_0/net37 vss 1.529713f
C664 sarlogic_0/_385_/a_36_68# vss 0.112263f
C665 sarlogic_0/FILLER_0_0_266/a_36_472# vss 0.417394f
C666 sarlogic_0/FILLER_0_0_266/a_124_375# vss 0.246306f
C667 sarlogic_0/net12 vss 1.263595f
C668 sarlogic_0/net22 vss 2.108509f
C669 sarlogic_0/FILLER_0_9_290/a_36_472# vss 0.417394f
C670 sarlogic_0/FILLER_0_9_290/a_124_375# vss 0.246306f
C671 sarlogic_0/_223_/a_36_160# vss 0.696445f
C672 sarlogic_0/FILLER_0_14_263/a_36_472# vss 0.417394f
C673 sarlogic_0/FILLER_0_14_263/a_124_375# vss 0.246306f
C674 sarlogic_0/_158_ vss 0.309522f
C675 sarlogic_0/_369_/a_36_68# vss 0.150048f
C676 sarlogic_0/net71 vss 1.420869f
C677 sarlogic_0/_438_/a_2560_156# vss 0.016968f
C678 sarlogic_0/_438_/a_2665_112# vss 0.62251f
C679 sarlogic_0/_438_/a_2248_156# vss 0.371662f
C680 sarlogic_0/_438_/a_1204_472# vss 0.012971f
C681 sarlogic_0/_438_/a_1000_472# vss 0.291735f
C682 sarlogic_0/_438_/a_796_472# vss 0.023206f
C683 sarlogic_0/_438_/a_1308_423# vss 0.279043f
C684 sarlogic_0/_438_/a_448_472# vss 0.684413f
C685 sarlogic_0/_438_/a_36_151# vss 1.43589f
C686 sarlogic_0/FILLER_0_23_274/a_36_472# vss 0.417394f
C687 sarlogic_0/FILLER_0_23_274/a_124_375# vss 0.246306f
C688 sarlogic_0/FILLER_0_17_282/a_36_472# vss 0.417394f
C689 sarlogic_0/FILLER_0_17_282/a_124_375# vss 0.246306f
C690 sarlogic_0/FILLER_0_5_198/a_484_472# vss 0.345058f
C691 sarlogic_0/FILLER_0_5_198/a_36_472# vss 0.404746f
C692 sarlogic_0/FILLER_0_5_198/a_572_375# vss 0.232991f
C693 sarlogic_0/FILLER_0_5_198/a_124_375# vss 0.185089f
C694 sarlogic_0/_163_ vss 1.03762f
C695 sarlogic_0/_169_ vss 0.245383f
C696 sarlogic_0/_386_/a_848_380# vss 0.40208f
C697 sarlogic_0/_386_/a_124_24# vss 0.591898f
C698 sarlogic_0/FILLER_0_20_2/a_484_472# vss 0.345058f
C699 sarlogic_0/FILLER_0_20_2/a_36_472# vss 0.404746f
C700 sarlogic_0/FILLER_0_20_2/a_572_375# vss 0.232991f
C701 sarlogic_0/FILLER_0_20_2/a_124_375# vss 0.185089f
C702 sarlogic_0/FILLER_0_16_154/a_1380_472# vss 0.345058f
C703 sarlogic_0/FILLER_0_16_154/a_932_472# vss 0.33241f
C704 sarlogic_0/FILLER_0_16_154/a_484_472# vss 0.33241f
C705 sarlogic_0/FILLER_0_16_154/a_36_472# vss 0.404746f
C706 sarlogic_0/FILLER_0_16_154/a_1468_375# vss 0.233029f
C707 sarlogic_0/FILLER_0_16_154/a_1020_375# vss 0.171606f
C708 sarlogic_0/FILLER_0_16_154/a_572_375# vss 0.171606f
C709 sarlogic_0/FILLER_0_16_154/a_124_375# vss 0.185399f
C710 sarlogic_0/FILLER_0_0_232/a_36_472# vss 0.417394f
C711 sarlogic_0/FILLER_0_0_232/a_124_375# vss 0.246306f
C712 sarlogic_0/FILLER_0_19_195/a_36_472# vss 0.417394f
C713 sarlogic_0/FILLER_0_19_195/a_124_375# vss 0.246306f
C714 sarlogic_0/_049_ vss 0.329957f
C715 sarlogic_0/net33 vss 1.934915f
C716 sarlogic_0/_207_/a_67_603# vss 0.345683f
C717 sarlogic_0/FILLER_0_3_54/a_36_472# vss 0.417394f
C718 sarlogic_0/FILLER_0_3_54/a_124_375# vss 0.246306f
C719 sarlogic_0/FILLER_0_2_101/a_36_472# vss 0.417394f
C720 sarlogic_0/FILLER_0_2_101/a_124_375# vss 0.246306f
C721 sarlogic_0/trim_mask\[0\] vss 0.605753f
C722 sarlogic_0/_439_/a_2560_156# vss 0.016968f
C723 sarlogic_0/_439_/a_2665_112# vss 0.62251f
C724 sarlogic_0/_439_/a_2248_156# vss 0.371662f
C725 sarlogic_0/_439_/a_1204_472# vss 0.012971f
C726 sarlogic_0/_439_/a_1000_472# vss 0.291735f
C727 sarlogic_0/_439_/a_796_472# vss 0.023206f
C728 sarlogic_0/_439_/a_1308_423# vss 0.279043f
C729 sarlogic_0/_439_/a_448_472# vss 0.684413f
C730 sarlogic_0/_439_/a_36_151# vss 1.43589f
C731 sarlogic_0/_066_ vss 0.333041f
C732 sarlogic_0/FILLER_0_23_44/a_1380_472# vss 0.345058f
C733 sarlogic_0/FILLER_0_23_44/a_932_472# vss 0.33241f
C734 sarlogic_0/FILLER_0_23_44/a_484_472# vss 0.33241f
C735 sarlogic_0/FILLER_0_23_44/a_36_472# vss 0.404746f
C736 sarlogic_0/FILLER_0_23_44/a_1468_375# vss 0.233029f
C737 sarlogic_0/FILLER_0_23_44/a_1020_375# vss 0.171606f
C738 sarlogic_0/FILLER_0_23_44/a_572_375# vss 0.171606f
C739 sarlogic_0/FILLER_0_23_44/a_124_375# vss 0.185399f
C740 sarlogic_0/FILLER_0_23_88/a_36_472# vss 0.417394f
C741 sarlogic_0/FILLER_0_23_88/a_124_375# vss 0.246306f
C742 sarlogic_0/FILLER_0_5_164/a_484_472# vss 0.345058f
C743 sarlogic_0/FILLER_0_5_164/a_36_472# vss 0.404746f
C744 sarlogic_0/FILLER_0_5_164/a_572_375# vss 0.232991f
C745 sarlogic_0/FILLER_0_5_164/a_124_375# vss 0.185089f
C746 sarlogic_0/_060_ vss 2.485177f
C747 sarlogic_0/_113_ vss 2.833205f
C748 sarlogic_0/_090_ vss 2.629271f
C749 sarlogic_0/_310_/a_49_472# vss 0.098072f
C750 sarlogic_0/_037_ vss 0.467089f
C751 sarlogic_0/_170_ vss 0.413995f
C752 sarlogic_0/_387_/a_36_113# vss 0.418095f
C753 sarlogic_0/_208_/a_36_160# vss 0.696445f
C754 sarlogic_0/FILLER_0_18_76/a_484_472# vss 0.345058f
C755 sarlogic_0/FILLER_0_18_76/a_36_472# vss 0.404746f
C756 sarlogic_0/FILLER_0_18_76/a_572_375# vss 0.232991f
C757 sarlogic_0/FILLER_0_18_76/a_124_375# vss 0.185089f
C758 sarlogic_0/_225_/a_36_160# vss 0.386641f
C759 sarlogic_0/FILLER_0_2_177/a_484_472# vss 0.345058f
C760 sarlogic_0/FILLER_0_2_177/a_36_472# vss 0.404746f
C761 sarlogic_0/FILLER_0_2_177/a_572_375# vss 0.232991f
C762 sarlogic_0/FILLER_0_2_177/a_124_375# vss 0.185089f
C763 sarlogic_0/FILLER_0_2_111/a_1380_472# vss 0.345058f
C764 sarlogic_0/FILLER_0_2_111/a_932_472# vss 0.33241f
C765 sarlogic_0/FILLER_0_2_111/a_484_472# vss 0.33241f
C766 sarlogic_0/FILLER_0_2_111/a_36_472# vss 0.404746f
C767 sarlogic_0/FILLER_0_2_111/a_1468_375# vss 0.233029f
C768 sarlogic_0/FILLER_0_2_111/a_1020_375# vss 0.171606f
C769 sarlogic_0/FILLER_0_2_111/a_572_375# vss 0.171606f
C770 sarlogic_0/FILLER_0_2_111/a_124_375# vss 0.185399f
C771 sarlogic_0/FILLER_0_15_228/a_36_472# vss 0.417394f
C772 sarlogic_0/FILLER_0_15_228/a_124_375# vss 0.246306f
C773 sarlogic_0/net47 vss 2.314376f
C774 sarlogic_0/_242_/a_36_160# vss 0.696445f
C775 sarlogic_0/_117_ vss 1.266251f
C776 sarlogic_0/_311_/a_66_473# vss 0.11665f
C777 sarlogic_0/_043_ vss 0.487279f
C778 sarlogic_0/_190_/a_36_160# vss 0.696445f
C779 sarlogic_0/FILLER_0_9_105/a_484_472# vss 0.345058f
C780 sarlogic_0/FILLER_0_9_105/a_36_472# vss 0.404746f
C781 sarlogic_0/FILLER_0_9_105/a_572_375# vss 0.232991f
C782 sarlogic_0/FILLER_0_9_105/a_124_375# vss 0.185089f
C783 sarlogic_0/FILLER_0_13_100/a_36_472# vss 0.417394f
C784 sarlogic_0/FILLER_0_13_100/a_124_375# vss 0.246306f
C785 sarlogic_0/FILLER_0_22_177/a_1380_472# vss 0.345058f
C786 sarlogic_0/FILLER_0_22_177/a_932_472# vss 0.33241f
C787 sarlogic_0/FILLER_0_22_177/a_484_472# vss 0.33241f
C788 sarlogic_0/FILLER_0_22_177/a_36_472# vss 0.404746f
C789 sarlogic_0/FILLER_0_22_177/a_1468_375# vss 0.233029f
C790 sarlogic_0/FILLER_0_22_177/a_1020_375# vss 0.171606f
C791 sarlogic_0/FILLER_0_22_177/a_572_375# vss 0.171606f
C792 sarlogic_0/FILLER_0_22_177/a_124_375# vss 0.185399f
C793 sarlogic_0/FILLER_0_15_2/a_484_472# vss 0.345058f
C794 sarlogic_0/FILLER_0_15_2/a_36_472# vss 0.404746f
C795 sarlogic_0/FILLER_0_15_2/a_572_375# vss 0.232991f
C796 sarlogic_0/FILLER_0_15_2/a_124_375# vss 0.185089f
C797 sarlogic_0/FILLER_0_15_10/a_36_472# vss 0.417394f
C798 sarlogic_0/FILLER_0_15_10/a_124_375# vss 0.246306f
C799 sarlogic_0/FILLER_0_19_171/a_1380_472# vss 0.345058f
C800 sarlogic_0/FILLER_0_19_171/a_932_472# vss 0.33241f
C801 sarlogic_0/FILLER_0_19_171/a_484_472# vss 0.33241f
C802 sarlogic_0/FILLER_0_19_171/a_36_472# vss 0.404746f
C803 sarlogic_0/FILLER_0_19_171/a_1468_375# vss 0.233029f
C804 sarlogic_0/FILLER_0_19_171/a_1020_375# vss 0.171606f
C805 sarlogic_0/FILLER_0_19_171/a_572_375# vss 0.171606f
C806 sarlogic_0/FILLER_0_19_171/a_124_375# vss 0.185399f
C807 sarlogic_0/net13 vss 1.176306f
C808 sarlogic_0/net23 vss 2.091399f
C809 sarlogic_0/FILLER_0_20_87/a_36_472# vss 0.417394f
C810 sarlogic_0/FILLER_0_20_87/a_124_375# vss 0.246306f
C811 sarlogic_0/FILLER_0_20_98/a_36_472# vss 0.417394f
C812 sarlogic_0/FILLER_0_20_98/a_124_375# vss 0.246306f
C813 sarlogic_0/_055_ vss 1.782885f
C814 sarlogic_0/FILLER_0_18_53/a_484_472# vss 0.345058f
C815 sarlogic_0/FILLER_0_18_53/a_36_472# vss 0.404746f
C816 sarlogic_0/FILLER_0_18_53/a_572_375# vss 0.232991f
C817 sarlogic_0/FILLER_0_18_53/a_124_375# vss 0.185089f
C818 sarlogic_0/FILLER_0_2_165/a_36_472# vss 0.417394f
C819 sarlogic_0/FILLER_0_2_165/a_124_375# vss 0.246306f
C820 sarlogic_0/FILLER_0_15_205/a_36_472# vss 0.417394f
C821 sarlogic_0/FILLER_0_15_205/a_124_375# vss 0.246306f
C822 sarlogic_0/FILLER_0_23_282/a_484_472# vss 0.345058f
C823 sarlogic_0/FILLER_0_23_282/a_36_472# vss 0.404746f
C824 sarlogic_0/FILLER_0_23_282/a_572_375# vss 0.232991f
C825 sarlogic_0/FILLER_0_23_282/a_124_375# vss 0.185089f
C826 sarlogic_0/net42 vss 1.067446f
C827 sarlogic_0/net17 vss 2.210219f
C828 sarlogic_0/_172_ vss 0.265782f
C829 sarlogic_0/_171_ vss 0.300355f
C830 sarlogic_0/_389_/a_36_148# vss 0.388358f
C831 sarlogic_0/_080_ vss 0.328202f
C832 sarlogic_0/_260_/a_36_68# vss 0.112263f
C833 sarlogic_0/FILLER_0_0_96/a_36_472# vss 0.417394f
C834 sarlogic_0/FILLER_0_0_96/a_124_375# vss 0.246306f
C835 sarlogic_0/FILLER_0_9_72/a_1380_472# vss 0.345058f
C836 sarlogic_0/FILLER_0_9_72/a_932_472# vss 0.33241f
C837 sarlogic_0/FILLER_0_9_72/a_484_472# vss 0.33241f
C838 sarlogic_0/FILLER_0_9_72/a_36_472# vss 0.404746f
C839 sarlogic_0/FILLER_0_9_72/a_1468_375# vss 0.233029f
C840 sarlogic_0/FILLER_0_9_72/a_1020_375# vss 0.171606f
C841 sarlogic_0/FILLER_0_9_72/a_572_375# vss 0.171606f
C842 sarlogic_0/FILLER_0_9_72/a_124_375# vss 0.185399f
C843 sarlogic_0/FILLER_0_20_31/a_36_472# vss 0.417394f
C844 sarlogic_0/FILLER_0_20_31/a_124_375# vss 0.246306f
C845 sarlogic_0/_227_/a_36_160# vss 0.386641f
C846 sarlogic_0/_120_ vss 1.533088f
C847 sarlogic_0/_313_/a_67_603# vss 0.345683f
C848 sarlogic_0/FILLER_0_5_172/a_36_472# vss 0.417394f
C849 sarlogic_0/FILLER_0_5_172/a_124_375# vss 0.246306f
C850 sarlogic_0/FILLER_0_12_20/a_484_472# vss 0.345058f
C851 sarlogic_0/FILLER_0_12_20/a_36_472# vss 0.404746f
C852 sarlogic_0/FILLER_0_12_20/a_572_375# vss 0.232991f
C853 sarlogic_0/FILLER_0_12_20/a_124_375# vss 0.185089f
C854 sarlogic_0/_134_ vss 0.365972f
C855 sarlogic_0/_062_ vss 1.717773f
C856 sarlogic_0/_059_ vss 1.686761f
C857 sarlogic_0/_261_/a_36_160# vss 0.386641f
C858 sarlogic_0/_044_ vss 0.388801f
C859 sarlogic_0/mask\[1\] vss 1.295078f
C860 sarlogic_0/_192_/a_67_603# vss 0.345683f
C861 sarlogic_0/FILLER_0_13_142/a_1380_472# vss 0.345058f
C862 sarlogic_0/FILLER_0_13_142/a_932_472# vss 0.33241f
C863 sarlogic_0/FILLER_0_13_142/a_484_472# vss 0.33241f
C864 sarlogic_0/FILLER_0_13_142/a_36_472# vss 0.404746f
C865 sarlogic_0/FILLER_0_13_142/a_1468_375# vss 0.233029f
C866 sarlogic_0/FILLER_0_13_142/a_1020_375# vss 0.171606f
C867 sarlogic_0/FILLER_0_13_142/a_572_375# vss 0.171606f
C868 sarlogic_0/FILLER_0_13_142/a_124_375# vss 0.185399f
C869 sarlogic_0/FILLER_0_9_60/a_484_472# vss 0.345058f
C870 sarlogic_0/FILLER_0_9_60/a_36_472# vss 0.404746f
C871 sarlogic_0/FILLER_0_9_60/a_572_375# vss 0.232991f
C872 sarlogic_0/FILLER_0_9_60/a_124_375# vss 0.185089f
C873 sarlogic_0/FILLER_0_7_233/a_36_472# vss 0.417394f
C874 sarlogic_0/FILLER_0_7_233/a_124_375# vss 0.246306f
C875 sarlogic_0/_228_/a_36_68# vss 0.69549f
C876 sarlogic_0/FILLER_0_21_206/a_36_472# vss 0.417394f
C877 sarlogic_0/FILLER_0_21_206/a_124_375# vss 0.246306f
C878 sarlogic_0/_067_ vss 0.851951f
C879 sarlogic_0/_135_ vss 0.339478f
C880 sarlogic_0/_193_/a_36_160# vss 0.696445f
C881 sarlogic_0/_180_ vss 0.390598f
C882 sarlogic_0/cal_count\[1\] vss 1.568289f
C883 sarlogic_0/FILLER_0_4_213/a_484_472# vss 0.345058f
C884 sarlogic_0/FILLER_0_4_213/a_36_472# vss 0.404746f
C885 sarlogic_0/FILLER_0_4_213/a_572_375# vss 0.232991f
C886 sarlogic_0/FILLER_0_4_213/a_124_375# vss 0.185089f
C887 sarlogic_0/FILLER_0_11_282/a_36_472# vss 0.417394f
C888 sarlogic_0/FILLER_0_11_282/a_124_375# vss 0.246306f
C889 sarlogic_0/FILLER_0_18_61/a_36_472# vss 0.417394f
C890 sarlogic_0/FILLER_0_18_61/a_124_375# vss 0.246306f
C891 sarlogic_0/FILLER_0_15_235/a_484_472# vss 0.345058f
C892 sarlogic_0/FILLER_0_15_235/a_36_472# vss 0.404746f
C893 sarlogic_0/FILLER_0_15_235/a_572_375# vss 0.232991f
C894 sarlogic_0/FILLER_0_15_235/a_124_375# vss 0.185089f
C895 sarlogic_0/FILLER_0_23_290/a_36_472# vss 0.417394f
C896 sarlogic_0/FILLER_0_23_290/a_124_375# vss 0.246306f
C897 sarlogic_0/_121_ vss 0.532847f
C898 sarlogic_0/_315_/a_36_68# vss 0.052951f
C899 sarlogic_0/_246_/a_36_68# vss 0.69549f
C900 sarlogic_0/FILLER_0_5_181/a_36_472# vss 0.417394f
C901 sarlogic_0/FILLER_0_5_181/a_124_375# vss 0.246306f
C902 sarlogic_0/_082_ vss 0.619901f
C903 sarlogic_0/net8 vss 1.163723f
C904 sarlogic_0/net18 vss 2.032159f
C905 sarlogic_0/_332_/a_36_472# vss 0.031137f
C906 sarlogic_0/_179_ vss 0.336984f
C907 sarlogic_0/_401_/a_36_68# vss 0.112263f
C908 sarlogic_0/FILLER_0_14_107/a_1380_472# vss 0.345058f
C909 sarlogic_0/FILLER_0_14_107/a_932_472# vss 0.33241f
C910 sarlogic_0/FILLER_0_14_107/a_484_472# vss 0.33241f
C911 sarlogic_0/FILLER_0_14_107/a_36_472# vss 0.404746f
C912 sarlogic_0/FILLER_0_14_107/a_1468_375# vss 0.233029f
C913 sarlogic_0/FILLER_0_14_107/a_1020_375# vss 0.171606f
C914 sarlogic_0/FILLER_0_14_107/a_572_375# vss 0.171606f
C915 sarlogic_0/FILLER_0_14_107/a_124_375# vss 0.185399f
C916 sarlogic_0/_097_ vss 0.592554f
C917 sarlogic_0/FILLER_0_1_204/a_36_472# vss 0.417394f
C918 sarlogic_0/FILLER_0_1_204/a_124_375# vss 0.246306f
C919 sarlogic_0/FILLER_0_15_72/a_484_472# vss 0.345058f
C920 sarlogic_0/FILLER_0_15_72/a_36_472# vss 0.404746f
C921 sarlogic_0/FILLER_0_15_72/a_572_375# vss 0.232991f
C922 sarlogic_0/FILLER_0_15_72/a_124_375# vss 0.185089f
C923 sarlogic_0/FILLER_0_17_104/a_1380_472# vss 0.345058f
C924 sarlogic_0/FILLER_0_17_104/a_932_472# vss 0.33241f
C925 sarlogic_0/FILLER_0_17_104/a_484_472# vss 0.33241f
C926 sarlogic_0/FILLER_0_17_104/a_36_472# vss 0.404746f
C927 sarlogic_0/FILLER_0_17_104/a_1468_375# vss 0.233029f
C928 sarlogic_0/FILLER_0_17_104/a_1020_375# vss 0.171606f
C929 sarlogic_0/FILLER_0_17_104/a_572_375# vss 0.171606f
C930 sarlogic_0/FILLER_0_17_104/a_124_375# vss 0.185399f
C931 sarlogic_0/FILLER_0_8_37/a_484_472# vss 0.345058f
C932 sarlogic_0/FILLER_0_8_37/a_36_472# vss 0.404746f
C933 sarlogic_0/FILLER_0_8_37/a_572_375# vss 0.232991f
C934 sarlogic_0/FILLER_0_8_37/a_124_375# vss 0.185089f
C935 sarlogic_0/FILLER_0_15_212/a_1380_472# vss 0.345058f
C936 sarlogic_0/FILLER_0_15_212/a_932_472# vss 0.33241f
C937 sarlogic_0/FILLER_0_15_212/a_484_472# vss 0.33241f
C938 sarlogic_0/FILLER_0_15_212/a_36_472# vss 0.404746f
C939 sarlogic_0/FILLER_0_15_212/a_1468_375# vss 0.233029f
C940 sarlogic_0/FILLER_0_15_212/a_1020_375# vss 0.171606f
C941 sarlogic_0/FILLER_0_15_212/a_572_375# vss 0.171606f
C942 sarlogic_0/FILLER_0_15_212/a_124_375# vss 0.185399f
C943 sarlogic_0/FILLER_0_23_60/a_36_472# vss 0.417394f
C944 sarlogic_0/FILLER_0_23_60/a_124_375# vss 0.246306f
C945 sarlogic_0/_123_ vss 0.344874f
C946 sarlogic_0/_122_ vss 0.600118f
C947 sarlogic_0/calibrate vss 1.343796f
C948 sarlogic_0/_316_/a_848_380# vss 0.40208f
C949 sarlogic_0/_316_/a_124_24# vss 0.591898f
C950 sarlogic_0/_247_/a_36_160# vss 0.696445f
C951 sarlogic_0/FILLER_0_12_50/a_36_472# vss 0.417394f
C952 sarlogic_0/FILLER_0_12_50/a_124_375# vss 0.246306f
C953 sarlogic_0/_084_ vss 0.296163f
C954 sarlogic_0/cal_itt\[0\] vss 1.831055f
C955 sarlogic_0/cal_itt\[1\] vss 1.705665f
C956 sarlogic_0/FILLER_0_11_109/a_36_472# vss 0.417394f
C957 sarlogic_0/FILLER_0_11_109/a_124_375# vss 0.246306f
C958 sarlogic_0/_182_ vss 0.34197f
C959 sarlogic_0/_402_/a_1948_68# vss 0.022025f
C960 sarlogic_0/_402_/a_718_527# vss 0.001795f
C961 sarlogic_0/_402_/a_56_567# vss 0.424713f
C962 sarlogic_0/_402_/a_728_93# vss 0.65929f
C963 sarlogic_0/_402_/a_1296_93# vss 0.317801f
C964 sarlogic_0/_045_ vss 0.349338f
C965 sarlogic_0/mask\[2\] vss 1.335688f
C966 sarlogic_0/_195_/a_67_603# vss 0.345683f
C967 sarlogic_0/_333_/a_36_160# vss 0.386641f
C968 sarlogic_0/_098_ vss 1.816151f
C969 sarlogic_0/_147_ vss 0.322539f
C970 sarlogic_0/_350_/a_49_472# vss 0.054843f
C971 sarlogic_0/FILLER_0_12_236/a_484_472# vss 0.345058f
C972 sarlogic_0/FILLER_0_12_236/a_36_472# vss 0.404746f
C973 sarlogic_0/FILLER_0_12_236/a_572_375# vss 0.232991f
C974 sarlogic_0/FILLER_0_12_236/a_124_375# vss 0.185089f
C975 sarlogic_0/FILLER_0_2_171/a_36_472# vss 0.417394f
C976 sarlogic_0/FILLER_0_2_171/a_124_375# vss 0.246306f
C977 sarlogic_0/_014_ vss 0.363432f
C978 sarlogic_0/_317_/a_36_113# vss 0.418095f
C979 sarlogic_0/_248_/a_36_68# vss 0.69549f
C980 sarlogic_0/FILLER_0_17_38/a_484_472# vss 0.345058f
C981 sarlogic_0/FILLER_0_17_38/a_36_472# vss 0.404746f
C982 sarlogic_0/FILLER_0_17_38/a_572_375# vss 0.232991f
C983 sarlogic_0/FILLER_0_17_38/a_124_375# vss 0.185089f
C984 sarlogic_0/_001_ vss 0.285216f
C985 sarlogic_0/_265_/a_244_68# vss 0.138666f
C986 sarlogic_0/_196_/a_36_160# vss 0.696445f
C987 sarlogic_0/FILLER_0_6_90/a_484_472# vss 0.345058f
C988 sarlogic_0/FILLER_0_6_90/a_36_472# vss 0.404746f
C989 sarlogic_0/FILLER_0_6_90/a_572_375# vss 0.232991f
C990 sarlogic_0/FILLER_0_6_90/a_124_375# vss 0.185089f
C991 sarlogic_0/_183_ vss 0.356629f
C992 sarlogic_0/_334_/a_36_160# vss 0.386641f
C993 sarlogic_0/_282_/a_36_160# vss 0.386641f
C994 sarlogic_0/_024_ vss 0.451815f
C995 sarlogic_0/_009_ vss 0.397943f
C996 sarlogic_0/_420_/a_2560_156# vss 0.016968f
C997 sarlogic_0/_420_/a_2665_112# vss 0.62251f
C998 sarlogic_0/_420_/a_2248_156# vss 0.371662f
C999 sarlogic_0/_420_/a_1204_472# vss 0.012971f
C1000 sarlogic_0/_420_/a_1000_472# vss 0.291735f
C1001 sarlogic_0/_420_/a_796_472# vss 0.023206f
C1002 sarlogic_0/_420_/a_1308_423# vss 0.279043f
C1003 sarlogic_0/_420_/a_448_472# vss 0.684413f
C1004 sarlogic_0/_420_/a_36_151# vss 1.43589f
C1005 clk vss 26.056288f
C1006 sarlogic_0/FILLER_0_8_2/a_36_472# vss 0.417394f
C1007 sarlogic_0/FILLER_0_8_2/a_124_375# vss 0.246306f
C1008 sarlogic_0/FILLER_0_8_24/a_484_472# vss 0.345058f
C1009 sarlogic_0/FILLER_0_8_24/a_36_472# vss 0.404746f
C1010 sarlogic_0/FILLER_0_8_24/a_572_375# vss 0.232991f
C1011 sarlogic_0/FILLER_0_8_24/a_124_375# vss 0.185089f
C1012 sarlogic_0/_124_ vss 0.294081f
C1013 sarlogic_0/_118_ vss 1.378735f
C1014 sarlogic_0/_071_ vss 1.600488f
C1015 sarlogic_0/net9 vss 1.13171f
C1016 sarlogic_0/net19 vss 1.889339f
C1017 sarlogic_0/_138_ vss 0.33132f
C1018 sarlogic_0/_137_ vss 1.178616f
C1019 sarlogic_0/_335_/a_49_472# vss 0.054843f
C1020 sarlogic_0/_404_/a_36_472# vss 0.031137f
C1021 sarlogic_0/FILLER_0_20_107/a_36_472# vss 0.417394f
C1022 sarlogic_0/FILLER_0_20_107/a_124_375# vss 0.246306f
C1023 sarlogic_0/FILLER_0_9_142/a_36_472# vss 0.417394f
C1024 sarlogic_0/FILLER_0_9_142/a_124_375# vss 0.246306f
C1025 sarlogic_0/_099_ vss 1.152785f
C1026 sarlogic_0/_283_/a_36_472# vss 0.031137f
C1027 sarlogic_0/mask\[7\] vss 1.478045f
C1028 sarlogic_0/_352_/a_49_472# vss 0.054843f
C1029 sarlogic_0/_010_ vss 0.377779f
C1030 sarlogic_0/_421_/a_2560_156# vss 0.016968f
C1031 sarlogic_0/_421_/a_2665_112# vss 0.62251f
C1032 sarlogic_0/_421_/a_2248_156# vss 0.371662f
C1033 sarlogic_0/_421_/a_1204_472# vss 0.012971f
C1034 sarlogic_0/_421_/a_1000_472# vss 0.291735f
C1035 sarlogic_0/_421_/a_796_472# vss 0.023206f
C1036 sarlogic_0/_421_/a_1308_423# vss 0.279043f
C1037 sarlogic_0/_421_/a_448_472# vss 0.684413f
C1038 sarlogic_0/_421_/a_36_151# vss 1.43589f
C1039 sarlogic_0/FILLER_0_1_212/a_36_472# vss 0.417394f
C1040 sarlogic_0/FILLER_0_1_212/a_124_375# vss 0.246306f
C1041 sarlogic_0/FILLER_0_8_239/a_36_472# vss 0.417394f
C1042 sarlogic_0/FILLER_0_8_239/a_124_375# vss 0.246306f
C1043 sarlogic_0/_125_ vss 1.526603f
C1044 sarlogic_0/_058_ vss 1.483584f
C1045 sarlogic_0/FILLER_0_6_177/a_484_472# vss 0.345058f
C1046 sarlogic_0/FILLER_0_6_177/a_36_472# vss 0.404746f
C1047 sarlogic_0/FILLER_0_6_177/a_572_375# vss 0.232991f
C1048 sarlogic_0/FILLER_0_6_177/a_124_375# vss 0.185089f
C1049 sarlogic_0/state\[1\] vss 2.652405f
C1050 sarlogic_0/_267_/a_36_472# vss 0.137725f
C1051 sarlogic_0/_184_ vss 0.350066f
C1052 sarlogic_0/cal_count\[2\] vss 1.971854f
C1053 sarlogic_0/_405_/a_67_603# vss 0.345683f
C1054 sarlogic_0/_018_ vss 0.358633f
C1055 sarlogic_0/_046_ vss 0.361963f
C1056 sarlogic_0/_198_/a_67_603# vss 0.345683f
C1057 sarlogic_0/_094_ vss 1.263877f
C1058 sarlogic_0/_100_ vss 0.333135f
C1059 sarlogic_0/net36 vss 2.262756f
C1060 sarlogic_0/FILLER_0_17_133/a_36_472# vss 0.417394f
C1061 sarlogic_0/FILLER_0_17_133/a_124_375# vss 0.246306f
C1062 sarlogic_0/_025_ vss 0.350324f
C1063 sarlogic_0/_148_ vss 0.325709f
C1064 sarlogic_0/_422_/a_2560_156# vss 0.016968f
C1065 sarlogic_0/_422_/a_2665_112# vss 0.62251f
C1066 sarlogic_0/_422_/a_2248_156# vss 0.371662f
C1067 sarlogic_0/_422_/a_1204_472# vss 0.012971f
C1068 sarlogic_0/_422_/a_1000_472# vss 0.291735f
C1069 sarlogic_0/_422_/a_796_472# vss 0.023206f
C1070 sarlogic_0/_422_/a_1308_423# vss 0.279043f
C1071 sarlogic_0/_422_/a_448_472# vss 0.684413f
C1072 sarlogic_0/_422_/a_36_151# vss 1.43589f
C1073 sarlogic_0/FILLER_0_1_266/a_484_472# vss 0.345058f
C1074 sarlogic_0/FILLER_0_1_266/a_36_472# vss 0.404746f
C1075 sarlogic_0/FILLER_0_1_266/a_572_375# vss 0.232991f
C1076 sarlogic_0/FILLER_0_1_266/a_124_375# vss 0.185089f
C1077 sarlogic_0/_152_ vss 0.918583f
C1078 sarlogic_0/_081_ vss 1.140656f
C1079 sarlogic_0/_370_/a_848_380# vss 0.40208f
C1080 sarlogic_0/_370_/a_124_24# vss 0.591898f
C1081 sarlogic_0/FILLER_0_24_274/a_1380_472# vss 0.345058f
C1082 sarlogic_0/FILLER_0_24_274/a_932_472# vss 0.33241f
C1083 sarlogic_0/FILLER_0_24_274/a_484_472# vss 0.33241f
C1084 sarlogic_0/FILLER_0_24_274/a_36_472# vss 0.404746f
C1085 sarlogic_0/FILLER_0_24_274/a_1468_375# vss 0.233029f
C1086 sarlogic_0/FILLER_0_24_274/a_1020_375# vss 0.171606f
C1087 sarlogic_0/FILLER_0_24_274/a_572_375# vss 0.171606f
C1088 sarlogic_0/FILLER_0_24_274/a_124_375# vss 0.185399f
C1089 sarlogic_0/_185_ vss 0.386917f
C1090 sarlogic_0/_406_/a_36_159# vss 0.374116f
C1091 sarlogic_0/_337_/a_49_472# vss 0.054843f
C1092 sarlogic_0/_199_/a_36_160# vss 0.696445f
C1093 sarlogic_0/_285_/a_36_472# vss 0.031137f
C1094 sarlogic_0/_354_/a_49_472# vss 0.054843f
C1095 sarlogic_0/_012_ vss 0.75195f
C1096 sarlogic_0/_423_/a_2560_156# vss 0.016968f
C1097 sarlogic_0/_423_/a_2665_112# vss 0.62251f
C1098 sarlogic_0/_423_/a_2248_156# vss 0.371662f
C1099 sarlogic_0/_423_/a_1204_472# vss 0.012971f
C1100 sarlogic_0/_423_/a_1000_472# vss 0.291735f
C1101 sarlogic_0/_423_/a_796_472# vss 0.023206f
C1102 sarlogic_0/_423_/a_1308_423# vss 0.279043f
C1103 sarlogic_0/_423_/a_448_472# vss 0.684413f
C1104 sarlogic_0/_423_/a_36_151# vss 1.43589f
C1105 sarlogic_0/FILLER_0_5_88/a_36_472# vss 0.417394f
C1106 sarlogic_0/FILLER_0_5_88/a_124_375# vss 0.246306f
C1107 sarlogic_0/trim_mask\[1\] vss 1.020743f
C1108 sarlogic_0/_029_ vss 0.308904f
C1109 sarlogic_0/_440_/a_2560_156# vss 0.016968f
C1110 sarlogic_0/_440_/a_2665_112# vss 0.62251f
C1111 sarlogic_0/_440_/a_2248_156# vss 0.371662f
C1112 sarlogic_0/_440_/a_1204_472# vss 0.012971f
C1113 sarlogic_0/_440_/a_1000_472# vss 0.291735f
C1114 sarlogic_0/_440_/a_796_472# vss 0.023206f
C1115 sarlogic_0/_440_/a_1308_423# vss 0.279043f
C1116 sarlogic_0/_440_/a_448_472# vss 0.684413f
C1117 sarlogic_0/_440_/a_36_151# vss 1.43589f
C1118 sarlogic_0/_159_ vss 0.351814f
C1119 sarlogic_0/_371_/a_36_113# vss 0.418095f
C1120 sarlogic_0/FILLER_0_17_56/a_484_472# vss 0.345058f
C1121 sarlogic_0/FILLER_0_17_56/a_36_472# vss 0.404746f
C1122 sarlogic_0/FILLER_0_17_56/a_572_375# vss 0.232991f
C1123 sarlogic_0/FILLER_0_17_56/a_124_375# vss 0.185089f
C1124 sarlogic_0/_083_ vss 0.527882f
C1125 sarlogic_0/_078_ vss 0.904554f
C1126 sarlogic_0/_269_/a_36_472# vss 0.031137f
C1127 sarlogic_0/_181_ vss 0.829168f
C1128 sarlogic_0/_407_/a_36_472# vss 0.031137f
C1129 sarlogic_0/_019_ vss 0.32907f
C1130 sarlogic_0/_139_ vss 0.346404f
C1131 sarlogic_0/FILLER_0_14_123/a_36_472# vss 0.417394f
C1132 sarlogic_0/FILLER_0_14_123/a_124_375# vss 0.246306f
C1133 sarlogic_0/_005_ vss 0.340993f
C1134 sarlogic_0/_101_ vss 0.280497f
C1135 sarlogic_0/_424_/a_2560_156# vss 0.016968f
C1136 sarlogic_0/_424_/a_2665_112# vss 0.62251f
C1137 sarlogic_0/_424_/a_2248_156# vss 0.371662f
C1138 sarlogic_0/_424_/a_1204_472# vss 0.012971f
C1139 sarlogic_0/_424_/a_1000_472# vss 0.291735f
C1140 sarlogic_0/_424_/a_796_472# vss 0.023206f
C1141 sarlogic_0/_424_/a_1308_423# vss 0.279043f
C1142 sarlogic_0/_424_/a_448_472# vss 0.684413f
C1143 sarlogic_0/_424_/a_36_151# vss 1.43589f
C1144 sarlogic_0/_026_ vss 0.320379f
C1145 sarlogic_0/_149_ vss 0.305496f
C1146 sarlogic_0/FILLER_0_5_54/a_1380_472# vss 0.345058f
C1147 sarlogic_0/FILLER_0_5_54/a_932_472# vss 0.33241f
C1148 sarlogic_0/FILLER_0_5_54/a_484_472# vss 0.33241f
C1149 sarlogic_0/FILLER_0_5_54/a_36_472# vss 0.404746f
C1150 sarlogic_0/FILLER_0_5_54/a_1468_375# vss 0.233029f
C1151 sarlogic_0/FILLER_0_5_54/a_1020_375# vss 0.171606f
C1152 sarlogic_0/FILLER_0_5_54/a_572_375# vss 0.171606f
C1153 sarlogic_0/FILLER_0_5_54/a_124_375# vss 0.185399f
C1154 sarlogic_0/FILLER_0_17_142/a_484_472# vss 0.345058f
C1155 sarlogic_0/FILLER_0_17_142/a_36_472# vss 0.404746f
C1156 sarlogic_0/FILLER_0_17_142/a_572_375# vss 0.232991f
C1157 sarlogic_0/FILLER_0_17_142/a_124_375# vss 0.185089f
C1158 sarlogic_0/_068_ vss 3.162692f
C1159 sarlogic_0/_076_ vss 3.812442f
C1160 sarlogic_0/_133_ vss 1.430901f
C1161 sarlogic_0/_070_ vss 3.115722f
C1162 sarlogic_0/_372_/a_170_472# vss 0.077257f
C1163 sarlogic_0/net49 vss 5.140563f
C1164 sarlogic_0/_030_ vss 0.307083f
C1165 sarlogic_0/net66 vss 1.472669f
C1166 sarlogic_0/_441_/a_2560_156# vss 0.016968f
C1167 sarlogic_0/_441_/a_2665_112# vss 0.62251f
C1168 sarlogic_0/_441_/a_2248_156# vss 0.371662f
C1169 sarlogic_0/_441_/a_1204_472# vss 0.012971f
C1170 sarlogic_0/_441_/a_1000_472# vss 0.291735f
C1171 sarlogic_0/_441_/a_796_472# vss 0.023206f
C1172 sarlogic_0/_441_/a_1308_423# vss 0.279043f
C1173 sarlogic_0/_441_/a_448_472# vss 0.684413f
C1174 sarlogic_0/_441_/a_36_151# vss 1.43589f
C1175 sarlogic_0/FILLER_0_5_206/a_36_472# vss 0.417394f
C1176 sarlogic_0/FILLER_0_5_206/a_124_375# vss 0.246306f
C1177 sarlogic_0/fanout49/a_36_160# vss 0.696445f
C1178 sarlogic_0/FILLER_0_8_247/a_1380_472# vss 0.345058f
C1179 sarlogic_0/FILLER_0_8_247/a_932_472# vss 0.33241f
C1180 sarlogic_0/FILLER_0_8_247/a_484_472# vss 0.33241f
C1181 sarlogic_0/FILLER_0_8_247/a_36_472# vss 0.404746f
C1182 sarlogic_0/FILLER_0_8_247/a_1468_375# vss 0.233029f
C1183 sarlogic_0/FILLER_0_8_247/a_1020_375# vss 0.171606f
C1184 sarlogic_0/FILLER_0_8_247/a_572_375# vss 0.171606f
C1185 sarlogic_0/FILLER_0_8_247/a_124_375# vss 0.185399f
C1186 sarlogic_0/FILLER_0_12_220/a_1380_472# vss 0.345058f
C1187 sarlogic_0/FILLER_0_12_220/a_932_472# vss 0.33241f
C1188 sarlogic_0/FILLER_0_12_220/a_484_472# vss 0.33241f
C1189 sarlogic_0/FILLER_0_12_220/a_36_472# vss 0.404746f
C1190 sarlogic_0/FILLER_0_12_220/a_1468_375# vss 0.233029f
C1191 sarlogic_0/FILLER_0_12_220/a_1020_375# vss 0.171606f
C1192 sarlogic_0/FILLER_0_12_220/a_572_375# vss 0.171606f
C1193 sarlogic_0/FILLER_0_12_220/a_124_375# vss 0.185399f
C1194 sarlogic_0/FILLER_0_21_286/a_484_472# vss 0.345058f
C1195 sarlogic_0/FILLER_0_21_286/a_36_472# vss 0.404746f
C1196 sarlogic_0/FILLER_0_21_286/a_572_375# vss 0.232991f
C1197 sarlogic_0/FILLER_0_21_286/a_124_375# vss 0.185089f
C1198 sarlogic_0/_140_ vss 1.276518f
C1199 sarlogic_0/_339_/a_36_160# vss 0.386641f
C1200 sarlogic_0/_095_ vss 2.689027f
C1201 sarlogic_0/_186_ vss 0.580923f
C1202 sarlogic_0/_408_/a_1936_472# vss 0.009918f
C1203 sarlogic_0/_408_/a_718_524# vss 0.005143f
C1204 sarlogic_0/_408_/a_56_524# vss 0.41096f
C1205 sarlogic_0/_408_/a_728_93# vss 0.654825f
C1206 sarlogic_0/_408_/a_1336_472# vss 0.316639f
C1207 sarlogic_0/FILLER_0_20_169/a_36_472# vss 0.417394f
C1208 sarlogic_0/FILLER_0_20_169/a_124_375# vss 0.246306f
C1209 sarlogic_0/_210_/a_67_603# vss 0.345683f
C1210 sarlogic_0/_425_/a_2560_156# vss 0.016968f
C1211 sarlogic_0/_425_/a_2665_112# vss 0.62251f
C1212 sarlogic_0/_425_/a_2248_156# vss 0.371662f
C1213 sarlogic_0/_425_/a_1204_472# vss 0.012971f
C1214 sarlogic_0/_425_/a_1000_472# vss 0.291735f
C1215 sarlogic_0/_425_/a_796_472# vss 0.023206f
C1216 sarlogic_0/_425_/a_1308_423# vss 0.279043f
C1217 sarlogic_0/_425_/a_448_472# vss 0.684413f
C1218 sarlogic_0/_425_/a_36_151# vss 1.43589f
C1219 sarlogic_0/net5 vss 0.610761f
C1220 sarlogic_0/input5/a_36_113# vss 0.418095f
C1221 sarlogic_0/FILLER_0_11_78/a_484_472# vss 0.345058f
C1222 sarlogic_0/FILLER_0_11_78/a_36_472# vss 0.404746f
C1223 sarlogic_0/FILLER_0_11_78/a_572_375# vss 0.232991f
C1224 sarlogic_0/FILLER_0_11_78/a_124_375# vss 0.185089f
C1225 sarlogic_0/_102_ vss 0.335308f
C1226 sarlogic_0/_287_/a_36_472# vss 0.031137f
C1227 sarlogic_0/mask\[9\] vss 1.383606f
C1228 sarlogic_0/_356_/a_36_472# vss 0.031137f
C1229 sarlogic_0/_031_ vss 0.417351f
C1230 sarlogic_0/net69 vss 1.020293f
C1231 sarlogic_0/_442_/a_2560_156# vss 0.016968f
C1232 sarlogic_0/_442_/a_2665_112# vss 0.62251f
C1233 sarlogic_0/_442_/a_2248_156# vss 0.371662f
C1234 sarlogic_0/_442_/a_1204_472# vss 0.012971f
C1235 sarlogic_0/_442_/a_1000_472# vss 0.291735f
C1236 sarlogic_0/_442_/a_796_472# vss 0.023206f
C1237 sarlogic_0/_442_/a_1308_423# vss 0.279043f
C1238 sarlogic_0/_442_/a_448_472# vss 0.684413f
C1239 sarlogic_0/_442_/a_36_151# vss 1.43589f
C1240 sarlogic_0/net64 vss 2.598514f
C1241 sarlogic_0/fanout59/a_36_160# vss 0.696445f
C1242 sarlogic_0/FILLER_0_14_99/a_36_472# vss 0.417394f
C1243 sarlogic_0/FILLER_0_14_99/a_124_375# vss 0.246306f
C1244 sarlogic_0/_038_ vss 0.362839f
C1245 sarlogic_0/_136_ vss 1.345638f
C1246 sarlogic_0/_390_/a_36_68# vss 0.150048f
C1247 sarlogic_0/FILLER_0_15_282/a_484_472# vss 0.345058f
C1248 sarlogic_0/FILLER_0_15_282/a_36_472# vss 0.404746f
C1249 sarlogic_0/FILLER_0_15_282/a_572_375# vss 0.232991f
C1250 sarlogic_0/FILLER_0_15_282/a_124_375# vss 0.185089f
C1251 sarlogic_0/FILLER_0_11_124/a_36_472# vss 0.417394f
C1252 sarlogic_0/FILLER_0_11_124/a_124_375# vss 0.246306f
C1253 sarlogic_0/FILLER_0_11_135/a_36_472# vss 0.417394f
C1254 sarlogic_0/FILLER_0_11_135/a_124_375# vss 0.246306f
C1255 sarlogic_0/_188_ vss 0.349407f
C1256 sarlogic_0/cal_count\[3\] vss 1.862896f
C1257 sarlogic_0/_050_ vss 0.622354f
C1258 sarlogic_0/_211_/a_36_160# vss 0.386641f
C1259 sarlogic_0/net4 vss 2.711508f
C1260 en vss 25.538645f
C1261 sarlogic_0/input4/a_36_68# vss 0.69549f
C1262 sarlogic_0/_426_/a_2560_156# vss 0.016968f
C1263 sarlogic_0/_426_/a_2665_112# vss 0.62251f
C1264 sarlogic_0/_426_/a_2248_156# vss 0.371662f
C1265 sarlogic_0/_426_/a_1204_472# vss 0.012971f
C1266 sarlogic_0/_426_/a_1000_472# vss 0.291735f
C1267 sarlogic_0/_426_/a_796_472# vss 0.023206f
C1268 sarlogic_0/_426_/a_1308_423# vss 0.279043f
C1269 sarlogic_0/_426_/a_448_472# vss 0.684413f
C1270 sarlogic_0/_426_/a_36_151# vss 1.43589f
C1271 sarlogic_0/_027_ vss 0.302949f
C1272 sarlogic_0/_150_ vss 0.320497f
C1273 sarlogic_0/FILLER_0_18_107/a_3172_472# vss 0.345058f
C1274 sarlogic_0/FILLER_0_18_107/a_2724_472# vss 0.33241f
C1275 sarlogic_0/FILLER_0_18_107/a_2276_472# vss 0.33241f
C1276 sarlogic_0/FILLER_0_18_107/a_1828_472# vss 0.33241f
C1277 sarlogic_0/FILLER_0_18_107/a_1380_472# vss 0.33241f
C1278 sarlogic_0/FILLER_0_18_107/a_932_472# vss 0.33241f
C1279 sarlogic_0/FILLER_0_18_107/a_484_472# vss 0.33241f
C1280 sarlogic_0/FILLER_0_18_107/a_36_472# vss 0.404746f
C1281 sarlogic_0/FILLER_0_18_107/a_3260_375# vss 0.233093f
C1282 sarlogic_0/FILLER_0_18_107/a_2812_375# vss 0.17167f
C1283 sarlogic_0/FILLER_0_18_107/a_2364_375# vss 0.17167f
C1284 sarlogic_0/FILLER_0_18_107/a_1916_375# vss 0.17167f
C1285 sarlogic_0/FILLER_0_18_107/a_1468_375# vss 0.17167f
C1286 sarlogic_0/FILLER_0_18_107/a_1020_375# vss 0.17167f
C1287 sarlogic_0/FILLER_0_18_107/a_572_375# vss 0.17167f
C1288 sarlogic_0/FILLER_0_18_107/a_124_375# vss 0.185915f
C1289 sarlogic_0/trim_mask\[4\] vss 0.987791f
C1290 sarlogic_0/_032_ vss 0.34876f
C1291 sarlogic_0/_443_/a_2560_156# vss 0.016968f
C1292 sarlogic_0/_443_/a_2665_112# vss 0.62251f
C1293 sarlogic_0/_443_/a_2248_156# vss 0.371662f
C1294 sarlogic_0/_443_/a_1204_472# vss 0.012971f
C1295 sarlogic_0/_443_/a_1000_472# vss 0.291735f
C1296 sarlogic_0/_443_/a_796_472# vss 0.023206f
C1297 sarlogic_0/_443_/a_1308_423# vss 0.279043f
C1298 sarlogic_0/_443_/a_448_472# vss 0.684413f
C1299 sarlogic_0/_443_/a_36_151# vss 1.43589f
C1300 sarlogic_0/_061_ vss 0.84986f
C1301 sarlogic_0/_056_ vss 2.393362f
C1302 sarlogic_0/_374_/a_36_68# vss 0.112263f
C1303 sarlogic_0/fanout58/a_36_160# vss 0.696445f
C1304 sarlogic_0/net74 vss 1.237373f
C1305 sarlogic_0/fanout69/a_36_113# vss 0.418095f
C1306 sarlogic_0/_173_ vss 0.339446f
C1307 sarlogic_0/FILLER_0_3_142/a_36_472# vss 0.417394f
C1308 sarlogic_0/FILLER_0_3_142/a_124_375# vss 0.246306f
C1309 sarlogic_0/FILLER_0_17_64/a_36_472# vss 0.417394f
C1310 sarlogic_0/FILLER_0_17_64/a_124_375# vss 0.246306f
C1311 sarlogic_0/FILLER_0_11_101/a_484_472# vss 0.345058f
C1312 sarlogic_0/FILLER_0_11_101/a_36_472# vss 0.404746f
C1313 sarlogic_0/FILLER_0_11_101/a_572_375# vss 0.232991f
C1314 sarlogic_0/FILLER_0_11_101/a_124_375# vss 0.185089f
C1315 sarlogic_0/FILLER_0_22_86/a_1380_472# vss 0.345058f
C1316 sarlogic_0/FILLER_0_22_86/a_932_472# vss 0.33241f
C1317 sarlogic_0/FILLER_0_22_86/a_484_472# vss 0.33241f
C1318 sarlogic_0/FILLER_0_22_86/a_36_472# vss 0.404746f
C1319 sarlogic_0/FILLER_0_22_86/a_1468_375# vss 0.233029f
C1320 sarlogic_0/FILLER_0_22_86/a_1020_375# vss 0.171606f
C1321 sarlogic_0/FILLER_0_22_86/a_572_375# vss 0.171606f
C1322 sarlogic_0/FILLER_0_22_86/a_124_375# vss 0.185399f
C1323 sarlogic_0/net24 vss 1.61895f
C1324 sarlogic_0/net3 vss 0.740676f
C1325 sarlogic_0/input3/a_36_113# vss 0.418095f
C1326 sarlogic_0/_103_ vss 0.350464f
C1327 sarlogic_0/_289_/a_36_472# vss 0.031137f
C1328 sarlogic_0/_151_ vss 0.300777f
C1329 sarlogic_0/_427_/a_2560_156# vss 0.016968f
C1330 sarlogic_0/_427_/a_2665_112# vss 0.91969f
C1331 sarlogic_0/_427_/a_2248_156# vss 0.30886f
C1332 sarlogic_0/_427_/a_1204_472# vss 0.012971f
C1333 sarlogic_0/_427_/a_1000_472# vss 0.291735f
C1334 sarlogic_0/_427_/a_796_472# vss 0.023206f
C1335 sarlogic_0/_427_/a_1308_423# vss 0.279043f
C1336 sarlogic_0/_427_/a_448_472# vss 0.684413f
C1337 sarlogic_0/_427_/a_36_151# vss 1.43587f
C1338 sarlogic_0/FILLER_0_17_161/a_36_472# vss 0.417394f
C1339 sarlogic_0/FILLER_0_17_161/a_124_375# vss 0.246306f
C1340 sarlogic_0/FILLER_0_18_139/a_1380_472# vss 0.345058f
C1341 sarlogic_0/FILLER_0_18_139/a_932_472# vss 0.33241f
C1342 sarlogic_0/FILLER_0_18_139/a_484_472# vss 0.33241f
C1343 sarlogic_0/FILLER_0_18_139/a_36_472# vss 0.404746f
C1344 sarlogic_0/FILLER_0_18_139/a_1468_375# vss 0.233029f
C1345 sarlogic_0/FILLER_0_18_139/a_1020_375# vss 0.171606f
C1346 sarlogic_0/FILLER_0_18_139/a_572_375# vss 0.171606f
C1347 sarlogic_0/FILLER_0_18_139/a_124_375# vss 0.185399f
C1348 sarlogic_0/_161_ vss 0.592909f
C1349 sarlogic_0/_162_ vss 0.597238f
C1350 sarlogic_0/_375_/a_36_68# vss 0.048026f
C1351 sarlogic_0/trim_val\[0\] vss 0.742779f
C1352 sarlogic_0/net67 vss 1.662327f
C1353 sarlogic_0/_444_/a_2560_156# vss 0.016968f
C1354 sarlogic_0/_444_/a_2665_112# vss 0.62251f
C1355 sarlogic_0/_444_/a_2248_156# vss 0.371662f
C1356 sarlogic_0/_444_/a_1204_472# vss 0.012971f
C1357 sarlogic_0/_444_/a_1000_472# vss 0.291735f
C1358 sarlogic_0/_444_/a_796_472# vss 0.023206f
C1359 sarlogic_0/_444_/a_1308_423# vss 0.279043f
C1360 sarlogic_0/_444_/a_448_472# vss 0.684413f
C1361 sarlogic_0/_444_/a_36_151# vss 1.43589f
C1362 sarlogic_0/net65 vss 0.804072f
C1363 sarlogic_0/fanout57/a_36_113# vss 0.418095f
C1364 sarlogic_0/fanout68/a_36_113# vss 0.418095f
C1365 sarlogic_0/FILLER_0_12_2/a_484_472# vss 0.345058f
C1366 sarlogic_0/FILLER_0_12_2/a_36_472# vss 0.404746f
C1367 sarlogic_0/FILLER_0_12_2/a_572_375# vss 0.232991f
C1368 sarlogic_0/FILLER_0_12_2/a_124_375# vss 0.185089f
C1369 sarlogic_0/net79 vss 1.584979f
C1370 sarlogic_0/fanout79/a_36_160# vss 0.386641f
C1371 sarlogic_0/_392_/a_36_68# vss 0.112263f
C1372 sarlogic_0/FILLER_0_13_228/a_36_472# vss 0.417394f
C1373 sarlogic_0/FILLER_0_13_228/a_124_375# vss 0.246306f
C1374 sarlogic_0/FILLER_0_13_206/a_36_472# vss 0.417394f
C1375 sarlogic_0/FILLER_0_13_206/a_124_375# vss 0.246306f
C1376 sarlogic_0/FILLER_0_20_177/a_1380_472# vss 0.345058f
C1377 sarlogic_0/FILLER_0_20_177/a_932_472# vss 0.33241f
C1378 sarlogic_0/FILLER_0_20_177/a_484_472# vss 0.33241f
C1379 sarlogic_0/FILLER_0_20_177/a_36_472# vss 0.404746f
C1380 sarlogic_0/FILLER_0_20_177/a_1468_375# vss 0.233029f
C1381 sarlogic_0/FILLER_0_20_177/a_1020_375# vss 0.171606f
C1382 sarlogic_0/FILLER_0_20_177/a_572_375# vss 0.171606f
C1383 sarlogic_0/FILLER_0_20_177/a_124_375# vss 0.185399f
C1384 sarlogic_0/_051_ vss 0.349381f
C1385 sarlogic_0/_213_/a_67_603# vss 0.345683f
C1386 sarlogic_0/net2 vss 0.461658f
C1387 sarlogic_0/input2/a_36_113# vss 0.418095f
C1388 sarlogic_0/_129_ vss 0.926508f
C1389 sarlogic_0/_131_ vss 1.734297f
C1390 sarlogic_0/_359_/a_36_488# vss 0.101145f
C1391 sarlogic_0/FILLER_0_11_64/a_36_472# vss 0.417394f
C1392 sarlogic_0/FILLER_0_11_64/a_124_375# vss 0.246306f
C1393 sarlogic_0/state\[2\] vss 0.607433f
C1394 sarlogic_0/net53 vss 4.483899f
C1395 sarlogic_0/_017_ vss 0.334329f
C1396 sarlogic_0/net70 vss 1.238296f
C1397 sarlogic_0/_428_/a_2560_156# vss 0.016968f
C1398 sarlogic_0/_428_/a_2665_112# vss 0.62251f
C1399 sarlogic_0/_428_/a_2248_156# vss 0.371662f
C1400 sarlogic_0/_428_/a_1204_472# vss 0.012971f
C1401 sarlogic_0/_428_/a_1000_472# vss 0.291735f
C1402 sarlogic_0/_428_/a_796_472# vss 0.023206f
C1403 sarlogic_0/_428_/a_1308_423# vss 0.279043f
C1404 sarlogic_0/_428_/a_448_472# vss 0.684413f
C1405 sarlogic_0/_428_/a_36_151# vss 1.43589f
C1406 sarlogic_0/FILLER_0_5_72/a_1380_472# vss 0.345058f
C1407 sarlogic_0/FILLER_0_5_72/a_932_472# vss 0.33241f
C1408 sarlogic_0/FILLER_0_5_72/a_484_472# vss 0.33241f
C1409 sarlogic_0/FILLER_0_5_72/a_36_472# vss 0.404746f
C1410 sarlogic_0/FILLER_0_5_72/a_1468_375# vss 0.233029f
C1411 sarlogic_0/FILLER_0_5_72/a_1020_375# vss 0.171606f
C1412 sarlogic_0/FILLER_0_5_72/a_572_375# vss 0.171606f
C1413 sarlogic_0/FILLER_0_5_72/a_124_375# vss 0.185399f
C1414 sarlogic_0/_376_/a_36_160# vss 0.386641f
C1415 sarlogic_0/trim_val\[1\] vss 0.683578f
C1416 sarlogic_0/_445_/a_2560_156# vss 0.016968f
C1417 sarlogic_0/_445_/a_2665_112# vss 0.62251f
C1418 sarlogic_0/_445_/a_2248_156# vss 0.371662f
C1419 sarlogic_0/_445_/a_1204_472# vss 0.012971f
C1420 sarlogic_0/_445_/a_1000_472# vss 0.291735f
C1421 sarlogic_0/_445_/a_796_472# vss 0.023206f
C1422 sarlogic_0/_445_/a_1308_423# vss 0.279043f
C1423 sarlogic_0/_445_/a_448_472# vss 0.684413f
C1424 sarlogic_0/_445_/a_36_151# vss 1.43589f
C1425 sarlogic_0/fanout67/a_36_160# vss 0.386641f
C1426 sarlogic_0/fanout56/a_36_113# vss 0.418095f
C1427 sarlogic_0/net78 vss 0.686263f
C1428 sarlogic_0/fanout78/a_36_113# vss 0.418095f
C1429 sarlogic_0/_174_ vss 0.979741f
C1430 sarlogic_0/FILLER_0_0_198/a_36_472# vss 0.417394f
C1431 sarlogic_0/FILLER_0_0_198/a_124_375# vss 0.246306f
C1432 sarlogic_0/FILLER_0_15_290/a_36_472# vss 0.417394f
C1433 sarlogic_0/FILLER_0_15_290/a_124_375# vss 0.246306f
C1434 sarlogic_0/FILLER_0_24_290/a_36_472# vss 0.417394f
C1435 sarlogic_0/FILLER_0_24_290/a_124_375# vss 0.246306f
C1436 sarlogic_0/FILLER_0_4_107/a_1380_472# vss 0.345058f
C1437 sarlogic_0/FILLER_0_4_107/a_932_472# vss 0.33241f
C1438 sarlogic_0/FILLER_0_4_107/a_484_472# vss 0.33241f
C1439 sarlogic_0/FILLER_0_4_107/a_36_472# vss 0.404746f
C1440 sarlogic_0/FILLER_0_4_107/a_1468_375# vss 0.233029f
C1441 sarlogic_0/FILLER_0_4_107/a_1020_375# vss 0.171606f
C1442 sarlogic_0/FILLER_0_4_107/a_572_375# vss 0.171606f
C1443 sarlogic_0/FILLER_0_4_107/a_124_375# vss 0.185399f
C1444 sarlogic_0/FILLER_0_7_104/a_1380_472# vss 0.345058f
C1445 sarlogic_0/FILLER_0_7_104/a_932_472# vss 0.33241f
C1446 sarlogic_0/FILLER_0_7_104/a_484_472# vss 0.33241f
C1447 sarlogic_0/FILLER_0_7_104/a_36_472# vss 0.404746f
C1448 sarlogic_0/FILLER_0_7_104/a_1468_375# vss 0.233029f
C1449 sarlogic_0/FILLER_0_7_104/a_1020_375# vss 0.171606f
C1450 sarlogic_0/FILLER_0_7_104/a_572_375# vss 0.171606f
C1451 sarlogic_0/FILLER_0_7_104/a_124_375# vss 0.185399f
C1452 sarlogic_0/_214_/a_36_160# vss 0.386641f
C1453 sarlogic_0/net1 vss 0.364811f
C1454 sarlogic_0/input1/a_36_113# vss 0.418095f
C1455 sarlogic_0/_429_/a_2560_156# vss 0.016968f
C1456 sarlogic_0/_429_/a_2665_112# vss 0.62251f
C1457 sarlogic_0/_429_/a_2248_156# vss 0.371662f
C1458 sarlogic_0/_429_/a_1204_472# vss 0.012971f
C1459 sarlogic_0/_429_/a_1000_472# vss 0.291735f
C1460 sarlogic_0/_429_/a_796_472# vss 0.023206f
C1461 sarlogic_0/_429_/a_1308_423# vss 0.279043f
C1462 sarlogic_0/_429_/a_448_472# vss 0.684413f
C1463 sarlogic_0/_429_/a_36_151# vss 1.43589f
C1464 sarlogic_0/_011_ vss 0.278979f
C1465 sarlogic_0/_377_/a_36_472# vss 0.031137f
C1466 sarlogic_0/fanout66/a_36_113# vss 0.418095f
C1467 sarlogic_0/_035_ vss 0.327801f
C1468 sarlogic_0/_446_/a_2560_156# vss 0.016968f
C1469 sarlogic_0/_446_/a_2665_112# vss 0.62251f
C1470 sarlogic_0/_446_/a_2248_156# vss 0.371662f
C1471 sarlogic_0/_446_/a_1204_472# vss 0.012971f
C1472 sarlogic_0/_446_/a_1000_472# vss 0.291735f
C1473 sarlogic_0/_446_/a_796_472# vss 0.023206f
C1474 sarlogic_0/_446_/a_1308_423# vss 0.279043f
C1475 sarlogic_0/_446_/a_448_472# vss 0.684413f
C1476 sarlogic_0/_446_/a_36_151# vss 1.43589f
C1477 sarlogic_0/fanout77/a_36_113# vss 0.418095f
C1478 sarlogic_0/FILLER_0_5_212/a_36_472# vss 0.417394f
C1479 sarlogic_0/FILLER_0_5_212/a_124_375# vss 0.246306f
C1480 sarlogic_0/fanout55/a_36_160# vss 0.696445f
C1481 sarlogic_0/_175_ vss 0.344159f
C1482 sarlogic_0/_394_/a_1936_472# vss 0.009918f
C1483 sarlogic_0/_394_/a_718_524# vss 0.005143f
C1484 sarlogic_0/_394_/a_56_524# vss 0.41096f
C1485 sarlogic_0/_394_/a_728_93# vss 0.654825f
C1486 sarlogic_0/_394_/a_1336_472# vss 0.316639f
C1487 sarlogic_0/FILLER_0_3_172/a_3172_472# vss 0.345058f
C1488 sarlogic_0/FILLER_0_3_172/a_2724_472# vss 0.33241f
C1489 sarlogic_0/FILLER_0_3_172/a_2276_472# vss 0.33241f
C1490 sarlogic_0/FILLER_0_3_172/a_1828_472# vss 0.33241f
C1491 sarlogic_0/FILLER_0_3_172/a_1380_472# vss 0.33241f
C1492 sarlogic_0/FILLER_0_3_172/a_932_472# vss 0.33241f
C1493 sarlogic_0/FILLER_0_3_172/a_484_472# vss 0.33241f
C1494 sarlogic_0/FILLER_0_3_172/a_36_472# vss 0.404746f
C1495 sarlogic_0/FILLER_0_3_172/a_3260_375# vss 0.233093f
C1496 sarlogic_0/FILLER_0_3_172/a_2812_375# vss 0.17167f
C1497 sarlogic_0/FILLER_0_3_172/a_2364_375# vss 0.17167f
C1498 sarlogic_0/FILLER_0_3_172/a_1916_375# vss 0.17167f
C1499 sarlogic_0/FILLER_0_3_172/a_1468_375# vss 0.17167f
C1500 sarlogic_0/FILLER_0_3_172/a_1020_375# vss 0.17167f
C1501 sarlogic_0/FILLER_0_3_172/a_572_375# vss 0.17167f
C1502 sarlogic_0/FILLER_0_3_172/a_124_375# vss 0.185915f
C1503 sarlogic_0/FILLER_0_17_72/a_3172_472# vss 0.345058f
C1504 sarlogic_0/FILLER_0_17_72/a_2724_472# vss 0.33241f
C1505 sarlogic_0/FILLER_0_17_72/a_2276_472# vss 0.33241f
C1506 sarlogic_0/FILLER_0_17_72/a_1828_472# vss 0.33241f
C1507 sarlogic_0/FILLER_0_17_72/a_1380_472# vss 0.33241f
C1508 sarlogic_0/FILLER_0_17_72/a_932_472# vss 0.33241f
C1509 sarlogic_0/FILLER_0_17_72/a_484_472# vss 0.33241f
C1510 sarlogic_0/FILLER_0_17_72/a_36_472# vss 0.404746f
C1511 sarlogic_0/FILLER_0_17_72/a_3260_375# vss 0.233093f
C1512 sarlogic_0/FILLER_0_17_72/a_2812_375# vss 0.17167f
C1513 sarlogic_0/FILLER_0_17_72/a_2364_375# vss 0.17167f
C1514 sarlogic_0/FILLER_0_17_72/a_1916_375# vss 0.17167f
C1515 sarlogic_0/FILLER_0_17_72/a_1468_375# vss 0.17167f
C1516 sarlogic_0/FILLER_0_17_72/a_1020_375# vss 0.17167f
C1517 sarlogic_0/FILLER_0_17_72/a_572_375# vss 0.17167f
C1518 sarlogic_0/FILLER_0_17_72/a_124_375# vss 0.185915f
C1519 sarlogic_0/FILLER_0_2_93/a_484_472# vss 0.345058f
C1520 sarlogic_0/FILLER_0_2_93/a_36_472# vss 0.404746f
C1521 sarlogic_0/FILLER_0_2_93/a_572_375# vss 0.232991f
C1522 sarlogic_0/FILLER_0_2_93/a_124_375# vss 0.185089f
C1523 sarlogic_0/FILLER_0_11_142/a_484_472# vss 0.345058f
C1524 sarlogic_0/FILLER_0_11_142/a_36_472# vss 0.404746f
C1525 sarlogic_0/FILLER_0_11_142/a_572_375# vss 0.232991f
C1526 sarlogic_0/FILLER_0_11_142/a_124_375# vss 0.185089f
C1527 sarlogic_0/net25 vss 1.803472f
C1528 sarlogic_0/_232_/a_67_603# vss 0.345683f
C1529 sarlogic_0/net35 vss 1.844415f
C1530 sarlogic_0/mask\[8\] vss 1.276233f
C1531 sarlogic_0/_301_/a_36_472# vss 0.031137f
C1532 sarlogic_0/_033_ vss 0.323682f
C1533 sarlogic_0/_165_ vss 0.331995f
C1534 sarlogic_0/FILLER_0_3_2/a_36_472# vss 0.417394f
C1535 sarlogic_0/FILLER_0_3_2/a_124_375# vss 0.246306f
C1536 sarlogic_0/trim_val\[3\] vss 0.719615f
C1537 sarlogic_0/_036_ vss 0.369206f
C1538 sarlogic_0/net68 vss 1.735004f
C1539 sarlogic_0/_447_/a_2560_156# vss 0.016968f
C1540 sarlogic_0/_447_/a_2665_112# vss 0.62251f
C1541 sarlogic_0/_447_/a_2248_156# vss 0.371662f
C1542 sarlogic_0/_447_/a_1204_472# vss 0.012971f
C1543 sarlogic_0/_447_/a_1000_472# vss 0.291735f
C1544 sarlogic_0/_447_/a_796_472# vss 0.023206f
C1545 sarlogic_0/_447_/a_1308_423# vss 0.279043f
C1546 sarlogic_0/_447_/a_448_472# vss 0.684413f
C1547 sarlogic_0/_447_/a_36_151# vss 1.43589f
C1548 sarlogic_0/FILLER_0_19_28/a_484_472# vss 0.345058f
C1549 sarlogic_0/FILLER_0_19_28/a_36_472# vss 0.404746f
C1550 sarlogic_0/FILLER_0_19_28/a_572_375# vss 0.232991f
C1551 sarlogic_0/FILLER_0_19_28/a_124_375# vss 0.185089f
C1552 sarlogic_0/fanout65/a_36_113# vss 0.418095f
C1553 sarlogic_0/fanout76/a_36_160# vss 0.386641f
C1554 sarlogic_0/net54 vss 5.456963f
C1555 sarlogic_0/fanout54/a_36_160# vss 0.696445f
C1556 sarlogic_0/FILLER_0_4_49/a_484_472# vss 0.345058f
C1557 sarlogic_0/FILLER_0_4_49/a_36_472# vss 0.404746f
C1558 sarlogic_0/FILLER_0_4_49/a_572_375# vss 0.232991f
C1559 sarlogic_0/FILLER_0_4_49/a_124_375# vss 0.185089f
C1560 sarlogic_0/_176_ vss 0.804011f
C1561 sarlogic_0/_085_ vss 2.280803f
C1562 sarlogic_0/_116_ vss 1.959915f
C1563 sarlogic_0/_395_/a_36_488# vss 0.101145f
C1564 sarlogic_0/FILLER_0_14_50/a_36_472# vss 0.417394f
C1565 sarlogic_0/FILLER_0_14_50/a_124_375# vss 0.246306f
C1566 sarlogic_0/FILLER_0_8_263/a_36_472# vss 0.417394f
C1567 sarlogic_0/FILLER_0_8_263/a_124_375# vss 0.246306f
C1568 sarlogic_0/FILLER_0_0_130/a_36_472# vss 0.417394f
C1569 sarlogic_0/FILLER_0_0_130/a_124_375# vss 0.246306f
C1570 sarlogic_0/FILLER_0_16_255/a_36_472# vss 0.417394f
C1571 sarlogic_0/FILLER_0_16_255/a_124_375# vss 0.246306f
C1572 sarlogic_0/FILLER_0_7_59/a_484_472# vss 0.345058f
C1573 sarlogic_0/FILLER_0_7_59/a_36_472# vss 0.404746f
C1574 sarlogic_0/FILLER_0_7_59/a_572_375# vss 0.232991f
C1575 sarlogic_0/FILLER_0_7_59/a_124_375# vss 0.185089f
C1576 sarlogic_0/output19/a_224_472# vss 2.38465f
C1577 sarlogic_0/FILLER_0_7_146/a_36_472# vss 0.417394f
C1578 sarlogic_0/FILLER_0_7_146/a_124_375# vss 0.246306f
C1579 sarlogic_0/_216_/a_67_603# vss 0.345683f
C1580 sarlogic_0/FILLER_0_15_116/a_484_472# vss 0.345058f
C1581 sarlogic_0/FILLER_0_15_116/a_36_472# vss 0.404746f
C1582 sarlogic_0/FILLER_0_15_116/a_572_375# vss 0.232991f
C1583 sarlogic_0/FILLER_0_15_116/a_124_375# vss 0.185089f
C1584 sarlogic_0/_063_ vss 0.370155f
C1585 sarlogic_0/_233_/a_36_160# vss 0.386641f
C1586 sarlogic_0/FILLER_0_21_28/a_3172_472# vss 0.345058f
C1587 sarlogic_0/FILLER_0_21_28/a_2724_472# vss 0.33241f
C1588 sarlogic_0/FILLER_0_21_28/a_2276_472# vss 0.33241f
C1589 sarlogic_0/FILLER_0_21_28/a_1828_472# vss 0.33241f
C1590 sarlogic_0/FILLER_0_21_28/a_1380_472# vss 0.33241f
C1591 sarlogic_0/FILLER_0_21_28/a_932_472# vss 0.33241f
C1592 sarlogic_0/FILLER_0_21_28/a_484_472# vss 0.33241f
C1593 sarlogic_0/FILLER_0_21_28/a_36_472# vss 0.404746f
C1594 sarlogic_0/FILLER_0_21_28/a_3260_375# vss 0.233093f
C1595 sarlogic_0/FILLER_0_21_28/a_2812_375# vss 0.17167f
C1596 sarlogic_0/FILLER_0_21_28/a_2364_375# vss 0.17167f
C1597 sarlogic_0/FILLER_0_21_28/a_1916_375# vss 0.17167f
C1598 sarlogic_0/FILLER_0_21_28/a_1468_375# vss 0.17167f
C1599 sarlogic_0/FILLER_0_21_28/a_1020_375# vss 0.17167f
C1600 sarlogic_0/FILLER_0_21_28/a_572_375# vss 0.17167f
C1601 sarlogic_0/FILLER_0_21_28/a_124_375# vss 0.185915f
C1602 sarlogic_0/_110_ vss 0.323912f
C1603 sarlogic_0/_379_/a_36_472# vss 0.031137f
C1604 sarlogic_0/trim_val\[4\] vss 0.662409f
C1605 sarlogic_0/net76 vss 1.454269f
C1606 sarlogic_0/_448_/a_2560_156# vss 0.016968f
C1607 sarlogic_0/_448_/a_2665_112# vss 0.62251f
C1608 sarlogic_0/_448_/a_2248_156# vss 0.371662f
C1609 sarlogic_0/_448_/a_1204_472# vss 0.012971f
C1610 sarlogic_0/_448_/a_1000_472# vss 0.291735f
C1611 sarlogic_0/_448_/a_796_472# vss 0.023206f
C1612 sarlogic_0/_448_/a_1308_423# vss 0.279043f
C1613 sarlogic_0/_448_/a_448_472# vss 0.684413f
C1614 sarlogic_0/_448_/a_36_151# vss 1.43589f
C1615 sarlogic_0/fanout64/a_36_160# vss 0.386641f
C1616 sarlogic_0/fanout75/a_36_113# vss 0.418095f
C1617 sarlogic_0/_250_/a_36_68# vss 0.69549f
C1618 sarlogic_0/net56 vss 0.843396f
C1619 sarlogic_0/fanout53/a_36_160# vss 0.696445f
C1620 sarlogic_0/_177_ vss 0.358286f
C1621 result[2] vss 24.971811f
C1622 sarlogic_0/net29 vss 1.802718f
C1623 sarlogic_0/output29/a_224_472# vss 2.38465f
C1624 sarlogic_0/output18/a_224_472# vss 2.38465f
C1625 sarlogic_0/FILLER_0_14_181/a_36_472# vss 0.417394f
C1626 sarlogic_0/FILLER_0_14_181/a_124_375# vss 0.246306f
C1627 sarlogic_0/_052_ vss 0.569133f
C1628 sarlogic_0/_217_/a_36_160# vss 0.386641f
C1629 sarlogic_0/net44 vss 1.407054f
C1630 sarlogic_0/_303_/a_36_472# vss 0.031137f
C1631 sarlogic_0/en_co_clk vss 0.346872f
C1632 sarlogic_0/net55 vss 5.119958f
C1633 sarlogic_0/net72 vss 1.366255f
C1634 sarlogic_0/_449_/a_2560_156# vss 0.016968f
C1635 sarlogic_0/_449_/a_2665_112# vss 0.62251f
C1636 sarlogic_0/_449_/a_2248_156# vss 0.371662f
C1637 sarlogic_0/_449_/a_1204_472# vss 0.012971f
C1638 sarlogic_0/_449_/a_1000_472# vss 0.291735f
C1639 sarlogic_0/_449_/a_796_472# vss 0.023206f
C1640 sarlogic_0/_449_/a_1308_423# vss 0.279043f
C1641 sarlogic_0/_449_/a_448_472# vss 0.684413f
C1642 sarlogic_0/_449_/a_36_151# vss 1.43589f
C1643 sarlogic_0/fanout52/a_36_160# vss 0.696445f
C1644 sarlogic_0/net82 vss 0.706042f
C1645 sarlogic_0/fanout74/a_36_113# vss 0.418095f
C1646 sarlogic_0/FILLER_0_10_28/a_36_472# vss 0.417394f
C1647 sarlogic_0/FILLER_0_10_28/a_124_375# vss 0.246306f
C1648 sarlogic_0/mask\[0\] vss 2.242948f
C1649 sarlogic_0/_320_/a_36_472# vss 0.137725f
C1650 sarlogic_0/fanout63/a_36_160# vss 0.696445f
C1651 sarlogic_0/FILLER_0_14_81/a_36_472# vss 0.417394f
C1652 sarlogic_0/FILLER_0_14_81/a_124_375# vss 0.246306f
C1653 sarlogic_0/_397_/a_36_472# vss 0.031137f
C1654 sarlogic_0/FILLER_0_13_212/a_1380_472# vss 0.345058f
C1655 sarlogic_0/FILLER_0_13_212/a_932_472# vss 0.33241f
C1656 sarlogic_0/FILLER_0_13_212/a_484_472# vss 0.33241f
C1657 sarlogic_0/FILLER_0_13_212/a_36_472# vss 0.404746f
C1658 sarlogic_0/FILLER_0_13_212/a_1468_375# vss 0.233029f
C1659 sarlogic_0/FILLER_0_13_212/a_1020_375# vss 0.171606f
C1660 sarlogic_0/FILLER_0_13_212/a_572_375# vss 0.171606f
C1661 sarlogic_0/FILLER_0_13_212/a_124_375# vss 0.185399f
C1662 sarlogic_0/net39 vss 1.445128f
C1663 sarlogic_0/output39/a_224_472# vss 2.38465f
C1664 result[1] vss 24.970469f
C1665 sarlogic_0/net28 vss 1.759728f
C1666 sarlogic_0/output28/a_224_472# vss 2.38465f
C1667 sarlogic_0/output17/a_224_472# vss 2.38465f
C1668 sarlogic_0/FILLER_0_16_37/a_36_472# vss 0.417394f
C1669 sarlogic_0/FILLER_0_16_37/a_124_375# vss 0.246306f
C1670 sarlogic_0/net26 vss 1.671545f
C1671 sarlogic_0/_064_ vss 0.581481f
C1672 sarlogic_0/trim_val\[2\] vss 0.65354f
C1673 sarlogic_0/trim_mask\[2\] vss 0.92551f
C1674 sarlogic_0/_235_/a_67_603# vss 0.345683f
C1675 sarlogic_0/_013_ vss 0.48783f
C1676 sarlogic_0/_111_ vss 0.369652f
C1677 sarlogic_0/FILLER_0_18_177/a_3172_472# vss 0.345058f
C1678 sarlogic_0/FILLER_0_18_177/a_2724_472# vss 0.33241f
C1679 sarlogic_0/FILLER_0_18_177/a_2276_472# vss 0.33241f
C1680 sarlogic_0/FILLER_0_18_177/a_1828_472# vss 0.33241f
C1681 sarlogic_0/FILLER_0_18_177/a_1380_472# vss 0.33241f
C1682 sarlogic_0/FILLER_0_18_177/a_932_472# vss 0.33241f
C1683 sarlogic_0/FILLER_0_18_177/a_484_472# vss 0.33241f
C1684 sarlogic_0/FILLER_0_18_177/a_36_472# vss 0.404746f
C1685 sarlogic_0/FILLER_0_18_177/a_3260_375# vss 0.233093f
C1686 sarlogic_0/FILLER_0_18_177/a_2812_375# vss 0.17167f
C1687 sarlogic_0/FILLER_0_18_177/a_2364_375# vss 0.17167f
C1688 sarlogic_0/FILLER_0_18_177/a_1916_375# vss 0.17167f
C1689 sarlogic_0/FILLER_0_18_177/a_1468_375# vss 0.17167f
C1690 sarlogic_0/FILLER_0_18_177/a_1020_375# vss 0.17167f
C1691 sarlogic_0/FILLER_0_18_177/a_572_375# vss 0.17167f
C1692 sarlogic_0/FILLER_0_18_177/a_124_375# vss 0.185915f
C1693 sarlogic_0/FILLER_0_18_100/a_36_472# vss 0.417394f
C1694 sarlogic_0/FILLER_0_18_100/a_124_375# vss 0.246306f
C1695 sarlogic_0/_073_ vss 0.953711f
C1696 sarlogic_0/_126_ vss 2.036767f
C1697 sarlogic_0/_069_ vss 2.034557f
C1698 sarlogic_0/_321_/a_170_472# vss 0.077257f
C1699 sarlogic_0/fanout51/a_36_113# vss 0.418095f
C1700 sarlogic_0/net62 vss 4.932099f
C1701 sarlogic_0/fanout62/a_36_160# vss 0.696445f
C1702 sarlogic_0/fanout73/a_36_113# vss 0.418095f
C1703 sarlogic_0/FILLER_0_19_47/a_484_472# vss 0.345058f
C1704 sarlogic_0/FILLER_0_19_47/a_36_472# vss 0.404746f
C1705 sarlogic_0/FILLER_0_19_47/a_572_375# vss 0.232991f
C1706 sarlogic_0/FILLER_0_19_47/a_124_375# vss 0.185089f
C1707 sarlogic_0/FILLER_0_14_91/a_484_472# vss 0.345058f
C1708 sarlogic_0/FILLER_0_14_91/a_36_472# vss 0.404746f
C1709 sarlogic_0/FILLER_0_14_91/a_572_375# vss 0.232991f
C1710 sarlogic_0/FILLER_0_14_91/a_124_375# vss 0.185089f
C1711 sarlogic_0/FILLER_0_10_214/a_36_472# vss 0.417394f
C1712 sarlogic_0/FILLER_0_10_214/a_124_375# vss 0.246306f
C1713 sarlogic_0/FILLER_0_10_247/a_36_472# vss 0.417394f
C1714 sarlogic_0/FILLER_0_10_247/a_124_375# vss 0.246306f
C1715 sarlogic_0/_178_ vss 1.252435f
C1716 sarlogic_0/_398_/a_36_113# vss 0.418095f
C1717 sarlogic_0/FILLER_0_16_241/a_36_472# vss 0.417394f
C1718 sarlogic_0/FILLER_0_16_241/a_124_375# vss 0.246306f
C1719 sarlogic_0/net38 vss 1.529392f
C1720 sarlogic_0/output38/a_224_472# vss 2.38465f
C1721 sarlogic_0/net16 vss 1.295744f
C1722 sarlogic_0/output16/a_224_472# vss 2.38465f
C1723 result[0] vss 29.692343f
C1724 sarlogic_0/output27/a_224_472# vss 2.38465f
C1725 sarlogic_0/_219_/a_36_160# vss 0.386641f
C1726 sarlogic_0/FILLER_0_20_193/a_484_472# vss 0.345058f
C1727 sarlogic_0/FILLER_0_20_193/a_36_472# vss 0.404746f
C1728 sarlogic_0/FILLER_0_20_193/a_572_375# vss 0.232991f
C1729 sarlogic_0/FILLER_0_20_193/a_124_375# vss 0.185089f
C1730 sarlogic_0/_236_/a_36_160# vss 0.696445f
C1731 sarlogic_0/_112_ vss 0.308886f
C1732 sarlogic_0/_305_/a_36_159# vss 0.374116f
C1733 sarlogic_0/_074_ vss 1.813232f
C1734 sarlogic_0/_253_/a_36_68# vss 0.061249f
C1735 sarlogic_0/net50 vss 4.486121f
C1736 sarlogic_0/net52 vss 3.536016f
C1737 sarlogic_0/fanout50/a_36_160# vss 0.696445f
C1738 sarlogic_0/FILLER_0_10_37/a_36_472# vss 0.417394f
C1739 sarlogic_0/FILLER_0_10_37/a_124_375# vss 0.246306f
C1740 sarlogic_0/fanout72/a_36_113# vss 0.418095f
C1741 sarlogic_0/fanout61/a_36_113# vss 0.418095f
C1742 sarlogic_0/_128_ vss 0.447252f
C1743 sarlogic_0/_127_ vss 1.291729f
C1744 sarlogic_0/_322_/a_848_380# vss 0.40208f
C1745 sarlogic_0/_322_/a_124_24# vss 0.591898f
C1746 sarlogic_0/_088_ vss 0.457961f
C1747 sarlogic_0/_079_ vss 1.114894f
C1748 sarlogic_0/_087_ vss 0.601674f
C1749 sarlogic_0/_270_/a_36_472# vss 0.031137f
C1750 sarlogic_0/FILLER_0_4_123/a_36_472# vss 0.417394f
C1751 sarlogic_0/FILLER_0_4_123/a_124_375# vss 0.246306f
C1752 sarlogic_0/FILLER_0_17_218/a_484_472# vss 0.345058f
C1753 sarlogic_0/FILLER_0_17_218/a_36_472# vss 0.404746f
C1754 sarlogic_0/FILLER_0_17_218/a_572_375# vss 0.232991f
C1755 sarlogic_0/FILLER_0_17_218/a_124_375# vss 0.185089f
C1756 sarlogic_0/output37/a_224_472# vss 2.38465f
C1757 valid vss 29.398195f
C1758 sarlogic_0/net48 vss 1.219262f
C1759 sarlogic_0/output48/a_224_472# vss 2.38465f
C1760 sarlogic_0/net15 vss 1.447491f
C1761 sarlogic_0/output15/a_224_472# vss 2.38465f
C1762 sarlogic_0/output26/a_224_472# vss 2.38465f
C1763 sarlogic_0/FILLER_0_16_57/a_1380_472# vss 0.345058f
C1764 sarlogic_0/FILLER_0_16_57/a_932_472# vss 0.33241f
C1765 sarlogic_0/FILLER_0_16_57/a_484_472# vss 0.33241f
C1766 sarlogic_0/FILLER_0_16_57/a_36_472# vss 0.404746f
C1767 sarlogic_0/FILLER_0_16_57/a_1468_375# vss 0.233029f
C1768 sarlogic_0/FILLER_0_16_57/a_1020_375# vss 0.171606f
C1769 sarlogic_0/FILLER_0_16_57/a_572_375# vss 0.171606f
C1770 sarlogic_0/FILLER_0_16_57/a_124_375# vss 0.185399f
C1771 sarlogic_0/_306_/a_36_68# vss 0.69549f
C1772 sarlogic_0/_072_ vss 2.604301f
C1773 sarlogic_0/fanout82/a_36_113# vss 0.418095f
C1774 sarlogic_0/_015_ vss 0.406653f
C1775 sarlogic_0/_323_/a_36_113# vss 0.418095f
C1776 sarlogic_0/net60 vss 5.024503f
C1777 sarlogic_0/net61 vss 1.666523f
C1778 sarlogic_0/fanout60/a_36_160# vss 0.696445f
C1779 sarlogic_0/fanout71/a_36_113# vss 0.418095f
C1780 sarlogic_0/FILLER_0_6_239/a_36_472# vss 0.417394f
C1781 sarlogic_0/FILLER_0_6_239/a_124_375# vss 0.246306f
C1782 sarlogic_0/FILLER_0_4_99/a_36_472# vss 0.417394f
C1783 sarlogic_0/FILLER_0_4_99/a_124_375# vss 0.246306f
C1784 sarlogic_0/net57 vss 1.383718f
C1785 sarlogic_0/FILLER_0_10_256/a_36_472# vss 0.417394f
C1786 sarlogic_0/FILLER_0_10_256/a_124_375# vss 0.246306f
C1787 sarlogic_0/cal_itt\[3\] vss 1.854962f
C1788 sarlogic_0/_340_/a_36_160# vss 0.386641f
C1789 sarlogic_0/FILLER_0_4_177/a_484_472# vss 0.345058f
C1790 sarlogic_0/FILLER_0_4_177/a_36_472# vss 0.404746f
C1791 sarlogic_0/FILLER_0_4_177/a_572_375# vss 0.232991f
C1792 sarlogic_0/FILLER_0_4_177/a_124_375# vss 0.185089f
C1793 sarlogic_0/FILLER_0_4_144/a_484_472# vss 0.345058f
C1794 sarlogic_0/FILLER_0_4_144/a_36_472# vss 0.404746f
C1795 sarlogic_0/FILLER_0_4_144/a_572_375# vss 0.232991f
C1796 sarlogic_0/FILLER_0_4_144/a_124_375# vss 0.185089f
C1797 sarlogic_0/output14/a_224_472# vss 2.38465f
C1798 result[9] vss 30.117216f
C1799 sarlogic_0/output36/a_224_472# vss 2.38465f
C1800 sarlogic_0/output47/a_224_472# vss 2.38465f
C1801 sarlogic_0/output25/a_224_472# vss 2.389677f
C1802 sarlogic_0/FILLER_0_12_136/a_1380_472# vss 0.345058f
C1803 sarlogic_0/FILLER_0_12_136/a_932_472# vss 0.33241f
C1804 sarlogic_0/FILLER_0_12_136/a_484_472# vss 0.33241f
C1805 sarlogic_0/FILLER_0_12_136/a_36_472# vss 0.404746f
C1806 sarlogic_0/FILLER_0_12_136/a_1468_375# vss 0.233029f
C1807 sarlogic_0/FILLER_0_12_136/a_1020_375# vss 0.171606f
C1808 sarlogic_0/FILLER_0_12_136/a_572_375# vss 0.171606f
C1809 sarlogic_0/FILLER_0_12_136/a_124_375# vss 0.185399f
C1810 sarlogic_0/FILLER_0_16_89/a_1380_472# vss 0.345058f
C1811 sarlogic_0/FILLER_0_16_89/a_932_472# vss 0.33241f
C1812 sarlogic_0/FILLER_0_16_89/a_484_472# vss 0.33241f
C1813 sarlogic_0/FILLER_0_16_89/a_36_472# vss 0.404746f
C1814 sarlogic_0/FILLER_0_16_89/a_1468_375# vss 0.233029f
C1815 sarlogic_0/FILLER_0_16_89/a_1020_375# vss 0.171606f
C1816 sarlogic_0/FILLER_0_16_89/a_572_375# vss 0.171606f
C1817 sarlogic_0/FILLER_0_16_89/a_124_375# vss 0.185399f
C1818 sarlogic_0/FILLER_0_21_125/a_484_472# vss 0.345058f
C1819 sarlogic_0/FILLER_0_21_125/a_36_472# vss 0.404746f
C1820 sarlogic_0/FILLER_0_21_125/a_572_375# vss 0.232991f
C1821 sarlogic_0/FILLER_0_21_125/a_124_375# vss 0.185089f
C1822 sarlogic_0/_238_/a_67_603# vss 0.345683f
C1823 sarlogic_0/_096_ vss 2.205532f
C1824 sarlogic_0/_093_ vss 1.893313f
C1825 sarlogic_0/FILLER_0_19_55/a_36_472# vss 0.417394f
C1826 sarlogic_0/FILLER_0_19_55/a_124_375# vss 0.246306f
C1827 sarlogic_0/net81 vss 1.738987f
C1828 sarlogic_0/fanout81/a_36_160# vss 0.386641f
C1829 sarlogic_0/_057_ vss 1.600886f
C1830 sarlogic_0/_255_/a_224_552# vss 1.31114f
C1831 sarlogic_0/net73 vss 1.058857f
C1832 sarlogic_0/fanout70/a_36_113# vss 0.418095f
C1833 sarlogic_0/_003_ vss 0.3064f
C1834 sarlogic_0/_089_ vss 0.36777f
C1835 sarlogic_0/_272_/a_36_472# vss 0.031137f
C1836 sarlogic_0/_187_ vss 0.311229f
C1837 sarlogic_0/_410_/a_36_68# vss 0.112263f
C1838 sarlogic_0/_141_ vss 1.249289f
C1839 sarlogic_0/mask\[3\] vss 1.26722f
C1840 sarlogic_0/_341_/a_49_472# vss 0.054843f
C1841 cal vss 25.534355f
C1842 sarlogic_0/FILLER_0_7_195/a_36_472# vss 0.417394f
C1843 sarlogic_0/FILLER_0_7_195/a_124_375# vss 0.246306f
C1844 sarlogic_0/FILLER_0_7_162/a_36_472# vss 0.417394f
C1845 sarlogic_0/FILLER_0_7_162/a_124_375# vss 0.246306f
C1846 sarlogic_0/output13/a_224_472# vss 2.391402f
C1847 sarlogic_0/FILLER_0_18_2/a_3172_472# vss 0.345058f
C1848 sarlogic_0/FILLER_0_18_2/a_2724_472# vss 0.33241f
C1849 sarlogic_0/FILLER_0_18_2/a_2276_472# vss 0.33241f
C1850 sarlogic_0/FILLER_0_18_2/a_1828_472# vss 0.33241f
C1851 sarlogic_0/FILLER_0_18_2/a_1380_472# vss 0.33241f
C1852 sarlogic_0/FILLER_0_18_2/a_932_472# vss 0.33241f
C1853 sarlogic_0/FILLER_0_18_2/a_484_472# vss 0.33241f
C1854 sarlogic_0/FILLER_0_18_2/a_36_472# vss 0.404746f
C1855 sarlogic_0/FILLER_0_18_2/a_3260_375# vss 0.233093f
C1856 sarlogic_0/FILLER_0_18_2/a_2812_375# vss 0.17167f
C1857 sarlogic_0/FILLER_0_18_2/a_2364_375# vss 0.17167f
C1858 sarlogic_0/FILLER_0_18_2/a_1916_375# vss 0.17167f
C1859 sarlogic_0/FILLER_0_18_2/a_1468_375# vss 0.17167f
C1860 sarlogic_0/FILLER_0_18_2/a_1020_375# vss 0.17167f
C1861 sarlogic_0/FILLER_0_18_2/a_572_375# vss 0.17167f
C1862 sarlogic_0/FILLER_0_18_2/a_124_375# vss 0.185915f
C1863 sarlogic_0/net46 vss 1.13395f
C1864 sarlogic_0/output46/a_224_472# vss 2.38465f
C1865 result[8] vss 25.736643f
C1866 sarlogic_0/output35/a_224_472# vss 2.38465f
C1867 sarlogic_0/output24/a_224_472# vss 2.38465f
C1868 sarlogic_0/FILLER_0_8_107/a_36_472# vss 0.417394f
C1869 sarlogic_0/FILLER_0_8_107/a_124_375# vss 0.246306f
C1870 sarlogic_0/FILLER_0_12_124/a_36_472# vss 0.417394f
C1871 sarlogic_0/FILLER_0_12_124/a_124_375# vss 0.246306f
C1872 sarlogic_0/net41 vss 1.746759f
C1873 sarlogic_0/_065_ vss 0.523724f
C1874 sarlogic_0/_239_/a_36_160# vss 0.696445f
C1875 sarlogic_0/FILLER_0_1_98/a_36_472# vss 0.417394f
C1876 sarlogic_0/FILLER_0_1_98/a_124_375# vss 0.246306f
C1877 sarlogic_0/_115_ vss 1.281516f
C1878 sarlogic_0/_114_ vss 2.293579f
C1879 sarlogic_0/_308_/a_848_380# vss 0.40208f
C1880 sarlogic_0/_308_/a_124_24# vss 0.591898f
C1881 sarlogic_0/_256_/a_36_68# vss 0.063181f
C1882 sarlogic_0/FILLER_0_10_78/a_1380_472# vss 0.345058f
C1883 sarlogic_0/FILLER_0_10_78/a_932_472# vss 0.33241f
C1884 sarlogic_0/FILLER_0_10_78/a_484_472# vss 0.33241f
C1885 sarlogic_0/FILLER_0_10_78/a_36_472# vss 0.404746f
C1886 sarlogic_0/FILLER_0_10_78/a_1468_375# vss 0.233029f
C1887 sarlogic_0/FILLER_0_10_78/a_1020_375# vss 0.171606f
C1888 sarlogic_0/FILLER_0_10_78/a_572_375# vss 0.171606f
C1889 sarlogic_0/FILLER_0_10_78/a_124_375# vss 0.185399f
C1890 sarlogic_0/_130_ vss 0.304085f
C1891 sarlogic_0/net80 vss 1.375599f
C1892 sarlogic_0/fanout80/a_36_113# vss 0.418095f
C1893 sarlogic_0/net58 vss 5.308423f
C1894 sarlogic_0/_000_ vss 0.382358f
C1895 sarlogic_0/net75 vss 1.474299f
C1896 sarlogic_0/_411_/a_2560_156# vss 0.016968f
C1897 sarlogic_0/_411_/a_2665_112# vss 0.62251f
C1898 sarlogic_0/_411_/a_2248_156# vss 0.371662f
C1899 sarlogic_0/_411_/a_1204_472# vss 0.012971f
C1900 sarlogic_0/_411_/a_1000_472# vss 0.291735f
C1901 sarlogic_0/_411_/a_796_472# vss 0.023206f
C1902 sarlogic_0/_411_/a_1308_423# vss 0.279043f
C1903 sarlogic_0/_411_/a_448_472# vss 0.684413f
C1904 sarlogic_0/_411_/a_36_151# vss 1.43589f
C1905 sarlogic_0/state\[0\] vss 0.680109f
C1906 sarlogic_0/_273_/a_36_68# vss 0.69549f
C1907 sarlogic_0/_142_ vss 0.324372f
C1908 sarlogic_0/FILLER_0_9_223/a_484_472# vss 0.345058f
C1909 sarlogic_0/FILLER_0_9_223/a_36_472# vss 0.404746f
C1910 sarlogic_0/FILLER_0_9_223/a_572_375# vss 0.232991f
C1911 sarlogic_0/FILLER_0_9_223/a_124_375# vss 0.185089f
C1912 sarlogic_0/FILLER_0_4_197/a_1380_472# vss 0.345058f
C1913 sarlogic_0/FILLER_0_4_197/a_932_472# vss 0.33241f
C1914 sarlogic_0/FILLER_0_4_197/a_484_472# vss 0.33241f
C1915 sarlogic_0/FILLER_0_4_197/a_36_472# vss 0.404746f
C1916 sarlogic_0/FILLER_0_4_197/a_1468_375# vss 0.233029f
C1917 sarlogic_0/FILLER_0_4_197/a_1020_375# vss 0.171606f
C1918 sarlogic_0/FILLER_0_4_197/a_572_375# vss 0.171606f
C1919 sarlogic_0/FILLER_0_4_197/a_124_375# vss 0.185399f
C1920 sarlogic_0/FILLER_0_17_226/a_36_472# vss 0.417394f
C1921 sarlogic_0/FILLER_0_17_226/a_124_375# vss 0.246306f
C1922 sarlogic_0/FILLER_0_5_109/a_484_472# vss 0.345058f
C1923 sarlogic_0/FILLER_0_5_109/a_36_472# vss 0.404746f
C1924 sarlogic_0/FILLER_0_5_109/a_572_375# vss 0.232991f
C1925 sarlogic_0/FILLER_0_5_109/a_124_375# vss 0.185089f
C1926 sarlogic_0/output12/a_224_472# vss 2.38465f
C1927 result[7] vss 24.988647f
C1928 sarlogic_0/net34 vss 1.724665f
C1929 sarlogic_0/output34/a_224_472# vss 2.38465f
C1930 sarlogic_0/net45 vss 1.12041f
C1931 sarlogic_0/output45/a_224_472# vss 2.38465f
C1932 sarlogic_0/output23/a_224_472# vss 2.390503f
C1933 sarlogic_0/FILLER_0_15_142/a_484_472# vss 0.345058f
C1934 sarlogic_0/FILLER_0_15_142/a_36_472# vss 0.404746f
C1935 sarlogic_0/FILLER_0_15_142/a_572_375# vss 0.232991f
C1936 sarlogic_0/FILLER_0_15_142/a_124_375# vss 0.185089f
C1937 sarlogic_0/_077_ vss 1.645892f
C1938 sarlogic_0/_075_ vss 0.374516f
C1939 sarlogic_0/_257_/a_36_472# vss 0.031137f
C1940 sarlogic_0/_326_/a_36_160# vss 0.696445f
C1941 sarlogic_0/_412_/a_2560_156# vss 0.016968f
C1942 sarlogic_0/_412_/a_2665_112# vss 0.62251f
C1943 sarlogic_0/_412_/a_2248_156# vss 0.371662f
C1944 sarlogic_0/_412_/a_1204_472# vss 0.012971f
C1945 sarlogic_0/_412_/a_1000_472# vss 0.291735f
C1946 sarlogic_0/_412_/a_796_472# vss 0.023206f
C1947 sarlogic_0/_412_/a_1308_423# vss 0.279043f
C1948 sarlogic_0/_412_/a_448_472# vss 0.684413f
C1949 sarlogic_0/_412_/a_36_151# vss 1.43589f
C1950 sarlogic_0/_091_ vss 1.841339f
C1951 sarlogic_0/_274_/a_36_68# vss 0.063181f
C1952 sarlogic_0/_143_ vss 0.329289f
C1953 sarlogic_0/mask\[4\] vss 1.300438f
C1954 sarlogic_0/_343_/a_49_472# vss 0.054843f
C1955 sarlogic_0/FILLER_0_13_65/a_36_472# vss 0.417394f
C1956 sarlogic_0/FILLER_0_13_65/a_124_375# vss 0.246306f
C1957 sarlogic_0/_360_/a_36_160# vss 0.386641f
C1958 sarlogic_0/FILLER_0_4_185/a_36_472# vss 0.417394f
C1959 sarlogic_0/FILLER_0_4_185/a_124_375# vss 0.246306f
C1960 sarlogic_0/FILLER_0_4_152/a_36_472# vss 0.417394f
C1961 sarlogic_0/FILLER_0_4_152/a_124_375# vss 0.246306f
C1962 sarlogic_0/_291_/a_36_160# vss 0.386641f
C1963 sarlogic_0/output9/a_224_472# vss 2.38465f
C1964 sarlogic_0/output11/a_224_472# vss 2.391497f
C1965 sarlogic_0/output44/a_224_472# vss 2.38465f
C1966 result[6] vss 24.936083f
C1967 sarlogic_0/output33/a_224_472# vss 2.38465f
C1968 sarlogic_0/output22/a_224_472# vss 2.38465f
C1969 sarlogic_0/FILLER_0_8_127/a_36_472# vss 0.417394f
C1970 sarlogic_0/FILLER_0_8_127/a_124_375# vss 0.246306f
C1971 sarlogic_0/FILLER_0_8_138/a_36_472# vss 0.417394f
C1972 sarlogic_0/FILLER_0_8_138/a_124_375# vss 0.246306f
C1973 sarlogic_0/FILLER_0_21_133/a_36_472# vss 0.417394f
C1974 sarlogic_0/FILLER_0_21_133/a_124_375# vss 0.246306f
C1975 sarlogic_0/FILLER_0_24_130/a_36_472# vss 0.417394f
C1976 sarlogic_0/FILLER_0_24_130/a_124_375# vss 0.246306f
C1977 sarlogic_0/FILLER_0_18_171/a_36_472# vss 0.417394f
C1978 sarlogic_0/FILLER_0_18_171/a_124_375# vss 0.246306f
C1979 sarlogic_0/_258_/a_36_160# vss 0.386641f
C1980 sarlogic_0/_016_ vss 0.314121f
C1981 sarlogic_0/_327_/a_36_472# vss 0.031137f
C1982 sarlogic_0/_189_/a_67_603# vss 0.345683f
C1983 sarlogic_0/FILLER_0_24_63/a_36_472# vss 0.417394f
C1984 sarlogic_0/FILLER_0_24_63/a_124_375# vss 0.246306f
C1985 sarlogic_0/FILLER_0_24_96/a_36_472# vss 0.417394f
C1986 sarlogic_0/FILLER_0_24_96/a_124_375# vss 0.246306f
C1987 sarlogic_0/cal_itt\[2\] vss 1.473514f
C1988 sarlogic_0/_002_ vss 0.289553f
C1989 sarlogic_0/_413_/a_2560_156# vss 0.016968f
C1990 sarlogic_0/_413_/a_2665_112# vss 0.62251f
C1991 sarlogic_0/_413_/a_2248_156# vss 0.371662f
C1992 sarlogic_0/_413_/a_1204_472# vss 0.012971f
C1993 sarlogic_0/_413_/a_1000_472# vss 0.291735f
C1994 sarlogic_0/_413_/a_796_472# vss 0.023206f
C1995 sarlogic_0/_413_/a_1308_423# vss 0.279043f
C1996 sarlogic_0/_413_/a_448_472# vss 0.684413f
C1997 sarlogic_0/_413_/a_36_151# vss 1.43589f
C1998 sarlogic_0/_092_ vss 0.680239f
C1999 sarlogic_0/FILLER_0_7_72/a_3172_472# vss 0.345058f
C2000 sarlogic_0/FILLER_0_7_72/a_2724_472# vss 0.33241f
C2001 sarlogic_0/FILLER_0_7_72/a_2276_472# vss 0.33241f
C2002 sarlogic_0/FILLER_0_7_72/a_1828_472# vss 0.33241f
C2003 sarlogic_0/FILLER_0_7_72/a_1380_472# vss 0.33241f
C2004 sarlogic_0/FILLER_0_7_72/a_932_472# vss 0.33241f
C2005 sarlogic_0/FILLER_0_7_72/a_484_472# vss 0.33241f
C2006 sarlogic_0/FILLER_0_7_72/a_36_472# vss 0.404746f
C2007 sarlogic_0/FILLER_0_7_72/a_3260_375# vss 0.233093f
C2008 sarlogic_0/FILLER_0_7_72/a_2812_375# vss 0.17167f
C2009 sarlogic_0/FILLER_0_7_72/a_2364_375# vss 0.17167f
C2010 sarlogic_0/FILLER_0_7_72/a_1916_375# vss 0.17167f
C2011 sarlogic_0/FILLER_0_7_72/a_1468_375# vss 0.17167f
C2012 sarlogic_0/FILLER_0_7_72/a_1020_375# vss 0.17167f
C2013 sarlogic_0/FILLER_0_7_72/a_572_375# vss 0.17167f
C2014 sarlogic_0/FILLER_0_7_72/a_124_375# vss 0.185915f
C2015 sarlogic_0/_086_ vss 2.45259f
C2016 sarlogic_0/_119_ vss 1.237181f
C2017 sarlogic_0/net63 vss 5.362473f
C2018 sarlogic_0/_430_/a_2560_156# vss 0.016968f
C2019 sarlogic_0/_430_/a_2665_112# vss 0.62251f
C2020 sarlogic_0/_430_/a_2248_156# vss 0.371662f
C2021 sarlogic_0/_430_/a_1204_472# vss 0.012971f
C2022 sarlogic_0/_430_/a_1000_472# vss 0.291735f
C2023 sarlogic_0/_430_/a_796_472# vss 0.023206f
C2024 sarlogic_0/_430_/a_1308_423# vss 0.279043f
C2025 sarlogic_0/_430_/a_448_472# vss 0.684413f
C2026 sarlogic_0/_430_/a_36_151# vss 1.43589f
C2027 sarlogic_0/_292_/a_36_160# vss 0.386641f
C2028 sarlogic_0/output8/a_224_472# vss 2.38465f
C2029 sarlogic_0/output10/a_224_472# vss 2.38465f
C2030 result[5] vss 24.947828f
C2031 sarlogic_0/net32 vss 1.789002f
C2032 sarlogic_0/output32/a_224_472# vss 2.38465f
C2033 sarlogic_0/output43/a_224_472# vss 2.38465f
C2034 sarlogic_0/output21/a_224_472# vss 2.39076f
C2035 sarlogic_0/_053_ vss 1.705161f
C2036 sarlogic_0/FILLER_0_16_107/a_484_472# vss 0.345058f
C2037 sarlogic_0/FILLER_0_16_107/a_36_472# vss 0.404746f
C2038 sarlogic_0/FILLER_0_16_107/a_572_375# vss 0.232991f
C2039 sarlogic_0/FILLER_0_16_107/a_124_375# vss 0.185089f
C2040 sarlogic_0/FILLER_0_3_204/a_36_472# vss 0.417394f
C2041 sarlogic_0/FILLER_0_3_204/a_124_375# vss 0.246306f
C2042 sarlogic_0/FILLER_0_9_28/a_3172_472# vss 0.345058f
C2043 sarlogic_0/FILLER_0_9_28/a_2724_472# vss 0.33241f
C2044 sarlogic_0/FILLER_0_9_28/a_2276_472# vss 0.33241f
C2045 sarlogic_0/FILLER_0_9_28/a_1828_472# vss 0.33241f
C2046 sarlogic_0/FILLER_0_9_28/a_1380_472# vss 0.33241f
C2047 sarlogic_0/FILLER_0_9_28/a_932_472# vss 0.33241f
C2048 sarlogic_0/FILLER_0_9_28/a_484_472# vss 0.33241f
C2049 sarlogic_0/FILLER_0_9_28/a_36_472# vss 0.404746f
C2050 sarlogic_0/FILLER_0_9_28/a_3260_375# vss 0.233093f
C2051 sarlogic_0/FILLER_0_9_28/a_2812_375# vss 0.17167f
C2052 sarlogic_0/FILLER_0_9_28/a_2364_375# vss 0.17167f
C2053 sarlogic_0/FILLER_0_9_28/a_1916_375# vss 0.17167f
C2054 sarlogic_0/FILLER_0_9_28/a_1468_375# vss 0.17167f
C2055 sarlogic_0/FILLER_0_9_28/a_1020_375# vss 0.17167f
C2056 sarlogic_0/FILLER_0_9_28/a_572_375# vss 0.17167f
C2057 sarlogic_0/FILLER_0_9_28/a_124_375# vss 0.185915f
C2058 sarlogic_0/_132_ vss 1.491425f
C2059 sarlogic_0/_328_/a_36_113# vss 0.418095f
C2060 sarlogic_0/_414_/a_2560_156# vss 0.016968f
C2061 sarlogic_0/_414_/a_2665_112# vss 0.62251f
C2062 sarlogic_0/_414_/a_2248_156# vss 0.371662f
C2063 sarlogic_0/_414_/a_1204_472# vss 0.012971f
C2064 sarlogic_0/_414_/a_1000_472# vss 0.291735f
C2065 sarlogic_0/_414_/a_796_472# vss 0.023206f
C2066 sarlogic_0/_414_/a_1308_423# vss 0.279043f
C2067 sarlogic_0/_414_/a_448_472# vss 0.684413f
C2068 sarlogic_0/_414_/a_36_151# vss 1.43589f
C2069 sarlogic_0/_276_/a_36_160# vss 0.386641f
C2070 sarlogic_0/_144_ vss 1.173846f
C2071 sarlogic_0/_345_/a_36_160# vss 0.386641f
C2072 sarlogic_0/_155_ vss 0.638535f
C2073 sarlogic_0/_020_ vss 0.316793f
C2074 sarlogic_0/_431_/a_2560_156# vss 0.016968f
C2075 sarlogic_0/_431_/a_2665_112# vss 0.62251f
C2076 sarlogic_0/_431_/a_2248_156# vss 0.371662f
C2077 sarlogic_0/_431_/a_1204_472# vss 0.012971f
C2078 sarlogic_0/_431_/a_1000_472# vss 0.291735f
C2079 sarlogic_0/_431_/a_796_472# vss 0.023206f
C2080 sarlogic_0/_431_/a_1308_423# vss 0.279043f
C2081 sarlogic_0/_431_/a_448_472# vss 0.684413f
C2082 sarlogic_0/_431_/a_36_151# vss 1.43589f
C2083 sarlogic_0/_105_ vss 1.21281f
C2084 sarlogic_0/_293_/a_36_472# vss 0.031137f
C2085 sarlogic_0/FILLER_0_5_128/a_484_472# vss 0.345058f
C2086 sarlogic_0/FILLER_0_5_128/a_36_472# vss 0.404746f
C2087 sarlogic_0/FILLER_0_5_128/a_572_375# vss 0.232991f
C2088 sarlogic_0/FILLER_0_5_128/a_124_375# vss 0.185089f
C2089 sarlogic_0/FILLER_0_5_117/a_36_472# vss 0.417394f
C2090 sarlogic_0/FILLER_0_5_117/a_124_375# vss 0.246306f
C2091 sarlogic_0/net7 vss 1.174913f
C2092 sarlogic_0/output7/a_224_472# vss 2.38465f
C2093 sarlogic_0/output42/a_224_472# vss 2.38465f
C2094 result[4] vss 24.779842f
C2095 sarlogic_0/net31 vss 1.912935f
C2096 sarlogic_0/output31/a_224_472# vss 2.38465f
C2097 sarlogic_0/output20/a_224_472# vss 2.38465f
C2098 sarlogic_0/FILLER_0_16_73/a_484_472# vss 0.345058f
C2099 sarlogic_0/FILLER_0_16_73/a_36_472# vss 0.404746f
C2100 sarlogic_0/FILLER_0_16_73/a_572_375# vss 0.232991f
C2101 sarlogic_0/FILLER_0_16_73/a_124_375# vss 0.185089f
C2102 sarlogic_0/FILLER_0_21_142/a_484_472# vss 0.345058f
C2103 sarlogic_0/FILLER_0_21_142/a_36_472# vss 0.404746f
C2104 sarlogic_0/FILLER_0_21_142/a_572_375# vss 0.232991f
C2105 sarlogic_0/FILLER_0_21_142/a_124_375# vss 0.185089f
C2106 sarlogic_0/FILLER_0_15_150/a_36_472# vss 0.417394f
C2107 sarlogic_0/FILLER_0_15_150/a_124_375# vss 0.246306f
C2108 sarlogic_0/FILLER_0_19_125/a_36_472# vss 0.417394f
C2109 sarlogic_0/FILLER_0_19_125/a_124_375# vss 0.246306f
C2110 sarlogic_0/net10 vss 1.481359f
C2111 sarlogic_0/net20 vss 2.034189f
C2112 sarlogic_0/_277_/a_36_160# vss 0.386641f
C2113 sarlogic_0/net27 vss 2.023744f
C2114 sarlogic_0/_004_ vss 0.390107f
C2115 sarlogic_0/_415_/a_2560_156# vss 0.016968f
C2116 sarlogic_0/_415_/a_2665_112# vss 0.62251f
C2117 sarlogic_0/_415_/a_2248_156# vss 0.371662f
C2118 sarlogic_0/_415_/a_1204_472# vss 0.012971f
C2119 sarlogic_0/_415_/a_1000_472# vss 0.291735f
C2120 sarlogic_0/_415_/a_796_472# vss 0.023206f
C2121 sarlogic_0/_415_/a_1308_423# vss 0.279043f
C2122 sarlogic_0/_415_/a_448_472# vss 0.684413f
C2123 sarlogic_0/_415_/a_36_151# vss 1.43589f
C2124 sarlogic_0/mask\[5\] vss 1.334568f
C2125 sarlogic_0/_346_/a_49_472# vss 0.054843f
C2126 sarlogic_0/_028_ vss 0.386029f
C2127 sarlogic_0/_363_/a_36_68# vss 0.150048f
C2128 sarlogic_0/_021_ vss 0.316776f
C2129 sarlogic_0/_432_/a_2560_156# vss 0.016968f
C2130 sarlogic_0/_432_/a_2665_112# vss 0.62251f
C2131 sarlogic_0/_432_/a_2248_156# vss 0.371662f
C2132 sarlogic_0/_432_/a_1204_472# vss 0.012971f
C2133 sarlogic_0/_432_/a_1000_472# vss 0.291735f
C2134 sarlogic_0/_432_/a_796_472# vss 0.023206f
C2135 sarlogic_0/_432_/a_1308_423# vss 0.279043f
C2136 sarlogic_0/_432_/a_448_472# vss 0.684413f
C2137 sarlogic_0/_432_/a_36_151# vss 1.43589f
C2138 sarlogic_0/_008_ vss 0.423631f
C2139 sarlogic_0/_104_ vss 1.435764f
C2140 sarlogic_0/_106_ vss 0.378703f
C2141 sarlogic_0/FILLER_0_17_200/a_484_472# vss 0.345058f
C2142 sarlogic_0/FILLER_0_17_200/a_36_472# vss 0.404746f
C2143 sarlogic_0/FILLER_0_17_200/a_572_375# vss 0.232991f
C2144 sarlogic_0/FILLER_0_17_200/a_124_375# vss 0.185089f
C2145 dacn_0/carray_n_0/n9 vss 14.559587f
C2146 dacn_0/out vss -0.682701p
C2147 dacn_0/carray_n_0/n8 vss 40.389835f
C2148 dacn_0/carray_n_0/n7 vss 57.16868f
C2149 dacn_0/carray_n_0/n6 vss 53.444874f
C2150 dacn_0/carray_n_0/n0 vss 17.398035f
C2151 dacn_0/carray_n_0/n1 vss 16.427063f
C2152 dacn_0/carray_n_0/n2 vss 30.239845f
C2153 dacn_0/carray_n_0/n3 vss 33.722244f
C2154 dacn_0/carray_n_0/n4 vss 39.983227f
C2155 dacn_0/carray_n_0/n5 vss 47.48966f
C2156 dacp_0/sample vss 0.104013p
C2157 dacn_0/bootstrapped_sw_n_0/vbsh vss 9.037161f
C2158 dacn_0/bootstrapped_sw_n_0/vbsl vss 8.446682f
C2159 dacn_0/bootstrapped_sw_n_0/vg vss 1.162193f
C2160 dacn_0/bootstrapped_sw_n_0/vs vss 0.065021f
C2161 dacn_0/bootstrapped_sw_n_0/enb vss 1.52928f
C2162 vinn vss 40.695953f
C2163 dacn_0/ctl9 vss 8.1548f
C2164 dacn_0/ctl8 vss 8.644266f
C2165 dacn_0/ctl7 vss 11.504689f
C2166 dacn_0/ctl6 vss 12.597453f
C2167 dacn_0/ctl5 vss 13.726896f
C2168 dacn_0/ctl4 vss 14.503242f
C2169 dacn_0/ctl3 vss 15.096921f
C2170 dacn_0/ctl1 vss 22.76591f
C2171 dacn_0/ctl10 vss 10.859402f
C2172 dacn_0/ctl2 vss 16.774553f
C2173 dacn_0/carray_n_0/ndum vss 14.881927f
C2174 latch_0/R vss 5.935133f
C2175 latch_0/S vss 7.551805f
C2176 comparator_0/trim_left_0/trim_switch_left_0/n0 vss 0.59175f
C2177 comparator_0/trim_left_0/trim_switch_left_0/n1 vss 0.614476f
C2178 comparator_0/trim_left_0/trim_switch_left_0/n4 vss 4.186667f
C2179 comparator_0/in vss -4.630677f
C2180 comparator_0/trim_left_0/trim_switch_left_0/n3 vss 3.310458f
C2181 comparator_0/trim_left_0/trim_switch_left_0/n2 vss 1.980191f
C2182 sarlogic_0/trim[0] vss 5.465488f
C2183 sarlogic_0/trim[1] vss 6.197476f
C2184 sarlogic_0/trim[2] vss 5.740468f
C2185 sarlogic_0/trim[3] vss 11.552049f
C2186 sarlogic_0/trim[4] vss 10.713926f
C2187 comparator_0/diff vss 0.155718f
C2188 buffer_0/out vss 7.9748f
C2189 sarlogic_0/trimb[4] vss 10.747439f
C2190 sarlogic_0/trimb[3] vss 10.092912f
C2191 sarlogic_0/trimb[2] vss 5.74902f
C2192 sarlogic_0/trimb[1] vss 5.811154f
C2193 sarlogic_0/trimb[0] vss 5.559114f
C2194 comparator_0/trim_right_0/trim_switch_right_0/XM0_trim_right_0/D vss 0.677622f
C2195 comparator_0/trim_right_0/trim_switch_right_0/XM1_trim_right_0/D vss 0.716105f
C2196 comparator_0/trim_right_0/trim_switch_right_0/XM4_trim_right_0/D vss 4.186667f
C2197 comparator_0/ip vss -4.6307f
C2198 comparator_0/trim_right_0/trim_switch_right_0/XM3_trim_right_0/D vss 3.310458f
C2199 comparator_0/trim_right_0/trim_switch_right_0/XM2_trim_right_0/D vss 1.980191f
C2200 dacp_0/carray_p_0/n2 vss 30.239845f
C2201 dacp_0/carray_p_0/n3 vss 33.722244f
C2202 dacp_0/carray_p_0/n4 vss 39.983227f
C2203 dacp_0/carray_p_0/n5 vss 47.48966f
C2204 dacp_0/carray_p_0/n9 vss 14.559587f
C2205 dacp_0/out vss -0.680742p
C2206 dacp_0/carray_p_0/n8 vss 40.389835f
C2207 dacp_0/carray_p_0/n7 vss 57.16868f
C2208 dacp_0/carray_p_0/n6 vss 53.444874f
C2209 dacp_0/carray_p_0/n0 vss 17.398035f
C2210 dacp_0/carray_p_0/n1 vss 16.427063f
C2211 dacp_0/bootstrapped_sw_p_0/vs vss 0.065021f
C2212 dacp_0/bootstrapped_sw_p_0/enb vss 1.52928f
C2213 dacp_0/bootstrapped_sw_p_0/vg vss 1.162193f
C2214 dacp_0/bootstrapped_sw_p_0/vbsh vss 9.037161f
C2215 dacp_0/bootstrapped_sw_p_0/vbsl vss 8.446682f
C2216 vinp vss 40.695305f
C2217 dacp_0/ctl9 vss 7.725754f
C2218 dacp_0/ctl8 vss 8.39172f
C2219 dacp_0/ctl7 vss 11.074413f
C2220 dacp_0/ctl6 vss 12.387031f
C2221 dacp_0/ctl5 vss 13.424606f
C2222 dacp_0/ctl4 vss 13.417045f
C2223 dacp_0/ctl3 vss 15.41302f
C2224 dacp_0/ctl1 vss 21.83176f
C2225 dacp_0/ctl10 vss 10.44588f
C2226 dacp_0/ctl2 vss 15.116745f
C2227 dacp_0/carray_p_0/ndum vss 14.881927f
C2228 buffer_0/middle vss 0.926667f
C2229 buffer_0/in vss 6.778908f
C2230 buffer_0/buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vss 0.17777f
C2231 latch_0/Qn vss 0.762147f
C2232 latch_0/Q vss 7.041345f
C2233 latch_0/tutyuu2 vss 0.613078f
C2234 latch_0/tutyuu1 vss 0.612955f
.ends

