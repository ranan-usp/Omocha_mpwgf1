* NGSPICE file created from saradc.ext - technology: gf180mcuD

.subckt XM2$3$1 a_n36_120# a_n116_n100# w_n460_n310# VSUBS
X0 w_n460_n310# a_n36_120# a_n116_n100# w_n460_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_n100# w_n460_n310# 0.09188f
C1 a_n36_120# w_n460_n310# 0.143803f
C2 a_n116_n100# a_n36_120# 0.001764f
C3 a_n116_n100# VSUBS 0.04225f
C4 a_n36_120# VSUBS 0.082818f
C5 w_n460_n310# VSUBS 1.56551f
.ends

.subckt XM1$3$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_28_n200# a_n36_20# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134096f
C2 a_n36_20# a_n254_n386# 0.226575f
.ends

.subckt x4 out in vdd vss
XXM2$3$1_0 in out vdd vss XM2$3$1
XXM1$3$1_0 in vss out XM1$3$1
C0 out in 0.057341f
C1 in vdd 0.039699f
C2 vss in 0.018605f
C3 out vdd 0.102755f
C4 out vss 0.048617f
C5 vss vdd 0.057876f
C6 vss 0 0.19553f
C7 vdd 0 1.704834f
C8 out 0 0.450443f
C9 in 0 0.431461f
.ends

.subckt XM2$1$3 a_n36_120# a_n116_n100# w_n278_n310# VSUBS
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 w_n278_n310# a_n36_120# 0.143685f
C1 w_n278_n310# a_n116_n100# 0.090454f
C2 a_n116_n100# a_n36_120# 0.001764f
C3 a_n116_n100# VSUBS 0.043675f
C4 a_n36_120# VSUBS 0.082818f
C5 w_n278_n310# VSUBS 1.57235f
.ends

.subckt XM1$1$3 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n36_20# a_28_n200# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134096f
C2 a_n36_20# a_n254_n386# 0.22648f
.ends

.subckt x2 out in vdd vss
XXM2$1$3_0 in out vdd vss XM2$1$3
XXM1$1$3_0 in vss out XM1$1$3
C0 vss vdd 0.057427f
C1 vdd in 0.039609f
C2 vss in 0.017815f
C3 out vdd 0.093301f
C4 out vss 0.045442f
C5 out in 0.057341f
C6 vss 0 0.200924f
C7 vdd 0 1.717231f
C8 out 0 0.463681f
C9 in 0 0.432083f
.ends

.subckt XM4$5 a_540_n1607# a_258_n1293# a_258_n1793# a_396_n1607# a_476_n1387#
X0 a_540_n1607# a_476_n1387# a_396_n1607# a_258_n1793# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_396_n1607# a_540_n1607# 0.06854f
C1 a_476_n1387# a_396_n1607# 0.001764f
C2 a_476_n1387# a_540_n1607# 0.001764f
C3 a_540_n1607# a_258_n1793# 0.065139f
C4 a_396_n1607# a_258_n1793# 0.065139f
C5 a_476_n1387# a_258_n1793# 0.220578f
.ends

.subckt XM3$5 a_n67_n1582# a_n349_n1268# a_n131_n1362# a_n211_n1582# a_n349_n1768#
X0 a_n67_n1582# a_n131_n1362# a_n211_n1582# a_n349_n1768# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n211_n1582# a_n67_n1582# 0.06854f
C1 a_n131_n1362# a_n211_n1582# 0.001764f
C2 a_n131_n1362# a_n67_n1582# 0.001764f
C3 a_n67_n1582# a_n349_n1768# 0.065139f
C4 a_n211_n1582# a_n349_n1768# 0.065139f
C5 a_n131_n1362# a_n349_n1768# 0.220578f
.ends

.subckt XM2$2$1 a_n36_120# a_n116_n100# w_n460_n310# VSUBS
X0 w_n460_n310# a_n36_120# a_n116_n100# w_n460_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_n100# w_n460_n310# 0.09188f
C1 a_n36_120# a_n116_n100# 0.001764f
C2 a_n36_120# w_n460_n310# 0.143803f
C3 a_n116_n100# VSUBS 0.04225f
C4 a_n36_120# VSUBS 0.082818f
C5 w_n460_n310# VSUBS 1.56551f
.ends

.subckt XM1$2$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_28_n200# a_n36_20# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134096f
C2 a_n36_20# a_n254_n386# 0.226575f
.ends

.subckt x3 out in vdd vss
XXM2$2$1_0 in out vdd vss XM2$2$1
XXM1$2$1_0 in vss out XM1$2$1
C0 in vdd 0.039699f
C1 in vss 0.018605f
C2 in out 0.057341f
C3 vdd vss 0.057622f
C4 out vdd 0.102755f
C5 out vss 0.048617f
C6 vss 0 0.194402f
C7 vdd 0 1.705041f
C8 out 0 0.450443f
C9 in 0 0.431461f
.ends

.subckt XM1$5 a_n36_20# a_n254_n386# a_n254_114# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_28_n200# a_n36_20# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134096f
C2 a_n36_20# a_n254_n386# 0.22648f
.ends

.subckt XM2$5 a_n36_120# a_n116_n100# w_n278_n310# VSUBS
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_n100# a_n36_120# 0.001764f
C1 a_n116_n100# w_n278_n310# 0.090454f
C2 w_n278_n310# a_n36_120# 0.143685f
C3 a_n116_n100# VSUBS 0.043675f
C4 a_n36_120# VSUBS 0.082818f
C5 w_n278_n310# VSUBS 1.57235f
.ends

.subckt x1 out in vdd XM1$5_0/a_n254_114# vss
XXM1$5_0 in vss XM1$5_0/a_n254_114# out XM1$5
XXM2$5_0 in out vdd vss XM2$5
C0 vdd out 0.093301f
C1 out in 0.057341f
C2 vss vdd 0.057306f
C3 vss in 0.017815f
C4 vdd in 0.039609f
C5 vss out 0.045442f
C6 vss 0 0.1996f
C7 out 0 0.463681f
C8 in 0 0.432083f
C9 vdd 0 1.717231f
.ends

.subckt latch Qn Q S R XM3$5_0/a_n211_n1582# x3_0/out x4_0/out XM4$5_0/a_540_n1607#
+ VSUBS
Xx4_0 x4_0/out S Q VSUBS x4
Xx2_0 Qn Q Q VSUBS x2
XXM4$5_0 XM4$5_0/a_540_n1607# VSUBS VSUBS Q x3_0/out XM4$5
XXM3$5_0 Qn VSUBS x4_0/out XM3$5_0/a_n211_n1582# VSUBS XM3$5
Xx3_0 x3_0/out R Q VSUBS x3
Xx1_0 Q Qn Q VSUBS VSUBS x1
C0 S VSUBS 0.033653f
C1 Q R 0.065254f
C2 S x4_0/out 0.115854f
C3 VSUBS x4_0/out 0.056312f
C4 S Q 0.053978f
C5 VSUBS Q 0.081616f
C6 x3_0/out XM4$5_0/a_540_n1607# 0.05058f
C7 x3_0/out R 0.115854f
C8 Qn XM4$5_0/a_540_n1607# 0.001478f
C9 Q x4_0/out 0.162322f
C10 VSUBS x3_0/out 0.056312f
C11 VSUBS XM3$5_0/a_n211_n1582# 0.004577f
C12 S Qn 0.011276f
C13 Qn VSUBS 0.201264f
C14 Q x3_0/out 0.210824f
C15 XM3$5_0/a_n211_n1582# x4_0/out 0.05058f
C16 Q XM3$5_0/a_n211_n1582# 0.002119f
C17 Qn x4_0/out 0.109327f
C18 Qn Q 1.569045f
C19 Qn x3_0/out 0.060761f
C20 VSUBS XM4$5_0/a_540_n1607# 0.004577f
C21 VSUBS R 0.033653f
C22 x3_0/out 0 0.589125f
C23 R 0 0.441972f
C24 XM3$5_0/a_n211_n1582# 0 0.065139f
C25 XM4$5_0/a_540_n1607# 0 0.065139f
C26 VSUBS 0 0.306028f
C27 Qn 0 0.639183f
C28 Q 0 6.695502f
C29 x4_0/out 0 0.589061f
C30 S 0 0.441972f
.ends

.subckt XM2$6 a_n36_120# a_n116_n100# w_n278_n310# VSUBS
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_n100# w_n278_n310# 0.090564f
C1 a_n36_120# w_n278_n310# 0.138578f
C2 a_n36_120# a_n116_n100# 0.001764f
C3 a_n116_n100# VSUBS 0.043675f
C4 a_n36_120# VSUBS 0.08816f
C5 w_n278_n310# VSUBS 1.2321f
.ends

.subckt XM1$6 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_28_n200# a_n36_20# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134177f
C2 a_n36_20# a_n254_n386# 0.22667f
.ends

.subckt inv$2 out in vdd vss
XXM2$6_0 in out vdd vss XM2$6
XXM1$6_0 in vss out XM1$6
C0 vss vdd 0.050184f
C1 vss out 0.056311f
C2 in vss 0.019395f
C3 out vdd 0.086562f
C4 in vdd 0.034991f
C5 in out 0.057341f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt buffer in out inv$2_1/in inv$2_1/vdd VSUBS
Xinv$2_0 inv$2_1/in in inv$2_1/vdd VSUBS inv$2
Xinv$2_1 out inv$2_1/in inv$2_1/vdd VSUBS inv$2
C0 VSUBS in 0.033849f
C1 inv$2_1/in in 0.118184f
C2 out VSUBS 0.027914f
C3 out inv$2_1/in 0.160621f
C4 inv$2_1/vdd VSUBS -0.035287f
C5 inv$2_1/vdd inv$2_1/in 0.122776f
C6 inv$2_1/vdd in 0.051816f
C7 VSUBS inv$2_1/in 0.084611f
C8 inv$2_1/vdd out 0.042403f
C9 out 0 0.544428f
C10 VSUBS 0 0.247812f
C11 inv$2_1/vdd 0 2.60626f
C12 inv$2_1/in 0 0.821157f
C13 in 0 0.478121f
.ends

.subckt XM3 a_n3152_1140# a_n3064_1048# w_n3314_932# a_n2964_1140# VSUBS
X0 a_n2964_1140# a_n3064_1048# a_n3152_1140# w_n3314_932# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 w_n3314_932# a_n2964_1140# 0.009117f
C1 a_n3064_1048# a_n3152_1140# 0.002993f
C2 a_n3152_1140# w_n3314_932# 0.008969f
C3 a_n3152_1140# a_n2964_1140# 0.103318f
C4 a_n3064_1048# w_n3314_932# 0.157732f
C5 a_n3064_1048# a_n2964_1140# 0.002993f
C6 a_n2964_1140# VSUBS 0.100353f
C7 a_n3152_1140# VSUBS 0.100353f
C8 a_n3064_1048# VSUBS 0.130702f
C9 w_n3314_932# VSUBS 1.4688f
.ends

.subckt XM1 a_912_4129# a_995_4229# a_811_3903# a_1507_3903# a_995_4041#
X0 a_995_4229# a_912_4129# a_995_4041# a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_995_4229# a_912_4129# 0.002993f
C1 a_912_4129# a_995_4041# 0.002993f
C2 a_995_4229# a_995_4041# 0.103318f
C3 a_995_4041# a_811_3903# 0.109266f
C4 a_912_4129# a_811_3903# 0.288275f
C5 a_995_4229# a_811_3903# 0.109266f
.ends

.subckt XMs a_1030_4680# a_1030_4868# a_947_4768# a_846_4542#
X0 a_1030_4868# a_947_4768# a_1030_4680# a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_947_4768# a_1030_4680# 0.002993f
C1 a_1030_4680# a_1030_4868# 0.103318f
C2 a_947_4768# a_1030_4868# 0.002993f
C3 a_1030_4680# a_846_4542# 0.387117f
C4 a_947_4768# a_846_4542# 0.288368f
C5 a_1030_4868# a_846_4542# 0.109266f
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668# VSUBS
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0_m4m5_noshield c_width=8u c_length=8u
C0 m4_n3440_n548# m4_n3800_n668# 0.646322f
C1 m4_n3440_n548# VSUBS 1.17298f
C2 m4_n3800_n668# VSUBS 1.64833f
.ends

.subckt sw_cap_unit in out VSUBS
Xcap_mim_2p0fF_8JNR63_0 out in VSUBS cap_mim_2p0fF_8JNR63
C0 out VSUBS 1.17298f
C1 in VSUBS 1.64833f
.ends

.subckt sw_cap out in VSUBS
Xsw_cap_unit_0 in out VSUBS sw_cap_unit
Xsw_cap_unit_1 in out VSUBS sw_cap_unit
Xsw_cap_unit_2 in out VSUBS sw_cap_unit
Xsw_cap_unit_3 in out VSUBS sw_cap_unit
Xsw_cap_unit_4 in out VSUBS sw_cap_unit
C0 out in 2.231591f
C1 out VSUBS 6.064711f
C2 in VSUBS 7.39096f
.ends

.subckt XMs1 a_n2529_n616# a_n2717_n616# a_n2629_n699# a_n2855_n800#
X0 a_n2529_n616# a_n2629_n699# a_n2717_n616# a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n2529_n616# a_n2629_n699# 0.002993f
C1 a_n2717_n616# a_n2629_n699# 0.002993f
C2 a_n2717_n616# a_n2529_n616# 0.103318f
C3 a_n2529_n616# a_n2855_n800# 0.109266f
C4 a_n2717_n616# a_n2855_n800# 0.177295f
C5 a_n2629_n699# a_n2855_n800# 0.288368f
.ends

.subckt XM4 a_n2550_442# a_n2362_442# w_n2712_234# a_n2462_359# VSUBS
X0 a_n2362_442# a_n2462_359# a_n2550_442# w_n2712_234# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n2362_442# w_n2712_234# 0.008969f
C1 a_n2550_442# a_n2362_442# 0.103318f
C2 a_n2462_359# a_n2362_442# 0.002993f
C3 a_n2550_442# w_n2712_234# 0.058295f
C4 a_n2462_359# w_n2712_234# 0.173648f
C5 a_n2462_359# a_n2550_442# 0.002993f
C6 a_n2362_442# VSUBS 0.100353f
C7 a_n2550_442# VSUBS 0.119847f
C8 a_n2462_359# VSUBS 0.147064f
C9 w_n2712_234# VSUBS 1.4688f
.ends

.subckt XM2_inv a_n36_120# a_n116_n100# w_n278_n310# VSUBS
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_n100# w_n278_n310# 0.090564f
C1 a_n36_120# w_n278_n310# 0.138578f
C2 a_n36_120# a_n116_n100# 0.001764f
C3 a_n116_n100# VSUBS 0.043675f
C4 a_n36_120# VSUBS 0.08816f
C5 w_n278_n310# VSUBS 1.2321f
.ends

.subckt XM1_inv a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_28_n200# a_n36_20# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134177f
C2 a_n36_20# a_n254_n386# 0.22667f
.ends

.subckt inv out in vdd vss
XXM2_inv_0 in out vdd vss XM2_inv
XXM1_inv_0 in vss out XM1_inv
C0 out vss 0.056311f
C1 in vss 0.019395f
C2 vss vdd 0.050184f
C3 in out 0.057341f
C4 out vdd 0.086562f
C5 in vdd 0.034991f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt XM2 a_912_3686# a_811_3460# a_995_3786# a_1507_3460# a_995_3598#
X0 a_995_3786# a_912_3686# a_995_3598# a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_912_3686# a_995_3786# 0.002993f
C1 a_995_3598# a_995_3786# 0.103318f
C2 a_995_3598# a_912_3686# 0.002993f
C3 a_995_3598# a_811_3460# 0.109266f
C4 a_912_3686# a_811_3460# 0.288275f
C5 a_995_3786# a_811_3460# 0.109266f
.ends

.subckt XMs2 a_n3762_561# a_n3988_469# a_n3662_653# a_n3850_653# a_n3988_1165#
X0 a_n3662_653# a_n3762_561# a_n3850_653# a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n3850_653# a_n3762_561# 0.002993f
C1 a_n3662_653# a_n3762_561# 0.002993f
C2 a_n3662_653# a_n3850_653# 0.103318f
C3 a_n3662_653# a_n3988_469# 0.109266f
C4 a_n3850_653# a_n3988_469# 0.109266f
C5 a_n3762_561# a_n3988_469# 0.288275f
.ends

.subckt bootstrapped_sw in vdd vss en enb out vs vg vbsh vbsl
XXM3_0 vbsh vg XM4_0/w_n2712_234# vdd vss XM3
XXM1_0 vg vbsl vss vss in XM1
XXMs_0 out in vg vss XMs
Xsw_cap_0 vbsh vbsl vss sw_cap
XXMs1_0 vs vg vdd vss XMs1
XXM4_0 vg vbsh XM4_0/w_n2712_234# enb vss XM4
Xinv_0 enb en vdd vss inv
XXM2_0 enb vss vss vss vbsl XM2
XXMs2_0 enb vss vss vs vss XMs2
C0 XM4_0/w_n2712_234# vdd 0.079362f
C1 vbsh out 0.100712f
C2 vs vbsl 0.001422f
C3 XM4_0/w_n2712_234# out 0.005706f
C4 vdd vg 0.447812f
C5 vbsh enb 0.052707f
C6 XM4_0/w_n2712_234# vbsh 0.101815f
C7 vbsl vdd 0.005409f
C8 vg out 0.04429f
C9 XM4_0/w_n2712_234# enb 0.041524f
C10 vbsh vg 0.144325f
C11 vbsl out 0.058082f
C12 in vbsh 0.008752f
C13 en vdd 0.065092f
C14 vg enb 0.612109f
C15 XM4_0/w_n2712_234# vg 0.080093f
C16 vbsl vbsh 0.025766f
C17 vbsl enb 0.017274f
C18 XM4_0/w_n2712_234# vbsl 0.009881f
C19 vs enb 0.00376f
C20 vdd out 0.017908f
C21 in vg 0.075595f
C22 vbsl vg 0.046114f
C23 vdd vbsh 0.168905f
C24 vs vg 0.01049f
C25 en enb 0.029269f
C26 in vbsl 0.299565f
C27 vdd enb 0.448382f
C28 out vss 1.088543f
C29 vs vss 0.072259f
C30 enb vss 1.595319f
C31 vdd vss 3.106074f
C32 en vss 0.642295f
C33 XM4_0/w_n2712_234# vss 1.968192f
C34 vbsh vss 7.100617f
C35 vbsl vss 8.368301f
C36 in vss 0.308876f
C37 vg vss 1.218873f
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VSS ZN 0.180794f
C1 VNW ZN 0.023676f
C2 VDD ZN 0.271625f
C3 VDD VSS 0.029045f
C4 VDD VNW 0.082022f
C5 VNW VSS 0.006277f
C6 I ZN 0.58604f
C7 VDD I 0.074838f
C8 VSS I 0.091531f
C9 VNW I 0.285482f
C10 VSS VPW 0.296769f
C11 ZN VPW 0.099188f
C12 VDD VPW 0.238483f
C13 I VPW 0.610668f
C14 VNW VPW 1.31158f
.ends

.subckt dummy VSS ZN I VDD VNW VPW
X0 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VDD ZN 0.271625f
C1 VNW ZN 0.026913f
C2 VSS ZN 0.180794f
C3 VDD VNW 0.108083f
C4 VDD VSS 0.035859f
C5 VNW VSS 0.011638f
C6 I ZN 0.58604f
C7 VDD I 0.075475f
C8 VNW I 0.291591f
C9 VSS I 0.092168f
C10 VSS VPW 0.337898f
C11 ZN VPW 0.095951f
C12 VDD VPW 0.258911f
C13 I VPW 0.604559f
C14 VNW VPW 1.53535f
.ends

.subckt inv_renketu dummy_1/I inv$1_8/I inv$1_1/I inv$1_3/I dummy_0/ZN inv$1_5/I dummy_0/I
+ inv$1_7/I inv$1_9/ZN inv$1_6/ZN inv$1_0/ZN inv$1_9/VNW inv$1_0/I inv$1_4/ZN inv$1_9/I
+ inv$1_2/I inv$1_10/I inv$1_7/ZN inv$1_1/ZN inv$1_3/ZN inv$1_4/I inv$1_8/ZN inv$1_9/VSS
+ inv$1_9/VDD inv$1_10/ZN VSUBS inv$1_6/I inv$1_2/ZN inv$1_5/ZN
Xinv$1_10 inv$1_9/VSS inv$1_10/ZN inv$1_10/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_0 inv$1_9/VSS inv$1_0/ZN inv$1_0/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_1 inv$1_9/VSS inv$1_1/ZN inv$1_1/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_2 inv$1_9/VSS inv$1_2/ZN inv$1_2/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_3 inv$1_9/VSS inv$1_3/ZN inv$1_3/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_4 inv$1_9/VSS inv$1_4/ZN inv$1_4/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_5 inv$1_9/VSS inv$1_5/ZN inv$1_5/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_6 inv$1_9/VSS inv$1_6/ZN inv$1_6/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_7 inv$1_9/VSS inv$1_7/ZN inv$1_7/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_8 inv$1_9/VSS inv$1_8/ZN inv$1_8/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xinv$1_9 inv$1_9/VSS inv$1_9/ZN inv$1_9/I inv$1_9/VDD inv$1_9/VNW VSUBS inv$1
Xdummy_0 inv$1_9/VSS dummy_0/ZN dummy_0/I inv$1_9/VDD inv$1_9/VNW VSUBS dummy
Xdummy_1 inv$1_9/VSS dummy_1/ZN dummy_1/I inv$1_9/VDD inv$1_9/VNW VSUBS dummy
C0 inv$1_9/ZN inv$1_8/ZN 0.161793f
C1 inv$1_9/VNW dummy_0/ZN -0.002275f
C2 inv$1_9/VNW inv$1_10/I 0.010403f
C3 inv$1_3/ZN inv$1_0/ZN 0.161792f
C4 inv$1_9/VSS inv$1_6/I 0.104553f
C5 inv$1_9/VNW inv$1_0/I 0.011179f
C6 inv$1_9/VNW inv$1_4/I 0.010403f
C7 inv$1_9/VDD inv$1_9/ZN 0.104396f
C8 inv$1_9/ZN inv$1_10/ZN 0.161792f
C9 inv$1_0/ZN inv$1_9/VSS 0.003829f
C10 inv$1_3/I inv$1_9/VDD 0.00333f
C11 inv$1_6/ZN inv$1_5/ZN 0.161792f
C12 inv$1_9/VDD inv$1_5/ZN 0.104396f
C13 inv$1_4/ZN inv$1_9/VDD 0.104396f
C14 inv$1_7/ZN inv$1_8/I 0.002086f
C15 inv$1_3/ZN inv$1_9/VNW 0.006066f
C16 inv$1_3/I inv$1_1/ZN 0.028928f
C17 inv$1_0/I dummy_0/I 0.017781f
C18 inv$1_9/VNW inv$1_9/VSS -0.005361f
C19 inv$1_9/ZN inv$1_10/I 0.002086f
C20 inv$1_1/ZN inv$1_4/ZN 0.161792f
C21 inv$1_8/ZN inv$1_7/I 0.028928f
C22 inv$1_8/ZN inv$1_9/I 0.002086f
C23 inv$1_6/I inv$1_7/ZN 0.028928f
C24 inv$1_3/I inv$1_0/I 0.084161f
C25 inv$1_6/ZN inv$1_7/I 0.002086f
C26 inv$1_9/VDD inv$1_7/I 0.00333f
C27 inv$1_4/I inv$1_5/ZN 0.028928f
C28 inv$1_9/I inv$1_10/ZN 0.028928f
C29 inv$1_9/VDD inv$1_9/I 0.00333f
C30 inv$1_5/I inv$1_6/ZN 0.028928f
C31 inv$1_4/I inv$1_4/ZN 0.031424f
C32 inv$1_5/I inv$1_9/VDD 0.00333f
C33 inv$1_9/VNW inv$1_8/I 0.010403f
C34 inv$1_2/I inv$1_9/VDD 0.00333f
C35 inv$1_3/ZN inv$1_3/I 0.031424f
C36 inv$1_2/I inv$1_10/ZN 0.002086f
C37 inv$1_9/VNW inv$1_1/I 0.010403f
C38 inv$1_9/VDD inv$1_8/ZN 0.104396f
C39 inv$1_9/VSS inv$1_9/ZN 0.003829f
C40 inv$1_9/VNW inv$1_7/ZN 0.006066f
C41 inv$1_3/I inv$1_9/VSS 0.104553f
C42 inv$1_2/I inv$1_2/ZN 0.031424f
C43 inv$1_9/VNW dummy_1/ZN -0.001925f
C44 inv$1_2/I dummy_1/I 0.021288f
C45 inv$1_9/VSS inv$1_5/ZN 0.003829f
C46 inv$1_9/VSS inv$1_4/ZN 0.003829f
C47 inv$1_9/VNW inv$1_6/I 0.010403f
C48 inv$1_9/I inv$1_10/I 0.084161f
C49 inv$1_9/VDD inv$1_6/ZN 0.104396f
C50 inv$1_2/I inv$1_10/I 0.084161f
C51 inv$1_9/VDD inv$1_10/ZN 0.104396f
C52 inv$1_9/VNW inv$1_0/ZN 0.008403f
C53 inv$1_5/I inv$1_4/I 0.084161f
C54 inv$1_9/ZN inv$1_8/I 0.028928f
C55 inv$1_2/ZN inv$1_9/VDD 0.107277f
C56 inv$1_2/ZN inv$1_10/ZN 0.161793f
C57 inv$1_3/I inv$1_1/I 0.084161f
C58 inv$1_1/ZN inv$1_9/VDD 0.104396f
C59 inv$1_1/I inv$1_4/ZN 0.028928f
C60 inv$1_9/VDD dummy_0/ZN 0.001671f
C61 inv$1_9/VDD inv$1_10/I 0.00333f
C62 inv$1_10/I inv$1_10/ZN 0.031424f
C63 inv$1_9/VSS inv$1_7/I 0.104553f
C64 inv$1_9/VSS inv$1_9/I 0.104553f
C65 inv$1_2/ZN dummy_1/I 0.003027f
C66 inv$1_5/I inv$1_9/VSS 0.104553f
C67 inv$1_0/I inv$1_9/VDD 0.00333f
C68 inv$1_9/VSS inv$1_2/I 0.107646f
C69 inv$1_0/ZN dummy_0/I 0.023262f
C70 inv$1_6/I inv$1_5/ZN 0.002086f
C71 inv$1_4/I inv$1_9/VDD 0.00333f
C72 inv$1_2/ZN inv$1_10/I 0.028928f
C73 inv$1_9/VSS inv$1_8/ZN 0.003829f
C74 inv$1_3/I inv$1_0/ZN 0.002086f
C75 inv$1_3/ZN inv$1_9/VDD 0.104396f
C76 inv$1_8/I inv$1_7/I 0.084161f
C77 inv$1_8/I inv$1_9/I 0.084161f
C78 inv$1_0/I dummy_0/ZN 0.002409f
C79 inv$1_4/I inv$1_1/ZN 0.002086f
C80 inv$1_9/VSS inv$1_6/ZN 0.003829f
C81 inv$1_9/VSS inv$1_10/ZN 0.003829f
C82 inv$1_9/VSS inv$1_9/VDD -0.006814f
C83 inv$1_9/VNW inv$1_9/ZN 0.006066f
C84 inv$1_9/VNW inv$1_3/I 0.010403f
C85 inv$1_3/ZN inv$1_1/ZN 0.161793f
C86 inv$1_7/ZN inv$1_7/I 0.031424f
C87 inv$1_8/ZN inv$1_8/I 0.031424f
C88 inv$1_9/VNW inv$1_5/ZN 0.006066f
C89 inv$1_9/VNW inv$1_4/ZN 0.006066f
C90 inv$1_9/VSS inv$1_2/ZN 0.003829f
C91 inv$1_6/I inv$1_7/I 0.084161f
C92 inv$1_2/I dummy_1/ZN 0.027478f
C93 inv$1_5/I inv$1_6/I 0.084161f
C94 inv$1_3/ZN inv$1_0/I 0.028928f
C95 inv$1_9/VSS inv$1_1/ZN 0.003829f
C96 inv$1_7/ZN inv$1_8/ZN 0.161792f
C97 inv$1_9/VSS dummy_0/ZN 0.001445f
C98 inv$1_9/VSS inv$1_10/I 0.104553f
C99 inv$1_9/VDD inv$1_8/I 0.00333f
C100 inv$1_9/VSS inv$1_0/I 0.108299f
C101 inv$1_1/I inv$1_9/VDD 0.00333f
C102 inv$1_4/I inv$1_9/VSS 0.104553f
C103 inv$1_6/ZN inv$1_7/ZN 0.161793f
C104 inv$1_9/VDD inv$1_7/ZN 0.104396f
C105 inv$1_9/VDD dummy_1/ZN 0.010249f
C106 inv$1_6/I inv$1_6/ZN 0.031424f
C107 inv$1_6/I inv$1_9/VDD 0.00333f
C108 inv$1_9/VNW inv$1_9/I 0.010403f
C109 inv$1_9/VNW inv$1_7/I 0.010403f
C110 inv$1_3/ZN inv$1_9/VSS 0.003829f
C111 inv$1_5/I inv$1_9/VNW 0.010403f
C112 inv$1_1/I inv$1_1/ZN 0.031424f
C113 inv$1_9/VNW inv$1_2/I 0.011789f
C114 inv$1_2/ZN dummy_1/ZN 0.022956f
C115 inv$1_4/ZN inv$1_5/ZN 0.161793f
C116 inv$1_0/ZN inv$1_9/VDD 0.107658f
C117 inv$1_9/VNW inv$1_8/ZN 0.006066f
C118 inv$1_4/I inv$1_1/I 0.084161f
C119 inv$1_9/VNW inv$1_6/ZN 0.006066f
C120 inv$1_3/ZN inv$1_1/I 0.002086f
C121 inv$1_9/VNW inv$1_10/ZN 0.006066f
C122 inv$1_9/VNW inv$1_9/VDD -0.157887f
C123 inv$1_0/ZN dummy_0/ZN 0.0229f
C124 inv$1_9/ZN inv$1_9/I 0.031424f
C125 inv$1_9/VSS inv$1_8/I 0.104553f
C126 inv$1_0/ZN inv$1_0/I 0.031424f
C127 inv$1_9/VSS inv$1_1/I 0.104553f
C128 inv$1_9/VNW inv$1_2/ZN 0.008692f
C129 inv$1_5/I inv$1_5/ZN 0.031424f
C130 inv$1_5/I inv$1_4/ZN 0.002086f
C131 inv$1_9/VNW inv$1_1/ZN 0.006066f
C132 inv$1_9/VSS inv$1_7/ZN 0.003829f
C133 dummy_1/ZN VSUBS 0.095951f
C134 dummy_1/I VSUBS 0.604559f
C135 dummy_0/ZN VSUBS 0.095951f
C136 dummy_0/I VSUBS 0.604559f
C137 inv$1_9/ZN VSUBS 0.260352f
C138 inv$1_9/I VSUBS 0.670517f
C139 inv$1_8/ZN VSUBS 0.260352f
C140 inv$1_8/I VSUBS 0.670517f
C141 inv$1_7/ZN VSUBS 0.260352f
C142 inv$1_7/I VSUBS 0.670517f
C143 inv$1_6/ZN VSUBS 0.260352f
C144 inv$1_6/I VSUBS 0.670517f
C145 inv$1_5/ZN VSUBS 0.260352f
C146 inv$1_5/I VSUBS 0.670517f
C147 inv$1_4/ZN VSUBS 0.260352f
C148 inv$1_4/I VSUBS 0.670517f
C149 inv$1_3/ZN VSUBS 0.260352f
C150 inv$1_3/I VSUBS 0.670517f
C151 inv$1_9/VSS VSUBS 2.848055f
C152 inv$1_2/ZN VSUBS 0.398879f
C153 inv$1_9/VDD VSUBS 2.113035f
C154 inv$1_2/I VSUBS 0.741957f
C155 inv$1_9/VNW VSUBS 14.066851f
C156 inv$1_1/ZN VSUBS 0.260352f
C157 inv$1_1/I VSUBS 0.670517f
C158 inv$1_0/ZN VSUBS 0.398674f
C159 inv$1_0/I VSUBS 0.735921f
C160 inv$1_10/ZN VSUBS 0.260352f
C161 inv$1_10/I VSUBS 0.670517f
.ends

.subckt dacp ctl0 in dum ctl2 ctl1 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 out ndum n1
+ n2 n3 n4 n5 n6 n7 n8 n9 sample bootstrapped_sw_0/vbsl bootstrapped_sw_0/vbsh n0
+ vdd vss
Xbootstrapped_sw_0 in vdd vss sample bootstrapped_sw_0/enb out bootstrapped_sw_0/vs
+ bootstrapped_sw_0/vg bootstrapped_sw_0/vbsh bootstrapped_sw_0/vbsl bootstrapped_sw
Xinv_renketu_0 inv_renketu_0/dummy_1/I ctl7 ctl2 ctl1 inv_renketu_0/dummy_0/ZN ctl4
+ inv_renketu_0/dummy_0/I ctl6 n8 n5 ndum inv_renketu_0/inv$1_9/VNW dum n3 ctl8 ctl0
+ ctl9 n6 n2 n1 ctl3 n7 inv_renketu_0/inv$1_9/VSS inv_renketu_0/inv$1_9/VDD n9 vss
+ ctl5 n0 n4 inv_renketu
C0 n0 inv_renketu_0/inv$1_9/VDD 0.008798f
C1 n9 n1 0.349226f
C2 n6 inv_renketu_0/inv$1_9/VDD 0.001148f
C3 inv_renketu_0/inv$1_9/VNW n0 0.002542f
C4 inv_renketu_0/inv$1_9/VDD ndum 0.001148f
C5 n7 n2 0.485327f
C6 bootstrapped_sw_0/vbsh out 0.137967f
C7 n5 n2 0.208084f
C8 inv_renketu_0/inv$1_9/VSS ctl0 0.002242f
C9 n9 n0 0.184985f
C10 n8 n4 2.84323f
C11 n9 n6 14.716789f
C12 n3 n2 22.840685f
C13 n7 n5 3.36878f
C14 sample inv_renketu_0/dummy_0/I 0.008276f
C15 inv_renketu_0/inv$1_9/VSS ctl1 0.002242f
C16 n9 ndum 0.127951f
C17 n2 out 6.640605f
C18 n3 n7 0.891504f
C19 n2 n1 16.604633f
C20 n3 n5 0.346757f
C21 n8 inv_renketu_0/inv$1_9/VDD 0.001148f
C22 ctl3 inv_renketu_0/inv$1_9/VSS 0.002242f
C23 n7 out 0.210031p
C24 n5 out 52.565514f
C25 n7 n1 0.212006f
C26 sample inv_renketu_0/inv$1_9/VSS 0.011446f
C27 n5 n1 0.141538f
C28 inv_renketu_0/inv$1_9/VSS ctl5 0.002242f
C29 n4 inv_renketu_0/inv$1_9/VDD 0.001148f
C30 sample ndum 0.046157f
C31 n3 out 13.201303f
C32 n2 n0 0.099287f
C33 ctl7 ctl8 0.076437f
C34 ctl6 ctl5 0.076437f
C35 n3 n1 0.144232f
C36 n6 n2 0.207962f
C37 n9 n8 87.102684f
C38 ctl1 ctl2 0.076437f
C39 n7 n0 0.06073f
C40 n1 out 3.367623f
C41 n5 n0 0.025424f
C42 n2 ndum 0.041162f
C43 n6 n7 34.326103f
C44 n6 n5 28.589401f
C45 ctl0 ctl9 0.076437f
C46 n9 n4 3.740573f
C47 ctl3 ctl2 0.076437f
C48 ctl3 ctl4 0.076437f
C49 n3 n0 0.051666f
C50 n7 ndum 0.06073f
C51 n5 ndum 0.025424f
C52 n3 n6 0.336612f
C53 inv_renketu_0/inv$1_9/VSS ctl7 0.002242f
C54 ctl5 ctl4 0.076437f
C55 out n0 1.745294f
C56 ctl6 ctl7 0.076437f
C57 n1 n0 8.476099f
C58 ctl1 dum 0.076437f
C59 n6 out 0.105055p
C60 n3 ndum 0.025424f
C61 n9 inv_renketu_0/inv$1_9/VDD 0.001148f
C62 n6 n1 0.141395f
C63 inv_renketu_0/inv$1_9/VSS ctl8 0.002242f
C64 n2 n8 0.770199f
C65 out ndum 1.640173f
C66 n1 ndum 8.161697f
C67 sample dum 0.00183f
C68 n7 n8 50.178104f
C69 n5 n8 5.60732f
C70 n2 n4 0.213181f
C71 n6 n0 0.025424f
C72 sample inv_renketu_0/inv$1_9/VDD 0.013129f
C73 inv_renketu_0/dummy_1/I n0 0.001307f
C74 n3 n8 1.46111f
C75 n7 n4 1.70387f
C76 n5 n4 27.491999f
C77 n6 ndum 0.025424f
C78 ctl6 inv_renketu_0/inv$1_9/VSS 0.002242f
C79 sample inv_renketu_0/inv$1_9/VNW 0.008949f
C80 n8 out 0.420151p
C81 n2 inv_renketu_0/inv$1_9/VDD 0.001148f
C82 n1 n8 0.285054f
C83 n3 n4 25.8929f
C84 n7 inv_renketu_0/inv$1_9/VDD 0.001148f
C85 out n4 26.32268f
C86 bootstrapped_sw_0/vbsl out 0.061234f
C87 n5 inv_renketu_0/inv$1_9/VDD 0.001148f
C88 n1 n4 0.141659f
C89 ctl9 ctl8 0.076437f
C90 n8 n0 0.097254f
C91 n9 n2 0.996653f
C92 n3 inv_renketu_0/inv$1_9/VDD 0.001148f
C93 n6 n8 11.2161f
C94 inv_renketu_0/inv$1_9/VSS ctl2 0.002242f
C95 inv_renketu_0/inv$1_9/VSS ctl4 0.002242f
C96 out inv_renketu_0/inv$1_9/VDD 0.007958f
C97 n9 n7 29.516087f
C98 n9 n5 7.399346f
C99 n1 inv_renketu_0/inv$1_9/VDD 0.001148f
C100 n8 ndum 0.097254f
C101 n0 n4 0.040502f
C102 sample inv_renketu_0/dummy_0/ZN 0.007127f
C103 n6 n4 0.614078f
C104 n3 n9 1.911224f
C105 inv_renketu_0/inv$1_9/VNW out 0.003912f
C106 inv_renketu_0/inv$1_9/VSS ctl9 0.002242f
C107 n4 ndum 0.025424f
C108 inv_renketu_0/inv$1_9/VSS dum 0.002242f
C109 n9 out 0.846163p
C110 inv_renketu_0/dummy_1/ZN vss 0.095951f
C111 inv_renketu_0/dummy_1/I vss 0.604559f
C112 inv_renketu_0/dummy_0/ZN vss 0.095951f
C113 inv_renketu_0/dummy_0/I vss 0.604559f
C114 ctl8 vss 0.863789f
C115 ctl7 vss 0.863789f
C116 ctl6 vss 0.863789f
C117 ctl5 vss 0.863789f
C118 ctl4 vss 0.863789f
C119 ctl3 vss 0.863789f
C120 ctl1 vss 0.863789f
C121 inv_renketu_0/inv$1_9/VSS vss 2.848055f
C122 inv_renketu_0/inv$1_9/VDD vss 2.113035f
C123 ctl0 vss 1.029175f
C124 inv_renketu_0/inv$1_9/VNW vss 14.066851f
C125 ctl2 vss 0.863789f
C126 ndum vss 13.878879f
C127 dum vss 1.023139f
C128 ctl9 vss 0.863789f
C129 n4 vss 39.311863f
C130 n5 vss 47.33512f
C131 n9 vss 14.292219f
C132 out vss -0.683569p
C133 n8 vss 39.909065f
C134 n7 vss 56.191708f
C135 n6 vss 52.976902f
C136 n0 vss 16.631123f
C137 n2 vss 30.111814f
C138 n1 vss 17.119806f
C139 n3 vss 33.594227f
C140 bootstrapped_sw_0/vs vss 0.065021f
C141 bootstrapped_sw_0/enb vss 1.523612f
C142 vdd vss 3.098478f
C143 sample vss 20.462025f
C144 bootstrapped_sw_0/XM4_0/w_n2712_234# vss 1.968192f
C145 bootstrapped_sw_0/vbsh vss 7.079245f
C146 bootstrapped_sw_0/vbsl vss 8.446682f
C147 in vss 0.297821f
C148 bootstrapped_sw_0/vg vss 1.1621f
.ends

.subckt inv$1$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 ZN I 0.58604f
C1 VNW VSS 0.006277f
C2 VNW ZN 0.023676f
C3 ZN VSS 0.180794f
C4 I VDD 0.074838f
C5 VNW VDD 0.082022f
C6 VSS VDD 0.029045f
C7 VNW I 0.285482f
C8 I VSS 0.091531f
C9 ZN VDD 0.271625f
C10 VSS VPW 0.296769f
C11 ZN VPW 0.099188f
C12 VDD VPW 0.238483f
C13 I VPW 0.610668f
C14 VNW VPW 1.31158f
.ends

.subckt dummy$1 VSS ZN I VDD VNW VPW
X0 VSS I ZN VPW nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 ZN I 0.58604f
C1 VNW VSS 0.011638f
C2 VNW ZN 0.026913f
C3 ZN VSS 0.180794f
C4 I VDD 0.075475f
C5 VNW VDD 0.108083f
C6 VSS VDD 0.035859f
C7 VNW I 0.291591f
C8 I VSS 0.092168f
C9 ZN VDD 0.271625f
C10 VSS VPW 0.337898f
C11 ZN VPW 0.095951f
C12 VDD VPW 0.258911f
C13 I VPW 0.604559f
C14 VNW VPW 1.53535f
.ends

.subckt inv_renketu$1 inv$1$1_7/I inv$1$1_6/ZN inv$1$1_9/ZN inv$1$1_0/I dummy$1_0/I
+ inv$1$1_10/I inv$1$1_0/ZN inv$1$1_4/I inv$1$1_6/I inv$1$1_8/ZN inv$1$1_5/ZN inv$1$1_8/I
+ inv$1$1_2/I dummy$1_0/ZN inv$1$1_9/VSS inv$1$1_9/VDD inv$1$1_2/ZN inv$1$1_1/I inv$1$1_9/I
+ inv$1$1_7/ZN inv$1$1_3/ZN inv$1$1_3/I inv$1$1_4/ZN inv$1$1_1/ZN dummy$1_1/I inv$1$1_9/VNW
+ inv$1$1_5/I inv$1$1_10/ZN VSUBS
Xinv$1$1_0 inv$1$1_9/VSS inv$1$1_0/ZN inv$1$1_0/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_1 inv$1$1_9/VSS inv$1$1_1/ZN inv$1$1_1/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_2 inv$1$1_9/VSS inv$1$1_2/ZN inv$1$1_2/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_3 inv$1$1_9/VSS inv$1$1_3/ZN inv$1$1_3/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_4 inv$1$1_9/VSS inv$1$1_4/ZN inv$1$1_4/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_5 inv$1$1_9/VSS inv$1$1_5/ZN inv$1$1_5/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_6 inv$1$1_9/VSS inv$1$1_6/ZN inv$1$1_6/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_7 inv$1$1_9/VSS inv$1$1_7/ZN inv$1$1_7/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xinv$1$1_8 inv$1$1_9/VSS inv$1$1_8/ZN inv$1$1_8/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xdummy$1_0 inv$1$1_9/VSS dummy$1_0/ZN dummy$1_0/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ dummy$1
Xinv$1$1_9 inv$1$1_9/VSS inv$1$1_9/ZN inv$1$1_9/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
Xdummy$1_1 inv$1$1_9/VSS dummy$1_1/ZN dummy$1_1/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ dummy$1
Xinv$1$1_10 inv$1$1_9/VSS inv$1$1_10/ZN inv$1$1_10/I inv$1$1_9/VDD inv$1$1_9/VNW VSUBS
+ inv$1$1
C0 inv$1$1_4/ZN inv$1$1_9/VSS 0.003829f
C1 inv$1$1_1/I inv$1$1_1/ZN 0.031424f
C2 inv$1$1_9/VNW inv$1$1_6/I 0.010403f
C3 inv$1$1_9/VNW inv$1$1_7/ZN 0.006066f
C4 inv$1$1_6/I inv$1$1_9/VDD 0.00333f
C5 inv$1$1_9/VDD inv$1$1_7/ZN 0.104396f
C6 inv$1$1_9/VNW inv$1$1_9/ZN 0.006066f
C7 inv$1$1_9/ZN inv$1$1_9/VDD 0.104396f
C8 inv$1$1_9/VSS inv$1$1_2/ZN 0.003829f
C9 inv$1$1_10/I inv$1$1_9/VNW 0.010403f
C10 inv$1$1_9/VSS inv$1$1_1/I 0.104553f
C11 inv$1$1_10/I inv$1$1_9/VDD 0.00333f
C12 inv$1$1_9/VNW inv$1$1_3/ZN 0.006066f
C13 inv$1$1_9/VSS inv$1$1_6/ZN 0.003829f
C14 inv$1$1_3/I inv$1$1_0/I 0.084161f
C15 inv$1$1_3/ZN inv$1$1_9/VDD 0.104396f
C16 inv$1$1_4/I inv$1$1_9/VNW 0.010403f
C17 inv$1$1_0/ZN inv$1$1_0/I 0.031424f
C18 inv$1$1_4/I inv$1$1_9/VDD 0.00333f
C19 inv$1$1_6/ZN inv$1$1_6/I 0.031424f
C20 inv$1$1_9/VNW inv$1$1_9/VDD -0.157887f
C21 inv$1$1_10/I inv$1$1_2/ZN 0.028928f
C22 inv$1$1_6/ZN inv$1$1_7/ZN 0.161793f
C23 inv$1$1_4/ZN inv$1$1_4/I 0.031424f
C24 inv$1$1_4/ZN inv$1$1_9/VNW 0.006066f
C25 inv$1$1_4/ZN inv$1$1_9/VDD 0.104396f
C26 inv$1$1_9/VSS inv$1$1_8/I 0.104553f
C27 inv$1$1_9/VNW inv$1$1_2/ZN 0.008692f
C28 inv$1$1_1/I inv$1$1_3/ZN 0.002086f
C29 inv$1$1_9/VDD inv$1$1_2/ZN 0.107277f
C30 inv$1$1_8/I inv$1$1_7/ZN 0.002086f
C31 inv$1$1_7/I inv$1$1_8/ZN 0.028928f
C32 dummy$1_1/I inv$1$1_2/ZN 0.003027f
C33 inv$1$1_10/ZN inv$1$1_9/I 0.028928f
C34 inv$1$1_1/I inv$1$1_4/I 0.084161f
C35 inv$1$1_1/I inv$1$1_9/VNW 0.010403f
C36 inv$1$1_9/ZN inv$1$1_8/I 0.028928f
C37 inv$1$1_9/VSS inv$1$1_0/I 0.108299f
C38 inv$1$1_1/I inv$1$1_9/VDD 0.00333f
C39 inv$1$1_9/VNW inv$1$1_6/ZN 0.006066f
C40 inv$1$1_4/ZN inv$1$1_1/I 0.028928f
C41 inv$1$1_6/ZN inv$1$1_9/VDD 0.104396f
C42 inv$1$1_9/I inv$1$1_8/ZN 0.002086f
C43 inv$1$1_9/VNW inv$1$1_8/I 0.010403f
C44 inv$1$1_2/I dummy$1_1/ZN 0.027478f
C45 inv$1$1_9/VDD inv$1$1_8/I 0.00333f
C46 inv$1$1_3/ZN inv$1$1_0/I 0.028928f
C47 inv$1$1_0/ZN dummy$1_0/I 0.023262f
C48 inv$1$1_9/VNW inv$1$1_0/I 0.011179f
C49 inv$1$1_9/VDD inv$1$1_0/I 0.00333f
C50 inv$1$1_5/I inv$1$1_5/ZN 0.031424f
C51 inv$1$1_10/ZN inv$1$1_2/I 0.002086f
C52 dummy$1_0/ZN inv$1$1_0/ZN 0.0229f
C53 inv$1$1_9/VSS inv$1$1_7/I 0.104553f
C54 inv$1$1_9/VSS inv$1$1_10/ZN 0.003829f
C55 inv$1$1_6/I inv$1$1_7/I 0.084161f
C56 inv$1$1_7/I inv$1$1_7/ZN 0.031424f
C57 dummy$1_0/ZN inv$1$1_9/VSS 0.001445f
C58 inv$1$1_10/ZN inv$1$1_9/ZN 0.161792f
C59 inv$1$1_9/VSS inv$1$1_9/I 0.104553f
C60 inv$1$1_9/VNW dummy$1_1/ZN -0.001925f
C61 inv$1$1_9/VSS inv$1$1_8/ZN 0.003829f
C62 inv$1$1_0/ZN inv$1$1_3/I 0.002086f
C63 dummy$1_1/ZN inv$1$1_9/VDD 0.010249f
C64 inv$1$1_10/I inv$1$1_10/ZN 0.031424f
C65 inv$1$1_9/VSS inv$1$1_5/ZN 0.003829f
C66 inv$1$1_9/I inv$1$1_9/ZN 0.031424f
C67 inv$1$1_1/ZN inv$1$1_3/I 0.028928f
C68 inv$1$1_7/ZN inv$1$1_8/ZN 0.161792f
C69 inv$1$1_9/VNW inv$1$1_7/I 0.010403f
C70 inv$1$1_9/ZN inv$1$1_8/ZN 0.161793f
C71 inv$1$1_5/I inv$1$1_9/VSS 0.104553f
C72 inv$1$1_9/VDD inv$1$1_7/I 0.00333f
C73 inv$1$1_5/ZN inv$1$1_6/I 0.002086f
C74 dummy$1_1/ZN inv$1$1_2/ZN 0.022956f
C75 inv$1$1_10/ZN inv$1$1_9/VNW 0.006066f
C76 inv$1$1_10/I inv$1$1_9/I 0.084161f
C77 inv$1$1_10/ZN inv$1$1_9/VDD 0.104396f
C78 inv$1$1_5/I inv$1$1_6/I 0.084161f
C79 inv$1$1_9/VSS inv$1$1_3/I 0.104553f
C80 dummy$1_0/ZN inv$1$1_9/VNW -0.002275f
C81 dummy$1_0/ZN inv$1$1_9/VDD 0.001671f
C82 inv$1$1_9/I inv$1$1_9/VNW 0.010403f
C83 inv$1$1_0/ZN inv$1$1_9/VSS 0.003829f
C84 inv$1$1_9/I inv$1$1_9/VDD 0.00333f
C85 inv$1$1_10/ZN inv$1$1_2/ZN 0.161793f
C86 inv$1$1_9/VNW inv$1$1_8/ZN 0.006066f
C87 inv$1$1_9/VDD inv$1$1_8/ZN 0.104396f
C88 inv$1$1_9/VSS inv$1$1_1/ZN 0.003829f
C89 inv$1$1_9/VSS inv$1$1_2/I 0.107646f
C90 inv$1$1_4/I inv$1$1_5/ZN 0.028928f
C91 inv$1$1_5/ZN inv$1$1_9/VNW 0.006066f
C92 inv$1$1_6/ZN inv$1$1_7/I 0.002086f
C93 inv$1$1_5/ZN inv$1$1_9/VDD 0.104396f
C94 inv$1$1_5/I inv$1$1_4/I 0.084161f
C95 inv$1$1_4/ZN inv$1$1_5/ZN 0.161793f
C96 inv$1$1_5/I inv$1$1_9/VNW 0.010403f
C97 inv$1$1_5/I inv$1$1_9/VDD 0.00333f
C98 inv$1$1_3/I inv$1$1_3/ZN 0.031424f
C99 inv$1$1_5/I inv$1$1_4/ZN 0.002086f
C100 inv$1$1_7/I inv$1$1_8/I 0.084161f
C101 inv$1$1_0/ZN inv$1$1_3/ZN 0.161792f
C102 inv$1$1_9/VNW inv$1$1_3/I 0.010403f
C103 inv$1$1_10/I inv$1$1_2/I 0.084161f
C104 inv$1$1_9/VSS inv$1$1_6/I 0.104553f
C105 inv$1$1_3/I inv$1$1_9/VDD 0.00333f
C106 inv$1$1_9/VSS inv$1$1_7/ZN 0.003829f
C107 inv$1$1_0/ZN inv$1$1_9/VNW 0.008403f
C108 inv$1$1_1/ZN inv$1$1_3/ZN 0.161793f
C109 inv$1$1_9/VSS inv$1$1_9/ZN 0.003829f
C110 inv$1$1_0/ZN inv$1$1_9/VDD 0.107658f
C111 inv$1$1_5/ZN inv$1$1_6/ZN 0.161792f
C112 inv$1$1_4/I inv$1$1_1/ZN 0.002086f
C113 inv$1$1_6/I inv$1$1_7/ZN 0.028928f
C114 inv$1$1_1/ZN inv$1$1_9/VNW 0.006066f
C115 inv$1$1_9/VNW inv$1$1_2/I 0.011789f
C116 inv$1$1_1/ZN inv$1$1_9/VDD 0.104396f
C117 inv$1$1_2/I inv$1$1_9/VDD 0.00333f
C118 inv$1$1_9/I inv$1$1_8/I 0.084161f
C119 inv$1$1_10/I inv$1$1_9/VSS 0.104553f
C120 dummy$1_0/I inv$1$1_0/I 0.017781f
C121 inv$1$1_5/I inv$1$1_6/ZN 0.028928f
C122 inv$1$1_4/ZN inv$1$1_1/ZN 0.161792f
C123 dummy$1_1/I inv$1$1_2/I 0.021288f
C124 inv$1$1_8/I inv$1$1_8/ZN 0.031424f
C125 inv$1$1_9/VSS inv$1$1_3/ZN 0.003829f
C126 inv$1$1_1/I inv$1$1_3/I 0.084161f
C127 dummy$1_0/ZN inv$1$1_0/I 0.002409f
C128 inv$1$1_9/VSS inv$1$1_4/I 0.104553f
C129 inv$1$1_10/I inv$1$1_9/ZN 0.002086f
C130 inv$1$1_9/VSS inv$1$1_9/VNW -0.005361f
C131 inv$1$1_2/I inv$1$1_2/ZN 0.031424f
C132 inv$1$1_9/VSS inv$1$1_9/VDD -0.006814f
C133 inv$1$1_10/ZN VSUBS 0.260352f
C134 inv$1$1_10/I VSUBS 0.670517f
C135 dummy$1_1/ZN VSUBS 0.095951f
C136 dummy$1_1/I VSUBS 0.604559f
C137 inv$1$1_9/ZN VSUBS 0.260352f
C138 inv$1$1_9/I VSUBS 0.670517f
C139 dummy$1_0/ZN VSUBS 0.095951f
C140 dummy$1_0/I VSUBS 0.604559f
C141 inv$1$1_8/ZN VSUBS 0.260352f
C142 inv$1$1_8/I VSUBS 0.670517f
C143 inv$1$1_7/ZN VSUBS 0.260352f
C144 inv$1$1_7/I VSUBS 0.670517f
C145 inv$1$1_6/ZN VSUBS 0.260352f
C146 inv$1$1_6/I VSUBS 0.670517f
C147 inv$1$1_5/ZN VSUBS 0.260352f
C148 inv$1$1_5/I VSUBS 0.670517f
C149 inv$1$1_4/ZN VSUBS 0.260352f
C150 inv$1$1_4/I VSUBS 0.670517f
C151 inv$1$1_3/ZN VSUBS 0.260352f
C152 inv$1$1_3/I VSUBS 0.670517f
C153 inv$1$1_9/VSS VSUBS 2.848055f
C154 inv$1$1_2/ZN VSUBS 0.398879f
C155 inv$1$1_9/VDD VSUBS 2.113035f
C156 inv$1$1_2/I VSUBS 0.741957f
C157 inv$1$1_9/VNW VSUBS 14.066851f
C158 inv$1$1_1/ZN VSUBS 0.260352f
C159 inv$1$1_1/I VSUBS 0.670517f
C160 inv$1$1_0/ZN VSUBS 0.398674f
C161 inv$1$1_0/I VSUBS 0.735921f
.ends

.subckt XMs$1 a_1030_4680# a_1030_4868# a_947_4768# a_846_4542#
X0 a_1030_4868# a_947_4768# a_1030_4680# a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_1030_4868# a_1030_4680# 0.103318f
C1 a_1030_4868# a_947_4768# 0.002993f
C2 a_1030_4680# a_947_4768# 0.002993f
C3 a_1030_4680# a_846_4542# 0.387117f
C4 a_947_4768# a_846_4542# 0.288368f
C5 a_1030_4868# a_846_4542# 0.109266f
.ends

.subckt XM3$4 a_n3152_1140# a_n3064_1048# w_n3314_932# a_n2964_1140# VSUBS
X0 a_n2964_1140# a_n3064_1048# a_n3152_1140# w_n3314_932# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 w_n3314_932# a_n3152_1140# 0.008969f
C1 a_n2964_1140# w_n3314_932# 0.009117f
C2 a_n2964_1140# a_n3152_1140# 0.103318f
C3 w_n3314_932# a_n3064_1048# 0.157732f
C4 a_n3152_1140# a_n3064_1048# 0.002993f
C5 a_n2964_1140# a_n3064_1048# 0.002993f
C6 a_n2964_1140# VSUBS 0.100353f
C7 a_n3152_1140# VSUBS 0.100353f
C8 a_n3064_1048# VSUBS 0.130702f
C9 w_n3314_932# VSUBS 1.4688f
.ends

.subckt XM2_inv$1 a_n36_120# a_n116_n100# w_n278_n310# VSUBS
X0 w_n278_n310# a_n36_120# a_n116_n100# w_n278_n310# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 w_n278_n310# a_n116_n100# 0.090564f
C1 w_n278_n310# a_n36_120# 0.138578f
C2 a_n116_n100# a_n36_120# 0.001764f
C3 a_n116_n100# VSUBS 0.043675f
C4 a_n36_120# VSUBS 0.08816f
C5 w_n278_n310# VSUBS 1.2321f
.ends

.subckt XM1_inv$1 a_n36_20# a_n254_n386# a_28_n200#
X0 a_28_n200# a_n36_20# a_n254_n386# a_n254_n386# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n36_20# a_28_n200# 0.001764f
C1 a_28_n200# a_n254_n386# 0.134177f
C2 a_n36_20# a_n254_n386# 0.22667f
.ends

.subckt inv$3 out in vdd vss
XXM2_inv$1_0 in out vdd vss XM2_inv$1
XXM1_inv$1_0 in vss out XM1_inv$1
C0 vss vdd 0.050184f
C1 vss in 0.019395f
C2 vdd in 0.034991f
C3 vss out 0.056311f
C4 vdd out 0.086562f
C5 out in 0.057341f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt XMs2$1 a_n3762_561# a_n3988_469# a_n3662_653# a_n3850_653# a_n3988_1165#
X0 a_n3662_653# a_n3762_561# a_n3850_653# a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n3662_653# a_n3762_561# 0.002993f
C1 a_n3850_653# a_n3762_561# 0.002993f
C2 a_n3662_653# a_n3850_653# 0.103318f
C3 a_n3662_653# a_n3988_469# 0.109266f
C4 a_n3850_653# a_n3988_469# 0.109266f
C5 a_n3762_561# a_n3988_469# 0.288275f
.ends

.subckt XM2$4 a_912_3686# a_811_3460# a_995_3786# a_1507_3460# a_995_3598#
X0 a_995_3786# a_912_3686# a_995_3598# a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_995_3598# a_995_3786# 0.103318f
C1 a_912_3686# a_995_3786# 0.002993f
C2 a_995_3598# a_912_3686# 0.002993f
C3 a_995_3598# a_811_3460# 0.109266f
C4 a_912_3686# a_811_3460# 0.288275f
C5 a_995_3786# a_811_3460# 0.109266f
.ends

.subckt cap_mim_2p0fF_8JNR63$1 m4_n3440_n548# m4_n3800_n668# VSUBS
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0_m4m5_noshield c_width=8u c_length=8u
C0 m4_n3800_n668# m4_n3440_n548# 0.646322f
C1 m4_n3440_n548# VSUBS 1.17298f
C2 m4_n3800_n668# VSUBS 1.64833f
.ends

.subckt sw_cap_unit$1 in out VSUBS
Xcap_mim_2p0fF_8JNR63_0 out in VSUBS cap_mim_2p0fF_8JNR63$1
C0 out VSUBS 1.17298f
C1 in VSUBS 1.64833f
.ends

.subckt sw_cap$1 out in VSUBS
Xsw_cap_unit$1_0 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_1 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_2 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_3 in out VSUBS sw_cap_unit$1
Xsw_cap_unit$1_4 in out VSUBS sw_cap_unit$1
C0 in out 2.231591f
C1 out VSUBS 6.064711f
C2 in VSUBS 7.39096f
.ends

.subckt XMs1$1 a_n2529_n616# a_n2717_n616# a_n2629_n699# a_n2855_n800#
X0 a_n2529_n616# a_n2629_n699# a_n2717_n616# a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n2629_n699# a_n2529_n616# 0.002993f
C1 a_n2717_n616# a_n2629_n699# 0.002993f
C2 a_n2717_n616# a_n2529_n616# 0.103318f
C3 a_n2529_n616# a_n2855_n800# 0.109266f
C4 a_n2717_n616# a_n2855_n800# 0.177295f
C5 a_n2629_n699# a_n2855_n800# 0.288368f
.ends

.subckt XM1$4 a_912_4129# a_995_4229# a_811_3903# a_1507_3903# a_995_4041#
X0 a_995_4229# a_912_4129# a_995_4041# a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_995_4041# a_995_4229# 0.103318f
C1 a_995_4229# a_912_4129# 0.002993f
C2 a_995_4041# a_912_4129# 0.002993f
C3 a_995_4041# a_811_3903# 0.109266f
C4 a_912_4129# a_811_3903# 0.288275f
C5 a_995_4229# a_811_3903# 0.109266f
.ends

.subckt XM4$4 a_n2550_442# a_n2362_442# w_n2712_234# a_n2462_359# VSUBS
X0 a_n2362_442# a_n2462_359# a_n2550_442# w_n2712_234# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 a_n2362_442# a_n2462_359# 0.002993f
C1 w_n2712_234# a_n2550_442# 0.058295f
C2 a_n2462_359# w_n2712_234# 0.173648f
C3 a_n2462_359# a_n2550_442# 0.002993f
C4 a_n2362_442# w_n2712_234# 0.008969f
C5 a_n2362_442# a_n2550_442# 0.103318f
C6 a_n2362_442# VSUBS 0.100353f
C7 a_n2550_442# VSUBS 0.119847f
C8 a_n2462_359# VSUBS 0.147064f
C9 w_n2712_234# VSUBS 1.4688f
.ends

.subckt bootstrapped_sw$1 in vdd vss en enb out vs vg vbsl vbsh
XXMs$1_0 out in vg vss XMs$1
XXM3$4_0 vbsh vg XM4$4_0/w_n2712_234# vdd vss XM3$4
Xinv$3_0 enb en vdd vss inv$3
XXMs2$1_0 enb vss vss vs vss XMs2$1
XXM2$4_0 enb vss vss vss vbsl XM2$4
Xsw_cap$1_0 vbsh vbsl vss sw_cap$1
XXMs1$1_0 vs vg vdd vss XMs1$1
XXM1$4_0 vg vbsl vss vss in XM1$4
XXM4$4_0 vg vbsh XM4$4_0/w_n2712_234# enb vss XM4$4
C0 enb XM4$4_0/w_n2712_234# 0.041524f
C1 vdd enb 0.448382f
C2 en enb 0.029269f
C3 vbsl vg 0.046114f
C4 vbsl out 0.058082f
C5 enb vs 0.00376f
C6 vg XM4$4_0/w_n2712_234# 0.080093f
C7 out XM4$4_0/w_n2712_234# 0.005706f
C8 vdd vg 0.447812f
C9 vbsl vbsh 0.025766f
C10 vdd out 0.017908f
C11 vg vs 0.01049f
C12 vbsh XM4$4_0/w_n2712_234# 0.101815f
C13 vdd vbsh 0.168905f
C14 in vg 0.075595f
C15 vbsl XM4$4_0/w_n2712_234# 0.009881f
C16 vg enb 0.612109f
C17 vbsl vdd 0.005409f
C18 in vbsh 0.008752f
C19 vbsl vs 0.001422f
C20 vdd XM4$4_0/w_n2712_234# 0.079362f
C21 enb vbsh 0.052707f
C22 vdd en 0.065092f
C23 out vg 0.04429f
C24 vg vbsh 0.144325f
C25 vbsl in 0.299565f
C26 out vbsh 0.100712f
C27 vbsl enb 0.017274f
C28 out vss 1.088543f
C29 XM4$4_0/w_n2712_234# vss 1.968192f
C30 in vss 0.308876f
C31 vbsh vss 7.100617f
C32 vbsl vss 8.368301f
C33 enb vss 1.595319f
C34 vs vss 0.072259f
C35 vdd vss 3.106074f
C36 en vss 0.642295f
C37 vg vss 1.218873f
.ends

.subckt dacn in dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl0 out ndum n1
+ n2 n3 n4 n5 n6 n7 n8 n9 n0 sample vdd bootstrapped_sw$1_0/vbsl bootstrapped_sw$1_0/vbsh
+ vss
Xinv_renketu$1_0 ctl6 n5 n8 dum inv_renketu$1_0/dummy$1_0/I ctl9 ndum ctl3 ctl5 n7
+ n4 ctl7 ctl0 inv_renketu$1_0/dummy$1_0/ZN inv_renketu$1_0/inv$1$1_9/VSS inv_renketu$1_0/inv$1$1_9/VDD
+ n0 ctl2 ctl8 n6 n1 ctl1 n3 n2 inv_renketu$1_0/dummy$1_1/I inv_renketu$1_0/inv$1$1_9/VNW
+ ctl4 n9 vss inv_renketu$1
Xbootstrapped_sw$1_0 in vdd vss sample bootstrapped_sw$1_0/enb out bootstrapped_sw$1_0/vs
+ bootstrapped_sw$1_0/vg bootstrapped_sw$1_0/vbsl bootstrapped_sw$1_0/vbsh bootstrapped_sw$1
C0 n8 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C1 ctl1 dum 0.076437f
C2 out inv_renketu$1_0/inv$1$1_9/VDD 0.007958f
C3 ctl7 ctl8 0.076437f
C4 n7 n1 0.212006f
C5 n9 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C6 inv_renketu$1_0/inv$1$1_9/VDD n0 0.008798f
C7 ndum sample 0.046157f
C8 n4 n1 0.141659f
C9 ndum n1 8.161697f
C10 inv_renketu$1_0/inv$1$1_9/VSS ctl0 0.002242f
C11 ctl2 ctl3 0.076437f
C12 n5 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C13 inv_renketu$1_0/dummy$1_0/ZN sample 0.007127f
C14 out bootstrapped_sw$1_0/vbsh 0.137967f
C15 n8 n3 1.46111f
C16 n2 n1 16.604633f
C17 inv_renketu$1_0/inv$1$1_9/VSS ctl2 0.002242f
C18 inv_renketu$1_0/inv$1$1_9/VSS ctl8 0.002242f
C19 out n3 13.201303f
C20 n9 n3 1.911224f
C21 n6 n1 0.141395f
C22 n3 n0 0.051666f
C23 n7 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C24 n5 n3 0.346757f
C25 n4 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C26 ctl0 ctl9 0.076437f
C27 ndum inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C28 out n8 0.420151p
C29 n9 n8 87.102684f
C30 n8 n0 0.097254f
C31 out n9 0.846163p
C32 out n0 1.745294f
C33 ctl8 ctl9 0.076437f
C34 n9 n0 0.184985f
C35 n2 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C36 ctl4 ctl3 0.076437f
C37 inv_renketu$1_0/inv$1$1_9/VNW sample 0.008949f
C38 n5 n8 5.60732f
C39 n7 n3 0.891504f
C40 n6 inv_renketu$1_0/inv$1$1_9/VDD 0.001148f
C41 out n5 52.565514f
C42 n4 n3 25.8929f
C43 n5 n9 7.399346f
C44 inv_renketu$1_0/inv$1$1_9/VSS ctl4 0.002242f
C45 ndum n3 0.025424f
C46 inv_renketu$1_0/inv$1$1_9/VSS ctl7 0.002242f
C47 ctl4 ctl5 0.076437f
C48 n5 n0 0.025424f
C49 inv_renketu$1_0/inv$1$1_9/VSS sample 0.011446f
C50 ctl7 ctl6 0.076437f
C51 n2 n3 22.840685f
C52 inv_renketu$1_0/inv$1$1_9/VSS ctl3 0.002242f
C53 n7 n8 50.178104f
C54 out bootstrapped_sw$1_0/vbsl 0.061234f
C55 n4 n8 2.84323f
C56 out n7 0.210031p
C57 n6 n3 0.336612f
C58 n7 n9 29.516087f
C59 ndum n8 0.097254f
C60 out n4 26.32268f
C61 n7 n0 0.06073f
C62 n4 n9 3.740573f
C63 out ndum 1.640173f
C64 inv_renketu$1_0/inv$1$1_9/VSS ctl5 0.002242f
C65 n4 n0 0.040502f
C66 ndum n9 0.127951f
C67 inv_renketu$1_0/dummy$1_1/I n0 0.001307f
C68 n5 n7 3.36878f
C69 sample dum 0.00183f
C70 n2 n8 0.770199f
C71 ctl2 ctl1 0.076437f
C72 inv_renketu$1_0/inv$1$1_9/VSS ctl6 0.002242f
C73 n5 n4 27.491999f
C74 ctl5 ctl6 0.076437f
C75 out n2 6.640605f
C76 inv_renketu$1_0/inv$1$1_9/VDD sample 0.013129f
C77 ndum n5 0.025424f
C78 n8 n6 11.2161f
C79 n2 n9 0.996653f
C80 inv_renketu$1_0/inv$1$1_9/VDD n1 0.001148f
C81 n2 n0 0.099287f
C82 out n6 0.105055p
C83 inv_renketu$1_0/inv$1$1_9/VSS dum 0.002242f
C84 n9 n6 14.716789f
C85 n6 n0 0.025424f
C86 n2 n5 0.208084f
C87 inv_renketu$1_0/inv$1$1_9/VSS ctl9 0.002242f
C88 n5 n6 28.589401f
C89 n7 n4 1.70387f
C90 ndum n7 0.06073f
C91 ndum n4 0.025424f
C92 inv_renketu$1_0/dummy$1_0/I sample 0.008276f
C93 n3 n1 0.144232f
C94 n2 n7 0.485327f
C95 n2 n4 0.213181f
C96 out inv_renketu$1_0/inv$1$1_9/VNW 0.003912f
C97 n7 n6 34.326103f
C98 n2 ndum 0.041162f
C99 inv_renketu$1_0/inv$1$1_9/VNW n0 0.002542f
C100 n4 n6 0.614078f
C101 ndum n6 0.025424f
C102 n8 n1 0.285054f
C103 out n1 3.367623f
C104 n9 n1 0.349226f
C105 n1 n0 8.476099f
C106 n2 n6 0.207962f
C107 inv_renketu$1_0/inv$1$1_9/VDD n3 0.001148f
C108 inv_renketu$1_0/inv$1$1_9/VSS ctl1 0.002242f
C109 n5 n1 0.141538f
C110 bootstrapped_sw$1_0/XM4$4_0/w_n2712_234# vss 1.968192f
C111 in vss 0.297821f
C112 bootstrapped_sw$1_0/vbsh vss 7.079245f
C113 bootstrapped_sw$1_0/vbsl vss 8.446682f
C114 bootstrapped_sw$1_0/enb vss 1.523612f
C115 bootstrapped_sw$1_0/vs vss 0.065021f
C116 vdd vss 3.098478f
C117 sample vss 20.462025f
C118 bootstrapped_sw$1_0/vg vss 1.1621f
C119 ctl9 vss 0.863789f
C120 inv_renketu$1_0/dummy$1_1/ZN vss 0.095951f
C121 inv_renketu$1_0/dummy$1_1/I vss 0.604559f
C122 ctl8 vss 0.863789f
C123 inv_renketu$1_0/dummy$1_0/ZN vss 0.095951f
C124 inv_renketu$1_0/dummy$1_0/I vss 0.604559f
C125 ctl7 vss 0.863789f
C126 ctl6 vss 0.863789f
C127 ctl5 vss 0.863789f
C128 ctl4 vss 0.863789f
C129 ctl3 vss 0.863789f
C130 ctl1 vss 0.863789f
C131 inv_renketu$1_0/inv$1$1_9/VSS vss 2.848055f
C132 inv_renketu$1_0/inv$1$1_9/VDD vss 2.113035f
C133 ctl0 vss 1.029175f
C134 inv_renketu$1_0/inv$1$1_9/VNW vss 14.066851f
C135 ctl2 vss 0.863789f
C136 ndum vss 13.878879f
C137 dum vss 1.023139f
C138 n0 vss 16.631123f
C139 n1 vss 17.119806f
C140 n4 vss 39.311863f
C141 n5 vss 47.33512f
C142 n2 vss 30.111814f
C143 n3 vss 33.594227f
C144 n9 vss 14.292219f
C145 out vss -0.683569p
C146 n8 vss 39.909065f
C147 n7 vss 56.191708f
C148 n6 vss 52.976902f
.ends

.subckt XMinn a_719_n1284# a_937_n880# a_857_n1100# a_719_n788# a_1001_n1100#
X0 a_1001_n1100# a_937_n880# a_857_n1100# a_719_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_1001_n1100# a_937_n880# 0.001764f
C1 a_937_n880# a_857_n1100# 0.001764f
C2 a_1001_n1100# a_857_n1100# 0.06854f
C3 a_1001_n1100# a_719_n1284# 0.057707f
C4 a_857_n1100# a_719_n1284# 0.057707f
C5 a_937_n880# a_719_n1284# 0.21851f
.ends

.subckt XM1$3 a_n1416_1000# a_n1336_908# a_n1272_1000# w_n1578_790# VSUBS
X0 a_n1272_1000# a_n1336_908# a_n1416_1000# w_n1578_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n1416_1000# w_n1578_790# 0.022441f
C1 a_n1272_1000# a_n1336_908# 0.001764f
C2 a_n1336_908# a_n1416_1000# 0.001764f
C3 a_n1272_1000# a_n1416_1000# 0.06854f
C4 a_n1336_908# w_n1578_790# 0.132558f
C5 a_n1272_1000# w_n1578_790# 0.021497f
C6 a_n1272_1000# VSUBS 0.043675f
C7 a_n1416_1000# VSUBS 0.043675f
C8 a_n1336_908# VSUBS 0.08816f
C9 w_n1578_790# VSUBS 1.17557f
.ends

.subckt XM3$2 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n496_n791# a_n336_n791# 0.131547f
C1 a_n240_n571# a_n176_n791# 0.005902f
C2 a_n640_n791# a_n496_n791# 0.131547f
C3 a_n400_n571# a_n336_n791# 0.005902f
C4 a_n640_n791# a_n336_n791# 0.040052f
C5 a_n176_n791# a_n16_n791# 0.131547f
C6 a_n400_n571# a_n240_n571# 0.043712f
C7 a_n240_n571# a_n336_n791# 0.005902f
C8 a_n496_n791# a_n560_n571# 0.005902f
C9 a_n80_n571# a_n240_n571# 0.043712f
C10 a_n400_n571# a_n560_n571# 0.043712f
C11 a_n176_n791# a_n336_n791# 0.131547f
C12 a_n16_n791# a_n336_n791# 0.040052f
C13 a_n640_n791# a_n560_n571# 0.005902f
C14 a_n80_n571# a_n176_n791# 0.005902f
C15 a_n496_n791# a_n400_n571# 0.005902f
C16 a_n80_n571# a_n16_n791# 0.005902f
C17 a_n16_n791# a_n778_n975# 0.182857f
C18 a_n176_n791# a_n778_n975# 0.043869f
C19 a_n336_n791# a_n778_n975# 0.097543f
C20 a_n496_n791# a_n778_n975# 0.043869f
C21 a_n640_n791# a_n778_n975# 0.277121f
C22 a_n80_n571# a_n778_n975# 0.191307f
C23 a_n240_n571# a_n778_n975# 0.164084f
C24 a_n400_n571# a_n778_n975# 0.16416f
C25 a_n560_n571# a_n778_n975# 0.198604f
.ends

.subckt XM2$2 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n157_n712# a_n237_n932# 0.005902f
C1 a_3_n712# a_n157_n712# 0.043712f
C2 a_n93_n932# a_n237_n932# 0.131547f
C3 a_n93_n932# a_3_n712# 0.005902f
C4 a_67_n932# a_n93_n932# 0.131547f
C5 a_n93_n932# a_n157_n712# 0.005902f
C6 a_67_n932# a_n237_n932# 0.040052f
C7 a_67_n932# a_3_n712# 0.005902f
C8 a_67_n932# a_n375_n1116# 0.182823f
C9 a_n93_n932# a_n375_n1116# 0.043869f
C10 a_n237_n932# a_n375_n1116# 0.182332f
C11 a_3_n712# a_n375_n1116# 0.191252f
C12 a_n157_n712# a_n375_n1116# 0.191252f
.ends

.subckt XM0$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n266_803# a_n202_583# 0.005902f
C1 a_n346_583# a_n266_803# 0.011845f
C2 a_n346_583# a_n202_583# 0.14243f
C3 a_n202_583# a_n484_399# 0.098801f
C4 a_n346_583# a_n484_399# 0.215099f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM1$2 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n266_803# a_n202_583# 0.011845f
C1 a_n346_583# a_n266_803# 0.001764f
C2 a_n346_583# a_n202_583# 0.075352f
C3 a_n202_583# a_n484_399# 0.24117f
C4 a_n346_583# a_n484_399# 0.057381f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM4$2 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_1674_n916# a_1834_n916# 0.131547f
C1 a_2090_n696# a_2250_n696# 0.043712f
C2 a_1610_n696# a_1450_n696# 0.043712f
C3 a_2250_n696# a_2314_n916# 0.005902f
C4 a_1610_n696# a_1514_n916# 0.005902f
C5 a_1930_n696# a_1834_n916# 0.005902f
C6 a_2090_n696# a_1994_n916# 0.005902f
C7 a_2410_n696# a_2250_n696# 0.043712f
C8 a_1994_n916# a_2314_n916# 0.040052f
C9 a_1210_n916# a_1354_n916# 0.131547f
C10 a_1354_n916# a_1290_n696# 0.005902f
C11 a_1674_n916# a_1770_n696# 0.005902f
C12 a_1450_n696# a_1354_n916# 0.005902f
C13 a_1610_n696# a_1674_n916# 0.005902f
C14 a_2410_n696# a_2314_n916# 0.005902f
C15 a_1354_n916# a_1514_n916# 0.131547f
C16 a_1930_n696# a_1770_n696# 0.043712f
C17 a_2154_n916# a_2250_n696# 0.005902f
C18 a_1674_n916# a_1354_n916# 0.040052f
C19 a_2090_n696# a_2154_n916# 0.005902f
C20 a_1210_n916# a_1290_n696# 0.005902f
C21 a_1450_n696# a_1290_n696# 0.043712f
C22 a_2154_n916# a_2314_n916# 0.131547f
C23 a_2474_n916# a_2314_n916# 0.131547f
C24 a_2154_n916# a_1994_n916# 0.131547f
C25 a_1770_n696# a_1834_n916# 0.005902f
C26 a_1450_n696# a_1514_n916# 0.005902f
C27 a_1674_n916# a_1994_n916# 0.040052f
C28 a_2474_n916# a_2410_n696# 0.005902f
C29 a_2090_n696# a_1930_n696# 0.043712f
C30 a_1930_n696# a_1994_n916# 0.005902f
C31 a_1674_n916# a_1514_n916# 0.131547f
C32 a_1610_n696# a_1770_n696# 0.043712f
C33 a_1994_n916# a_1834_n916# 0.131547f
C34 a_2474_n916# a_1072_n1100# 0.19427f
C35 a_2314_n916# a_1072_n1100# 0.126868f
C36 a_2154_n916# a_1072_n1100# 0.043869f
C37 a_1994_n916# a_1072_n1100# 0.097543f
C38 a_1834_n916# a_1072_n1100# 0.043869f
C39 a_1674_n916# a_1072_n1100# 0.097543f
C40 a_1514_n916# a_1072_n1100# 0.043869f
C41 a_1354_n916# a_1072_n1100# 0.126868f
C42 a_1210_n916# a_1072_n1100# 0.099481f
C43 a_2410_n696# a_1072_n1100# 0.198604f
C44 a_2250_n696# a_1072_n1100# 0.16416f
C45 a_2090_n696# a_1072_n1100# 0.164084f
C46 a_1930_n696# a_1072_n1100# 0.164049f
C47 a_1770_n696# a_1072_n1100# 0.164031f
C48 a_1610_n696# a_1072_n1100# 0.16402f
C49 a_1450_n696# a_1072_n1100# 0.164014f
C50 a_1290_n696# a_1072_n1100# 0.191268f
.ends

.subckt trim_switch$1 m1_n149_n1117# m1_n1378_n1819# m1_711_n1117# m1_n2738_n1819#
+ m1_n447_n1117# m1_n2669_n1117# XM1$2_0/a_n202_583# XM0$1_0/a_n346_583# m1_n1309_n1117#
+ m1_802_n1819# VSUBS
XXM3$2_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$2
XXM2$2_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$2
XXM0$1_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0$1_0/a_n346_583# XM0$1
XXM1$2_0 VSUBS XM1$2_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$2
XXM4$2_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$2
C0 m1_n447_n1117# m1_n1309_n1117# 0.041018f
C1 m1_711_n1117# m1_802_n1819# 0.272119f
C2 XM0$1_0/a_n346_583# XM1$2_0/a_n202_583# 0.027386f
C3 m1_n1378_n1819# m1_n1309_n1117# 0.014034f
C4 m1_n2669_n1117# m1_n1309_n1117# 0.027949f
C5 m1_n447_n1117# XM0$1_0/a_n346_583# 0.07096f
C6 m1_n1378_n1819# m1_n2738_n1819# 0.040124f
C7 m1_n2669_n1117# m1_n2738_n1819# 0.092062f
C8 m1_n149_n1117# XM1$2_0/a_n202_583# 0.07096f
C9 m1_n1378_n1819# XM0$1_0/a_n346_583# 0.039382f
C10 m1_n149_n1117# m1_711_n1117# 0.02663f
C11 XM1$2_0/a_n202_583# m1_802_n1819# 0.00859f
C12 m1_n149_n1117# m1_n447_n1117# 0.123582f
C13 m1_802_n1819# VSUBS 1.278621f
C14 m1_711_n1117# VSUBS 1.959711f
C15 XM1$2_0/a_n202_583# VSUBS 0.42776f
C16 m1_n149_n1117# VSUBS 0.407201f
C17 XM0$1_0/a_n346_583# VSUBS 0.314559f
C18 m1_n447_n1117# VSUBS 0.388025f
C19 m1_n1378_n1819# VSUBS 0.604021f
C20 m1_n1309_n1117# VSUBS 0.637566f
C21 m1_n2738_n1819# VSUBS 1.12292f
C22 m1_n2669_n1117# VSUBS 1.128649f
.ends

.subckt trim drain d_4 d_1 d_0 d_2 d_3 n1 n0 n3 n4 n2 VSUBS
Xtrim_switch$1_0 d_1 n2 d_4 n3 d_0 d_3 n1 n0 d_2 n4 VSUBS trim_switch$1
C0 n3 n0 0.087807f
C1 n4 n3 1.600479f
C2 n3 n1 0.087807f
C3 n2 d_0 0.002632f
C4 n1 d_1 0.003099f
C5 n2 d_4 0.00312f
C6 drain n2 3.213024f
C7 drain n3 6.427485f
C8 n2 n3 0.58337f
C9 n2 d_1 0.003137f
C10 n4 n0 0.166348f
C11 n1 n0 0.520979f
C12 n4 n1 0.169398f
C13 n0 d_0 0.004139f
C14 drain n0 1.60623f
C15 n2 n0 0.103368f
C16 drain n4 12.877382f
C17 n4 n2 0.596682f
C18 drain n1 1.60623f
C19 n2 n1 0.081094f
C20 n4 VSUBS 4.367046f
C21 drain VSUBS -5.906306f
C22 n3 VSUBS 3.463842f
C23 n2 VSUBS 2.03715f
C24 n0 VSUBS 0.689164f
C25 n1 VSUBS 0.727243f
C26 d_4 VSUBS 1.64786f
C27 d_1 VSUBS 0.345562f
C28 d_0 VSUBS 0.33412f
C29 d_2 VSUBS 0.513348f
C30 d_3 VSUBS 0.927186f
.ends

.subckt XMl4 a_44_908# a_108_1000# a_n36_1000# w_n198_790# VSUBS
X0 a_108_1000# a_44_908# a_n36_1000# w_n198_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n36_1000# a_44_908# 0.001764f
C1 a_44_908# w_n198_790# 0.131025f
C2 a_n36_1000# w_n198_790# 0.008358f
C3 a_44_908# a_108_1000# 0.001764f
C4 a_n36_1000# a_108_1000# 0.06854f
C5 a_108_1000# w_n198_790# 0.010275f
C6 a_108_1000# VSUBS 0.047486f
C7 a_n36_1000# VSUBS 0.049403f
C8 a_44_908# VSUBS 0.087507f
C9 w_n198_790# VSUBS 1.54752f
.ends

.subckt XM4$3 a_1264_908# a_1328_1000# w_1022_790# a_1184_1000# VSUBS
X0 a_1328_1000# a_1264_908# a_1184_1000# w_1022_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_1184_1000# a_1264_908# 0.001764f
C1 a_1264_908# w_1022_790# 0.132558f
C2 a_1184_1000# w_1022_790# 0.021497f
C3 a_1264_908# a_1328_1000# 0.001764f
C4 a_1184_1000# a_1328_1000# 0.06854f
C5 a_1328_1000# w_1022_790# 0.022441f
C6 a_1328_1000# VSUBS 0.043675f
C7 a_1184_1000# VSUBS 0.043675f
C8 a_1264_908# VSUBS 0.08816f
C9 w_1022_790# VSUBS 1.17557f
.ends

.subckt XMl2 a_33_n1100# a_n111_n1100# a_n31_n880# a_n249_n1284#
X0 a_33_n1100# a_n31_n880# a_n111_n1100# a_n249_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_33_n1100# a_n111_n1100# 0.06854f
C1 a_n111_n1100# a_n31_n880# 0.001764f
C2 a_33_n1100# a_n31_n880# 0.001764f
C3 a_33_n1100# a_n249_n1284# 0.066395f
C4 a_n111_n1100# a_n249_n1284# 0.057707f
C5 a_n31_n880# a_n249_n1284# 0.218606f
.ends

.subckt XM3$3 a_n71_n882# a_73_n882# a_9_n662# w_n509_n1092# VSUBS
X0 a_73_n882# a_9_n662# a_n71_n882# w_n509_n1092# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n71_n882# a_9_n662# 0.001764f
C1 a_9_n662# w_n509_n1092# 0.131025f
C2 a_n71_n882# w_n509_n1092# 0.010275f
C3 a_9_n662# a_73_n882# 0.001764f
C4 a_n71_n882# a_73_n882# 0.06854f
C5 a_73_n882# w_n509_n1092# 0.008358f
C6 a_73_n882# VSUBS 0.049403f
C7 a_n71_n882# VSUBS 0.047486f
C8 a_9_n662# VSUBS 0.087507f
C9 w_n509_n1092# VSUBS 1.54752f
.ends

.subckt XMdiff a_721_n1097# a_817_n1189# a_439_n1281# a_657_n1189# a_577_n1097# a_881_n1097#
X0 a_721_n1097# a_657_n1189# a_577_n1097# a_439_n1281# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_881_n1097# a_817_n1189# a_721_n1097# a_439_n1281# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_881_n1097# a_817_n1189# 0.001764f
C1 a_881_n1097# a_721_n1097# 0.06854f
C2 a_817_n1189# a_657_n1189# 0.043712f
C3 a_577_n1097# a_657_n1189# 0.001764f
C4 a_817_n1189# a_721_n1097# 0.001764f
C5 a_577_n1097# a_721_n1097# 0.06854f
C6 a_721_n1097# a_657_n1189# 0.001764f
C7 a_881_n1097# a_439_n1281# 0.115307f
C8 a_721_n1097# a_439_n1281# 0.02923f
C9 a_577_n1097# a_439_n1281# 0.115307f
C10 a_817_n1189# a_439_n1281# 0.191347f
C11 a_657_n1189# a_439_n1281# 0.191347f
.ends

.subckt XMl3 a_n116_908# w_n634_790# a_n196_1000# a_n52_1000# VSUBS
X0 a_n52_1000# a_n116_908# a_n196_1000# w_n634_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n196_1000# a_n116_908# 0.001764f
C1 a_n116_908# w_n634_790# 0.139286f
C2 a_n196_1000# w_n634_790# 0.024248f
C3 a_n116_908# a_n52_1000# 0.001764f
C4 a_n196_1000# a_n52_1000# 0.06854f
C5 a_n52_1000# w_n634_790# 0.021497f
C6 a_n52_1000# VSUBS 0.043675f
C7 a_n196_1000# VSUBS 0.041759f
C8 a_n116_908# VSUBS 0.081314f
C9 w_n634_790# VSUBS 1.68331f
.ends

.subckt XM4$1 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_1354_n916# a_1290_n696# 0.005902f
C1 a_1674_n916# a_1994_n916# 0.040052f
C2 a_2090_n696# a_2154_n916# 0.005902f
C3 a_2090_n696# a_1930_n696# 0.043712f
C4 a_2090_n696# a_1994_n916# 0.005902f
C5 a_1930_n696# a_1834_n916# 0.005902f
C6 a_1994_n916# a_1834_n916# 0.131547f
C7 a_2314_n916# a_2250_n696# 0.005902f
C8 a_1930_n696# a_1770_n696# 0.043712f
C9 a_2154_n916# a_2250_n696# 0.005902f
C10 a_2154_n916# a_2314_n916# 0.131547f
C11 a_1994_n916# a_2314_n916# 0.040052f
C12 a_1514_n916# a_1450_n696# 0.005902f
C13 a_2154_n916# a_1994_n916# 0.131547f
C14 a_1514_n916# a_1674_n916# 0.131547f
C15 a_1210_n916# a_1290_n696# 0.005902f
C16 a_1610_n696# a_1514_n916# 0.005902f
C17 a_1610_n696# a_1450_n696# 0.043712f
C18 a_1930_n696# a_1994_n916# 0.005902f
C19 a_2314_n916# a_2474_n916# 0.131547f
C20 a_2410_n696# a_2250_n696# 0.043712f
C21 a_1610_n696# a_1674_n916# 0.005902f
C22 a_1450_n696# a_1290_n696# 0.043712f
C23 a_2410_n696# a_2314_n916# 0.005902f
C24 a_1674_n916# a_1834_n916# 0.131547f
C25 a_1210_n916# a_1354_n916# 0.131547f
C26 a_1674_n916# a_1770_n696# 0.005902f
C27 a_1610_n696# a_1770_n696# 0.043712f
C28 a_1354_n916# a_1514_n916# 0.131547f
C29 a_1354_n916# a_1450_n696# 0.005902f
C30 a_2410_n696# a_2474_n916# 0.005902f
C31 a_1834_n916# a_1770_n696# 0.005902f
C32 a_1354_n916# a_1674_n916# 0.040052f
C33 a_2090_n696# a_2250_n696# 0.043712f
C34 a_2474_n916# a_1072_n1100# 0.19427f
C35 a_2314_n916# a_1072_n1100# 0.126868f
C36 a_2154_n916# a_1072_n1100# 0.043869f
C37 a_1994_n916# a_1072_n1100# 0.097543f
C38 a_1834_n916# a_1072_n1100# 0.043869f
C39 a_1674_n916# a_1072_n1100# 0.097543f
C40 a_1514_n916# a_1072_n1100# 0.043869f
C41 a_1354_n916# a_1072_n1100# 0.126868f
C42 a_1210_n916# a_1072_n1100# 0.099481f
C43 a_2410_n696# a_1072_n1100# 0.198604f
C44 a_2250_n696# a_1072_n1100# 0.16416f
C45 a_2090_n696# a_1072_n1100# 0.164084f
C46 a_1930_n696# a_1072_n1100# 0.164049f
C47 a_1770_n696# a_1072_n1100# 0.164031f
C48 a_1610_n696# a_1072_n1100# 0.16402f
C49 a_1450_n696# a_1072_n1100# 0.164014f
C50 a_1290_n696# a_1072_n1100# 0.191268f
.ends

.subckt XM2$1$1 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n237_n932# a_n93_n932# 0.131547f
C1 a_3_n712# a_67_n932# 0.005902f
C2 a_n93_n932# a_67_n932# 0.131547f
C3 a_3_n712# a_n157_n712# 0.043712f
C4 a_n157_n712# a_n93_n932# 0.005902f
C5 a_n237_n932# a_67_n932# 0.040052f
C6 a_3_n712# a_n93_n932# 0.005902f
C7 a_n237_n932# a_n157_n712# 0.005902f
C8 a_67_n932# a_n375_n1116# 0.182823f
C9 a_n93_n932# a_n375_n1116# 0.043869f
C10 a_n237_n932# a_n375_n1116# 0.182332f
C11 a_3_n712# a_n375_n1116# 0.191252f
C12 a_n157_n712# a_n375_n1116# 0.191252f
.ends

.subckt XM1$1$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n202_583# a_n346_583# 0.075352f
C1 a_n346_583# a_n266_803# 0.001764f
C2 a_n202_583# a_n266_803# 0.011845f
C3 a_n202_583# a_n484_399# 0.24117f
C4 a_n346_583# a_n484_399# 0.057381f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM3$1 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n240_n571# a_n176_n791# 0.005902f
C1 a_n80_n571# a_n240_n571# 0.043712f
C2 a_n176_n791# a_n336_n791# 0.131547f
C3 a_n16_n791# a_n336_n791# 0.040052f
C4 a_n400_n571# a_n496_n791# 0.005902f
C5 a_n16_n791# a_n176_n791# 0.131547f
C6 a_n80_n571# a_n176_n791# 0.005902f
C7 a_n80_n571# a_n16_n791# 0.005902f
C8 a_n496_n791# a_n560_n571# 0.005902f
C9 a_n640_n791# a_n496_n791# 0.131547f
C10 a_n496_n791# a_n336_n791# 0.131547f
C11 a_n240_n571# a_n400_n571# 0.043712f
C12 a_n400_n571# a_n560_n571# 0.043712f
C13 a_n640_n791# a_n560_n571# 0.005902f
C14 a_n400_n571# a_n336_n791# 0.005902f
C15 a_n240_n571# a_n336_n791# 0.005902f
C16 a_n640_n791# a_n336_n791# 0.040052f
C17 a_n16_n791# a_n778_n975# 0.182857f
C18 a_n176_n791# a_n778_n975# 0.043869f
C19 a_n336_n791# a_n778_n975# 0.097543f
C20 a_n496_n791# a_n778_n975# 0.043869f
C21 a_n640_n791# a_n778_n975# 0.277121f
C22 a_n80_n571# a_n778_n975# 0.191307f
C23 a_n240_n571# a_n778_n975# 0.164084f
C24 a_n400_n571# a_n778_n975# 0.16416f
C25 a_n560_n571# a_n778_n975# 0.198604f
.ends

.subckt XM0 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n346_583# a_n202_583# 0.14243f
C1 a_n346_583# a_n266_803# 0.011845f
C2 a_n266_803# a_n202_583# 0.005902f
C3 a_n202_583# a_n484_399# 0.098801f
C4 a_n346_583# a_n484_399# 0.215099f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt trim_switch m1_n149_n1117# XM0_0/a_n346_583# m1_711_n1117# m1_n447_n1117#
+ m1_n2669_n1117# m1_n1378_n1819# m1_802_n1819# m1_n1309_n1117# XM1$1$1_0/a_n202_583#
+ m1_n2738_n1819# VSUBS
XXM4$1_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$1
XXM2$1$1_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$1$1
XXM1$1$1_0 VSUBS XM1$1$1_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$1$1
XXM3$1_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$1
XXM0_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0_0/a_n346_583# XM0
C0 m1_n2669_n1117# m1_n1309_n1117# 0.027949f
C1 m1_n447_n1117# XM0_0/a_n346_583# 0.07096f
C2 XM0_0/a_n346_583# XM1$1$1_0/a_n202_583# 0.027386f
C3 m1_n2669_n1117# m1_n2738_n1819# 0.092062f
C4 m1_711_n1117# m1_802_n1819# 0.272119f
C5 m1_n1309_n1117# m1_n1378_n1819# 0.014034f
C6 m1_n1378_n1819# m1_n2738_n1819# 0.040124f
C7 m1_802_n1819# XM1$1$1_0/a_n202_583# 0.00859f
C8 m1_711_n1117# m1_n149_n1117# 0.02663f
C9 XM0_0/a_n346_583# m1_n1378_n1819# 0.039382f
C10 m1_n447_n1117# m1_n149_n1117# 0.123582f
C11 m1_n149_n1117# XM1$1$1_0/a_n202_583# 0.07096f
C12 m1_n447_n1117# m1_n1309_n1117# 0.041018f
C13 XM0_0/a_n346_583# VSUBS 0.314559f
C14 m1_n447_n1117# VSUBS 0.388025f
C15 m1_n2738_n1819# VSUBS 1.12292f
C16 m1_n2669_n1117# VSUBS 1.128649f
C17 XM1$1$1_0/a_n202_583# VSUBS 0.42776f
C18 m1_n149_n1117# VSUBS 0.407201f
C19 m1_n1378_n1819# VSUBS 0.604021f
C20 m1_n1309_n1117# VSUBS 0.637566f
C21 m1_802_n1819# VSUBS 1.278621f
C22 m1_711_n1117# VSUBS 1.959711f
.ends

.subckt trimb d_4 d_1 d_0 d_2 d_3 n1 n0 n3 drain n4 n2 VSUBS
Xtrim_switch_0 d_1 n0 d_4 d_0 d_3 n2 n4 d_2 n1 n3 VSUBS trim_switch
C0 n3 n4 1.600479f
C1 n2 n1 0.081094f
C2 n4 drain 12.877382f
C3 n0 n3 0.087807f
C4 n0 drain 1.60623f
C5 n3 drain 6.427485f
C6 n1 n4 0.169398f
C7 n2 d_1 0.003137f
C8 n1 n0 0.520979f
C9 n1 n3 0.087807f
C10 n1 drain 1.60623f
C11 n2 d_0 0.002632f
C12 n0 d_0 0.004139f
C13 n2 d_4 0.00312f
C14 n2 n4 0.596682f
C15 d_1 n1 0.003099f
C16 n2 n0 0.103368f
C17 n2 n3 0.58337f
C18 n2 drain 3.213024f
C19 n0 n4 0.166348f
C20 n2 VSUBS 2.03715f
C21 n0 VSUBS 0.689164f
C22 n1 VSUBS 0.727243f
C23 n4 VSUBS 4.367046f
C24 drain VSUBS -5.906306f
C25 n3 VSUBS 3.463842f
C26 d_0 VSUBS 0.33412f
C27 d_3 VSUBS 0.927186f
C28 d_1 VSUBS 0.345562f
C29 d_2 VSUBS 0.513348f
C30 d_4 VSUBS 1.64786f
.ends

.subckt XM2$3 a_69_n911# w_n237_n1121# a_5_n691# a_n75_n911# VSUBS
X0 a_69_n911# a_5_n691# a_n75_n911# w_n237_n1121# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 w_n237_n1121# a_5_n691# 0.131025f
C1 a_n75_n911# a_69_n911# 0.06854f
C2 a_69_n911# w_n237_n1121# 0.010275f
C3 a_n75_n911# w_n237_n1121# 0.008358f
C4 a_69_n911# a_5_n691# 0.001764f
C5 a_n75_n911# a_5_n691# 0.001764f
C6 a_69_n911# VSUBS 0.047486f
C7 a_n75_n911# VSUBS 0.049403f
C8 a_5_n691# VSUBS 0.087507f
C9 w_n237_n1121# VSUBS 1.54752f
.ends

.subckt XMl1 a_1362_n1100# a_1442_n880# a_1506_n1100# a_1224_n1284#
X0 a_1506_n1100# a_1442_n880# a_1362_n1100# a_1224_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_1442_n880# a_1362_n1100# 0.001764f
C1 a_1506_n1100# a_1442_n880# 0.001764f
C2 a_1506_n1100# a_1362_n1100# 0.06854f
C3 a_1506_n1100# a_1224_n1284# 0.057707f
C4 a_1362_n1100# a_1224_n1284# 0.066395f
C5 a_1442_n880# a_1224_n1284# 0.218606f
.ends

.subckt XMinp a_251_n1284# a_389_n1100# a_251_n788# a_469_n880# a_533_n1100#
X0 a_533_n1100# a_469_n880# a_389_n1100# a_251_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_389_n1100# a_533_n1100# 0.06854f
C1 a_533_n1100# a_469_n880# 0.001764f
C2 a_389_n1100# a_469_n880# 0.001764f
C3 a_533_n1100# a_251_n1284# 0.057707f
C4 a_389_n1100# a_251_n1284# 0.057707f
C5 a_469_n880# a_251_n1284# 0.21851f
.ends

.subckt comparator vdd vp vn trimb0 diff ip trimb_0/n3 outn clkc trim4 outp trim3
+ trim2 trim_0/n3 trim1 trim0 in trimb4 trim_0/n4 trimb3 trimb_0/n2 trim_0/n2 trimb2
+ trimb_0/n4 vss trimb1
XXMinn_0 vss vn in vss diff XMinn
XXM1$3_0 in clkc vdd vdd vss XM1$3
Xtrim_0 in trim4 trim1 trim0 trim2 trim3 trim_0/n1 trim_0/n0 trim_0/n3 trim_0/n4 trim_0/n2
+ vss trim
XXMl4_0 outn outp vdd vdd vss XMl4
XXM4$3_0 clkc ip vdd vdd vss XM4$3
XXMl2_0 outp ip outn vss XMl2
XXM3$3_0 outp vdd clkc vdd vss XM3$3
XXMdiff_0 diff clkc vss clkc vss vss XMdiff
XXMl3_0 outp vdd outn vdd vss XMl3
Xtrimb_0 trimb4 trimb1 trimb0 trimb2 trimb3 trimb_0/n1 trimb_0/n0 trimb_0/n3 ip trimb_0/n4
+ trimb_0/n2 vss trimb
XXM2$3_0 outn vdd clkc vdd vss XM2$3
XXMl1_0 outn outp in vss XMl1
XXMinp_0 vss diff vss vp ip XMinp
C0 vn outn 0.196568f
C1 trimb_0/n4 trimb_0/n0 0.032158f
C2 diff outp 0.006112f
C3 trim_0/n0 trim_0/n4 0.032158f
C4 trim_0/n2 trim_0/n4 0.128631f
C5 diff ip 0.133902f
C6 vp vn 0.180638f
C7 trim1 trim4 0.420884f
C8 diff in 0.133902f
C9 ip trimb_0/n0 1.606993f
C10 trimb_0/n4 trimb_0/n2 0.128631f
C11 trim2 trim0 0.78245f
C12 outp clkc 0.22388f
C13 outp outn 1.248977f
C14 trim_0/n1 in 1.606993f
C15 vdd clkc 0.233505f
C16 trimb_0/n4 trimb_0/n3 0.241184f
C17 ip clkc 0.46748f
C18 vdd outn 0.464524f
C19 trim0 trim4 0.001193f
C20 ip outn 0.016739f
C21 ip trimb_0/n2 3.21681f
C22 outp vp 0.243335f
C23 in clkc 0.467511f
C24 in outn 0.120156f
C25 trim_0/n0 in 1.606993f
C26 vp vdd 0.059928f
C27 trim_0/n2 in 3.21681f
C28 ip vp 0.542294f
C29 trim_0/n4 trim_0/n3 0.241184f
C30 ip trimb_0/n3 6.427209f
C31 trimb0 trimb1 0.720503f
C32 trim3 trim2 0.919951f
C33 trimb_0/n4 trimb_0/n1 0.032158f
C34 outp vn 0.223138f
C35 trimb0 trimb4 0.001193f
C36 vn vdd 0.059928f
C37 diff clkc 0.071648f
C38 trim0 trim1 0.720503f
C39 trimb3 trimb2 0.919951f
C40 diff outn 0.003297f
C41 trimb_0/n4 trimb1 0.001374f
C42 vn in 0.542295f
C43 ip trimb_0/n1 1.606993f
C44 trimb_0/n4 trimb4 0.002224f
C45 trim_0/n0 trim_0/n1 0.032158f
C46 trim_0/n4 trim4 0.002224f
C47 trimb0 trimb2 0.78245f
C48 diff vp 0.004194f
C49 trim_0/n4 in 12.853658f
C50 trimb4 trimb1 0.420884f
C51 ip trimb_0/n4 12.853658f
C52 trim_0/n3 in 6.427209f
C53 clkc outn 0.223756f
C54 outp vdd 0.441033f
C55 outp ip 0.120151f
C56 diff vn 0.004194f
C57 outp in 0.016739f
C58 ip vdd 0.088929f
C59 vp clkc 0.104841f
C60 vp outn 0.197573f
C61 trim_0/n4 trim1 0.001374f
C62 vdd in 0.088929f
C63 trim_0/n1 trim_0/n4 0.032158f
C64 trimb_0/n0 trimb_0/n1 0.032158f
C65 vn clkc 0.104842f
C66 vp vss 1.116181f
C67 outn vss 2.443821f
C68 vdd vss 7.878819f
C69 trimb_0/n2 vss 1.980196f
C70 trimb_0/n0 vss 0.677622f
C71 trimb_0/n1 vss 0.716105f
C72 trimb_0/n4 vss 4.199544f
C73 ip vss -4.381578f
C74 trimb_0/n3 vss 3.31053f
C75 trimb0 vss 0.985146f
C76 trimb3 vss 2.983196f
C77 trimb1 vss 0.99849f
C78 trimb2 vss 1.41065f
C79 trimb4 vss 2.263372f
C80 clkc vss 4.180552f
C81 outp vss 2.478554f
C82 trim_0/n4 vss 4.199544f
C83 in vss -4.381556f
C84 trim_0/n3 vss 3.31053f
C85 trim_0/n2 vss 1.980196f
C86 trim_0/n0 vss 0.677622f
C87 trim_0/n1 vss 0.716105f
C88 trim4 vss 2.263372f
C89 trim1 vss 0.99849f
C90 trim0 vss 0.985146f
C91 trim2 vss 1.41065f
C92 trim3 vss 2.983196f
C93 diff vss 0.21339f
C94 vn vss 1.131981f
.ends

.subckt cap_mim_2p0fF_RCWXT2$1 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
C0 m4_n3120_n3000# m4_n3240_n3120# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30_flip cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$1
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_RCWXT2 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
C0 m4_n3120_n3000# m4_n3240_n3120# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap1 m5_n86730_51500# m5_n11730_51500# m5_n33870_51500# m5_86130_51500#
+ m5_14520_n66196# m5_n18870_51500# m5_44520_n66196# m5_n30480_n66196# m5_74520_n66196#
+ m5_33270_51500# m5_11130_51500# m5_n480_n66196# m5_n60480_n66196# m5_18270_51500#
+ m5_n90480_n66196# m5_104520_n66196# m5_n41730_51500# m5_n63870_51500# m5_n26730_51500#
+ m5_n48870_51500# m5_n3870_51500# m5_n105480_n66196# m5_n101730_51500# m5_63270_51500#
+ m5_n108870_51500# m5_48270_51500# m5_41130_51500# m5_29520_n66196# m5_26130_51500#
+ m5_n15480_n66196# m5_n93870_51500# m5_59520_n66196# m5_3270_51500# m5_n71730_51500#
+ m5_n78870_51500# m5_n45480_n66196# m5_n56730_51500# m5_89520_n66196# m5_n75480_n66196#
+ m5_93270_51500# m5_71130_51500# m5_101130_51500# m5_78270_51500# m5_56130_51500#
+ m5_108270_51500# VSUBS
Xmim_cap_30_30_flip_233 m5_89520_n66196# mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_222 m5_14520_n66196# mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_200 m5_44520_n66196# mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_211 m5_n480_n66196# mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_68 m5_n45480_n66196# mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_57 m5_n15480_n66196# mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_79 m5_n75480_n66196# mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_13 m5_44520_n66196# mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_24 m5_44520_n66196# mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_46 m5_89520_n66196# mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_35 m5_29520_n66196# mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_213 m5_29520_n66196# m5_26130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_224 m5_104520_n66196# mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_202 m5_29520_n66196# mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_235 m5_59520_n66196# mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_212 m5_44520_n66196# m5_48270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_234 m5_74520_n66196# mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_223 m5_n480_n66196# mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_201 m5_29520_n66196# mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_58 m5_n30480_n66196# mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_69 m5_n30480_n66196# mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_14 m5_29520_n66196# mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_25 m5_29520_n66196# mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_47 m5_74520_n66196# mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_36 m5_104520_n66196# mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_214 m5_14520_n66196# m5_11130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_225 m5_89520_n66196# mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_203 m5_14520_n66196# mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_236 m5_59520_n66196# mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_224 m5_104520_n66196# m5_108270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_213 m5_29520_n66196# m5_33270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_235 m5_59520_n66196# mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_202 m5_14520_n66196# mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_59 m5_n45480_n66196# mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_15 m5_14520_n66196# mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_48 m5_59520_n66196# mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_26 m5_14520_n66196# mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_37 m5_104520_n66196# mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_226 m5_74520_n66196# mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_204 m5_14520_n66196# mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_237 m5_59520_n66196# mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_215 m5_44520_n66196# mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_225 m5_89520_n66196# m5_93270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_214 m5_14520_n66196# m5_18270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_236 m5_104520_n66196# mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_203 m5_n480_n66196# mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_16 m5_29520_n66196# mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_49 m5_59520_n66196# mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_38 m5_89520_n66196# mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_27 m5_14520_n66196# mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_227 m5_89520_n66196# mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_238 m5_59520_n66196# mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_205 m5_44520_n66196# mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_216 m5_29520_n66196# mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_226 m5_74520_n66196# m5_78270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_215 m5_n480_n66196# m5_3270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_237 m5_89520_n66196# mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_204 m5_44520_n66196# mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_17 m5_44520_n66196# mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_28 m5_44520_n66196# mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_39 m5_74520_n66196# mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_228 m5_104520_n66196# mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_217 m5_44520_n66196# mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_239 m5_59520_n66196# mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_206 m5_29520_n66196# mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_227 m5_59520_n66196# m5_63270_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_216 m5_44520_n66196# mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_238 m5_74520_n66196# mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_205 m5_29520_n66196# mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_18 m5_29520_n66196# mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_29 m5_29520_n66196# mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_229 m5_89520_n66196# mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_218 m5_29520_n66196# mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_207 m5_14520_n66196# mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_228 m5_104520_n66196# mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_217 m5_29520_n66196# mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_206 m5_14520_n66196# mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_239 m5_59520_n66196# mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_19 m5_14520_n66196# mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_219 m5_44520_n66196# mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_208 m5_29520_n66196# mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_229 m5_89520_n66196# mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_218 m5_14520_n66196# mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_207 m5_n480_n66196# mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_209 m5_14520_n66196# mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_219 m5_n480_n66196# mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_208 m5_44520_n66196# mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_190 m5_74520_n66196# mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_209 m5_29520_n66196# mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_90 m5_n90480_n66196# mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_180 m5_n30480_n66196# mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_191 m5_74520_n66196# mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_80 m5_n75480_n66196# mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_91 m5_n90480_n66196# mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_190 m5_74520_n66196# mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_170 m5_n45480_n66196# m5_n48870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_181 m5_n45480_n66196# mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_192 m5_104520_n66196# mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_81 m5_n90480_n66196# mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_70 m5_n15480_n66196# mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_92 m5_n75480_n66196# mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_0 m5_59520_n66196# mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_191 m5_59520_n66196# mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_180 m5_104520_n66196# mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_0 m5_89520_n66196# mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_160 m5_n105480_n66196# mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_193 m5_89520_n66196# mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_182 m5_n45480_n66196# mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_171 m5_n480_n66196# mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_60 m5_59520_n66196# mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_82 m5_n75480_n66196# mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_71 m5_n30480_n66196# mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_93 m5_n90480_n66196# mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_1 m5_104520_n66196# mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_170 m5_n60480_n66196# mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_192 m5_44520_n66196# mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_181 m5_89520_n66196# mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_1 m5_74520_n66196# mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_183 m5_n480_n66196# m5_n3870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_172 m5_n480_n66196# mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_150 m5_n60480_n66196# mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_194 m5_74520_n66196# mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_161 m5_n90480_n66196# mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_83 m5_n90480_n66196# mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_72 m5_n45480_n66196# mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_94 m5_n75480_n66196# mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_50 m5_74520_n66196# mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_61 m5_104520_n66196# mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_2 m5_89520_n66196# mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_160 m5_n30480_n66196# mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_193 m5_29520_n66196# mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_182 m5_74520_n66196# mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_171 m5_n60480_n66196# mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_2 m5_104520_n66196# mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_173 m5_n15480_n66196# mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_162 m5_n60480_n66196# mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_184 m5_89520_n66196# mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_195 m5_104520_n66196# mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_140 m5_n105480_n66196# mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_151 m5_n105480_n66196# mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_73 m5_n15480_n66196# mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_84 m5_n75480_n66196# mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_95 m5_n90480_n66196# mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_51 m5_59520_n66196# mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_40 m5_44520_n66196# mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_62 m5_89520_n66196# mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_3 m5_104520_n66196# mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_161 m5_n45480_n66196# mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_172 m5_n60480_n66196# mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_194 m5_14520_n66196# mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_183 m5_59520_n66196# mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_150 m5_n105480_n66196# mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_3 m5_89520_n66196# mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_174 m5_n30480_n66196# mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_152 m5_n75480_n66196# mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_141 m5_n105480_n66196# mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_196 m5_44520_n66196# mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_130 m5_n15480_n66196# mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_185 m5_104520_n66196# mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_163 m5_n105480_n66196# mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_30 m5_29520_n66196# mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_74 m5_n30480_n66196# mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_85 m5_n90480_n66196# mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_52 m5_104520_n66196# mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_96 m5_n105480_n66196# mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_41 m5_29520_n66196# mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_63 m5_74520_n66196# mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_4 m5_89520_n66196# mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_151 m5_n105480_n66196# mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_162 m5_n15480_n66196# mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_140 m5_n75480_n66196# mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_173 m5_n60480_n66196# mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_184 m5_104520_n66196# mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_195 m5_n480_n66196# mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_4 m5_74520_n66196# mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_131 m5_n30480_n66196# mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_120 m5_n30480_n66196# mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_153 m5_n90480_n66196# mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_186 m5_89520_n66196# mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_142 m5_n60480_n66196# mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_197 m5_44520_n66196# mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_164 m5_n60480_n66196# mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_175 m5_n15480_n66196# mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_31 m5_14520_n66196# mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_75 m5_n45480_n66196# mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_20 m5_29520_n66196# mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_64 m5_n15480_n66196# mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_86 m5_n75480_n66196# mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_42 m5_44520_n66196# mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_53 m5_89520_n66196# mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_97 m5_n105480_n66196# mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_5 m5_74520_n66196# mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_152 m5_n105480_n66196# m5_n101730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_163 m5_n30480_n66196# mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_141 m5_n90480_n66196# mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_174 m5_n60480_n66196# mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_130 m5_n45480_n66196# mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_196 m5_44520_n66196# mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_185 m5_89520_n66196# mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_5 m5_104520_n66196# mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_154 m5_n60480_n66196# m5_n63870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_176 m5_n45480_n66196# mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_165 m5_n60480_n66196# mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_110 m5_n480_n66196# mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_132 m5_n480_n66196# mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_121 m5_n45480_n66196# mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_143 m5_n75480_n66196# mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_198 m5_29520_n66196# mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_187 m5_104520_n66196# mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_76 m5_n105480_n66196# mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_21 m5_14520_n66196# mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_65 m5_n30480_n66196# mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_10 m5_104520_n66196# mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_32 m5_44520_n66196# mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_43 m5_29520_n66196# mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_54 m5_74520_n66196# mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_87 m5_n90480_n66196# mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_98 m5_n105480_n66196# mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_6 m5_59520_n66196# mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_153 m5_n75480_n66196# mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_164 m5_n45480_n66196# mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_175 m5_n60480_n66196# mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_131 m5_n15480_n66196# mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_142 m5_n75480_n66196# mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_120 m5_n15480_n66196# mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_197 m5_29520_n66196# mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_186 m5_74520_n66196# mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_6 m5_89520_n66196# mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_155 m5_n75480_n66196# m5_n78870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_166 m5_n75480_n66196# mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_111 m5_n15480_n66196# mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_100 m5_n105480_n66196# mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_133 m5_n15480_n66196# mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_144 m5_n90480_n66196# mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_122 m5_n30480_n66196# mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_199 m5_14520_n66196# mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_188 m5_89520_n66196# mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_177 m5_n30480_n66196# mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_77 m5_n105480_n66196# mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_22 m5_n480_n66196# mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_66 m5_n45480_n66196# mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_11 m5_89520_n66196# mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_99 m5_n105480_n66196# mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_33 m5_29520_n66196# mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_44 m5_14520_n66196# mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_55 m5_59520_n66196# mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_88 m5_n75480_n66196# mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_7 m5_74520_n66196# mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_110 m5_n30480_n66196# mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_121 m5_n30480_n66196# mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_154 m5_n90480_n66196# mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_176 m5_104520_n66196# mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_143 m5_n90480_n66196# mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_198 m5_14520_n66196# mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_187 m5_59520_n66196# mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_132 m5_n105480_n66196# mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_165 m5_n15480_n66196# mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_7 m5_104520_n66196# mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_156 m5_n90480_n66196# m5_n93870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_167 m5_n90480_n66196# mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_178 m5_n480_n66196# mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_101 m5_n105480_n66196# mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_112 m5_n30480_n66196# mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_145 m5_n75480_n66196# mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_123 m5_n45480_n66196# mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_189 m5_74520_n66196# mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_134 m5_n480_n66196# mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_23 m5_14520_n66196# mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_67 m5_n15480_n66196# mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_78 m5_n105480_n66196# mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_12 m5_74520_n66196# mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_34 m5_14520_n66196# mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_56 m5_104520_n66196# mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_45 m5_n480_n66196# mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_89 m5_n75480_n66196# mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_8 m5_59520_n66196# mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_100 m5_n45480_n66196# mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_111 m5_n15480_n66196# mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_177 m5_89520_n66196# mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_188 m5_104520_n66196# mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_133 m5_n105480_n66196# mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_122 m5_n45480_n66196# mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_199 m5_n480_n66196# mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_144 m5_n90480_n66196# mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_155 m5_n75480_n66196# mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_166 m5_n30480_n66196# mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_8 m5_89520_n66196# mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_168 m5_n15480_n66196# m5_n18870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_157 m5_n105480_n66196# m5_n108870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_179 m5_n15480_n66196# mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_102 m5_n105480_n66196# mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_113 m5_n45480_n66196# mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_135 m5_n45480_n66196# mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_146 m5_n60480_n66196# mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_124 m5_n15480_n66196# mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_68 m5_n30480_n66196# mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_79 m5_n105480_n66196# mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_24 m5_44520_n66196# mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_13 m5_59520_n66196# mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_35 m5_n480_n66196# mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_57 m5_89520_n66196# mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_46 m5_14520_n66196# mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_9 m5_104520_n66196# mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_156 m5_n15480_n66196# m5_n11730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_145 m5_n75480_n66196# mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_101 m5_n15480_n66196# mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_112 m5_n60480_n66196# mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_123 m5_n30480_n66196# mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_178 m5_74520_n66196# mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_134 m5_n105480_n66196# mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_189 m5_89520_n66196# mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_167 m5_n45480_n66196# mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_9 m5_74520_n66196# mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_103 m5_n105480_n66196# mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_114 m5_n480_n66196# mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_136 m5_n105480_n66196# mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_147 m5_n75480_n66196# mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_125 m5_n30480_n66196# mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_169 m5_n30480_n66196# m5_n33870_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_158 m5_n105480_n66196# mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_14 m5_89520_n66196# mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_69 m5_n45480_n66196# mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_25 m5_29520_n66196# mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_58 m5_74520_n66196# mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_36 m5_44520_n66196# mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_47 m5_n480_n66196# mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_157 m5_n30480_n66196# m5_n26730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_168 m5_n60480_n66196# m5_n56730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_146 m5_n90480_n66196# mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_113 m5_n60480_n66196# mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_102 m5_n30480_n66196# mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_135 m5_n105480_n66196# mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_124 m5_n45480_n66196# mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_179 m5_59520_n66196# mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_104 m5_n30480_n66196# mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_115 m5_n15480_n66196# mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_137 m5_n60480_n66196# mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_148 m5_n90480_n66196# mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_126 m5_n45480_n66196# mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_159 m5_n75480_n66196# mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_15 m5_74520_n66196# mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_26 m5_14520_n66196# mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_59 m5_59520_n66196# mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_37 m5_29520_n66196# mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_48 m5_104520_n66196# mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_158 m5_n45480_n66196# m5_n41730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_147 m5_n75480_n66196# m5_n71730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_169 m5_n60480_n66196# mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_114 m5_n60480_n66196# mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_103 m5_n45480_n66196# mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_136 m5_n75480_n66196# mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_125 m5_n15480_n66196# mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_105 m5_n45480_n66196# mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_116 m5_n30480_n66196# mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_149 m5_n90480_n66196# mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_138 m5_n75480_n66196# mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_127 m5_n480_n66196# mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_16 m5_n480_n66196# mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_27 m5_n480_n66196# mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_38 m5_14520_n66196# mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_49 m5_89520_n66196# mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_115 m5_n60480_n66196# mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_104 m5_n15480_n66196# mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_137 m5_n90480_n66196# mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_126 m5_n30480_n66196# mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_148 m5_n90480_n66196# m5_n86730_51500# VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_159 m5_n15480_n66196# mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_117 m5_n45480_n66196# mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_106 m5_n480_n66196# mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_139 m5_n90480_n66196# mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_128 m5_n15480_n66196# mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_17 m5_44520_n66196# mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_28 m5_n480_n66196# mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_39 m5_n480_n66196# mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_149 m5_n105480_n66196# mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_116 m5_n60480_n66196# mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_105 m5_n30480_n66196# mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_138 m5_n75480_n66196# mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_127 m5_n45480_n66196# mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_118 m5_n480_n66196# mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_107 m5_n15480_n66196# mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_129 m5_n480_n66196# mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_90 m5_n60480_n66196# mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_29 m5_44520_n66196# mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_18 m5_29520_n66196# mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_117 m5_n60480_n66196# mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_106 m5_n45480_n66196# mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_139 m5_n90480_n66196# mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_128 m5_n15480_n66196# mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_119 m5_n15480_n66196# mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_108 m5_n30480_n66196# mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_80 m5_n90480_n66196# mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_91 m5_n75480_n66196# mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_19 m5_44520_n66196# mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_118 m5_n60480_n66196# mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_107 m5_n15480_n66196# mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_129 m5_n30480_n66196# mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_109 m5_n45480_n66196# mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_70 m5_n45480_n66196# mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_81 m5_n60480_n66196# mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_92 m5_n90480_n66196# mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_119 m5_n60480_n66196# mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_108 m5_n30480_n66196# mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_82 m5_n75480_n66196# mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_60 m5_n30480_n66196# mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_71 m5_n15480_n66196# mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_93 m5_n60480_n66196# mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_109 m5_n45480_n66196# mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_50 m5_59520_n66196# mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_83 m5_n90480_n66196# mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_72 m5_n60480_n66196# mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_61 m5_n45480_n66196# mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_94 m5_n75480_n66196# mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_73 m5_n75480_n66196# mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_84 m5_n105480_n66196# mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_62 m5_n480_n66196# mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_95 m5_n90480_n66196# mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_51 m5_59520_n66196# mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_40 m5_89520_n66196# mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_74 m5_n90480_n66196# mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_52 m5_59520_n66196# mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_85 m5_n105480_n66196# mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_63 m5_n480_n66196# mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_96 m5_n75480_n66196# mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_30 m5_44520_n66196# mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_41 m5_74520_n66196# mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_230 m5_74520_n66196# mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_75 m5_n60480_n66196# mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_20 m5_29520_n66196# mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_64 m5_n15480_n66196# mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_86 m5_n105480_n66196# mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_53 m5_59520_n66196# mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_31 m5_29520_n66196# mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_42 m5_104520_n66196# mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_97 m5_n60480_n66196# mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_220 m5_104520_n66196# m5_101130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_231 m5_74520_n66196# mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_230 m5_74520_n66196# mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_65 m5_n480_n66196# mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_76 m5_n75480_n66196# mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_10 m5_74520_n66196# mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_54 m5_59520_n66196# mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_21 m5_14520_n66196# mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_87 m5_n105480_n66196# mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_32 m5_14520_n66196# mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_43 m5_89520_n66196# mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_98 m5_n75480_n66196# mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_221 m5_89520_n66196# m5_86130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_232 m5_59520_n66196# m5_56130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_210 m5_14520_n66196# mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_231 m5_59520_n66196# mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_220 m5_44520_n66196# mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_66 m5_n15480_n66196# mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_77 m5_n90480_n66196# mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_11 m5_104520_n66196# mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_22 m5_14520_n66196# mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_88 m5_n90480_n66196# mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_44 m5_74520_n66196# mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_99 m5_n90480_n66196# mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_33 m5_14520_n66196# mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_55 m5_59520_n66196# mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_222 m5_74520_n66196# m5_71130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_233 m5_59520_n66196# mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_200 m5_29520_n66196# mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_211 m5_14520_n66196# mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_232 m5_104520_n66196# mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_221 m5_29520_n66196# mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_210 m5_14520_n66196# mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_67 m5_n30480_n66196# mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_12 m5_44520_n66196# mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_23 m5_44520_n66196# mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_56 m5_n480_n66196# mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_78 m5_n60480_n66196# mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_89 m5_n60480_n66196# mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_45 m5_104520_n66196# mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_34 m5_44520_n66196# mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_212 m5_44520_n66196# m5_41130_51500# VSUBS mim_cap_30_30
Xmim_cap_30_30_234 m5_59520_n66196# mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_223 m5_104520_n66196# mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
Xmim_cap_30_30_201 m5_44520_n66196# mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS mim_cap_30_30
C0 mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C1 m5_n45480_n66196# m5_n41730_51500# 0.222064f
C2 mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C3 mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C4 mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C5 m5_n480_n66196# m5_n3870_51500# 0.222064f
C6 mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C7 m5_63270_51500# mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C8 mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C9 mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C10 m5_78270_51500# m5_74520_n66196# 0.222064f
C11 m5_n30480_n66196# m5_n15480_n66196# 5.150949f
C12 mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C13 mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C14 mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C15 mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C16 mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C17 mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C18 mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C19 mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C20 mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C21 mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C22 mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C23 mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C24 mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C25 mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C26 mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C27 mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C28 m5_44520_n66196# m5_29520_n66196# 5.150949f
C29 mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C30 mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C31 m5_n3870_51500# mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C32 mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C33 mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C34 mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C35 mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C36 mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C37 mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C38 mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C39 mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C40 mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C41 mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C42 mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C43 mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C44 m5_3270_51500# mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C45 mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C46 m5_n56730_51500# m5_n60480_n66196# 0.222064f
C47 m5_14520_n66196# m5_18270_51500# 0.222064f
C48 mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C49 mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C50 mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C51 mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C52 mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C53 mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C54 m5_n60480_n66196# m5_n75480_n66196# 5.150949f
C55 mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C56 mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C57 mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C58 mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C59 mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C60 mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C61 mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C62 mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C63 mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C64 mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C65 mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C66 mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C67 mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C68 m5_56130_51500# mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C69 mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C70 mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C71 mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C72 mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C73 mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C74 mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C75 mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C76 m5_26130_51500# mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C77 mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C78 mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C79 mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_101130_51500# 0.592904f
C80 mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C81 mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C82 m5_29520_n66196# m5_33270_51500# 0.222065f
C83 mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C84 m5_33270_51500# mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C85 mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C86 mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C87 mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C88 mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C89 mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C90 m5_n26730_51500# m5_n30480_n66196# 0.222064f
C91 m5_86130_51500# m5_89520_n66196# 0.222064f
C92 mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C93 mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C94 mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C95 m5_n45480_n66196# m5_n30480_n66196# 5.150949f
C96 mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C97 m5_n15480_n66196# m5_n18870_51500# 0.222064f
C98 mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C99 mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C100 mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C101 mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C102 mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C103 mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C104 mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C105 m5_74520_n66196# m5_89520_n66196# 5.150949f
C106 mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C107 mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C108 mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C109 mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C110 mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C111 mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C112 mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C113 mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C114 mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C115 mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C116 m5_89520_n66196# m5_104520_n66196# 2.575473f
C117 mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C118 mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C119 mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C120 mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C121 mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C122 mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C123 mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C124 mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C125 mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C126 mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C127 mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C128 mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C129 mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_18270_51500# 0.592904f
C130 m5_n11730_51500# mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C131 mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C132 mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C133 mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C134 mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C135 mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C136 mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C137 mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C138 mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C139 mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C140 mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C141 mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C142 mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C143 mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C144 mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C145 mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C146 mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C147 mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C148 mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C149 mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_108270_51500# 0.592904f
C150 mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C151 mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C152 mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C153 mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C154 mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C155 mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C156 mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C157 mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C158 mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C159 mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C160 mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C161 mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C162 mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C163 mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C164 mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C165 mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C166 mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C167 mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C168 mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C169 mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C170 mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C171 mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C172 mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C173 m5_14520_n66196# m5_11130_51500# 0.222064f
C174 mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C175 m5_101130_51500# m5_104520_n66196# 0.222064f
C176 mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C177 mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C178 m5_48270_51500# mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C179 mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C180 mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C181 mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C182 mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C183 mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C184 mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C185 m5_n75480_n66196# m5_n71730_51500# 0.222065f
C186 mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C187 mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C188 mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C189 mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C190 mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C191 mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C192 mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n71730_51500# 0.592904f
C193 mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C194 mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C195 mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C196 mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C197 mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C198 mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C199 mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C200 mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n93870_51500# 0.592904f
C201 mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C202 mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C203 mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C204 mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C205 mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C206 m5_108270_51500# m5_104520_n66196# 0.222064f
C207 mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C208 mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C209 mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C210 mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C211 m5_n78870_51500# m5_n75480_n66196# 0.222064f
C212 mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C213 m5_14520_n66196# m5_n480_n66196# 5.150949f
C214 mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C215 m5_n101730_51500# mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C216 mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C217 mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C218 mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C219 m5_44520_n66196# m5_59520_n66196# 5.150949f
C220 mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C221 mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_11130_51500# 0.592904f
C222 m5_n480_n66196# m5_n15480_n66196# 2.575473f
C223 mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C224 mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_86130_51500# 0.592904f
C225 mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n86730_51500# 0.592904f
C226 mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C227 mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C228 mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C229 mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C230 mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C231 mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C232 mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C233 mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C234 mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C235 mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C236 mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C237 mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C238 mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C239 mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C240 mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C241 mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C242 m5_56130_51500# m5_59520_n66196# 0.222064f
C243 mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C244 mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C245 mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C246 mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C247 mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C248 mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C249 mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C250 m5_n90480_n66196# m5_n75480_n66196# 5.150949f
C251 mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C252 mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C253 mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C254 m5_74520_n66196# m5_71130_51500# 0.222064f
C255 mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C256 mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C257 mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C258 mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C259 mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C260 mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C261 mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C262 mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C263 mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C264 mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C265 mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C266 mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C267 mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C268 mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C269 m5_63270_51500# m5_59520_n66196# 0.222064f
C270 mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C271 mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C272 mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C273 mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C274 mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C275 m5_n48870_51500# mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C276 mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C277 mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C278 mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C279 mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C280 mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C281 mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C282 mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C283 mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C284 m5_n45480_n66196# m5_n60480_n66196# 5.150949f
C285 mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C286 m5_n33870_51500# m5_n30480_n66196# 0.222064f
C287 mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C288 mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C289 m5_n26730_51500# mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C290 mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C291 m5_41130_51500# mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C292 mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C293 mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C294 mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C295 mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C296 mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C297 mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C298 mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C299 mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C300 mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C301 mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C302 mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C303 mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C304 mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C305 mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C306 mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C307 mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C308 m5_n105480_n66196# m5_n90480_n66196# 5.150949f
C309 mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C310 mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C311 mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C312 m5_93270_51500# mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C313 mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C314 mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C315 mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C316 mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C317 mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C318 mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C319 mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C320 mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C321 mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C322 mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C323 mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C324 mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C325 mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n33870_51500# 0.592904f
C326 mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C327 mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C328 mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C329 mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C330 mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C331 mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C332 mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C333 mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C334 mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C335 mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C336 mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C337 m5_93270_51500# m5_89520_n66196# 0.222064f
C338 mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C339 mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C340 mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C341 mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C342 mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C343 mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C344 mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C345 m5_n90480_n66196# m5_n93870_51500# 0.222064f
C346 mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C347 mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C348 mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C349 mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C350 mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C351 m5_44520_n66196# m5_48270_51500# 0.222064f
C352 mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C353 mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C354 m5_n63870_51500# m5_n60480_n66196# 0.222064f
C355 mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C356 mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C357 mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C358 mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C359 mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C360 mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C361 m5_n105480_n66196# m5_n108870_51500# 0.222064f
C362 mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C363 mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C364 mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C365 mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C366 mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C367 mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C368 mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C369 mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C370 mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C371 mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C372 m5_29520_n66196# m5_26130_51500# 0.222064f
C373 mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C374 mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C375 mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C376 mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C377 mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C378 mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C379 mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C380 mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C381 mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C382 mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C383 mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C384 mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C385 mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C386 m5_n90480_n66196# m5_n86730_51500# 0.222064f
C387 mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C388 mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C389 mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C390 mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C391 mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n108870_51500# 0.592904f
C392 mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C393 m5_n56730_51500# mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C394 mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C395 mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C396 mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C397 mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C398 mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C399 mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C400 mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C401 mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C402 mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C403 mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C404 mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C405 mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C406 mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C407 mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C408 mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C409 mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C410 mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C411 m5_n105480_n66196# m5_n101730_51500# 0.222064f
C412 mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C413 mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n78870_51500# 0.592904f
C414 m5_78270_51500# mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C415 mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C416 mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C417 mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C418 m5_44520_n66196# m5_41130_51500# 0.222064f
C419 mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C420 mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C421 mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C422 mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C423 mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C424 mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C425 mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C426 mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C427 m5_14520_n66196# m5_29520_n66196# 5.150949f
C428 mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C429 mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C430 mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C431 mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C432 mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C433 mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C434 mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C435 mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C436 mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C437 mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C438 mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C439 mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C440 mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C441 mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n18870_51500# 0.592904f
C442 mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C443 m5_3270_51500# m5_n480_n66196# 0.222064f
C444 mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C445 mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C446 mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C447 mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C448 mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C449 mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C450 mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C451 mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C452 mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C453 mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C454 mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C455 mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C456 mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C457 mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C458 mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C459 mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C460 mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C461 mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C462 mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_71130_51500# 0.592904f
C463 mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C464 mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C465 mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C466 m5_n15480_n66196# m5_n11730_51500# 0.222064f
C467 mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C468 mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C469 mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n41730_51500# 0.592904f
C470 mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C471 mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C472 mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C473 mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C474 mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C475 mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# m5_n63870_51500# 0.592904f
C476 mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C477 mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C478 mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C479 mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C480 mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C481 mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C482 m5_n45480_n66196# m5_n48870_51500# 0.222064f
C483 mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C484 mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C485 mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C486 m5_59520_n66196# m5_74520_n66196# 5.150949f
C487 mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C488 mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C489 mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C490 mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C491 mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C492 mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C493 mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# 0.592904f
C494 mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C495 mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C496 mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C497 m5_41130_51500# VSUBS 11.35416f
C498 mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C499 mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C500 mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C501 mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C502 mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C503 mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C504 m5_44520_n66196# VSUBS 0.145007p
C505 mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C506 mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C507 mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C508 mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C509 mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C510 mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C511 mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C512 mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C513 m5_71130_51500# VSUBS 11.35416f
C514 mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C515 mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C516 mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C517 mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C518 mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C519 mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C520 m5_14520_n66196# VSUBS 0.145007p
C521 mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C522 m5_104520_n66196# VSUBS 0.145007p
C523 mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C524 mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C525 mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C526 mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C527 mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C528 m5_56130_51500# VSUBS 11.35416f
C529 m5_86130_51500# VSUBS 11.35416f
C530 mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C531 mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C532 mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C533 mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C534 m5_n105480_n66196# VSUBS 0.145007p
C535 mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C536 mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C537 m5_59520_n66196# VSUBS 0.145007p
C538 mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C539 m5_74520_n66196# VSUBS 0.145007p
C540 mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C541 mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C542 mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C543 mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C544 m5_101130_51500# VSUBS 11.35416f
C545 mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C546 mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C547 mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C548 mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C549 mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C550 mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C551 m5_n15480_n66196# VSUBS 0.145007p
C552 mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C553 mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C554 mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C555 mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C556 mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C557 mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C558 mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C559 m5_n480_n66196# VSUBS 0.145007p
C560 mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C561 mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C562 mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C563 mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C564 mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C565 mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C566 mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C567 mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C568 mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C569 mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C570 mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C571 mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C572 mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C573 m5_n90480_n66196# VSUBS 0.145007p
C574 mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C575 mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C576 mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C577 mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C578 mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C579 mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C580 m5_n75480_n66196# VSUBS 0.145007p
C581 mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C582 mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C583 mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C584 mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C585 m5_n60480_n66196# VSUBS 0.145007p
C586 mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C587 m5_n45480_n66196# VSUBS 0.145007p
C588 mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C589 mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C590 mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C591 mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C592 mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C593 mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C594 mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C595 mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C596 mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C597 mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C598 mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C599 mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C600 mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C601 mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C602 mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C603 mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C604 mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C605 mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C606 mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C607 mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C608 mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C609 mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C610 mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C611 mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C612 mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C613 mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C614 mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C615 mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C616 mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C617 mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C618 mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C619 mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C620 m5_n86730_51500# VSUBS 11.35416f
C621 mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C622 mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C623 mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C624 mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C625 mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C626 mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C627 mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C628 mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C629 mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C630 mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C631 mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C632 mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C633 mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C634 mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C635 mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C636 mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C637 mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C638 mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C639 m5_n71730_51500# VSUBS 11.35416f
C640 m5_n41730_51500# VSUBS 11.35416f
C641 mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C642 mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C643 mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C644 mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C645 mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C646 mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C647 mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C648 mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C649 mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C650 mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C651 mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C652 mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C653 mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C654 mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C655 mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C656 mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C657 mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C658 m5_n56730_51500# VSUBS 11.35416f
C659 m5_n26730_51500# VSUBS 11.35416f
C660 mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C661 mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C662 mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C663 mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C664 mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C665 mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C666 mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C667 m5_n33870_51500# VSUBS 11.35416f
C668 mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C669 mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C670 mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C671 mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C672 mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C673 mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C674 mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C675 mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C676 mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C677 mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C678 mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C679 mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C680 mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C681 mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C682 m5_n11730_51500# VSUBS 11.35416f
C683 mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C684 mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C685 mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C686 mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C687 mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C688 mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C689 mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C690 mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C691 mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C692 mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C693 mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C694 mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C695 mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C696 mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C697 m5_n108870_51500# VSUBS 11.35416f
C698 m5_n18870_51500# VSUBS 11.35416f
C699 mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C700 mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C701 mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C702 mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C703 mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C704 mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C705 mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C706 mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C707 mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C708 mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C709 mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C710 mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C711 mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C712 mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C713 mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C714 mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C715 mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C716 mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C717 mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C718 mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C719 mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C720 mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C721 mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C722 mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C723 mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C724 mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C725 mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C726 mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C727 m5_n93870_51500# VSUBS 11.35416f
C728 mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C729 mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C730 mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C731 mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C732 mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C733 mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C734 mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C735 mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C736 mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C737 mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C738 mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C739 mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C740 mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C741 mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C742 mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C743 mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C744 mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C745 mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C746 mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C747 mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C748 mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C749 mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C750 mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C751 mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C752 mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C753 mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C754 mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C755 mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C756 mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C757 m5_n78870_51500# VSUBS 11.35416f
C758 mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C759 m5_89520_n66196# VSUBS 0.145007p
C760 mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C761 mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C762 mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C763 mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C764 mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C765 mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C766 mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C767 mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C768 mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C769 mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C770 mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C771 mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C772 mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C773 mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C774 mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C775 mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C776 mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C777 mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C778 mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C779 mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C780 mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C781 mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C782 mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C783 mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C784 mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C785 mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C786 m5_n63870_51500# VSUBS 11.35416f
C787 mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C788 mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C789 mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C790 mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C791 mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C792 mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C793 mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C794 m5_n101730_51500# VSUBS 11.35416f
C795 mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C796 mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C797 mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C798 mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C799 mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C800 mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C801 mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C802 mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C803 mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C804 mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C805 mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C806 mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C807 mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C808 mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C809 mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C810 mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C811 mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C812 mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C813 mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C814 mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C815 mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C816 mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C817 mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C818 mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C819 mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C820 mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C821 mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C822 mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C823 mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C824 mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C825 mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C826 mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C827 mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C828 mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C829 mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C830 mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C831 mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C832 mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C833 mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C834 mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C835 mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C836 mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C837 mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C838 mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C839 mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C840 mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C841 mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C842 mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C843 mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C844 mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C845 mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C846 mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C847 mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C848 mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C849 mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C850 mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C851 mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C852 mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C853 mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C854 mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C855 mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C856 mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C857 mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C858 mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C859 mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C860 mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C861 mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C862 mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C863 mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C864 mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C865 mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C866 mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C867 mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C868 m5_n3870_51500# VSUBS 11.35416f
C869 mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C870 mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C871 mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C872 mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C873 mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C874 mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C875 mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C876 mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C877 mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C878 mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C879 mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C880 mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C881 mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C882 mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C883 mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C884 mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C885 mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C886 mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C887 mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C888 mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C889 mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C890 mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C891 m5_n48870_51500# VSUBS 11.35416f
C892 mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C893 mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C894 mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C895 mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C896 mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C897 mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C898 mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C899 mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C900 mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C901 mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C902 mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C903 mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C904 mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C905 mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C906 mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C907 mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C908 mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C909 mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C910 mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C911 mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C912 mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C913 mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C914 mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C915 mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C916 mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C917 mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C918 mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C919 mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C920 mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C921 m5_63270_51500# VSUBS 11.35416f
C922 mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C923 mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C924 mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C925 mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C926 mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C927 mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C928 mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C929 mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C930 mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C931 m5_3270_51500# VSUBS 11.35416f
C932 m5_78270_51500# VSUBS 11.35416f
C933 mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C934 mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C935 mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C936 mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C937 mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C938 mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C939 mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C940 mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C941 m5_29520_n66196# VSUBS 0.145007p
C942 mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C943 mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C944 m5_18270_51500# VSUBS 11.35416f
C945 m5_93270_51500# VSUBS 11.35416f
C946 mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C947 mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C948 mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C949 mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C950 mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C951 mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C952 mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C953 mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C954 mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C955 mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C956 mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C957 m5_33270_51500# VSUBS 11.35416f
C958 m5_108270_51500# VSUBS 11.35416f
C959 mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C960 mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C961 mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C962 m5_11130_51500# VSUBS 11.35416f
C963 mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C964 mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C965 mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C966 mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C967 mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C968 m5_n30480_n66196# VSUBS 0.145007p
C969 mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C970 mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C971 mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C972 mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C973 m5_48270_51500# VSUBS 11.35416f
C974 mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C975 mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C976 mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C977 m5_26130_51500# VSUBS 11.35416f
C978 mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C979 mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C980 mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C981 mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C982 mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C983 mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C984 mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C985 mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C986 mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C987 mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C988 mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
.ends

.subckt cap_mim_2p0fF_DMYL6H m4_n114303_n17580# m4_n114183_n17460# VSUBS
X0 m4_n114183_n17460# m4_n114303_n17580# cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
C0 m4_n114183_n17460# m4_n114303_n17580# 8.5013f
C1 m4_n114183_n17460# VSUBS 85.381996f
C2 m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS cap_mim_2p0fF_DMYL6H
C0 cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt cap_mim_2p0fF_RCWXT2$2 m4_n3148_n3000# m4_n3268_n3120# VSUBS
X0 m4_n3148_n3000# m4_n3268_n3120# cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
C0 m4_n3148_n3000# m4_n3268_n3120# 2.57661f
C1 m4_n3148_n3000# VSUBS 9.60519f
C2 m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30$1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_DMYL6H$1 m4_93823_n2660# m4_93943_n2540# VSUBS
X0 m4_93943_n2540# m4_93823_n2660# cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
C0 m4_93943_n2540# m4_93823_n2660# 8.5013f
C1 m4_93943_n2540# VSUBS 85.381996f
C2 m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100$1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS cap_mim_2p0fF_DMYL6H$1
C0 cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap2 vdd vss VSUBS
Xmim_cap_100_100_0 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_1 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_2 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_20 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_0 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_3 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_21 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_22 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_1 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_10 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_11 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_4 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_23 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_2 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_12 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_24 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_3 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_13 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_4 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_14 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_5 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_6 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_15 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_16 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_7 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_8 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_17 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_9 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_18 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_19 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100$1_0 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_1 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_2 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_3 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_4 vss vdd VSUBS mim_cap_100_100$1
C0 vdd vss 0.270043p
C1 vdd VSUBS 1.380468p
C2 vss VSUBS 0.670421p
.ends

.subckt mim_cap_boss vss vdd VSUBS
Xmim_cap1_0 vdd vdd vdd vdd vss vdd vss vss vss vdd vdd vss vss vdd vss vss vdd vdd
+ vdd vdd vdd vss vdd vdd vdd vdd vdd vss vdd vss vdd vss vdd vdd vdd vss vdd vss
+ vss vdd vdd vdd vdd vdd vdd VSUBS mim_cap1
Xmim_cap2_0 vdd vss VSUBS mim_cap2
C0 vss vdd 0.664748p
C1 vdd VSUBS 3.062432p
C2 vss VSUBS 3.110667p
C3 mim_cap1_0/mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C4 mim_cap1_0/mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C5 mim_cap1_0/mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C6 mim_cap1_0/mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C7 mim_cap1_0/mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C8 mim_cap1_0/mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C9 mim_cap1_0/mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C10 mim_cap1_0/mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C11 mim_cap1_0/mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C12 mim_cap1_0/mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C13 mim_cap1_0/mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C14 mim_cap1_0/mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C15 mim_cap1_0/mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C16 mim_cap1_0/mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C17 mim_cap1_0/mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C18 mim_cap1_0/mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C19 mim_cap1_0/mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C20 mim_cap1_0/mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C21 mim_cap1_0/mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C22 mim_cap1_0/mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C23 mim_cap1_0/mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C24 mim_cap1_0/mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C25 mim_cap1_0/mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C26 mim_cap1_0/mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C27 mim_cap1_0/mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C28 mim_cap1_0/mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C29 mim_cap1_0/mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C30 mim_cap1_0/mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C31 mim_cap1_0/mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C32 mim_cap1_0/mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C33 mim_cap1_0/mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C34 mim_cap1_0/mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C35 mim_cap1_0/mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C36 mim_cap1_0/mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C37 mim_cap1_0/mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C38 mim_cap1_0/mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C39 mim_cap1_0/mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C40 mim_cap1_0/mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C41 mim_cap1_0/mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C42 mim_cap1_0/mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C43 mim_cap1_0/mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C44 mim_cap1_0/mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C45 mim_cap1_0/mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C46 mim_cap1_0/mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C47 mim_cap1_0/mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C48 mim_cap1_0/mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C49 mim_cap1_0/mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C50 mim_cap1_0/mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C51 mim_cap1_0/mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C52 mim_cap1_0/mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C53 mim_cap1_0/mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C54 mim_cap1_0/mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C55 mim_cap1_0/mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C56 mim_cap1_0/mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C57 mim_cap1_0/mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C58 mim_cap1_0/mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C59 mim_cap1_0/mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C60 mim_cap1_0/mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C61 mim_cap1_0/mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C62 mim_cap1_0/mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C63 mim_cap1_0/mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C64 mim_cap1_0/mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C65 mim_cap1_0/mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C66 mim_cap1_0/mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C67 mim_cap1_0/mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C68 mim_cap1_0/mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C69 mim_cap1_0/mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C70 mim_cap1_0/mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C71 mim_cap1_0/mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C72 mim_cap1_0/mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C73 mim_cap1_0/mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C74 mim_cap1_0/mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C75 mim_cap1_0/mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C76 mim_cap1_0/mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C77 mim_cap1_0/mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C78 mim_cap1_0/mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C79 mim_cap1_0/mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C80 mim_cap1_0/mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C81 mim_cap1_0/mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C82 mim_cap1_0/mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C83 mim_cap1_0/mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C84 mim_cap1_0/mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C85 mim_cap1_0/mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C86 mim_cap1_0/mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C87 mim_cap1_0/mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C88 mim_cap1_0/mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C89 mim_cap1_0/mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C90 mim_cap1_0/mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C91 mim_cap1_0/mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C92 mim_cap1_0/mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C93 mim_cap1_0/mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C94 mim_cap1_0/mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C95 mim_cap1_0/mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C96 mim_cap1_0/mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C97 mim_cap1_0/mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C98 mim_cap1_0/mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C99 mim_cap1_0/mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C100 mim_cap1_0/mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C101 mim_cap1_0/mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C102 mim_cap1_0/mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C103 mim_cap1_0/mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C104 mim_cap1_0/mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C105 mim_cap1_0/mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C106 mim_cap1_0/mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C107 mim_cap1_0/mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C108 mim_cap1_0/mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C109 mim_cap1_0/mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C110 mim_cap1_0/mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C111 mim_cap1_0/mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C112 mim_cap1_0/mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C113 mim_cap1_0/mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C114 mim_cap1_0/mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C115 mim_cap1_0/mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C116 mim_cap1_0/mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C117 mim_cap1_0/mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C118 mim_cap1_0/mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C119 mim_cap1_0/mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C120 mim_cap1_0/mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C121 mim_cap1_0/mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C122 mim_cap1_0/mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C123 mim_cap1_0/mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C124 mim_cap1_0/mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C125 mim_cap1_0/mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C126 mim_cap1_0/mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C127 mim_cap1_0/mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C128 mim_cap1_0/mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C129 mim_cap1_0/mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C130 mim_cap1_0/mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C131 mim_cap1_0/mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C132 mim_cap1_0/mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C133 mim_cap1_0/mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C134 mim_cap1_0/mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C135 mim_cap1_0/mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C136 mim_cap1_0/mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C137 mim_cap1_0/mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C138 mim_cap1_0/mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C139 mim_cap1_0/mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C140 mim_cap1_0/mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C141 mim_cap1_0/mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C142 mim_cap1_0/mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C143 mim_cap1_0/mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C144 mim_cap1_0/mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C145 mim_cap1_0/mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C146 mim_cap1_0/mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C147 mim_cap1_0/mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C148 mim_cap1_0/mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C149 mim_cap1_0/mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C150 mim_cap1_0/mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C151 mim_cap1_0/mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C152 mim_cap1_0/mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C153 mim_cap1_0/mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C154 mim_cap1_0/mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C155 mim_cap1_0/mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C156 mim_cap1_0/mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C157 mim_cap1_0/mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C158 mim_cap1_0/mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C159 mim_cap1_0/mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C160 mim_cap1_0/mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C161 mim_cap1_0/mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C162 mim_cap1_0/mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C163 mim_cap1_0/mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C164 mim_cap1_0/mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C165 mim_cap1_0/mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C166 mim_cap1_0/mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C167 mim_cap1_0/mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C168 mim_cap1_0/mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C169 mim_cap1_0/mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C170 mim_cap1_0/mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C171 mim_cap1_0/mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C172 mim_cap1_0/mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C173 mim_cap1_0/mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C174 mim_cap1_0/mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C175 mim_cap1_0/mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C176 mim_cap1_0/mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C177 mim_cap1_0/mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C178 mim_cap1_0/mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C179 mim_cap1_0/mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C180 mim_cap1_0/mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C181 mim_cap1_0/mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C182 mim_cap1_0/mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C183 mim_cap1_0/mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C184 mim_cap1_0/mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C185 mim_cap1_0/mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C186 mim_cap1_0/mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C187 mim_cap1_0/mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C188 mim_cap1_0/mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C189 mim_cap1_0/mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C190 mim_cap1_0/mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C191 mim_cap1_0/mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C192 mim_cap1_0/mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C193 mim_cap1_0/mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C194 mim_cap1_0/mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C195 mim_cap1_0/mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C196 mim_cap1_0/mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C197 mim_cap1_0/mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C198 mim_cap1_0/mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C199 mim_cap1_0/mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C200 mim_cap1_0/mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C201 mim_cap1_0/mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C202 mim_cap1_0/mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C203 mim_cap1_0/mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C204 mim_cap1_0/mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C205 mim_cap1_0/mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C206 mim_cap1_0/mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C207 mim_cap1_0/mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C208 mim_cap1_0/mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C209 mim_cap1_0/mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C210 mim_cap1_0/mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C211 mim_cap1_0/mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C212 mim_cap1_0/mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C213 mim_cap1_0/mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C214 mim_cap1_0/mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C215 mim_cap1_0/mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C216 mim_cap1_0/mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C217 mim_cap1_0/mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C218 mim_cap1_0/mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C219 mim_cap1_0/mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C220 mim_cap1_0/mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C221 mim_cap1_0/mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C222 mim_cap1_0/mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C223 mim_cap1_0/mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C224 mim_cap1_0/mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C225 mim_cap1_0/mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C226 mim_cap1_0/mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C227 mim_cap1_0/mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C228 mim_cap1_0/mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C229 mim_cap1_0/mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C230 mim_cap1_0/mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C231 mim_cap1_0/mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C232 mim_cap1_0/mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C233 mim_cap1_0/mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C234 mim_cap1_0/mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C235 mim_cap1_0/mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C236 mim_cap1_0/mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C237 mim_cap1_0/mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C238 mim_cap1_0/mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C239 mim_cap1_0/mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C240 mim_cap1_0/mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C241 mim_cap1_0/mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C242 mim_cap1_0/mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C243 mim_cap1_0/mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C244 mim_cap1_0/mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C245 mim_cap1_0/mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C246 mim_cap1_0/mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C247 mim_cap1_0/mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C248 mim_cap1_0/mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C249 mim_cap1_0/mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C250 mim_cap1_0/mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C251 mim_cap1_0/mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C252 mim_cap1_0/mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C253 mim_cap1_0/mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C254 mim_cap1_0/mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C255 mim_cap1_0/mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C256 mim_cap1_0/mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C257 mim_cap1_0/mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C258 mim_cap1_0/mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C259 mim_cap1_0/mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C260 mim_cap1_0/mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C261 mim_cap1_0/mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C262 mim_cap1_0/mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C263 mim_cap1_0/mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C264 mim_cap1_0/mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C265 mim_cap1_0/mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C266 mim_cap1_0/mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C267 mim_cap1_0/mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C268 mim_cap1_0/mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C269 mim_cap1_0/mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C270 mim_cap1_0/mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C271 mim_cap1_0/mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C272 mim_cap1_0/mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C273 mim_cap1_0/mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C274 mim_cap1_0/mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C275 mim_cap1_0/mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C276 mim_cap1_0/mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C277 mim_cap1_0/mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C278 mim_cap1_0/mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C279 mim_cap1_0/mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C280 mim_cap1_0/mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C281 mim_cap1_0/mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C282 mim_cap1_0/mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C283 mim_cap1_0/mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C284 mim_cap1_0/mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C285 mim_cap1_0/mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C286 mim_cap1_0/mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C287 mim_cap1_0/mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C288 mim_cap1_0/mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C289 mim_cap1_0/mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C290 mim_cap1_0/mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C291 mim_cap1_0/mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C292 mim_cap1_0/mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C293 mim_cap1_0/mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C294 mim_cap1_0/mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C295 mim_cap1_0/mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C296 mim_cap1_0/mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C297 mim_cap1_0/mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C298 mim_cap1_0/mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C299 mim_cap1_0/mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C300 mim_cap1_0/mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C301 mim_cap1_0/mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C302 mim_cap1_0/mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C303 mim_cap1_0/mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C304 mim_cap1_0/mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C305 mim_cap1_0/mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C306 mim_cap1_0/mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C307 mim_cap1_0/mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C308 mim_cap1_0/mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C309 mim_cap1_0/mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C310 mim_cap1_0/mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C311 mim_cap1_0/mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C312 mim_cap1_0/mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C313 mim_cap1_0/mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C314 mim_cap1_0/mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C315 mim_cap1_0/mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C316 mim_cap1_0/mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C317 mim_cap1_0/mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C318 mim_cap1_0/mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C319 mim_cap1_0/mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C320 mim_cap1_0/mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C321 mim_cap1_0/mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C322 mim_cap1_0/mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C323 mim_cap1_0/mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C324 mim_cap1_0/mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C325 mim_cap1_0/mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C326 mim_cap1_0/mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C327 mim_cap1_0/mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C328 mim_cap1_0/mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C329 mim_cap1_0/mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C330 mim_cap1_0/mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C331 mim_cap1_0/mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C332 mim_cap1_0/mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C333 mim_cap1_0/mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C334 mim_cap1_0/mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C335 mim_cap1_0/mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C336 mim_cap1_0/mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C337 mim_cap1_0/mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C338 mim_cap1_0/mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C339 mim_cap1_0/mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C340 mim_cap1_0/mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C341 mim_cap1_0/mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C342 mim_cap1_0/mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C343 mim_cap1_0/mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C344 mim_cap1_0/mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C345 mim_cap1_0/mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C346 mim_cap1_0/mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C347 mim_cap1_0/mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C348 mim_cap1_0/mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C349 mim_cap1_0/mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C350 mim_cap1_0/mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C351 mim_cap1_0/mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C352 mim_cap1_0/mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C353 mim_cap1_0/mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C354 mim_cap1_0/mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C355 mim_cap1_0/mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C356 mim_cap1_0/mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C357 mim_cap1_0/mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C358 mim_cap1_0/mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C359 mim_cap1_0/mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C360 mim_cap1_0/mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C361 mim_cap1_0/mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C362 mim_cap1_0/mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C363 mim_cap1_0/mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C364 mim_cap1_0/mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C365 mim_cap1_0/mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C366 mim_cap1_0/mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C367 mim_cap1_0/mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C368 mim_cap1_0/mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C369 mim_cap1_0/mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C370 mim_cap1_0/mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C371 mim_cap1_0/mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C372 mim_cap1_0/mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C373 mim_cap1_0/mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C374 mim_cap1_0/mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C375 mim_cap1_0/mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C376 mim_cap1_0/mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C377 mim_cap1_0/mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C378 mim_cap1_0/mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C379 mim_cap1_0/mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C380 mim_cap1_0/mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C381 mim_cap1_0/mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C382 mim_cap1_0/mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C383 mim_cap1_0/mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C384 mim_cap1_0/mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C385 mim_cap1_0/mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C386 mim_cap1_0/mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C387 mim_cap1_0/mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C388 mim_cap1_0/mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C389 mim_cap1_0/mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C390 mim_cap1_0/mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C391 mim_cap1_0/mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C392 mim_cap1_0/mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C393 mim_cap1_0/mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C394 mim_cap1_0/mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C395 mim_cap1_0/mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C396 mim_cap1_0/mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C397 mim_cap1_0/mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C398 mim_cap1_0/mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C399 mim_cap1_0/mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C400 mim_cap1_0/mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C401 mim_cap1_0/mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C402 mim_cap1_0/mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C403 mim_cap1_0/mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C404 mim_cap1_0/mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C405 mim_cap1_0/mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C406 mim_cap1_0/mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C407 mim_cap1_0/mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C408 mim_cap1_0/mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C409 mim_cap1_0/mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C410 mim_cap1_0/mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C411 mim_cap1_0/mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C412 mim_cap1_0/mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C413 mim_cap1_0/mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C414 mim_cap1_0/mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C415 mim_cap1_0/mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C416 mim_cap1_0/mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C417 mim_cap1_0/mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C418 mim_cap1_0/mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C419 mim_cap1_0/mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C420 mim_cap1_0/mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C421 mim_cap1_0/mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C422 mim_cap1_0/mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C423 mim_cap1_0/mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C424 mim_cap1_0/mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C425 mim_cap1_0/mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C426 mim_cap1_0/mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C427 mim_cap1_0/mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C428 mim_cap1_0/mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C429 mim_cap1_0/mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C430 mim_cap1_0/mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C431 mim_cap1_0/mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C432 mim_cap1_0/mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C433 mim_cap1_0/mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C434 mim_cap1_0/mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C435 mim_cap1_0/mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C436 mim_cap1_0/mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C437 mim_cap1_0/mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C438 mim_cap1_0/mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C439 mim_cap1_0/mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C440 mim_cap1_0/mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C441 mim_cap1_0/mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C442 mim_cap1_0/mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C443 mim_cap1_0/mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C444 mim_cap1_0/mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C445 mim_cap1_0/mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C446 mim_cap1_0/mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C447 mim_cap1_0/mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C448 mim_cap1_0/mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C449 mim_cap1_0/mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C450 mim_cap1_0/mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C451 mim_cap1_0/mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C452 mim_cap1_0/mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW a_36_472# a_572_375# a_124_375#
+ a_484_472#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VDD a_484_472# 0.179463f
C1 a_36_472# a_484_472# 0.013276f
C2 a_484_472# VSS 0.148682f
C3 VDD a_124_375# 0.12673f
C4 a_36_472# a_124_375# 0.285629f
C5 a_124_375# VSS 0.136476f
C6 VDD VNW 0.11314f
C7 VSS VNW 0.008822f
C8 a_36_472# VNW 0.025611f
C9 a_484_472# a_572_375# 0.285629f
C10 a_124_375# a_572_375# 0.012222f
C11 a_572_375# VNW 0.18122f
C12 a_124_375# a_484_472# 0.086742f
C13 a_484_472# VNW 0.024396f
C14 a_124_375# VNW 0.180172f
C15 a_36_472# VDD 0.093681f
C16 VDD VSS 0.013184f
C17 a_36_472# VSS 0.151218f
C18 VDD a_572_375# 0.129266f
C19 VSS a_572_375# 0.082563f
C20 VSS VPW 0.360066f
C21 VDD VPW 0.286281f
C22 VNW VPW 1.65967f
C23 a_484_472# VPW 0.345058f
C24 a_36_472# VPW 0.404746f
C25 a_572_375# VPW 0.232991f
C26 a_124_375# VPW 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VNW VPW
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 VDD VNW 0.048519f
C1 VDD I 0.017439f
C2 I VNW 0.027206f
C3 VDD VSS 0.009725f
C4 VSS VNW 0.007461f
C5 I VSS 0.031625f
C6 VSS VPW 0.12617f
C7 VDD VPW 0.087026f
C8 I VPW 0.139667f
C9 VNW VPW 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW a_224_472#
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 VNW VDD 0.093678f
C1 A1 VDD 0.028041f
C2 VSS VDD 0.023219f
C3 A2 VNW 0.128798f
C4 ZN VDD 0.117921f
C5 ZN a_224_472# 0.023693f
C6 A2 A1 0.037814f
C7 VSS A2 0.043352f
C8 VDD a_224_472# 0.013964f
C9 A2 ZN 0.378409f
C10 VNW A1 0.136915f
C11 VSS VNW 0.010571f
C12 VSS A1 0.168633f
C13 A2 VDD 0.255318f
C14 A2 a_224_472# 0.008979f
C15 VNW ZN 0.019783f
C16 A1 ZN 0.579732f
C17 VSS ZN 0.08687f
C18 VSS VPW 0.331491f
C19 ZN VPW 0.058886f
C20 VDD VPW 0.218051f
C21 A1 VPW 0.331856f
C22 A2 VPW 0.334514f
C23 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VNW VPW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_1456_156#
+ a_1288_156# a_2248_156# a_2560_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VPW nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 VNW a_2665_112# 0.354715f
C1 RN a_2665_112# 0.336469f
C2 VNW a_2248_156# 0.212431f
C3 RN a_2248_156# 0.094336f
C4 a_1204_472# VNW 0.016269f
C5 RN a_1204_472# 0.021039f
C6 VNW VDD 0.503557f
C7 RN VDD 0.034984f
C8 a_2248_156# a_1000_472# 0.001232f
C9 VSS VNW 0.010602f
C10 VSS RN 0.441968f
C11 a_1204_472# a_1000_472# 0.66083f
C12 a_1000_472# VDD 0.119211f
C13 VSS a_1000_472# 0.04356f
C14 RN a_3041_156# 0.01068f
C15 a_796_472# D 0.082858f
C16 a_448_472# a_1456_156# 0.00227f
C17 a_2560_156# a_448_472# 0.277491f
C18 RN VNW 0.329494f
C19 a_796_472# a_448_472# 0.401636f
C20 a_2560_156# a_36_151# 0.003674f
C21 VNW a_1000_472# 0.241357f
C22 RN a_1000_472# 0.0832f
C23 a_448_472# a_1308_423# 0.882105f
C24 a_796_472# a_36_151# 0.011851f
C25 a_36_151# a_1308_423# 0.05539f
C26 a_448_472# a_2665_112# 0.020455f
C27 CLK VDD 0.02303f
C28 a_1288_156# VSS 0.001702f
C29 D VDD 0.009367f
C30 VSS CLK 0.021952f
C31 VSS D 0.064618f
C32 a_448_472# a_2248_156# 0.510371f
C33 a_36_151# a_2665_112# 0.019043f
C34 a_448_472# a_1204_472# 0.008996f
C35 a_448_472# VDD 0.456269f
C36 a_2248_156# a_36_151# 0.042802f
C37 VSS a_448_472# 1.20207f
C38 a_1204_472# a_36_151# 0.006996f
C39 a_36_151# VDD 0.417088f
C40 CLK VNW 0.137037f
C41 VSS a_36_151# 0.291264f
C42 VNW D 0.128231f
C43 a_448_472# VNW 0.341284f
C44 a_448_472# RN 0.078731f
C45 VNW a_36_151# 1.28833f
C46 a_448_472# a_1000_472# 0.361958f
C47 RN a_36_151# 0.080102f
C48 Q a_2665_112# 0.109436f
C49 a_1000_472# a_36_151# 0.08126f
C50 a_2560_156# a_2665_112# 0.116059f
C51 a_2248_156# Q 0.014355f
C52 a_2560_156# a_2248_156# 0.119687f
C53 Q VDD 0.149344f
C54 VSS Q 0.113401f
C55 a_2560_156# VDD 0.00217f
C56 VSS a_1456_156# 0.001901f
C57 VSS a_2560_156# 0.128503f
C58 a_2248_156# a_1308_423# 0.056721f
C59 VSS a_796_472# 0.05215f
C60 a_1204_472# a_1308_423# 0.026665f
C61 a_1288_156# a_448_472# 0.002067f
C62 a_1308_423# VDD 0.094185f
C63 a_448_472# CLK 0.002757f
C64 VSS a_1308_423# 0.013866f
C65 a_448_472# D 0.328788f
C66 VNW Q 0.034443f
C67 a_2248_156# a_2665_112# 0.633318f
C68 a_2560_156# VNW 0.020165f
C69 CLK a_36_151# 0.669598f
C70 a_2560_156# RN 0.038779f
C71 a_2665_112# VDD 0.102046f
C72 D a_36_151# 0.094113f
C73 a_796_472# VNW 0.010232f
C74 VSS a_2665_112# 0.184997f
C75 a_2248_156# VDD 1.11667f
C76 a_448_472# a_36_151# 0.536965f
C77 a_1204_472# VDD 0.282626f
C78 VNW a_1308_423# 0.149014f
C79 a_3041_156# a_2665_112# 0.001774f
C80 VSS a_2248_156# 0.030473f
C81 a_796_472# a_1000_472# 0.048436f
C82 RN a_1308_423# 0.079294f
C83 VSS VDD 0.01338f
C84 a_1000_472# a_1308_423# 0.934191f
C85 Q VPW 0.114762f
C86 VSS VPW 1.26186f
C87 RN VPW 1.36673f
C88 D VPW 0.253406f
C89 VDD VPW 0.79945f
C90 CLK VPW 0.291241f
C91 VNW VPW 6.1377f
C92 a_2560_156# VPW 0.016968f
C93 a_2665_112# VPW 0.62251f
C94 a_2248_156# VPW 0.371662f
C95 a_1204_472# VPW 0.012971f
C96 a_1000_472# VPW 0.291735f
C97 a_796_472# VPW 0.023206f
C98 a_1308_423# VPW 0.279043f
C99 a_448_472# VPW 0.684413f
C100 a_36_151# VPW 1.43589f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VNW VPW a_36_68# a_244_472#
+ a_692_472#
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 B2 VDD 0.246452f
C1 B2 a_244_472# 0.002003f
C2 VSS B1 0.025138f
C3 a_36_68# B1 0.437534f
C4 VNW VSS 0.010714f
C5 a_36_68# a_692_472# 0.015646f
C6 a_36_68# VNW 0.040298f
C7 VNW B1 0.125926f
C8 VSS ZN 0.085273f
C9 VSS A1 0.084232f
C10 a_36_68# ZN 0.419486f
C11 a_36_68# A1 0.160084f
C12 VSS VDD 0.011512f
C13 VSS A2 0.087422f
C14 a_36_68# VDD 0.787847f
C15 a_36_68# A2 0.340509f
C16 a_36_68# a_244_472# 0.027448f
C17 B1 ZN 0.079f
C18 A1 B1 0.163724f
C19 a_692_472# ZN 0.011665f
C20 VNW ZN 0.010694f
C21 VNW A1 0.115376f
C22 B1 VDD 0.014643f
C23 a_692_472# VDD 0.004194f
C24 VNW VDD 0.139306f
C25 VNW A2 0.125671f
C26 a_244_472# B1 0.003598f
C27 A1 ZN 0.430191f
C28 VDD ZN 0.004634f
C29 A2 ZN 0.390894f
C30 A1 VDD 0.014671f
C31 A1 A2 0.038725f
C32 B2 VSS 0.025295f
C33 a_36_68# B2 0.369561f
C34 A2 VDD 0.019572f
C35 a_244_472# VDD 0.00636f
C36 B2 B1 0.036483f
C37 VNW B2 0.133721f
C38 a_36_68# VSS 0.392965f
C39 VSS VPW 0.383233f
C40 ZN VPW 0.012598f
C41 VDD VPW 0.318857f
C42 A2 VPW 0.2826f
C43 A1 VPW 0.258579f
C44 B1 VPW 0.257485f
C45 B2 VPW 0.309037f
C46 VNW VPW 2.00777f
C47 a_36_68# VPW 0.150048f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW a_49_472#
+ a_665_69# a_257_69#
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
C0 VNW VSS 0.011011f
C1 ZN VNW 0.017894f
C2 VSS a_665_69# 0.003829f
C3 ZN a_665_69# 0.001059f
C4 A2 VSS 0.150463f
C5 VDD VNW 0.112326f
C6 VSS a_257_69# 0.00576f
C7 A2 ZN 0.102518f
C8 VSS a_49_472# 0.02154f
C9 ZN a_49_472# 0.239204f
C10 VSS B2 0.06757f
C11 ZN B2 0.001886f
C12 VDD A2 0.013575f
C13 VNW A1 0.10965f
C14 VDD a_49_472# 0.887006f
C15 A1 a_665_69# 0.002008f
C16 VDD B2 0.026097f
C17 A2 A1 0.392541f
C18 A1 a_49_472# 0.021757f
C19 VSS B1 0.095385f
C20 ZN B1 0.367665f
C21 VDD B1 0.017923f
C22 A1 B1 0.041046f
C23 A2 VNW 0.131727f
C24 VNW a_49_472# 0.026629f
C25 A2 a_665_69# 0.006702f
C26 VNW B2 0.129409f
C27 A2 a_49_472# 0.075759f
C28 B2 a_257_69# 0.003563f
C29 a_49_472# B2 0.151151f
C30 ZN VSS 0.071892f
C31 VNW B1 0.109456f
C32 VDD VSS 0.00787f
C33 VDD ZN 0.004108f
C34 B1 a_257_69# 0.003901f
C35 a_49_472# B1 0.069833f
C36 B1 B2 0.18297f
C37 A1 VSS 0.087393f
C38 ZN A1 0.447732f
C39 VDD A1 0.013859f
C40 VSS VPW 0.39457f
C41 ZN VPW 0.021794f
C42 VDD VPW 0.243433f
C43 A2 VPW 0.322629f
C44 A1 VPW 0.250967f
C45 B1 VPW 0.261124f
C46 B2 VPW 0.322244f
C47 VNW VPW 1.83372f
C48 a_49_472# VPW 0.054843f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VNW VPW a_36_160#
X0 Z a_36_160# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VPW nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VDD I 0.02612f
C1 VNW VDD 0.087464f
C2 Z VDD 0.128274f
C3 VSS VDD 0.009574f
C4 a_36_160# I 0.545454f
C5 a_36_160# VNW 0.170864f
C6 Z a_36_160# 0.281838f
C7 VSS a_36_160# 0.074156f
C8 a_36_160# VDD 0.2736f
C9 VNW I 0.2276f
C10 Z I 0.041707f
C11 VSS I 0.12329f
C12 Z VNW 0.030347f
C13 VSS VNW 0.009324f
C14 VSS Z 0.146199f
C15 VSS VPW 0.28275f
C16 Z VPW 0.10469f
C17 VDD VPW 0.178615f
C18 I VPW 0.323491f
C19 VNW VPW 1.31158f
C20 a_36_160# VPW 0.386641f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 ZN VDD 0.098026f
C1 I ZN 0.47009f
C2 VSS ZN 0.077008f
C3 VNW ZN 0.031181f
C4 I VDD 0.157124f
C5 VSS VDD 0.025441f
C6 VSS I 0.058937f
C7 VNW VDD 0.076212f
C8 VNW I 0.135368f
C9 VNW VSS 0.011085f
C10 VSS VPW 0.242183f
C11 ZN VPW 0.095505f
C12 VDD VPW 0.182097f
C13 I VPW 0.355642f
C14 VNW VPW 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 ZN VDD 0.137375f
C1 I ZN 0.262199f
C2 VSS ZN 0.115297f
C3 VNW ZN 0.022202f
C4 I VDD 0.041847f
C5 VSS VDD 0.025626f
C6 VSS I 0.0533f
C7 VNW VDD 0.076257f
C8 VNW I 0.137757f
C9 VNW VSS 0.011339f
C10 VSS VPW 0.2316f
C11 ZN VPW 0.113404f
C12 VDD VPW 0.181139f
C13 I VPW 0.341982f
C14 VNW VPW 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW a_36_472# a_124_375#
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VDD VNW 0.061035f
C1 VSS VDD 0.006592f
C2 a_36_472# VDD 0.093681f
C3 a_124_375# VNW 0.179924f
C4 VSS a_124_375# 0.082879f
C5 a_36_472# a_124_375# 0.285629f
C6 a_124_375# VDD 0.126034f
C7 VSS VNW 0.004411f
C8 a_36_472# VNW 0.025989f
C9 a_36_472# VSS 0.150876f
C10 VSS VPW 0.218985f
C11 VDD VPW 0.182777f
C12 VNW VPW 0.96348f
C13 a_36_472# VPW 0.417394f
C14 a_124_375# VPW 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VNW VPW a_224_472#
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 VDD I 0.1311f
C1 VNW VDD 0.305516f
C2 Z VDD 0.819024f
C3 VSS VDD 0.031131f
C4 a_224_472# I 0.796069f
C5 a_224_472# VNW 1.14633f
C6 Z a_224_472# 2.29481f
C7 VSS a_224_472# 0.659695f
C8 a_224_472# VDD 0.74621f
C9 VNW I 0.55539f
C10 Z I 0.001907f
C11 VSS I 0.158668f
C12 Z VNW 0.038011f
C13 VSS VNW 0.01282f
C14 VSS Z 0.70427f
C15 VSS VPW 0.910368f
C16 Z VPW 0.18914f
C17 VDD VPW 0.724491f
C18 I VPW 1.16773f
C19 VNW VPW 4.79254f
C20 a_224_472# VPW 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW a_36_472# a_244_68#
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
C0 VSS ZN 0.304078f
C1 A2 VDD 0.015143f
C2 A2 VNW 0.128282f
C3 A1 A2 0.047589f
C4 a_36_472# VDD 0.581285f
C5 a_36_472# VNW 0.013943f
C6 A1 a_36_472# 0.104556f
C7 B a_36_472# 0.01027f
C8 VDD ZN 0.003129f
C9 VSS VDD 0.01275f
C10 VNW ZN 0.014655f
C11 VSS VNW 0.009145f
C12 A1 ZN 0.245346f
C13 B ZN 0.00761f
C14 A1 VSS 0.021732f
C15 B VSS 0.080416f
C16 a_244_68# ZN 0.008784f
C17 a_244_68# VSS 0.00255f
C18 a_36_472# A2 0.10395f
C19 VNW VDD 0.11216f
C20 A2 ZN 0.248411f
C21 VSS A2 0.069479f
C22 A1 VDD 0.0167f
C23 B VDD 0.071777f
C24 A1 VNW 0.122087f
C25 B VNW 0.137038f
C26 a_36_472# ZN 0.088503f
C27 a_36_472# VSS 0.004325f
C28 B A1 0.157699f
C29 VSS VPW 0.361309f
C30 VDD VPW 0.259458f
C31 ZN VPW 0.040013f
C32 B VPW 0.378232f
C33 A1 VPW 0.264815f
C34 A2 VPW 0.3189f
C35 VNW VPW 1.65967f
C36 a_36_472# VPW 0.031137f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW a_36_113#
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 a_36_113# VSS 0.11114f
C1 I a_36_113# 0.476912f
C2 VDD Z 0.085355f
C3 VNW VSS 0.009307f
C4 VNW I 0.152645f
C5 Z a_36_113# 0.191876f
C6 VDD a_36_113# 0.278283f
C7 I VSS 0.070302f
C8 Z VNW 0.030118f
C9 VDD VNW 0.088196f
C10 Z VSS 0.136942f
C11 VDD VSS 0.009561f
C12 VNW a_36_113# 0.160792f
C13 Z I 0.031362f
C14 VDD I 0.028968f
C15 VSS VPW 0.283681f
C16 Z VPW 0.117185f
C17 VDD VPW 0.180237f
C18 I VPW 0.336876f
C19 VNW VPW 1.31158f
C20 a_36_113# VPW 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW a_1916_375# a_1380_472#
+ a_3260_375# a_36_472# a_932_472# a_2812_375# a_2276_472# a_1828_472# a_3172_472#
+ a_572_375# a_2724_472# a_124_375# a_1468_375# a_1020_375# a_484_472# a_2364_375#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_2724_472# VDD 0.179463f
C1 VNW a_1916_375# 0.181468f
C2 a_3260_375# a_3172_472# 0.285629f
C3 a_2364_375# VDD 0.129962f
C4 a_1916_375# VDD 0.129962f
C5 a_2724_472# a_3172_472# 0.013276f
C6 VNW a_124_375# 0.180172f
C7 VSS a_1828_472# 0.142721f
C8 a_1020_375# VSS 0.131736f
C9 a_484_472# VNW 0.024018f
C10 a_2276_472# VSS 0.142721f
C11 a_932_472# a_484_472# 0.013276f
C12 VDD a_124_375# 0.12673f
C13 a_484_472# VDD 0.179463f
C14 a_2364_375# a_2724_472# 0.087174f
C15 VSS a_2812_375# 0.131736f
C16 a_124_375# a_36_472# 0.285629f
C17 a_2276_472# a_1828_472# 0.013276f
C18 a_484_472# a_36_472# 0.013276f
C19 a_1916_375# a_2364_375# 0.013103f
C20 a_572_375# a_124_375# 0.013103f
C21 a_484_472# a_572_375# 0.285629f
C22 a_1468_375# VSS 0.131736f
C23 VNW VSS 0.035286f
C24 a_1020_375# a_1468_375# 0.013103f
C25 a_1468_375# a_1828_472# 0.087174f
C26 a_932_472# VSS 0.142721f
C27 VNW a_1020_375# 0.181468f
C28 VNW a_1828_472# 0.024018f
C29 VSS VDD 0.052737f
C30 VSS a_1380_472# 0.142721f
C31 a_932_472# a_1020_375# 0.285629f
C32 VSS a_36_472# 0.142026f
C33 VNW a_2276_472# 0.024018f
C34 a_1020_375# VDD 0.129962f
C35 VDD a_1828_472# 0.179463f
C36 a_1020_375# a_1380_472# 0.087174f
C37 a_1380_472# a_1828_472# 0.013276f
C38 VNW a_2812_375# 0.181468f
C39 a_572_375# VSS 0.131736f
C40 a_3260_375# VSS 0.081304f
C41 VSS a_3172_472# 0.139489f
C42 a_2276_472# VDD 0.179463f
C43 a_572_375# a_1020_375# 0.013103f
C44 VDD a_2812_375# 0.129962f
C45 VNW a_1468_375# 0.181468f
C46 a_2724_472# VSS 0.142721f
C47 a_484_472# a_124_375# 0.087174f
C48 a_2364_375# VSS 0.131736f
C49 a_1468_375# VDD 0.129962f
C50 a_932_472# VNW 0.024018f
C51 a_1916_375# VSS 0.131736f
C52 a_1468_375# a_1380_472# 0.285629f
C53 a_3260_375# a_2812_375# 0.013103f
C54 a_2812_375# a_3172_472# 0.087174f
C55 VNW VDD 0.425768f
C56 VNW a_1380_472# 0.024018f
C57 a_2276_472# a_2724_472# 0.013276f
C58 VNW a_36_472# 0.025611f
C59 a_1916_375# a_1828_472# 0.285629f
C60 a_932_472# VDD 0.179463f
C61 a_2364_375# a_2276_472# 0.285629f
C62 a_932_472# a_1380_472# 0.013276f
C63 a_2724_472# a_2812_375# 0.285629f
C64 VDD a_1380_472# 0.179463f
C65 a_572_375# VNW 0.181468f
C66 a_1916_375# a_2276_472# 0.087174f
C67 a_3260_375# VNW 0.18122f
C68 VNW a_3172_472# 0.024396f
C69 a_2364_375# a_2812_375# 0.013103f
C70 VSS a_124_375# 0.131736f
C71 VDD a_36_472# 0.093681f
C72 a_484_472# VSS 0.142721f
C73 a_932_472# a_572_375# 0.087174f
C74 a_572_375# VDD 0.129962f
C75 a_3260_375# VDD 0.129266f
C76 VDD a_3172_472# 0.179463f
C77 VNW a_2724_472# 0.024018f
C78 VNW a_2364_375# 0.181468f
C79 a_1916_375# a_1468_375# 0.013103f
C80 VSS VPW 1.20585f
C81 VDD VPW 0.907304f
C82 VNW VPW 5.83682f
C83 a_3172_472# VPW 0.345058f
C84 a_2724_472# VPW 0.33241f
C85 a_2276_472# VPW 0.33241f
C86 a_1828_472# VPW 0.33241f
C87 a_1380_472# VPW 0.33241f
C88 a_932_472# VPW 0.33241f
C89 a_484_472# VPW 0.33241f
C90 a_36_472# VPW 0.404746f
C91 a_3260_375# VPW 0.233093f
C92 a_2812_375# VPW 0.17167f
C93 a_2364_375# VPW 0.17167f
C94 a_1916_375# VPW 0.17167f
C95 a_1468_375# VPW 0.17167f
C96 a_1020_375# VPW 0.17167f
C97 a_572_375# VPW 0.17167f
C98 a_124_375# VPW 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_455_68# a_271_68#
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 VSS VNW 0.008577f
C1 ZN a_271_68# 0.001916f
C2 VDD A3 0.079999f
C3 VDD A2 0.023177f
C4 VDD ZN 0.33173f
C5 VSS A3 0.07804f
C6 VSS A2 0.104901f
C7 VSS ZN 0.064021f
C8 VSS a_455_68# 0.006909f
C9 A3 VNW 0.148237f
C10 A2 VNW 0.121191f
C11 VNW ZN 0.034322f
C12 A1 VDD 0.022021f
C13 A1 VSS 0.084906f
C14 A1 VNW 0.12917f
C15 A3 A2 0.117566f
C16 A3 ZN 0.008403f
C17 A2 ZN 0.078589f
C18 a_455_68# A2 0.005127f
C19 a_455_68# ZN 0.002926f
C20 VSS a_271_68# 0.006038f
C21 A1 A2 0.133044f
C22 A1 ZN 0.384588f
C23 A1 a_455_68# 0.004981f
C24 VSS VDD 0.008734f
C25 VDD VNW 0.112537f
C26 A2 a_271_68# 0.004027f
C27 VSS VPW 0.307914f
C28 ZN VPW 0.133449f
C29 VDD VPW 0.241872f
C30 A1 VPW 0.287469f
C31 A2 VPW 0.25736f
C32 A3 VPW 0.326833f
C33 VNW VPW 1.48562f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW a_245_68#
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
C0 VSS a_245_68# 0.002295f
C1 ZN VSS 0.098328f
C2 A1 VSS 0.131667f
C3 A2 VDD 0.039698f
C4 VSS VNW 0.006174f
C5 ZN VDD 0.240333f
C6 A1 VDD 0.027485f
C7 ZN A2 0.038658f
C8 A1 A2 0.226398f
C9 VDD VNW 0.084263f
C10 A1 a_245_68# 0.008831f
C11 ZN A1 0.351362f
C12 VSS VDD 0.017706f
C13 A2 VNW 0.125396f
C14 A2 VSS 0.051087f
C15 ZN VNW 0.02653f
C16 A1 VNW 0.119756f
C17 VSS VPW 0.238729f
C18 ZN VPW 0.105772f
C19 VDD VPW 0.243067f
C20 A1 VPW 0.290957f
C21 A2 VPW 0.314823f
C22 VNW VPW 1.13753f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW a_255_603# a_67_603#
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VSS A2 0.025748f
C1 VNW a_67_603# 0.157241f
C2 VDD a_255_603# 0.005359f
C3 VDD A1 0.01431f
C4 a_255_603# A2 0.001961f
C5 A1 A2 0.062395f
C6 VNW Z 0.033884f
C7 VDD VNW 0.11771f
C8 Z a_67_603# 0.181586f
C9 VDD a_67_603# 0.307039f
C10 VSS A1 0.050738f
C11 VNW A2 0.216313f
C12 A2 a_67_603# 0.505374f
C13 VSS VNW 0.010039f
C14 VSS a_67_603# 0.250493f
C15 VDD Z 0.196046f
C16 Z A2 0.027598f
C17 VDD A2 0.147628f
C18 VSS Z 0.158265f
C19 VSS VDD 0.008648f
C20 VNW A1 0.220003f
C21 a_255_603# a_67_603# 0.007617f
C22 A1 a_67_603# 0.540888f
C23 VSS VPW 0.359722f
C24 Z VPW 0.102754f
C25 VDD VPW 0.233025f
C26 A2 VPW 0.313441f
C27 A1 VPW 0.39469f
C28 VNW VPW 1.65967f
C29 a_67_603# VPW 0.345683f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VNW VPW a_36_68# a_1612_497#
+ a_2124_68# a_244_497# a_2960_68# a_3368_68# a_2552_68# a_1164_497# a_716_497#
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
C0 A2 ZN 1.2828f
C1 VSS VNW 0.004483f
C2 a_36_68# A1 0.065645f
C3 a_2960_68# B 0.002626f
C4 a_1164_497# ZN 0.021094f
C5 VSS VDD 0.005699f
C6 A1 ZN 1.37575f
C7 a_3368_68# VSS 0.004815f
C8 a_1612_497# VDD 0.009792f
C9 VSS A2 0.060501f
C10 a_36_68# B 1.37417f
C11 A2 a_1612_497# 0.010709f
C12 ZN B 0.426118f
C13 C VNW 0.636287f
C14 a_244_497# ZN 0.009475f
C15 a_36_68# a_2960_68# 0.009506f
C16 a_716_497# ZN 0.027752f
C17 a_36_68# ZN 1.98502f
C18 C VDD 0.095093f
C19 VSS A1 0.060963f
C20 VSS B 0.072527f
C21 a_36_68# a_2124_68# 0.012118f
C22 VSS a_2960_68# 0.002422f
C23 VNW VDD 0.366897f
C24 VSS a_36_68# 3.64719f
C25 B a_2552_68# 0.002588f
C26 A2 VNW 0.590323f
C27 VSS ZN 0.006216f
C28 ZN a_1612_497# 0.024559f
C29 C B 1.73339f
C30 A2 VDD 0.15752f
C31 a_36_68# a_2552_68# 0.009506f
C32 VSS a_2124_68# 0.004133f
C33 a_36_68# C 0.105844f
C34 A1 VNW 0.51833f
C35 C ZN 0.514613f
C36 VNW B 0.600992f
C37 a_1164_497# VDD 0.008664f
C38 A1 VDD 0.078657f
C39 a_1164_497# A2 0.009095f
C40 A1 A2 1.73987f
C41 B VDD 0.100578f
C42 VSS a_2552_68# 0.002422f
C43 A2 B 0.037299f
C44 a_36_68# VNW 0.004654f
C45 ZN VNW 0.056895f
C46 VSS C 0.092809f
C47 a_244_497# VDD 0.020528f
C48 a_244_497# A2 0.01347f
C49 a_716_497# VDD 0.008599f
C50 a_36_68# VDD 0.021485f
C51 a_3368_68# a_36_68# 0.007478f
C52 a_716_497# A2 0.00653f
C53 a_36_68# A2 0.108262f
C54 ZN VDD 2.06829f
C55 VSS VPW 1.08055f
C56 ZN VPW 0.051826f
C57 VDD VPW 0.846798f
C58 C VPW 1.06351f
C59 B VPW 1.11555f
C60 A1 VPW 1.1956f
C61 A2 VPW 1.16629f
C62 VNW VPW 5.892971f
C63 a_36_68# VPW 0.063181f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW a_36_160#
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
C0 I VSS 0.178818f
C1 VNW VSS 0.00834f
C2 I a_36_160# 0.564508f
C3 VNW a_36_160# 0.302514f
C4 VSS a_36_160# 0.114407f
C5 Z I 0.016176f
C6 Z VNW 0.021185f
C7 I VDD 0.028233f
C8 VDD VNW 0.111398f
C9 Z VSS 0.111496f
C10 VDD VSS 0.01316f
C11 Z a_36_160# 0.426617f
C12 VDD a_36_160# 0.31851f
C13 Z VDD 0.161733f
C14 I VNW 0.1633f
C15 VSS VPW 0.397291f
C16 Z VPW 0.097163f
C17 VDD VPW 0.238155f
C18 I VPW 0.333888f
C19 VNW VPW 1.65967f
C20 a_36_160# VPW 0.696445f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW a_1380_472# a_36_472#
+ a_932_472# a_572_375# a_124_375# a_1468_375# a_1020_375# a_484_472#
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_1020_375# a_932_472# 0.285629f
C1 VNW a_1380_472# 0.024396f
C2 a_124_375# VSS 0.134699f
C3 a_484_472# VSS 0.148077f
C4 a_36_472# VSS 0.147381f
C5 VNW VSS 0.017643f
C6 a_572_375# VSS 0.134699f
C7 a_1468_375# VNW 0.18122f
C8 a_1020_375# VNW 0.181468f
C9 a_572_375# a_1020_375# 0.012552f
C10 VDD a_1380_472# 0.179463f
C11 a_484_472# a_932_472# 0.013276f
C12 a_932_472# VNW 0.024018f
C13 a_572_375# a_932_472# 0.086905f
C14 a_484_472# a_124_375# 0.086905f
C15 a_36_472# a_124_375# 0.285629f
C16 VNW a_124_375# 0.180172f
C17 VDD VSS 0.026369f
C18 a_572_375# a_124_375# 0.012552f
C19 a_1468_375# VDD 0.129266f
C20 a_1020_375# VDD 0.129962f
C21 a_484_472# a_36_472# 0.013276f
C22 a_484_472# VNW 0.024018f
C23 a_36_472# VNW 0.025611f
C24 a_484_472# a_572_375# 0.285629f
C25 a_1380_472# VSS 0.144845f
C26 VDD a_932_472# 0.179463f
C27 a_1468_375# a_1380_472# 0.285629f
C28 a_572_375# VNW 0.181468f
C29 a_1020_375# a_1380_472# 0.086905f
C30 a_932_472# a_1380_472# 0.013276f
C31 VDD a_124_375# 0.12673f
C32 a_484_472# VDD 0.179463f
C33 a_1468_375# VSS 0.082091f
C34 a_1020_375# VSS 0.134699f
C35 a_36_472# VDD 0.093681f
C36 a_1468_375# a_1020_375# 0.012552f
C37 VDD VNW 0.217349f
C38 a_572_375# VDD 0.129962f
C39 a_932_472# VSS 0.148077f
C40 VSS VPW 0.642184f
C41 VDD VPW 0.493288f
C42 VNW VPW 3.05206f
C43 a_1380_472# VPW 0.345058f
C44 a_932_472# VPW 0.33241f
C45 a_484_472# VPW 0.33241f
C46 a_36_472# VPW 0.404746f
C47 a_1468_375# VPW 0.233029f
C48 a_1020_375# VPW 0.171606f
C49 a_572_375# VPW 0.171606f
C50 a_124_375# VPW 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW a_36_68#
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 Z VDD 0.172592f
C1 a_36_68# VNW 0.296832f
C2 VSS VNW 0.009972f
C3 VSS a_36_68# 0.156367f
C4 VNW I 0.133333f
C5 a_36_68# I 0.731677f
C6 VDD VNW 0.114912f
C7 Z VNW 0.023138f
C8 VSS I 0.128735f
C9 a_36_68# VDD 0.271105f
C10 a_36_68# Z 0.432914f
C11 VSS VDD 0.014283f
C12 VSS Z 0.133443f
C13 VDD I 0.029139f
C14 Z I 0.018906f
C15 VSS VPW 0.338876f
C16 Z VPW 0.103236f
C17 VDD VPW 0.234026f
C18 I VPW 0.298844f
C19 VNW VPW 1.65967f
C20 a_36_68# VPW 0.69549f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW a_848_380# a_1084_68#
+ a_124_24# a_1152_472# a_692_472#
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
C0 VSS Z 0.129676f
C1 a_124_24# I1 0.564972f
C2 VDD I1 0.227359f
C3 VNW Z 0.020389f
C4 S a_692_472# 0.002582f
C5 I0 a_848_380# 0.082224f
C6 VSS a_848_380# 0.130064f
C7 S a_124_24# 0.245829f
C8 VDD S 0.056165f
C9 VSS I1 0.026996f
C10 a_848_380# a_1152_472# 0.007362f
C11 a_124_24# a_692_472# 0.033243f
C12 VDD a_692_472# 0.009663f
C13 VNW a_848_380# 0.174516f
C14 VNW I1 0.127749f
C15 VDD a_124_24# 0.309232f
C16 I0 S 0.533789f
C17 VSS S 0.081531f
C18 S VNW 0.253706f
C19 I0 a_124_24# 0.004772f
C20 VSS a_124_24# 0.501844f
C21 VDD I0 0.028914f
C22 Z I1 0.027341f
C23 VSS VDD 0.028952f
C24 a_124_24# a_1152_472# 0.00128f
C25 VDD a_1152_472# 0.00645f
C26 VNW a_124_24# 0.277682f
C27 S a_1084_68# 0.001644f
C28 VDD VNW 0.182986f
C29 a_124_24# a_692_68# 0.006853f
C30 a_124_24# a_1084_68# 0.002839f
C31 a_848_380# I1 0.013444f
C32 VSS I0 0.124513f
C33 I0 VNW 0.103064f
C34 VSS VNW 0.009598f
C35 a_124_24# Z 0.219295f
C36 VDD Z 0.20273f
C37 S a_848_380# 0.754833f
C38 VSS a_692_68# 0.001982f
C39 I0 a_1084_68# 0.00492f
C40 VSS a_1084_68# 0.009508f
C41 a_692_472# a_848_380# 0.003985f
C42 S I1 0.042269f
C43 a_692_472# I1 0.001219f
C44 a_124_24# a_848_380# 0.302602f
C45 VDD a_848_380# 0.319708f
C46 VSS VPW 0.565512f
C47 Z VPW 0.047467f
C48 VDD VPW 0.424967f
C49 I0 VPW 0.267152f
C50 S VPW 0.549493f
C51 I1 VPW 0.247562f
C52 VNW VPW 2.87801f
C53 a_848_380# VPW 0.40208f
C54 a_124_24# VPW 0.591898f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW a_36_68# a_244_472#
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 A1 A2 0.038725f
C1 VNW B 0.163023f
C2 ZN a_244_472# 0.014146f
C3 A1 VSS 0.090903f
C4 a_36_68# VDD 0.753239f
C5 VNW a_36_68# 0.038286f
C6 A1 B 0.034707f
C7 a_36_68# ZN 0.56857f
C8 VNW VDD 0.117098f
C9 ZN VDD 0.006004f
C10 VNW ZN 0.011308f
C11 A2 VSS 0.083821f
C12 A1 a_36_68# 0.292244f
C13 A1 VDD 0.014914f
C14 A1 VNW 0.117811f
C15 A1 ZN 0.496662f
C16 B VSS 0.198567f
C17 a_36_68# A2 0.489122f
C18 A2 VDD 0.017122f
C19 VNW A2 0.122386f
C20 a_36_68# VSS 0.117681f
C21 ZN A2 0.400775f
C22 VDD VSS 0.004855f
C23 a_36_68# B 0.389329f
C24 a_36_68# a_244_472# 0.013419f
C25 VNW VSS 0.0064f
C26 B VDD 0.07579f
C27 ZN VSS 0.088946f
C28 VDD a_244_472# 0.004051f
C29 VSS VPW 0.342662f
C30 ZN VPW 0.011384f
C31 VDD VPW 0.256635f
C32 B VPW 0.339176f
C33 A1 VPW 0.256004f
C34 A2 VPW 0.28395f
C35 VNW VPW 1.65967f
C36 a_36_68# VPW 0.112263f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW a_224_552#
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
C0 VNW Z 0.027266f
C1 VNW VSS 0.009226f
C2 VNW VDD 0.176912f
C3 VNW I 0.376531f
C4 a_224_552# Z 1.17071f
C5 a_224_552# VSS 0.331404f
C6 a_224_552# VDD 0.347549f
C7 I a_224_552# 0.421587f
C8 VSS Z 0.275062f
C9 VDD Z 0.356369f
C10 I Z 0.002319f
C11 VSS VDD 0.030201f
C12 I VSS 0.061715f
C13 VNW a_224_552# 0.5926f
C14 I VDD 0.069894f
C15 VSS VPW 0.628617f
C16 Z VPW 0.102362f
C17 VDD VPW 0.415149f
C18 I VPW 0.471574f
C19 VNW VPW 2.70396f
C20 a_224_552# VPW 1.31114f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW a_234_472# a_672_472#
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 VDD a_672_472# 0.005379f
C1 a_234_472# ZN 0.003154f
C2 A2 a_672_472# 0.0147f
C3 A1 ZN 0.274601f
C4 VDD ZN 0.517479f
C5 VSS ZN 0.460527f
C6 A2 ZN 0.509001f
C7 VNW ZN 0.03148f
C8 a_234_472# VDD 0.0121f
C9 a_234_472# A2 0.018681f
C10 VDD A1 0.037494f
C11 a_672_472# ZN 0.023475f
C12 VSS A1 0.052992f
C13 VDD VSS 0.023993f
C14 A2 A1 0.636124f
C15 VNW A1 0.25895f
C16 VDD A2 0.13595f
C17 VNW VDD 0.137685f
C18 VSS A2 0.07211f
C19 VNW VSS 0.010681f
C20 VNW A2 0.275679f
C21 VSS VPW 0.451405f
C22 ZN VPW 0.138491f
C23 VDD VPW 0.322159f
C24 A1 VPW 0.557317f
C25 A2 VPW 0.617688f
C26 VNW VPW 2.00777f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_448_472# a_244_472#
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
C0 VSS ZN 0.283414f
C1 VNW VDD 0.11801f
C2 VSS VDD 0.01583f
C3 A2 A3 0.416588f
C4 A2 A1 0.145555f
C5 A2 a_244_472# 0.003952f
C6 VNW A3 0.136756f
C7 VNW A1 0.127941f
C8 VSS A3 0.058214f
C9 VSS A1 0.025677f
C10 ZN a_448_472# 0.006209f
C11 VDD a_448_472# 0.013539f
C12 ZN VDD 0.116419f
C13 VNW A2 0.116878f
C14 VSS A2 0.027728f
C15 A1 a_448_472# 0.012619f
C16 ZN A3 0.035547f
C17 ZN A1 0.499849f
C18 VDD A3 0.201466f
C19 VDD A1 0.095023f
C20 ZN a_244_472# 0.001803f
C21 a_244_472# VDD 0.006513f
C22 VSS VNW 0.008407f
C23 a_244_472# A3 0.019089f
C24 A2 a_448_472# 0.012315f
C25 ZN A2 0.096665f
C26 A2 VDD 0.09496f
C27 ZN VNW 0.040402f
C28 VSS VPW 0.367618f
C29 ZN VPW 0.134331f
C30 VDD VPW 0.264623f
C31 A1 VPW 0.311038f
C32 A2 VPW 0.285534f
C33 A3 VPW 0.334053f
C34 VNW VPW 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VNW VPW a_36_68# a_1732_68#
+ a_244_68# a_1100_68# a_1528_68# a_672_68#
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
C0 a_244_68# a_36_68# 0.009768f
C1 a_1732_68# ZN 0.002613f
C2 A2 A1 0.077487f
C3 A3 A1 0.001696f
C4 A2 ZN 1.77619f
C5 A3 ZN 0.150755f
C6 VSS a_672_68# 0.003125f
C7 a_36_68# VSS 2.77545f
C8 VDD A2 0.124271f
C9 VDD A3 0.107959f
C10 a_36_68# a_1528_68# 0.012072f
C11 A2 VNW 0.630933f
C12 A1 VSS 0.065524f
C13 A3 VNW 0.599629f
C14 ZN VSS 0.00864f
C15 a_36_68# a_672_68# 0.012389f
C16 VDD VSS 0.004708f
C17 a_1100_68# A3 0.003385f
C18 A3 A2 1.65768f
C19 VSS VNW 0.003704f
C20 a_36_68# A1 0.118844f
C21 a_36_68# ZN 0.885472f
C22 VDD a_36_68# 0.029088f
C23 a_1100_68# VSS 0.003125f
C24 a_1732_68# VSS 0.002237f
C25 A1 ZN 1.266f
C26 A2 VSS 0.070822f
C27 A3 VSS 0.09506f
C28 a_36_68# VNW 0.007741f
C29 VDD A1 0.115489f
C30 VDD ZN 1.57207f
C31 a_244_68# VSS 0.006268f
C32 a_1100_68# a_36_68# 0.012396f
C33 a_1732_68# a_36_68# 0.011094f
C34 A1 VNW 0.700258f
C35 ZN VNW 0.095885f
C36 A3 a_672_68# 0.003442f
C37 a_36_68# A2 0.223434f
C38 A3 a_36_68# 1.03106f
C39 VDD VNW 0.292073f
C40 VSS a_1528_68# 0.003775f
C41 VSS VPW 0.861061f
C42 ZN VPW 0.103891f
C43 VDD VPW 0.701563f
C44 A1 VPW 1.27704f
C45 A3 VPW 1.11693f
C46 A2 VPW 1.08692f
C47 VNW VPW 4.73584f
C48 a_36_68# VPW 0.061249f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW a_36_159#
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
C0 VSS Z 0.102819f
C1 a_36_159# A1 0.377122f
C2 VNW a_36_159# 0.162496f
C3 a_36_159# Z 0.215269f
C4 A1 A2 0.061431f
C5 a_36_159# VSS 0.244357f
C6 a_244_159# VSS 0.001449f
C7 VDD A1 0.04397f
C8 VNW A2 0.20463f
C9 VNW VDD 0.125609f
C10 A2 Z 0.020174f
C11 VDD Z 0.158212f
C12 a_244_159# a_36_159# 0.003343f
C13 VSS A2 0.011099f
C14 VSS VDD 0.014131f
C15 a_36_159# A2 0.472781f
C16 a_36_159# VDD 0.130189f
C17 VNW A1 0.206765f
C18 VNW Z 0.032842f
C19 VDD A2 0.184025f
C20 VSS A1 0.010276f
C21 VNW VSS 0.007925f
C22 VSS VPW 0.35312f
C23 Z VPW 0.096476f
C24 VDD VPW 0.251252f
C25 A2 VPW 0.262264f
C26 A1 VPW 0.321274f
C27 VNW VPW 1.65967f
C28 a_36_159# VPW 0.374116f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VNW VPW a_2590_472#
+ a_170_472# a_1602_69# a_786_69# a_3126_472# a_1194_69# a_3662_472# a_2034_472# a_358_69#
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VPW nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VPW nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VPW nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
C0 VDD A2 0.052548f
C1 a_3126_472# a_170_472# 0.01307f
C2 a_1602_69# ZN 0.008113f
C3 B a_3662_472# 0.007338f
C4 VNW C 0.61926f
C5 VSS a_170_472# 0.00801f
C6 VSS A1 0.087217f
C7 VNW ZN 0.045695f
C8 a_3126_472# VDD 0.00779f
C9 B C 1.34577f
C10 A1 a_170_472# 0.0698f
C11 a_786_69# ZN 0.008749f
C12 VSS VDD 0.016824f
C13 B ZN 0.231932f
C14 VDD a_170_472# 2.96356f
C15 VDD A1 0.051939f
C16 VSS a_358_69# 0.005318f
C17 A1 a_358_69# 0.001641f
C18 B a_2590_472# 0.007345f
C19 A2 ZN 1.83822f
C20 VNW B 0.617219f
C21 a_1194_69# ZN 0.00847f
C22 B a_2034_472# 0.008709f
C23 a_170_472# a_3662_472# 0.013628f
C24 VSS C 0.088883f
C25 VNW A2 0.513788f
C26 VSS ZN 1.77446f
C27 C a_170_472# 0.075372f
C28 VDD a_3662_472# 0.007223f
C29 A1 C 0.001754f
C30 B A2 0.05388f
C31 a_170_472# ZN 0.818521f
C32 A1 ZN 1.40746f
C33 VDD C 0.089678f
C34 VDD ZN 0.008843f
C35 VSS a_1602_69# 0.005669f
C36 a_358_69# ZN 0.011344f
C37 a_170_472# a_2590_472# 0.013379f
C38 VNW VSS 0.012025f
C39 a_3126_472# B 0.007345f
C40 VSS a_786_69# 0.003966f
C41 VNW a_170_472# 0.018375f
C42 VSS B 0.119454f
C43 VNW A1 0.480244f
C44 VDD a_2590_472# 0.007681f
C45 B a_170_472# 2.12702f
C46 a_786_69# A1 0.001203f
C47 B A1 0.001644f
C48 VNW VDD 0.393677f
C49 a_170_472# a_2034_472# 0.020753f
C50 B VDD 0.110239f
C51 VDD a_2034_472# 0.008673f
C52 VSS A2 0.104058f
C53 A2 a_170_472# 0.109943f
C54 a_1194_69# VSS 0.005069f
C55 A2 A1 1.72617f
C56 C ZN 1.79111f
C57 VSS VPW 1.33264f
C58 VDD VPW 0.809429f
C59 ZN VPW 0.171181f
C60 C VPW 1.26656f
C61 B VPW 1.19887f
C62 A1 VPW 1.12703f
C63 A2 VPW 1.09165f
C64 VNW VPW 6.53302f
C65 a_170_472# VPW 0.077257f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW a_1792_472# a_224_472#
+ a_1568_472# a_36_472# a_1120_472# a_672_472#
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
C0 a_1568_472# A1 0.002055f
C1 A2 A1 0.085569f
C2 a_1792_472# A1 0.006624f
C3 a_1120_472# A2 0.002647f
C4 ZN A2 0.250963f
C5 ZN a_1792_472# 0.004144f
C6 a_672_472# VDD 0.01105f
C7 VDD VSS 0.012739f
C8 a_224_472# a_36_472# 0.01823f
C9 a_36_472# VNW 0.031928f
C10 a_36_472# A3 0.100976f
C11 VDD A1 0.054887f
C12 VNW A3 0.478769f
C13 a_1120_472# VDD 0.011157f
C14 VSS A1 0.115774f
C15 ZN VDD 0.005367f
C16 ZN VSS 2.18568f
C17 a_224_472# A2 0.002647f
C18 a_1568_472# a_36_472# 0.025433f
C19 A2 a_36_472# 0.993181f
C20 A2 VNW 0.539636f
C21 a_1792_472# a_36_472# 0.022081f
C22 A2 A3 1.6562f
C23 ZN A1 1.56829f
C24 a_224_472# VDD 0.010911f
C25 A2 a_1568_472# 0.004974f
C26 a_36_472# VDD 1.90933f
C27 VDD VNW 0.286001f
C28 VDD A3 0.09322f
C29 a_672_472# a_36_472# 0.01823f
C30 a_36_472# VSS 0.020716f
C31 VNW VSS 0.009996f
C32 VSS A3 0.10353f
C33 a_36_472# A1 0.174868f
C34 VNW A1 0.520086f
C35 a_1568_472# VDD 0.005385f
C36 a_1120_472# a_36_472# 0.01951f
C37 A1 A3 0.008795f
C38 A2 VDD 0.082489f
C39 a_1792_472# VDD 0.002998f
C40 ZN a_36_472# 0.362263f
C41 ZN VNW 0.046016f
C42 a_672_472# A2 0.002647f
C43 ZN A3 1.42151f
C44 A2 VSS 0.128956f
C45 VSS VPW 0.918064f
C46 ZN VPW 0.159858f
C47 VDD VPW 0.61695f
C48 A1 VPW 1.35739f
C49 A3 VPW 1.33073f
C50 A2 VPW 1.29013f
C51 VNW VPW 4.79254f
C52 a_36_472# VPW 0.137725f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW a_468_472# a_244_472#
+ a_1130_472# a_906_472#
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 VSS ZN 1.3936f
C1 A3 a_1130_472# 0.016495f
C2 A3 VNW 0.28584f
C3 ZN a_468_472# 0.015602f
C4 A1 VSS 0.044587f
C5 VDD a_1130_472# 0.011629f
C6 VDD VNW 0.178574f
C7 A3 A2 0.624599f
C8 A3 a_906_472# 0.017829f
C9 a_244_472# ZN 0.019831f
C10 VDD A2 0.038421f
C11 VDD a_906_472# 0.011614f
C12 A2 VNW 0.241313f
C13 A3 ZN 1.03634f
C14 A3 A1 0.292395f
C15 VDD ZN 0.579119f
C16 a_1130_472# ZN 0.001342f
C17 VNW ZN 0.031771f
C18 VDD A1 0.038139f
C19 A3 VSS 0.0525f
C20 A1 VNW 0.254404f
C21 A3 a_468_472# 0.010018f
C22 A2 ZN 0.694728f
C23 VDD VSS 0.009106f
C24 a_906_472# ZN 0.002855f
C25 VSS VNW 0.007164f
C26 A2 A1 0.570018f
C27 VDD a_468_472# 0.00502f
C28 A3 a_244_472# 0.010666f
C29 A2 VSS 0.043139f
C30 A1 ZN 0.084783f
C31 VDD a_244_472# 0.00632f
C32 VDD A3 0.178286f
C33 VSS VPW 0.509614f
C34 ZN VPW 0.172636f
C35 VDD VPW 0.441158f
C36 A1 VPW 0.622214f
C37 A2 VPW 0.627317f
C38 A3 VPW 0.692739f
C39 VNW VPW 2.70396f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VNW VPW a_1492_488#
+ a_244_68# a_1044_488# a_636_68# a_36_488#
X0 VSS B ZN VPW nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VPW nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VPW nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VPW nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
C0 B C 0.560408f
C1 VSS B 0.089442f
C2 a_244_68# ZN 0.001328f
C3 A1 VSS 0.090485f
C4 a_36_488# VNW 0.010653f
C5 ZN VNW 0.028815f
C6 A2 a_36_488# 0.076279f
C7 VDD VNW 0.191798f
C8 A2 ZN 0.752866f
C9 A2 VDD 0.02614f
C10 B a_1492_488# 0.007233f
C11 VSS C 0.05406f
C12 a_36_488# B 0.80489f
C13 B ZN 0.413891f
C14 VDD B 0.04259f
C15 A1 a_36_488# 0.031215f
C16 A1 ZN 0.372797f
C17 A1 VDD 0.026261f
C18 a_1044_488# a_36_488# 0.018358f
C19 A2 VNW 0.280457f
C20 a_1044_488# VDD 0.004195f
C21 A1 a_244_68# 0.003444f
C22 VSS a_636_68# 0.002222f
C23 a_36_488# C 0.041645f
C24 B VNW 0.298561f
C25 VSS a_36_488# 0.005331f
C26 ZN C 0.191881f
C27 VSS ZN 0.708286f
C28 VDD C 0.040747f
C29 A2 B 0.036672f
C30 VSS VDD 0.009527f
C31 A1 VNW 0.25321f
C32 A1 A2 0.652956f
C33 VSS a_244_68# 0.004878f
C34 a_36_488# a_1492_488# 0.017313f
C35 VDD a_1492_488# 0.00909f
C36 a_636_68# ZN 0.00593f
C37 C VNW 0.268332f
C38 VSS VNW 0.008434f
C39 a_1044_488# B 0.012375f
C40 a_36_488# ZN 0.459425f
C41 VSS A2 0.077665f
C42 a_36_488# VDD 1.67897f
C43 VDD ZN 0.004894f
C44 VSS VPW 0.653933f
C45 VDD VPW 0.406726f
C46 ZN VPW 0.089692f
C47 C VPW 0.626227f
C48 B VPW 0.654892f
C49 A1 VPW 0.552174f
C50 A2 VPW 0.559992f
C51 VNW VPW 3.2261f
C52 a_36_488# VPW 0.101145f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VNW VPW a_244_524# a_2215_68#
+ a_56_524# a_718_524# a_728_93# a_1936_472# a_1336_472#
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
C0 VSS VDD 0.013872f
C1 A2 a_56_524# 0.908796f
C2 VDD VNW 0.360391f
C3 a_1936_472# VDD 0.595117f
C4 VDD Z 0.01058f
C5 a_728_93# a_56_524# 0.016741f
C6 a_1524_472# a_728_93# 0.007139f
C7 A1 a_56_524# 0.569057f
C8 VDD A2 0.208821f
C9 VDD a_728_93# 0.575073f
C10 a_1336_472# a_1524_472# 0.001046f
C11 A1 VDD 0.018915f
C12 a_2215_68# VSS 0.004309f
C13 a_1336_472# VDD 0.033982f
C14 a_718_524# VNW 0.020055f
C15 a_2215_68# Z 0.008507f
C16 A2 a_244_524# 0.004824f
C17 a_718_524# A2 0.107911f
C18 a_718_524# a_728_93# 0.329834f
C19 A1 a_718_524# 0.026418f
C20 A3 VSS 0.056027f
C21 VDD a_56_524# 0.049641f
C22 A3 VNW 0.268193f
C23 a_1936_472# A3 0.018144f
C24 A3 Z 0.259021f
C25 VSS VNW 0.007756f
C26 VSS Z 0.277351f
C27 a_1936_472# VNW 0.004015f
C28 VNW Z 0.028011f
C29 A3 a_728_93# 0.720358f
C30 a_1936_472# Z 0.337902f
C31 VSS A2 0.047538f
C32 A2 VNW 0.369075f
C33 VSS a_728_93# 0.709567f
C34 a_728_93# VNW 0.346549f
C35 a_1336_472# A3 0.490376f
C36 a_718_524# a_56_524# 0.009198f
C37 a_1936_472# a_728_93# 0.105997f
C38 A1 VSS 0.139902f
C39 a_728_93# Z 0.402606f
C40 A1 VNW 0.293766f
C41 a_728_93# a_952_93# 0.00421f
C42 VDD a_244_524# 0.004322f
C43 A2 a_728_93# 0.416172f
C44 a_1336_472# VSS 0.326133f
C45 VDD a_718_524# 0.554575f
C46 a_1336_472# VNW 0.144065f
C47 a_1936_472# a_1336_472# 0.004622f
C48 A1 A2 0.321942f
C49 a_1336_472# Z 0.021039f
C50 A1 a_728_93# 0.12992f
C51 a_1336_472# A2 0.001757f
C52 a_1336_472# a_728_93# 0.62718f
C53 A3 VDD 0.028848f
C54 VSS a_56_524# 0.214447f
C55 VNW a_56_524# 0.188846f
C56 VSS VPW 0.861752f
C57 Z VPW 0.085787f
C58 A1 VPW 0.602985f
C59 A2 VPW 0.640744f
C60 VDD VPW 0.543474f
C61 A3 VPW 0.593976f
C62 VNW VPW 4.270391f
C63 a_1936_472# VPW 0.009918f
C64 a_718_524# VPW 0.005143f
C65 a_56_524# VPW 0.41096f
C66 a_728_93# VPW 0.654825f
C67 a_1336_472# VPW 0.316639f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VNW VPW a_652_68# a_244_68#
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
C0 A2 VNW 0.277885f
C1 a_244_68# A1 0.004867f
C2 VSS VNW 0.008805f
C3 A2 VSS 0.057292f
C4 ZN A1 0.363066f
C5 ZN VDD 0.409997f
C6 VNW A1 0.232646f
C7 A2 A1 0.708017f
C8 VSS A1 0.115936f
C9 VNW VDD 0.123338f
C10 A2 VDD 0.070487f
C11 ZN a_244_68# 0.001926f
C12 VSS VDD 0.020712f
C13 ZN a_652_68# 0.008436f
C14 A1 VDD 0.050088f
C15 VSS a_244_68# 0.006834f
C16 ZN VNW 0.033841f
C17 A2 ZN 0.891023f
C18 VSS a_652_68# 0.003855f
C19 ZN VSS 0.2597f
C20 VSS VPW 0.385688f
C21 ZN VPW 0.120217f
C22 VDD VPW 0.305683f
C23 A1 VPW 0.522064f
C24 A2 VPW 0.568932f
C25 VNW VPW 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VNW VPW a_36_68# a_1612_497#
+ a_692_497# a_1388_497# a_960_497#
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
C0 a_692_497# A3 0.019827f
C1 A1 a_36_68# 0.158235f
C2 a_960_497# A3 0.014254f
C3 a_692_497# ZN 0.018589f
C4 a_960_497# ZN 0.012124f
C5 a_692_497# VDD 0.00542f
C6 a_36_68# A3 0.036843f
C7 A1 A2 0.703324f
C8 a_960_497# VDD 0.003264f
C9 ZN a_36_68# 1.49222f
C10 a_1612_497# A2 0.006056f
C11 A2 A3 1.11591f
C12 a_36_68# B 0.184521f
C13 a_36_68# VDD 0.001802f
C14 ZN A2 0.152712f
C15 VDD A2 0.030601f
C16 a_36_68# VNW 0.001442f
C17 VNW A2 0.281901f
C18 A1 VSS 0.032188f
C19 VSS A3 0.03178f
C20 VSS ZN 0.006088f
C21 a_692_497# A2 0.001398f
C22 VSS B 0.047409f
C23 VSS VDD 0.010407f
C24 a_960_497# A2 0.003506f
C25 a_36_68# A2 0.032025f
C26 VSS VNW 0.008187f
C27 a_1388_497# A3 0.02079f
C28 ZN a_1388_497# 0.001168f
C29 a_1388_497# VDD 0.005409f
C30 VSS a_36_68# 2.0408f
C31 VSS A2 0.030287f
C32 A1 a_1612_497# 0.003158f
C33 A1 A3 0.206693f
C34 A1 ZN 0.619225f
C35 a_1612_497# A3 0.030605f
C36 A1 VDD 0.091309f
C37 ZN A3 1.02771f
C38 a_1388_497# A2 0.008156f
C39 a_1612_497# VDD 0.009412f
C40 B A3 0.036798f
C41 VDD A3 0.555327f
C42 A1 VNW 0.279057f
C43 ZN B 0.244028f
C44 ZN VDD 1.08837f
C45 VDD B 0.119783f
C46 VNW A3 0.297068f
C47 ZN VNW 0.025446f
C48 VNW B 0.309147f
C49 VNW VDD 0.248379f
C50 VSS VPW 0.663038f
C51 ZN VPW 0.080495f
C52 VDD VPW 0.512998f
C53 A1 VPW 0.643779f
C54 A2 VPW 0.561227f
C55 A3 VPW 0.573818f
C56 B VPW 0.585725f
C57 VNW VPW 3.48825f
C58 a_36_68# VPW 0.048026f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VNW VPW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_2248_156#
+ a_2560_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VPW nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VPW nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 a_1308_423# VDD 0.094185f
C1 VNW a_36_151# 1.28833f
C2 VDD a_36_151# 0.417101f
C3 a_1000_472# VNW 0.241357f
C4 a_1308_423# a_448_472# 0.882105f
C5 VDD a_1000_472# 0.119211f
C6 Q VNW 0.026596f
C7 a_1308_423# a_2248_156# 0.056721f
C8 VNW a_796_472# 0.010232f
C9 Q VDD 0.260055f
C10 a_448_472# a_36_151# 0.536965f
C11 RN VNW 0.304626f
C12 a_2248_156# a_36_151# 0.042802f
C13 a_2665_112# a_3041_156# 0.001841f
C14 VDD RN 0.035003f
C15 a_1000_472# a_448_472# 0.361958f
C16 CLK a_36_151# 0.669598f
C17 a_1308_423# VSS 0.013866f
C18 a_2248_156# a_1000_472# 0.001232f
C19 a_796_472# a_448_472# 0.401636f
C20 Q a_2248_156# 0.013765f
C21 VSS a_36_151# 0.291264f
C22 a_2560_156# a_36_151# 0.003674f
C23 RN a_448_472# 0.078731f
C24 a_2248_156# RN 0.080362f
C25 VSS a_1000_472# 0.04356f
C26 a_1308_423# a_1204_472# 0.026665f
C27 Q VSS 0.170514f
C28 VSS a_796_472# 0.05215f
C29 VDD VNW 0.546785f
C30 a_1204_472# a_36_151# 0.006996f
C31 VSS RN 0.436942f
C32 RN a_2560_156# 0.038779f
C33 a_1456_156# a_448_472# 0.00227f
C34 a_1204_472# a_1000_472# 0.66083f
C35 a_1288_156# a_448_472# 0.002067f
C36 D a_36_151# 0.094113f
C37 VNW a_448_472# 0.341284f
C38 VDD a_448_472# 0.456269f
C39 a_2248_156# VNW 0.181292f
C40 CLK VNW 0.137037f
C41 RN a_1204_472# 0.021039f
C42 a_2248_156# VDD 1.12036f
C43 VSS a_1456_156# 0.001901f
C44 a_796_472# D 0.082858f
C45 VDD CLK 0.02303f
C46 VSS a_1288_156# 0.001702f
C47 VSS VNW 0.012596f
C48 a_2560_156# VNW 0.019282f
C49 a_2248_156# a_448_472# 0.510371f
C50 a_2665_112# a_36_151# 0.019033f
C51 VSS VDD 0.02167f
C52 VDD a_2560_156# 0.00302f
C53 CLK a_448_472# 0.002757f
C54 RN a_3041_156# 0.014924f
C55 Q a_2665_112# 0.263315f
C56 a_1204_472# VNW 0.016269f
C57 VSS a_448_472# 1.20207f
C58 a_2560_156# a_448_472# 0.277491f
C59 VDD a_1204_472# 0.282626f
C60 VSS a_2248_156# 0.030372f
C61 a_2248_156# a_2560_156# 0.119687f
C62 a_2665_112# RN 0.322698f
C63 VSS CLK 0.021952f
C64 VNW D 0.128231f
C65 VDD D 0.009367f
C66 a_1204_472# a_448_472# 0.008996f
C67 VSS a_2560_156# 0.128503f
C68 a_1308_423# a_36_151# 0.05539f
C69 a_448_472# D 0.328788f
C70 a_1308_423# a_1000_472# 0.934191f
C71 a_2665_112# VNW 0.486803f
C72 a_2665_112# VDD 0.152571f
C73 a_1000_472# a_36_151# 0.08126f
C74 VSS D 0.064618f
C75 a_1308_423# RN 0.079294f
C76 a_796_472# a_36_151# 0.011851f
C77 a_2665_112# a_448_472# 0.020455f
C78 VSS a_3041_156# 0.004935f
C79 a_1000_472# a_796_472# 0.048436f
C80 RN a_36_151# 0.080119f
C81 a_2248_156# a_2665_112# 0.63615f
C82 RN a_1000_472# 0.0832f
C83 VSS a_2665_112# 0.21484f
C84 a_2665_112# a_2560_156# 0.116229f
C85 a_1308_423# VNW 0.149014f
C86 Q VPW 0.061347f
C87 VSS VPW 1.33519f
C88 RN VPW 1.37098f
C89 D VPW 0.253406f
C90 VDD VPW 0.859994f
C91 CLK VPW 0.291241f
C92 VNW VPW 6.48579f
C93 a_2560_156# VPW 0.016968f
C94 a_2665_112# VPW 0.91969f
C95 a_2248_156# VPW 0.30886f
C96 a_1204_472# VPW 0.012971f
C97 a_1000_472# VPW 0.291735f
C98 a_796_472# VPW 0.023206f
C99 a_1308_423# VPW 0.279043f
C100 a_448_472# VPW 0.684413f
C101 a_36_151# VPW 1.43587f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW a_438_68#
+ a_244_68# a_1254_68# a_1060_68# a_632_68# a_1458_68#
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
C0 ZN A3 0.881941f
C1 A4 VSS 0.056757f
C2 A4 VNW 0.388525f
C3 a_632_68# VSS 0.005832f
C4 A4 VDD 0.047422f
C5 A4 A3 0.297972f
C6 A4 ZN 1.94271f
C7 VSS a_244_68# 0.007139f
C8 a_632_68# A3 0.0083f
C9 A1 A2 0.516286f
C10 VSS a_1458_68# 0.002548f
C11 a_632_68# ZN 0.001673f
C12 VSS A2 0.036637f
C13 A3 a_244_68# 0.007f
C14 VNW A2 0.317841f
C15 a_1254_68# VSS 0.002331f
C16 VDD A2 0.041932f
C17 A1 VSS 0.037456f
C18 A3 A2 0.40854f
C19 ZN a_1458_68# 0.01082f
C20 ZN A2 0.068627f
C21 A1 VNW 0.345207f
C22 A1 VDD 0.044019f
C23 a_1254_68# A3 0.004873f
C24 A1 A3 0.831807f
C25 VNW VSS 0.006403f
C26 ZN a_1254_68# 0.008913f
C27 a_1060_68# VSS 0.001868f
C28 VDD VSS 0.004026f
C29 A1 ZN 0.071728f
C30 A3 VSS 0.248503f
C31 A4 A2 0.762551f
C32 a_438_68# VSS 0.00542f
C33 ZN VSS 0.89636f
C34 VDD VNW 0.1769f
C35 A3 VNW 0.300046f
C36 a_1060_68# A3 0.004303f
C37 VDD A3 0.040467f
C38 ZN VNW 0.062752f
C39 A1 A4 0.451294f
C40 a_1060_68# ZN 0.007219f
C41 A3 a_438_68# 0.007312f
C42 ZN VDD 1.39778f
C43 VSS VPW 0.597574f
C44 VDD VPW 0.397078f
C45 ZN VPW 0.12583f
C46 A1 VPW 0.558392f
C47 A2 VPW 0.513744f
C48 A3 VPW 0.547819f
C49 A4 VPW 0.580825f
C50 VNW VPW 3.05206f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
C0 ZN VNW 0.025997f
C1 VDD I 0.164681f
C2 VSS I 0.071429f
C3 VNW I 0.283715f
C4 ZN I 0.614595f
C5 VDD VSS 0.022662f
C6 VDD VNW 0.103267f
C7 VDD ZN 0.24022f
C8 VSS VNW 0.01054f
C9 ZN VSS 0.15979f
C10 VSS VPW 0.345063f
C11 ZN VPW 0.094435f
C12 VDD VPW 0.235951f
C13 I VPW 0.642286f
C14 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VNW VPW a_468_472#
+ a_224_472# a_244_68# a_916_472#
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
C0 a_224_472# A3 0.012212f
C1 a_224_472# VDD 0.016257f
C2 B2 VNW 0.125762f
C3 ZN a_916_472# 0.008827f
C4 A1 A2 0.038953f
C5 A1 ZN 0.164807f
C6 a_244_68# A2 0.356992f
C7 A2 VSS 0.030842f
C8 a_244_68# ZN 0.2576f
C9 ZN VSS 0.069913f
C10 A3 A2 0.129823f
C11 A2 VDD 0.071137f
C12 ZN VDD 0.006472f
C13 ZN B1 0.457921f
C14 a_244_68# a_916_472# 0.018012f
C15 VNW A2 0.121626f
C16 a_916_472# VDD 0.004169f
C17 a_468_472# A2 0.002382f
C18 VNW ZN 0.012941f
C19 a_244_68# A1 0.480797f
C20 A1 VSS 0.029231f
C21 A1 VDD 0.015114f
C22 B2 ZN 0.371232f
C23 a_244_68# VSS 0.329999f
C24 a_244_68# A3 0.010697f
C25 a_244_68# VDD 0.520053f
C26 A1 B1 0.13457f
C27 A3 VSS 0.046517f
C28 VSS VDD 0.027141f
C29 a_244_68# B1 0.212448f
C30 A3 VDD 0.236688f
C31 B1 VSS 0.072063f
C32 a_224_472# A2 0.014544f
C33 VNW A1 0.125824f
C34 B1 VDD 0.015317f
C35 A1 a_468_472# 0.001494f
C36 a_244_68# VNW 0.043485f
C37 VNW VSS 0.013582f
C38 a_244_68# a_468_472# 0.022611f
C39 VNW A3 0.13805f
C40 VNW VDD 0.158216f
C41 a_468_472# VDD 0.005594f
C42 a_244_68# B2 0.29062f
C43 VNW B1 0.116377f
C44 B2 VSS 0.072128f
C45 B2 VDD 0.018546f
C46 B2 B1 0.038725f
C47 a_244_68# a_224_472# 0.004752f
C48 a_224_472# VSS 0.00124f
C49 VSS VPW 0.474343f
C50 ZN VPW 0.00986f
C51 VDD VPW 0.363224f
C52 B2 VPW 0.282623f
C53 B1 VPW 0.257203f
C54 A1 VPW 0.255736f
C55 A2 VPW 0.254473f
C56 A3 VPW 0.308666f
C57 VNW VPW 2.35586f
C58 a_244_68# VPW 0.138666f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VNW VPW a_244_567# a_718_527#
+ a_2172_497# a_56_567# a_1948_68# a_728_93# a_1296_93#
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VPW nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
C0 VDD a_244_567# 0.006111f
C1 a_1296_93# ZN 0.029802f
C2 VDD a_728_93# 0.78216f
C3 a_56_567# A1 0.368741f
C4 ZN A3 0.033406f
C5 a_1296_93# a_1948_68# 0.005923f
C6 VNW ZN 0.032895f
C7 VSS ZN 0.004739f
C8 ZN a_2172_497# 0.03345f
C9 a_1948_68# A3 0.069927f
C10 VNW a_1948_68# 0.002346f
C11 VSS a_1948_68# 0.719859f
C12 VNW a_718_527# 0.020227f
C13 ZN a_728_93# 0.663929f
C14 VDD A1 0.022573f
C15 a_718_527# A2 0.141128f
C16 a_1948_68# a_728_93# 0.02618f
C17 a_56_567# VDD 0.056918f
C18 a_718_527# a_728_93# 0.21558f
C19 a_1296_93# A3 0.356198f
C20 a_1296_93# VNW 0.155715f
C21 a_1296_93# VSS 0.379749f
C22 a_718_527# A1 0.023145f
C23 VNW A3 0.298581f
C24 a_1296_93# A2 0.002759f
C25 VSS A3 0.047056f
C26 VSS VNW 0.009921f
C27 a_56_567# a_718_527# 0.00772f
C28 a_1504_93# a_1296_93# 0.003723f
C29 VNW A2 0.388997f
C30 VSS A2 0.051212f
C31 a_1296_93# a_728_93# 0.624643f
C32 VDD ZN 0.47211f
C33 a_1504_93# VSS 0.003902f
C34 a_244_567# A2 0.004089f
C35 a_728_93# A3 0.721889f
C36 VDD a_1948_68# 0.001604f
C37 VNW a_728_93# 0.385878f
C38 VSS a_728_93# 0.328386f
C39 a_728_93# a_2172_497# 0.010602f
C40 a_728_93# A2 0.516752f
C41 VDD a_718_527# 0.618394f
C42 VSS a_952_93# 0.003841f
C43 a_1948_68# ZN 0.381585f
C44 VNW A1 0.342048f
C45 VSS A1 0.0538f
C46 a_952_93# a_728_93# 0.003723f
C47 A1 A2 0.757944f
C48 a_56_567# VNW 0.187311f
C49 a_56_567# VSS 0.400197f
C50 a_56_567# A2 0.174541f
C51 a_56_567# a_244_567# 0.00105f
C52 a_728_93# A1 0.281966f
C53 a_1296_93# VDD 0.030892f
C54 a_56_567# a_728_93# 0.070648f
C55 VDD A3 0.022483f
C56 VNW VDD 0.370487f
C57 VSS VDD 0.011823f
C58 VDD a_2172_497# 0.010751f
C59 VDD A2 0.210416f
C60 VSS VPW 0.875791f
C61 ZN VPW 0.08517f
C62 A1 VPW 0.604039f
C63 A2 VPW 0.633287f
C64 VDD VPW 0.584594f
C65 A3 VPW 0.573218f
C66 VNW VPW 4.42794f
C67 a_1948_68# VPW 0.022025f
C68 a_718_527# VPW 0.001795f
C69 a_56_567# VPW 0.424713f
C70 a_728_93# VPW 0.65929f
C71 a_1296_93# VPW 0.317801f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VNW VPW a_36_68# a_244_497#
+ a_1657_68# a_1229_68# a_716_497#
X0 a_1229_68# B a_36_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
C0 VDD A2 0.147417f
C1 VSS a_1229_68# 0.002856f
C2 VSS A2 0.030494f
C3 A2 A1 0.722847f
C4 a_1229_68# a_36_68# 0.011792f
C5 a_36_68# A2 0.091399f
C6 VSS VDD 0.007619f
C7 a_244_497# A2 0.020646f
C8 VDD A1 0.033883f
C9 a_36_68# VDD 0.019083f
C10 a_716_497# ZN 0.025301f
C11 C VNW 0.309331f
C12 a_244_497# VDD 0.016799f
C13 VSS A1 0.031008f
C14 C ZN 0.501479f
C15 a_1657_68# B 0.002626f
C16 VSS a_36_68# 2.1107f
C17 ZN VNW 0.042076f
C18 C B 0.698524f
C19 a_36_68# A1 0.039393f
C20 B VNW 0.311256f
C21 B ZN 0.3603f
C22 a_716_497# A2 0.010693f
C23 A2 VNW 0.30827f
C24 a_716_497# VDD 0.008883f
C25 ZN A2 1.02528f
C26 a_1229_68# B 0.003462f
C27 B A2 0.037237f
C28 C VDD 0.056662f
C29 VDD VNW 0.219901f
C30 a_1657_68# VSS 0.002208f
C31 ZN VDD 0.761655f
C32 C VSS 0.04168f
C33 B VDD 0.089771f
C34 a_1657_68# a_36_68# 0.009002f
C35 VSS VNW 0.005994f
C36 VSS ZN 0.004788f
C37 C a_36_68# 0.055076f
C38 A1 VNW 0.269127f
C39 VSS B 0.032629f
C40 a_36_68# VNW 0.00468f
C41 ZN A1 0.622246f
C42 ZN a_36_68# 0.528658f
C43 B a_36_68# 0.587375f
C44 a_244_497# ZN 0.006285f
C45 VSS VPW 0.620026f
C46 ZN VPW 0.062404f
C47 VDD VPW 0.531064f
C48 C VPW 0.529789f
C49 B VPW 0.589191f
C50 A1 VPW 0.58772f
C51 A2 VPW 0.613706f
C52 VNW VPW 3.34705f
C53 a_36_68# VPW 0.052951f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW a_428_148# a_36_148#
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
C0 A3 A2 0.340591f
C1 VNW VSS 0.007319f
C2 A3 Z 0.001054f
C3 VDD VSS 0.012823f
C4 a_428_148# A3 0.001335f
C5 VNW A2 0.189332f
C6 A3 VNW 0.213241f
C7 VDD A2 0.022493f
C8 VNW Z 0.033257f
C9 A1 a_36_148# 0.205722f
C10 A3 VDD 0.022574f
C11 VDD Z 0.164783f
C12 VNW VDD 0.134134f
C13 A1 VSS 0.00434f
C14 a_36_148# VSS 0.798993f
C15 A1 A2 0.307806f
C16 a_36_148# A2 0.141951f
C17 A3 a_36_148# 0.477475f
C18 a_36_148# Z 0.156534f
C19 a_428_148# a_36_148# 0.007047f
C20 A1 VNW 0.214361f
C21 A1 a_244_148# 0.002081f
C22 VNW a_36_148# 0.194548f
C23 A2 VSS 0.004456f
C24 A1 VDD 0.021719f
C25 a_244_148# a_36_148# 0.004781f
C26 A3 VSS 0.005273f
C27 a_36_148# VDD 0.556761f
C28 Z VSS 0.093779f
C29 VSS VPW 0.415001f
C30 Z VPW 0.095371f
C31 VDD VPW 0.277732f
C32 A3 VPW 0.275015f
C33 A2 VPW 0.257076f
C34 A1 VPW 0.330738f
C35 VNW VPW 2.00777f
C36 a_36_148# VPW 0.388358f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW a_1044_68# a_452_68#
+ a_276_68# a_860_68#
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 ZN A1 0.430404f
C1 VDD VNW 0.172362f
C2 VDD A1 0.041745f
C3 a_276_68# VSS 0.003438f
C4 ZN a_276_68# 0.007178f
C5 A2 VSS 0.130985f
C6 ZN A2 0.082264f
C7 A1 a_452_68# 0.001247f
C8 A2 a_860_68# 0.003842f
C9 VDD A2 0.041181f
C10 A1 VNW 0.280755f
C11 A3 VSS 0.074424f
C12 ZN A3 1.24554f
C13 A2 VNW 0.279783f
C14 A2 A1 0.708241f
C15 VDD A3 0.099291f
C16 a_1044_68# VSS 0.00861f
C17 a_1044_68# ZN 0.001223f
C18 VNW A3 0.347673f
C19 ZN VSS 0.476547f
C20 A1 A3 0.037905f
C21 a_860_68# VSS 0.005864f
C22 ZN a_860_68# 0.001808f
C23 VDD VSS 0.009236f
C24 ZN VDD 0.550625f
C25 A2 A3 1.13496f
C26 a_452_68# VSS 0.003244f
C27 ZN a_452_68# 0.007752f
C28 a_1044_68# A2 0.006328f
C29 VNW VSS 0.007349f
C30 ZN VNW 0.034063f
C31 A1 VSS 0.050488f
C32 VSS VPW 0.511432f
C33 ZN VPW 0.112753f
C34 VDD VPW 0.407724f
C35 A1 VPW 0.540441f
C36 A2 VPW 0.524145f
C37 A3 VPW 0.582222f
C38 VNW VPW 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW a_692_473#
+ a_254_473# a_66_473# a_2700_473# a_1660_473# a_3220_473# a_1212_473# a_2180_473#
+ a_3740_473# a_1920_473#
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VPW nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
C0 a_692_473# a_66_473# 0.022803f
C1 A2 VDD 0.054912f
C2 a_66_473# VDD 3.19476f
C3 a_1920_473# a_66_473# 0.023791f
C4 A2 VNW 0.584134f
C5 a_66_473# VNW 0.040351f
C6 a_254_473# a_66_473# 0.016207f
C7 a_66_473# A4 0.100571f
C8 a_2180_473# ZN 0.018904f
C9 VDD ZN 0.007051f
C10 a_1920_473# ZN 0.017667f
C11 ZN VNW 0.038639f
C12 a_1660_473# VDD 0.008572f
C13 ZN A4 1.44735f
C14 a_66_473# a_3220_473# 0.021354f
C15 a_66_473# A2 0.182327f
C16 A3 VSS 0.078892f
C17 VSS A1 0.093176f
C18 a_3740_473# VDD 0.003118f
C19 a_3220_473# ZN 0.019778f
C20 a_2700_473# VDD 0.003457f
C21 A2 ZN 2.14591f
C22 a_66_473# ZN 0.956309f
C23 a_1660_473# a_66_473# 0.035002f
C24 A3 VDD 0.086829f
C25 VSS VDD 0.009708f
C26 VDD A1 0.055928f
C27 A3 VNW 0.567739f
C28 VSS VNW 0.006947f
C29 A1 VNW 0.553741f
C30 A3 A4 1.96796f
C31 VSS A4 0.099821f
C32 a_1660_473# ZN 0.00216f
C33 a_3740_473# A2 0.010293f
C34 a_3740_473# a_66_473# 0.028219f
C35 a_66_473# a_2700_473# 0.021497f
C36 a_2180_473# VDD 0.00368f
C37 VDD a_1212_473# 0.014305f
C38 a_692_473# VDD 0.017923f
C39 a_3740_473# ZN 0.004594f
C40 a_2700_473# ZN 0.019492f
C41 a_1920_473# VDD 0.004058f
C42 VDD VNW 0.394018f
C43 a_254_473# VDD 0.012952f
C44 VDD A4 0.110338f
C45 A3 A2 0.0303f
C46 A2 VSS 0.076134f
C47 A3 a_66_473# 1.66251f
C48 A2 A1 2.13585f
C49 a_66_473# VSS 0.01197f
C50 a_66_473# A1 0.077909f
C51 A4 VNW 0.513548f
C52 A3 ZN 0.417545f
C53 VSS ZN 4.39577f
C54 ZN A1 1.60655f
C55 a_3220_473# VDD 0.003326f
C56 a_66_473# a_2180_473# 0.020817f
C57 A3 a_1660_473# 0.0054f
C58 a_66_473# a_1212_473# 0.018664f
C59 VSS VPW 1.3434f
C60 ZN VPW 0.240026f
C61 VDD VPW 0.844436f
C62 A1 VPW 1.40024f
C63 A2 VPW 1.30271f
C64 A4 VPW 1.33565f
C65 A3 VPW 1.29175f
C66 VNW VPW 6.70706f
C67 a_66_473# VPW 0.11665f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VNW VPW a_49_472# a_1133_69#
+ a_741_69#
X0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VPW nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VPW nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
C0 ZN A1 0.182845f
C1 VDD VNW 0.151549f
C2 a_741_69# VSS 0.002035f
C3 A2 VDD 0.029358f
C4 ZN a_1133_69# 0.001193f
C5 VNW VSS 0.0086f
C6 ZN VDD 0.008463f
C7 a_1133_69# A1 0.003427f
C8 A2 VSS 0.047574f
C9 VDD A1 0.028601f
C10 a_49_472# VNW 0.012852f
C11 ZN VSS 0.784804f
C12 A2 a_49_472# 0.086717f
C13 A1 VSS 0.129775f
C14 VNW B 0.260678f
C15 ZN a_49_472# 0.475008f
C16 A2 B 0.029994f
C17 a_49_472# A1 0.03417f
C18 a_1133_69# VSS 0.00441f
C19 ZN B 0.20884f
C20 VDD VSS 0.009099f
C21 a_49_472# VDD 1.09818f
C22 a_49_472# VSS 0.01207f
C23 VDD B 0.045174f
C24 A2 a_741_69# 0.001142f
C25 ZN a_741_69# 0.006341f
C26 A2 VNW 0.272677f
C27 VSS B 0.061328f
C28 ZN VNW 0.025755f
C29 a_49_472# B 0.234399f
C30 A1 VNW 0.241301f
C31 ZN A2 0.800412f
C32 A2 A1 0.809974f
C33 VSS VPW 0.510011f
C34 ZN VPW 0.070911f
C35 VDD VPW 0.327438f
C36 A1 VPW 0.556927f
C37 A2 VPW 0.56333f
C38 B VPW 0.662515f
C39 VNW VPW 2.52991f
C40 a_49_472# VPW 0.098072f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2$1 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VNW I 0.285482f
C1 VNW ZN 0.027829f
C2 VNW VDD 0.097124f
C3 VNW VSS 0.010163f
C4 ZN I 0.58604f
C5 VDD I 0.074838f
C6 VSS I 0.091531f
C7 ZN VDD 0.266247f
C8 ZN VSS 0.179304f
C9 VDD VSS 0.023187f
C10 VSS VPW 0.308828f
C11 ZN VPW 0.100523f
C12 VDD VPW 0.240805f
C13 I VPW 0.610668f
C14 VNW VPW 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VNW VPW a_448_472#
+ a_36_151# a_1293_527# a_3081_151# a_1284_156# a_1040_527# a_1353_112# a_836_156#
+ a_1697_156# a_2449_156# a_3129_107# a_2225_156#
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VPW nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VPW nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VPW nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VPW nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VPW nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VPW nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VPW nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
C0 a_36_151# a_2225_156# 0.153684f
C1 a_448_472# a_2449_156# 0.056679f
C2 VDD a_1353_112# 0.016257f
C3 a_836_156# VNW 0.01368f
C4 a_1040_527# VNW 0.223863f
C5 VSS D 0.067877f
C6 a_2225_156# a_1353_112# 0.152869f
C7 CLK a_448_472# 0.001313f
C8 VNW SETN 0.811046f
C9 SETN a_3129_107# 0.089288f
C10 VDD a_1040_527# 0.039677f
C11 a_448_472# a_36_151# 0.473132f
C12 VNW VSS 0.009462f
C13 VDD SETN 0.127822f
C14 a_36_151# a_2449_156# 0.005967f
C15 VSS a_3129_107# 0.136769f
C16 SETN a_2225_156# 0.070597f
C17 VDD VSS 0.013814f
C18 VNW D 0.1615f
C19 a_448_472# a_1353_112# 0.317251f
C20 a_448_472# a_1697_156# 0.007618f
C21 VSS a_2225_156# 1.18908f
C22 CLK a_36_151# 0.700974f
C23 VDD D 0.004944f
C24 a_448_472# a_836_156# 0.427756f
C25 VSS a_1284_156# 0.003637f
C26 VNW a_3129_107# 0.323464f
C27 a_448_472# a_1040_527# 0.869605f
C28 a_448_472# SETN 0.083903f
C29 VDD VNW 0.539099f
C30 VDD a_3129_107# 0.351307f
C31 SETN a_2449_156# 0.302222f
C32 a_36_151# a_1353_112# 0.840879f
C33 a_448_472# VSS 1.07431f
C34 VNW a_2225_156# 0.209033f
C35 a_2225_156# a_3129_107# 0.514036f
C36 a_448_472# D 0.400104f
C37 a_836_156# a_36_151# 0.015697f
C38 VDD a_2225_156# 0.073415f
C39 a_3081_151# a_2225_156# 0.004129f
C40 a_1040_527# a_36_151# 0.206392f
C41 a_36_151# a_1293_527# 0.008379f
C42 a_1697_156# a_1353_112# 0.002752f
C43 SETN a_36_151# 0.077775f
C44 CLK VSS 0.021941f
C45 a_448_472# VNW 0.400964f
C46 Q VSS 0.131272f
C47 VSS a_36_151# 0.286331f
C48 a_1040_527# a_1353_112# 0.387423f
C49 VNW a_2449_156# 0.043816f
C50 a_2449_156# a_3129_107# 0.00955f
C51 a_448_472# VDD 0.624585f
C52 SETN a_1353_112# 0.072983f
C53 a_36_151# D 0.092705f
C54 VDD a_2449_156# 0.208631f
C55 a_3081_151# a_2449_156# 0.001203f
C56 a_836_156# a_1040_527# 0.068207f
C57 a_448_472# a_2225_156# 0.153996f
C58 VSS a_1353_112# 0.027348f
C59 CLK VNW 0.136589f
C60 a_2225_156# a_2449_156# 0.569174f
C61 Q VNW 0.031621f
C62 a_1040_527# a_1293_527# 0.00215f
C63 a_448_472# a_1284_156# 0.002691f
C64 Q a_3129_107# 0.179468f
C65 a_1040_527# SETN 0.063241f
C66 VNW a_36_151# 0.909435f
C67 a_836_156# VSS 0.050008f
C68 CLK VDD 0.022091f
C69 Q VDD 0.282179f
C70 a_1040_527# VSS 0.060221f
C71 VDD a_36_151# 1.41468f
C72 VSS SETN 0.008083f
C73 a_836_156# D 0.108102f
C74 VNW a_1353_112# 0.219511f
C75 Q VPW 0.105566f
C76 VSS VPW 1.35707f
C77 SETN VPW 0.710246f
C78 D VPW 0.247102f
C79 VDD VPW 0.833181f
C80 CLK VPW 0.290467f
C81 VNW VPW 6.44257f
C82 a_2449_156# VPW 0.049992f
C83 a_2225_156# VPW 0.434082f
C84 a_3129_107# VPW 0.58406f
C85 a_836_156# VPW 0.019766f
C86 a_1040_527# VPW 0.302082f
C87 a_1353_112# VPW 0.286513f
C88 a_448_472# VPW 1.21246f
C89 a_36_151# VPW 1.31409f
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[8] ctlp[0]
+ ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8] ctlp[9] cal clk
+ clkc comp en result[0] result[1] result[2] result[3] result[4] result[5] result[6]
+ result[7] result[8] result[9] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4]
+ trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] valid output13/a_224_472# output23/a_224_472#
+ net27 output25/a_224_472# cal_itt\[1\] ctln[7] net15 net59 ctln[9] output10/a_224_472#
+ net24 output11/a_224_472# output21/a_224_472# net14 output12/a_224_472# output22/a_224_472#
+ vdd net62 net20 vss
XFILLER_0_17_200 vdd vss vdd vss FILLER_0_17_200/a_36_472# FILLER_0_17_200/a_572_375#
+ FILLER_0_17_200/a_124_375# FILLER_0_17_200/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_294_ vdd vss _008_ _104_ _106_ vdd vss _294_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_432_ _021_ mask\[3\] net63 vss net80 vdd vdd vss _432_/a_2665_112# _432_/a_448_472#
+ _432_/a_796_472# _432_/a_36_151# _432_/a_1204_472# _432_/a_3041_156# _432_/a_1000_472#
+ _432_/a_1308_423# _432_/a_1456_156# _432_/a_1288_156# _432_/a_2248_156# _432_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ vdd vss _363_/a_36_68# _363_/a_244_472#
+ _363_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ vdd vss _346_/a_49_472# _346_/a_665_69#
+ _346_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd vdd vss _415_/a_2665_112# _415_/a_448_472#
+ _415_/a_796_472# _415_/a_36_151# _415_/a_1204_472# _415_/a_3041_156# _415_/a_1000_472#
+ _415_/a_1308_423# _415_/a_1456_156# _415_/a_1288_156# _415_/a_2248_156# _415_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd vdd vss _277_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss vdd vss FILLER_0_19_125/a_36_472# FILLER_0_19_125/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss vdd vss FILLER_0_15_150/a_36_472# FILLER_0_15_150/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss vdd vss FILLER_0_21_142/a_36_472# FILLER_0_21_142/a_572_375#
+ FILLER_0_21_142/a_124_375# FILLER_0_21_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss vdd vss FILLER_0_16_73/a_36_472# FILLER_0_16_73/a_572_375#
+ FILLER_0_16_73/a_124_375# FILLER_0_16_73/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss vdd vss output20/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss vdd vss output31/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss vdd vss output42/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 ctln[0] net7 vdd vss vdd vss output7/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss vdd vss FILLER_0_5_117/a_36_472# FILLER_0_5_117/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss vdd vss FILLER_0_5_128/a_36_472# FILLER_0_5_128/a_572_375#
+ FILLER_0_5_128/a_124_375# FILLER_0_5_128/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_293_ net31 vdd vss _106_ mask\[4\] _105_ vdd vss _293_/a_36_472# _293_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_431_ _020_ mask\[2\] net53 vss net70 vdd vdd vss _431_/a_2665_112# _431_/a_448_472#
+ _431_/a_796_472# _431_/a_36_151# _431_/a_1204_472# _431_/a_3041_156# _431_/a_1000_472#
+ _431_/a_1308_423# _431_/a_1456_156# _431_/a_1288_156# _431_/a_2248_156# _431_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_362_ vdd vss trim_mask\[1\] _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_345_ vss _144_ _132_ vdd vdd vss _345_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ vss _093_ _092_ vdd vdd vss _276_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd vdd vss _414_/a_2665_112# _414_/a_448_472#
+ _414_/a_796_472# _414_/a_36_151# _414_/a_1204_472# _414_/a_3041_156# _414_/a_1000_472#
+ _414_/a_1308_423# _414_/a_1456_156# _414_/a_1288_156# _414_/a_2248_156# _414_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd vdd vss _328_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss vdd vss FILLER_0_9_28/a_1916_375# FILLER_0_9_28/a_1380_472#
+ FILLER_0_9_28/a_3260_375# FILLER_0_9_28/a_36_472# FILLER_0_9_28/a_932_472# FILLER_0_9_28/a_2812_375#
+ FILLER_0_9_28/a_2276_472# FILLER_0_9_28/a_1828_472# FILLER_0_9_28/a_3172_472# FILLER_0_9_28/a_572_375#
+ FILLER_0_9_28/a_2724_472# FILLER_0_9_28/a_124_375# FILLER_0_9_28/a_1468_375# FILLER_0_9_28/a_1020_375#
+ FILLER_0_9_28/a_484_472# FILLER_0_9_28/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_204 vdd vss vdd vss FILLER_0_3_204/a_36_472# FILLER_0_3_204/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _078_ vdd vss _080_ _073_ _076_ vdd vss _259_/a_455_68# _259_/a_271_68# gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd vss vdd vss FILLER_0_16_107/a_36_472# FILLER_0_16_107/a_572_375#
+ FILLER_0_16_107/a_124_375# FILLER_0_16_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss vdd vss output21/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss vdd vss output43/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss vdd vss output32/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss vdd vss output10/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss vdd vss output8/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ vss _105_ _098_ vdd vdd vss _292_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_430_ _019_ mask\[1\] net63 vss net80 vdd vdd vss _430_/a_2665_112# _430_/a_448_472#
+ _430_/a_796_472# _430_/a_36_151# _430_/a_1204_472# _430_/a_3041_156# _430_/a_1000_472#
+ _430_/a_1308_423# _430_/a_1456_156# _430_/a_1288_156# _430_/a_2248_156# _430_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_361_ vdd vss _154_ _086_ _119_ vdd vss _361_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss vdd vss FILLER_0_7_72/a_1916_375# FILLER_0_7_72/a_1380_472#
+ FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472# FILLER_0_7_72/a_932_472# FILLER_0_7_72/a_2812_375#
+ FILLER_0_7_72/a_2276_472# FILLER_0_7_72/a_1828_472# FILLER_0_7_72/a_3172_472# FILLER_0_7_72/a_572_375#
+ FILLER_0_7_72/a_2724_472# FILLER_0_7_72/a_124_375# FILLER_0_7_72/a_1468_375# FILLER_0_7_72/a_1020_375#
+ FILLER_0_7_72/a_484_472# FILLER_0_7_72/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ vdd vss _275_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__191__I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd vdd vss _413_/a_2665_112# _413_/a_448_472#
+ _413_/a_796_472# _413_/a_36_151# _413_/a_1204_472# _413_/a_3041_156# _413_/a_1000_472#
+ _413_/a_1308_423# _413_/a_1456_156# _413_/a_1288_156# _413_/a_2248_156# _413_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_96 vdd vss vdd vss FILLER_0_24_96/a_36_472# FILLER_0_24_96/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss vdd vss FILLER_0_24_63/a_36_472# FILLER_0_24_63/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ vdd vss _043_ net27 mask\[0\] vdd vss _189_/a_255_603# _189_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_327_ _131_ vdd vss _016_ _127_ _130_ vdd vss _327_/a_36_472# _327_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ vss _079_ _078_ vdd vdd vss _258_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss vdd vss FILLER_0_18_171/a_36_472# FILLER_0_18_171/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss vdd vss FILLER_0_24_130/a_36_472# FILLER_0_24_130/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss vdd vss FILLER_0_21_133/a_36_472# FILLER_0_21_133/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss vdd vss FILLER_0_8_138/a_36_472# FILLER_0_8_138/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss vdd vss FILLER_0_8_127/a_36_472# FILLER_0_8_127/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 ctlp[5] net22 vdd vss vdd vss output22/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 result[6] net33 vdd vss vdd vss output33/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss vdd vss output44/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss vdd vss output11/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss vdd vss output9/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd vdd vss _291_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss vdd vss FILLER_0_4_152/a_36_472# FILLER_0_4_152/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss vdd vss FILLER_0_4_185/a_36_472# FILLER_0_4_185/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd vdd vss _360_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss vdd vss FILLER_0_13_65/a_36_472# FILLER_0_13_65/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ vdd vss _343_/a_49_472# _343_/a_665_69#
+ _343_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ vdd vss _274_/a_36_68# _274_/a_1612_497#
+ _274_/a_2124_68# _274_/a_244_497# _274_/a_2960_68# _274_/a_3368_68# _274_/a_2552_68#
+ _274_/a_1164_497# _274_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd vdd vss _412_/a_2665_112# _412_/a_448_472#
+ _412_/a_796_472# _412_/a_36_151# _412_/a_1204_472# _412_/a_3041_156# _412_/a_1000_472#
+ _412_/a_1308_423# _412_/a_1456_156# _412_/a_1288_156# _412_/a_2248_156# _412_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__292__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ vdd vss _326_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ vdd vss _257_/a_36_472# _257_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__301__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss vdd vss FILLER_0_15_142/a_36_472# FILLER_0_15_142/a_572_375#
+ FILLER_0_15_142/a_124_375# FILLER_0_15_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 ctlp[6] net23 vdd vss vdd vss output23/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss vdd vss output45/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss vdd vss output34/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss vdd vss output12/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss vdd vss FILLER_0_5_109/a_36_472# FILLER_0_5_109/a_572_375#
+ FILLER_0_5_109/a_124_375# FILLER_0_5_109/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss vdd vss FILLER_0_17_226/a_36_472# FILLER_0_17_226/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss vdd vss FILLER_0_4_197/a_1380_472# FILLER_0_4_197/a_36_472#
+ FILLER_0_4_197/a_932_472# FILLER_0_4_197/a_572_375# FILLER_0_4_197/a_124_375# FILLER_0_4_197/a_1468_375#
+ FILLER_0_4_197/a_1020_375# FILLER_0_4_197/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ vdd vss _290_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss vdd vss FILLER_0_9_223/a_36_472# FILLER_0_9_223/a_572_375#
+ FILLER_0_9_223/a_124_375# FILLER_0_9_223/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_273_ vss _090_ state\[0\] vdd vdd vss _273_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd vdd vss _411_/a_2665_112# _411_/a_448_472#
+ _411_/a_796_472# _411_/a_36_151# _411_/a_1204_472# _411_/a_3041_156# _411_/a_1000_472#
+ _411_/a_1308_423# _411_/a_1456_156# _411_/a_1288_156# _411_/a_2248_156# _411_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout80 vss net80 net81 vdd vdd vss fanout80/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_325_ vdd vss _130_ _118_ _129_ vdd vss _325_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd vss vdd vss FILLER_0_10_78/a_1380_472# FILLER_0_10_78/a_36_472#
+ FILLER_0_10_78/a_932_472# FILLER_0_10_78/a_572_375# FILLER_0_10_78/a_124_375# FILLER_0_10_78/a_1468_375#
+ FILLER_0_10_78/a_1020_375# FILLER_0_10_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ vdd vss _256_/a_36_68# _256_/a_1612_497#
+ _256_/a_2124_68# _256_/a_244_497# _256_/a_2960_68# _256_/a_3368_68# _256_/a_2552_68#
+ _256_/a_1164_497# _256_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ vdd vss _308_/a_848_380# _308_/a_1084_68#
+ _308_/a_124_24# _308_/a_1152_472# _308_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss vdd vss FILLER_0_1_98/a_36_472# FILLER_0_1_98/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ vdd vss _239_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss vdd vss FILLER_0_12_124/a_36_472# FILLER_0_12_124/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss vdd vss FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 ctlp[7] net24 vdd vss vdd vss output24/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss vdd vss output35/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss vdd vss output46/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss vdd vss FILLER_0_18_2/a_1916_375# FILLER_0_18_2/a_1380_472#
+ FILLER_0_18_2/a_3260_375# FILLER_0_18_2/a_36_472# FILLER_0_18_2/a_932_472# FILLER_0_18_2/a_2812_375#
+ FILLER_0_18_2/a_2276_472# FILLER_0_18_2/a_1828_472# FILLER_0_18_2/a_3172_472# FILLER_0_18_2/a_572_375#
+ FILLER_0_18_2/a_2724_472# FILLER_0_18_2/a_124_375# FILLER_0_18_2/a_1468_375# FILLER_0_18_2/a_1020_375#
+ FILLER_0_18_2/a_484_472# FILLER_0_18_2/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 ctln[6] net13 vdd vss vdd vss output13/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss vdd vss FILLER_0_7_162/a_36_472# FILLER_0_7_162/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss vdd vss FILLER_0_7_195/a_36_472# FILLER_0_7_195/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ vdd vss _341_/a_49_472# _341_/a_665_69#
+ _341_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss vdd vss _410_/a_36_68# _410_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ vdd vss _272_/a_36_472# _272_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd vdd vss fanout70/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ _076_ vss vdd _057_ vdd vss _255_/a_224_552# gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_324_ vdd vss _129_ calibrate _062_ vdd vss _324_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output40_I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 vss net81 net82 vdd vdd vss fanout81/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_55 vdd vss vdd vss FILLER_0_19_55/a_36_472# FILLER_0_19_55/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_307_ vdd vss _114_ _113_ _096_ vdd vss _307_/a_234_472# _307_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] vdd vss _238_/a_255_603# _238_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss vdd vss FILLER_0_21_125/a_36_472# FILLER_0_21_125/a_572_375#
+ FILLER_0_21_125/a_124_375# FILLER_0_21_125/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss vdd vss FILLER_0_16_89/a_1380_472# FILLER_0_16_89/a_36_472#
+ FILLER_0_16_89/a_932_472# FILLER_0_16_89/a_572_375# FILLER_0_16_89/a_124_375# FILLER_0_16_89/a_1468_375#
+ FILLER_0_16_89/a_1020_375# FILLER_0_16_89/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss vdd vss FILLER_0_12_136/a_1380_472# FILLER_0_12_136/a_36_472#
+ FILLER_0_12_136/a_932_472# FILLER_0_12_136/a_572_375# FILLER_0_12_136/a_124_375#
+ FILLER_0_12_136/a_1468_375# FILLER_0_12_136/a_1020_375# FILLER_0_12_136/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 ctlp[8] net25 vdd vss vdd vss output25/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss vdd vss output47/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 result[9] net36 vdd vss vdd vss output36/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss vdd vss output14/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss vdd vss FILLER_0_4_144/a_36_472# FILLER_0_4_144/a_572_375#
+ FILLER_0_4_144/a_124_375# FILLER_0_4_144/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss vdd vss FILLER_0_4_177/a_36_472# FILLER_0_4_177/a_572_375#
+ FILLER_0_4_177/a_124_375# FILLER_0_4_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd vdd vss _340_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss vdd vss FILLER_0_10_256/a_36_472# FILLER_0_10_256/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__200__I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_99 vdd vss vdd vss FILLER_0_4_99/a_36_472# FILLER_0_4_99/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss vdd vss FILLER_0_6_239/a_36_472# FILLER_0_6_239/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout71 vss net71 net73 vdd vdd vss fanout71/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 net60 vss vdd net61 vdd vss fanout60/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_323_ vss _015_ _128_ vdd vdd vss _323_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd vdd vss fanout82/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ vdd vss _254_/a_448_472# _254_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_237_ vdd vss net40 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_306_ vss _113_ _057_ vdd vdd vss _306_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_57 vdd vss vdd vss FILLER_0_16_57/a_1380_472# FILLER_0_16_57/a_36_472#
+ FILLER_0_16_57/a_932_472# FILLER_0_16_57/a_572_375# FILLER_0_16_57/a_124_375# FILLER_0_16_57/a_1468_375#
+ FILLER_0_16_57/a_1020_375# FILLER_0_16_57/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss vdd vss output26/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss vdd vss output15/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss vdd vss output48/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss vdd vss output37/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss vdd vss FILLER_0_17_218/a_36_472# FILLER_0_17_218/a_572_375#
+ FILLER_0_17_218/a_124_375# FILLER_0_17_218/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss vdd vss FILLER_0_4_123/a_36_472# FILLER_0_4_123/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ vdd vss _270_/a_36_472# _270_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ vdd vss _399_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ vdd vss _322_/a_848_380# _322_/a_1084_68# _322_/a_124_24#
+ _322_/a_1152_472# _322_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd vdd vss fanout61/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd vdd vss fanout72/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd vss vdd vss FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net50 vss vdd net52 vdd vss fanout50/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] vdd vss _253_/a_36_68#
+ _253_/a_1732_68# _253_/a_244_68# _253_/a_1100_68# _253_/a_1528_68# _253_/a_672_68#
+ gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_305_ vdd vss _112_ net1 _081_ vdd vss _305_/a_36_159# gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ net40 vss vdd _064_ vdd vss _236_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss vdd vss FILLER_0_20_193/a_36_472# FILLER_0_20_193/a_572_375#
+ FILLER_0_20_193/a_124_375# FILLER_0_20_193/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd vdd vss _219_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss vdd vss output27/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss vdd vss output16/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss vdd vss output38/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss vdd vss FILLER_0_16_241/a_36_472# FILLER_0_16_241/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd vdd vss _398_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vss vdd vss FILLER_0_10_247/a_36_472# FILLER_0_10_247/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_214 vdd vss vdd vss FILLER_0_10_214/a_36_472# FILLER_0_10_214/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_91 vdd vss vdd vss FILLER_0_14_91/a_36_472# FILLER_0_14_91/a_572_375#
+ FILLER_0_14_91/a_124_375# FILLER_0_14_91/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__209__I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I vss net19 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss vdd vss FILLER_0_19_47/a_36_472# FILLER_0_19_47/a_572_375#
+ FILLER_0_19_47/a_124_375# FILLER_0_19_47/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd vdd vss fanout73/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 net62 vss vdd net64 vdd vss fanout62/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vss net51 net52 vdd vdd vss fanout51/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ vdd vss _321_/a_2590_472# _321_/a_170_472#
+ _321_/a_1602_69# _321_/a_786_69# _321_/a_3126_472# _321_/a_1194_69# _321_/a_3662_472#
+ _321_/a_2034_472# _321_/a_358_69# gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_252_ vdd vss cal_itt\[0\] _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_100 vdd vss vdd vss FILLER_0_18_100/a_36_472# FILLER_0_18_100/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss vdd vss FILLER_0_18_177/a_1916_375# FILLER_0_18_177/a_1380_472#
+ FILLER_0_18_177/a_3260_375# FILLER_0_18_177/a_36_472# FILLER_0_18_177/a_932_472#
+ FILLER_0_18_177/a_2812_375# FILLER_0_18_177/a_2276_472# FILLER_0_18_177/a_1828_472#
+ FILLER_0_18_177/a_3172_472# FILLER_0_18_177/a_572_375# FILLER_0_18_177/a_2724_472#
+ FILLER_0_18_177/a_124_375# FILLER_0_18_177/a_1468_375# FILLER_0_18_177/a_1020_375#
+ FILLER_0_18_177/a_484_472# FILLER_0_18_177/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ vdd vss _304_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] vdd vss _235_/a_255_603# _235_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss vdd vss FILLER_0_16_37/a_36_472# FILLER_0_16_37/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss vdd vss output17/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss vdd vss output28/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss vdd vss output39/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss vdd vss FILLER_0_13_212/a_1380_472# FILLER_0_13_212/a_36_472#
+ FILLER_0_13_212/a_932_472# FILLER_0_13_212/a_572_375# FILLER_0_13_212/a_124_375#
+ FILLER_0_13_212/a_1468_375# FILLER_0_13_212/a_1020_375# FILLER_0_13_212/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ vdd vss _397_/a_36_472# _397_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss vdd vss FILLER_0_14_81/a_36_472# FILLER_0_14_81/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout63 net63 vss vdd net64 vdd vss fanout63/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ vdd vss _320_/a_1792_472# _320_/a_224_472#
+ _320_/a_1568_472# _320_/a_36_472# _320_/a_1120_472# _320_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_28 vdd vss vdd vss FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 vss net74 net82 vdd vdd vss fanout74/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net52 vss vdd net57 vdd vss fanout52/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ vdd vss _251_/a_468_472# _251_/a_244_472# _251_/a_1130_472#
+ _251_/a_906_472# gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_449_ _038_ en_co_clk net55 vss net72 vdd vdd vss _449_/a_2665_112# _449_/a_448_472#
+ _449_/a_796_472# _449_/a_36_151# _449_/a_1204_472# _449_/a_3041_156# _449_/a_1000_472#
+ _449_/a_1308_423# _449_/a_1456_156# _449_/a_1288_156# _449_/a_2248_156# _449_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ vdd vss _303_/a_36_472# _303_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_217_ vss net26 _052_ vdd vdd vss _217_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_181 vdd vss vdd vss FILLER_0_14_181/a_36_472# FILLER_0_14_181/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 ctlp[1] net18 vdd vss vdd vss output18/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss vdd vss output29/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ vdd vss _396_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout53 net53 vss vdd net56 vdd vss fanout53/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_250_ vss _072_ _071_ vdd vdd vss _250_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 vss net75 net76 vdd vdd vss fanout75/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd vdd vss fanout64/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd vdd vss _448_/a_2665_112# _448_/a_448_472#
+ _448_/a_796_472# _448_/a_36_151# _448_/a_1204_472# _448_/a_3041_156# _448_/a_1000_472#
+ _448_/a_1308_423# _448_/a_1456_156# _448_/a_1288_156# _448_/a_2248_156# _448_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ vdd vss _379_/a_36_472# _379_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_302_ vdd vss _012_ _093_ _110_ vdd vss _302_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss vdd vss FILLER_0_21_28/a_1916_375# FILLER_0_21_28/a_1380_472#
+ FILLER_0_21_28/a_3260_375# FILLER_0_21_28/a_36_472# FILLER_0_21_28/a_932_472# FILLER_0_21_28/a_2812_375#
+ FILLER_0_21_28/a_2276_472# FILLER_0_21_28/a_1828_472# FILLER_0_21_28/a_3172_472#
+ FILLER_0_21_28/a_572_375# FILLER_0_21_28/a_2724_472# FILLER_0_21_28/a_124_375# FILLER_0_21_28/a_1468_375#
+ FILLER_0_21_28/a_1020_375# FILLER_0_21_28/a_484_472# FILLER_0_21_28/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__216__A2 vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ vss net39 _063_ vdd vdd vss _233_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss vdd vss FILLER_0_15_116/a_36_472# FILLER_0_15_116/a_572_375#
+ FILLER_0_15_116/a_124_375# FILLER_0_15_116/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_216_ vdd vss _052_ mask\[9\] net36 vdd vss _216_/a_255_603# _216_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_146 vdd vss vdd vss FILLER_0_7_146/a_36_472# FILLER_0_7_146/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 ctlp[2] net19 vdd vss vdd vss output19/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss vdd vss FILLER_0_7_59/a_36_472# FILLER_0_7_59/a_572_375# FILLER_0_7_59/a_124_375#
+ FILLER_0_7_59/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss vdd vss FILLER_0_16_255/a_36_472# FILLER_0_16_255/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss vdd vss FILLER_0_0_130/a_36_472# FILLER_0_0_130/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss vdd vss FILLER_0_8_263/a_36_472# FILLER_0_8_263/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss vdd vss FILLER_0_14_50/a_36_472# FILLER_0_14_50/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ vdd vss _395_/a_1492_488# _395_/a_244_68#
+ _395_/a_1044_488# _395_/a_636_68# _395_/a_36_488# gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss vdd vss FILLER_0_4_49/a_36_472# FILLER_0_4_49/a_572_375# FILLER_0_4_49/a_124_375#
+ FILLER_0_4_49/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 vdd vss fanout54/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd vdd vss fanout76/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd vdd vss fanout65/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss vdd vss FILLER_0_19_28/a_36_472# FILLER_0_19_28/a_572_375#
+ FILLER_0_19_28/a_124_375# FILLER_0_19_28/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd vdd vss _447_/a_2665_112# _447_/a_448_472#
+ _447_/a_796_472# _447_/a_36_151# _447_/a_1204_472# _447_/a_3041_156# _447_/a_1000_472#
+ _447_/a_1308_423# _447_/a_1456_156# _447_/a_1288_156# _447_/a_2248_156# _447_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_2 vdd vss vdd vss FILLER_0_3_2/a_36_472# FILLER_0_3_2/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ vdd vss _033_ _160_ _165_ vdd vss _378_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ vdd vss _301_/a_36_472# _301_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] vdd vss _232_/a_255_603# _232_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss vdd vss FILLER_0_11_142/a_36_472# FILLER_0_11_142/a_572_375#
+ FILLER_0_11_142/a_124_375# FILLER_0_11_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss vdd vss FILLER_0_2_93/a_36_472# FILLER_0_2_93/a_572_375# FILLER_0_2_93/a_124_375#
+ FILLER_0_2_93/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss vdd vss FILLER_0_17_72/a_1916_375# FILLER_0_17_72/a_1380_472#
+ FILLER_0_17_72/a_3260_375# FILLER_0_17_72/a_36_472# FILLER_0_17_72/a_932_472# FILLER_0_17_72/a_2812_375#
+ FILLER_0_17_72/a_2276_472# FILLER_0_17_72/a_1828_472# FILLER_0_17_72/a_3172_472#
+ FILLER_0_17_72/a_572_375# FILLER_0_17_72/a_2724_472# FILLER_0_17_72/a_124_375# FILLER_0_17_72/a_1468_375#
+ FILLER_0_17_72/a_1020_375# FILLER_0_17_72/a_484_472# FILLER_0_17_72/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss vdd vss FILLER_0_3_172/a_1916_375# FILLER_0_3_172/a_1380_472#
+ FILLER_0_3_172/a_3260_375# FILLER_0_3_172/a_36_472# FILLER_0_3_172/a_932_472# FILLER_0_3_172/a_2812_375#
+ FILLER_0_3_172/a_2276_472# FILLER_0_3_172/a_1828_472# FILLER_0_3_172/a_3172_472#
+ FILLER_0_3_172/a_572_375# FILLER_0_3_172/a_2724_472# FILLER_0_3_172/a_124_375# FILLER_0_3_172/a_1468_375#
+ FILLER_0_3_172/a_1020_375# FILLER_0_3_172/a_484_472# FILLER_0_3_172/a_2364_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] vdd vss _394_/a_244_524# _394_/a_2215_68#
+ _394_/a_56_524# _394_/a_718_524# _394_/a_728_93# _394_/a_1936_472# _394_/a_1336_472#
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 vdd vss fanout55/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss vdd vss FILLER_0_5_212/a_36_472# FILLER_0_5_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd vdd vss fanout77/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd vdd vss _446_/a_2665_112# _446_/a_448_472#
+ _446_/a_796_472# _446_/a_36_151# _446_/a_1204_472# _446_/a_3041_156# _446_/a_1000_472#
+ _446_/a_1308_423# _446_/a_1456_156# _446_/a_1288_156# _446_/a_2248_156# _446_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout66 vss net66 net68 vdd vdd vss fanout66/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ vdd vss _377_/a_36_472# _377_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd vss _011_ _104_ _109_ vdd vss _300_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ vdd vss _231_/a_652_68# _231_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd vdd vss _429_/a_2665_112# _429_/a_448_472#
+ _429_/a_796_472# _429_/a_36_151# _429_/a_1204_472# _429_/a_3041_156# _429_/a_1000_472#
+ _429_/a_1308_423# _429_/a_1456_156# _429_/a_1288_156# _429_/a_2248_156# _429_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd vdd vss input1/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd vdd vss _214_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss vdd vss FILLER_0_7_104/a_1380_472# FILLER_0_7_104/a_36_472#
+ FILLER_0_7_104/a_932_472# FILLER_0_7_104/a_572_375# FILLER_0_7_104/a_124_375# FILLER_0_7_104/a_1468_375#
+ FILLER_0_7_104/a_1020_375# FILLER_0_7_104/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss vdd vss FILLER_0_4_107/a_1380_472# FILLER_0_4_107/a_36_472#
+ FILLER_0_4_107/a_932_472# FILLER_0_4_107/a_572_375# FILLER_0_4_107/a_124_375# FILLER_0_4_107/a_1468_375#
+ FILLER_0_4_107/a_1020_375# FILLER_0_4_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss vdd vss FILLER_0_24_290/a_36_472# FILLER_0_24_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss vdd vss FILLER_0_15_290/a_36_472# FILLER_0_15_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss vdd vss FILLER_0_0_198/a_36_472# FILLER_0_0_198/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd vdd vss fanout78/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd vdd vss fanout56/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd vdd vss fanout67/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd vdd vss _445_/a_2665_112# _445_/a_448_472#
+ _445_/a_796_472# _445_/a_36_151# _445_/a_1204_472# _445_/a_3041_156# _445_/a_1000_472#
+ _445_/a_1308_423# _445_/a_1456_156# _445_/a_1288_156# _445_/a_2248_156# _445_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vss _164_ _163_ vdd vdd vss _376_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd vss _062_ _060_ _061_ vdd vss _230_/a_652_68# _230_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vss vdd vss FILLER_0_5_72/a_1380_472# FILLER_0_5_72/a_36_472# FILLER_0_5_72/a_932_472#
+ FILLER_0_5_72/a_572_375# FILLER_0_5_72/a_124_375# FILLER_0_5_72/a_1468_375# FILLER_0_5_72/a_1020_375#
+ FILLER_0_5_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ _017_ state\[2\] net53 vss net70 vdd vdd vss _428_/a_2665_112# _428_/a_448_472#
+ _428_/a_796_472# _428_/a_36_151# _428_/a_1204_472# _428_/a_3041_156# _428_/a_1000_472#
+ _428_/a_1308_423# _428_/a_1456_156# _428_/a_1288_156# _428_/a_2248_156# _428_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd vss vdd vss FILLER_0_11_64/a_36_472# FILLER_0_11_64/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ vdd vss _359_/a_1492_488# _359_/a_244_68#
+ _359_/a_1044_488# _359_/a_636_68# _359_/a_36_488# gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vss net2 clk vdd vdd vss input2/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output22_I vss net22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 vdd vss _213_/a_255_603# _213_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_177 vdd vss vdd vss FILLER_0_20_177/a_1380_472# FILLER_0_20_177/a_36_472#
+ FILLER_0_20_177/a_932_472# FILLER_0_20_177/a_572_375# FILLER_0_20_177/a_124_375#
+ FILLER_0_20_177/a_1468_375# FILLER_0_20_177/a_1020_375# FILLER_0_20_177/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_206 vdd vss vdd vss FILLER_0_13_206/a_36_472# FILLER_0_13_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss vdd vss FILLER_0_13_228/a_36_472# FILLER_0_13_228/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss vdd vss _392_/a_36_68# _392_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__282__I vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 vss net79 net81 vdd vdd vss fanout79/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_2 vdd vss vdd vss FILLER_0_12_2/a_36_472# FILLER_0_12_2/a_572_375# FILLER_0_12_2/a_124_375#
+ FILLER_0_12_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout68 vss net68 net69 vdd vdd vss fanout68/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 vss net57 net65 vdd vdd vss fanout57/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd vdd vss _444_/a_2665_112# _444_/a_448_472#
+ _444_/a_796_472# _444_/a_36_151# _444_/a_1204_472# _444_/a_3041_156# _444_/a_1000_472#
+ _444_/a_1308_423# _444_/a_1456_156# _444_/a_1288_156# _444_/a_2248_156# _444_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] vdd vss _375_/a_36_68# _375_/a_1612_497#
+ _375_/a_692_497# _375_/a_1388_497# _375_/a_960_497# gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__277__I vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd vss vdd vss FILLER_0_18_139/a_1380_472# FILLER_0_18_139/a_36_472#
+ FILLER_0_18_139/a_932_472# FILLER_0_18_139/a_572_375# FILLER_0_18_139/a_124_375#
+ FILLER_0_18_139/a_1468_375# FILLER_0_18_139/a_1020_375# FILLER_0_18_139/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_161 vdd vss vdd vss FILLER_0_17_161/a_36_472# FILLER_0_17_161/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ _016_ state\[1\] net53 vdd vss net70 vdd vss _427_/a_2665_112# _427_/a_448_472#
+ _427_/a_796_472# _427_/a_36_151# _427_/a_1204_472# _427_/a_3041_156# _427_/a_1000_472#
+ _427_/a_1308_423# _427_/a_2248_156# _427_/a_2560_156# gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_358_ vdd vss _053_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ vdd vss _289_/a_36_472# _289_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd vdd vss input3/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss vdd vss FILLER_0_22_86/a_1380_472# FILLER_0_22_86/a_36_472#
+ FILLER_0_22_86/a_932_472# FILLER_0_22_86/a_572_375# FILLER_0_22_86/a_124_375# FILLER_0_22_86/a_1468_375#
+ FILLER_0_22_86/a_1020_375# FILLER_0_22_86/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss vdd vss FILLER_0_11_101/a_36_472# FILLER_0_11_101/a_572_375#
+ FILLER_0_11_101/a_124_375# FILLER_0_11_101/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss vdd vss FILLER_0_17_64/a_36_472# FILLER_0_17_64/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss vdd vss FILLER_0_3_142/a_36_472# FILLER_0_3_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ vdd vss _391_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 vss net69 net74 vdd vdd vss fanout69/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net58 vss vdd net59 vdd vss fanout58/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_374_ vdd _061_ _056_ _162_ calibrate vss vdd vss _374_/a_36_68# _374_/a_244_472#
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd vdd vss _443_/a_2665_112# _443_/a_448_472#
+ _443_/a_796_472# _443_/a_36_151# _443_/a_1204_472# _443_/a_3041_156# _443_/a_1000_472#
+ _443_/a_1308_423# _443_/a_1456_156# _443_/a_1288_156# _443_/a_2248_156# _443_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_107 vdd vss vdd vss FILLER_0_18_107/a_1916_375# FILLER_0_18_107/a_1380_472#
+ FILLER_0_18_107/a_3260_375# FILLER_0_18_107/a_36_472# FILLER_0_18_107/a_932_472#
+ FILLER_0_18_107/a_2812_375# FILLER_0_18_107/a_2276_472# FILLER_0_18_107/a_1828_472#
+ FILLER_0_18_107/a_3172_472# FILLER_0_18_107/a_572_375# FILLER_0_18_107/a_2724_472#
+ FILLER_0_18_107/a_124_375# FILLER_0_18_107/a_1468_375# FILLER_0_18_107/a_1020_375#
+ FILLER_0_18_107/a_484_472# FILLER_0_18_107/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ vdd vss _288_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ _015_ state\[0\] net64 vss net81 vdd vdd vss _426_/a_2665_112# _426_/a_448_472#
+ _426_/a_796_472# _426_/a_36_151# _426_/a_1204_472# _426_/a_3041_156# _426_/a_1000_472#
+ _426_/a_1308_423# _426_/a_1456_156# _426_/a_1288_156# _426_/a_2248_156# _426_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 vss net4 en vdd vdd vss input4/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_211_ vss net24 _050_ vdd vdd vss _211_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ vdd vss _409_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd vss vdd vss FILLER_0_11_135/a_36_472# FILLER_0_11_135/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vss vdd vss FILLER_0_11_124/a_36_472# FILLER_0_11_124/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss vdd vss FILLER_0_15_282/a_36_472# FILLER_0_15_282/a_572_375#
+ FILLER_0_15_282/a_124_375# FILLER_0_15_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ vdd vss _390_/a_36_68# _390_/a_244_472#
+ _390_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss vdd vss FILLER_0_14_99/a_36_472# FILLER_0_14_99/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 vdd vss fanout59/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ vdd vss _373_/a_438_68# _373_/a_244_68#
+ _373_/a_1254_68# _373_/a_1060_68# _373_/a_632_68# _373_/a_1458_68# gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd vdd vss _442_/a_2665_112# _442_/a_448_472#
+ _442_/a_796_472# _442_/a_36_151# _442_/a_1204_472# _442_/a_3041_156# _442_/a_1000_472#
+ _442_/a_1308_423# _442_/a_1456_156# _442_/a_1288_156# _442_/a_2248_156# _442_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ vdd vss _356_/a_36_472# _356_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ vdd vss _287_/a_36_472# _287_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss vdd vss FILLER_0_11_78/a_36_472# FILLER_0_11_78/a_572_375#
+ FILLER_0_11_78/a_124_375# FILLER_0_11_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd vdd vss input5/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd vdd vss _425_/a_2665_112# _425_/a_448_472#
+ _425_/a_796_472# _425_/a_36_151# _425_/a_1204_472# _425_/a_3041_156# _425_/a_1000_472#
+ _425_/a_1308_423# _425_/a_1456_156# _425_/a_1288_156# _425_/a_2248_156# _425_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 vdd vss _210_/a_255_603# _210_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss vdd vss FILLER_0_20_169/a_36_472# FILLER_0_20_169/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] vdd vss _408_/a_244_524# _408_/a_2215_68#
+ _408_/a_56_524# _408_/a_718_524# _408_/a_728_93# _408_/a_1936_472# _408_/a_1336_472#
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd vdd vss _339_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss vdd vss FILLER_0_21_286/a_36_472# FILLER_0_21_286/a_572_375#
+ FILLER_0_21_286/a_124_375# FILLER_0_21_286/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss vdd vss FILLER_0_12_220/a_1380_472# FILLER_0_12_220/a_36_472#
+ FILLER_0_12_220/a_932_472# FILLER_0_12_220/a_572_375# FILLER_0_12_220/a_124_375#
+ FILLER_0_12_220/a_1468_375# FILLER_0_12_220/a_1020_375# FILLER_0_12_220/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss vdd vss FILLER_0_8_247/a_1380_472# FILLER_0_8_247/a_36_472#
+ FILLER_0_8_247/a_932_472# FILLER_0_8_247/a_572_375# FILLER_0_8_247/a_124_375# FILLER_0_8_247/a_1468_375#
+ FILLER_0_8_247/a_1020_375# FILLER_0_8_247/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 net49 vss vdd net50 vdd vss fanout49/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_206 vdd vss vdd vss FILLER_0_5_206/a_36_472# FILLER_0_5_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd vdd vss _441_/a_2665_112# _441_/a_448_472#
+ _441_/a_796_472# _441_/a_36_151# _441_/a_1204_472# _441_/a_3041_156# _441_/a_1000_472#
+ _441_/a_1308_423# _441_/a_1456_156# _441_/a_1288_156# _441_/a_2248_156# _441_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ vdd vss _372_/a_2590_472# _372_/a_170_472#
+ _372_/a_1602_69# _372_/a_786_69# _372_/a_3126_472# _372_/a_1194_69# _372_/a_3662_472#
+ _372_/a_2034_472# _372_/a_358_69# gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__303__A2 vss _098_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vss vdd vss FILLER_0_17_142/a_36_472# FILLER_0_17_142/a_572_375#
+ FILLER_0_17_142/a_124_375# FILLER_0_17_142/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_54 vdd vss vdd vss FILLER_0_5_54/a_1380_472# FILLER_0_5_54/a_36_472# FILLER_0_5_54/a_932_472#
+ FILLER_0_5_54/a_572_375# FILLER_0_5_54/a_124_375# FILLER_0_5_54/a_1468_375# FILLER_0_5_54/a_1020_375#
+ FILLER_0_5_54/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_355_ vdd vss _149_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd vdd vss _424_/a_2665_112# _424_/a_448_472#
+ _424_/a_796_472# _424_/a_36_151# _424_/a_1204_472# _424_/a_3041_156# _424_/a_1000_472#
+ _424_/a_1308_423# _424_/a_1456_156# _424_/a_1288_156# _424_/a_2248_156# _424_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ vdd vss _005_ _094_ _101_ vdd vss _286_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_123 vdd vss vdd vss FILLER_0_14_123/a_36_472# FILLER_0_14_123/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ vdd vss _407_/a_36_472# _407_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ vdd vss _269_/a_36_472# _269_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss vdd vss FILLER_0_17_56/a_36_472# FILLER_0_17_56/a_572_375#
+ FILLER_0_17_56/a_124_375# FILLER_0_17_56/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vss _032_ _159_ vdd vdd vss _371_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd vdd vss _440_/a_2665_112# _440_/a_448_472#
+ _440_/a_796_472# _440_/a_36_151# _440_/a_1204_472# _440_/a_3041_156# _440_/a_1000_472#
+ _440_/a_1308_423# _440_/a_1456_156# _440_/a_1288_156# _440_/a_2248_156# _440_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd vss vdd vss FILLER_0_5_88/a_36_472# FILLER_0_5_88/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ _012_ net35 net55 vss net72 vdd vdd vss _423_/a_2665_112# _423_/a_448_472#
+ _423_/a_796_472# _423_/a_36_151# _423_/a_1204_472# _423_/a_3041_156# _423_/a_1000_472#
+ _423_/a_1308_423# _423_/a_1456_156# _423_/a_1288_156# _423_/a_2248_156# _423_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ vdd vss _354_/a_49_472# _354_/a_665_69#
+ _354_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_285_ net28 vdd vss _101_ mask\[1\] _099_ vdd vss _285_/a_36_472# _285_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_199_ net20 vss vdd _046_ vdd vss _199_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ vdd vss _337_/a_49_472# _337_/a_665_69#
+ _337_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] vdd vss _406_/a_36_159# gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ vdd vss _268_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss vdd vss FILLER_0_24_274/a_1380_472# FILLER_0_24_274/a_36_472#
+ FILLER_0_24_274/a_932_472# FILLER_0_24_274/a_572_375# FILLER_0_24_274/a_124_375#
+ FILLER_0_24_274/a_1468_375# FILLER_0_24_274/a_1020_375# FILLER_0_24_274/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ vdd vss _370_/a_848_380# _370_/a_1084_68#
+ _370_/a_124_24# _370_/a_1152_472# _370_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss vdd vss FILLER_0_1_266/a_36_472# FILLER_0_1_266/a_572_375#
+ FILLER_0_1_266/a_124_375# FILLER_0_1_266/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_422_ _011_ net34 net61 vss net78 vdd vdd vss _422_/a_2665_112# _422_/a_448_472#
+ _422_/a_796_472# _422_/a_36_151# _422_/a_1204_472# _422_/a_3041_156# _422_/a_1000_472#
+ _422_/a_1308_423# _422_/a_1456_156# _422_/a_1288_156# _422_/a_2248_156# _422_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_353_ vdd vss _148_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss vdd vss FILLER_0_17_133/a_36_472# FILLER_0_17_133/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output36_I vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_284_ vdd vss _004_ _094_ _100_ vdd vss _284_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_198_ vdd vss _046_ mask\[3\] net30 vdd vss _198_/a_255_603# _198_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_336_ vdd vss _138_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] vdd vss _405_/a_255_603# _405_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] vdd vss _267_/a_1792_472# _267_/a_224_472#
+ _267_/a_1568_472# _267_/a_36_472# _267_/a_1120_472# _267_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss vdd vss FILLER_0_6_177/a_36_472# FILLER_0_6_177/a_572_375#
+ FILLER_0_6_177/a_124_375# FILLER_0_6_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ vdd vss _319_/a_234_472# _319_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss vdd vss FILLER_0_8_239/a_36_472# FILLER_0_8_239/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss vdd vss FILLER_0_1_212/a_36_472# FILLER_0_1_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd vdd vss _421_/a_2665_112# _421_/a_448_472#
+ _421_/a_796_472# _421_/a_36_151# _421_/a_1204_472# _421_/a_3041_156# _421_/a_1000_472#
+ _421_/a_1308_423# _421_/a_1456_156# _421_/a_1288_156# _421_/a_2248_156# _421_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ vdd vss _352_/a_49_472# _352_/a_665_69#
+ _352_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ vdd vss _283_/a_36_472# _283_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vdd vss vdd vss FILLER_0_9_142/a_36_472# FILLER_0_9_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vss vdd vss FILLER_0_20_107/a_36_472# FILLER_0_20_107/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ vdd vss _404_/a_36_472# _404_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ vdd vss _335_/a_49_472# _335_/a_665_69#
+ _335_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_266_ vdd vss _055_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_197_ vdd vss net19 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd vss _124_ _115_ _118_ vdd vss _318_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd vss vdd vss FILLER_0_8_24/a_36_472# FILLER_0_8_24/a_572_375# FILLER_0_8_24/a_124_375#
+ FILLER_0_8_24/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss vdd vss FILLER_0_8_2/a_36_472# FILLER_0_8_2/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd vdd vss _420_/a_2665_112# _420_/a_448_472#
+ _420_/a_796_472# _420_/a_36_151# _420_/a_1204_472# _420_/a_3041_156# _420_/a_1000_472#
+ _420_/a_1308_423# _420_/a_1456_156# _420_/a_1288_156# _420_/a_2248_156# _420_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd vdd vss _282_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_334_ vss _137_ _132_ vdd vdd vss _334_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_403_ vdd vss _183_ cal_count\[2\] _176_ vdd vss _403_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vss vdd vss FILLER_0_6_90/a_36_472# FILLER_0_6_90/a_572_375# FILLER_0_6_90/a_124_375#
+ FILLER_0_6_90/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net19 vss vdd _045_ vdd vss _196_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ vdd vss _265_/a_468_472# _265_/a_224_472#
+ _265_/a_244_68# _265_/a_916_472# gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd vss vdd vss FILLER_0_17_38/a_36_472# FILLER_0_17_38/a_572_375#
+ FILLER_0_17_38/a_124_375# FILLER_0_17_38/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_248_ vss _070_ _069_ vdd vdd vss _248_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__409__A2 vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd vdd vss _317_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss vdd vss FILLER_0_2_171/a_36_472# FILLER_0_2_171/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss vdd vss FILLER_0_12_236/a_36_472# FILLER_0_12_236/a_572_375#
+ FILLER_0_12_236/a_124_375# FILLER_0_12_236/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ vdd vss _350_/a_49_472# _350_/a_665_69#
+ _350_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ vdd vss _281_/a_234_472# _281_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd vdd vss _333_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 vdd vss _195_/a_255_603# _195_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] vdd vss _402_/a_244_567# _402_/a_718_527#
+ _402_/a_2172_497# _402_/a_56_567# _402_/a_1948_68# _402_/a_728_93# _402_/a_1296_93#
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss vdd vss FILLER_0_11_109/a_36_472# FILLER_0_11_109/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] vdd vss _264_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss vdd vss FILLER_0_12_50/a_36_472# FILLER_0_12_50/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ vdd vss _247_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate vdd vss _316_/a_848_380# _316_/a_1084_68#
+ _316_/a_124_24# _316_/a_1152_472# _316_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_60 vdd vss vdd vss FILLER_0_23_60/a_36_472# FILLER_0_23_60/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vss vdd vss FILLER_0_15_212/a_1380_472# FILLER_0_15_212/a_36_472#
+ FILLER_0_15_212/a_932_472# FILLER_0_15_212/a_572_375# FILLER_0_15_212/a_124_375#
+ FILLER_0_15_212/a_1468_375# FILLER_0_15_212/a_1020_375# FILLER_0_15_212/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vss vdd vss FILLER_0_8_37/a_36_472# FILLER_0_8_37/a_572_375# FILLER_0_8_37/a_124_375#
+ FILLER_0_8_37/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss vdd vss FILLER_0_17_104/a_1380_472# FILLER_0_17_104/a_36_472#
+ FILLER_0_17_104/a_932_472# FILLER_0_17_104/a_572_375# FILLER_0_17_104/a_124_375#
+ FILLER_0_17_104/a_1468_375# FILLER_0_17_104/a_1020_375# FILLER_0_17_104/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_72 vdd vss vdd vss FILLER_0_15_72/a_36_472# FILLER_0_15_72/a_572_375#
+ FILLER_0_15_72/a_124_375# FILLER_0_15_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd vss vdd vss FILLER_0_1_204/a_36_472# FILLER_0_1_204/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ vdd vss _280_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss vdd vss FILLER_0_14_107/a_1380_472# FILLER_0_14_107/a_36_472#
+ FILLER_0_14_107/a_932_472# FILLER_0_14_107/a_572_375# FILLER_0_14_107/a_124_375#
+ FILLER_0_14_107/a_1468_375# FILLER_0_14_107/a_1020_375# FILLER_0_14_107/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ vdd _180_ _179_ _181_ _174_ vss vdd vss _401_/a_36_68# _401_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_332_ _126_ vdd vss _017_ _127_ _135_ vdd vss _332_/a_36_472# _332_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_194_ vss net8 net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ vdd vss _263_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss vdd vss FILLER_0_5_181/a_36_472# FILLER_0_5_181/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_246_ vss _068_ _055_ vdd vdd vss _246_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss vdd vss _315_/a_36_68# _315_/a_244_497#
+ _315_/a_1657_68# _315_/a_1229_68# _315_/a_716_497# gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_290 vdd vss vdd vss FILLER_0_23_290/a_36_472# FILLER_0_23_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss vdd vss FILLER_0_15_235/a_36_472# FILLER_0_15_235/a_572_375#
+ FILLER_0_15_235/a_124_375# FILLER_0_15_235/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ vdd vss _229_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss vdd vss FILLER_0_18_61/a_36_472# FILLER_0_18_61/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss vdd vss FILLER_0_11_282/a_36_472# FILLER_0_11_282/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss vdd vss FILLER_0_4_213/a_36_472# FILLER_0_4_213/a_572_375#
+ FILLER_0_4_213/a_124_375# FILLER_0_4_213/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ vdd vss _180_ cal_count\[1\] _178_ vdd vss _400_/a_245_68# gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_193_ net18 vss vdd _044_ vdd vss _193_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_331_ _134_ vdd vss _135_ _086_ _132_ vdd vss _331_/a_448_472# _331_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ vdd vss _121_ _085_ _069_ vdd vss _314_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_245_ vdd vss net6 _067_ net67 vdd vss _245_/a_234_472# _245_/a_672_472# gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_206 vdd vss vdd vss FILLER_0_21_206/a_36_472# FILLER_0_21_206/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd vdd vss _228_/a_36_68# gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss vdd vss FILLER_0_7_233/a_36_472# FILLER_0_7_233/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss vdd vss FILLER_0_9_60/a_36_472# FILLER_0_9_60/a_572_375# FILLER_0_9_60/a_124_375#
+ FILLER_0_9_60/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vss vdd vss FILLER_0_13_142/a_1380_472# FILLER_0_13_142/a_36_472#
+ FILLER_0_13_142/a_932_472# FILLER_0_13_142/a_572_375# FILLER_0_13_142/a_124_375#
+ FILLER_0_13_142/a_1468_375# FILLER_0_13_142/a_1020_375# FILLER_0_13_142/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ vdd vss _044_ mask\[1\] net28 vdd vss _192_/a_255_603# _192_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
X_261_ vss _081_ _059_ vdd vdd vss _261_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_330_ vdd vss _134_ _133_ _062_ vdd vss _330_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss vdd vss FILLER_0_12_20/a_36_472# FILLER_0_12_20/a_572_375#
+ FILLER_0_12_20/a_124_375# FILLER_0_12_20/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss vdd vss FILLER_0_5_172/a_36_472# FILLER_0_5_172/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ vdd vss en_co_clk _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__190__I vss _043_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_313_ vdd vss _120_ _059_ _119_ vdd vss _313_/a_255_603# _313_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__257__A1 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd vdd vss _227_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss vdd vss FILLER_0_20_31/a_36_472# FILLER_0_20_31/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss vdd vss FILLER_0_9_72/a_1380_472# FILLER_0_9_72/a_36_472# FILLER_0_9_72/a_932_472#
+ FILLER_0_9_72/a_572_375# FILLER_0_9_72/a_124_375# FILLER_0_9_72/a_1468_375# FILLER_0_9_72/a_1020_375#
+ FILLER_0_9_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss vdd vss FILLER_0_0_96/a_36_472# FILLER_0_0_96/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss vdd vss _260_/a_36_68# _260_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ vdd vss _389_/a_428_148# _389_/a_36_148# gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ vdd vss _312_/a_234_472# _312_/a_672_472#
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd vss net47 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd vss vdd vss FILLER_0_23_282/a_36_472# FILLER_0_23_282/a_572_375#
+ FILLER_0_23_282/a_124_375# FILLER_0_23_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss vdd vss FILLER_0_15_205/a_36_472# FILLER_0_15_205/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss vdd vss FILLER_0_2_165/a_36_472# FILLER_0_2_165/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss vdd vss FILLER_0_18_53/a_36_472# FILLER_0_18_53/a_572_375#
+ FILLER_0_18_53/a_124_375# FILLER_0_18_53/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ vdd vss _226_/a_1044_68# _226_/a_452_68# _226_/a_276_68#
+ _226_/a_860_68# gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_98 vdd vss vdd vss FILLER_0_20_98/a_36_472# FILLER_0_20_98/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_87 vdd vss vdd vss FILLER_0_20_87/a_36_472# FILLER_0_20_87/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss vdd vss FILLER_0_19_171/a_1380_472# FILLER_0_19_171/a_36_472#
+ FILLER_0_19_171/a_932_472# FILLER_0_19_171/a_572_375# FILLER_0_19_171/a_124_375#
+ FILLER_0_19_171/a_1468_375# FILLER_0_19_171/a_1020_375# FILLER_0_19_171/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss vdd vss FILLER_0_15_10/a_36_472# FILLER_0_15_10/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss vdd vss FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_572_375# FILLER_0_15_2/a_124_375#
+ FILLER_0_15_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss vdd vss FILLER_0_22_177/a_1380_472# FILLER_0_22_177/a_36_472#
+ FILLER_0_22_177/a_932_472# FILLER_0_22_177/a_572_375# FILLER_0_22_177/a_124_375#
+ FILLER_0_22_177/a_1468_375# FILLER_0_22_177/a_1020_375# FILLER_0_22_177/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss vdd vss FILLER_0_13_100/a_36_472# FILLER_0_13_100/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss vdd vss FILLER_0_9_105/a_36_472# FILLER_0_9_105/a_572_375#
+ FILLER_0_9_105/a_124_375# FILLER_0_9_105/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ vdd vss _190_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ vdd vss _311_/a_692_473# _311_/a_254_473#
+ _311_/a_66_473# _311_/a_2700_473# _311_/a_1660_473# _311_/a_3220_473# _311_/a_1212_473#
+ _311_/a_2180_473# _311_/a_3740_473# _311_/a_1920_473# gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_242_ net47 vss vdd _066_ vdd vss _242_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_228 vdd vss vdd vss FILLER_0_15_228/a_36_472# FILLER_0_15_228/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss vdd vss FILLER_0_2_111/a_1380_472# FILLER_0_2_111/a_36_472#
+ FILLER_0_2_111/a_932_472# FILLER_0_2_111/a_572_375# FILLER_0_2_111/a_124_375# FILLER_0_2_111/a_1468_375#
+ FILLER_0_2_111/a_1020_375# FILLER_0_2_111/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss vdd vss FILLER_0_2_177/a_36_472# FILLER_0_2_177/a_572_375#
+ FILLER_0_2_177/a_124_375# FILLER_0_2_177/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd vdd vss _225_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss vdd vss FILLER_0_18_76/a_36_472# FILLER_0_18_76/a_572_375#
+ FILLER_0_18_76/a_124_375# FILLER_0_18_76/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ vdd vss _208_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd vdd vss _387_/a_36_113# gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_310_ _090_ vdd vss _117_ _060_ _113_ vdd vss _310_/a_49_472# _310_/a_1133_69# _310_/a_741_69#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_164 vdd vss vdd vss FILLER_0_5_164/a_36_472# FILLER_0_5_164/a_572_375#
+ FILLER_0_5_164/a_124_375# FILLER_0_5_164/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd vss vdd vss FILLER_0_23_88/a_36_472# FILLER_0_23_88/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss vdd vss FILLER_0_23_44/a_1380_472# FILLER_0_23_44/a_36_472#
+ FILLER_0_23_44/a_932_472# FILLER_0_23_44/a_572_375# FILLER_0_23_44/a_124_375# FILLER_0_23_44/a_1468_375#
+ FILLER_0_23_44/a_1020_375# FILLER_0_23_44/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] vdd vss _241_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd vdd vss _439_/a_2665_112# _439_/a_448_472#
+ _439_/a_796_472# _439_/a_36_151# _439_/a_1204_472# _439_/a_3041_156# _439_/a_1000_472#
+ _439_/a_1308_423# _439_/a_1456_156# _439_/a_1288_156# _439_/a_2248_156# _439_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd vss vdd vss FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss vdd vss FILLER_0_3_54/a_36_472# FILLER_0_3_54/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2$1
X_207_ vdd vss _049_ mask\[6\] net33 vdd vss _207_/a_255_603# _207_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss vdd vss FILLER_0_19_195/a_36_472# FILLER_0_19_195/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss vdd vss FILLER_0_0_232/a_36_472# FILLER_0_0_232/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss vdd vss FILLER_0_16_154/a_1380_472# FILLER_0_16_154/a_36_472#
+ FILLER_0_16_154/a_932_472# FILLER_0_16_154/a_572_375# FILLER_0_16_154/a_124_375#
+ FILLER_0_16_154/a_1468_375# FILLER_0_16_154/a_1020_375# FILLER_0_16_154/a_484_472#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss vdd vss FILLER_0_20_2/a_36_472# FILLER_0_20_2/a_572_375# FILLER_0_20_2/a_124_375#
+ FILLER_0_20_2/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ vdd vss _386_/a_848_380# _386_/a_1084_68#
+ _386_/a_124_24# _386_/a_1152_472# _386_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss vdd vss FILLER_0_5_198/a_36_472# FILLER_0_5_198/a_572_375#
+ FILLER_0_5_198/a_124_375# FILLER_0_5_198/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_240_ vdd vss net41 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_282 vdd vss vdd vss FILLER_0_17_282/a_36_472# FILLER_0_17_282/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_274 vdd vss vdd vss FILLER_0_23_274/a_36_472# FILLER_0_23_274/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd vdd vss _438_/a_2665_112# _438_/a_448_472#
+ _438_/a_796_472# _438_/a_36_151# _438_/a_1204_472# _438_/a_3041_156# _438_/a_1000_472#
+ _438_/a_1308_423# _438_/a_1456_156# _438_/a_1288_156# _438_/a_2248_156# _438_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ vdd vss _369_/a_36_68# _369_/a_244_472#
+ _369_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss vdd vss FILLER_0_14_263/a_36_472# FILLER_0_14_263/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] vdd vss _223_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss vdd vss FILLER_0_9_290/a_36_472# FILLER_0_9_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss vdd vss FILLER_0_0_266/a_36_472# FILLER_0_0_266/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss vdd vss _385_/a_36_68# _385_/a_244_472# gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ vdd vss _299_/a_36_472# _299_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd vdd vss _437_/a_2665_112# _437_/a_448_472#
+ _437_/a_796_472# _437_/a_36_151# _437_/a_1204_472# _437_/a_3041_156# _437_/a_1000_472#
+ _437_/a_1308_423# _437_/a_1456_156# _437_/a_1288_156# _437_/a_2248_156# _437_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_78 vdd vss vdd vss FILLER_0_3_78/a_36_472# FILLER_0_3_78/a_572_375# FILLER_0_3_78/a_124_375#
+ FILLER_0_3_78/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_368_ vdd vss trim_mask\[4\] _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_222_ vdd vss net38 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ vdd vss _205_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss vdd vss FILLER_0_19_142/a_36_472# FILLER_0_19_142/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd vdd vss _453_/a_2665_112# _453_/a_448_472#
+ _453_/a_796_472# _453_/a_36_151# _453_/a_1204_472# _453_/a_3041_156# _453_/a_1000_472#
+ _453_/a_1308_423# _453_/a_1456_156# _453_/a_1288_156# _453_/a_2248_156# _453_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ vdd vss _384_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss vdd vss FILLER_0_10_107/a_36_472# FILLER_0_10_107/a_572_375#
+ FILLER_0_10_107/a_124_375# FILLER_0_10_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ vdd vss _298_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd vdd vss _436_/a_2665_112# _436_/a_448_472#
+ _436_/a_796_472# _436_/a_36_151# _436_/a_1204_472# _436_/a_3041_156# _436_/a_1000_472#
+ _436_/a_1308_423# _436_/a_1456_156# _436_/a_1288_156# _436_/a_2248_156# _436_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ vdd vss _367_/a_36_68# _367_/a_244_472#
+ _367_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss vdd vss FILLER_0_13_80/a_36_472# FILLER_0_13_80/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss vdd vss FILLER_0_1_192/a_36_472# FILLER_0_1_192/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd vss vdd vss FILLER_0_9_270/a_36_472# FILLER_0_9_270/a_572_375#
+ FILLER_0_9_270/a_124_375# FILLER_0_9_270/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vss net38 _054_ vdd vdd vss _221_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ _008_ net31 net60 vss net77 vdd vdd vss _419_/a_2665_112# _419_/a_448_472#
+ _419_/a_796_472# _419_/a_36_151# _419_/a_1204_472# _419_/a_3041_156# _419_/a_1000_472#
+ _419_/a_1308_423# _419_/a_1456_156# _419_/a_1288_156# _419_/a_2248_156# _419_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 vdd vss _204_/a_255_603# _204_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss vdd vss FILLER_0_20_15/a_1380_472# FILLER_0_20_15/a_36_472#
+ FILLER_0_20_15/a_932_472# FILLER_0_20_15/a_572_375# FILLER_0_20_15/a_124_375# FILLER_0_20_15/a_1468_375#
+ FILLER_0_20_15/a_1020_375# FILLER_0_20_15/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss vdd vss FILLER_0_19_187/a_36_472# FILLER_0_19_187/a_572_375#
+ FILLER_0_19_187/a_124_375# FILLER_0_19_187/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss vdd vss FILLER_0_3_221/a_1380_472# FILLER_0_3_221/a_36_472#
+ FILLER_0_3_221/a_932_472# FILLER_0_3_221/a_572_375# FILLER_0_3_221/a_124_375# FILLER_0_3_221/a_1468_375#
+ FILLER_0_3_221/a_1020_375# FILLER_0_3_221/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss vdd vss FILLER_0_15_59/a_36_472# FILLER_0_15_59/a_572_375#
+ FILLER_0_15_59/a_124_375# FILLER_0_15_59/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd vss vdd vss FILLER_0_6_79/a_36_472# FILLER_0_6_79/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 vdd vss _452_/a_448_472# _452_/a_36_151#
+ _452_/a_1293_527# _452_/a_3081_151# _452_/a_1284_156# _452_/a_1040_527# _452_/a_1353_112#
+ _452_/a_836_156# _452_/a_1697_156# _452_/a_2449_156# _452_/a_3129_107# _452_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ vdd vss _383_/a_36_472# _383_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ vdd vss _297_/a_36_472# _297_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd vdd vss _435_/a_2665_112# _435_/a_448_472#
+ _435_/a_796_472# _435_/a_36_151# _435_/a_1204_472# _435_/a_3041_156# _435_/a_1000_472#
+ _435_/a_1308_423# _435_/a_1456_156# _435_/a_1288_156# _435_/a_2248_156# _435_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A2 vss cal_count\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ vdd vss trim_mask\[3\] _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_127 vdd vss vdd vss FILLER_0_2_127/a_36_472# FILLER_0_2_127/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vss vdd vss FILLER_0_18_37/a_1380_472# FILLER_0_18_37/a_36_472#
+ FILLER_0_18_37/a_932_472# FILLER_0_18_37/a_572_375# FILLER_0_18_37/a_124_375# FILLER_0_18_37/a_1468_375#
+ FILLER_0_18_37/a_1020_375# FILLER_0_18_37/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vss vdd vss FILLER_0_9_282/a_36_472# FILLER_0_9_282/a_572_375#
+ FILLER_0_9_282/a_124_375# FILLER_0_9_282/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd vss _054_ trim_val\[0\] _053_ vdd vss _220_/a_255_603# _220_/a_67_603#
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_349_ vdd vss _146_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _007_ net30 net60 vss net77 vdd vdd vss _418_/a_2665_112# _418_/a_448_472#
+ _418_/a_796_472# _418_/a_36_151# _418_/a_1204_472# _418_/a_3041_156# _418_/a_1000_472#
+ _418_/a_1308_423# _418_/a_1456_156# _418_/a_1288_156# _418_/a_2248_156# _418_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output21_I vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss vdd vss FILLER_0_19_155/a_36_472# FILLER_0_19_155/a_572_375#
+ FILLER_0_19_155/a_124_375# FILLER_0_19_155/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss vdd vss FILLER_0_19_111/a_36_472# FILLER_0_19_111/a_572_375#
+ FILLER_0_19_111/a_124_375# FILLER_0_19_111/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss vdd vss FILLER_0_22_128/a_1916_375# FILLER_0_22_128/a_1380_472#
+ FILLER_0_22_128/a_3260_375# FILLER_0_22_128/a_36_472# FILLER_0_22_128/a_932_472#
+ FILLER_0_22_128/a_2812_375# FILLER_0_22_128/a_2276_472# FILLER_0_22_128/a_1828_472#
+ FILLER_0_22_128/a_3172_472# FILLER_0_22_128/a_572_375# FILLER_0_22_128/a_2724_472#
+ FILLER_0_22_128/a_124_375# FILLER_0_22_128/a_1468_375# FILLER_0_22_128/a_1020_375#
+ FILLER_0_22_128/a_484_472# FILLER_0_22_128/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss vdd vss FILLER_0_15_180/a_36_472# FILLER_0_15_180/a_572_375#
+ FILLER_0_15_180/a_124_375# FILLER_0_15_180/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss vdd vss FILLER_0_21_150/a_36_472# FILLER_0_21_150/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss vdd vss FILLER_0_6_47/a_1916_375# FILLER_0_6_47/a_1380_472#
+ FILLER_0_6_47/a_3260_375# FILLER_0_6_47/a_36_472# FILLER_0_6_47/a_932_472# FILLER_0_6_47/a_2812_375#
+ FILLER_0_6_47/a_2276_472# FILLER_0_6_47/a_1828_472# FILLER_0_6_47/a_3172_472# FILLER_0_6_47/a_572_375#
+ FILLER_0_6_47/a_2724_472# FILLER_0_6_47/a_124_375# FILLER_0_6_47/a_1468_375# FILLER_0_6_47/a_1020_375#
+ FILLER_0_6_47/a_484_472# FILLER_0_6_47/a_2364_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 vdd vss _451_/a_448_472# _451_/a_36_151#
+ _451_/a_1293_527# _451_/a_3081_151# _451_/a_1284_156# _451_/a_1040_527# _451_/a_1353_112#
+ _451_/a_836_156# _451_/a_1697_156# _451_/a_2449_156# _451_/a_3129_107# _451_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_28 vdd vss vdd vss FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd vss _035_ _160_ _167_ vdd vss _382_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss vdd vss FILLER_0_18_209/a_36_472# FILLER_0_18_209/a_572_375#
+ FILLER_0_18_209/a_124_375# FILLER_0_18_209/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss vdd vss FILLER_0_5_136/a_36_472# FILLER_0_5_136/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ vdd vss _296_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd vdd vss _434_/a_2665_112# _434_/a_448_472#
+ _434_/a_796_472# _434_/a_36_151# _434_/a_1204_472# _434_/a_3041_156# _434_/a_1000_472#
+ _434_/a_1308_423# _434_/a_1456_156# _434_/a_1288_156# _434_/a_2248_156# _434_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ vdd vss _365_/a_36_68# _365_/a_244_472#
+ _365_/a_692_472# gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ vdd vss _348_/a_49_472# _348_/a_665_69#
+ _348_/a_257_69# gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd vdd vss _417_/a_2665_112# _417_/a_448_472#
+ _417_/a_796_472# _417_/a_36_151# _417_/a_1204_472# _417_/a_3041_156# _417_/a_1000_472#
+ _417_/a_1308_423# _417_/a_1456_156# _417_/a_1288_156# _417_/a_2248_156# _417_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_279_ vdd vss _096_ _090_ state\[1\] vdd vss _279_/a_652_68# _279_/a_244_68# gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_231 vdd vss vdd vss FILLER_0_6_231/a_36_472# FILLER_0_6_231/a_572_375#
+ FILLER_0_6_231/a_124_375# FILLER_0_6_231/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ vdd vss _202_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output14_I vss net14 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd vss vdd vss FILLER_0_4_91/a_36_472# FILLER_0_4_91/a_572_375# FILLER_0_4_91/a_124_375#
+ FILLER_0_4_91/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_94 vdd vss vdd vss FILLER_0_10_94/a_36_472# FILLER_0_10_94/a_572_375#
+ FILLER_0_10_94/a_124_375# FILLER_0_10_94/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss vdd vss FILLER_0_3_212/a_36_472# FILLER_0_3_212/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss vdd vss FILLER_0_19_134/a_36_472# FILLER_0_19_134/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss vdd vss FILLER_0_16_115/a_36_472# FILLER_0_16_115/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss vdd vss FILLER_0_22_107/a_36_472# FILLER_0_22_107/a_572_375#
+ FILLER_0_22_107/a_124_375# FILLER_0_22_107/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss vdd vss FILLER_0_21_60/a_36_472# FILLER_0_21_60/a_572_375#
+ FILLER_0_21_60/a_124_375# FILLER_0_21_60/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss vdd vss FILLER_0_6_37/a_36_472# FILLER_0_6_37/a_124_375# gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd vss vdd vss FILLER_0_8_156/a_36_472# FILLER_0_8_156/a_572_375#
+ FILLER_0_8_156/a_124_375# FILLER_0_8_156/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I vss rstn vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__243__I vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 vdd vss _450_/a_448_472# _450_/a_36_151#
+ _450_/a_1293_527# _450_/a_3081_151# _450_/a_1284_156# _450_/a_1040_527# _450_/a_1353_112#
+ _450_/a_836_156# _450_/a_1697_156# _450_/a_2449_156# _450_/a_3129_107# _450_/a_2225_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xoutput40 trim[2] net40 vdd vss vdd vss output40/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ vdd vss _381_/a_36_472# _381_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_148 vdd vss vdd vss FILLER_0_5_148/a_36_472# FILLER_0_5_148/a_572_375#
+ FILLER_0_5_148/a_124_375# FILLER_0_5_148/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd vdd vss _433_/a_2665_112# _433_/a_448_472#
+ _433_/a_796_472# _433_/a_36_151# _433_/a_1204_472# _433_/a_3041_156# _433_/a_1000_472#
+ _433_/a_1308_423# _433_/a_1456_156# _433_/a_1288_156# _433_/a_2248_156# _433_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ vdd vss _295_/a_36_472# _295_/a_244_68#
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss vdd vss FILLER_0_14_235/a_36_472# FILLER_0_14_235/a_572_375#
+ FILLER_0_14_235/a_124_375# FILLER_0_14_235/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss vdd vss FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_572_375#
+ FILLER_0_13_72/a_124_375# FILLER_0_13_72/a_484_472# gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_347_ vdd vss _145_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 vdd vss _278_/a_36_160# gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_290 vdd vss vdd vss FILLER_0_13_290/a_36_472# FILLER_0_13_290/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ _005_ net28 net62 vss net79 vdd vdd vss _416_/a_2665_112# _416_/a_448_472#
+ _416_/a_796_472# _416_/a_36_151# _416_/a_1204_472# _416_/a_3041_156# _416_/a_1000_472#
+ _416_/a_1308_423# _416_/a_1456_156# _416_/a_1288_156# _416_/a_2248_156# _416_/a_2560_156#
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_201_ vdd vss _047_ mask\[4\] net31 vdd vss _201_/a_255_603# _201_/a_67_603# gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 result[3] net30 vdd vss vdd vss output30/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_196 vdd vss vdd vss FILLER_0_12_196/a_36_472# FILLER_0_12_196/a_124_375#
+ gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 clkc net6 vdd vss vdd vss output6/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss vdd vss output41/a_224_472# gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ vdd vss _380_/a_224_472# gf180mcu_fd_sc_mcu7t5v0__nor2_1
C0 FILLER_0_5_128/a_124_375# _360_/a_36_160# 0.005705f
C1 fanout81/a_36_160# vss 0.02458f
C2 net50 FILLER_0_7_59/a_572_375# 0.009554f
C3 _422_/a_36_151# vdd 0.177717f
C4 _028_ _439_/a_1000_472# 0.003267f
C5 net63 FILLER_0_17_218/a_36_472# 0.003889f
C6 cal_count\[1\] _043_ 0.002223f
C7 net44 FILLER_0_15_10/a_124_375# 0.009108f
C8 _062_ _060_ 0.032472f
C9 _426_/a_796_472# vdd 0.007178f
C10 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_36_472# 0.012267f
C11 _265_/a_244_68# cal_itt\[0\] 0.003127f
C12 ctlp[2] mask\[7\] 0.036719f
C13 _093_ FILLER_0_18_107/a_124_375# 0.008393f
C14 _131_ _182_ 0.113302f
C15 trim_mask\[1\] net14 0.024935f
C16 _087_ FILLER_0_3_172/a_1916_375# 0.001223f
C17 FILLER_0_15_282/a_124_375# vdd 0.011964f
C18 _446_/a_1204_472# net40 0.026414f
C19 _178_ vss 0.150839f
C20 _086_ FILLER_0_5_181/a_36_472# 0.013437f
C21 _081_ cal_itt\[1\] 0.009747f
C22 FILLER_0_11_101/a_572_375# vdd 0.023482f
C23 _132_ _451_/a_448_472# 0.001197f
C24 _064_ net49 0.377675f
C25 FILLER_0_19_47/a_36_472# _012_ 0.001667f
C26 _185_ cal_count\[1\] 0.001949f
C27 net69 _441_/a_36_151# 0.035817f
C28 _120_ _389_/a_36_148# 0.022887f
C29 FILLER_0_17_104/a_1380_472# FILLER_0_16_115/a_124_375# 0.001723f
C30 trim_mask\[3\] _157_ 0.052956f
C31 net52 FILLER_0_3_142/a_124_375# 0.002239f
C32 _447_/a_2248_156# _030_ 0.001588f
C33 ctln[4] net75 0.00718f
C34 _003_ FILLER_0_5_181/a_124_375# 0.009929f
C35 _305_/a_36_159# net59 0.007898f
C36 _064_ net68 0.059889f
C37 trim_val\[2\] _036_ 0.279133f
C38 output8/a_224_472# net82 0.002936f
C39 vss _022_ 0.067509f
C40 _321_/a_170_472# _121_ 0.007364f
C41 _176_ _055_ 0.001694f
C42 net71 _437_/a_448_472# 0.060858f
C43 net63 FILLER_0_15_212/a_124_375# 0.001597f
C44 _064_ _445_/a_1204_472# 0.007445f
C45 FILLER_0_15_235/a_36_472# FILLER_0_15_228/a_36_472# 0.002765f
C46 _447_/a_796_472# _036_ 0.006511f
C47 _306_/a_36_68# _055_ 0.006686f
C48 cal_itt\[3\] vss 0.15522f
C49 FILLER_0_16_154/a_1380_472# vss 0.003609f
C50 _175_ cal_count\[1\] 0.203153f
C51 FILLER_0_3_172/a_3260_375# net21 0.049606f
C52 _408_/a_728_93# net40 0.084147f
C53 output34/a_224_472# _099_ 0.001498f
C54 FILLER_0_5_109/a_484_472# _153_ 0.071582f
C55 _152_ vdd 0.354509f
C56 _081_ vss 0.733408f
C57 _414_/a_1308_423# net22 0.011978f
C58 net75 FILLER_0_8_247/a_932_472# 0.006746f
C59 result[9] FILLER_0_24_274/a_36_472# 0.009425f
C60 _079_ _001_ 0.082209f
C61 result[4] net61 0.023257f
C62 _325_/a_224_472# _130_ 0.001685f
C63 FILLER_0_7_104/a_1380_472# vdd 0.011752f
C64 FILLER_0_21_142/a_36_472# vdd 0.111749f
C65 FILLER_0_12_136/a_1468_375# state\[2\] 0.035275f
C66 FILLER_0_3_78/a_124_375# _164_ 0.023555f
C67 fanout82/a_36_113# net82 0.003741f
C68 FILLER_0_17_56/a_124_375# _041_ 0.001489f
C69 FILLER_0_14_99/a_36_472# net14 0.036527f
C70 _053_ FILLER_0_7_146/a_36_472# 0.001014f
C71 net73 FILLER_0_18_107/a_1828_472# 0.01544f
C72 output42/a_224_472# _236_/a_36_160# 0.001892f
C73 net75 _426_/a_796_472# 0.003146f
C74 _318_/a_224_472# vdd 0.001873f
C75 _081_ FILLER_0_6_177/a_36_472# 0.00483f
C76 _043_ FILLER_0_13_72/a_124_375# 0.013517f
C77 FILLER_0_16_73/a_484_472# FILLER_0_17_72/a_572_375# 0.001723f
C78 _074_ _312_/a_234_472# 0.005755f
C79 FILLER_0_18_107/a_484_472# vdd 0.035309f
C80 FILLER_0_18_107/a_36_472# vss 0.003245f
C81 _420_/a_36_151# FILLER_0_23_290/a_124_375# 0.026277f
C82 _070_ _385_/a_36_68# 0.049178f
C83 _014_ FILLER_0_7_233/a_124_375# 0.00143f
C84 FILLER_0_19_195/a_36_472# _202_/a_36_160# 0.002647f
C85 net52 FILLER_0_9_72/a_1380_472# 0.003507f
C86 FILLER_0_20_2/a_572_375# net43 0.051705f
C87 _115_ _129_ 0.021405f
C88 _116_ _061_ 0.04837f
C89 net27 FILLER_0_12_236/a_36_472# 0.005414f
C90 net54 FILLER_0_22_128/a_36_472# 0.020739f
C91 _149_ _437_/a_36_151# 0.037766f
C92 FILLER_0_18_139/a_36_472# _145_ 0.002415f
C93 FILLER_0_18_37/a_1380_472# vss 0.002042f
C94 trim_val\[0\] vdd 0.056059f
C95 FILLER_0_16_89/a_932_472# vdd 0.002218f
C96 FILLER_0_16_89/a_484_472# vss -0.001894f
C97 _421_/a_448_472# net77 0.003958f
C98 _014_ vdd 0.035382f
C99 net15 FILLER_0_23_60/a_124_375# 0.038706f
C100 net69 _367_/a_244_472# 0.001708f
C101 _442_/a_2248_156# _153_ 0.0011f
C102 net74 FILLER_0_2_127/a_124_375# 0.001389f
C103 _086_ vss 0.615299f
C104 _010_ _419_/a_1000_472# 0.001598f
C105 _187_ _392_/a_36_68# 0.058263f
C106 _425_/a_796_472# calibrate 0.025807f
C107 net52 fanout52/a_36_160# 0.036543f
C108 _253_/a_36_68# net82 0.016638f
C109 _063_ _164_ 0.326812f
C110 ctln[7] _442_/a_2560_156# 0.001742f
C111 _414_/a_36_151# _072_ 0.033026f
C112 FILLER_0_20_169/a_124_375# _098_ 0.019219f
C113 _089_ vss 0.018272f
C114 _003_ vdd 0.032367f
C115 mask\[3\] _069_ 0.025564f
C116 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_124_375# 0.001597f
C117 net34 _199_/a_36_160# 0.026709f
C118 _011_ _422_/a_1000_472# 0.005583f
C119 _136_ vdd 1.020301f
C120 _119_ vss 0.22921f
C121 _000_ FILLER_0_3_221/a_1380_472# 0.025567f
C122 _086_ FILLER_0_6_177/a_36_472# 0.064045f
C123 _057_ _267_/a_1120_472# 0.001833f
C124 net21 vdd 1.653552f
C125 _070_ FILLER_0_7_233/a_124_375# 0.004917f
C126 trim_mask\[4\] _241_/a_224_472# 0.009431f
C127 net7 _447_/a_36_151# 0.002494f
C128 _430_/a_36_151# vss 0.011779f
C129 _133_ _134_ 0.015205f
C130 fanout53/a_36_160# fanout56/a_36_113# 0.001636f
C131 FILLER_0_22_177/a_1468_375# mask\[6\] 0.002149f
C132 _242_/a_36_160# _169_ 0.051038f
C133 _004_ result[1] 0.005653f
C134 _005_ vss 0.01812f
C135 net18 _416_/a_1204_472# 0.027218f
C136 mask\[5\] net31 0.017182f
C137 FILLER_0_9_28/a_1380_472# _120_ 0.00154f
C138 _070_ vdd 1.546772f
C139 _449_/a_1308_423# vss 0.027539f
C140 net50 FILLER_0_6_90/a_572_375# 0.010099f
C141 FILLER_0_6_239/a_124_375# _074_ 0.010359f
C142 result[0] net64 0.09782f
C143 net31 FILLER_0_18_209/a_572_375# 0.001813f
C144 _176_ _315_/a_36_68# 0.003811f
C145 FILLER_0_12_220/a_932_472# vss 0.003677f
C146 FILLER_0_12_220/a_1380_472# vdd 0.002025f
C147 _356_/a_36_472# vdd 0.016338f
C148 net55 FILLER_0_18_37/a_484_472# 0.006153f
C149 _322_/a_692_472# net74 0.003192f
C150 net75 _014_ 0.204357f
C151 FILLER_0_17_72/a_2364_375# vdd 0.002455f
C152 FILLER_0_17_72/a_1916_375# vss 0.001345f
C153 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_1020_375# 0.026339f
C154 net23 FILLER_0_16_154/a_484_472# 0.001369f
C155 output29/a_224_472# _416_/a_2665_112# 0.011048f
C156 FILLER_0_24_96/a_124_375# ctlp[7] 0.004486f
C157 output36/a_224_472# _045_ 0.041236f
C158 FILLER_0_8_247/a_1020_375# calibrate 0.008393f
C159 _398_/a_36_113# net3 0.099638f
C160 _142_ net23 0.037306f
C161 net16 FILLER_0_18_53/a_36_472# 0.001532f
C162 _077_ _059_ 0.020736f
C163 _061_ _117_ 0.046662f
C164 FILLER_0_22_86/a_1020_375# vdd 0.008761f
C165 net38 _450_/a_1293_527# 0.001307f
C166 net52 _443_/a_448_472# 0.050192f
C167 ctlp[1] vss 0.32843f
C168 _419_/a_1000_472# vdd 0.004107f
C169 _033_ FILLER_0_6_47/a_36_472# 0.001185f
C170 net57 _163_ 0.759175f
C171 _140_ _348_/a_257_69# 0.001089f
C172 result[4] output31/a_224_472# 0.049147f
C173 net80 FILLER_0_22_177/a_932_472# 0.002472f
C174 _104_ _291_/a_36_160# 0.006129f
C175 _091_ net36 0.067629f
C176 fanout81/a_36_160# net4 0.002848f
C177 FILLER_0_9_142/a_36_472# vdd 0.107619f
C178 FILLER_0_9_142/a_124_375# vss 0.006851f
C179 _453_/a_1308_423# _042_ 0.001778f
C180 _453_/a_448_472# net51 0.006397f
C181 FILLER_0_24_63/a_124_375# output26/a_224_472# 0.00515f
C182 _402_/a_1296_93# cal_count\[1\] 0.004472f
C183 _348_/a_49_472# _146_ 0.001552f
C184 _411_/a_448_472# net8 0.04545f
C185 _326_/a_36_160# vdd 0.066545f
C186 net53 vss 0.426484f
C187 _115_ _219_/a_36_160# 0.001218f
C188 FILLER_0_4_107/a_124_375# net47 0.004586f
C189 FILLER_0_24_96/a_124_375# net25 0.008342f
C190 _057_ _074_ 0.013823f
C191 net34 net23 0.058486f
C192 net15 _441_/a_796_472# 0.021664f
C193 net34 FILLER_0_22_128/a_1916_375# 0.04185f
C194 FILLER_0_1_266/a_36_472# net9 0.041635f
C195 _045_ vdd 0.246567f
C196 _437_/a_2248_156# vdd 0.054674f
C197 output37/a_224_472# net64 0.110037f
C198 _449_/a_796_472# net72 0.00138f
C199 _449_/a_36_151# net55 0.003388f
C200 _431_/a_2665_112# vss 0.033886f
C201 FILLER_0_9_223/a_36_472# _246_/a_36_68# 0.006596f
C202 net15 _447_/a_36_151# 0.001598f
C203 FILLER_0_4_177/a_572_375# net76 0.009573f
C204 FILLER_0_4_213/a_36_472# vss 0.003969f
C205 FILLER_0_4_213/a_484_472# vdd 0.007084f
C206 _053_ _414_/a_2560_156# 0.008732f
C207 _390_/a_36_68# net14 0.010844f
C208 _448_/a_36_151# FILLER_0_1_192/a_36_472# 0.008172f
C209 state\[0\] _128_ 0.228492f
C210 net63 _434_/a_36_151# 0.005153f
C211 net54 _436_/a_2560_156# 0.010748f
C212 net55 FILLER_0_17_72/a_1020_375# 0.049648f
C213 ctlp[8] mask\[8\] 0.001554f
C214 _412_/a_2665_112# fanout59/a_36_160# 0.016426f
C215 _446_/a_1000_472# net66 0.006158f
C216 net47 FILLER_0_5_148/a_36_472# 0.004409f
C217 _413_/a_2560_156# net21 0.002416f
C218 _192_/a_67_603# vdd 0.027014f
C219 fanout80/a_36_113# FILLER_0_15_205/a_36_472# 0.010419f
C220 net27 FILLER_0_9_290/a_36_472# 0.006729f
C221 net31 net30 0.130396f
C222 _413_/a_796_472# net65 0.006888f
C223 FILLER_0_5_72/a_124_375# net49 0.001158f
C224 _430_/a_2665_112# fanout63/a_36_160# 0.010365f
C225 net4 _081_ 0.02226f
C226 net54 _433_/a_2665_112# 0.047439f
C227 net54 FILLER_0_18_139/a_1020_375# 0.003589f
C228 _077_ _453_/a_2248_156# 0.013877f
C229 _056_ _310_/a_49_472# 0.003286f
C230 _340_/a_36_160# _140_ 0.062613f
C231 FILLER_0_4_185/a_124_375# _087_ 0.120668f
C232 _043_ FILLER_0_15_180/a_124_375# 0.003099f
C233 FILLER_0_21_125/a_36_472# vss 0.00143f
C234 FILLER_0_21_125/a_484_472# vdd 0.002728f
C235 mask\[4\] _291_/a_36_160# 0.00591f
C236 FILLER_0_19_47/a_124_375# _052_ 0.019401f
C237 FILLER_0_11_78/a_124_375# vss 0.006233f
C238 FILLER_0_11_78/a_572_375# vdd -0.006646f
C239 FILLER_0_20_193/a_36_472# _098_ 0.006652f
C240 FILLER_0_5_72/a_484_472# _029_ 0.004625f
C241 FILLER_0_5_72/a_1020_375# trim_mask\[1\] 0.010728f
C242 net15 FILLER_0_6_47/a_2724_472# 0.006158f
C243 FILLER_0_6_47/a_1468_375# vss 0.003462f
C244 FILLER_0_6_47/a_1916_375# vdd -0.014642f
C245 _343_/a_665_69# mask\[3\] 0.001405f
C246 output10/a_224_472# net19 0.037774f
C247 net19 _009_ 0.055383f
C248 net26 _423_/a_796_472# 0.001077f
C249 FILLER_0_4_123/a_36_472# net69 0.001015f
C250 output16/a_224_472# vss 0.009875f
C251 _444_/a_36_151# _054_ 0.011342f
C252 FILLER_0_13_206/a_36_472# net21 0.00171f
C253 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1380_472# 0.013276f
C254 _104_ _108_ 0.02837f
C255 _301_/a_36_472# vss 0.003975f
C256 FILLER_0_12_50/a_124_375# vss 0.004123f
C257 FILLER_0_12_50/a_36_472# vdd 0.012805f
C258 vdd _450_/a_2449_156# 0.003646f
C259 _016_ _095_ 0.034744f
C260 FILLER_0_5_128/a_124_375# _159_ 0.003644f
C261 _059_ net37 0.011845f
C262 _091_ FILLER_0_20_169/a_36_472# 0.007537f
C263 output48/a_224_472# net37 0.095886f
C264 FILLER_0_17_218/a_124_375# _069_ 0.003162f
C265 _188_ _453_/a_36_151# 0.03354f
C266 _422_/a_1308_423# _108_ 0.019345f
C267 _021_ vdd 0.022473f
C268 _256_/a_36_68# _072_ 0.027152f
C269 FILLER_0_21_286/a_124_375# net18 0.015582f
C270 _413_/a_796_472# net59 0.006163f
C271 _115_ FILLER_0_10_107/a_572_375# 0.040198f
C272 _396_/a_224_472# net36 0.00114f
C273 _098_ FILLER_0_16_154/a_1020_375# 0.003386f
C274 _419_/a_36_151# net77 0.163616f
C275 FILLER_0_9_60/a_484_472# vss 0.005321f
C276 _449_/a_448_472# FILLER_0_11_64/a_36_472# 0.001462f
C277 _204_/a_67_603# vss 0.010366f
C278 _091_ _432_/a_2248_156# 0.007123f
C279 fanout72/a_36_113# vss 0.053396f
C280 net62 FILLER_0_15_290/a_36_472# 0.009046f
C281 net28 _195_/a_67_603# 0.012984f
C282 ctln[7] output15/a_224_472# 0.00838f
C283 _072_ _395_/a_36_488# 0.024944f
C284 net3 cal_count\[2\] 0.119728f
C285 net34 net33 0.509436f
C286 ctlp[4] ctlp[3] 0.027598f
C287 _030_ _160_ 0.063581f
C288 net66 _034_ 0.139638f
C289 net49 _166_ 0.007445f
C290 net76 net22 0.118787f
C291 FILLER_0_23_282/a_572_375# vdd -0.013698f
C292 FILLER_0_23_282/a_124_375# vss 0.005048f
C293 FILLER_0_4_197/a_1380_472# net59 0.022002f
C294 net74 _062_ 0.062376f
C295 FILLER_0_18_2/a_2276_472# net38 0.002313f
C296 net20 output11/a_224_472# 0.036556f
C297 net58 _264_/a_224_472# 0.001803f
C298 net48 cal_itt\[0\] 0.006171f
C299 FILLER_0_21_28/a_2276_472# _012_ 0.023696f
C300 output47/a_224_472# vss 0.002843f
C301 result[8] _011_ 0.001294f
C302 _431_/a_2248_156# FILLER_0_17_142/a_572_375# 0.006739f
C303 _445_/a_1308_423# _034_ 0.002494f
C304 net27 FILLER_0_10_247/a_36_472# 0.016681f
C305 _433_/a_448_472# _022_ 0.074451f
C306 FILLER_0_11_109/a_36_472# vss 0.003131f
C307 _150_ net36 0.108945f
C308 trimb[1] net40 0.00126f
C309 FILLER_0_4_49/a_124_375# _232_/a_67_603# 0.002082f
C310 _414_/a_2248_156# net21 0.00415f
C311 FILLER_0_12_136/a_484_472# _127_ 0.005549f
C312 FILLER_0_2_93/a_572_375# vss 0.055237f
C313 _311_/a_254_473# net21 0.003733f
C314 FILLER_0_11_135/a_36_472# vss 0.006739f
C315 _072_ _228_/a_36_68# 0.005788f
C316 _437_/a_36_151# net14 0.014361f
C317 _448_/a_1204_472# vdd 0.002228f
C318 FILLER_0_10_78/a_1380_472# FILLER_0_10_94/a_36_472# 0.013277f
C319 output33/a_224_472# net33 0.151281f
C320 _176_ FILLER_0_15_72/a_572_375# 0.005529f
C321 net38 FILLER_0_20_2/a_484_472# 0.006727f
C322 FILLER_0_14_107/a_36_472# vss 0.003706f
C323 FILLER_0_14_107/a_484_472# vdd 0.030114f
C324 net52 _176_ 0.004215f
C325 net72 FILLER_0_12_50/a_36_472# 0.002007f
C326 valid vdd 0.148392f
C327 FILLER_0_22_177/a_36_472# vss 0.002984f
C328 FILLER_0_22_177/a_484_472# vdd 0.006974f
C329 mask\[2\] net23 0.431197f
C330 trim[4] output6/a_224_472# 0.004337f
C331 FILLER_0_12_136/a_572_375# FILLER_0_11_142/a_36_472# 0.001543f
C332 output44/a_224_472# _452_/a_1353_112# 0.001321f
C333 cal_itt\[3\] FILLER_0_5_198/a_124_375# 0.01268f
C334 net4 FILLER_0_12_220/a_932_472# 0.050731f
C335 _100_ _094_ 0.031066f
C336 _053_ _028_ 0.891578f
C337 _423_/a_36_151# FILLER_0_23_44/a_1468_375# 0.059049f
C338 _431_/a_448_472# fanout70/a_36_113# 0.001157f
C339 FILLER_0_7_104/a_484_472# _058_ 0.006506f
C340 net36 FILLER_0_15_212/a_484_472# 0.007742f
C341 FILLER_0_3_221/a_484_472# vss 0.005602f
C342 FILLER_0_3_221/a_932_472# vdd 0.005654f
C343 _064_ net47 0.110169f
C344 FILLER_0_15_116/a_124_375# net36 0.003055f
C345 _427_/a_448_472# _095_ 0.063616f
C346 _161_ vss 0.134214f
C347 net68 FILLER_0_5_54/a_572_375# 0.040374f
C348 _004_ _094_ 0.213913f
C349 net19 cal_itt\[0\] 0.111163f
C350 FILLER_0_9_28/a_2812_375# vdd 0.016637f
C351 net81 fanout79/a_36_160# 0.057526f
C352 mask\[0\] cal_count\[3\] 0.002612f
C353 _451_/a_36_151# vss 0.028073f
C354 _451_/a_448_472# vdd 0.04463f
C355 FILLER_0_5_54/a_932_472# _029_ 0.014976f
C356 FILLER_0_5_54/a_1468_375# trim_mask\[1\] 0.010901f
C357 FILLER_0_5_212/a_36_472# net37 0.007858f
C358 _104_ mask\[3\] 0.078406f
C359 _304_/a_224_472# _013_ 0.002769f
C360 _072_ calibrate 0.539702f
C361 FILLER_0_24_130/a_36_472# vdd 0.050082f
C362 _093_ _438_/a_1000_472# 0.001556f
C363 net50 net49 0.238748f
C364 _441_/a_36_151# _440_/a_448_472# 0.002538f
C365 _137_ FILLER_0_15_180/a_484_472# 0.046411f
C366 net52 _442_/a_2560_156# 0.008682f
C367 _294_/a_224_472# mask\[2\] 0.001715f
C368 FILLER_0_16_89/a_1020_375# _040_ 0.004252f
C369 fanout50/a_36_160# trim_val\[3\] 0.017252f
C370 net52 _036_ 0.013473f
C371 net50 net68 0.224698f
C372 fanout79/a_36_160# _060_ 0.005814f
C373 _429_/a_2248_156# _043_ 0.001001f
C374 FILLER_0_3_142/a_36_472# _081_ 0.001386f
C375 _257_/a_36_472# _068_ 0.002986f
C376 FILLER_0_18_177/a_3260_375# vss 0.055219f
C377 FILLER_0_18_177/a_36_472# vdd 0.110153f
C378 net20 net62 0.058892f
C379 output24/a_224_472# _025_ 0.010601f
C380 _115_ _322_/a_124_24# 0.019655f
C381 net9 vdd 0.190349f
C382 _076_ FILLER_0_8_156/a_484_472# 0.008487f
C383 net76 _076_ 0.003124f
C384 _013_ FILLER_0_18_53/a_484_472# 0.012916f
C385 _432_/a_796_472# _021_ 0.001666f
C386 net75 valid 0.002077f
C387 _053_ trim_mask\[0\] 0.007667f
C388 FILLER_0_23_88/a_36_472# vss 0.003481f
C389 _136_ _337_/a_49_472# 0.058704f
C390 _095_ _451_/a_2449_156# 0.001843f
C391 FILLER_0_16_57/a_124_375# vdd 0.008567f
C392 _440_/a_36_151# FILLER_0_6_47/a_1828_472# 0.001512f
C393 _417_/a_2560_156# _006_ 0.007804f
C394 FILLER_0_13_212/a_572_375# _070_ 0.003986f
C395 FILLER_0_5_128/a_36_472# _160_ 0.006214f
C396 FILLER_0_3_2/a_124_375# net66 0.027628f
C397 FILLER_0_7_72/a_484_472# net50 0.059395f
C398 net20 _199_/a_36_160# 0.05178f
C399 _287_/a_36_472# vdd 0.072871f
C400 FILLER_0_11_124/a_124_375# _135_ 0.004831f
C401 net25 _012_ 0.001747f
C402 trimb[0] net43 0.109028f
C403 net60 net30 0.001168f
C404 _171_ _172_ 0.104216f
C405 _089_ FILLER_0_5_198/a_124_375# 0.001517f
C406 FILLER_0_4_107/a_484_472# _031_ 0.002521f
C407 net65 _074_ 0.002666f
C408 _131_ FILLER_0_9_105/a_484_472# 0.004364f
C409 _002_ _087_ 0.00636f
C410 en fanout59/a_36_160# 0.242369f
C411 mask\[4\] mask\[3\] 1.118454f
C412 mask\[3\] net22 0.036607f
C413 _012_ net36 0.053654f
C414 net47 _153_ 0.755476f
C415 _412_/a_1204_472# net1 0.019647f
C416 FILLER_0_21_125/a_36_472# mask\[7\] 0.00344f
C417 _345_/a_36_160# _132_ 0.078243f
C418 net53 _427_/a_2248_156# 0.038716f
C419 _444_/a_2665_112# net67 0.03521f
C420 FILLER_0_5_72/a_1020_375# _164_ 0.018398f
C421 _015_ FILLER_0_8_247/a_1020_375# 0.006994f
C422 output17/a_224_472# net17 0.09023f
C423 FILLER_0_1_204/a_124_375# net11 0.01048f
C424 vss _201_/a_67_603# 0.012925f
C425 _077_ _134_ 0.043815f
C426 net81 _283_/a_36_472# 0.032292f
C427 output10/a_224_472# cal_itt\[0\] 0.008003f
C428 _091_ FILLER_0_16_154/a_1468_375# 0.003056f
C429 _114_ FILLER_0_13_142/a_1468_375# 0.001931f
C430 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_572_375# 0.001597f
C431 FILLER_0_8_127/a_124_375# vss 0.019066f
C432 _415_/a_2665_112# _416_/a_36_151# 0.001602f
C433 net57 _067_ 0.018966f
C434 _095_ FILLER_0_13_72/a_484_472# 0.027852f
C435 net75 net9 0.006945f
C436 _008_ _418_/a_2560_156# 0.006651f
C437 trim_mask\[2\] FILLER_0_2_93/a_572_375# 0.002818f
C438 _127_ vss 0.343764f
C439 _420_/a_36_151# net18 0.001426f
C440 FILLER_0_12_50/a_36_472# cal_count\[0\] 0.001857f
C441 _176_ _172_ 0.043154f
C442 _098_ _437_/a_36_151# 0.092841f
C443 _016_ net74 0.568682f
C444 _074_ net59 0.030221f
C445 FILLER_0_18_2/a_2276_472# net55 0.006033f
C446 net36 FILLER_0_15_235/a_484_472# 0.019725f
C447 FILLER_0_16_107/a_572_375# _040_ 0.001244f
C448 net65 FILLER_0_3_172/a_1020_375# 0.006035f
C449 output47/a_224_472# input3/a_36_113# 0.001371f
C450 _250_/a_36_68# _427_/a_2665_112# 0.002152f
C451 FILLER_0_7_104/a_572_375# _131_ 0.003031f
C452 net36 _438_/a_448_472# 0.034338f
C453 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1380_472# 0.013276f
C454 _274_/a_36_68# _070_ 0.032424f
C455 FILLER_0_14_91/a_36_472# en_co_clk 0.007733f
C456 FILLER_0_18_2/a_932_472# _452_/a_2225_156# 0.001256f
C457 FILLER_0_8_107/a_124_375# vss 0.031335f
C458 FILLER_0_12_136/a_1380_472# vss 0.031524f
C459 output35/a_224_472# net32 0.072991f
C460 ctln[4] _413_/a_2665_112# 0.001394f
C461 FILLER_0_16_57/a_124_375# net72 0.052543f
C462 _402_/a_1948_68# vdd 0.001429f
C463 _385_/a_244_472# net37 0.001593f
C464 FILLER_0_18_2/a_484_472# trimb[1] 0.009245f
C465 FILLER_0_21_142/a_572_375# _140_ 0.018708f
C466 _437_/a_2665_112# _436_/a_36_151# 0.001466f
C467 net70 _040_ 0.018254f
C468 _423_/a_2560_156# _012_ 0.004165f
C469 FILLER_0_15_142/a_36_472# net36 0.015456f
C470 net20 _429_/a_448_472# 0.002244f
C471 FILLER_0_16_89/a_124_375# _131_ 0.017319f
C472 net81 FILLER_0_14_235/a_124_375# 0.01391f
C473 _114_ FILLER_0_11_101/a_36_472# 0.00501f
C474 fanout68/a_36_113# _065_ 0.005586f
C475 FILLER_0_9_28/a_1020_375# net50 0.001512f
C476 net82 FILLER_0_3_221/a_124_375# 0.015932f
C477 net79 _005_ 1.006306f
C478 FILLER_0_8_138/a_36_472# _076_ 0.016628f
C479 net67 _160_ 0.003659f
C480 _410_/a_36_68# _453_/a_36_151# 0.002326f
C481 _071_ vss 0.126519f
C482 FILLER_0_19_111/a_484_472# vss 0.003811f
C483 net27 _100_ 0.006783f
C484 _023_ vss 0.114191f
C485 net79 FILLER_0_12_220/a_932_472# 0.005532f
C486 FILLER_0_19_187/a_36_472# vss 0.001951f
C487 FILLER_0_19_187/a_484_472# vdd 0.011023f
C488 ctlp[9] vdd 0.17413f
C489 net17 output6/a_224_472# 0.047757f
C490 FILLER_0_14_91/a_572_375# net14 0.005527f
C491 _446_/a_2665_112# _034_ 0.002484f
C492 _395_/a_36_488# state\[1\] 0.002702f
C493 _116_ _267_/a_36_472# 0.029316f
C494 FILLER_0_1_192/a_124_375# vdd 0.017212f
C495 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_36_472# 0.086635f
C496 net14 FILLER_0_10_94/a_484_472# 0.020589f
C497 _004_ net27 0.080285f
C498 _122_ _059_ 0.190023f
C499 FILLER_0_15_142/a_484_472# net36 0.012033f
C500 _174_ FILLER_0_15_59/a_572_375# 0.007123f
C501 FILLER_0_16_241/a_124_375# mask\[2\] 0.027201f
C502 ctlp[3] _422_/a_2560_156# 0.001006f
C503 net38 vss 0.633752f
C504 FILLER_0_16_73/a_484_472# vdd 0.003462f
C505 output11/a_224_472# vss 0.083244f
C506 _405_/a_67_603# cal_count\[2\] 0.021962f
C507 _030_ _156_ 0.153053f
C508 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1380_472# 0.013277f
C509 FILLER_0_21_28/a_2364_375# vdd -0.011393f
C510 FILLER_0_20_169/a_124_375# FILLER_0_19_171/a_36_472# 0.001543f
C511 FILLER_0_3_172/a_1380_472# vdd 0.043045f
C512 FILLER_0_21_125/a_484_472# _433_/a_36_151# 0.001723f
C513 _414_/a_36_151# vdd 0.166006f
C514 _053_ cal_itt\[3\] 0.471909f
C515 _077_ _229_/a_224_472# 0.001293f
C516 _442_/a_36_151# FILLER_0_2_127/a_36_472# 0.012873f
C517 ctlp[1] net79 0.002676f
C518 _131_ cal_count\[2\] 0.044147f
C519 FILLER_0_21_28/a_36_472# net17 0.00347f
C520 _427_/a_448_472# net74 0.051943f
C521 net4 FILLER_0_3_221/a_484_472# 0.043027f
C522 _438_/a_2665_112# net14 0.026903f
C523 output27/a_224_472# FILLER_0_8_263/a_124_375# 0.011584f
C524 state\[1\] _228_/a_36_68# 0.024977f
C525 net20 _294_/a_224_472# 0.008053f
C526 _093_ FILLER_0_18_107/a_3172_472# 0.008787f
C527 _076_ _083_ 0.006023f
C528 _359_/a_1492_488# _133_ 0.003815f
C529 _068_ _078_ 0.002973f
C530 net16 _173_ 0.029412f
C531 FILLER_0_22_177/a_1020_375# net33 0.013731f
C532 _091_ FILLER_0_18_209/a_484_472# 0.001212f
C533 _053_ _081_ 0.698311f
C534 _414_/a_2560_156# cal_itt\[3\] 0.007141f
C535 _132_ _040_ 0.023821f
C536 net57 _121_ 0.004182f
C537 _414_/a_36_151# FILLER_0_6_177/a_572_375# 0.073306f
C538 output15/a_224_472# net52 0.007862f
C539 net15 fanout50/a_36_160# 0.029852f
C540 _091_ FILLER_0_12_220/a_1020_375# 0.001598f
C541 FILLER_0_10_214/a_36_472# vss 0.008006f
C542 _005_ _416_/a_2665_112# 0.014205f
C543 _442_/a_1308_423# _031_ 0.003679f
C544 _053_ FILLER_0_7_104/a_932_472# 0.002529f
C545 _131_ FILLER_0_11_124/a_36_472# 0.015445f
C546 _412_/a_1000_472# net1 0.027748f
C547 _155_ FILLER_0_6_90/a_572_375# 0.001562f
C548 _414_/a_2560_156# _081_ 0.008322f
C549 result[0] FILLER_0_9_290/a_36_472# 0.020103f
C550 result[7] _108_ 0.063624f
C551 FILLER_0_5_72/a_124_375# net47 0.006974f
C552 _350_/a_49_472# _147_ 0.016114f
C553 _084_ vdd 0.134578f
C554 _413_/a_3041_156# net59 0.001022f
C555 net31 _277_/a_36_160# 0.053915f
C556 FILLER_0_8_127/a_36_472# _125_ 0.003088f
C557 FILLER_0_10_256/a_124_375# vss 0.006036f
C558 FILLER_0_10_256/a_36_472# vdd 0.025204f
C559 net22 _435_/a_2665_112# 0.004214f
C560 net58 net76 0.700034f
C561 FILLER_0_7_162/a_124_375# net47 0.030995f
C562 mask\[0\] _429_/a_2665_112# 0.016053f
C563 FILLER_0_7_162/a_36_472# vss 0.006392f
C564 _086_ _053_ 0.091538f
C565 _003_ _414_/a_796_472# 0.006511f
C566 net63 FILLER_0_22_177/a_1468_375# 0.005028f
C567 net24 FILLER_0_22_86/a_1020_375# 0.022658f
C568 _140_ _207_/a_67_603# 0.014923f
C569 net68 _054_ 0.08092f
C570 FILLER_0_12_136/a_484_472# net23 0.002172f
C571 net16 _444_/a_36_151# 0.010514f
C572 _325_/a_224_472# _118_ 0.004845f
C573 FILLER_0_20_177/a_1380_472# _098_ 0.00679f
C574 FILLER_0_4_107/a_124_375# vdd 0.036972f
C575 FILLER_0_5_212/a_36_472# _122_ 0.002272f
C576 _077_ _439_/a_1308_423# 0.022235f
C577 _103_ _418_/a_2248_156# 0.012186f
C578 net62 vss 1.17087f
C579 _119_ _053_ 0.038651f
C580 _144_ _437_/a_2665_112# 0.001186f
C581 _046_ mask\[2\] 0.003147f
C582 _430_/a_1308_423# mask\[2\] 0.020226f
C583 FILLER_0_16_241/a_36_472# _282_/a_36_160# 0.006647f
C584 _376_/a_36_160# FILLER_0_6_90/a_36_472# 0.195478f
C585 _085_ FILLER_0_13_142/a_1468_375# 0.001153f
C586 FILLER_0_9_105/a_484_472# FILLER_0_10_107/a_124_375# 0.001543f
C587 net47 _166_ 0.034342f
C588 net52 _449_/a_448_472# 0.001042f
C589 _010_ net77 0.009534f
C590 _297_/a_36_472# _108_ 0.011437f
C591 _093_ FILLER_0_17_72/a_1380_472# 0.008517f
C592 FILLER_0_9_28/a_1916_375# _042_ 0.002352f
C593 _413_/a_2665_112# net21 0.002828f
C594 vss FILLER_0_5_148/a_572_375# 0.042687f
C595 vdd FILLER_0_5_148/a_36_472# 0.001227f
C596 _233_/a_36_160# vss 0.01649f
C597 _079_ FILLER_0_6_231/a_572_375# 0.002768f
C598 output33/a_224_472# net18 0.110644f
C599 _162_ _058_ 0.015239f
C600 FILLER_0_17_72/a_572_375# FILLER_0_15_72/a_484_472# 0.001512f
C601 _199_/a_36_160# vss 0.004608f
C602 net75 _084_ 0.045583f
C603 net74 FILLER_0_13_72/a_484_472# 0.007142f
C604 _126_ _390_/a_36_68# 0.044675f
C605 net50 FILLER_0_8_37/a_36_472# 0.059367f
C606 _246_/a_36_68# vss 0.024639f
C607 net75 FILLER_0_10_256/a_36_472# 0.010024f
C608 _177_ _131_ 0.058938f
C609 _077_ FILLER_0_10_78/a_932_472# 0.002503f
C610 _415_/a_2665_112# result[1] 0.010555f
C611 ctln[5] net59 0.030363f
C612 _432_/a_2665_112# mask\[3\] 0.011428f
C613 net82 _159_ 0.001393f
C614 _077_ _311_/a_66_473# 0.002605f
C615 _217_/a_36_160# FILLER_0_19_28/a_484_472# 0.006053f
C616 _408_/a_728_93# _043_ 0.029183f
C617 net23 _386_/a_124_24# 0.010805f
C618 _176_ FILLER_0_11_101/a_572_375# 0.00389f
C619 output38/a_224_472# _064_ 0.017666f
C620 _428_/a_796_472# _017_ 0.025239f
C621 _116_ _113_ 0.179616f
C622 FILLER_0_21_28/a_2364_375# _424_/a_36_151# 0.059049f
C623 FILLER_0_19_155/a_572_375# vdd 0.01384f
C624 FILLER_0_19_155/a_124_375# vss 0.00336f
C625 net63 mask\[6\] 0.146994f
C626 FILLER_0_16_57/a_1380_472# cal_count\[1\] 0.001568f
C627 _096_ _055_ 0.047639f
C628 _098_ _438_/a_2665_112# 0.004321f
C629 FILLER_0_5_54/a_572_375# net47 0.009717f
C630 net14 FILLER_0_4_91/a_124_375# 0.009573f
C631 FILLER_0_2_111/a_932_472# _158_ 0.00264f
C632 output38/a_224_472# output41/a_224_472# 0.00607f
C633 _432_/a_448_472# vdd 0.035246f
C634 output29/a_224_472# _005_ 0.021351f
C635 net29 _101_ 0.007132f
C636 _114_ state\[2\] 0.528838f
C637 FILLER_0_0_198/a_124_375# vdd 0.04491f
C638 net82 FILLER_0_3_172/a_2364_375# 0.010439f
C639 net55 vss 0.947665f
C640 net73 FILLER_0_17_142/a_124_375# 0.003021f
C641 _452_/a_2225_156# vdd 0.005612f
C642 _452_/a_3129_107# vss 0.00145f
C643 _412_/a_796_472# net2 0.00566f
C644 FILLER_0_4_123/a_36_472# net74 0.001578f
C645 _165_ trim_mask\[1\] 0.002231f
C646 _369_/a_36_68# vss 0.002343f
C647 output28/a_224_472# vdd 0.044767f
C648 net17 _452_/a_1697_156# 0.001184f
C649 _039_ output6/a_224_472# 0.012051f
C650 net20 FILLER_0_16_241/a_124_375# 0.002327f
C651 net50 net47 0.040157f
C652 _394_/a_56_524# _095_ 0.10007f
C653 net18 _419_/a_448_472# 0.037373f
C654 _137_ FILLER_0_16_154/a_1020_375# 0.010692f
C655 _081_ FILLER_0_5_164/a_36_472# 0.001603f
C656 FILLER_0_12_2/a_124_375# clkc 0.003601f
C657 net71 _436_/a_36_151# 0.03535f
C658 _028_ FILLER_0_7_104/a_932_472# 0.003084f
C659 net76 FILLER_0_5_172/a_124_375# 0.001526f
C660 FILLER_0_4_185/a_36_472# _087_ 0.008805f
C661 _127_ _332_/a_36_472# 0.00288f
C662 trim[0] trim[1] 0.001567f
C663 output21/a_224_472# mask\[6\] 0.013037f
C664 _072_ _069_ 0.265737f
C665 net81 fanout82/a_36_113# 0.061162f
C666 net81 _425_/a_448_472# 0.056225f
C667 FILLER_0_2_171/a_36_472# FILLER_0_2_165/a_36_472# 0.003468f
C668 _340_/a_36_160# _098_ 0.019601f
C669 output30/a_224_472# net30 0.043557f
C670 output27/a_224_472# FILLER_0_9_282/a_484_472# 0.001711f
C671 net77 vdd 0.526632f
C672 FILLER_0_18_107/a_1020_375# FILLER_0_17_104/a_1380_472# 0.001597f
C673 _429_/a_448_472# vss 0.035246f
C674 net64 FILLER_0_14_235/a_124_375# 0.046554f
C675 _176_ _318_/a_224_472# 0.003019f
C676 _116_ _118_ 0.054068f
C677 _136_ _171_ 0.008792f
C678 _423_/a_36_151# vdd 0.088377f
C679 net52 _032_ 0.009879f
C680 _415_/a_448_472# net19 0.03569f
C681 FILLER_0_16_107/a_124_375# _093_ 0.003941f
C682 _088_ _073_ 0.001254f
C683 FILLER_0_14_50/a_36_472# _180_ 0.153222f
C684 FILLER_0_9_28/a_1020_375# _054_ 0.002273f
C685 mask\[8\] _050_ 0.001479f
C686 _093_ FILLER_0_16_115/a_124_375# 0.003988f
C687 _395_/a_36_488# vdd 0.066813f
C688 state\[1\] FILLER_0_12_196/a_36_472# 0.030132f
C689 ctlp[6] ctlp[7] 0.002504f
C690 _443_/a_36_151# trim_mask\[4\] 0.002625f
C691 calibrate _385_/a_36_68# 0.001996f
C692 mask\[3\] _008_ 0.799138f
C693 trim_mask\[3\] _156_ 0.002638f
C694 _132_ _428_/a_1204_472# 0.025555f
C695 trimb[3] output17/a_224_472# 0.047604f
C696 _427_/a_2248_156# _071_ 0.001131f
C697 FILLER_0_17_72/a_36_472# net36 0.001121f
C698 _086_ _028_ 0.011526f
C699 FILLER_0_10_214/a_124_375# _055_ 0.001419f
C700 _042_ net51 0.026776f
C701 _441_/a_36_151# FILLER_0_3_78/a_36_472# 0.001723f
C702 ctlp[1] FILLER_0_21_286/a_36_472# 0.014043f
C703 _423_/a_36_151# FILLER_0_23_60/a_36_472# 0.001723f
C704 mask\[1\] FILLER_0_15_180/a_484_472# 0.003594f
C705 _182_ cal_count\[1\] 0.166348f
C706 _442_/a_1308_423# FILLER_0_2_111/a_1468_375# 0.001048f
C707 FILLER_0_22_128/a_1916_375# vss 0.018094f
C708 FILLER_0_22_128/a_2364_375# vdd 0.015888f
C709 net23 vss 1.922425f
C710 _075_ _414_/a_2665_112# 0.050503f
C711 FILLER_0_20_107/a_124_375# vdd 0.04384f
C712 _060_ _223_/a_36_160# 0.002922f
C713 _424_/a_1000_472# vdd 0.002952f
C714 FILLER_0_23_290/a_36_472# vdd 0.089567f
C715 FILLER_0_23_290/a_124_375# vss 0.033011f
C716 _070_ _171_ 0.084342f
C717 fanout51/a_36_113# cal_count\[3\] 0.054567f
C718 _441_/a_2665_112# vss 0.005169f
C719 _064_ vdd 0.874293f
C720 mask\[5\] FILLER_0_20_177/a_1468_375# 0.013222f
C721 _059_ _160_ 0.037235f
C722 net75 output28/a_224_472# 0.00151f
C723 net55 _452_/a_836_156# 0.010887f
C724 _228_/a_36_68# vdd 0.036391f
C725 net69 _164_ 0.040362f
C726 _053_ FILLER_0_6_47/a_1468_375# 0.008103f
C727 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_484_472# 0.001723f
C728 _061_ _247_/a_36_160# 0.009993f
C729 mask\[3\] FILLER_0_18_177/a_932_472# 0.005654f
C730 _447_/a_1204_472# vdd 0.001085f
C731 _117_ _113_ 0.09166f
C732 fanout74/a_36_113# vss 0.048756f
C733 _320_/a_36_472# _090_ 0.001941f
C734 _187_ _186_ 0.032149f
C735 _176_ _136_ 0.114837f
C736 vdd output41/a_224_472# 0.003282f
C737 net50 FILLER_0_9_60/a_124_375# 0.001715f
C738 net63 FILLER_0_19_187/a_572_375# 0.049706f
C739 _035_ net49 0.018245f
C740 FILLER_0_20_193/a_572_375# _434_/a_2665_112# 0.002362f
C741 _439_/a_2248_156# vss 0.003954f
C742 _439_/a_2665_112# vdd 0.015979f
C743 _104_ _421_/a_448_472# 0.001106f
C744 _294_/a_224_472# vss 0.001022f
C745 _136_ _335_/a_49_472# 0.039074f
C746 _345_/a_36_160# vdd 0.100094f
C747 fanout49/a_36_160# _030_ 0.017759f
C748 calibrate FILLER_0_7_233/a_124_375# 0.011958f
C749 fanout64/a_36_160# _425_/a_2665_112# 0.005704f
C750 output21/a_224_472# _009_ 0.004164f
C751 output17/a_224_472# ctlp[0] 0.018696f
C752 mask\[9\] FILLER_0_18_76/a_36_472# 0.002584f
C753 ctln[2] net18 0.106494f
C754 trim_val\[4\] FILLER_0_3_172/a_36_472# 0.006208f
C755 net76 FILLER_0_3_172/a_2276_472# 0.002531f
C756 trim_val\[4\] _386_/a_124_24# 0.001172f
C757 _426_/a_36_151# FILLER_0_8_247/a_1380_472# 0.001723f
C758 net72 _423_/a_36_151# 0.024965f
C759 output34/a_224_472# net19 0.001308f
C760 net20 _046_ 0.194455f
C761 _116_ _068_ 0.011673f
C762 _176_ _070_ 0.467961f
C763 _320_/a_36_472# net22 0.005964f
C764 net56 FILLER_0_18_139/a_932_472# 0.011079f
C765 _070_ FILLER_0_5_164/a_572_375# 0.001083f
C766 calibrate vdd 0.857987f
C767 net32 _094_ 0.027571f
C768 result[6] _421_/a_448_472# 0.038671f
C769 FILLER_0_9_28/a_2724_472# _453_/a_36_151# 0.013806f
C770 FILLER_0_15_290/a_36_472# net18 0.002452f
C771 _025_ vss 0.016676f
C772 net56 FILLER_0_16_154/a_1020_375# 0.002321f
C773 fanout53/a_36_160# FILLER_0_16_154/a_484_472# 0.014774f
C774 net52 FILLER_0_2_93/a_124_375# 0.007787f
C775 FILLER_0_5_128/a_484_472# net74 0.025425f
C776 ctlp[1] ctlp[2] 0.002331f
C777 FILLER_0_17_72/a_2724_472# net14 0.007133f
C778 mask\[5\] FILLER_0_19_171/a_484_472# 0.007647f
C779 _118_ _117_ 0.032074f
C780 FILLER_0_15_10/a_36_472# vss 0.002605f
C781 cal_count\[3\] net51 0.042416f
C782 _105_ output35/a_224_472# 0.013092f
C783 output42/a_224_472# net40 0.003278f
C784 net55 _424_/a_448_472# 0.005273f
C785 _311_/a_1920_473# vdd 0.007492f
C786 _143_ FILLER_0_17_161/a_36_472# 0.00363f
C787 _430_/a_36_151# FILLER_0_17_200/a_36_472# 0.001723f
C788 FILLER_0_2_101/a_124_375# _367_/a_36_68# 0.001176f
C789 result[8] output19/a_224_472# 0.001465f
C790 net33 vss 0.674927f
C791 _431_/a_1308_423# vss 0.003472f
C792 cal_itt\[2\] _088_ 0.010847f
C793 _431_/a_448_472# _093_ 0.002095f
C794 _153_ vdd 0.672318f
C795 net34 _109_ 0.001298f
C796 _154_ _365_/a_36_68# 0.02267f
C797 _144_ net71 0.039862f
C798 _412_/a_1308_423# net65 0.024499f
C799 _232_/a_67_603# FILLER_0_5_54/a_36_472# 0.025312f
C800 _079_ _253_/a_36_68# 0.002433f
C801 _112_ FILLER_0_8_247/a_932_472# 0.001185f
C802 net4 _246_/a_36_68# 0.003771f
C803 net17 FILLER_0_20_15/a_124_375# 0.005919f
C804 net18 FILLER_0_17_282/a_36_472# 0.036965f
C805 _077_ FILLER_0_9_72/a_932_472# 0.006408f
C806 _321_/a_3662_472# net74 0.00253f
C807 _056_ vss 0.193804f
C808 _427_/a_2560_156# vss 0.003576f
C809 FILLER_0_12_124/a_36_472# _017_ 0.004641f
C810 _103_ _102_ 0.392644f
C811 _136_ FILLER_0_17_133/a_124_375# 0.001315f
C812 _424_/a_36_151# _423_/a_36_151# 0.006746f
C813 trim_val\[1\] _160_ 0.024279f
C814 output8/a_224_472# _411_/a_36_151# 0.12978f
C815 _053_ _161_ 0.001047f
C816 FILLER_0_14_81/a_36_472# _394_/a_728_93# 0.005826f
C817 FILLER_0_11_78/a_572_375# _171_ 0.001028f
C818 _287_/a_36_472# _099_ 0.030964f
C819 _093_ FILLER_0_18_177/a_2724_472# 0.003036f
C820 FILLER_0_14_263/a_36_472# output30/a_224_472# 0.002002f
C821 net75 calibrate 0.101912f
C822 _322_/a_1152_472# _129_ 0.002978f
C823 net41 _095_ 0.641184f
C824 net51 net40 0.060626f
C825 _002_ FILLER_0_3_172/a_2724_472# 0.006713f
C826 FILLER_0_17_56/a_124_375# vdd 0.008529f
C827 trim_val\[4\] vss 0.192567f
C828 net5 net8 0.001288f
C829 net38 _444_/a_796_472# 0.002641f
C830 _392_/a_36_68# vss 0.002019f
C831 _091_ net80 0.23053f
C832 FILLER_0_8_37/a_36_472# _054_ 0.015053f
C833 net16 _041_ 0.029736f
C834 FILLER_0_14_99/a_36_472# _095_ 0.011772f
C835 _214_/a_36_160# FILLER_0_23_88/a_124_375# 0.005398f
C836 _411_/a_1308_423# vss 0.0013f
C837 _412_/a_1308_423# net59 0.00291f
C838 _165_ _164_ 0.351097f
C839 output38/a_224_472# _446_/a_448_472# 0.007649f
C840 _258_/a_36_160# net59 0.003167f
C841 _449_/a_2560_156# _067_ 0.007511f
C842 cal_itt\[3\] _081_ 0.03503f
C843 output45/a_224_472# vdd -0.026726f
C844 net62 FILLER_0_13_212/a_1020_375# 0.001597f
C845 FILLER_0_13_212/a_36_472# vss 0.005259f
C846 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_36_472# 0.026657f
C847 net58 FILLER_0_8_263/a_124_375# 0.001876f
C848 _394_/a_56_524# net74 0.005616f
C849 _012_ FILLER_0_23_44/a_1020_375# 0.002827f
C850 _436_/a_1204_472# vdd 0.003143f
C851 _080_ net37 0.005467f
C852 net42 output6/a_224_472# 0.009273f
C853 _068_ _117_ 0.011659f
C854 FILLER_0_9_28/a_1828_472# _054_ 0.003145f
C855 trimb[4] FILLER_0_15_2/a_36_472# 0.006046f
C856 mask\[2\] FILLER_0_15_235/a_572_375# 0.003879f
C857 _040_ vdd 0.065702f
C858 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3172_472# 0.013277f
C859 _000_ net8 0.021422f
C860 mask\[5\] _434_/a_2665_112# 0.003849f
C861 net60 _418_/a_2665_112# 0.042307f
C862 _176_ FILLER_0_11_78/a_572_375# 0.013887f
C863 _125_ vdd 0.218505f
C864 net54 mask\[9\] 0.094381f
C865 net20 net18 0.025322f
C866 _030_ _440_/a_36_151# 0.001187f
C867 net52 FILLER_0_6_79/a_36_472# 0.012286f
C868 _394_/a_56_524# cal_count\[1\] 0.022487f
C869 mask\[8\] _423_/a_2665_112# 0.004281f
C870 net35 _423_/a_2248_156# 0.003899f
C871 _103_ _198_/a_67_603# 0.005362f
C872 ctln[6] ctln[7] 0.00499f
C873 output10/a_224_472# net10 0.012455f
C874 ctlp[1] _420_/a_1308_423# 0.001418f
C875 _440_/a_1000_472# _029_ 0.004334f
C876 mask\[7\] FILLER_0_22_128/a_1916_375# 0.007718f
C877 mask\[7\] net23 0.225177f
C878 FILLER_0_16_241/a_124_375# vss 0.04897f
C879 FILLER_0_16_241/a_36_472# vdd 0.012388f
C880 net47 _054_ 0.171966f
C881 _422_/a_2665_112# _107_ 0.005055f
C882 output10/a_224_472# FILLER_0_0_232/a_124_375# 0.00363f
C883 _168_ _160_ 0.03261f
C884 FILLER_0_5_212/a_124_375# FILLER_0_3_212/a_36_472# 0.001512f
C885 _086_ cal_itt\[3\] 0.046874f
C886 net54 FILLER_0_22_86/a_1380_472# 0.059367f
C887 _254_/a_448_472# _074_ 0.002163f
C888 _077_ _114_ 0.047702f
C889 output6/a_224_472# clkc 0.017846f
C890 _069_ state\[1\] 0.003884f
C891 net35 FILLER_0_22_128/a_1380_472# 0.016004f
C892 trim_mask\[2\] _381_/a_36_472# 0.034251f
C893 output39/a_224_472# net66 0.009679f
C894 _092_ _069_ 0.040267f
C895 net36 _451_/a_836_156# 0.007104f
C896 FILLER_0_2_111/a_124_375# trim_mask\[3\] 0.004993f
C897 net72 FILLER_0_17_56/a_124_375# 0.018942f
C898 trim_val\[4\] FILLER_0_2_165/a_124_375# 0.009193f
C899 net16 net49 0.055931f
C900 _089_ cal_itt\[3\] 0.049851f
C901 vdd FILLER_0_12_196/a_36_472# 0.019648f
C902 vss FILLER_0_12_196/a_124_375# 0.042104f
C903 _086_ _081_ 0.033115f
C904 _367_/a_36_68# net14 0.055776f
C905 _363_/a_36_68# vss 0.043707f
C906 _119_ cal_itt\[3\] 0.010152f
C907 net16 net68 0.275467f
C908 net64 FILLER_0_9_282/a_572_375# 0.002322f
C909 _136_ FILLER_0_16_154/a_932_472# 0.008185f
C910 trim_mask\[1\] FILLER_0_6_47/a_36_472# 0.004319f
C911 _174_ vdd 0.18623f
C912 output39/a_224_472# _445_/a_1308_423# 0.010408f
C913 FILLER_0_1_266/a_484_472# net18 0.010423f
C914 FILLER_0_1_266/a_572_375# net8 0.016292f
C915 _089_ _081_ 0.002206f
C916 net27 mask\[0\] 0.067038f
C917 _207_/a_67_603# FILLER_0_22_128/a_3260_375# 0.00744f
C918 fanout68/a_36_113# net66 0.042828f
C919 _086_ FILLER_0_7_104/a_932_472# 0.001786f
C920 net20 FILLER_0_15_212/a_1468_375# 0.006824f
C921 net64 _223_/a_36_160# 0.007842f
C922 FILLER_0_21_142/a_572_375# _098_ 0.006558f
C923 _052_ FILLER_0_18_37/a_572_375# 0.00706f
C924 _444_/a_2248_156# vdd 0.041347f
C925 _115_ cal_count\[3\] 0.004426f
C926 FILLER_0_13_80/a_36_472# _451_/a_3129_107# 0.001115f
C927 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1380_472# 0.013276f
C928 net40 net6 0.00772f
C929 FILLER_0_8_138/a_124_375# _129_ 0.006506f
C930 FILLER_0_12_220/a_572_375# _060_ 0.00145f
C931 _446_/a_448_472# vdd 0.006805f
C932 ctlp[1] _421_/a_1000_472# 0.007039f
C933 _427_/a_2248_156# net23 0.033973f
C934 net53 FILLER_0_13_142/a_572_375# 0.001597f
C935 FILLER_0_5_72/a_124_375# vdd -0.005497f
C936 output14/a_224_472# _442_/a_36_151# 0.172111f
C937 net62 net79 1.615103f
C938 _446_/a_1000_472# net17 0.031119f
C939 net63 _429_/a_36_151# 0.0144f
C940 FILLER_0_4_144/a_36_472# _370_/a_848_380# 0.15783f
C941 _316_/a_124_24# _123_ 0.009391f
C942 _053_ FILLER_0_8_107/a_124_375# 0.002386f
C943 _394_/a_1336_472# FILLER_0_13_72/a_36_472# 0.008136f
C944 _394_/a_728_93# FILLER_0_13_72/a_572_375# 0.001064f
C945 _009_ _296_/a_224_472# 0.001278f
C946 net20 fanout75/a_36_113# 0.001027f
C947 _063_ _444_/a_36_151# 0.030369f
C948 FILLER_0_4_91/a_572_375# _160_ 0.007391f
C949 _431_/a_2560_156# _136_ 0.013111f
C950 FILLER_0_3_204/a_36_472# FILLER_0_4_197/a_932_472# 0.026657f
C951 result[6] _419_/a_36_151# 0.001968f
C952 _148_ _025_ 0.007252f
C953 net35 FILLER_0_22_107/a_572_375# 0.010438f
C954 mask\[8\] FILLER_0_22_107/a_36_472# 0.017159f
C955 _089_ _270_/a_36_472# 0.00437f
C956 _055_ _311_/a_1212_473# 0.004259f
C957 _211_/a_36_160# _050_ 0.010927f
C958 FILLER_0_7_162/a_124_375# vdd 0.011809f
C959 _072_ _090_ 0.091468f
C960 _169_ _163_ 0.013133f
C961 FILLER_0_21_142/a_572_375# _433_/a_2248_156# 0.006739f
C962 _417_/a_1000_472# net30 0.004556f
C963 FILLER_0_16_89/a_36_472# _136_ 0.00722f
C964 FILLER_0_17_104/a_572_375# _451_/a_36_151# 0.001619f
C965 FILLER_0_17_104/a_124_375# _451_/a_448_472# 0.001718f
C966 net65 _163_ 0.013462f
C967 _372_/a_2590_472# _062_ 0.0012f
C968 FILLER_0_18_177/a_124_375# FILLER_0_20_177/a_36_472# 0.0027f
C969 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_572_375# 0.086635f
C970 FILLER_0_12_136/a_1020_375# _126_ 0.012732f
C971 mask\[7\] net33 0.02491f
C972 _415_/a_2248_156# _416_/a_36_151# 0.001495f
C973 _098_ FILLER_0_15_228/a_36_472# 0.022074f
C974 _119_ _086_ 0.419383f
C975 net54 _352_/a_49_472# 0.003941f
C976 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_572_375# 0.007947f
C977 _176_ _451_/a_448_472# 0.007191f
C978 _451_/a_1697_156# net14 0.001298f
C979 input1/a_36_113# en 0.036849f
C980 net70 FILLER_0_11_101/a_484_472# 0.001474f
C981 net82 net76 0.061682f
C982 net15 _449_/a_36_151# 0.020788f
C983 _292_/a_36_160# net32 0.011466f
C984 _094_ _418_/a_1204_472# 0.009231f
C985 net54 net35 0.114666f
C986 FILLER_0_18_107/a_1020_375# mask\[9\] 0.005758f
C987 net72 _174_ 0.199504f
C988 _046_ vss 0.088886f
C989 _430_/a_1308_423# vss 0.003054f
C990 _072_ net22 0.147672f
C991 mask\[0\] _043_ 0.929722f
C992 _307_/a_234_472# _126_ 0.00204f
C993 net26 _052_ 0.100927f
C994 trim[4] _236_/a_36_160# 0.004514f
C995 _415_/a_2665_112# net27 0.030051f
C996 vdd _166_ 0.108744f
C997 _315_/a_716_497# net23 0.004725f
C998 FILLER_0_15_282/a_484_472# result[3] 0.026996f
C999 _056_ net4 0.002408f
C1000 net62 _416_/a_2665_112# 0.037195f
C1001 _420_/a_36_151# FILLER_0_23_282/a_36_472# 0.001723f
C1002 output12/a_224_472# _413_/a_36_151# 0.006251f
C1003 net17 _034_ 0.020793f
C1004 FILLER_0_12_20/a_124_375# net6 0.003726f
C1005 _141_ FILLER_0_19_155/a_124_375# 0.029562f
C1006 _431_/a_36_151# net70 0.031018f
C1007 _410_/a_244_472# _042_ 0.003902f
C1008 _149_ FILLER_0_20_87/a_36_472# 0.001938f
C1009 _061_ _311_/a_66_473# 0.030169f
C1010 _073_ _260_/a_36_68# 0.079772f
C1011 net7 output7/a_224_472# 0.01565f
C1012 net50 FILLER_0_4_91/a_36_472# 0.058499f
C1013 _413_/a_1000_472# net21 0.041643f
C1014 FILLER_0_9_28/a_36_472# output42/a_224_472# 0.010684f
C1015 FILLER_0_9_28/a_484_472# vdd 0.010868f
C1016 _140_ FILLER_0_22_128/a_2724_472# 0.004196f
C1017 _170_ _241_/a_224_472# 0.001199f
C1018 FILLER_0_15_290/a_36_472# _417_/a_36_151# 0.027236f
C1019 net58 FILLER_0_9_282/a_484_472# 0.091905f
C1020 net15 FILLER_0_15_59/a_36_472# 0.00464f
C1021 FILLER_0_16_57/a_124_375# _176_ 0.015872f
C1022 _095_ cal_count\[2\] 0.270066f
C1023 _345_/a_36_160# _433_/a_36_151# 0.015565f
C1024 FILLER_0_18_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001684f
C1025 FILLER_0_0_232/a_36_472# vss 0.007185f
C1026 FILLER_0_9_270/a_572_375# vdd 0.02345f
C1027 _015_ vdd 0.27747f
C1028 _290_/a_224_472# net18 0.00868f
C1029 FILLER_0_16_255/a_36_472# _094_ 0.005892f
C1030 FILLER_0_5_109/a_124_375# FILLER_0_4_107/a_484_472# 0.001684f
C1031 FILLER_0_12_20/a_572_375# net40 0.007477f
C1032 FILLER_0_20_193/a_572_375# net35 0.002196f
C1033 FILLER_0_9_28/a_1020_375# net16 0.012909f
C1034 FILLER_0_21_125/a_36_472# _022_ 0.002295f
C1035 FILLER_0_17_200/a_484_472# mask\[3\] 0.014805f
C1036 _025_ _436_/a_1308_423# 0.006243f
C1037 net70 FILLER_0_18_107/a_1380_472# 0.00116f
C1038 FILLER_0_3_142/a_36_472# net23 0.043034f
C1039 _058_ _055_ 0.070216f
C1040 _428_/a_1204_472# vdd 0.001231f
C1041 result[7] _421_/a_448_472# 0.018021f
C1042 _031_ FILLER_0_2_127/a_124_375# 0.013811f
C1043 _032_ _152_ 0.001206f
C1044 FILLER_0_5_54/a_572_375# vdd 0.004086f
C1045 _413_/a_36_151# FILLER_0_3_204/a_36_472# 0.001723f
C1046 FILLER_0_12_220/a_484_472# _070_ 0.004091f
C1047 _432_/a_1000_472# net80 0.033803f
C1048 cal_count\[3\] _389_/a_428_148# 0.001072f
C1049 _077_ _187_ 0.058967f
C1050 result[8] FILLER_0_24_274/a_1468_375# 0.00726f
C1051 fanout51/a_36_113# _120_ 0.014349f
C1052 output43/a_224_472# vdd -0.032713f
C1053 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_572_375# 0.086635f
C1054 cal_itt\[1\] net18 0.026586f
C1055 FILLER_0_17_282/a_36_472# _417_/a_36_151# 0.001723f
C1056 FILLER_0_15_72/a_484_472# vdd 0.002283f
C1057 FILLER_0_15_72/a_36_472# vss 0.038986f
C1058 FILLER_0_9_28/a_36_472# net51 0.002082f
C1059 fanout74/a_36_113# FILLER_0_3_142/a_36_472# 0.016516f
C1060 _412_/a_1308_423# output9/a_224_472# 0.001352f
C1061 net50 vdd 0.661261f
C1062 FILLER_0_17_72/a_2724_472# _131_ 0.004095f
C1063 _053_ FILLER_0_7_162/a_36_472# 0.004888f
C1064 _074_ _375_/a_960_497# 0.004175f
C1065 _035_ net47 0.101683f
C1066 FILLER_0_22_177/a_36_472# _434_/a_448_472# 0.012285f
C1067 _440_/a_448_472# _164_ 0.0036f
C1068 _196_/a_36_160# FILLER_0_14_263/a_36_472# 0.004828f
C1069 _443_/a_1000_472# vss 0.031435f
C1070 _305_/a_36_159# _316_/a_124_24# 0.003478f
C1071 _431_/a_36_151# _132_ 0.051016f
C1072 output36/a_224_472# net29 0.077505f
C1073 _033_ FILLER_0_6_37/a_36_472# 0.017695f
C1074 FILLER_0_19_28/a_124_375# net40 0.047489f
C1075 mask\[3\] FILLER_0_17_161/a_124_375# 0.032905f
C1076 _155_ net47 0.009532f
C1077 _058_ _313_/a_67_603# 0.010094f
C1078 _141_ net23 0.782974f
C1079 output28/a_224_472# _416_/a_2248_156# 0.023576f
C1080 result[1] _416_/a_448_472# 0.008784f
C1081 FILLER_0_4_197/a_36_472# _079_ 0.002448f
C1082 sample net18 0.103617f
C1083 _072_ _076_ 0.068172f
C1084 FILLER_0_5_72/a_1020_375# _440_/a_2248_156# 0.001068f
C1085 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_124_375# 0.012001f
C1086 net75 _015_ 0.025217f
C1087 net18 vss 1.110302f
C1088 _164_ FILLER_0_6_47/a_36_472# 0.047981f
C1089 _077_ _251_/a_906_472# 0.001076f
C1090 trimb[3] FILLER_0_20_15/a_124_375# 0.001391f
C1091 _067_ FILLER_0_13_72/a_572_375# 0.001874f
C1092 FILLER_0_17_64/a_36_472# net36 0.00195f
C1093 _091_ _106_ 0.001188f
C1094 _174_ cal_count\[0\] 0.009645f
C1095 _132_ FILLER_0_18_107/a_1380_472# 0.034976f
C1096 net16 FILLER_0_18_37/a_36_472# 0.001132f
C1097 _144_ FILLER_0_22_128/a_2812_375# 0.001601f
C1098 _069_ vdd 0.985405f
C1099 net46 FILLER_0_21_28/a_484_472# 0.001795f
C1100 cal_itt\[2\] _260_/a_36_68# 0.004081f
C1101 _076_ net47 0.00115f
C1102 net15 FILLER_0_9_60/a_572_375# 0.047331f
C1103 net29 vdd 0.611195f
C1104 FILLER_0_7_146/a_124_375# calibrate 0.014163f
C1105 FILLER_0_12_2/a_124_375# net67 0.003339f
C1106 net62 output29/a_224_472# 0.138536f
C1107 _371_/a_36_113# FILLER_0_2_127/a_124_375# 0.002437f
C1108 FILLER_0_5_164/a_124_375# _066_ 0.006762f
C1109 _120_ net51 1.716752f
C1110 ctlp[1] _419_/a_796_472# 0.001178f
C1111 FILLER_0_17_72/a_1916_375# net53 0.001657f
C1112 net82 _083_ 0.010347f
C1113 _177_ _095_ 0.004392f
C1114 _093_ FILLER_0_17_142/a_484_472# 0.011974f
C1115 FILLER_0_10_78/a_484_472# FILLER_0_9_72/a_1020_375# 0.001543f
C1116 net52 FILLER_0_2_165/a_36_472# 0.002601f
C1117 _448_/a_448_472# net22 0.085004f
C1118 FILLER_0_8_107/a_36_472# _219_/a_36_160# 0.002767f
C1119 net9 _082_ 0.001006f
C1120 _434_/a_1308_423# mask\[6\] 0.022677f
C1121 net65 _073_ 0.775972f
C1122 output11/a_224_472# ctln[3] 0.068614f
C1123 FILLER_0_16_73/a_484_472# _176_ 0.010681f
C1124 ctln[6] net52 0.1064f
C1125 FILLER_0_7_72/a_1916_375# _376_/a_36_160# 0.001925f
C1126 FILLER_0_16_57/a_124_375# _183_ 0.005825f
C1127 net69 _159_ 0.010086f
C1128 FILLER_0_10_37/a_36_472# net16 0.012905f
C1129 net16 _408_/a_1936_472# 0.022235f
C1130 result[7] FILLER_0_24_274/a_484_472# 0.006641f
C1131 FILLER_0_4_99/a_36_472# _153_ 0.066147f
C1132 cal_itt\[3\] _161_ 0.20195f
C1133 FILLER_0_9_28/a_2364_375# _220_/a_67_603# 0.002082f
C1134 FILLER_0_15_212/a_1468_375# vss 0.060206f
C1135 FILLER_0_15_212/a_36_472# vdd 0.105575f
C1136 _093_ FILLER_0_18_76/a_36_472# 0.129892f
C1137 _440_/a_2665_112# _160_ 0.008418f
C1138 state\[0\] _426_/a_2665_112# 0.017088f
C1139 FILLER_0_22_86/a_484_472# _437_/a_448_472# 0.008036f
C1140 FILLER_0_6_90/a_572_375# net14 0.031929f
C1141 _091_ fanout56/a_36_113# 0.001254f
C1142 _422_/a_36_151# net19 0.033614f
C1143 _227_/a_36_160# FILLER_0_8_156/a_124_375# 0.005398f
C1144 FILLER_0_24_274/a_932_472# FILLER_0_23_282/a_36_472# 0.05841f
C1145 net16 _184_ 0.028159f
C1146 _020_ _136_ 0.022753f
C1147 state\[0\] _060_ 0.047136f
C1148 FILLER_0_5_164/a_124_375# net37 0.008158f
C1149 valid fanout64/a_36_160# 0.001811f
C1150 mask\[5\] net35 0.003646f
C1151 net31 net36 0.00943f
C1152 _415_/a_2248_156# result[1] 0.010922f
C1153 net79 _056_ 0.022406f
C1154 _118_ _059_ 0.022651f
C1155 FILLER_0_10_78/a_1020_375# net52 0.001158f
C1156 net66 net40 0.124825f
C1157 _124_ FILLER_0_10_107/a_484_472# 0.00438f
C1158 state\[1\] _090_ 0.087906f
C1159 net39 _034_ 0.004367f
C1160 _073_ net59 0.028673f
C1161 result[5] result[4] 0.090472f
C1162 _397_/a_36_472# net55 0.039732f
C1163 _086_ FILLER_0_11_135/a_36_472# 0.004074f
C1164 _431_/a_2665_112# net53 0.004057f
C1165 net16 FILLER_0_8_37/a_36_472# 0.012905f
C1166 cal_count\[3\] _067_ 0.478427f
C1167 FILLER_0_4_91/a_572_375# _156_ 0.004958f
C1168 _420_/a_796_472# _009_ 0.012395f
C1169 net34 FILLER_0_22_177/a_932_472# 0.003953f
C1170 _445_/a_1308_423# net40 0.046345f
C1171 net74 _390_/a_36_68# 0.008011f
C1172 net80 _434_/a_1204_472# 0.003997f
C1173 _144_ _049_ 0.100508f
C1174 mask\[4\] FILLER_0_18_177/a_1916_375# 0.013466f
C1175 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_124_375# 0.026339f
C1176 net48 _014_ 0.276733f
C1177 _308_/a_848_380# FILLER_0_9_105/a_124_375# 0.005599f
C1178 _443_/a_36_151# net13 0.001896f
C1179 _443_/a_1308_423# net23 0.034115f
C1180 FILLER_0_20_177/a_124_375# vdd 0.001964f
C1181 mask\[3\] _098_ 0.026156f
C1182 FILLER_0_17_226/a_124_375# mask\[3\] 0.010642f
C1183 net50 _441_/a_1000_472# 0.02354f
C1184 net52 _441_/a_2248_156# 0.023959f
C1185 FILLER_0_9_28/a_1828_472# net16 0.001946f
C1186 trimb[4] cal_count\[2\] 0.146942f
C1187 _442_/a_2665_112# _157_ 0.001587f
C1188 net38 _221_/a_36_160# 0.029767f
C1189 FILLER_0_4_49/a_36_472# net66 0.012791f
C1190 FILLER_0_13_212/a_36_472# net79 0.006158f
C1191 FILLER_0_12_136/a_1380_472# FILLER_0_13_142/a_572_375# 0.001684f
C1192 _053_ net23 0.031487f
C1193 ctln[6] _387_/a_36_113# 0.007687f
C1194 _086_ _161_ 0.077837f
C1195 _430_/a_1000_472# mask\[2\] 0.00785f
C1196 FILLER_0_16_89/a_36_472# _451_/a_448_472# 0.011974f
C1197 net50 _447_/a_448_472# 0.001219f
C1198 state\[1\] net22 0.007096f
C1199 _096_ _320_/a_1568_472# 0.001632f
C1200 net63 _432_/a_36_151# 0.001392f
C1201 mask\[4\] _092_ 0.072581f
C1202 FILLER_0_18_61/a_36_472# vss 0.00605f
C1203 _092_ net22 0.010937f
C1204 net73 FILLER_0_17_104/a_1380_472# 0.003206f
C1205 FILLER_0_16_255/a_124_375# net30 0.001055f
C1206 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_124_375# 0.012001f
C1207 net40 _167_ 0.020177f
C1208 FILLER_0_10_78/a_484_472# _115_ 0.005678f
C1209 net50 _439_/a_796_472# 0.002389f
C1210 net52 _439_/a_1204_472# 0.027632f
C1211 _070_ FILLER_0_11_109/a_124_375# 0.002358f
C1212 FILLER_0_17_104/a_1468_375# vss 0.001786f
C1213 FILLER_0_17_104/a_36_472# vdd 0.095484f
C1214 FILLER_0_5_54/a_484_472# FILLER_0_6_47/a_1380_472# 0.026657f
C1215 FILLER_0_5_54/a_1468_375# FILLER_0_6_47/a_2276_472# 0.001597f
C1216 _425_/a_1000_472# net37 0.002879f
C1217 _067_ net40 0.040115f
C1218 result[7] _419_/a_36_151# 0.001036f
C1219 net28 net36 0.002537f
C1220 cal_count\[2\] cal_count\[1\] 0.067712f
C1221 _434_/a_448_472# _023_ 0.03093f
C1222 net41 FILLER_0_21_28/a_484_472# 0.060027f
C1223 net16 net47 0.089651f
C1224 net74 FILLER_0_11_124/a_36_472# 0.020589f
C1225 _053_ _439_/a_2248_156# 0.002486f
C1226 FILLER_0_21_286/a_572_375# net77 0.044323f
C1227 ctlp[1] FILLER_0_23_282/a_124_375# 0.00324f
C1228 mask\[8\] _437_/a_36_151# 0.005179f
C1229 ctln[1] FILLER_0_3_221/a_1020_375# 0.001554f
C1230 net15 _453_/a_2560_156# 0.049334f
C1231 _422_/a_36_151# _009_ 0.015085f
C1232 _030_ FILLER_0_3_78/a_572_375# 0.007667f
C1233 net49 FILLER_0_3_78/a_124_375# 0.001597f
C1234 cal_itt\[2\] net65 0.514538f
C1235 _068_ _059_ 0.255081f
C1236 _012_ FILLER_0_23_60/a_124_375# 0.002827f
C1237 net69 FILLER_0_2_111/a_932_472# 0.011453f
C1238 _031_ FILLER_0_2_111/a_36_472# 0.034656f
C1239 net48 _070_ 0.264809f
C1240 FILLER_0_5_109/a_572_375# _153_ 0.03228f
C1241 FILLER_0_4_49/a_36_472# _167_ 0.063278f
C1242 _004_ fanout79/a_36_160# 0.048599f
C1243 net44 _452_/a_2225_156# 0.044858f
C1244 _429_/a_36_151# FILLER_0_15_212/a_1020_375# 0.035849f
C1245 net65 net1 0.035488f
C1246 _077_ FILLER_0_8_239/a_124_375# 0.001772f
C1247 _069_ FILLER_0_13_206/a_36_472# 0.005793f
C1248 FILLER_0_20_15/a_1468_375# net40 0.030032f
C1249 FILLER_0_19_171/a_1020_375# vdd 0.025918f
C1250 FILLER_0_20_87/a_36_472# net14 0.001471f
C1251 _091_ FILLER_0_13_212/a_124_375# 0.025558f
C1252 FILLER_0_4_123/a_36_472# _370_/a_124_24# 0.003595f
C1253 _205_/a_36_160# net21 0.020847f
C1254 ctlp[5] vss 0.032166f
C1255 FILLER_0_15_235/a_572_375# vss 0.002683f
C1256 FILLER_0_15_235/a_36_472# vdd 0.019127f
C1257 _114_ _311_/a_2180_473# 0.00515f
C1258 trim_val\[3\] vss 0.249446f
C1259 net78 _421_/a_36_151# 0.001368f
C1260 FILLER_0_4_177/a_572_375# FILLER_0_5_181/a_124_375# 0.05841f
C1261 FILLER_0_18_177/a_2812_375# net21 0.048071f
C1262 output42/a_224_472# FILLER_0_8_24/a_124_375# 0.001168f
C1263 _115_ _120_ 0.076035f
C1264 _093_ net54 0.003211f
C1265 _438_/a_36_151# vdd 0.111691f
C1266 _144_ _433_/a_1204_472# 0.009472f
C1267 _412_/a_36_151# net65 0.015454f
C1268 net52 _154_ 0.001512f
C1269 _307_/a_672_472# _113_ 0.006607f
C1270 _104_ _010_ 0.252687f
C1271 _063_ net49 0.002854f
C1272 _079_ FILLER_0_5_212/a_124_375# 0.005363f
C1273 result[2] FILLER_0_13_290/a_124_375# 0.015011f
C1274 ctln[7] net52 0.06558f
C1275 _322_/a_848_380# _062_ 0.001872f
C1276 mask\[5\] FILLER_0_18_177/a_2276_472# 0.001063f
C1277 cal_itt\[2\] net59 0.014956f
C1278 cal_count\[3\] _121_ 0.011368f
C1279 FILLER_0_14_91/a_572_375# _095_ 0.011885f
C1280 _114_ _061_ 0.123371f
C1281 _424_/a_2665_112# net36 0.028938f
C1282 FILLER_0_0_130/a_36_472# vdd 0.050082f
C1283 FILLER_0_0_130/a_124_375# vss 0.018073f
C1284 _322_/a_1084_68# _118_ 0.002515f
C1285 FILLER_0_14_81/a_124_375# _177_ 0.002725f
C1286 net21 mask\[6\] 0.634881f
C1287 net4 net18 0.034592f
C1288 net1 net59 0.920133f
C1289 _054_ vdd 0.360345f
C1290 _008_ _419_/a_36_151# 0.014476f
C1291 _431_/a_2248_156# _427_/a_36_151# 0.001081f
C1292 net38 _178_ 0.123812f
C1293 _415_/a_1308_423# FILLER_0_9_270/a_124_375# 0.001064f
C1294 _017_ FILLER_0_14_107/a_484_472# 0.004583f
C1295 result[6] _010_ 0.056004f
C1296 _354_/a_49_472# net71 0.010421f
C1297 net70 FILLER_0_14_107/a_1380_472# 0.003355f
C1298 _106_ _293_/a_36_472# 0.04279f
C1299 FILLER_0_20_98/a_36_472# vss 0.00206f
C1300 _230_/a_244_68# net21 0.00165f
C1301 _360_/a_36_160# net74 0.001912f
C1302 FILLER_0_16_57/a_36_472# cal_count\[2\] 0.001952f
C1303 _067_ FILLER_0_12_20/a_124_375# 0.017026f
C1304 _123_ FILLER_0_6_231/a_572_375# 0.00487f
C1305 _412_/a_36_151# net59 0.003938f
C1306 FILLER_0_10_78/a_1380_472# _308_/a_124_24# 0.037778f
C1307 _086_ _127_ 0.042698f
C1308 _074_ _062_ 0.005012f
C1309 _420_/a_1000_472# vss 0.002146f
C1310 result[9] _421_/a_1308_423# 0.011854f
C1311 _292_/a_36_160# _105_ 0.027405f
C1312 output25/a_224_472# _051_ 0.019651f
C1313 _431_/a_1204_472# _137_ 0.005886f
C1314 _100_ _283_/a_36_472# 0.033597f
C1315 _430_/a_448_472# net81 0.003775f
C1316 net53 _451_/a_36_151# 0.030715f
C1317 net70 _451_/a_1040_527# 0.002679f
C1318 _084_ _082_ 0.044645f
C1319 _115_ FILLER_0_9_105/a_572_375# 0.003191f
C1320 _109_ vss 0.023215f
C1321 FILLER_0_8_127/a_124_375# _119_ 0.013315f
C1322 ctln[1] FILLER_0_1_266/a_36_472# 0.002068f
C1323 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_572_375# 0.086635f
C1324 net20 _419_/a_1204_472# 0.006482f
C1325 _230_/a_244_68# _070_ 0.001641f
C1326 FILLER_0_16_241/a_36_472# _099_ 0.158391f
C1327 net19 _419_/a_1000_472# 0.012949f
C1328 _442_/a_2248_156# _158_ 0.001288f
C1329 mask\[9\] _438_/a_2248_156# 0.036436f
C1330 _093_ FILLER_0_18_139/a_484_472# 0.008683f
C1331 _236_/a_36_160# net39 0.052649f
C1332 FILLER_0_18_209/a_124_375# _047_ 0.006317f
C1333 FILLER_0_5_181/a_124_375# net22 0.00205f
C1334 _395_/a_36_488# _176_ 0.010116f
C1335 _395_/a_1044_488# _085_ 0.00391f
C1336 FILLER_0_24_130/a_124_375# _050_ 0.007643f
C1337 output36/a_224_472# FILLER_0_15_282/a_36_472# 0.008834f
C1338 _376_/a_36_160# FILLER_0_6_79/a_124_375# 0.004736f
C1339 _177_ cal_count\[1\] 0.03631f
C1340 FILLER_0_3_172/a_3260_375# net22 0.015274f
C1341 _434_/a_1000_472# vdd 0.032431f
C1342 ctln[8] _168_ 0.001145f
C1343 _427_/a_36_151# _043_ 0.002267f
C1344 FILLER_0_13_142/a_36_472# vdd 0.104785f
C1345 fanout53/a_36_160# vss 0.006674f
C1346 FILLER_0_13_142/a_1468_375# vss 0.00614f
C1347 FILLER_0_4_177/a_124_375# vss 0.002462f
C1348 FILLER_0_4_177/a_572_375# vdd 0.001622f
C1349 net57 FILLER_0_8_156/a_36_472# 0.001544f
C1350 FILLER_0_21_133/a_36_472# vss 0.004298f
C1351 _417_/a_36_151# vss 0.040392f
C1352 _429_/a_796_472# _018_ 0.002291f
C1353 net67 output6/a_224_472# 0.070024f
C1354 FILLER_0_4_99/a_124_375# _160_ 0.005563f
C1355 FILLER_0_5_128/a_124_375# net47 0.011156f
C1356 FILLER_0_12_124/a_124_375# vdd -0.00168f
C1357 _077_ _449_/a_36_151# 0.002475f
C1358 net7 vss 0.117948f
C1359 _086_ _071_ 0.041029f
C1360 _104_ vdd 0.662413f
C1361 FILLER_0_8_247/a_1380_472# vss 0.001338f
C1362 _322_/a_1084_68# _068_ 0.001022f
C1363 _052_ FILLER_0_18_53/a_572_375# 0.001631f
C1364 _095_ _402_/a_56_567# 0.010012f
C1365 _421_/a_2665_112# vdd 0.029293f
C1366 _415_/a_1308_423# net18 0.010051f
C1367 _132_ FILLER_0_14_107/a_1380_472# 0.049391f
C1368 net49 net14 0.00344f
C1369 _239_/a_36_160# _064_ 0.001292f
C1370 state\[0\] net64 0.01679f
C1371 FILLER_0_21_142/a_124_375# vss 0.009345f
C1372 _442_/a_2248_156# net14 0.025334f
C1373 output27/a_224_472# vdd 0.070751f
C1374 _067_ FILLER_0_13_80/a_124_375# 0.001857f
C1375 _096_ _136_ 0.022182f
C1376 net50 FILLER_0_7_59/a_484_472# 0.011974f
C1377 _130_ _114_ 0.002404f
C1378 _422_/a_1308_423# vdd 0.004083f
C1379 FILLER_0_5_128/a_484_472# _370_/a_124_24# 0.00171f
C1380 _115_ _227_/a_36_160# 0.00124f
C1381 _426_/a_1204_472# vdd 0.003412f
C1382 output38/a_224_472# _035_ 0.091395f
C1383 _265_/a_244_68# _084_ 0.016463f
C1384 _093_ FILLER_0_18_107/a_1020_375# 0.006376f
C1385 _359_/a_36_488# _129_ 0.002527f
C1386 _098_ FILLER_0_20_87/a_36_472# 0.016138f
C1387 FILLER_0_15_282/a_572_375# vss 0.058168f
C1388 FILLER_0_15_282/a_36_472# vdd 0.10628f
C1389 net81 _415_/a_36_151# 0.046145f
C1390 result[6] vdd 0.513079f
C1391 _446_/a_2665_112# net40 0.027712f
C1392 net19 _192_/a_67_603# 0.003106f
C1393 net36 FILLER_0_15_205/a_36_472# 0.005101f
C1394 FILLER_0_11_101/a_484_472# vdd 0.009482f
C1395 FILLER_0_11_101/a_36_472# vss 0.001641f
C1396 mask\[5\] FILLER_0_21_206/a_36_472# 0.019416f
C1397 output24/a_224_472# net71 0.001495f
C1398 _090_ vdd 0.751973f
C1399 net69 _441_/a_1308_423# 0.016223f
C1400 _185_ _180_ 0.001053f
C1401 fanout61/a_36_113# vdd 0.108255f
C1402 FILLER_0_9_223/a_36_472# _077_ 0.005511f
C1403 _072_ _128_ 0.072191f
C1404 _064_ _036_ 0.003286f
C1405 trim_mask\[2\] trim_val\[3\] 0.003342f
C1406 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_124_375# 0.012222f
C1407 FILLER_0_4_49/a_572_375# _164_ 0.005532f
C1408 net71 _437_/a_796_472# 0.006933f
C1409 FILLER_0_7_162/a_36_472# _081_ 0.002493f
C1410 net63 FILLER_0_15_212/a_1020_375# 0.001012f
C1411 _445_/a_448_472# net66 0.010949f
C1412 _064_ _445_/a_2665_112# 0.004701f
C1413 _053_ _363_/a_36_68# 0.021227f
C1414 net66 trim[3] 0.00567f
C1415 cal_count\[3\] FILLER_0_11_124/a_124_375# 0.002147f
C1416 net46 FILLER_0_20_15/a_572_375# 0.029486f
C1417 output12/a_224_472# vss 0.013728f
C1418 _127_ FILLER_0_9_142/a_124_375# 0.005447f
C1419 _413_/a_1204_472# vdd 0.001027f
C1420 ctlp[2] net33 0.004972f
C1421 output25/a_224_472# vdd 0.03413f
C1422 _431_/a_36_151# vdd 0.145005f
C1423 _420_/a_448_472# net77 0.001276f
C1424 _132_ _140_ 0.019255f
C1425 mask\[4\] vdd 0.794539f
C1426 FILLER_0_18_100/a_36_472# _136_ 0.003419f
C1427 _127_ net53 0.00917f
C1428 net22 vdd 1.920713f
C1429 _029_ trim_mask\[1\] 1.002118f
C1430 net20 _274_/a_716_497# 0.001321f
C1431 result[9] FILLER_0_24_274/a_932_472# 0.001826f
C1432 _439_/a_2248_156# trim_mask\[0\] 0.005416f
C1433 result[4] net60 0.244453f
C1434 _274_/a_36_68# _069_ 0.02257f
C1435 FILLER_0_8_24/a_572_375# net40 0.038492f
C1436 _068_ _247_/a_36_160# 0.003213f
C1437 fanout70/a_36_113# net73 0.21211f
C1438 _091_ _323_/a_36_113# 0.001651f
C1439 ctlp[5] mask\[7\] 0.131468f
C1440 FILLER_0_17_56/a_36_472# _041_ 0.004881f
C1441 FILLER_0_3_78/a_36_472# _164_ 0.022063f
C1442 net73 FILLER_0_18_107/a_2724_472# 0.02814f
C1443 _081_ FILLER_0_5_148/a_572_375# 0.01425f
C1444 net75 _426_/a_1204_472# 0.001592f
C1445 output32/a_224_472# _418_/a_448_472# 0.008149f
C1446 net32 _011_ 0.072502f
C1447 _043_ FILLER_0_13_72/a_36_472# 0.017766f
C1448 net26 net40 0.001136f
C1449 _093_ FILLER_0_18_209/a_572_375# 0.064723f
C1450 FILLER_0_2_101/a_36_472# trim_mask\[3\] 0.013363f
C1451 fanout67/a_36_160# _220_/a_67_603# 0.005474f
C1452 net15 vss 1.330044f
C1453 FILLER_0_18_107/a_1380_472# vdd 0.009462f
C1454 _076_ _385_/a_36_68# 0.006512f
C1455 FILLER_0_7_72/a_932_472# _077_ 0.001315f
C1456 _406_/a_36_159# _278_/a_36_160# 0.001331f
C1457 net79 net18 0.222939f
C1458 _217_/a_36_160# vdd 0.092586f
C1459 FILLER_0_20_2/a_484_472# net43 0.005543f
C1460 _208_/a_36_160# FILLER_0_22_128/a_3260_375# 0.001948f
C1461 _049_ FILLER_0_22_128/a_3172_472# 0.01125f
C1462 FILLER_0_18_100/a_36_472# _356_/a_36_472# 0.010679f
C1463 FILLER_0_14_107/a_36_472# _451_/a_36_151# 0.001723f
C1464 FILLER_0_3_204/a_36_472# vss 0.003572f
C1465 net54 FILLER_0_22_128/a_932_472# 0.014735f
C1466 _026_ _437_/a_36_151# 0.012193f
C1467 _149_ _437_/a_1308_423# 0.015677f
C1468 net10 FILLER_0_0_232/a_124_375# 0.022977f
C1469 _292_/a_36_160# _047_ 0.001291f
C1470 FILLER_0_16_89/a_1380_472# vss 0.005351f
C1471 FILLER_0_10_214/a_124_375# _070_ 0.017713f
C1472 output43/a_224_472# output46/a_224_472# 0.292611f
C1473 fanout77/a_36_113# net77 0.031558f
C1474 _275_/a_224_472# mask\[3\] 0.002528f
C1475 _035_ vdd 0.215473f
C1476 net69 _367_/a_36_68# 0.008893f
C1477 FILLER_0_13_142/a_572_375# net23 0.009573f
C1478 _119_ FILLER_0_7_162/a_36_472# 0.005739f
C1479 _119_ _324_/a_224_472# 0.00368f
C1480 _425_/a_1204_472# calibrate 0.009749f
C1481 _413_/a_36_151# FILLER_0_1_192/a_36_472# 0.046516f
C1482 _155_ vdd 0.193832f
C1483 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_572_375# 0.001597f
C1484 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_36_472# 0.026657f
C1485 FILLER_0_7_72/a_3172_472# FILLER_0_7_104/a_36_472# 0.013276f
C1486 _204_/a_67_603# _201_/a_67_603# 0.001129f
C1487 FILLER_0_5_117/a_36_472# _163_ 0.007418f
C1488 _087_ FILLER_0_6_177/a_124_375# 0.001151f
C1489 _038_ vdd 0.043998f
C1490 FILLER_0_21_133/a_124_375# _140_ 0.018383f
C1491 valid net19 0.00646f
C1492 mask\[5\] output35/a_224_472# 0.003461f
C1493 net11 vdd 0.330644f
C1494 net20 FILLER_0_3_221/a_1380_472# 0.008749f
C1495 FILLER_0_5_117/a_124_375# FILLER_0_4_107/a_1380_472# 0.001684f
C1496 _057_ _267_/a_1792_472# 0.003005f
C1497 _408_/a_56_524# FILLER_0_12_20/a_572_375# 0.009967f
C1498 _077_ FILLER_0_9_60/a_572_375# 0.018665f
C1499 FILLER_0_16_255/a_124_375# _417_/a_2665_112# 0.003856f
C1500 _186_ vss 0.0718f
C1501 _413_/a_36_151# FILLER_0_3_172/a_1828_472# 0.001723f
C1502 mask\[7\] _109_ 0.028117f
C1503 ctln[1] vdd 0.825166f
C1504 FILLER_0_22_177/a_484_472# mask\[6\] 0.006573f
C1505 FILLER_0_22_177/a_124_375# _146_ 0.001864f
C1506 _074_ _316_/a_124_24# 0.018608f
C1507 result[9] _419_/a_448_472# 0.015767f
C1508 _176_ _040_ 0.272465f
C1509 _132_ _149_ 0.087289f
C1510 _176_ _125_ 0.089769f
C1511 net73 mask\[9\] 0.383862f
C1512 net62 _005_ 0.097739f
C1513 _187_ _181_ 0.001158f
C1514 _325_/a_224_472# _129_ 0.003137f
C1515 _114_ _428_/a_2248_156# 0.004516f
C1516 net54 FILLER_0_22_107/a_124_375# 0.003502f
C1517 _432_/a_2560_156# _091_ 0.001542f
C1518 output48/a_224_472# net2 0.06309f
C1519 _133_ vss 0.18326f
C1520 _076_ vdd 0.806117f
C1521 net81 FILLER_0_15_228/a_36_472# 0.003953f
C1522 _449_/a_1000_472# vss 0.029565f
C1523 net50 FILLER_0_6_90/a_484_472# 0.012286f
C1524 _067_ _120_ 0.031156f
C1525 net72 _217_/a_36_160# 0.068583f
C1526 FILLER_0_21_133/a_36_472# mask\[7\] 0.003404f
C1527 _091_ FILLER_0_17_218/a_572_375# 0.001927f
C1528 _430_/a_2248_156# net36 0.001198f
C1529 FILLER_0_5_109/a_124_375# _151_ 0.003377f
C1530 net55 FILLER_0_18_37/a_1380_472# 0.007432f
C1531 _151_ _163_ 0.501188f
C1532 _450_/a_36_151# net6 0.035997f
C1533 _450_/a_1040_527# output6/a_224_472# 0.005581f
C1534 trim_mask\[4\] _386_/a_124_24# 0.040347f
C1535 net2 net5 0.47659f
C1536 FILLER_0_17_72/a_3260_375# vdd 0.007427f
C1537 _376_/a_36_160# vss 0.03081f
C1538 _093_ net30 0.001859f
C1539 _127_ FILLER_0_11_135/a_36_472# 0.044488f
C1540 _009_ FILLER_0_23_282/a_572_375# 0.016879f
C1541 FILLER_0_8_247/a_36_472# calibrate 0.008647f
C1542 net19 net9 0.342451f
C1543 _028_ _363_/a_36_68# 0.015609f
C1544 _421_/a_2248_156# mask\[7\] 0.016229f
C1545 _053_ FILLER_0_5_54/a_124_375# 0.001571f
C1546 _081_ net23 0.081773f
C1547 net27 _415_/a_2248_156# 0.022666f
C1548 net60 _421_/a_36_151# 0.224039f
C1549 FILLER_0_22_86/a_36_472# vdd -0.001506f
C1550 FILLER_0_22_86/a_1468_375# vss 0.013146f
C1551 _418_/a_36_151# vss 0.041728f
C1552 _090_ _279_/a_244_68# 0.001986f
C1553 net33 _434_/a_448_472# 0.003049f
C1554 _422_/a_448_472# mask\[7\] 0.048658f
C1555 output32/a_224_472# result[7] 0.063135f
C1556 net52 _443_/a_796_472# 0.004334f
C1557 _419_/a_2248_156# vdd 0.040646f
C1558 _450_/a_448_472# net40 0.00222f
C1559 net72 _038_ 0.013821f
C1560 _426_/a_448_472# calibrate 0.002745f
C1561 _176_ _174_ 0.00677f
C1562 net29 _099_ 0.358926f
C1563 _411_/a_2248_156# net8 0.06032f
C1564 FILLER_0_21_142/a_36_472# FILLER_0_22_128/a_1468_375# 0.001543f
C1565 FILLER_0_13_206/a_36_472# net22 0.053292f
C1566 mask\[5\] FILLER_0_19_195/a_36_472# 0.007596f
C1567 net75 ctln[1] 0.159105f
C1568 cal net5 0.039735f
C1569 _453_/a_1000_472# _042_ 0.004985f
C1570 fanout53/a_36_160# _427_/a_2248_156# 0.027388f
C1571 net74 _159_ 0.129233f
C1572 FILLER_0_16_89/a_1020_375# net14 0.029702f
C1573 _348_/a_665_69# _146_ 0.001153f
C1574 result[7] _010_ 0.054533f
C1575 state\[2\] vss 0.185787f
C1576 FILLER_0_4_107/a_1020_375# net47 0.011446f
C1577 _217_/a_36_160# _424_/a_36_151# 0.035111f
C1578 net15 _441_/a_1204_472# 0.005939f
C1579 net34 FILLER_0_22_128/a_2812_375# 0.005158f
C1580 _178_ FILLER_0_15_10/a_36_472# 0.001356f
C1581 net15 trim_mask\[2\] 0.026132f
C1582 FILLER_0_4_99/a_124_375# _156_ 0.081915f
C1583 net15 FILLER_0_11_64/a_124_375# 0.047331f
C1584 _437_/a_2665_112# vss 0.002056f
C1585 _437_/a_2560_156# vdd 0.0026f
C1586 sample fanout59/a_36_160# 0.001854f
C1587 output47/a_224_472# net38 0.082174f
C1588 _449_/a_1308_423# net55 0.001985f
C1589 output19/a_224_472# _107_ 0.005034f
C1590 _131_ _041_ 0.035642f
C1591 _429_/a_36_151# _136_ 0.001188f
C1592 _105_ _422_/a_2665_112# 0.011125f
C1593 FILLER_0_8_239/a_36_472# calibrate 0.008683f
C1594 mask\[5\] _346_/a_49_472# 0.037629f
C1595 _086_ net23 0.037804f
C1596 _429_/a_36_151# net21 0.054289f
C1597 FILLER_0_4_177/a_484_472# net76 0.006746f
C1598 ctln[0] vdd 0.051631f
C1599 FILLER_0_17_282/a_124_375# _006_ 0.004694f
C1600 net20 _077_ 0.094476f
C1601 fanout59/a_36_160# vss 0.010949f
C1602 _415_/a_1204_472# vdd 0.00108f
C1603 fanout62/a_36_160# net64 0.052109f
C1604 FILLER_0_7_72/a_36_472# _439_/a_448_472# 0.008036f
C1605 net63 _434_/a_1308_423# 0.003686f
C1606 FILLER_0_17_56/a_124_375# _183_ 0.019253f
C1607 net50 FILLER_0_5_88/a_124_375# 0.03181f
C1608 _068_ _229_/a_224_472# 0.002601f
C1609 _131_ FILLER_0_14_123/a_36_472# 0.029747f
C1610 net15 _439_/a_1000_472# 0.001798f
C1611 FILLER_0_22_177/a_36_472# _023_ 0.007019f
C1612 FILLER_0_17_72/a_2276_472# mask\[9\] 0.006767f
C1613 _029_ _164_ 0.031781f
C1614 _446_/a_2248_156# net66 0.002766f
C1615 _063_ net47 0.142088f
C1616 _430_/a_1000_472# vss 0.001626f
C1617 net52 _387_/a_36_113# 0.02405f
C1618 trim_mask\[4\] vss 0.641217f
C1619 _062_ _226_/a_452_68# 0.001697f
C1620 _112_ calibrate 0.024557f
C1621 mask\[3\] _137_ 0.231419f
C1622 FILLER_0_18_171/a_124_375# mask\[3\] 0.001156f
C1623 FILLER_0_5_72/a_1020_375# net49 0.002208f
C1624 _415_/a_36_151# net64 0.001735f
C1625 _119_ net23 0.0245f
C1626 _443_/a_36_151# _170_ 0.014771f
C1627 fanout64/a_36_160# calibrate 0.001117f
C1628 _077_ _453_/a_2560_156# 0.001286f
C1629 output32/a_224_472# _008_ 0.074809f
C1630 _043_ FILLER_0_15_180/a_36_472# 0.001219f
C1631 _414_/a_2248_156# net22 0.062122f
C1632 net76 FILLER_0_3_172/a_124_375# 0.001186f
C1633 FILLER_0_7_72/a_1468_375# vdd 0.001135f
C1634 en_co_clk FILLER_0_13_100/a_36_472# 0.001752f
C1635 _256_/a_1612_497# vss 0.004265f
C1636 FILLER_0_10_78/a_124_375# _453_/a_2665_112# 0.006271f
C1637 FILLER_0_19_47/a_36_472# _052_ 0.015772f
C1638 FILLER_0_11_78/a_36_472# vss 0.00471f
C1639 FILLER_0_11_78/a_484_472# vdd 0.001756f
C1640 _121_ _120_ 0.069685f
C1641 ctln[2] FILLER_0_0_266/a_124_375# 0.041898f
C1642 net81 net76 0.236554f
C1643 fanout49/a_36_160# _440_/a_2665_112# 0.00631f
C1644 FILLER_0_5_72/a_36_472# trim_mask\[1\] 0.015775f
C1645 FILLER_0_5_72/a_1380_472# _029_ 0.007385f
C1646 net80 _146_ 0.021227f
C1647 FILLER_0_6_47/a_2364_375# vss 0.008275f
C1648 FILLER_0_6_47/a_2812_375# vdd 0.002455f
C1649 output10/a_224_472# net9 0.003212f
C1650 _261_/a_36_160# _163_ 0.002002f
C1651 net26 _423_/a_1204_472# 0.001069f
C1652 output29/a_224_472# net18 0.010345f
C1653 _444_/a_1308_423# _054_ 0.005457f
C1654 net16 vdd 2.255325f
C1655 cal_itt\[3\] _056_ 0.023192f
C1656 _411_/a_2665_112# vss 0.00238f
C1657 FILLER_0_12_20/a_124_375# _450_/a_448_472# 0.001597f
C1658 output39/a_224_472# net17 0.041253f
C1659 FILLER_0_18_171/a_36_472# _432_/a_36_151# 0.059367f
C1660 net43 vss 0.132286f
C1661 net34 net61 0.037731f
C1662 _414_/a_1000_472# _074_ 0.00222f
C1663 output44/a_224_472# vss 0.014054f
C1664 FILLER_0_17_218/a_36_472# _069_ 0.001246f
C1665 FILLER_0_7_104/a_1380_472# _154_ 0.002799f
C1666 _118_ _311_/a_66_473# 0.008528f
C1667 _432_/a_2665_112# vdd 0.009104f
C1668 cal_count\[3\] _453_/a_1000_472# 0.001123f
C1669 FILLER_0_21_286/a_36_472# net18 0.18097f
C1670 _422_/a_1000_472# _108_ 0.027806f
C1671 cal FILLER_0_1_266/a_572_375# 0.001707f
C1672 FILLER_0_21_142/a_124_375# _433_/a_448_472# 0.006782f
C1673 _115_ FILLER_0_10_107/a_484_472# 0.017642f
C1674 fanout68/a_36_113# net17 0.001252f
C1675 FILLER_0_16_107/a_36_472# net36 0.001245f
C1676 _077_ FILLER_0_7_72/a_2724_472# 0.004635f
C1677 result[7] vdd 0.500292f
C1678 FILLER_0_13_100/a_124_375# net14 0.041373f
C1679 FILLER_0_16_107/a_572_375# net14 0.002308f
C1680 _210_/a_67_603# _436_/a_2665_112# 0.007103f
C1681 _055_ net21 0.025995f
C1682 _072_ _395_/a_1492_488# 0.003088f
C1683 net32 _102_ 0.038622f
C1684 ctln[3] FILLER_0_0_232/a_36_472# 0.015594f
C1685 net34 _049_ 0.048403f
C1686 net57 net36 0.087967f
C1687 FILLER_0_23_282/a_36_472# vss 0.003317f
C1688 _069_ FILLER_0_15_212/a_124_375# 0.039975f
C1689 FILLER_0_24_63/a_124_375# vss 0.03143f
C1690 FILLER_0_21_28/a_3172_472# _012_ 0.018785f
C1691 _390_/a_244_472# _067_ 0.004031f
C1692 trim_mask\[4\] FILLER_0_2_165/a_124_375# 0.011181f
C1693 output33/a_224_472# net61 0.04987f
C1694 _320_/a_1792_472# net79 0.002091f
C1695 _174_ _183_ 0.008231f
C1696 fanout69/a_36_113# vss 0.002239f
C1697 cal_itt\[1\] FILLER_0_3_221/a_1380_472# 0.004939f
C1698 _445_/a_1000_472# _034_ 0.007034f
C1699 _445_/a_2665_112# _166_ 0.002292f
C1700 _062_ FILLER_0_8_156/a_124_375# 0.008116f
C1701 _394_/a_728_93# _043_ 0.00355f
C1702 _433_/a_796_472# _022_ 0.025882f
C1703 ctlp[1] FILLER_0_23_290/a_124_375# 0.053745f
C1704 _027_ net36 0.185347f
C1705 _408_/a_56_524# _067_ 0.003678f
C1706 net45 vdd 0.087369f
C1707 net70 net14 0.106631f
C1708 FILLER_0_12_136/a_1380_472# _127_ 0.001432f
C1709 FILLER_0_15_142/a_124_375# _136_ 0.001706f
C1710 net20 net37 0.039674f
C1711 FILLER_0_2_93/a_484_472# vss 0.003689f
C1712 _070_ _055_ 0.516713f
C1713 _411_/a_2560_156# vdd 0.001315f
C1714 net55 FILLER_0_11_78/a_124_375# 0.001597f
C1715 net41 _408_/a_728_93# 0.058816f
C1716 net47 net14 0.033547f
C1717 _086_ _056_ 0.043494f
C1718 _437_/a_1308_423# net14 0.085815f
C1719 _448_/a_2248_156# vss 0.003807f
C1720 _448_/a_2665_112# vdd 0.005876f
C1721 _119_ _313_/a_255_603# 0.001151f
C1722 net53 net23 0.501857f
C1723 net16 net72 0.367221f
C1724 net79 _417_/a_36_151# 0.082646f
C1725 _255_/a_224_552# vdd 0.082462f
C1726 _176_ FILLER_0_15_72/a_484_472# 0.00753f
C1727 _152_ _058_ 0.00259f
C1728 FILLER_0_14_107/a_1380_472# vdd 0.002511f
C1729 net58 vdd 0.929215f
C1730 _115_ FILLER_0_10_94/a_572_375# 0.00887f
C1731 FILLER_0_22_177/a_932_472# vss -0.001894f
C1732 FILLER_0_22_177/a_1380_472# vdd 0.007188f
C1733 _114_ _267_/a_36_472# 0.011923f
C1734 net20 result[9] 1.593573f
C1735 FILLER_0_19_125/a_124_375# net73 0.005414f
C1736 _079_ net76 2.404004f
C1737 FILLER_0_12_136/a_1020_375# FILLER_0_11_142/a_484_472# 0.001543f
C1738 _043_ FILLER_0_13_80/a_36_472# 0.016194f
C1739 _119_ _056_ 0.008929f
C1740 FILLER_0_22_177/a_572_375# _435_/a_36_151# 0.059049f
C1741 cal_itt\[3\] FILLER_0_5_198/a_36_472# 0.07099f
C1742 mask\[3\] net56 0.002632f
C1743 net66 FILLER_0_5_54/a_932_472# 0.001419f
C1744 FILLER_0_12_136/a_572_375# cal_count\[3\] 0.005006f
C1745 _423_/a_36_151# FILLER_0_23_44/a_484_472# 0.001723f
C1746 FILLER_0_3_221/a_1380_472# vss 0.002804f
C1747 FILLER_0_18_2/a_3172_472# FILLER_0_19_28/a_124_375# 0.001684f
C1748 net36 FILLER_0_15_212/a_1380_472# 0.006416f
C1749 _068_ _311_/a_66_473# 0.071325f
C1750 _394_/a_728_93# _175_ 0.010801f
C1751 FILLER_0_15_116/a_36_472# net36 0.013546f
C1752 _427_/a_796_472# _095_ 0.007281f
C1753 _297_/a_36_472# vdd 0.042391f
C1754 _255_/a_224_552# FILLER_0_6_177/a_572_375# 0.001776f
C1755 _008_ vdd 0.284571f
C1756 _334_/a_36_160# FILLER_0_17_104/a_1380_472# 0.004111f
C1757 _070_ _313_/a_67_603# 0.004265f
C1758 net9 cal_itt\[0\] 0.110446f
C1759 _216_/a_67_603# FILLER_0_18_61/a_124_375# 0.014522f
C1760 _451_/a_1040_527# vdd 0.004038f
C1761 FILLER_0_5_54/a_484_472# trim_mask\[1\] 0.013584f
C1762 _093_ _438_/a_2248_156# 0.004221f
C1763 FILLER_0_12_136/a_1380_472# _071_ 0.004003f
C1764 net61 _419_/a_448_472# 0.024246f
C1765 trim[4] net40 0.017911f
C1766 net79 FILLER_0_15_282/a_572_375# 0.01043f
C1767 net57 _116_ 0.069858f
C1768 net50 _036_ 0.002727f
C1769 _374_/a_36_68# _076_ 0.026674f
C1770 FILLER_0_16_89/a_36_472# _040_ 0.015634f
C1771 output47/a_224_472# net55 0.160037f
C1772 FILLER_0_11_124/a_124_375# _120_ 0.012164f
C1773 output47/a_224_472# _452_/a_3129_107# 0.018181f
C1774 net62 _285_/a_36_472# 0.001288f
C1775 net63 net21 0.278824f
C1776 _048_ vss 0.056146f
C1777 mask\[1\] FILLER_0_15_228/a_36_472# 0.02055f
C1778 FILLER_0_5_128/a_124_375# vdd 0.008803f
C1779 _411_/a_2560_156# net75 0.007047f
C1780 FILLER_0_4_49/a_124_375# trim_val\[1\] 0.024557f
C1781 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_572_375# 0.007947f
C1782 _069_ _176_ 0.766885f
C1783 net27 FILLER_0_9_282/a_124_375# 0.003572f
C1784 FILLER_0_18_177/a_484_472# vss -0.001894f
C1785 FILLER_0_18_177/a_932_472# vdd 0.029926f
C1786 _140_ vdd 0.598538f
C1787 _115_ _322_/a_692_472# 0.00171f
C1788 ctlp[1] net33 0.11288f
C1789 mask\[0\] _283_/a_36_472# 0.004645f
C1790 net16 _424_/a_36_151# 0.002969f
C1791 ctln[4] net10 0.1323f
C1792 _411_/a_1000_472# ctln[1] 0.040782f
C1793 mask\[5\] FILLER_0_20_193/a_124_375# 0.015793f
C1794 net58 net75 0.061787f
C1795 trimb[2] net17 0.007637f
C1796 output32/a_224_472# _006_ 0.001009f
C1797 _136_ _337_/a_665_69# 0.001794f
C1798 _058_ net21 0.004383f
C1799 ctln[4] FILLER_0_0_232/a_124_375# 0.002726f
C1800 net16 _447_/a_448_472# 0.063057f
C1801 _105_ _011_ 0.003998f
C1802 FILLER_0_16_57/a_1020_375# vdd 0.004428f
C1803 FILLER_0_16_57/a_572_375# vss 0.00372f
C1804 _440_/a_36_151# FILLER_0_6_47/a_2724_472# 0.001653f
C1805 _439_/a_1308_423# FILLER_0_6_47/a_3260_375# 0.001224f
C1806 net60 result[3] 0.001124f
C1807 _383_/a_36_472# trim_mask\[3\] 0.003193f
C1808 _089_ FILLER_0_5_198/a_36_472# 0.001314f
C1809 FILLER_0_21_150/a_124_375# vss 0.013882f
C1810 FILLER_0_21_150/a_36_472# vdd 0.092128f
C1811 output21/a_224_472# net21 0.011791f
C1812 _002_ _088_ 0.003969f
C1813 _086_ _363_/a_36_68# 0.007567f
C1814 _186_ _407_/a_244_68# 0.001153f
C1815 FILLER_0_5_198/a_572_375# net21 0.023563f
C1816 _066_ _386_/a_124_24# 0.059053f
C1817 net71 vss 0.335256f
C1818 _065_ _441_/a_36_151# 0.00701f
C1819 _070_ _058_ 0.07307f
C1820 net53 _427_/a_2560_156# 0.004594f
C1821 FILLER_0_4_123/a_36_472# FILLER_0_2_111/a_1468_375# 0.00189f
C1822 _015_ FILLER_0_8_247/a_36_472# 0.005458f
C1823 FILLER_0_17_56/a_572_375# FILLER_0_15_59/a_36_472# 0.001188f
C1824 _070_ _315_/a_36_68# 0.031892f
C1825 output39/a_224_472# net39 0.129913f
C1826 _286_/a_224_472# _094_ 0.008468f
C1827 net80 _147_ 0.022618f
C1828 mask\[0\] FILLER_0_14_235/a_124_375# 0.009674f
C1829 _256_/a_1612_497# net4 0.002497f
C1830 FILLER_0_18_2/a_2364_375# vdd 0.002983f
C1831 net47 FILLER_0_5_136/a_124_375# 0.010674f
C1832 FILLER_0_24_290/a_124_375# vss 0.034103f
C1833 FILLER_0_24_290/a_36_472# vdd 0.089567f
C1834 _016_ _427_/a_36_151# 0.00483f
C1835 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_484_472# 0.026657f
C1836 FILLER_0_5_172/a_124_375# vdd 0.028449f
C1837 FILLER_0_6_239/a_36_472# _316_/a_124_24# 0.002228f
C1838 FILLER_0_20_87/a_36_472# _438_/a_1308_423# 0.010224f
C1839 _426_/a_36_151# FILLER_0_9_270/a_36_472# 0.008172f
C1840 _077_ vss 1.071923f
C1841 _323_/a_36_113# _426_/a_2248_156# 0.001661f
C1842 _015_ _426_/a_448_472# 0.035938f
C1843 net16 cal_count\[0\] 0.152321f
C1844 trim_mask\[2\] FILLER_0_2_93/a_484_472# 0.001424f
C1845 FILLER_0_10_78/a_124_375# vdd -0.011193f
C1846 _128_ vdd 0.217501f
C1847 FILLER_0_21_142/a_484_472# net54 0.038728f
C1848 _098_ _437_/a_1308_423# 0.005568f
C1849 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_124_375# 0.016748f
C1850 net65 FILLER_0_3_172/a_1916_375# 0.003745f
C1851 _413_/a_448_472# net76 0.029504f
C1852 output25/a_224_472# net24 0.002325f
C1853 _402_/a_1948_68# _401_/a_36_68# 0.012664f
C1854 FILLER_0_7_104/a_1468_375# _131_ 0.029718f
C1855 net80 _435_/a_448_472# 0.005274f
C1856 net41 FILLER_0_17_38/a_124_375# 0.001109f
C1857 FILLER_0_5_181/a_36_472# net37 0.010376f
C1858 net36 _438_/a_796_472# 0.016855f
C1859 output36/a_224_472# _006_ 0.022685f
C1860 _386_/a_124_24# net37 0.00431f
C1861 output28/a_224_472# net19 0.101711f
C1862 _067_ _043_ 0.189767f
C1863 result[8] _108_ 0.007884f
C1864 _144_ FILLER_0_18_107/a_1828_472# 0.001169f
C1865 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_124_375# 0.009654f
C1866 FILLER_0_16_57/a_1020_375# net72 0.002937f
C1867 _126_ _320_/a_36_472# 0.026216f
C1868 _412_/a_2248_156# net65 0.039861f
C1869 FILLER_0_11_142/a_124_375# vss 0.008766f
C1870 FILLER_0_11_142/a_572_375# vdd 0.014107f
C1871 _149_ vdd 0.379674f
C1872 FILLER_0_18_2/a_36_472# trimb[4] 0.001673f
C1873 ctln[4] FILLER_0_1_212/a_36_472# 0.006408f
C1874 FILLER_0_10_78/a_36_472# FILLER_0_9_72/a_572_375# 0.001543f
C1875 _432_/a_36_151# _136_ 0.004543f
C1876 _015_ FILLER_0_8_239/a_36_472# 0.002627f
C1877 _013_ vss 0.163674f
C1878 _326_/a_36_160# _058_ 0.003897f
C1879 FILLER_0_16_89/a_1020_375# _131_ 0.015706f
C1880 net81 FILLER_0_14_235/a_36_472# 0.002571f
C1881 _088_ _078_ 0.047558f
C1882 _079_ _083_ 0.872842f
C1883 FILLER_0_12_236/a_124_375# vdd 0.005169f
C1884 cal_count\[3\] net17 0.068527f
C1885 _114_ _113_ 0.201729f
C1886 net33 _204_/a_67_603# 0.022193f
C1887 net82 FILLER_0_3_221/a_1020_375# 0.010208f
C1888 _074_ FILLER_0_6_231/a_572_375# 0.009029f
C1889 output47/a_224_472# FILLER_0_15_10/a_36_472# 0.038484f
C1890 FILLER_0_3_172/a_1916_375# net59 0.001221f
C1891 FILLER_0_4_177/a_36_472# FILLER_0_2_177/a_124_375# 0.001512f
C1892 _444_/a_2665_112# FILLER_0_8_37/a_484_472# 0.001167f
C1893 FILLER_0_7_146/a_36_472# _133_ 0.009796f
C1894 FILLER_0_7_146/a_124_375# _076_ 0.00688f
C1895 FILLER_0_10_78/a_36_472# cal_count\[3\] 0.266339f
C1896 _066_ vss 0.08113f
C1897 _093_ _277_/a_36_160# 0.018101f
C1898 _085_ _267_/a_36_472# 0.034055f
C1899 _006_ vdd 0.632993f
C1900 net36 _196_/a_36_160# 0.024527f
C1901 FILLER_0_1_192/a_36_472# vss 0.004422f
C1902 _094_ _195_/a_67_603# 0.043278f
C1903 net44 _054_ 0.003562f
C1904 _132_ _098_ 0.038463f
C1905 _408_/a_728_93# cal_count\[2\] 0.001568f
C1906 _140_ _024_ 0.00287f
C1907 net57 _225_/a_36_160# 0.022745f
C1908 net48 calibrate 0.482314f
C1909 _412_/a_2248_156# net59 0.008792f
C1910 _062_ _163_ 0.001206f
C1911 trim[0] vss 0.132654f
C1912 _094_ net30 0.188507f
C1913 _405_/a_67_603# _184_ 0.010046f
C1914 vdd output40/a_224_472# 0.079607f
C1915 _162_ calibrate 0.228839f
C1916 FILLER_0_21_28/a_3260_375# vdd -0.001166f
C1917 FILLER_0_3_172/a_2276_472# vdd 0.00806f
C1918 fanout71/a_36_113# vss 0.007654f
C1919 net79 _418_/a_36_151# 0.059124f
C1920 _414_/a_1204_472# _053_ 0.003935f
C1921 net73 _093_ 0.350073f
C1922 FILLER_0_8_2/a_124_375# vss 0.003001f
C1923 FILLER_0_8_2/a_36_472# vdd 0.104141f
C1924 net17 net40 1.095167f
C1925 fanout57/a_36_113# vdd 0.005473f
C1926 _427_/a_796_472# net74 0.020124f
C1927 net4 FILLER_0_3_221/a_1380_472# 0.003953f
C1928 cal_itt\[0\] _084_ 0.061227f
C1929 net81 FILLER_0_8_263/a_124_375# 0.026195f
C1930 net37 vss 0.666835f
C1931 _114_ _118_ 0.074399f
C1932 FILLER_0_22_177/a_36_472# net33 0.013661f
C1933 net68 _453_/a_36_151# 0.039234f
C1934 _282_/a_36_160# _098_ 0.00388f
C1935 net57 FILLER_0_16_154/a_1468_375# 0.217874f
C1936 net15 FILLER_0_15_72/a_124_375# 0.006566f
C1937 _414_/a_36_151# FILLER_0_6_177/a_484_472# 0.006095f
C1938 output15/a_224_472# net50 0.00515f
C1939 ctln[8] fanout50/a_36_160# 0.004838f
C1940 net69 net49 0.051235f
C1941 _157_ vss 0.039512f
C1942 _091_ FILLER_0_12_220/a_36_472# 0.003655f
C1943 _255_/a_224_552# _374_/a_36_68# 0.00191f
C1944 net16 _407_/a_36_472# 0.027354f
C1945 FILLER_0_17_72/a_572_375# _131_ 0.006224f
C1946 _442_/a_1000_472# _031_ 0.004174f
C1947 FILLER_0_17_64/a_124_375# vdd 0.027957f
C1948 FILLER_0_16_255/a_36_472# _102_ 0.004641f
C1949 _432_/a_2665_112# _337_/a_49_472# 0.001051f
C1950 _155_ FILLER_0_6_90/a_484_472# 0.005297f
C1951 net20 _122_ 0.046817f
C1952 net68 net69 0.053856f
C1953 result[9] vss 0.348416f
C1954 result[6] FILLER_0_21_286/a_572_375# 0.015047f
C1955 FILLER_0_3_142/a_36_472# trim_mask\[4\] 0.008297f
C1956 FILLER_0_5_72/a_1020_375# net47 0.006974f
C1957 net20 net61 0.014444f
C1958 _059_ FILLER_0_5_136/a_36_472# 0.001755f
C1959 net19 calibrate 0.043159f
C1960 ctlp[2] _109_ 0.059999f
C1961 _053_ net15 0.041871f
C1962 FILLER_0_8_37/a_484_472# _160_ 0.001767f
C1963 fanout61/a_36_113# FILLER_0_21_286/a_572_375# 0.015816f
C1964 _161_ _056_ 0.065732f
C1965 FILLER_0_16_107/a_572_375# _131_ 0.015859f
C1966 net32 output19/a_224_472# 0.101682f
C1967 _127_ net23 0.069001f
C1968 _009_ net77 0.001183f
C1969 FILLER_0_21_133/a_124_375# _098_ 0.006462f
C1970 FILLER_0_20_177/a_124_375# _434_/a_36_151# 0.059049f
C1971 net80 FILLER_0_17_161/a_36_472# 0.003342f
C1972 _077_ FILLER_0_11_64/a_124_375# 0.013507f
C1973 FILLER_0_10_214/a_36_472# _246_/a_36_68# 0.001844f
C1974 FILLER_0_0_266/a_36_472# vdd 0.05043f
C1975 FILLER_0_0_266/a_124_375# vss 0.007654f
C1976 FILLER_0_10_78/a_1468_375# _389_/a_36_148# 0.001699f
C1977 net38 net55 0.10956f
C1978 _042_ _039_ 0.003075f
C1979 net38 _452_/a_3129_107# 0.005269f
C1980 net63 FILLER_0_22_177/a_484_472# 0.059367f
C1981 _430_/a_448_472# _019_ 0.019666f
C1982 mask\[3\] net64 0.002654f
C1983 FILLER_0_3_78/a_124_375# vdd 0.002419f
C1984 FILLER_0_12_136/a_1380_472# net23 0.011488f
C1985 _179_ vss 0.089947f
C1986 _452_/a_36_151# net40 0.012138f
C1987 net16 _444_/a_1308_423# 0.002172f
C1988 FILLER_0_13_228/a_124_375# vdd -0.007362f
C1989 net70 _131_ 0.57653f
C1990 _405_/a_67_603# net47 0.004116f
C1991 cal_count\[3\] FILLER_0_12_28/a_124_375# 0.013328f
C1992 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_124_375# 0.001597f
C1993 _137_ _333_/a_36_160# 0.022811f
C1994 FILLER_0_2_101/a_124_375# vdd 0.044073f
C1995 FILLER_0_4_107/a_1020_375# vdd 0.025121f
C1996 _077_ _439_/a_1000_472# 0.030609f
C1997 _103_ _418_/a_2560_156# 0.002179f
C1998 _360_/a_36_160# FILLER_0_5_117/a_124_375# 0.004736f
C1999 net2 en 0.067828f
C2000 fanout78/a_36_113# net77 0.036366f
C2001 _009_ FILLER_0_23_290/a_36_472# 0.002345f
C2002 trimb[1] FILLER_0_20_15/a_36_472# 0.001292f
C2003 _435_/a_36_151# vdd 0.059103f
C2004 FILLER_0_19_111/a_124_375# net14 0.001837f
C2005 FILLER_0_12_20/a_124_375# net17 0.002167f
C2006 _013_ _424_/a_448_472# 0.043803f
C2007 FILLER_0_9_72/a_572_375# _439_/a_36_151# 0.059049f
C2008 _114_ _068_ 1.097353f
C2009 _091_ mask\[2\] 2.252217f
C2010 FILLER_0_7_195/a_124_375# _062_ 0.001983f
C2011 output19/a_224_472# _422_/a_2248_156# 0.011418f
C2012 ctlp[2] _422_/a_448_472# 0.011383f
C2013 _093_ _143_ 0.003295f
C2014 _071_ net23 0.027895f
C2015 _093_ FILLER_0_17_72/a_2276_472# 0.017114f
C2016 net72 FILLER_0_17_64/a_124_375# 0.002236f
C2017 vss FILLER_0_5_148/a_484_472# 0.009015f
C2018 _412_/a_448_472# en 0.011052f
C2019 _063_ vdd 0.201806f
C2020 FILLER_0_24_96/a_124_375# output24/a_224_472# 0.00363f
C2021 output31/a_224_472# FILLER_0_17_282/a_36_472# 0.008834f
C2022 _079_ FILLER_0_6_231/a_484_472# 0.008159f
C2023 FILLER_0_21_28/a_1468_375# _423_/a_36_151# 0.001543f
C2024 vdd FILLER_0_21_60/a_124_375# 0.014029f
C2025 fanout75/a_36_113# _081_ 0.015843f
C2026 fanout70/a_36_113# net36 0.007807f
C2027 net63 FILLER_0_18_177/a_36_472# 0.015187f
C2028 fanout62/a_36_160# FILLER_0_9_290/a_36_472# 0.001961f
C2029 _053_ _133_ 0.288819f
C2030 _077_ net4 0.656292f
C2031 _021_ _432_/a_36_151# 0.033849f
C2032 FILLER_0_19_47/a_124_375# _182_ 0.001771f
C2033 _139_ vdd 0.085044f
C2034 cal en 0.482495f
C2035 _164_ FILLER_0_6_37/a_36_472# 0.001049f
C2036 _052_ net36 0.005689f
C2037 net20 FILLER_0_13_212/a_932_472# 0.003007f
C2038 FILLER_0_12_28/a_124_375# net40 0.047331f
C2039 _005_ net18 0.073455f
C2040 net16 _404_/a_36_472# 0.001126f
C2041 mask\[5\] _292_/a_36_160# 0.007486f
C2042 net20 _288_/a_224_472# 0.003019f
C2043 net67 FILLER_0_6_37/a_124_375# 0.002918f
C2044 _053_ _376_/a_36_160# 0.005109f
C2045 FILLER_0_7_72/a_3172_472# vss 0.002425f
C2046 _176_ FILLER_0_11_101/a_484_472# 0.001777f
C2047 _236_/a_36_160# net67 0.009332f
C2048 _428_/a_1204_472# _017_ 0.005148f
C2049 _085_ _113_ 0.084246f
C2050 FILLER_0_21_28/a_3260_375# _424_/a_36_151# 0.035849f
C2051 FILLER_0_19_155/a_36_472# vss 0.004125f
C2052 FILLER_0_19_155/a_484_472# vdd 0.003341f
C2053 _235_/a_67_603# net40 0.001273f
C2054 _132_ _131_ 0.444097f
C2055 _140_ _433_/a_36_151# 0.020943f
C2056 FILLER_0_5_54/a_1468_375# net47 0.005049f
C2057 cal_count\[3\] _039_ 0.004827f
C2058 net14 FILLER_0_4_91/a_36_472# 0.005793f
C2059 FILLER_0_0_198/a_36_472# vss 0.00344f
C2060 net82 FILLER_0_3_172/a_3260_375# 0.007693f
C2061 en_co_clk vss 0.014954f
C2062 net68 _165_ 0.002748f
C2063 net73 FILLER_0_17_142/a_36_472# 0.002925f
C2064 FILLER_0_12_136/a_572_375# _120_ 0.001584f
C2065 _158_ vdd 0.131365f
C2066 ctlp[1] net18 0.088706f
C2067 _110_ vss 0.131865f
C2068 net18 _419_/a_796_472# 0.006586f
C2069 _137_ FILLER_0_16_154/a_36_472# 0.005011f
C2070 trim_mask\[2\] _157_ 0.002951f
C2071 trimb[2] trimb[3] 0.369908f
C2072 FILLER_0_5_164/a_572_375# net22 0.002238f
C2073 net64 FILLER_0_11_282/a_36_472# 0.003938f
C2074 net20 output31/a_224_472# 0.004424f
C2075 _376_/a_36_160# FILLER_0_5_88/a_36_472# 0.001448f
C2076 FILLER_0_17_200/a_484_472# vdd 0.008335f
C2077 _253_/a_36_68# _074_ 0.026327f
C2078 _093_ FILLER_0_19_142/a_124_375# 0.00346f
C2079 _075_ net21 0.012335f
C2080 FILLER_0_16_73/a_572_375# _040_ 0.014453f
C2081 _126_ FILLER_0_13_100/a_124_375# 0.00134f
C2082 _414_/a_36_151# _055_ 0.001987f
C2083 mask\[9\] FILLER_0_20_87/a_124_375# 0.004793f
C2084 FILLER_0_15_150/a_124_375# _427_/a_448_472# 0.008952f
C2085 _072_ _126_ 0.012566f
C2086 FILLER_0_19_55/a_124_375# _052_ 0.053626f
C2087 _122_ FILLER_0_5_181/a_36_472# 0.003016f
C2088 net39 net40 0.279259f
C2089 _028_ net15 0.223301f
C2090 output30/a_224_472# result[3] 0.019025f
C2091 _359_/a_1044_488# net74 0.005311f
C2092 result[0] FILLER_0_9_282/a_124_375# 0.00283f
C2093 _007_ vdd 0.129966f
C2094 net33 _023_ 0.015172f
C2095 net64 FILLER_0_14_235/a_36_472# 0.067888f
C2096 net62 _429_/a_448_472# 0.002713f
C2097 _136_ _172_ 0.024344f
C2098 _423_/a_1308_423# vdd 0.00335f
C2099 _423_/a_448_472# vss 0.002481f
C2100 _039_ net40 0.036781f
C2101 mask\[9\] net36 1.116767f
C2102 net73 FILLER_0_19_125/a_36_472# 0.004017f
C2103 net38 FILLER_0_15_10/a_36_472# 0.020589f
C2104 vdd net14 2.23064f
C2105 _316_/a_1084_68# net37 0.001574f
C2106 _075_ _070_ 0.009314f
C2107 _365_/a_244_472# net14 0.001257f
C2108 FILLER_0_17_72/a_932_472# net36 0.00356f
C2109 _106_ net31 0.035117f
C2110 _095_ _041_ 0.002104f
C2111 FILLER_0_17_161/a_124_375# vdd 0.014253f
C2112 _182_ _180_ 0.090106f
C2113 _129_ _059_ 0.005414f
C2114 net4 net37 0.021795f
C2115 net13 vss 0.071697f
C2116 FILLER_0_22_128/a_2812_375# vss 0.004347f
C2117 FILLER_0_22_128/a_3260_375# vdd 0.005207f
C2118 result[8] _435_/a_2665_112# 0.001855f
C2119 FILLER_0_20_107/a_36_472# vss 0.004557f
C2120 _424_/a_2248_156# vdd -0.005751f
C2121 _095_ FILLER_0_14_123/a_36_472# 0.014431f
C2122 _024_ _435_/a_36_151# 0.10993f
C2123 _070_ _172_ 0.237178f
C2124 _190_/a_36_160# net47 0.001489f
C2125 result[6] _420_/a_448_472# 0.017262f
C2126 _098_ FILLER_0_19_111/a_124_375# 0.001331f
C2127 mask\[5\] FILLER_0_20_177/a_484_472# 0.016114f
C2128 net55 _452_/a_3129_107# 0.006395f
C2129 _053_ FILLER_0_6_47/a_2364_375# 0.007053f
C2130 mask\[3\] FILLER_0_18_177/a_1828_472# 0.004274f
C2131 _447_/a_2248_156# vss 0.003961f
C2132 _447_/a_2665_112# vdd 0.022038f
C2133 net23 FILLER_0_5_148/a_572_375# 0.039975f
C2134 FILLER_0_18_107/a_124_375# _438_/a_2665_112# 0.029834f
C2135 net82 vdd 1.014512f
C2136 _320_/a_224_472# _113_ 0.00871f
C2137 _176_ _038_ 0.039948f
C2138 _051_ _098_ 0.006332f
C2139 net50 FILLER_0_9_60/a_36_472# 0.001914f
C2140 FILLER_0_13_142/a_1380_472# _225_/a_36_160# 0.004111f
C2141 net63 FILLER_0_19_187/a_484_472# 0.020823f
C2142 FILLER_0_10_78/a_572_375# _115_ 0.004573f
C2143 _439_/a_2560_156# vss 0.001309f
C2144 FILLER_0_8_138/a_124_375# _120_ 0.12254f
C2145 FILLER_0_8_263/a_124_375# net64 0.004793f
C2146 _445_/a_448_472# net17 0.038794f
C2147 FILLER_0_9_28/a_36_472# net17 0.012954f
C2148 net3 vdd 0.118499f
C2149 FILLER_0_15_116/a_572_375# net70 0.050592f
C2150 net17 trim[3] 0.001664f
C2151 _181_ _402_/a_2172_497# 0.001555f
C2152 mask\[5\] FILLER_0_18_177/a_124_375# 0.002726f
C2153 _431_/a_36_151# FILLER_0_17_133/a_124_375# 0.059049f
C2154 mask\[2\] FILLER_0_15_212/a_484_472# 0.001641f
C2155 net1 _001_ 0.300335f
C2156 _028_ _133_ 0.007084f
C2157 ctln[2] net8 0.057281f
C2158 trim_val\[4\] FILLER_0_3_172/a_932_472# 0.001407f
C2159 FILLER_0_10_37/a_36_472# _453_/a_36_151# 0.003462f
C2160 FILLER_0_7_195/a_36_472# _074_ 0.008706f
C2161 _141_ FILLER_0_21_150/a_124_375# 0.02192f
C2162 _176_ _076_ 0.046873f
C2163 net23 FILLER_0_19_155/a_124_375# 0.001347f
C2164 trimb[1] cal_count\[2\] 0.003178f
C2165 _070_ FILLER_0_5_164/a_484_472# 0.003424f
C2166 _122_ vss 0.750387f
C2167 _091_ net20 0.0557f
C2168 result[6] _421_/a_796_472# 0.004697f
C2169 _091_ _339_/a_36_160# 0.031941f
C2170 _008_ _099_ 0.006163f
C2171 _028_ _376_/a_36_160# 0.026437f
C2172 _132_ _126_ 0.247838f
C2173 result[6] fanout77/a_36_113# 0.001469f
C2174 net61 vss 0.254538f
C2175 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_124_375# 0.012552f
C2176 net50 FILLER_0_2_93/a_124_375# 0.007132f
C2177 net52 FILLER_0_2_93/a_36_472# 0.009026f
C2178 _412_/a_36_151# _001_ 0.006762f
C2179 FILLER_0_12_20/a_124_375# _039_ 0.004669f
C2180 net35 _435_/a_2248_156# 0.001854f
C2181 _159_ _370_/a_124_24# 0.021983f
C2182 mask\[5\] FILLER_0_19_171/a_1380_472# 0.007596f
C2183 _144_ _146_ 0.333799f
C2184 ctlp[2] _300_/a_224_472# 0.002954f
C2185 _188_ net51 0.044278f
C2186 _083_ _260_/a_244_472# 0.00134f
C2187 FILLER_0_5_109/a_36_472# _363_/a_36_68# 0.001024f
C2188 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_572_375# 0.086635f
C2189 output31/a_224_472# _289_/a_36_472# 0.00101f
C2190 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001723f
C2191 input1/a_36_113# vss 0.05331f
C2192 _251_/a_906_472# _068_ 0.001762f
C2193 FILLER_0_4_107/a_124_375# _154_ 0.00183f
C2194 FILLER_0_19_142/a_36_472# _145_ 0.010377f
C2195 _430_/a_36_151# FILLER_0_17_200/a_124_375# 0.059049f
C2196 _341_/a_49_472# mask\[3\] 0.00631f
C2197 net75 net82 0.214597f
C2198 _049_ vss 0.026036f
C2199 _412_/a_36_151# output37/a_224_472# 0.006358f
C2200 fanout54/a_36_160# vss 0.061573f
C2201 _310_/a_49_472# _113_ 0.020387f
C2202 _153_ _365_/a_36_68# 0.056496f
C2203 net35 net25 0.129685f
C2204 FILLER_0_13_65/a_36_472# _043_ 0.013651f
C2205 FILLER_0_4_197/a_1020_375# net22 0.040565f
C2206 _426_/a_2248_156# FILLER_0_8_239/a_124_375# 0.001068f
C2207 _072_ _267_/a_224_472# 0.004269f
C2208 net17 FILLER_0_20_15/a_1020_375# 0.039975f
C2209 _132_ FILLER_0_15_116/a_572_375# 0.003964f
C2210 _061_ vss 0.046487f
C2211 FILLER_0_17_142/a_36_472# FILLER_0_19_142/a_124_375# 0.001512f
C2212 FILLER_0_10_78/a_36_472# _120_ 0.004669f
C2213 FILLER_0_15_205/a_124_375# vdd 0.015886f
C2214 FILLER_0_5_136/a_124_375# vdd 0.035814f
C2215 trim_val\[1\] _034_ 0.001535f
C2216 _424_/a_36_151# _423_/a_1308_423# 0.001722f
C2217 _135_ _134_ 0.038135f
C2218 FILLER_0_5_198/a_124_375# net37 0.009149f
C2219 output27/a_224_472# fanout64/a_36_160# 0.027335f
C2220 FILLER_0_19_125/a_124_375# _334_/a_36_160# 0.001633f
C2221 FILLER_0_14_263/a_124_375# net30 0.016642f
C2222 _098_ vdd 2.272938f
C2223 _408_/a_728_93# _402_/a_56_567# 0.001359f
C2224 _322_/a_1084_68# _129_ 0.00419f
C2225 FILLER_0_17_226/a_124_375# vdd 0.026497f
C2226 _086_ FILLER_0_4_177/a_124_375# 0.024433f
C2227 _429_/a_2665_112# FILLER_0_15_228/a_124_375# 0.001077f
C2228 FILLER_0_17_56/a_572_375# vss 0.05884f
C2229 FILLER_0_17_56/a_36_472# vdd 0.040007f
C2230 FILLER_0_3_54/a_124_375# _160_ 0.004602f
C2231 _414_/a_1204_472# cal_itt\[3\] 0.052432f
C2232 net23 FILLER_0_22_128/a_1916_375# 0.004205f
C2233 net38 _444_/a_1204_472# 0.018432f
C2234 net65 _002_ 0.042811f
C2235 _056_ _246_/a_36_68# 0.017953f
C2236 _277_/a_36_160# _094_ 0.007538f
C2237 _448_/a_36_151# _037_ 0.012725f
C2238 ctln[4] net21 0.009947f
C2239 _413_/a_2560_156# net82 0.00101f
C2240 _269_/a_36_472# _083_ 0.015096f
C2241 FILLER_0_13_212/a_932_472# vss 0.022933f
C2242 net62 FILLER_0_13_212/a_36_472# 0.015187f
C2243 mask\[3\] _103_ 0.055796f
C2244 _436_/a_2665_112# vdd 0.007946f
C2245 _436_/a_2248_156# vss 0.002799f
C2246 _441_/a_36_151# net66 0.057618f
C2247 fanout74/a_36_113# net23 0.005294f
C2248 _308_/a_848_380# _115_ 0.00763f
C2249 net73 FILLER_0_18_139/a_36_472# 0.002491f
C2250 mask\[2\] FILLER_0_15_235/a_484_472# 0.004683f
C2251 _028_ FILLER_0_6_47/a_2364_375# 0.016593f
C2252 _121_ _062_ 0.001616f
C2253 vdd _433_/a_2248_156# 0.008127f
C2254 net76 FILLER_0_5_206/a_36_472# 0.00169f
C2255 _176_ FILLER_0_11_78/a_484_472# 0.008724f
C2256 _395_/a_36_488# _055_ 0.002775f
C2257 FILLER_0_18_139/a_572_375# vdd 0.004039f
C2258 FILLER_0_18_139/a_124_375# vss 0.006869f
C2259 net49 _440_/a_448_472# 0.049861f
C2260 FILLER_0_7_72/a_1020_375# FILLER_0_6_79/a_124_375# 0.026339f
C2261 comp FILLER_0_12_2/a_124_375# 0.007468f
C2262 net50 FILLER_0_6_79/a_36_472# 0.001614f
C2263 FILLER_0_15_116/a_124_375# FILLER_0_14_107/a_1020_375# 0.026339f
C2264 FILLER_0_7_146/a_36_472# net37 0.00208f
C2265 _411_/a_2665_112# ctln[3] 0.003037f
C2266 _394_/a_718_524# cal_count\[1\] 0.009499f
C2267 net68 _440_/a_448_472# 0.02254f
C2268 _132_ FILLER_0_17_104/a_932_472# 0.006091f
C2269 _002_ net59 0.016205f
C2270 _181_ vss 0.003673f
C2271 _239_/a_36_160# net16 0.003137f
C2272 net42 net40 0.007686f
C2273 ctlp[1] _420_/a_1000_472# 0.001106f
C2274 mask\[7\] FILLER_0_22_128/a_2812_375# 0.001476f
C2275 _105_ output19/a_224_472# 0.107668f
C2276 _275_/a_224_472# _092_ 0.002138f
C2277 output31/a_224_472# vss -0.003316f
C2278 _132_ _137_ 0.023462f
C2279 _126_ state\[1\] 1.191746f
C2280 net35 FILLER_0_22_128/a_2276_472# 0.014483f
C2281 _130_ vss 0.090346f
C2282 _178_ _186_ 0.020123f
C2283 _174_ _401_/a_36_68# 0.033989f
C2284 net29 net19 0.305661f
C2285 net36 _451_/a_3129_107# 0.013154f
C2286 net72 FILLER_0_17_56/a_36_472# 0.008058f
C2287 FILLER_0_10_78/a_484_472# _439_/a_36_151# 0.00271f
C2288 _115_ FILLER_0_9_72/a_1468_375# 0.025664f
C2289 _004_ _415_/a_36_151# 0.013592f
C2290 _432_/a_448_472# net63 0.002757f
C2291 net73 FILLER_0_18_107/a_572_375# 0.008889f
C2292 _138_ _043_ 0.005826f
C2293 _139_ _337_/a_49_472# 0.024331f
C2294 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_124_375# 0.003732f
C2295 net68 FILLER_0_6_47/a_36_472# 0.001248f
C2296 net64 FILLER_0_9_282/a_484_472# 0.005717f
C2297 net16 _036_ 0.637538f
C2298 trim_mask\[1\] FILLER_0_6_47/a_932_472# 0.007542f
C2299 _189_/a_255_603# net64 0.002455f
C2300 net39 _445_/a_448_472# 0.014537f
C2301 _372_/a_170_472# _385_/a_36_68# 0.009691f
C2302 FILLER_0_1_266/a_484_472# net8 0.016327f
C2303 net16 _445_/a_2665_112# 0.061595f
C2304 FILLER_0_24_96/a_36_472# output25/a_224_472# 0.010475f
C2305 _053_ _077_ 0.123663f
C2306 FILLER_0_11_101/a_572_375# _070_ 0.011557f
C2307 _052_ FILLER_0_18_37/a_1468_375# 0.001585f
C2308 _444_/a_2665_112# vss 0.002271f
C2309 _444_/a_2560_156# vdd 0.025035f
C2310 FILLER_0_12_220/a_1468_375# _060_ 0.001429f
C2311 FILLER_0_12_220/a_484_472# _090_ 0.006993f
C2312 _155_ FILLER_0_7_104/a_484_472# 0.003068f
C2313 input5/a_36_113# net5 0.061819f
C2314 _021_ FILLER_0_18_171/a_36_472# 0.103755f
C2315 ctlp[1] _421_/a_2248_156# 0.012937f
C2316 _427_/a_2560_156# net23 0.042069f
C2317 calibrate _055_ 0.006584f
C2318 state\[2\] FILLER_0_13_142/a_572_375# 0.007511f
C2319 _072_ _248_/a_36_68# 0.001683f
C2320 fanout53/a_36_160# net53 0.014917f
C2321 net53 FILLER_0_13_142/a_1468_375# 0.002334f
C2322 _425_/a_36_151# _316_/a_124_24# 0.036238f
C2323 FILLER_0_5_72/a_1020_375# vdd 0.009501f
C2324 FILLER_0_5_72/a_572_375# vss 0.006023f
C2325 _446_/a_2248_156# net17 0.008375f
C2326 output11/a_224_472# FILLER_0_0_232/a_36_472# 0.023414f
C2327 _394_/a_728_93# FILLER_0_13_72/a_484_472# 0.018997f
C2328 FILLER_0_15_142/a_572_375# net56 0.001809f
C2329 net61 mask\[7\] 0.071542f
C2330 net80 net57 0.002913f
C2331 _076_ FILLER_0_8_239/a_36_472# 0.029514f
C2332 FILLER_0_16_57/a_1380_472# _394_/a_728_93# 0.001627f
C2333 _057_ _116_ 0.028033f
C2334 FILLER_0_12_236/a_572_375# FILLER_0_14_235/a_484_472# 0.001026f
C2335 FILLER_0_4_91/a_484_472# _160_ 0.009925f
C2336 _432_/a_796_472# _098_ 0.038458f
C2337 _078_ net59 0.168928f
C2338 _070_ _152_ 0.114651f
C2339 _133_ _081_ 0.002847f
C2340 net4 _122_ 0.03487f
C2341 net35 FILLER_0_22_107/a_484_472# 0.008026f
C2342 trim_val\[4\] net23 0.014503f
C2343 _072_ _060_ 0.080908f
C2344 output22/a_224_472# vdd 0.111234f
C2345 _256_/a_36_68# _058_ 0.001402f
C2346 _144_ _147_ 0.057955f
C2347 _417_/a_2248_156# net30 0.048831f
C2348 FILLER_0_16_89/a_932_472# _136_ 0.045229f
C2349 FILLER_0_7_104/a_932_472# _133_ 0.019721f
C2350 _414_/a_2665_112# net22 0.004067f
C2351 _372_/a_3662_472# _062_ 0.0012f
C2352 _408_/a_56_524# net17 0.048018f
C2353 FILLER_0_18_177/a_572_375# FILLER_0_20_177/a_484_472# 0.0027f
C2354 FILLER_0_12_136/a_932_472# _069_ 0.002161f
C2355 FILLER_0_12_136/a_36_472# _126_ 0.014981f
C2356 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_484_472# 0.013277f
C2357 mask\[7\] _049_ 0.234746f
C2358 trim_val\[1\] FILLER_0_6_37/a_124_375# 0.007292f
C2359 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_484_472# 0.001963f
C2360 calibrate _313_/a_67_603# 0.021436f
C2361 _405_/a_67_603# vdd 0.034681f
C2362 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_572_375# 0.001597f
C2363 _436_/a_2665_112# FILLER_0_22_128/a_572_375# 0.001092f
C2364 _436_/a_2560_156# FILLER_0_22_128/a_124_375# 0.001178f
C2365 net1 input4/a_36_68# 0.056389f
C2366 _372_/a_170_472# vdd 0.031606f
C2367 net15 _449_/a_1308_423# 0.015651f
C2368 _094_ _418_/a_2665_112# 0.035668f
C2369 _131_ vdd 1.344823f
C2370 _120_ _039_ 0.148356f
C2371 FILLER_0_4_197/a_1468_375# net22 0.009108f
C2372 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_124_375# 0.012552f
C2373 FILLER_0_8_24/a_124_375# net17 0.039695f
C2374 FILLER_0_10_78/a_1380_472# _114_ 0.011079f
C2375 mask\[3\] _019_ 0.001403f
C2376 _091_ vss 0.56693f
C2377 _411_/a_448_472# net65 0.006279f
C2378 FILLER_0_20_177/a_124_375# mask\[6\] 0.001158f
C2379 result[7] _420_/a_448_472# 0.003274f
C2380 _443_/a_2248_156# _386_/a_124_24# 0.001257f
C2381 FILLER_0_5_128/a_484_472# _163_ 0.009861f
C2382 _136_ net21 0.022198f
C2383 net41 _065_ 0.001765f
C2384 FILLER_0_9_28/a_2276_472# _042_ 0.002496f
C2385 vss _160_ 1.119894f
C2386 _185_ _402_/a_728_93# 0.007151f
C2387 net16 _183_ 0.001103f
C2388 _086_ _133_ 0.035637f
C2389 fanout66/a_36_113# net69 0.001345f
C2390 _154_ _153_ 0.719561f
C2391 FILLER_0_12_20/a_36_472# net6 0.007073f
C2392 _141_ FILLER_0_19_155/a_36_472# 0.05777f
C2393 net7 output16/a_224_472# 0.001321f
C2394 _026_ FILLER_0_20_87/a_36_472# 0.004568f
C2395 _199_/a_36_160# _046_ 0.017122f
C2396 _410_/a_36_68# net51 0.014342f
C2397 net76 _123_ 0.003431f
C2398 _053_ net37 0.080949f
C2399 FILLER_0_24_96/a_124_375# vss 0.017357f
C2400 valid _425_/a_2665_112# 0.001839f
C2401 _165_ FILLER_0_6_47/a_124_375# 0.014312f
C2402 _136_ _070_ 0.010577f
C2403 _119_ _133_ 0.038875f
C2404 _449_/a_448_472# _038_ 0.064169f
C2405 _093_ _334_/a_36_160# 0.014676f
C2406 _058_ _439_/a_2665_112# 0.001029f
C2407 FILLER_0_16_57/a_1020_375# _176_ 0.006334f
C2408 _095_ _184_ 0.265966f
C2409 _136_ _356_/a_36_472# 0.004667f
C2410 _070_ net21 0.03068f
C2411 _267_/a_224_472# state\[1\] 0.001937f
C2412 FILLER_0_18_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001684f
C2413 _326_/a_36_160# FILLER_0_7_104/a_1380_472# 0.002051f
C2414 FILLER_0_15_142/a_36_472# fanout73/a_36_113# 0.009544f
C2415 net34 _419_/a_2665_112# 0.001468f
C2416 FILLER_0_9_270/a_36_472# vss 0.001642f
C2417 FILLER_0_9_270/a_484_472# vdd 0.006354f
C2418 net57 _385_/a_244_472# 0.001506f
C2419 mask\[7\] _436_/a_2248_156# 0.003615f
C2420 FILLER_0_12_20/a_484_472# net40 0.003391f
C2421 FILLER_0_17_72/a_2364_375# _136_ 0.047331f
C2422 FILLER_0_18_171/a_36_472# FILLER_0_18_177/a_36_472# 0.003468f
C2423 FILLER_0_22_128/a_3172_472# _146_ 0.008065f
C2424 _025_ _436_/a_1000_472# 0.061189f
C2425 FILLER_0_12_2/a_572_375# _450_/a_36_151# 0.001597f
C2426 _057_ _117_ 0.120323f
C2427 _428_/a_2665_112# vdd 0.004735f
C2428 _120_ FILLER_0_8_156/a_36_472# 0.005842f
C2429 trim_mask\[4\] _081_ 0.111668f
C2430 FILLER_0_5_54/a_1020_375# vss 0.003196f
C2431 FILLER_0_5_54/a_1468_375# vdd 0.014683f
C2432 trimb[1] FILLER_0_20_2/a_124_375# 0.003431f
C2433 FILLER_0_4_99/a_36_472# net14 0.022408f
C2434 _058_ calibrate 0.075294f
C2435 _170_ _386_/a_124_24# 0.008511f
C2436 FILLER_0_21_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001723f
C2437 net72 _131_ 0.186396f
C2438 clk vdd 0.053789f
C2439 FILLER_0_10_214/a_124_375# _069_ 0.014379f
C2440 result[8] FILLER_0_24_274/a_484_472# 0.005458f
C2441 _077_ _028_ 0.017713f
C2442 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_484_472# 0.013277f
C2443 cal_itt\[1\] net8 0.040042f
C2444 FILLER_0_7_72/a_1020_375# vss 0.004851f
C2445 _095_ FILLER_0_13_100/a_124_375# 0.001989f
C2446 _431_/a_2248_156# net73 0.003228f
C2447 net82 FILLER_0_3_142/a_124_375# 0.018696f
C2448 FILLER_0_5_172/a_124_375# FILLER_0_5_164/a_572_375# 0.012001f
C2449 _074_ _375_/a_1612_497# 0.004567f
C2450 _281_/a_672_472# _098_ 0.002084f
C2451 _122_ FILLER_0_5_198/a_124_375# 0.001352f
C2452 _443_/a_2248_156# vss 0.008696f
C2453 _443_/a_2665_112# vdd 0.011824f
C2454 _128_ _176_ 0.180252f
C2455 FILLER_0_10_78/a_124_375# _176_ 0.002785f
C2456 output36/a_224_472# result[2] 0.002356f
C2457 _308_/a_692_472# _115_ 0.001485f
C2458 _369_/a_244_472# _160_ 0.00146f
C2459 FILLER_0_19_28/a_36_472# net40 0.020968f
C2460 vss FILLER_0_3_212/a_124_375# 0.009048f
C2461 vdd FILLER_0_3_212/a_36_472# 0.110132f
C2462 net58 _082_ 0.004276f
C2463 _431_/a_36_151# _020_ 0.023081f
C2464 _093_ net36 0.214976f
C2465 net20 _420_/a_2248_156# 0.003737f
C2466 net70 _095_ 0.222423f
C2467 FILLER_0_5_72/a_1468_375# _440_/a_2665_112# 0.001077f
C2468 net15 FILLER_0_6_47/a_1468_375# 0.007439f
C2469 FILLER_0_9_223/a_36_472# _068_ 0.076678f
C2470 output22/a_224_472# _024_ 0.029795f
C2471 net8 vss 0.171128f
C2472 net62 net18 0.089041f
C2473 _164_ FILLER_0_6_47/a_932_472# 0.004272f
C2474 _057_ _225_/a_36_160# 0.026341f
C2475 net19 _420_/a_1204_472# 0.001828f
C2476 FILLER_0_15_142/a_572_375# _095_ 0.003935f
C2477 net15 output16/a_224_472# 0.013768f
C2478 _095_ net47 0.508892f
C2479 _116_ cal_count\[3\] 0.384121f
C2480 FILLER_0_16_73/a_124_375# _131_ 0.015859f
C2481 output35/a_224_472# _435_/a_2248_156# 0.019736f
C2482 net44 FILLER_0_8_2/a_36_472# 0.005851f
C2483 FILLER_0_4_144/a_124_375# net47 0.012023f
C2484 _132_ FILLER_0_18_107/a_2276_472# 0.006713f
C2485 output39/a_224_472# net67 0.008957f
C2486 net41 net51 0.031531f
C2487 net16 FILLER_0_18_37/a_932_472# 0.008749f
C2488 _326_/a_36_160# _070_ 0.018037f
C2489 _098_ _433_/a_36_151# 0.023263f
C2490 _126_ vdd 0.682779f
C2491 net17 _450_/a_36_151# 0.006157f
C2492 FILLER_0_9_28/a_3172_472# net51 0.047897f
C2493 _077_ trim_mask\[0\] 0.090587f
C2494 net24 net14 0.172253f
C2495 FILLER_0_9_28/a_36_472# net42 0.038355f
C2496 _150_ vss 0.016993f
C2497 _190_/a_36_160# vdd 0.031799f
C2498 _140_ _434_/a_36_151# 0.025956f
C2499 net15 FILLER_0_9_60/a_484_472# 0.020589f
C2500 net36 FILLER_0_15_180/a_572_375# 0.002531f
C2501 result[2] vdd 0.18482f
C2502 net15 fanout72/a_36_113# 0.010284f
C2503 net74 _370_/a_1084_68# 0.001301f
C2504 FILLER_0_5_164/a_36_472# _066_ 0.00611f
C2505 net61 net79 0.159f
C2506 ctlp[1] _419_/a_1204_472# 0.007338f
C2507 net17 _043_ 0.571818f
C2508 FILLER_0_6_239/a_124_375# _317_/a_36_113# 0.002437f
C2509 FILLER_0_18_2/a_1468_375# net38 0.016983f
C2510 _170_ vss 0.280383f
C2511 _053_ FILLER_0_7_72/a_3172_472# 0.032946f
C2512 result[1] FILLER_0_11_282/a_124_375# 0.018322f
C2513 _056_ FILLER_0_12_196/a_124_375# 0.027077f
C2514 net56 state\[1\] 0.007364f
C2515 _065_ _164_ 0.006953f
C2516 trim_val\[2\] _166_ 0.014514f
C2517 trim_mask\[2\] _160_ 0.367302f
C2518 _005_ _192_/a_255_603# 0.001058f
C2519 _101_ mask\[1\] 0.033941f
C2520 _323_/a_36_113# FILLER_0_10_247/a_124_375# 0.001846f
C2521 net64 FILLER_0_12_220/a_1468_375# 0.01836f
C2522 _434_/a_1000_472# mask\[6\] 0.021582f
C2523 _104_ net19 0.159483f
C2524 _111_ _438_/a_36_151# 0.003619f
C2525 net82 fanout52/a_36_160# 0.026154f
C2526 _185_ net17 0.270086f
C2527 FILLER_0_0_96/a_124_375# trim_mask\[3\] 0.006277f
C2528 _421_/a_2665_112# net19 0.01849f
C2529 _305_/a_36_159# net76 0.010842f
C2530 net16 _408_/a_2215_68# 0.002096f
C2531 result[7] FILLER_0_24_274/a_1380_472# 0.006454f
C2532 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_124_375# 0.012222f
C2533 FILLER_0_15_212/a_932_472# vdd 0.001767f
C2534 net62 FILLER_0_15_212/a_1468_375# 0.001106f
C2535 FILLER_0_18_2/a_3172_472# net17 0.002402f
C2536 FILLER_0_15_116/a_572_375# vdd 0.017636f
C2537 FILLER_0_6_90/a_484_472# net14 0.014785f
C2538 net20 _426_/a_2248_156# 0.007902f
C2539 _058_ _125_ 0.016525f
C2540 _132_ _095_ 0.042874f
C2541 _227_/a_36_160# FILLER_0_8_156/a_36_472# 0.006647f
C2542 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_124_375# 0.012221f
C2543 FILLER_0_24_274/a_1380_472# FILLER_0_23_282/a_484_472# 0.058411f
C2544 result[9] ctlp[2] 0.105977f
C2545 net58 fanout64/a_36_160# 0.002438f
C2546 ctlp[6] output24/a_224_472# 0.004288f
C2547 FILLER_0_5_164/a_36_472# net37 0.008378f
C2548 _141_ _049_ 0.0035f
C2549 result[6] net19 0.834308f
C2550 net53 state\[2\] 0.001982f
C2551 _134_ FILLER_0_10_107/a_572_375# 0.047331f
C2552 net55 _216_/a_255_603# 0.001011f
C2553 _030_ net40 0.002509f
C2554 state\[1\] _060_ 0.003973f
C2555 _188_ _067_ 0.001554f
C2556 FILLER_0_4_91/a_484_472# _156_ 0.009828f
C2557 FILLER_0_10_107/a_124_375# vdd 0.045066f
C2558 _091_ net4 0.125608f
C2559 _420_/a_1204_472# _009_ 0.009314f
C2560 _093_ _432_/a_2248_156# 0.012955f
C2561 _445_/a_1000_472# net40 0.015508f
C2562 net22 _205_/a_36_160# 0.109939f
C2563 _293_/a_36_472# vss 0.014842f
C2564 FILLER_0_4_197/a_124_375# _088_ 0.024641f
C2565 mask\[4\] FILLER_0_18_177/a_2812_375# 0.013557f
C2566 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_36_472# 0.001723f
C2567 trim_mask\[1\] _163_ 0.166315f
C2568 _308_/a_848_380# FILLER_0_9_105/a_36_472# 0.15783f
C2569 cal_count\[3\] _117_ 0.00114f
C2570 FILLER_0_18_177/a_2812_375# net22 0.010501f
C2571 _443_/a_1308_423# net13 0.004098f
C2572 _443_/a_1000_472# net23 0.034596f
C2573 FILLER_0_20_177/a_1020_375# vdd 0.005483f
C2574 net52 _441_/a_2560_156# 0.004721f
C2575 net50 _441_/a_2248_156# 0.027849f
C2576 _440_/a_448_472# net47 0.016997f
C2577 FILLER_0_13_212/a_932_472# net79 0.006824f
C2578 FILLER_0_4_49/a_572_375# net49 0.004345f
C2579 ctln[3] FILLER_0_0_266/a_124_375# 0.002726f
C2580 _333_/a_36_160# _097_ 0.001332f
C2581 _069_ _429_/a_36_151# 0.010076f
C2582 _443_/a_36_151# _442_/a_36_151# 0.06169f
C2583 FILLER_0_4_49/a_572_375# net68 0.023227f
C2584 FILLER_0_18_2/a_3172_472# _452_/a_36_151# 0.059367f
C2585 net22 mask\[6\] 0.612004f
C2586 net74 _372_/a_1194_69# 0.002006f
C2587 net82 _443_/a_448_472# 0.007335f
C2588 net52 _439_/a_2665_112# 0.00117f
C2589 _095_ FILLER_0_14_107/a_572_375# 0.01418f
C2590 _012_ vss 0.454371f
C2591 FILLER_0_17_104/a_932_472# vdd 0.020019f
C2592 _044_ net30 0.005104f
C2593 _050_ FILLER_0_22_107/a_572_375# 0.001825f
C2594 FILLER_0_17_56/a_36_472# _404_/a_36_472# 0.004546f
C2595 FILLER_0_13_290/a_36_472# output30/a_224_472# 0.0323f
C2596 FILLER_0_5_54/a_932_472# FILLER_0_6_47/a_1828_472# 0.026657f
C2597 _425_/a_2248_156# net37 0.01491f
C2598 _371_/a_36_113# _159_ 0.021612f
C2599 _104_ _009_ 0.284256f
C2600 vss _156_ 0.089339f
C2601 result[7] _419_/a_1308_423# 0.015718f
C2602 _131_ _331_/a_448_472# 0.007271f
C2603 _010_ _420_/a_2665_112# 0.029378f
C2604 _136_ _451_/a_448_472# 0.047841f
C2605 cal_count\[2\] _180_ 0.153207f
C2606 _434_/a_796_472# _023_ 0.002118f
C2607 _365_/a_692_472# _156_ 0.001127f
C2608 _071_ FILLER_0_13_142/a_1468_375# 0.007453f
C2609 _267_/a_36_472# vss 0.001495f
C2610 _105_ output18/a_224_472# 0.105478f
C2611 net79 _284_/a_224_472# 0.009327f
C2612 FILLER_0_21_286/a_484_472# net77 0.02147f
C2613 FILLER_0_18_171/a_124_375# vdd 0.021417f
C2614 _137_ vdd 0.945976f
C2615 ctlp[1] FILLER_0_23_282/a_36_472# 0.003169f
C2616 mask\[8\] _437_/a_1308_423# 0.001928f
C2617 net49 FILLER_0_3_78/a_36_472# 0.059367f
C2618 _030_ FILLER_0_3_78/a_484_472# 0.007736f
C2619 _422_/a_1308_423# _009_ 0.008875f
C2620 _453_/a_36_151# vdd 0.164654f
C2621 _031_ FILLER_0_2_111/a_932_472# 0.017509f
C2622 _413_/a_2665_112# net82 0.004306f
C2623 net48 _076_ 0.077031f
C2624 _108_ _107_ 0.018045f
C2625 _173_ _408_/a_728_93# 0.022838f
C2626 _328_/a_36_113# net70 0.00292f
C2627 _077_ cal_itt\[3\] 0.009816f
C2628 _036_ FILLER_0_3_78/a_124_375# 0.00215f
C2629 _429_/a_36_151# FILLER_0_15_212/a_36_472# 0.001723f
C2630 net74 FILLER_0_13_100/a_124_375# 0.005049f
C2631 net36 FILLER_0_18_76/a_572_375# 0.005153f
C2632 _126_ FILLER_0_13_206/a_36_472# 0.026561f
C2633 net54 _050_ 0.040506f
C2634 result[6] _009_ 0.095754f
C2635 FILLER_0_19_171/a_1468_375# vss 0.054352f
C2636 FILLER_0_19_171/a_36_472# vdd 0.004762f
C2637 net34 _146_ 0.004718f
C2638 _091_ FILLER_0_13_212/a_1020_375# 0.00799f
C2639 _162_ _076_ 0.008623f
C2640 net57 fanout56/a_36_113# 0.079542f
C2641 net69 vdd 1.102677f
C2642 net82 FILLER_0_2_177/a_572_375# 0.003837f
C2643 FILLER_0_15_235/a_484_472# vss 0.003614f
C2644 _114_ _311_/a_3220_473# 0.003283f
C2645 net62 FILLER_0_15_235/a_572_375# 0.001315f
C2646 _053_ _122_ 0.368823f
C2647 net78 _421_/a_1308_423# 0.015694f
C2648 FILLER_0_17_282/a_36_472# _418_/a_1308_423# 0.001295f
C2649 _438_/a_448_472# vss 0.00615f
C2650 FILLER_0_7_72/a_3172_472# _028_ 0.001873f
C2651 _213_/a_67_603# _051_ 0.015959f
C2652 _144_ _433_/a_2665_112# 0.030413f
C2653 _099_ _098_ 0.018316f
C2654 net4 FILLER_0_3_212/a_124_375# 0.001739f
C2655 _096_ _090_ 0.026104f
C2656 FILLER_0_17_72/a_2364_375# _451_/a_448_472# 0.001512f
C2657 net70 net74 0.017928f
C2658 net5 rstn 0.101356f
C2659 _069_ _055_ 0.741952f
C2660 net55 FILLER_0_18_61/a_36_472# 0.022296f
C2661 cal_count\[1\] FILLER_0_15_59/a_572_375# 0.008797f
C2662 FILLER_0_14_91/a_484_472# _095_ 0.011772f
C2663 FILLER_0_18_2/a_1468_375# net55 0.007169f
C2664 ctln[1] net19 0.001327f
C2665 FILLER_0_15_142/a_572_375# net74 0.001652f
C2666 net74 net47 0.030815f
C2667 _095_ state\[1\] 0.069906f
C2668 net4 net8 0.00647f
C2669 FILLER_0_15_142/a_36_472# vss 0.006166f
C2670 FILLER_0_10_37/a_124_375# _042_ 0.002437f
C2671 net16 _450_/a_3129_107# 0.064714f
C2672 _428_/a_36_151# _135_ 0.030608f
C2673 _063_ _445_/a_2665_112# 0.009759f
C2674 _450_/a_36_151# _039_ 0.018559f
C2675 net64 _282_/a_36_160# 0.014431f
C2676 _171_ net14 0.020479f
C2677 _132_ mask\[8\] 0.029292f
C2678 FILLER_0_17_64/a_124_375# _183_ 0.001236f
C2679 net57 _311_/a_66_473# 0.013777f
C2680 net18 net33 0.001671f
C2681 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1380_472# 0.013277f
C2682 _067_ FILLER_0_12_20/a_36_472# 0.015608f
C2683 _043_ _039_ 0.001161f
C2684 _114_ _135_ 0.018715f
C2685 _123_ FILLER_0_6_231/a_484_472# 0.001396f
C2686 _086_ _077_ 0.058673f
C2687 ctln[1] input2/a_36_113# 0.05197f
C2688 net72 _453_/a_36_151# 0.001607f
C2689 _328_/a_36_113# _132_ 0.006002f
C2690 _081_ _066_ 0.061358f
C2691 _420_/a_2248_156# vss -0.001f
C2692 _420_/a_2665_112# vdd 0.024431f
C2693 mask\[4\] FILLER_0_19_187/a_572_375# 0.00553f
C2694 _274_/a_244_497# net64 0.004085f
C2695 result[9] _421_/a_1000_472# 0.012144f
C2696 FILLER_0_15_142/a_484_472# vss 0.029611f
C2697 FILLER_0_7_72/a_3172_472# trim_mask\[0\] 0.001438f
C2698 net53 _451_/a_1353_112# 0.028324f
C2699 _115_ FILLER_0_9_105/a_484_472# 0.004075f
C2700 _263_/a_224_472# net59 0.002558f
C2701 _119_ _077_ 2.584241f
C2702 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_484_472# 0.013276f
C2703 _325_/a_224_472# _120_ 0.00233f
C2704 _414_/a_1308_423# _074_ 0.005458f
C2705 _013_ FILLER_0_18_37/a_1380_472# 0.01384f
C2706 net19 _419_/a_2248_156# 0.012726f
C2707 FILLER_0_17_104/a_124_375# net14 0.010099f
C2708 _086_ FILLER_0_11_142/a_124_375# 0.009046f
C2709 FILLER_0_10_214/a_124_375# _090_ 0.072741f
C2710 net44 net3 0.195171f
C2711 mask\[9\] _438_/a_2560_156# 0.008709f
C2712 _093_ FILLER_0_18_139/a_1380_472# 0.007013f
C2713 _236_/a_36_160# trim[1] 0.003604f
C2714 FILLER_0_18_209/a_36_472# _047_ 0.002672f
C2715 FILLER_0_7_146/a_124_375# _372_/a_170_472# 0.001188f
C2716 _176_ net14 0.031922f
C2717 FILLER_0_3_172/a_484_472# net22 0.012284f
C2718 cal_itt\[3\] net37 0.03677f
C2719 _434_/a_2248_156# vdd 0.019386f
C2720 _386_/a_848_380# net22 0.00429f
C2721 _075_ calibrate 0.022901f
C2722 _132_ net74 0.031741f
C2723 net56 vdd 0.277166f
C2724 FILLER_0_13_142/a_484_472# vss 0.024835f
C2725 FILLER_0_4_177/a_484_472# vdd 0.010663f
C2726 FILLER_0_4_177/a_36_472# vss 0.001806f
C2727 output8/a_224_472# _073_ 0.043098f
C2728 _091_ net79 0.052824f
C2729 _417_/a_1308_423# vss 0.002064f
C2730 net62 _417_/a_36_151# 0.044051f
C2731 _424_/a_448_472# _012_ 0.007299f
C2732 FILLER_0_16_57/a_484_472# FILLER_0_15_59/a_124_375# 0.001543f
C2733 FILLER_0_8_127/a_124_375# _133_ 0.001928f
C2734 _081_ net37 1.274337f
C2735 _213_/a_67_603# vdd 0.014901f
C2736 FILLER_0_1_266/a_572_375# rstn 0.00328f
C2737 _095_ _402_/a_718_527# 0.002109f
C2738 FILLER_0_8_24/a_124_375# net42 0.032303f
C2739 _091_ _141_ 0.010074f
C2740 _177_ _451_/a_2225_156# 0.031347f
C2741 net35 FILLER_0_22_177/a_124_375# 0.0073f
C2742 _044_ FILLER_0_14_263/a_36_472# 0.002013f
C2743 FILLER_0_22_86/a_572_375# net71 0.002239f
C2744 _248_/a_36_68# vdd 0.038887f
C2745 net63 _069_ 0.04528f
C2746 ctln[6] FILLER_0_0_130/a_36_472# 0.023355f
C2747 trim_mask\[2\] _156_ 0.018332f
C2748 FILLER_0_8_127/a_36_472# net74 0.063481f
C2749 net44 _245_/a_672_472# 0.001285f
C2750 FILLER_0_3_172/a_124_375# vdd 0.010886f
C2751 FILLER_0_16_107/a_484_472# net36 0.003765f
C2752 _178_ _179_ 0.063494f
C2753 output10/a_224_472# ctln[1] 0.083631f
C2754 _422_/a_1000_472# vdd 0.005284f
C2755 net81 vdd 1.658963f
C2756 _163_ _164_ 0.021311f
C2757 _165_ vdd 0.168803f
C2758 _131_ _404_/a_36_472# 0.031567f
C2759 _412_/a_2248_156# output37/a_224_472# 0.001141f
C2760 net67 net40 0.886781f
C2761 FILLER_0_8_107/a_124_375# _133_ 0.048874f
C2762 _426_/a_2248_156# vss 0.002303f
C2763 _426_/a_2665_112# vdd 0.008893f
C2764 FILLER_0_15_212/a_124_375# FILLER_0_15_205/a_124_375# 0.004426f
C2765 _087_ FILLER_0_5_181/a_36_472# 0.154469f
C2766 _033_ net17 0.028529f
C2767 _265_/a_224_472# net59 0.001052f
C2768 _088_ FILLER_0_3_172/a_2812_375# 0.002239f
C2769 ctlp[5] net23 0.025206f
C2770 FILLER_0_15_282/a_484_472# vss 0.005507f
C2771 net62 FILLER_0_15_282/a_572_375# 0.007699f
C2772 net61 ctlp[2] 0.022612f
C2773 ctlp[1] FILLER_0_24_290/a_124_375# 0.050488f
C2774 _060_ vdd 0.349556f
C2775 _098_ FILLER_0_15_212/a_124_375# 0.008125f
C2776 _113_ vss 0.147905f
C2777 FILLER_0_1_192/a_124_375# net21 0.067765f
C2778 net69 _441_/a_1000_472# 0.018209f
C2779 _304_/a_224_472# mask\[9\] 0.003125f
C2780 _093_ FILLER_0_16_89/a_572_375# 0.002889f
C2781 fanout50/a_36_160# _383_/a_36_472# 0.096296f
C2782 FILLER_0_21_125/a_572_375# _140_ 0.01659f
C2783 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_36_472# 0.086742f
C2784 FILLER_0_4_49/a_484_472# _164_ 0.003258f
C2785 _414_/a_36_151# _003_ 0.021191f
C2786 _069_ _315_/a_36_68# 0.002242f
C2787 _102_ net30 0.043037f
C2788 FILLER_0_16_37/a_36_472# _402_/a_1296_93# 0.001477f
C2789 _447_/a_448_472# net69 0.001694f
C2790 _086_ net37 0.039329f
C2791 ctln[4] FILLER_0_0_198/a_124_375# 0.015879f
C2792 _415_/a_2665_112# fanout62/a_36_160# 0.016426f
C2793 net63 FILLER_0_15_212/a_36_472# 0.059367f
C2794 net49 _029_ 0.004408f
C2795 _122_ FILLER_0_5_164/a_36_472# 0.002232f
C2796 trimb[1] FILLER_0_18_2/a_36_472# 0.010728f
C2797 _089_ net37 0.0326f
C2798 _414_/a_36_151# net21 0.007791f
C2799 net68 _029_ 0.094915f
C2800 _253_/a_36_68# _073_ 0.027664f
C2801 net52 FILLER_0_5_72/a_124_375# 0.029702f
C2802 FILLER_0_4_197/a_1380_472# net76 0.003767f
C2803 net12 vdd 0.082923f
C2804 _053_ _444_/a_2665_112# 0.001698f
C2805 _048_ _204_/a_67_603# 0.004547f
C2806 FILLER_0_20_107/a_124_375# FILLER_0_20_98/a_124_375# 0.003228f
C2807 FILLER_0_2_111/a_572_375# vdd 0.012666f
C2808 FILLER_0_8_24/a_484_472# net40 0.004383f
C2809 FILLER_0_6_79/a_124_375# FILLER_0_6_47/a_3260_375# 0.012001f
C2810 _330_/a_224_472# vdd 0.001701f
C2811 net75 net81 0.420021f
C2812 net20 _256_/a_244_497# 0.005033f
C2813 FILLER_0_12_136/a_1380_472# state\[2\] 0.005779f
C2814 net34 _147_ 0.144404f
C2815 _372_/a_358_69# _163_ 0.001427f
C2816 _116_ _120_ 0.005759f
C2817 result[7] net19 0.087363f
C2818 _428_/a_448_472# _131_ 0.041178f
C2819 _360_/a_36_160# FILLER_0_4_123/a_124_375# 0.013555f
C2820 _081_ FILLER_0_5_148/a_484_472# 0.016132f
C2821 _255_/a_224_552# _162_ 0.010564f
C2822 _057_ _375_/a_36_68# 0.003063f
C2823 _118_ vss 0.217218f
C2824 FILLER_0_7_72/a_36_472# vdd 0.106377f
C2825 _093_ FILLER_0_18_209/a_484_472# 0.014737f
C2826 ctln[8] vss 0.351742f
C2827 net26 FILLER_0_21_28/a_1828_472# 0.010367f
C2828 FILLER_0_18_107/a_2276_472# vdd 0.004405f
C2829 ctln[2] net2 0.004284f
C2830 output8/a_224_472# cal_itt\[2\] 0.05561f
C2831 FILLER_0_2_171/a_36_472# net22 0.081357f
C2832 net41 net66 0.08664f
C2833 FILLER_0_9_28/a_1380_472# net68 0.008573f
C2834 net78 _419_/a_448_472# 0.0122f
C2835 net36 _094_ 0.086414f
C2836 _016_ FILLER_0_12_136/a_572_375# 0.00332f
C2837 _026_ _437_/a_1308_423# 0.018479f
C2838 _149_ _437_/a_1000_472# 0.019115f
C2839 net54 FILLER_0_22_128/a_1828_472# 0.009504f
C2840 net28 _426_/a_36_151# 0.004878f
C2841 net67 FILLER_0_12_20/a_124_375# 0.007044f
C2842 net34 _435_/a_448_472# 0.013341f
C2843 _087_ vss 0.09895f
C2844 _079_ vdd 0.476075f
C2845 FILLER_0_8_107/a_36_472# _062_ 0.001832f
C2846 fanout82/a_36_113# _425_/a_36_151# 0.030783f
C2847 net34 net31 0.080525f
C2848 state\[2\] _071_ 0.04575f
C2849 _198_/a_67_603# net30 0.017304f
C2850 FILLER_0_13_142/a_1468_375# net23 0.011746f
C2851 fanout53/a_36_160# net23 0.007461f
C2852 ctln[1] cal_itt\[0\] 0.003349f
C2853 fanout49/a_36_160# vss 0.025717f
C2854 _425_/a_2665_112# calibrate 0.029064f
C2855 _077_ FILLER_0_12_50/a_124_375# 0.008485f
C2856 _018_ FILLER_0_15_205/a_36_472# 0.00273f
C2857 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_484_472# 0.026657f
C2858 _335_/a_49_472# _098_ 0.001047f
C2859 fanout52/a_36_160# _443_/a_2665_112# 0.007884f
C2860 _155_ _365_/a_36_68# 0.053708f
C2861 net80 net35 0.028982f
C2862 ctln[2] cal 0.009784f
C2863 result[5] _419_/a_448_472# 0.00232f
C2864 net58 net19 0.044785f
C2865 FILLER_0_2_165/a_36_472# net22 0.028367f
C2866 _077_ FILLER_0_9_60/a_484_472# 0.024249f
C2867 _142_ FILLER_0_17_142/a_124_375# 0.011387f
C2868 _053_ _160_ 0.0539f
C2869 _095_ vdd 1.051346f
C2870 _413_/a_36_151# FILLER_0_3_172/a_2724_472# 0.001723f
C2871 ctln[6] net22 0.014307f
C2872 ctln[7] FILLER_0_0_130/a_36_472# 0.012298f
C2873 output33/a_224_472# net31 0.005087f
C2874 net82 _082_ 0.286003f
C2875 _008_ net19 0.027093f
C2876 net41 _067_ 0.033696f
C2877 FILLER_0_4_144/a_124_375# vdd 0.005512f
C2878 FILLER_0_22_177/a_1380_472# mask\[6\] 0.006573f
C2879 FILLER_0_16_73/a_36_472# vdd 0.08735f
C2880 result[9] ctlp[1] 0.074012f
C2881 FILLER_0_17_64/a_124_375# FILLER_0_15_59/a_484_472# 0.001188f
C2882 net27 FILLER_0_11_282/a_124_375# 0.002857f
C2883 net63 FILLER_0_19_171/a_1020_375# 0.004794f
C2884 net18 _416_/a_1288_156# 0.001147f
C2885 net54 FILLER_0_22_107/a_36_472# 0.043792f
C2886 _068_ vss 0.547532f
C2887 FILLER_0_4_197/a_1020_375# net82 0.00123f
C2888 net15 net55 1.200864f
C2889 _449_/a_2248_156# vss 0.008071f
C2890 _449_/a_2665_112# vdd 0.012848f
C2891 _297_/a_36_472# mask\[6\] 0.02557f
C2892 cal_itt\[2\] _253_/a_36_68# 0.010756f
C2893 _429_/a_36_151# net22 0.020582f
C2894 _360_/a_36_160# _163_ 0.008593f
C2895 net75 _079_ 0.071974f
C2896 _337_/a_49_472# _137_ 0.046633f
C2897 result[7] _009_ 0.697145f
C2898 _450_/a_1353_112# net6 0.054189f
C2899 _450_/a_36_151# clkc 0.033095f
C2900 FILLER_0_17_72/a_36_472# vss 0.036865f
C2901 net27 FILLER_0_14_235/a_572_375# 0.006429f
C2902 FILLER_0_14_181/a_124_375# _098_ 0.005696f
C2903 FILLER_0_4_49/a_572_375# net47 0.00654f
C2904 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_932_472# 0.001723f
C2905 _425_/a_36_151# FILLER_0_8_247/a_124_375# 0.001597f
C2906 _009_ FILLER_0_23_282/a_484_472# 0.009744f
C2907 result[2] _416_/a_2248_156# 0.001396f
C2908 FILLER_0_8_247/a_932_472# calibrate 0.008694f
C2909 _142_ FILLER_0_17_161/a_36_472# 0.00657f
C2910 _430_/a_2665_112# _091_ 0.016404f
C2911 net52 net50 0.702793f
C2912 mask\[8\] _051_ 0.003475f
C2913 net60 _421_/a_1308_423# 0.020693f
C2914 FILLER_0_22_86/a_932_472# vdd 0.001826f
C2915 net62 _418_/a_36_151# 0.029844f
C2916 _418_/a_1308_423# vss 0.001913f
C2917 _113_ _279_/a_652_68# 0.001425f
C2918 _422_/a_796_472# mask\[7\] 0.001755f
C2919 _432_/a_448_472# _136_ 0.001892f
C2920 net38 _450_/a_1284_156# 0.001291f
C2921 net38 net43 0.016358f
C2922 net52 _443_/a_1204_472# 0.005165f
C2923 _411_/a_36_151# vdd 0.077963f
C2924 _419_/a_2560_156# vdd 0.003021f
C2925 _419_/a_2665_112# vss 0.004064f
C2926 output44/a_224_472# net38 0.106923f
C2927 _091_ FILLER_0_15_212/a_572_375# 0.022582f
C2928 net57 _428_/a_36_151# 0.023215f
C2929 net39 _033_ 0.607942f
C2930 _140_ mask\[6\] 0.605898f
C2931 cal_count\[2\] FILLER_0_15_2/a_572_375# 0.015401f
C2932 output15/a_224_472# net14 0.003312f
C2933 FILLER_0_0_198/a_124_375# net21 0.004256f
C2934 _000_ _260_/a_36_68# 0.004354f
C2935 FILLER_0_7_72/a_1020_375# _053_ 0.014569f
C2936 _077_ _161_ 0.023053f
C2937 _055_ _090_ 0.040233f
C2938 FILLER_0_19_125/a_36_472# FILLER_0_18_107/a_1916_375# 0.001684f
C2939 net72 _095_ 0.136566f
C2940 FILLER_0_4_152/a_124_375# net47 0.009228f
C2941 _114_ net57 0.22998f
C2942 result[8] vdd 0.590386f
C2943 ctlp[6] vss 0.115894f
C2944 _028_ FILLER_0_5_72/a_572_375# 0.00123f
C2945 net58 output10/a_224_472# 0.025878f
C2946 _074_ net76 0.026801f
C2947 FILLER_0_4_107/a_36_472# net47 0.002982f
C2948 _086_ _395_/a_1044_488# 0.001091f
C2949 _343_/a_257_69# _093_ 0.001043f
C2950 _413_/a_448_472# vdd 0.016117f
C2951 _098_ _434_/a_36_151# 0.019342f
C2952 net57 _443_/a_36_151# 0.003322f
C2953 net66 _164_ 0.093385f
C2954 cal_itt\[3\] _122_ 0.03282f
C2955 _449_/a_1000_472# net55 0.001617f
C2956 _259_/a_455_68# _076_ 0.002372f
C2957 _055_ net22 0.084669f
C2958 mask\[5\] output19/a_224_472# 0.092961f
C2959 _187_ _408_/a_1336_472# 0.002191f
C2960 net63 _434_/a_1000_472# 0.002404f
C2961 net64 vdd 1.155692f
C2962 FILLER_0_17_56/a_36_472# _183_ 0.056523f
C2963 _440_/a_448_472# vdd 0.007263f
C2964 _440_/a_36_151# vss 0.016458f
C2965 _081_ _122_ 2.557248f
C2966 _152_ calibrate 0.020369f
C2967 FILLER_0_24_96/a_36_472# net14 0.002882f
C2968 _446_/a_2560_156# net66 0.002649f
C2969 net32 _108_ 0.035815f
C2970 mask\[1\] vdd 0.741266f
C2971 _062_ _226_/a_1044_68# 0.001944f
C2972 trim_mask\[2\] fanout49/a_36_160# 0.12844f
C2973 _256_/a_36_68# _070_ 0.019259f
C2974 net54 FILLER_0_18_139/a_932_472# 0.003365f
C2975 _411_/a_36_151# net75 0.033786f
C2976 _443_/a_1308_423# _170_ 0.043472f
C2977 _104_ net63 0.005363f
C2978 net76 FILLER_0_3_172/a_1020_375# 0.007439f
C2979 _131_ FILLER_0_17_104/a_124_375# 0.006681f
C2980 FILLER_0_11_64/a_36_472# _038_ 0.001822f
C2981 FILLER_0_5_72/a_932_472# trim_mask\[1\] 0.014619f
C2982 mask\[5\] FILLER_0_20_169/a_124_375# 0.011078f
C2983 net65 _448_/a_36_151# 0.001983f
C2984 _395_/a_36_488# _070_ 0.005165f
C2985 _176_ _131_ 1.798819f
C2986 FILLER_0_6_47/a_36_472# vdd 0.090192f
C2987 FILLER_0_6_47/a_3260_375# vss 0.061766f
C2988 FILLER_0_13_212/a_572_375# _248_/a_36_68# 0.030745f
C2989 _164_ _167_ 0.311625f
C2990 _152_ _153_ 0.002954f
C2991 _444_/a_1000_472# _054_ 0.002998f
C2992 mask\[4\] _343_/a_49_472# 0.036987f
C2993 ctln[9] vdd 0.221231f
C2994 cal_itt\[3\] _061_ 0.001311f
C2995 _228_/a_36_68# net21 0.055313f
C2996 FILLER_0_12_20/a_36_472# _450_/a_448_472# 0.058631f
C2997 net65 output48/a_224_472# 0.015306f
C2998 mask\[8\] vdd 0.423606f
C2999 _431_/a_2248_156# net36 0.001441f
C3000 FILLER_0_12_2/a_124_375# vss 0.002871f
C3001 en_co_clk net53 0.001712f
C3002 _014_ calibrate 0.403103f
C3003 _422_/a_2248_156# _108_ 0.019477f
C3004 _086_ _122_ 0.033097f
C3005 FILLER_0_18_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001684f
C3006 net65 net5 0.004409f
C3007 _098_ FILLER_0_16_154/a_932_472# 0.001701f
C3008 _328_/a_36_113# vdd 0.136098f
C3009 FILLER_0_14_81/a_124_375# vdd 0.023163f
C3010 _419_/a_1000_472# net77 0.001113f
C3011 _413_/a_1000_472# net82 0.002029f
C3012 net20 net78 1.100401f
C3013 state\[1\] _097_ 0.004171f
C3014 _104_ output21/a_224_472# 0.002459f
C3015 _089_ _122_ 0.006163f
C3016 net75 net64 0.037337f
C3017 FILLER_0_22_86/a_124_375# net14 0.003962f
C3018 FILLER_0_8_127/a_124_375# _077_ 0.005095f
C3019 net19 _006_ 0.090449f
C3020 net41 _446_/a_2665_112# 0.004501f
C3021 _256_/a_244_497# vss 0.001274f
C3022 net73 _427_/a_448_472# 0.00132f
C3023 _448_/a_36_151# net59 0.062656f
C3024 _119_ _122_ 0.155432f
C3025 calibrate net21 0.036773f
C3026 net58 fanout58/a_36_160# 0.013794f
C3027 _086_ _311_/a_2180_473# 0.001744f
C3028 net58 cal_itt\[0\] 0.229955f
C3029 trimb[4] vdd 0.081023f
C3030 _390_/a_36_68# _067_ 0.029588f
C3031 net63 net22 0.223664f
C3032 mask\[4\] net63 0.043339f
C3033 output48/a_224_472# net59 0.039277f
C3034 FILLER_0_7_72/a_1828_472# _163_ 0.002095f
C3035 output33/a_224_472# net60 0.002526f
C3036 FILLER_0_4_197/a_124_375# net59 0.001026f
C3037 net65 _000_ 0.093773f
C3038 _178_ _181_ 0.188669f
C3039 _077_ FILLER_0_8_107/a_124_375# 0.010439f
C3040 _433_/a_1204_472# _022_ 0.005308f
C3041 net74 vdd 1.451847f
C3042 trim_mask\[4\] _369_/a_36_68# 0.00407f
C3043 _095_ cal_count\[0\] 0.005211f
C3044 _408_/a_718_524# _067_ 0.006516f
C3045 _017_ net14 0.014743f
C3046 _155_ _154_ 0.18488f
C3047 _076_ _055_ 0.056585f
C3048 net20 result[5] 0.045364f
C3049 net71 FILLER_0_19_111/a_484_472# 0.004544f
C3050 net55 FILLER_0_11_78/a_36_472# 0.059367f
C3051 net5 net59 0.923076f
C3052 _274_/a_36_68# net81 0.014689f
C3053 _086_ _061_ 0.152228f
C3054 _127_ FILLER_0_11_142/a_124_375# 0.00205f
C3055 _070_ calibrate 0.675125f
C3056 _132_ _145_ 0.010994f
C3057 FILLER_0_7_72/a_1020_375# _028_ 0.003837f
C3058 _437_/a_1000_472# net14 0.028506f
C3059 state\[2\] net23 0.331644f
C3060 net68 _220_/a_67_603# 0.030878f
C3061 cal_count\[1\] vdd 0.516859f
C3062 net7 _446_/a_36_151# 0.001237f
C3063 FILLER_0_17_38/a_124_375# _041_ 0.009172f
C3064 net4 _068_ 0.040977f
C3065 _126_ _171_ 0.01633f
C3066 _115_ FILLER_0_10_94/a_484_472# 0.015061f
C3067 FILLER_0_4_123/a_124_375# _159_ 0.023643f
C3068 net41 FILLER_0_8_24/a_572_375# 0.003909f
C3069 _114_ _267_/a_672_472# 0.001566f
C3070 _274_/a_36_68# _060_ 0.02117f
C3071 net44 _190_/a_36_160# 0.015628f
C3072 output44/a_224_472# net55 0.011586f
C3073 _402_/a_728_93# _182_ 0.00263f
C3074 _399_/a_224_472# _179_ 0.002288f
C3075 _432_/a_448_472# _021_ 0.032563f
C3076 _119_ _061_ 0.132725f
C3077 FILLER_0_22_177/a_1468_375# _435_/a_36_151# 0.059049f
C3078 FILLER_0_12_136/a_1468_375# cal_count\[3\] 0.004337f
C3079 _423_/a_36_151# FILLER_0_23_44/a_1380_472# 0.001723f
C3080 FILLER_0_7_104/a_1380_472# _125_ 0.001279f
C3081 output21/a_224_472# net22 0.022576f
C3082 _068_ _311_/a_692_473# 0.002377f
C3083 _427_/a_1204_472# _095_ 0.006692f
C3084 net41 net26 0.057852f
C3085 net68 FILLER_0_5_54/a_484_472# 0.047601f
C3086 _000_ net59 0.004356f
C3087 _074_ _083_ 0.035769f
C3088 FILLER_0_5_198/a_572_375# net22 0.029657f
C3089 _076_ _313_/a_67_603# 0.024219f
C3090 trim_mask\[4\] net23 0.180803f
C3091 FILLER_0_5_54/a_1380_472# trim_mask\[1\] 0.01205f
C3092 net65 FILLER_0_1_266/a_572_375# 0.002969f
C3093 ctln[3] net8 0.003753f
C3094 _445_/a_36_151# net47 0.002364f
C3095 _118_ _315_/a_716_497# 0.001968f
C3096 _029_ net47 2.210804f
C3097 net61 ctlp[1] 2.770871f
C3098 net61 _419_/a_796_472# 0.00438f
C3099 net60 _419_/a_448_472# 0.05959f
C3100 _095_ _281_/a_672_472# 0.00134f
C3101 net79 FILLER_0_15_282/a_484_472# 0.006575f
C3102 net57 _085_ 0.211414f
C3103 net82 FILLER_0_4_213/a_572_375# 0.00123f
C3104 net57 FILLER_0_5_164/a_124_375# 0.040872f
C3105 _277_/a_36_160# _102_ 0.061995f
C3106 FILLER_0_16_89/a_932_472# _040_ 0.00702f
C3107 _443_/a_448_472# net69 0.068491f
C3108 net79 _113_ 0.002432f
C3109 FILLER_0_9_142/a_124_375# _122_ 0.004711f
C3110 net20 FILLER_0_13_228/a_36_472# 0.020589f
C3111 ctlp[6] mask\[7\] 0.011418f
C3112 _131_ _183_ 0.227229f
C3113 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_484_472# 0.001963f
C3114 _126_ _176_ 0.057877f
C3115 fanout74/a_36_113# trim_mask\[4\] 0.026261f
C3116 net82 _032_ 0.014269f
C3117 net72 net74 0.035298f
C3118 _104_ output34/a_224_472# 0.112239f
C3119 net2 cal_itt\[1\] 0.284695f
C3120 _033_ net42 0.002707f
C3121 net27 FILLER_0_9_282/a_36_472# 0.002962f
C3122 net34 output23/a_224_472# 0.021474f
C3123 FILLER_0_18_177/a_1380_472# vss -0.001894f
C3124 FILLER_0_18_177/a_1828_472# vdd 0.004845f
C3125 _072_ _311_/a_3740_473# 0.005483f
C3126 _306_/a_36_68# _126_ 0.01893f
C3127 output34/a_224_472# _421_/a_2665_112# 0.00151f
C3128 _116_ _043_ 0.002037f
C3129 net35 FILLER_0_22_128/a_124_375# 0.010439f
C3130 ctln[5] net76 0.001707f
C3131 net20 net31 0.238809f
C3132 _093_ net80 0.818824f
C3133 net52 FILLER_0_0_130/a_36_472# 0.002743f
C3134 FILLER_0_5_212/a_36_472# net59 0.058827f
C3135 _136_ _040_ 0.788826f
C3136 net16 trim_val\[2\] 0.124462f
C3137 output32/a_224_472# _103_ 0.090957f
C3138 mask\[5\] FILLER_0_20_193/a_36_472# 0.013533f
C3139 _025_ _437_/a_2665_112# 0.001245f
C3140 vdd FILLER_0_13_72/a_124_375# -0.004549f
C3141 net72 cal_count\[1\] 0.13509f
C3142 output16/a_224_472# _447_/a_2248_156# 0.001937f
C3143 ctln[9] _447_/a_448_472# 0.003564f
C3144 net16 _447_/a_796_472# 0.003278f
C3145 _412_/a_448_472# cal_itt\[1\] 0.043203f
C3146 _013_ FILLER_0_21_28/a_1916_375# 0.006025f
C3147 FILLER_0_16_57/a_1468_375# vss 0.062643f
C3148 FILLER_0_16_57/a_36_472# vdd 0.088011f
C3149 _146_ vss 0.078821f
C3150 _379_/a_36_472# trim_val\[1\] 0.00909f
C3151 _086_ _130_ 0.008816f
C3152 net2 vss 0.213737f
C3153 FILLER_0_22_86/a_124_375# _098_ 0.011864f
C3154 _093_ _304_/a_224_472# 0.002907f
C3155 cal cal_itt\[1\] 0.036277f
C3156 fanout71/a_36_113# FILLER_0_19_111/a_484_472# 0.007864f
C3157 FILLER_0_5_198/a_484_472# net21 0.051161f
C3158 _066_ _386_/a_692_472# 0.001958f
C3159 net54 _437_/a_36_151# 0.019307f
C3160 _088_ _080_ 0.003418f
C3161 output17/a_224_472# vss 0.009426f
C3162 _070_ _125_ 0.125523f
C3163 _076_ _058_ 0.912225f
C3164 _428_/a_2665_112# FILLER_0_13_142/a_124_375# 0.003325f
C3165 FILLER_0_2_93/a_124_375# net14 0.007439f
C3166 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_572_375# 0.086635f
C3167 _015_ FILLER_0_8_247/a_932_472# 0.005458f
C3168 FILLER_0_5_72/a_932_472# _164_ 0.011079f
C3169 _068_ _315_/a_716_497# 0.00217f
C3170 _076_ _315_/a_36_68# 0.001568f
C3171 _070_ _315_/a_1657_68# 0.001601f
C3172 net41 FILLER_0_23_44/a_124_375# 0.001526f
C3173 output39/a_224_472# trim[1] 0.061797f
C3174 _101_ _100_ 0.012073f
C3175 mask\[0\] FILLER_0_14_235/a_36_472# 0.287093f
C3176 FILLER_0_18_2/a_1020_375# net44 0.009108f
C3177 net21 FILLER_0_12_196/a_36_472# 0.001298f
C3178 net81 _099_ 0.140011f
C3179 mask\[4\] output34/a_224_472# 0.001777f
C3180 _126_ FILLER_0_14_181/a_124_375# 0.004632f
C3181 mask\[2\] FILLER_0_15_205/a_36_472# 0.001204f
C3182 _091_ FILLER_0_16_154/a_1380_472# 0.00133f
C3183 _341_/a_49_472# vdd 0.026636f
C3184 FILLER_0_5_172/a_36_472# vss 0.003406f
C3185 _004_ _101_ 0.001514f
C3186 FILLER_0_21_28/a_124_375# net40 0.060428f
C3187 _015_ _426_/a_796_472# 0.007696f
C3188 cal vss 0.424638f
C3189 _176_ FILLER_0_10_107/a_124_375# 0.013408f
C3190 _098_ _437_/a_1000_472# 0.007963f
C3191 _067_ _450_/a_1353_112# 0.007106f
C3192 net65 FILLER_0_3_172/a_2812_375# 0.003745f
C3193 FILLER_0_14_50/a_124_375# vdd 0.026996f
C3194 output10/a_224_472# FILLER_0_0_266/a_36_472# 0.023414f
C3195 FILLER_0_7_104/a_484_472# _131_ 0.00432f
C3196 FILLER_0_10_78/a_1468_375# _115_ 0.032403f
C3197 net41 FILLER_0_17_38/a_36_472# 0.001308f
C3198 _359_/a_36_488# _062_ 0.005596f
C3199 FILLER_0_9_72/a_124_375# vdd -0.003896f
C3200 net36 _438_/a_1204_472# 0.012234f
C3201 _081_ _160_ 0.00816f
C3202 cal_count\[3\] _134_ 0.011364f
C3203 FILLER_0_16_57/a_572_375# net55 0.004559f
C3204 FILLER_0_16_57/a_36_472# net72 0.040135f
C3205 _269_/a_36_472# vdd 0.03432f
C3206 _126_ _320_/a_672_472# 0.003662f
C3207 FILLER_0_11_142/a_484_472# vdd 0.006641f
C3208 FILLER_0_11_142/a_36_472# vss 0.008744f
C3209 _026_ vdd 0.15542f
C3210 _290_/a_224_472# result[5] 0.001638f
C3211 _077_ _246_/a_36_68# 0.006077f
C3212 trim_val\[4\] trim_mask\[4\] 0.152123f
C3213 net18 _417_/a_36_151# 0.020548f
C3214 _273_/a_36_68# FILLER_0_9_223/a_36_472# 0.015795f
C3215 _326_/a_36_160# _125_ 0.050008f
C3216 FILLER_0_16_89/a_36_472# _131_ 0.013616f
C3217 FILLER_0_12_236/a_36_472# vdd 0.086431f
C3218 FILLER_0_12_236/a_572_375# vss 0.025768f
C3219 FILLER_0_21_206/a_124_375# vdd 0.038521f
C3220 FILLER_0_21_125/a_572_375# _098_ 0.006462f
C3221 net82 FILLER_0_3_221/a_36_472# 0.015923f
C3222 _097_ vdd 0.191424f
C3223 _105_ _291_/a_36_160# 0.002075f
C3224 _074_ FILLER_0_6_231/a_484_472# 0.004409f
C3225 vss output6/a_224_472# 0.004205f
C3226 FILLER_0_4_177/a_484_472# FILLER_0_2_177/a_572_375# 0.001512f
C3227 FILLER_0_7_146/a_36_472# _068_ 0.012745f
C3228 output25/a_224_472# _214_/a_36_160# 0.027335f
C3229 _103_ vdd 0.590261f
C3230 net60 FILLER_0_17_282/a_36_472# 0.009978f
C3231 fanout66/a_36_113# _029_ 0.001684f
C3232 _085_ _267_/a_672_472# 0.006682f
C3233 _116_ _267_/a_1568_472# 0.001147f
C3234 net78 vss 0.167812f
C3235 _086_ _160_ 0.007038f
C3236 _370_/a_124_24# net47 0.017609f
C3237 FILLER_0_23_88/a_124_375# net14 0.002894f
C3238 _408_/a_728_93# _184_ 0.001389f
C3239 FILLER_0_24_274/a_36_472# FILLER_0_23_274/a_36_472# 0.05841f
C3240 valid calibrate 0.002363f
C3241 _232_/a_67_603# trim_mask\[1\] 0.022808f
C3242 FILLER_0_6_239/a_36_472# net76 0.011803f
C3243 _130_ net53 0.00399f
C3244 _335_/a_49_472# _137_ 0.03139f
C3245 FILLER_0_15_282/a_572_375# net18 0.00298f
C3246 _352_/a_49_472# _436_/a_36_151# 0.005127f
C3247 net51 FILLER_0_12_28/a_36_472# 0.005661f
C3248 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_124_375# 0.026339f
C3249 FILLER_0_7_162/a_36_472# net37 0.090785f
C3250 net52 net22 0.017993f
C3251 _119_ _160_ 0.037232f
C3252 FILLER_0_21_28/a_484_472# vdd 0.011209f
C3253 _432_/a_2665_112# net63 0.067487f
C3254 FILLER_0_3_172/a_3172_472# vdd 0.003804f
C3255 _211_/a_36_160# vdd 0.030216f
C3256 net35 _436_/a_36_151# 0.014669f
C3257 _057_ _311_/a_66_473# 0.042545f
C3258 _043_ _225_/a_36_160# 0.007958f
C3259 trimb[0] trimb[2] 0.00878f
C3260 _430_/a_36_151# _091_ 0.02228f
C3261 net82 net19 1.14585f
C3262 _427_/a_1204_472# net74 0.003057f
C3263 _314_/a_224_472# vss 0.001399f
C3264 net23 FILLER_0_21_150/a_124_375# 0.045928f
C3265 output9/a_224_472# net5 0.005189f
C3266 cal_itt\[2\] FILLER_0_3_221/a_124_375# 0.006217f
C3267 FILLER_0_10_78/a_1380_472# vss 0.002096f
C3268 result[5] vss 0.307366f
C3269 _059_ _120_ 0.0127f
C3270 _274_/a_36_68# net64 0.036017f
C3271 FILLER_0_22_177/a_932_472# net33 0.014021f
C3272 mask\[8\] _433_/a_36_151# 0.001402f
C3273 net68 _453_/a_1308_423# 0.002195f
C3274 _144_ mask\[9\] 0.001909f
C3275 net10 net11 0.007522f
C3276 FILLER_0_7_104/a_1020_375# _151_ 0.002336f
C3277 net57 FILLER_0_16_154/a_484_472# 0.001532f
C3278 net15 FILLER_0_15_72/a_36_472# 0.007185f
C3279 _013_ net55 0.239055f
C3280 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_124_375# 0.003228f
C3281 _091_ FILLER_0_12_220/a_932_472# 0.001638f
C3282 FILLER_0_17_72/a_1468_375# _131_ 0.006871f
C3283 FILLER_0_17_64/a_36_472# vss 0.006428f
C3284 FILLER_0_4_49/a_572_375# vdd 0.005972f
C3285 net10 ctln[1] 0.029592f
C3286 ctlp[2] _420_/a_2248_156# 0.001156f
C3287 _036_ net69 0.353233f
C3288 result[9] net62 0.339372f
C3289 net81 FILLER_0_15_212/a_124_375# 0.005049f
C3290 FILLER_0_5_72/a_36_472# net47 0.003953f
C3291 result[6] FILLER_0_21_286/a_484_472# 0.011149f
C3292 net20 net60 0.033919f
C3293 net50 trim_val\[0\] 0.390586f
C3294 mask\[5\] output18/a_224_472# 0.00133f
C3295 _105_ _108_ 0.548284f
C3296 FILLER_0_14_181/a_124_375# _137_ 0.006021f
C3297 _077_ net23 0.0245f
C3298 ctln[1] FILLER_0_0_232/a_124_375# 0.012033f
C3299 _161_ _061_ 0.026347f
C3300 output34/a_224_472# _419_/a_2248_156# 0.022045f
C3301 FILLER_0_15_180/a_124_375# vdd 0.016985f
C3302 _448_/a_2248_156# trim_val\[4\] 0.001534f
C3303 FILLER_0_2_177/a_484_472# net22 0.001324f
C3304 _415_/a_2248_156# fanout62/a_36_160# 0.007753f
C3305 FILLER_0_20_177/a_1020_375# _434_/a_36_151# 0.059049f
C3306 _428_/a_448_472# _095_ 0.008804f
C3307 _430_/a_2248_156# mask\[2\] 0.009336f
C3308 _412_/a_2665_112# net59 0.055415f
C3309 net33 _048_ 0.017633f
C3310 FILLER_0_5_117/a_124_375# net47 0.011773f
C3311 _147_ vss 0.006333f
C3312 net15 _216_/a_255_603# 0.002146f
C3313 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1468_375# 0.016748f
C3314 net52 _038_ 0.001152f
C3315 net63 FILLER_0_22_177/a_1380_472# 0.062289f
C3316 net38 _452_/a_2449_156# 0.058386f
C3317 FILLER_0_4_152/a_124_375# vdd -0.001403f
C3318 ctlp[3] vss 0.037106f
C3319 FILLER_0_17_133/a_124_375# _137_ 0.009198f
C3320 FILLER_0_3_78/a_36_472# vdd 0.082597f
C3321 FILLER_0_3_78/a_572_375# vss 0.04008f
C3322 _189_/a_67_603# net20 0.011939f
C3323 net55 FILLER_0_21_28/a_2812_375# 0.004005f
C3324 _452_/a_1353_112# net40 0.003745f
C3325 _321_/a_170_472# vss 0.024882f
C3326 _017_ _131_ 0.005879f
C3327 ctlp[8] net25 0.055914f
C3328 FILLER_0_13_228/a_36_472# vss 0.006491f
C3329 FILLER_0_11_142/a_124_375# net23 0.002992f
C3330 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_572_375# 0.001597f
C3331 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_124_375# 0.012001f
C3332 FILLER_0_2_101/a_36_472# vss 0.004743f
C3333 FILLER_0_4_107/a_36_472# vdd 0.119007f
C3334 FILLER_0_4_107/a_1468_375# vss 0.055184f
C3335 _077_ _439_/a_2248_156# 0.038814f
C3336 net67 _450_/a_36_151# 0.067819f
C3337 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1468_375# 0.001597f
C3338 net2 net4 0.854661f
C3339 fanout78/a_36_113# _007_ 0.003126f
C3340 _395_/a_1044_488# _071_ 0.001198f
C3341 _025_ net71 0.030824f
C3342 _435_/a_1308_423# vdd 0.012856f
C3343 trimb[1] FILLER_0_20_15/a_932_472# 0.001069f
C3344 FILLER_0_19_111/a_36_472# net14 0.00143f
C3345 _255_/a_224_552# _058_ 0.06267f
C3346 _412_/a_1308_423# net76 0.023786f
C3347 _254_/a_244_472# _072_ 0.001552f
C3348 _013_ _424_/a_796_472# 0.032857f
C3349 FILLER_0_9_72/a_1468_375# _439_/a_36_151# 0.005577f
C3350 net31 vss 0.562041f
C3351 _258_/a_36_160# net76 0.015203f
C3352 net67 _043_ 0.003726f
C3353 _098_ _205_/a_36_160# 0.033853f
C3354 FILLER_0_18_2/a_1380_472# net17 0.003603f
C3355 _074_ _251_/a_468_472# 0.001217f
C3356 _093_ FILLER_0_17_72/a_3172_472# 0.012002f
C3357 net23 _066_ 0.031928f
C3358 _075_ net22 0.180274f
C3359 _128_ _055_ 1.887595f
C3360 sample FILLER_0_9_290/a_124_375# 0.00195f
C3361 _369_/a_36_68# _157_ 0.068266f
C3362 vss FILLER_0_21_60/a_572_375# 0.021222f
C3363 vdd FILLER_0_21_60/a_36_472# 0.08419f
C3364 result[4] _417_/a_2248_156# 0.001436f
C3365 FILLER_0_19_171/a_36_472# _434_/a_36_151# 0.00271f
C3366 net54 _438_/a_2665_112# 0.032855f
C3367 _451_/a_448_472# _040_ 0.026819f
C3368 net63 FILLER_0_18_177/a_932_472# 0.063742f
C3369 _030_ _384_/a_224_472# 0.003019f
C3370 FILLER_0_9_290/a_36_472# vdd 0.094552f
C3371 FILLER_0_9_290/a_124_375# vss 0.033914f
C3372 _053_ _068_ 0.066662f
C3373 _069_ net21 0.032615f
C3374 FILLER_0_5_206/a_36_472# vdd 0.090007f
C3375 FILLER_0_5_206/a_124_375# vss 0.050652f
C3376 _019_ vdd 0.015401f
C3377 cal net4 0.026084f
C3378 _098_ mask\[6\] 0.297837f
C3379 net26 FILLER_0_23_44/a_572_375# 0.003172f
C3380 FILLER_0_13_290/a_36_472# _416_/a_36_151# 0.001723f
C3381 _077_ _311_/a_1660_473# 0.001653f
C3382 _144_ _352_/a_49_472# 0.00176f
C3383 FILLER_0_16_57/a_124_375# FILLER_0_17_56/a_124_375# 0.026339f
C3384 fanout67/a_36_160# _439_/a_36_151# 0.00246f
C3385 FILLER_0_18_100/a_36_472# net14 0.046864f
C3386 _106_ _093_ 0.045972f
C3387 _059_ _227_/a_36_160# 0.099735f
C3388 _428_/a_2248_156# net53 0.001188f
C3389 _144_ net35 0.036236f
C3390 vdd _145_ 0.082579f
C3391 net64 _099_ 0.007017f
C3392 net23 net37 0.01763f
C3393 _069_ _070_ 0.257147f
C3394 FILLER_0_19_195/a_124_375# vdd 0.03587f
C3395 net41 _402_/a_728_93# 0.032823f
C3396 FILLER_0_5_54/a_484_472# net47 0.006652f
C3397 _188_ _039_ 0.002071f
C3398 output38/a_224_472# _445_/a_36_151# 0.199812f
C3399 _099_ mask\[1\] 0.19135f
C3400 _242_/a_36_160# net47 0.028264f
C3401 _077_ _056_ 1.777574f
C3402 _389_/a_36_148# vdd 0.039639f
C3403 net82 FILLER_0_3_172/a_484_472# 0.008052f
C3404 output34/a_224_472# result[7] 0.057094f
C3405 _020_ _131_ 0.011012f
C3406 net78 mask\[7\] 0.001437f
C3407 _173_ net51 0.016607f
C3408 net18 _418_/a_36_151# 0.017941f
C3409 FILLER_0_17_142/a_124_375# vss 0.008753f
C3410 FILLER_0_17_142/a_572_375# vdd 0.012885f
C3411 net57 FILLER_0_13_100/a_36_472# 0.077963f
C3412 net28 vss 0.185012f
C3413 _137_ FILLER_0_16_154/a_932_472# 0.004753f
C3414 _320_/a_36_472# mask\[0\] 0.001026f
C3415 net46 net17 0.791341f
C3416 _253_/a_672_68# _074_ 0.001857f
C3417 _232_/a_67_603# _164_ 0.076123f
C3418 output42/a_224_472# _444_/a_36_151# 0.002701f
C3419 _077_ _392_/a_36_68# 0.055912f
C3420 output27/a_224_472# _425_/a_2665_112# 0.021504f
C3421 FILLER_0_18_76/a_124_375# vdd 0.019258f
C3422 trim[1] net40 0.043114f
C3423 FILLER_0_18_107/a_36_472# FILLER_0_17_104/a_484_472# 0.026657f
C3424 _131_ FILLER_0_11_109/a_124_375# 0.001048f
C3425 _429_/a_2248_156# vdd -0.006752f
C3426 _429_/a_1204_472# vss 0.002428f
C3427 _038_ _172_ 0.050158f
C3428 _423_/a_1000_472# vdd 0.001833f
C3429 mask\[4\] FILLER_0_19_171/a_124_375# 0.001988f
C3430 FILLER_0_18_2/a_2812_375# vdd 0.021655f
C3431 FILLER_0_10_247/a_124_375# vss 0.006235f
C3432 FILLER_0_10_247/a_36_472# vdd 0.111658f
C3433 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_124_375# 0.001597f
C3434 _069_ FILLER_0_9_142/a_36_472# 0.035528f
C3435 net82 cal_itt\[0\] 0.063072f
C3436 FILLER_0_19_28/a_572_375# _452_/a_36_151# 0.0027f
C3437 FILLER_0_14_181/a_36_472# _113_ 0.004214f
C3438 net57 mask\[2\] 0.022012f
C3439 FILLER_0_17_226/a_36_472# _106_ 0.050907f
C3440 FILLER_0_7_72/a_1468_375# net52 0.003576f
C3441 _365_/a_36_68# net14 0.017522f
C3442 _111_ _098_ 0.014998f
C3443 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_36_472# 0.086635f
C3444 _126_ _017_ 0.071134f
C3445 FILLER_0_17_72/a_1828_472# net36 0.028046f
C3446 mask\[4\] FILLER_0_18_171/a_36_472# 0.01222f
C3447 net65 en 0.001469f
C3448 _421_/a_2248_156# _109_ 0.001349f
C3449 _431_/a_2560_156# _137_ 0.002967f
C3450 trim_mask\[2\] FILLER_0_3_78/a_572_375# 0.011713f
C3451 FILLER_0_17_161/a_36_472# vss 0.003343f
C3452 _131_ FILLER_0_14_107/a_1468_375# 0.051201f
C3453 fanout59/a_36_160# net18 0.003981f
C3454 net52 FILLER_0_6_47/a_2812_375# 0.018463f
C3455 FILLER_0_22_128/a_36_472# vss 0.001309f
C3456 FILLER_0_22_128/a_484_472# vdd 0.002467f
C3457 _281_/a_672_472# _097_ 0.002131f
C3458 net32 _421_/a_448_472# 0.022214f
C3459 _096_ _098_ 0.00638f
C3460 _422_/a_448_472# _109_ 0.006344f
C3461 _424_/a_2665_112# vss 0.013462f
C3462 _024_ _435_/a_1308_423# 0.002661f
C3463 result[6] _420_/a_796_472# 0.002296f
C3464 _098_ FILLER_0_19_111/a_36_472# 0.003915f
C3465 _144_ FILLER_0_19_125/a_124_375# 0.012834f
C3466 _128_ _315_/a_36_68# 0.04902f
C3467 net29 _045_ 0.344478f
C3468 _086_ _267_/a_36_472# 0.070088f
C3469 mask\[5\] FILLER_0_20_177/a_1380_472# 0.016114f
C3470 _442_/a_448_472# vdd 0.006758f
C3471 _442_/a_36_151# vss 0.021278f
C3472 _260_/a_36_68# _080_ 0.001888f
C3473 net55 _452_/a_2449_156# 0.015878f
C3474 trim_val\[4\] _066_ 0.015621f
C3475 _053_ FILLER_0_6_47/a_3260_375# 0.002746f
C3476 net15 trim_val\[3\] 0.068273f
C3477 _447_/a_2560_156# vss 0.00126f
C3478 net23 FILLER_0_5_148/a_484_472# 0.047258f
C3479 _430_/a_2248_156# net20 0.001893f
C3480 _413_/a_1308_423# vdd 0.002686f
C3481 _126_ _250_/a_36_68# 0.022134f
C3482 _445_/a_36_151# vdd 0.052935f
C3483 _029_ vdd 0.223076f
C3484 _029_ _365_/a_244_472# 0.001956f
C3485 FILLER_0_15_290/a_36_472# output30/a_224_472# 0.001711f
C3486 _428_/a_448_472# net74 0.019814f
C3487 mask\[7\] _147_ 0.295801f
C3488 FILLER_0_15_116/a_484_472# net70 0.049569f
C3489 _176_ _095_ 0.064978f
C3490 FILLER_0_15_116/a_124_375# net53 0.009286f
C3491 _130_ _127_ 0.195571f
C3492 net29 _192_/a_67_603# 0.017997f
C3493 _377_/a_36_472# trim_mask\[1\] 0.001763f
C3494 en net59 0.490893f
C3495 _123_ FILLER_0_7_233/a_124_375# 0.007717f
C3496 ctlp[3] mask\[7\] 0.103955f
C3497 mask\[5\] FILLER_0_18_177/a_1020_375# 0.001604f
C3498 net81 _082_ 0.001633f
C3499 FILLER_0_15_282/a_572_375# _417_/a_36_151# 0.001597f
C3500 _306_/a_36_68# _095_ 0.001366f
C3501 _104_ _422_/a_36_151# 0.032235f
C3502 mask\[2\] FILLER_0_15_212/a_1380_472# 0.001225f
C3503 _141_ _146_ 0.020044f
C3504 FILLER_0_16_73/a_36_472# _176_ 0.013449f
C3505 net47 FILLER_0_6_37/a_36_472# 0.001161f
C3506 net75 FILLER_0_10_247/a_36_472# 0.001184f
C3507 _422_/a_36_151# _421_/a_2665_112# 0.001725f
C3508 net55 _423_/a_448_472# 0.00206f
C3509 net82 FILLER_0_2_171/a_36_472# 0.001777f
C3510 _072_ _375_/a_692_497# 0.001113f
C3511 net23 FILLER_0_19_155/a_36_472# 0.019429f
C3512 _123_ vdd 0.214703f
C3513 _449_/a_2665_112# _176_ 0.048319f
C3514 _431_/a_1000_472# _020_ 0.009685f
C3515 result[6] _421_/a_1204_472# 0.005361f
C3516 mask\[7\] _435_/a_448_472# 0.064472f
C3517 trim_val\[4\] net37 0.003661f
C3518 net60 vss 0.382678f
C3519 trim_val\[0\] _054_ 0.010002f
C3520 net61 net62 0.874859f
C3521 _136_ _438_/a_36_151# 0.030558f
C3522 net81 _426_/a_448_472# 0.003907f
C3523 FILLER_0_15_212/a_124_375# mask\[1\] 0.007876f
C3524 net50 FILLER_0_2_93/a_36_472# 0.008147f
C3525 FILLER_0_12_20/a_36_472# _039_ 0.007881f
C3526 net56 FILLER_0_16_154/a_932_472# 0.001401f
C3527 FILLER_0_9_28/a_1380_472# vdd 0.01306f
C3528 _062_ _117_ 0.042699f
C3529 _057_ _114_ 0.30288f
C3530 net52 _448_/a_2665_112# 0.039348f
C3531 FILLER_0_16_73/a_484_472# _040_ 0.004877f
C3532 FILLER_0_7_59/a_124_375# fanout67/a_36_160# 0.001597f
C3533 _134_ _120_ 0.047627f
C3534 net58 fanout76/a_36_160# 0.055026f
C3535 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_484_472# 0.013277f
C3536 net41 net17 0.911377f
C3537 FILLER_0_2_101/a_124_375# _154_ 0.003932f
C3538 FILLER_0_4_107/a_124_375# _153_ 0.073219f
C3539 FILLER_0_4_107/a_1020_375# _154_ 0.013746f
C3540 FILLER_0_16_73/a_572_375# _131_ 0.011479f
C3541 _413_/a_2248_156# vdd -0.006767f
C3542 net36 FILLER_0_16_115/a_36_472# 0.003805f
C3543 _189_/a_67_603# vss 0.004088f
C3544 FILLER_0_18_2/a_3260_375# _452_/a_36_151# 0.001597f
C3545 FILLER_0_20_15/a_572_375# vdd 0.003301f
C3546 _356_/a_36_472# _438_/a_36_151# 0.004432f
C3547 FILLER_0_13_65/a_124_375# _095_ 0.002035f
C3548 FILLER_0_14_181/a_124_375# _095_ 0.005538f
C3549 net17 FILLER_0_20_15/a_36_472# 0.004375f
C3550 _132_ FILLER_0_15_116/a_484_472# 0.010148f
C3551 FILLER_0_9_223/a_572_375# _223_/a_36_160# 0.001177f
C3552 _431_/a_2560_156# net56 0.001258f
C3553 FILLER_0_3_221/a_36_472# FILLER_0_3_212/a_36_472# 0.001963f
C3554 FILLER_0_15_205/a_36_472# vss 0.003239f
C3555 FILLER_0_5_136/a_36_472# vss 0.007658f
C3556 net79 FILLER_0_12_236/a_572_375# 0.010684f
C3557 _126_ FILLER_0_11_135/a_124_375# 0.008245f
C3558 net58 _412_/a_1456_156# 0.001045f
C3559 FILLER_0_5_198/a_36_472# net37 0.0114f
C3560 net75 _123_ 0.173358f
C3561 _086_ FILLER_0_4_177/a_36_472# 0.001464f
C3562 mask\[5\] _340_/a_36_160# 0.031249f
C3563 FILLER_0_17_56/a_484_472# vss 0.006298f
C3564 net23 net13 0.018808f
C3565 _135_ vss 0.097337f
C3566 net23 FILLER_0_22_128/a_2812_375# 0.050811f
C3567 FILLER_0_18_53/a_124_375# FILLER_0_18_37/a_1468_375# 0.012222f
C3568 _079_ _082_ 0.709481f
C3569 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_124_375# 0.012001f
C3570 net78 net79 0.009641f
C3571 cal_count\[2\] _402_/a_728_93# 0.036871f
C3572 _134_ FILLER_0_9_105/a_572_375# 0.02163f
C3573 _141_ _346_/a_665_69# 0.002048f
C3574 ctln[4] net11 0.194506f
C3575 _448_/a_2665_112# _387_/a_36_113# 0.010064f
C3576 _448_/a_1308_423# _037_ 0.034533f
C3577 _444_/a_448_472# net40 0.055844f
C3578 net63 _435_/a_36_151# 0.017194f
C3579 trim[0] _446_/a_36_151# 0.044586f
C3580 net38 _446_/a_1308_423# 0.010331f
C3581 FILLER_0_9_28/a_3260_375# fanout67/a_36_160# 0.001925f
C3582 net34 _422_/a_1204_472# 0.001029f
C3583 fanout54/a_36_160# FILLER_0_19_155/a_124_375# 0.005705f
C3584 net62 FILLER_0_13_212/a_932_472# 0.059367f
C3585 FILLER_0_19_55/a_124_375# FILLER_0_19_47/a_572_375# 0.012001f
C3586 net41 _452_/a_36_151# 0.036301f
C3587 _033_ net67 0.148585f
C3588 _012_ FILLER_0_23_44/a_932_472# 0.001572f
C3589 _441_/a_36_151# _030_ 0.005324f
C3590 FILLER_0_9_105/a_124_375# vdd 0.029831f
C3591 vdd _202_/a_36_160# 0.06338f
C3592 ctln[4] ctln[1] 0.002283f
C3593 _256_/a_36_68# calibrate 0.02084f
C3594 _398_/a_36_113# net17 0.002702f
C3595 input2/a_36_113# clk 0.021981f
C3596 _335_/a_49_472# mask\[1\] 0.032497f
C3597 mask\[0\] FILLER_0_12_220/a_1468_375# 0.001484f
C3598 _028_ FILLER_0_6_47/a_3260_375# 0.013006f
C3599 vss _433_/a_2665_112# 0.035903f
C3600 FILLER_0_14_91/a_124_375# _177_ 0.00134f
C3601 FILLER_0_18_139/a_1020_375# vss 0.032606f
C3602 FILLER_0_18_139/a_1468_375# vdd 0.015542f
C3603 FILLER_0_1_204/a_36_472# net59 0.067975f
C3604 net41 FILLER_0_16_37/a_36_472# 0.009425f
C3605 trimb[4] net44 0.127019f
C3606 net49 _440_/a_796_472# 0.003597f
C3607 FILLER_0_18_2/a_1468_375# output44/a_224_472# 0.032639f
C3608 _158_ _154_ 0.008872f
C3609 _410_/a_36_68# _039_ 0.016062f
C3610 result[5] net79 0.036275f
C3611 FILLER_0_15_116/a_572_375# FILLER_0_14_107/a_1468_375# 0.026339f
C3612 FILLER_0_15_116/a_36_472# FILLER_0_14_107/a_1020_375# 0.001723f
C3613 _086_ _113_ 0.072034f
C3614 _394_/a_1936_472# cal_count\[1\] 0.008364f
C3615 net63 _139_ 0.003073f
C3616 net68 _440_/a_796_472# 0.021463f
C3617 FILLER_0_15_142/a_36_472# net53 0.080484f
C3618 _032_ net69 0.347645f
C3619 output23/a_224_472# vss 0.075684f
C3620 _142_ FILLER_0_18_107/a_2724_472# 0.001549f
C3621 _100_ vdd 0.212037f
C3622 _273_/a_36_68# vss 0.095582f
C3623 FILLER_0_24_130/a_124_375# vdd 0.027763f
C3624 _370_/a_124_24# vdd 0.018613f
C3625 FILLER_0_7_104/a_1020_375# _062_ 0.003073f
C3626 cal_itt\[3\] _087_ 0.002881f
C3627 mask\[7\] FILLER_0_22_128/a_36_472# 0.013408f
C3628 _122_ net23 0.276617f
C3629 _080_ net59 0.038227f
C3630 _079_ _265_/a_244_68# 0.021777f
C3631 _004_ vdd 0.448886f
C3632 FILLER_0_21_142/a_572_375# net54 0.043619f
C3633 output31/a_224_472# net62 0.030092f
C3634 _427_/a_36_151# FILLER_0_14_123/a_36_472# 0.004032f
C3635 _305_/a_36_159# vdd 0.017293f
C3636 _067_ FILLER_0_12_28/a_36_472# 0.0127f
C3637 _148_ FILLER_0_22_128/a_36_472# 0.010386f
C3638 FILLER_0_15_116/a_124_375# _451_/a_36_151# 0.006111f
C3639 _072_ _074_ 2.017168f
C3640 _090_ net21 0.038093f
C3641 net35 FILLER_0_22_128/a_3172_472# 0.014415f
C3642 _261_/a_36_160# _059_ 0.004993f
C3643 _430_/a_1204_472# net63 0.013728f
C3644 FILLER_0_14_81/a_124_375# _176_ 0.001549f
C3645 _087_ _081_ 0.002169f
C3646 net41 FILLER_0_12_28/a_124_375# 0.003909f
C3647 net32 _419_/a_36_151# 0.006506f
C3648 result[2] net19 0.065763f
C3649 FILLER_0_2_111/a_36_472# trim_mask\[3\] 0.007915f
C3650 net36 _451_/a_2449_156# 0.016229f
C3651 net55 FILLER_0_17_56/a_572_375# 0.020564f
C3652 _256_/a_1164_497# _076_ 0.001871f
C3653 FILLER_0_14_91/a_36_472# _043_ 0.001779f
C3654 net73 FILLER_0_18_107/a_1468_375# 0.024898f
C3655 net58 _412_/a_2560_156# 0.005111f
C3656 _154_ net14 0.02512f
C3657 net68 FILLER_0_6_47/a_932_472# 0.014935f
C3658 _079_ _112_ 0.004464f
C3659 FILLER_0_10_78/a_124_375# net52 0.008557f
C3660 _020_ _137_ 0.228674f
C3661 FILLER_0_15_142/a_484_472# net53 0.044267f
C3662 net38 _160_ 0.00247f
C3663 ctln[7] net14 0.197449f
C3664 _418_/a_36_151# _417_/a_36_151# 0.005373f
C3665 FILLER_0_18_107/a_124_375# vdd 0.030961f
C3666 _180_ _041_ 0.00244f
C3667 FILLER_0_14_181/a_124_375# mask\[1\] 0.044784f
C3668 trim_mask\[1\] FILLER_0_6_47/a_1828_472# 0.007542f
C3669 net39 _445_/a_796_472# 0.002296f
C3670 _383_/a_36_472# vss 0.002794f
C3671 net23 _049_ 0.215528f
C3672 _431_/a_36_151# _136_ 0.03371f
C3673 _429_/a_36_151# FILLER_0_15_205/a_124_375# 0.059049f
C3674 _103_ _099_ 0.025799f
C3675 net29 _287_/a_36_472# 0.002936f
C3676 _413_/a_1204_472# net21 0.011236f
C3677 FILLER_0_11_101/a_484_472# _070_ 0.017841f
C3678 fanout54/a_36_160# net23 0.05522f
C3679 _433_/a_36_151# _145_ 0.004437f
C3680 net20 FILLER_0_15_212/a_1380_472# 0.001449f
C3681 _070_ _090_ 0.369847f
C3682 net17 _164_ 0.007595f
C3683 net24 _211_/a_36_160# 0.021941f
C3684 _052_ FILLER_0_18_37/a_484_472# 0.003861f
C3685 FILLER_0_17_200/a_484_472# net63 0.003767f
C3686 _073_ net76 0.040554f
C3687 _377_/a_36_472# _164_ 0.03259f
C3688 _074_ net47 0.012724f
C3689 _086_ _118_ 0.166544f
C3690 FILLER_0_12_220/a_484_472# _060_ 0.003379f
C3691 net22 net21 1.937266f
C3692 mask\[4\] net21 0.049513f
C3693 _114_ cal_count\[3\] 0.081644f
C3694 _176_ net74 0.067915f
C3695 FILLER_0_13_228/a_36_472# net79 0.006824f
C3696 FILLER_0_4_99/a_36_472# FILLER_0_4_107/a_36_472# 0.002296f
C3697 ctlp[1] _421_/a_2560_156# 0.001062f
C3698 _065_ net49 0.001576f
C3699 FILLER_0_11_282/a_36_472# _416_/a_448_472# 0.011962f
C3700 FILLER_0_24_274/a_124_375# vdd 0.012632f
C3701 fanout82/a_36_113# _316_/a_848_380# 0.001292f
C3702 state\[2\] FILLER_0_13_142/a_1468_375# 0.018691f
C3703 net53 FILLER_0_13_142/a_484_472# 0.059444f
C3704 _091_ FILLER_0_10_214/a_36_472# 0.001357f
C3705 FILLER_0_5_72/a_36_472# vdd 0.107678f
C3706 FILLER_0_5_72/a_1468_375# vss 0.057097f
C3707 net3 FILLER_0_15_10/a_124_375# 0.035504f
C3708 _446_/a_2560_156# net17 0.00101f
C3709 _270_/a_36_472# _087_ 0.02676f
C3710 _065_ net68 0.194392f
C3711 net60 mask\[7\] 0.001053f
C3712 FILLER_0_7_72/a_2724_472# _219_/a_36_160# 0.001448f
C3713 _119_ _118_ 0.001596f
C3714 _086_ _087_ 0.015938f
C3715 net54 FILLER_0_19_142/a_36_472# 0.07544f
C3716 _057_ _085_ 0.543871f
C3717 FILLER_0_9_28/a_1916_375# net68 0.050307f
C3718 _303_/a_36_472# net36 0.006675f
C3719 _176_ cal_count\[1\] 0.297763f
C3720 _070_ net22 0.032551f
C3721 _102_ net36 0.003446f
C3722 _076_ _152_ 0.063574f
C3723 _068_ _081_ 0.006663f
C3724 _430_/a_2248_156# vss 0.030251f
C3725 net75 _004_ 0.003999f
C3726 net75 _305_/a_36_159# 0.049563f
C3727 _089_ _087_ 0.002217f
C3728 net41 net39 0.003649f
C3729 FILLER_0_4_197/a_932_472# _088_ 0.014643f
C3730 FILLER_0_6_90/a_572_375# _163_ 0.007844f
C3731 FILLER_0_5_117/a_124_375# vdd 0.035079f
C3732 _408_/a_1336_472# vss 0.001022f
C3733 _408_/a_728_93# vdd 0.024163f
C3734 _417_/a_2560_156# net30 0.049334f
C3735 FILLER_0_2_93/a_124_375# net69 0.015032f
C3736 output9/a_224_472# en 0.011047f
C3737 vdd _107_ 0.038236f
C3738 _408_/a_718_524# net17 0.012884f
C3739 net41 _039_ 0.030362f
C3740 FILLER_0_18_177/a_1020_375# FILLER_0_20_177/a_932_472# 0.0027f
C3741 FILLER_0_12_136/a_932_472# _126_ 0.014483f
C3742 FILLER_0_19_134/a_124_375# _145_ 0.023167f
C3743 net61 net33 0.043271f
C3744 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_484_472# 0.026657f
C3745 _161_ _267_/a_36_472# 0.043279f
C3746 _432_/a_1204_472# net80 0.009362f
C3747 _058_ net14 0.40635f
C3748 _129_ vss 0.141494f
C3749 net15 _449_/a_1000_472# 0.056791f
C3750 cal_count\[2\] net17 0.074204f
C3751 FILLER_0_8_24/a_36_472# net17 0.045619f
C3752 FILLER_0_10_78/a_932_472# _120_ 0.003672f
C3753 _136_ _038_ 0.061274f
C3754 FILLER_0_22_128/a_484_472# _433_/a_36_151# 0.001653f
C3755 FILLER_0_15_142/a_572_375# FILLER_0_15_150/a_36_472# 0.086635f
C3756 _091_ net62 0.019946f
C3757 FILLER_0_13_65/a_124_375# net74 0.020091f
C3758 _426_/a_448_472# net64 0.054931f
C3759 _096_ _126_ 0.258912f
C3760 vss _034_ 0.008249f
C3761 net21 net11 0.10869f
C3762 _086_ _068_ 0.080666f
C3763 FILLER_0_23_274/a_124_375# vdd 0.014998f
C3764 FILLER_0_16_57/a_572_375# FILLER_0_18_61/a_36_472# 0.001512f
C3765 output20/a_224_472# _108_ 0.022243f
C3766 _187_ _042_ 0.009526f
C3767 net57 FILLER_0_3_172/a_36_472# 0.001007f
C3768 net58 _425_/a_2665_112# 0.069807f
C3769 net28 net79 0.116857f
C3770 net57 _386_/a_124_24# 0.037058f
C3771 _038_ _070_ 0.075667f
C3772 _119_ _068_ 0.040944f
C3773 _449_/a_796_472# _038_ 0.018626f
C3774 mask\[9\] _354_/a_49_472# 0.032687f
C3775 FILLER_0_16_57/a_36_472# _176_ 0.075537f
C3776 output38/a_224_472# FILLER_0_3_2/a_36_472# 0.035046f
C3777 _220_/a_67_603# vdd 0.020078f
C3778 FILLER_0_18_2/a_932_472# trimb[1] 0.011513f
C3779 _076_ net21 0.031683f
C3780 _412_/a_1204_472# cal_itt\[1\] 0.001547f
C3781 FILLER_0_9_142/a_124_375# _118_ 0.06224f
C3782 net64 FILLER_0_8_239/a_36_472# 0.002666f
C3783 ctlp[7] _050_ 0.153673f
C3784 _056_ _061_ 0.445098f
C3785 net76 net1 0.059026f
C3786 _436_/a_36_151# FILLER_0_22_107/a_124_375# 0.026916f
C3787 net65 FILLER_0_2_177/a_124_375# 0.018094f
C3788 _025_ _436_/a_2248_156# 0.001054f
C3789 FILLER_0_12_2/a_484_472# _450_/a_36_151# 0.059367f
C3790 result[7] _421_/a_1204_472# 0.014927f
C3791 _432_/a_2560_156# _093_ 0.007613f
C3792 FILLER_0_7_59/a_124_375# trim_mask\[1\] 0.001548f
C3793 net74 FILLER_0_13_142/a_124_375# 0.002722f
C3794 FILLER_0_5_54/a_36_472# vss 0.001756f
C3795 FILLER_0_5_54/a_484_472# vdd 0.003166f
C3796 trimb[1] FILLER_0_20_2/a_36_472# 0.003628f
C3797 cal_count\[2\] _452_/a_36_151# 0.006982f
C3798 FILLER_0_10_247/a_124_375# net79 0.00498f
C3799 FILLER_0_20_31/a_36_472# net40 0.045181f
C3800 result[9] net18 0.019413f
C3801 _242_/a_36_160# vdd 0.007995f
C3802 _070_ _076_ 0.198272f
C3803 net52 FILLER_0_3_78/a_124_375# 0.017889f
C3804 fanout64/a_36_160# net64 0.043709f
C3805 _093_ FILLER_0_17_218/a_572_375# 0.0029f
C3806 _441_/a_448_472# _164_ 0.016938f
C3807 FILLER_0_10_28/a_124_375# output6/a_224_472# 0.002633f
C3808 _413_/a_36_151# _088_ 0.001289f
C3809 _412_/a_36_151# net76 0.001169f
C3810 net68 net51 0.008885f
C3811 result[8] FILLER_0_24_274/a_1380_472# 0.005458f
C3812 net3 _278_/a_36_160# 0.014154f
C3813 net52 FILLER_0_2_101/a_124_375# 0.007787f
C3814 _173_ _067_ 0.011854f
C3815 output23/a_224_472# mask\[7\] 0.046766f
C3816 FILLER_0_16_37/a_36_472# cal_count\[2\] 0.008691f
C3817 _346_/a_49_472# _144_ 0.036821f
C3818 vss output30/a_224_472# 0.030732f
C3819 _064_ _446_/a_448_472# 0.01156f
C3820 _122_ FILLER_0_5_198/a_36_472# 0.00305f
C3821 _443_/a_2560_156# vss 0.002467f
C3822 net63 FILLER_0_15_205/a_124_375# 0.001597f
C3823 _088_ FILLER_0_4_213/a_124_375# 0.016013f
C3824 _073_ _083_ 0.097365f
C3825 _369_/a_36_68# _160_ 0.015312f
C3826 _273_/a_36_68# net4 0.06843f
C3827 _432_/a_36_151# FILLER_0_17_161/a_124_375# 0.035117f
C3828 _141_ FILLER_0_17_161/a_36_472# 0.011708f
C3829 FILLER_0_2_177/a_124_375# net59 0.005212f
C3830 net28 _416_/a_2665_112# 0.008877f
C3831 _408_/a_718_524# FILLER_0_12_28/a_124_375# 0.001192f
C3832 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_124_375# 0.004426f
C3833 net63 _098_ 0.055686f
C3834 _021_ mask\[4\] 0.018108f
C3835 FILLER_0_17_226/a_124_375# net63 0.00507f
C3836 net17 FILLER_0_23_44/a_572_375# 0.001332f
C3837 _013_ FILLER_0_18_61/a_36_472# 0.01628f
C3838 _017_ _095_ 0.002789f
C3839 _187_ cal_count\[3\] 0.031898f
C3840 net15 FILLER_0_6_47/a_2364_375# 0.022624f
C3841 FILLER_0_19_47/a_36_472# FILLER_0_18_37/a_1020_375# 0.001684f
C3842 _091_ _429_/a_448_472# 0.034713f
C3843 net19 _420_/a_2665_112# 0.012322f
C3844 ctln[8] output16/a_224_472# 0.006971f
C3845 net57 vss 0.818311f
C3846 _132_ _124_ 0.005668f
C3847 _085_ cal_count\[3\] 0.653405f
C3848 _076_ FILLER_0_9_142/a_36_472# 0.038562f
C3849 _068_ FILLER_0_9_142/a_124_375# 0.008226f
C3850 ctlp[2] net78 0.369805f
C3851 _340_/a_36_160# _348_/a_49_472# 0.001528f
C3852 _144_ FILLER_0_19_125/a_36_472# 0.153815f
C3853 FILLER_0_17_38/a_124_375# vdd 0.01443f
C3854 FILLER_0_4_144/a_36_472# net47 0.008498f
C3855 fanout75/a_36_113# net37 0.010418f
C3856 result[2] _193_/a_36_160# 0.040932f
C3857 _219_/a_36_160# vss 0.00157f
C3858 _098_ _433_/a_1308_423# 0.010653f
C3859 net16 trim_val\[0\] 0.00463f
C3860 _057_ _310_/a_49_472# 0.015839f
C3861 FILLER_0_3_2/a_124_375# vss 0.007235f
C3862 FILLER_0_3_2/a_36_472# vdd 0.106665f
C3863 result[0] net5 0.001104f
C3864 net34 net35 2.497277f
C3865 mask\[0\] state\[1\] 0.064758f
C3866 output8/a_224_472# _078_ 0.001267f
C3867 _027_ vss 0.011873f
C3868 _020_ FILLER_0_18_107/a_2276_472# 0.004069f
C3869 net36 FILLER_0_15_180/a_484_472# 0.00702f
C3870 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_572_375# 0.086635f
C3871 net23 _160_ 0.030085f
C3872 ctlp[1] _419_/a_2665_112# 0.009197f
C3873 net60 net79 0.113281f
C3874 _037_ vss 0.051886f
C3875 _274_/a_1612_497# state\[0\] 0.001071f
C3876 _267_/a_36_472# _071_ 0.001682f
C3877 _161_ _113_ 0.201931f
C3878 FILLER_0_5_109/a_484_472# _163_ 0.005054f
C3879 _327_/a_36_472# _126_ 0.011444f
C3880 _448_/a_1204_472# net22 0.002283f
C3881 _434_/a_2248_156# mask\[6\] 0.022666f
C3882 mask\[8\] _354_/a_257_69# 0.003809f
C3883 FILLER_0_7_162/a_124_375# calibrate 0.014255f
C3884 FILLER_0_21_28/a_1916_375# _012_ 0.023886f
C3885 _443_/a_2665_112# FILLER_0_2_165/a_36_472# 0.007491f
C3886 net52 _158_ 0.001338f
C3887 FILLER_0_16_57/a_36_472# _183_ 0.004107f
C3888 _413_/a_796_472# vdd 0.001569f
C3889 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_36_472# 0.086743f
C3890 FILLER_0_15_212/a_1380_472# vss 0.007595f
C3891 _432_/a_2665_112# _136_ 0.002691f
C3892 FILLER_0_15_116/a_484_472# vdd 0.006111f
C3893 _408_/a_728_93# cal_count\[0\] 0.007633f
C3894 _189_/a_67_603# net79 0.008944f
C3895 vss FILLER_0_6_37/a_124_375# 0.030885f
C3896 vdd FILLER_0_6_37/a_36_472# 0.138008f
C3897 net81 net19 0.786284f
C3898 FILLER_0_11_135/a_36_472# _118_ 0.002496f
C3899 _432_/a_2665_112# net21 0.005773f
C3900 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_36_472# 0.086743f
C3901 _059_ _062_ 0.161331f
C3902 _412_/a_1000_472# cal_itt\[1\] 0.012926f
C3903 output48/a_224_472# output37/a_224_472# 0.005147f
C3904 net57 FILLER_0_2_165/a_124_375# 0.007153f
C3905 FILLER_0_4_197/a_1380_472# vdd 0.00581f
C3906 _149_ FILLER_0_20_98/a_124_375# 0.020028f
C3907 _134_ FILLER_0_10_107/a_484_472# 0.020725f
C3908 net72 FILLER_0_17_38/a_124_375# 0.041464f
C3909 FILLER_0_14_181/a_124_375# _097_ 0.001668f
C3910 _375_/a_36_68# _062_ 0.012855f
C3911 net52 net14 0.072003f
C3912 cal_itt\[2\] _083_ 0.10423f
C3913 fanout70/a_36_113# fanout73/a_36_113# 0.001578f
C3914 fanout81/a_36_160# net2 0.044793f
C3915 output37/a_224_472# net5 0.072504f
C3916 _120_ FILLER_0_9_72/a_932_472# 0.001709f
C3917 _161_ _118_ 0.023939f
C3918 FILLER_0_10_107/a_36_472# vdd 0.117291f
C3919 FILLER_0_10_107/a_572_375# vss 0.017711f
C3920 _420_/a_2665_112# _009_ 0.001752f
C3921 _445_/a_2248_156# net40 0.004545f
C3922 net1 _083_ 0.30074f
C3923 ctlp[3] ctlp[2] 0.006764f
C3924 net48 _079_ 0.012855f
C3925 input5/a_36_113# vss 0.005833f
C3926 FILLER_0_5_128/a_124_375# _152_ 0.017496f
C3927 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_124_375# 0.012001f
C3928 mask\[4\] FILLER_0_18_177/a_36_472# 0.018019f
C3929 _131_ _154_ 0.019221f
C3930 ctln[2] rstn 0.017812f
C3931 _272_/a_36_472# net76 0.04597f
C3932 _432_/a_36_151# _098_ 0.00957f
C3933 FILLER_0_20_177/a_1468_375# vss 0.053913f
C3934 FILLER_0_20_177/a_36_472# vdd 0.114932f
C3935 output8/a_224_472# _411_/a_448_472# 0.010723f
C3936 net28 output29/a_224_472# 0.028512f
C3937 net50 _441_/a_2560_156# 0.008865f
C3938 _440_/a_796_472# net47 0.002508f
C3939 _230_/a_244_68# _060_ 0.002039f
C3940 _412_/a_448_472# fanout81/a_36_160# 0.00998f
C3941 mask\[8\] FILLER_0_22_86/a_124_375# 0.014263f
C3942 FILLER_0_4_49/a_484_472# net49 0.006499f
C3943 net82 fanout76/a_36_160# 0.001033f
C3944 output46/a_224_472# FILLER_0_20_15/a_572_375# 0.00135f
C3945 FILLER_0_16_89/a_1380_472# _451_/a_1353_112# 0.010457f
C3946 _015_ calibrate 0.105287f
C3947 _069_ _429_/a_1308_423# 0.027468f
C3948 net52 net82 0.108202f
C3949 FILLER_0_4_49/a_484_472# net68 0.027016f
C3950 FILLER_0_21_142/a_36_472# _140_ 0.009261f
C3951 net70 FILLER_0_16_115/a_124_375# 0.025173f
C3952 _321_/a_2034_472# _176_ 0.002722f
C3953 _069_ _395_/a_36_488# 0.042974f
C3954 net82 _443_/a_796_472# 0.00219f
C3955 net50 _439_/a_2665_112# 0.007973f
C3956 net63 output22/a_224_472# 0.017997f
C3957 _095_ FILLER_0_14_107/a_1468_375# 0.010523f
C3958 output32/a_224_472# net32 0.014826f
C3959 FILLER_0_17_104/a_1380_472# vss 0.001141f
C3960 _044_ result[3] 0.00251f
C3961 FILLER_0_5_54/a_1380_472# FILLER_0_6_47/a_2276_472# 0.026657f
C3962 _425_/a_2560_156# net37 0.002508f
C3963 _415_/a_1000_472# net18 0.006558f
C3964 ctln[5] _448_/a_448_472# 0.010887f
C3965 result[7] _419_/a_1000_472# 0.015362f
C3966 _308_/a_124_24# FILLER_0_9_72/a_1468_375# 0.007188f
C3967 _136_ _451_/a_1040_527# 0.00497f
C3968 trimb[1] vdd 0.225206f
C3969 net20 _088_ 0.001704f
C3970 _255_/a_224_552# _070_ 0.001333f
C3971 _141_ _433_/a_2665_112# 0.013144f
C3972 _384_/a_224_472# _168_ 0.003461f
C3973 mask\[8\] _437_/a_1000_472# 0.00112f
C3974 vdd FILLER_0_10_94/a_124_375# 0.020076f
C3975 _422_/a_1000_472# _009_ 0.007191f
C3976 _453_/a_1308_423# vdd 0.002896f
C3977 _453_/a_448_472# vss 0.00396f
C3978 FILLER_0_16_57/a_572_375# net15 0.013085f
C3979 mask\[4\] _201_/a_255_603# 0.002111f
C3980 _328_/a_36_113# _017_ 0.006485f
C3981 mask\[3\] FILLER_0_16_154/a_572_375# 0.027873f
C3982 net65 fanout65/a_36_113# 0.019148f
C3983 net25 _423_/a_2665_112# 0.007096f
C3984 mask\[5\] _108_ 0.036539f
C3985 _429_/a_36_151# FILLER_0_15_212/a_932_472# 0.001723f
C3986 _389_/a_36_148# _171_ 0.023988f
C3987 net36 FILLER_0_18_76/a_484_472# 0.005765f
C3988 net23 _170_ 0.107532f
C3989 _069_ _228_/a_36_68# 0.001676f
C3990 FILLER_0_19_171/a_932_472# vdd 0.011399f
C3991 FILLER_0_19_171/a_484_472# vss 0.001913f
C3992 FILLER_0_20_15/a_1380_472# net40 0.014911f
C3993 _091_ FILLER_0_13_212/a_36_472# 0.007355f
C3994 FILLER_0_14_181/a_124_375# FILLER_0_15_180/a_124_375# 0.026339f
C3995 _161_ _068_ 0.026092f
C3996 FILLER_0_9_223/a_572_375# state\[0\] 0.079258f
C3997 net73 _438_/a_2665_112# 0.001708f
C3998 _031_ vdd 0.327674f
C3999 comp FILLER_0_15_2/a_124_375# 0.034135f
C4000 FILLER_0_13_206/a_124_375# _043_ 0.014212f
C4001 net82 FILLER_0_2_177/a_484_472# 0.001777f
C4002 fanout77/a_36_113# _103_ 0.006045f
C4003 cal_count\[3\] _310_/a_49_472# 0.00277f
C4004 net78 _421_/a_1000_472# 0.022212f
C4005 _438_/a_796_472# vss 0.001171f
C4006 net70 _427_/a_36_151# 0.029237f
C4007 _131_ _058_ 0.031061f
C4008 _114_ _120_ 0.334426f
C4009 _029_ FILLER_0_5_88/a_124_375# 0.006771f
C4010 output13/a_224_472# vss 0.108144f
C4011 FILLER_0_15_142/a_572_375# _427_/a_36_151# 0.059049f
C4012 _017_ net74 0.041246f
C4013 FILLER_0_16_107/a_124_375# _132_ 0.003315f
C4014 FILLER_0_17_72/a_1020_375# _451_/a_3129_107# 0.001202f
C4015 FILLER_0_4_177/a_124_375# net37 0.00459f
C4016 net61 net18 0.71051f
C4017 _126_ _055_ 0.01647f
C4018 FILLER_0_15_282/a_124_375# _006_ 0.002249f
C4019 cal_count\[1\] FILLER_0_15_59/a_484_472# 0.006408f
C4020 FILLER_0_17_200/a_572_375# _093_ 0.002355f
C4021 _132_ FILLER_0_16_115/a_124_375# 0.033245f
C4022 _127_ _118_ 0.141388f
C4023 _077_ net15 0.238832f
C4024 _333_/a_36_160# FILLER_0_15_180/a_36_472# 0.016014f
C4025 FILLER_0_10_37/a_36_472# net51 0.002346f
C4026 FILLER_0_3_204/a_124_375# _088_ 0.00269f
C4027 net55 _012_ 0.060122f
C4028 _322_/a_124_24# vss 0.003731f
C4029 _322_/a_848_380# vdd 0.067623f
C4030 _214_/a_36_160# _098_ 0.001496f
C4031 _450_/a_1353_112# _039_ 0.019843f
C4032 _176_ _389_/a_36_148# 0.060256f
C4033 _008_ _419_/a_1000_472# 0.003267f
C4034 output44/a_224_472# net43 0.001041f
C4035 input1/a_36_113# net18 0.004922f
C4036 net74 _032_ 0.208799f
C4037 fanout69/a_36_113# trim_mask\[4\] 0.027938f
C4038 _074_ FILLER_0_7_233/a_124_375# 0.003081f
C4039 _369_/a_36_68# _156_ 0.001359f
C4040 _449_/a_36_151# FILLER_0_13_72/a_572_375# 0.035849f
C4041 _004_ _416_/a_2248_156# 0.001078f
C4042 mask\[4\] FILLER_0_19_187/a_484_472# 0.004669f
C4043 _431_/a_448_472# net70 0.002293f
C4044 output43/a_224_472# output45/a_224_472# 0.246888f
C4045 trim_val\[4\] _443_/a_2248_156# 0.050943f
C4046 net15 _013_ 0.152142f
C4047 _100_ _099_ 0.03589f
C4048 net57 _427_/a_2248_156# 0.002706f
C4049 net53 _451_/a_836_156# 0.006521f
C4050 mask\[0\] vdd 0.181371f
C4051 _074_ vdd 1.221102f
C4052 net32 vdd 0.50705f
C4053 output42/a_224_472# net47 0.083794f
C4054 net19 _419_/a_2560_156# 0.003213f
C4055 FILLER_0_17_104/a_1020_375# net14 0.002226f
C4056 _128_ net21 0.03068f
C4057 FILLER_0_5_128/a_572_375# net47 0.010055f
C4058 net81 fanout58/a_36_160# 0.005575f
C4059 _086_ FILLER_0_11_142/a_36_472# 0.006774f
C4060 _371_/a_36_113# vdd 0.007666f
C4061 ctln[6] net69 0.003695f
C4062 net81 cal_itt\[0\] 0.001048f
C4063 FILLER_0_3_172/a_1380_472# net22 0.012284f
C4064 _414_/a_36_151# net22 0.014398f
C4065 _434_/a_2560_156# vdd 0.002922f
C4066 _434_/a_2665_112# vss 0.00127f
C4067 FILLER_0_9_28/a_1828_472# net51 0.001502f
C4068 _435_/a_36_151# _434_/a_1308_423# 0.001518f
C4069 FILLER_0_13_142/a_1380_472# vss 0.004953f
C4070 FILLER_0_20_31/a_124_375# FILLER_0_20_15/a_1468_375# 0.012001f
C4071 _417_/a_1000_472# vss 0.001822f
C4072 net62 _417_/a_1308_423# 0.006676f
C4073 result[7] FILLER_0_23_282/a_572_375# 0.015853f
C4074 _074_ FILLER_0_6_177/a_572_375# 0.012642f
C4075 fanout67/a_36_160# net67 0.017633f
C4076 _142_ _093_ 0.492191f
C4077 _275_/a_224_472# net63 0.002538f
C4078 FILLER_0_16_57/a_932_472# FILLER_0_15_59/a_572_375# 0.001543f
C4079 _411_/a_1308_423# net8 0.0176f
C4080 fanout75/a_36_113# _122_ 0.001035f
C4081 _247_/a_36_160# _062_ 0.011327f
C4082 _077_ _133_ 0.003921f
C4083 _127_ _068_ 0.052712f
C4084 _128_ _070_ 1.279188f
C4085 FILLER_0_8_24/a_36_472# net42 0.010665f
C4086 _267_/a_36_472# net23 0.001178f
C4087 net35 FILLER_0_22_177/a_1020_375# 0.008333f
C4088 FILLER_0_22_86/a_1468_375# net71 0.010224f
C4089 result[8] mask\[6\] 0.111221f
C4090 FILLER_0_3_172/a_1020_375# vdd 0.009809f
C4091 _422_/a_2248_156# vdd 0.005833f
C4092 _443_/a_36_151# _370_/a_848_380# 0.001568f
C4093 net47 net51 0.007412f
C4094 net64 net19 0.029763f
C4095 trim_val\[4\] _170_ 0.281942f
C4096 FILLER_0_11_64/a_36_472# _453_/a_36_151# 0.001723f
C4097 FILLER_0_13_212/a_124_375# _043_ 0.011912f
C4098 _093_ FILLER_0_18_107/a_2812_375# 0.00626f
C4099 _095_ _280_/a_224_472# 0.001416f
C4100 input4/a_36_68# net5 0.004765f
C4101 _402_/a_56_567# _452_/a_36_151# 0.001915f
C4102 _096_ _095_ 0.086147f
C4103 _087_ FILLER_0_3_172/a_932_472# 0.001947f
C4104 _431_/a_448_472# _132_ 0.003024f
C4105 net62 FILLER_0_15_282/a_484_472# 0.009524f
C4106 _143_ _340_/a_36_160# 0.001064f
C4107 net75 _074_ 1.343862f
C4108 net66 net49 0.657679f
C4109 _449_/a_36_151# cal_count\[3\] 0.018365f
C4110 _098_ FILLER_0_15_212/a_1020_375# 0.00918f
C4111 FILLER_0_1_192/a_124_375# net11 0.003537f
C4112 net34 _093_ 0.005701f
C4113 _091_ _430_/a_1308_423# 0.023198f
C4114 FILLER_0_15_150/a_36_472# vdd 0.088307f
C4115 net69 _441_/a_2248_156# 0.036635f
C4116 _093_ FILLER_0_16_89/a_1468_375# 0.003988f
C4117 FILLER_0_4_197/a_36_472# _002_ 0.006574f
C4118 _086_ _314_/a_224_472# 0.003715f
C4119 FILLER_0_21_125/a_484_472# _140_ 0.013936f
C4120 net68 net66 0.81104f
C4121 net71 _437_/a_2665_112# 0.039687f
C4122 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_36_472# 0.001723f
C4123 _415_/a_2665_112# vdd 0.017004f
C4124 output31/a_224_472# net18 0.009938f
C4125 net63 FILLER_0_15_212/a_932_472# 0.002269f
C4126 net50 _444_/a_2248_156# 0.005539f
C4127 FILLER_0_0_130/a_124_375# net13 0.009149f
C4128 FILLER_0_3_172/a_2276_472# net21 0.003603f
C4129 FILLER_0_5_109/a_572_375# FILLER_0_5_117/a_124_375# 0.012001f
C4130 _128_ FILLER_0_9_142/a_36_472# 0.005101f
C4131 mask\[9\] FILLER_0_19_111/a_572_375# 0.027695f
C4132 _363_/a_244_472# _053_ 0.001236f
C4133 FILLER_0_20_98/a_124_375# net14 0.05242f
C4134 net20 FILLER_0_6_239/a_124_375# 0.004897f
C4135 FILLER_0_22_86/a_124_375# _026_ 0.001024f
C4136 net52 FILLER_0_5_72/a_1020_375# 0.00799f
C4137 _326_/a_36_160# _128_ 0.02761f
C4138 output10/a_224_472# _411_/a_36_151# 0.001362f
C4139 FILLER_0_4_123/a_124_375# net47 0.011322f
C4140 net79 output30/a_224_472# 0.078502f
C4141 _062_ _134_ 0.024038f
C4142 ctlp[4] _108_ 0.002002f
C4143 _079_ cal_itt\[0\] 0.018495f
C4144 _187_ _120_ 0.144679f
C4145 net57 FILLER_0_3_142/a_36_472# 0.002298f
C4146 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_36_472# 0.001963f
C4147 FILLER_0_2_111/a_1468_375# vdd 0.011806f
C4148 net49 _167_ 0.031111f
C4149 net58 valid 0.149817f
C4150 mask\[3\] net30 0.451388f
C4151 _372_/a_1194_69# _163_ 0.001328f
C4152 net34 output35/a_224_472# 0.0731f
C4153 _085_ _120_ 0.032964f
C4154 _414_/a_448_472# net76 0.002346f
C4155 _412_/a_2665_112# output37/a_224_472# 0.002025f
C4156 _124_ vdd 0.040228f
C4157 FILLER_0_15_142/a_484_472# net23 0.002884f
C4158 net68 _167_ 0.001302f
C4159 FILLER_0_9_60/a_124_375# net51 0.002346f
C4160 FILLER_0_18_107/a_2724_472# vss 0.003148f
C4161 FILLER_0_18_107/a_3172_472# vdd 0.004296f
C4162 _343_/a_49_472# _137_ 0.001419f
C4163 ctlp[1] net78 0.025929f
C4164 net78 _419_/a_796_472# 0.00376f
C4165 _052_ vss 0.077815f
C4166 FILLER_0_4_197/a_932_472# net59 0.003599f
C4167 trimb[1] FILLER_0_18_2/a_572_375# 0.010125f
C4168 FILLER_0_15_142/a_572_375# FILLER_0_15_150/a_124_375# 0.012001f
C4169 FILLER_0_18_100/a_124_375# mask\[9\] 0.005751f
C4170 FILLER_0_5_206/a_124_375# _081_ 0.031751f
C4171 _149_ _437_/a_2248_156# 0.031905f
C4172 _026_ _437_/a_1000_472# 0.042316f
C4173 net63 FILLER_0_20_177/a_1020_375# 0.005919f
C4174 net67 FILLER_0_12_20/a_36_472# 0.054453f
C4175 _086_ _321_/a_170_472# 0.046783f
C4176 _092_ _105_ 0.006701f
C4177 _256_/a_1612_497# _077_ 0.002724f
C4178 net34 _435_/a_796_472# 0.002288f
C4179 FILLER_0_17_56/a_572_375# FILLER_0_18_61/a_36_472# 0.001597f
C4180 _088_ vss 0.326434f
C4181 _093_ FILLER_0_17_72/a_1020_375# 0.001994f
C4182 mask\[0\] FILLER_0_13_206/a_36_472# 0.012766f
C4183 FILLER_0_13_142/a_484_472# net23 0.006746f
C4184 net69 _154_ 0.05211f
C4185 fanout55/a_36_160# _095_ 0.00409f
C4186 mask\[4\] FILLER_0_19_155/a_572_375# 0.020261f
C4187 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_36_472# 0.086635f
C4188 net47 net6 0.23883f
C4189 _155_ FILLER_0_4_107/a_124_375# 0.00162f
C4190 net81 _429_/a_36_151# 0.018551f
C4191 _072_ _163_ 0.016226f
C4192 output12/a_224_472# FILLER_0_0_198/a_36_472# 0.023414f
C4193 _441_/a_36_151# _168_ 0.033578f
C4194 _053_ _129_ 0.003479f
C4195 _053_ _372_/a_2034_472# 0.00181f
C4196 _045_ _006_ 0.00216f
C4197 fanout68/a_36_113# FILLER_0_3_54/a_124_375# 0.015816f
C4198 _063_ trim_val\[0\] 0.001978f
C4199 _119_ FILLER_0_4_107/a_1468_375# 0.001695f
C4200 _095_ _401_/a_36_68# 0.001398f
C4201 result[6] net77 0.111093f
C4202 net58 net9 0.018829f
C4203 net27 _323_/a_36_113# 0.010949f
C4204 _096_ mask\[1\] 0.010488f
C4205 _098_ FILLER_0_19_171/a_124_375# 0.040575f
C4206 net63 _137_ 0.006317f
C4207 fanout61/a_36_113# net77 0.052643f
C4208 _142_ FILLER_0_17_142/a_36_472# 0.011216f
C4209 FILLER_0_16_89/a_124_375# net36 0.011956f
C4210 trim_mask\[4\] _066_ 0.396509f
C4211 FILLER_0_18_107/a_3260_375# _145_ 0.00346f
C4212 net75 _411_/a_1204_472# 0.008304f
C4213 FILLER_0_5_109/a_124_375# net47 0.010784f
C4214 _098_ FILLER_0_15_235/a_124_375# 0.012702f
C4215 _413_/a_36_151# net65 0.033028f
C4216 FILLER_0_4_144/a_36_472# vdd 0.004289f
C4217 FILLER_0_4_144/a_572_375# vss 0.072463f
C4218 FILLER_0_22_177/a_36_472# _146_ 0.002f
C4219 net47 _163_ 0.64626f
C4220 result[9] _419_/a_1204_472# 0.019627f
C4221 FILLER_0_18_171/a_36_472# _098_ 0.020038f
C4222 FILLER_0_2_111/a_124_375# _369_/a_36_68# 0.001176f
C4223 ctln[5] vdd 0.256793f
C4224 _256_/a_36_68# net22 0.019035f
C4225 _449_/a_2560_156# vss 0.002544f
C4226 _093_ mask\[2\] 0.009354f
C4227 mask\[9\] vss 0.649041f
C4228 _136_ _139_ 0.394888f
C4229 cal_itt\[2\] _253_/a_672_68# 0.0016f
C4230 _429_/a_1308_423# net22 0.001856f
C4231 _414_/a_2248_156# _074_ 0.013023f
C4232 net73 _431_/a_1204_472# 0.026905f
C4233 net52 FILLER_0_5_54/a_1468_375# 0.003649f
C4234 FILLER_0_22_128/a_36_472# _022_ 0.001541f
C4235 _139_ net21 0.004991f
C4236 net15 _110_ 0.016359f
C4237 net17 _452_/a_448_472# 0.043154f
C4238 FILLER_0_17_72/a_932_472# vss 0.002754f
C4239 FILLER_0_17_72/a_1380_472# vdd 0.001762f
C4240 net27 FILLER_0_14_235/a_484_472# 0.010072f
C4241 _228_/a_36_68# _090_ 0.018462f
C4242 FILLER_0_4_49/a_484_472# net47 0.002964f
C4243 vss rstn 0.149553f
C4244 _076_ FILLER_0_5_148/a_36_472# 0.011563f
C4245 _098_ FILLER_0_20_98/a_124_375# 0.012779f
C4246 _053_ FILLER_0_5_54/a_36_472# 0.003309f
C4247 _413_/a_36_151# net59 0.02781f
C4248 _068_ _246_/a_36_68# 0.059106f
C4249 net60 _421_/a_1000_472# 0.035511f
C4250 _363_/a_244_472# _028_ 0.002693f
C4251 _418_/a_1000_472# vss 0.001193f
C4252 _430_/a_1204_472# net21 0.006991f
C4253 output27/a_224_472# calibrate 0.010614f
C4254 net15 _423_/a_448_472# 0.004833f
C4255 _422_/a_1204_472# mask\[7\] 0.025592f
C4256 _426_/a_2665_112# _055_ 0.00142f
C4257 _449_/a_36_151# _394_/a_1336_472# 0.001582f
C4258 net52 _443_/a_2665_112# 0.05031f
C4259 _074_ _374_/a_36_68# 0.001447f
C4260 net57 _428_/a_1308_423# 0.018725f
C4261 _091_ FILLER_0_15_212/a_1468_375# 0.002531f
C4262 trim[1] _033_ 0.015549f
C4263 net61 _422_/a_448_472# 0.006042f
C4264 cal_count\[2\] FILLER_0_15_2/a_484_472# 0.015036f
C4265 output7/a_224_472# net40 0.009154f
C4266 FILLER_0_0_198/a_124_375# net11 0.071885f
C4267 _426_/a_1204_472# calibrate 0.00182f
C4268 FILLER_0_18_107/a_484_472# net14 0.002472f
C4269 net20 _260_/a_36_68# 0.033776f
C4270 net31 ctlp[1] 0.050993f
C4271 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_36_472# 0.002765f
C4272 _228_/a_36_68# net22 0.052558f
C4273 _055_ _060_ 0.181186f
C4274 FILLER_0_4_213/a_124_375# net59 0.039014f
C4275 _118_ net23 0.108864f
C4276 net82 _152_ 0.001896f
C4277 _453_/a_2665_112# net51 0.046426f
C4278 net56 _427_/a_2665_112# 0.012193f
C4279 ctln[2] net65 0.113266f
C4280 _276_/a_36_160# _093_ 0.019339f
C4281 FILLER_0_16_89/a_932_472# net14 0.014714f
C4282 _028_ FILLER_0_5_72/a_1468_375# 0.00123f
C4283 _428_/a_36_151# _043_ 0.027757f
C4284 FILLER_0_17_200/a_484_472# net21 0.017997f
C4285 FILLER_0_7_195/a_124_375# _072_ 0.012244f
C4286 net17 FILLER_0_12_28/a_36_472# 0.012286f
C4287 FILLER_0_4_107/a_932_472# net47 0.008252f
C4288 FILLER_0_12_20/a_572_375# net47 0.00139f
C4289 _052_ _424_/a_448_472# 0.017551f
C4290 _078_ FILLER_0_3_221/a_124_375# 0.002694f
C4291 _098_ _434_/a_1308_423# 0.007057f
C4292 net27 FILLER_0_8_263/a_36_472# 0.003956f
C4293 _030_ _164_ 0.036025f
C4294 _449_/a_2248_156# net55 0.052445f
C4295 _114_ _043_ 0.071339f
C4296 net28 _005_ 0.080653f
C4297 net15 _447_/a_2248_156# 0.01843f
C4298 FILLER_0_8_239/a_36_472# _123_ 0.011767f
C4299 mask\[3\] FILLER_0_18_177/a_572_375# 0.002924f
C4300 FILLER_0_4_177/a_36_472# trim_val\[4\] 0.001889f
C4301 _053_ net57 0.037224f
C4302 FILLER_0_16_255/a_36_472# vdd 0.044615f
C4303 net63 _434_/a_2248_156# 0.063346f
C4304 _136_ net14 0.417108f
C4305 calibrate net22 0.036525f
C4306 _440_/a_1308_423# vss 0.028595f
C4307 net55 FILLER_0_17_72/a_36_472# 0.020422f
C4308 _446_/a_2665_112# net49 0.006979f
C4309 output29/a_224_472# output30/a_224_472# 0.005147f
C4310 _064_ _035_ 0.02225f
C4311 net18 net8 0.072251f
C4312 _053_ _219_/a_36_160# 0.005244f
C4313 net54 _210_/a_67_603# 0.001108f
C4314 _432_/a_36_151# _137_ 0.051293f
C4315 FILLER_0_18_171/a_124_375# _432_/a_36_151# 0.001597f
C4316 FILLER_0_20_87/a_124_375# _437_/a_36_151# 0.059049f
C4317 ctln[2] net59 0.009218f
C4318 net67 trim_mask\[1\] 0.01761f
C4319 _256_/a_36_68# _076_ 0.079206f
C4320 FILLER_0_21_133/a_36_472# _436_/a_2248_156# 0.001148f
C4321 _443_/a_1000_472# _170_ 0.012879f
C4322 _056_ _113_ 0.052362f
C4323 net1 _265_/a_468_472# 0.002612f
C4324 FILLER_0_12_124/a_36_472# _131_ 0.028609f
C4325 FILLER_0_19_47/a_124_375# vdd 0.025971f
C4326 FILLER_0_16_107/a_124_375# vdd 0.026251f
C4327 _035_ output41/a_224_472# 0.002168f
C4328 net76 FILLER_0_3_172/a_1916_375# 0.019901f
C4329 _131_ FILLER_0_17_104/a_1020_375# 0.006574f
C4330 net36 _437_/a_36_151# 0.002694f
C4331 vdd FILLER_0_16_115/a_124_375# 0.020393f
C4332 result[9] FILLER_0_23_282/a_36_472# 0.001324f
C4333 FILLER_0_6_47/a_932_472# vdd 0.003435f
C4334 _070_ net14 0.536953f
C4335 output37/a_224_472# en 0.003788f
C4336 _444_/a_2248_156# _054_ 0.002637f
C4337 FILLER_0_21_206/a_124_375# _205_/a_36_160# 0.03126f
C4338 _356_/a_36_472# net14 0.001801f
C4339 net35 vss 0.434438f
C4340 net82 net21 0.037271f
C4341 _062_ _311_/a_66_473# 0.027039f
C4342 _068_ net23 0.432092f
C4343 FILLER_0_6_239/a_124_375# vss 0.017355f
C4344 FILLER_0_6_239/a_36_472# vdd 0.092399f
C4345 net65 FILLER_0_3_221/a_1468_375# 0.001695f
C4346 fanout68/a_36_113# vss 0.006152f
C4347 _422_/a_2560_156# _108_ 0.008253f
C4348 FILLER_0_18_177/a_1828_472# FILLER_0_19_187/a_572_375# 0.001684f
C4349 _177_ net36 0.371814f
C4350 _081_ FILLER_0_5_136/a_36_472# 0.0028f
C4351 _152_ FILLER_0_5_136/a_124_375# 0.039558f
C4352 FILLER_0_14_81/a_36_472# vss 0.007047f
C4353 _088_ net4 0.096522f
C4354 output31/a_224_472# _417_/a_36_151# 0.07368f
C4355 net41 net67 0.03408f
C4356 _103_ net19 0.047895f
C4357 FILLER_0_21_206/a_124_375# mask\[6\] 0.008881f
C4358 fanout55/a_36_160# net74 0.016856f
C4359 FILLER_0_22_86/a_1020_375# net14 0.047331f
C4360 _091_ FILLER_0_19_171/a_572_375# 0.013568f
C4361 FILLER_0_5_212/a_124_375# _078_ 0.002018f
C4362 _065_ vdd 0.646511f
C4363 _431_/a_2665_112# FILLER_0_17_142/a_124_375# 0.004834f
C4364 _448_/a_1308_423# net59 0.014899f
C4365 _105_ vdd 0.565719f
C4366 _056_ _118_ 0.028015f
C4367 _095_ _055_ 0.002933f
C4368 _023_ _146_ 0.006636f
C4369 FILLER_0_9_28/a_1916_375# vdd 0.01295f
C4370 _069_ FILLER_0_15_212/a_36_472# 0.046864f
C4371 FILLER_0_0_96/a_124_375# vss 0.008342f
C4372 FILLER_0_0_96/a_36_472# vdd 0.047982f
C4373 net58 _084_ 0.141836f
C4374 _427_/a_36_151# vdd 0.107344f
C4375 FILLER_0_21_142/a_36_472# _098_ 0.002964f
C4376 _287_/a_36_472# _006_ 0.00121f
C4377 fanout55/a_36_160# cal_count\[1\] 0.007256f
C4378 net20 net65 0.335083f
C4379 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_36_472# 0.086635f
C4380 _408_/a_1936_472# _067_ 0.003007f
C4381 _093_ FILLER_0_18_177/a_2364_375# 0.001989f
C4382 _155_ _153_ 0.033366f
C4383 FILLER_0_9_223/a_124_375# vss 0.009569f
C4384 net20 _093_ 0.398457f
C4385 _127_ FILLER_0_11_142/a_36_472# 0.004538f
C4386 _401_/a_36_68# cal_count\[1\] 0.006747f
C4387 _095_ FILLER_0_15_10/a_124_375# 0.023187f
C4388 vdd FILLER_0_8_156/a_124_375# 0.005213f
C4389 _076_ calibrate 1.005804f
C4390 ctlp[6] net23 0.006951f
C4391 net15 FILLER_0_17_56/a_572_375# 0.007386f
C4392 _437_/a_2248_156# net14 0.023718f
C4393 _002_ FILLER_0_3_172/a_2364_375# 0.016984f
C4394 net81 _415_/a_448_472# 0.004045f
C4395 _430_/a_2665_112# FILLER_0_15_212/a_1380_472# 0.021761f
C4396 FILLER_0_15_142/a_124_375# _095_ 0.003935f
C4397 net75 FILLER_0_6_239/a_36_472# 0.009325f
C4398 _057_ vss 0.169369f
C4399 mask\[9\] _148_ 0.01635f
C4400 _180_ vdd 0.176915f
C4401 _429_/a_36_151# mask\[1\] 0.001021f
C4402 FILLER_0_17_38/a_36_472# _041_ 0.003805f
C4403 _126_ _172_ 0.017618f
C4404 _327_/a_36_472# net74 0.009344f
C4405 _142_ FILLER_0_16_154/a_124_375# 0.004001f
C4406 fanout51/a_36_113# vdd 0.013496f
C4407 _113_ FILLER_0_12_196/a_124_375# 0.001597f
C4408 _090_ FILLER_0_12_196/a_36_472# 0.002321f
C4409 FILLER_0_22_177/a_484_472# _435_/a_36_151# 0.001723f
C4410 _114_ FILLER_0_10_94/a_572_375# 0.008375f
C4411 _033_ _444_/a_448_472# 0.047424f
C4412 FILLER_0_12_136/a_484_472# cal_count\[3\] 0.007275f
C4413 _086_ _135_ 0.005637f
C4414 net66 net47 0.238874f
C4415 _068_ _311_/a_1660_473# 0.003542f
C4416 FILLER_0_19_125/a_124_375# vss 0.001974f
C4417 fanout71/a_36_113# net71 0.087994f
C4418 _443_/a_36_151# FILLER_0_2_127/a_124_375# 0.073306f
C4419 FILLER_0_15_205/a_124_375# net21 0.002912f
C4420 _427_/a_2665_112# _095_ 0.039612f
C4421 _258_/a_36_160# FILLER_0_7_233/a_124_375# 0.001633f
C4422 _431_/a_448_472# vdd 0.001932f
C4423 net20 net59 0.045227f
C4424 FILLER_0_9_28/a_484_472# _054_ 0.002831f
C4425 FILLER_0_5_198/a_484_472# net22 0.012457f
C4426 _068_ _313_/a_255_603# 0.001149f
C4427 _136_ _098_ 0.049635f
C4428 _451_/a_2225_156# vdd 0.012404f
C4429 _451_/a_3129_107# vss 0.01f
C4430 net65 FILLER_0_1_266/a_484_472# 0.004635f
C4431 output42/a_224_472# vdd 0.04917f
C4432 net61 _418_/a_36_151# 0.042401f
C4433 FILLER_0_5_128/a_572_375# vdd 0.008326f
C4434 _420_/a_36_151# FILLER_0_23_274/a_36_472# 0.001723f
C4435 _098_ net21 0.133694f
C4436 FILLER_0_3_54/a_124_375# net40 0.005766f
C4437 net60 ctlp[1] 0.073021f
C4438 net60 _419_/a_796_472# 0.003097f
C4439 net61 _419_/a_1204_472# 0.012025f
C4440 FILLER_0_3_204/a_124_375# net65 0.003831f
C4441 net52 net69 0.372114f
C4442 _412_/a_1308_423# vdd 0.003842f
C4443 _305_/a_36_159# _112_ 0.001664f
C4444 _258_/a_36_160# vdd 0.00617f
C4445 net82 FILLER_0_4_213/a_484_472# 0.002255f
C4446 net57 FILLER_0_5_164/a_36_472# 0.032208f
C4447 _056_ _068_ 0.127175f
C4448 comp _043_ 0.003867f
C4449 FILLER_0_12_124/a_36_472# _126_ 0.056268f
C4450 _032_ _442_/a_448_472# 0.001977f
C4451 _443_/a_448_472# _031_ 0.001143f
C4452 _443_/a_796_472# net69 0.020234f
C4453 ctln[0] output41/a_224_472# 0.001583f
C4454 _070_ FILLER_0_5_136/a_124_375# 0.001083f
C4455 _187_ _043_ 0.011995f
C4456 _280_/a_224_472# _097_ 0.007508f
C4457 _096_ _097_ 0.038778f
C4458 FILLER_0_18_177/a_2724_472# vdd 0.002749f
C4459 _077_ net37 0.003374f
C4460 FILLER_0_12_28/a_36_472# _039_ 0.007926f
C4461 result[7] net77 0.005269f
C4462 _044_ FILLER_0_13_290/a_36_472# 0.001194f
C4463 net35 FILLER_0_22_128/a_1020_375# 0.010202f
C4464 mask\[0\] _099_ 0.00418f
C4465 net47 _167_ 0.003019f
C4466 trimb[2] vss 0.102375f
C4467 FILLER_0_4_49/a_572_375# FILLER_0_3_54/a_36_472# 0.001597f
C4468 net16 _064_ 0.121797f
C4469 _079_ FILLER_0_5_198/a_572_375# 0.011369f
C4470 _088_ FILLER_0_5_198/a_124_375# 0.001374f
C4471 net50 _054_ 0.131493f
C4472 net64 _055_ 0.00384f
C4473 _289_/a_244_68# _103_ 0.001153f
C4474 _067_ net47 0.0609f
C4475 _308_/a_848_380# _134_ 0.001299f
C4476 _042_ vss 0.008272f
C4477 net51 vdd 0.692054f
C4478 vdd FILLER_0_13_72/a_36_472# 0.108152f
C4479 vss FILLER_0_13_72/a_572_375# 0.061657f
C4480 net16 _447_/a_1204_472# 0.00194f
C4481 net72 _180_ 0.040135f
C4482 FILLER_0_16_57/a_484_472# vss 0.004107f
C4483 FILLER_0_16_57/a_932_472# vdd 0.005518f
C4484 FILLER_0_3_204/a_124_375# net59 0.007104f
C4485 _018_ _043_ 0.0022f
C4486 FILLER_0_18_107/a_3172_472# FILLER_0_19_134/a_124_375# 0.001723f
C4487 net70 FILLER_0_14_99/a_124_375# 0.002922f
C4488 _114_ FILLER_0_12_136/a_124_375# 0.006974f
C4489 fanout68/a_36_113# trim_mask\[2\] 0.003509f
C4490 _164_ trim_mask\[3\] 0.016366f
C4491 net38 output6/a_224_472# 0.060017f
C4492 _260_/a_36_68# vss 0.030324f
C4493 output7/a_224_472# trim[3] 0.103375f
C4494 result[7] FILLER_0_23_290/a_36_472# 0.013403f
C4495 net67 _164_ 0.030648f
C4496 _186_ _181_ 0.018817f
C4497 _444_/a_36_151# net17 0.001435f
C4498 _219_/a_36_160# trim_mask\[0\] 0.395762f
C4499 _076_ _125_ 0.009254f
C4500 FILLER_0_2_93/a_36_472# net14 0.005108f
C4501 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_484_472# 0.013276f
C4502 _071_ _314_/a_224_472# 0.001359f
C4503 _352_/a_49_472# mask\[7\] 0.001066f
C4504 FILLER_0_1_98/a_36_472# FILLER_0_0_96/a_124_375# 0.001684f
C4505 _065_ _447_/a_448_472# 0.049072f
C4506 _066_ net37 0.006164f
C4507 FILLER_0_12_2/a_36_472# clkc 0.004826f
C4508 vdd _047_ 0.175913f
C4509 _093_ FILLER_0_19_111/a_572_375# 0.002743f
C4510 _073_ FILLER_0_3_221/a_1020_375# 0.002563f
C4511 _140_ FILLER_0_19_155/a_572_375# 0.040109f
C4512 _095_ _278_/a_36_160# 0.030448f
C4513 _148_ _352_/a_49_472# 0.003082f
C4514 net35 mask\[7\] 0.954332f
C4515 output27/a_224_472# FILLER_0_9_270/a_572_375# 0.00135f
C4516 _446_/a_448_472# _035_ 0.018273f
C4517 FILLER_0_14_50/a_124_375# _401_/a_36_68# 0.001129f
C4518 net31 _201_/a_67_603# 0.015773f
C4519 _127_ _321_/a_170_472# 0.023836f
C4520 _372_/a_170_472# _152_ 0.037088f
C4521 _131_ _152_ 0.002949f
C4522 FILLER_0_4_123/a_124_375# vdd 0.027816f
C4523 net35 _148_ 0.114816f
C4524 _214_/a_36_160# _213_/a_67_603# 0.002505f
C4525 _015_ _426_/a_1204_472# 0.008883f
C4526 FILLER_0_7_72/a_1380_472# vss 0.001117f
C4527 _008_ net77 0.029049f
C4528 _386_/a_124_24# _169_ 0.02709f
C4529 _176_ FILLER_0_10_107/a_36_472# 0.009019f
C4530 net63 result[8] 0.013631f
C4531 _098_ _437_/a_2248_156# 0.008669f
C4532 FILLER_0_14_50/a_36_472# vss 0.002954f
C4533 trimb[1] net44 0.089379f
C4534 output9/a_224_472# ctln[2] 0.080206f
C4535 net65 FILLER_0_3_172/a_36_472# 0.014671f
C4536 FILLER_0_7_104/a_1380_472# _131_ 0.043557f
C4537 input4/a_36_68# en 0.064323f
C4538 FILLER_0_9_72/a_1020_375# vdd -0.014642f
C4539 FILLER_0_9_72/a_572_375# vss 0.007993f
C4540 FILLER_0_4_144/a_36_472# FILLER_0_3_142/a_124_375# 0.001543f
C4541 net27 _426_/a_36_151# 0.008613f
C4542 _163_ _385_/a_36_68# 0.012699f
C4543 _451_/a_448_472# net14 0.04399f
C4544 _072_ _121_ 0.041039f
C4545 net81 fanout76/a_36_160# 0.041089f
C4546 FILLER_0_16_57/a_1468_375# net55 0.006307f
C4547 FILLER_0_16_57/a_932_472# net72 0.004262f
C4548 _093_ FILLER_0_18_100/a_124_375# 0.011632f
C4549 FILLER_0_5_128/a_36_472# _360_/a_36_160# 0.195479f
C4550 output8/a_224_472# FILLER_0_3_221/a_572_375# 0.03228f
C4551 FILLER_0_4_185/a_124_375# net76 0.053929f
C4552 _173_ FILLER_0_12_28/a_124_375# 0.009218f
C4553 FILLER_0_15_150/a_124_375# vdd 0.026143f
C4554 _132_ net54 0.016007f
C4555 net63 net64 0.002181f
C4556 cal_count\[3\] vss 1.35143f
C4557 _147_ _023_ 0.004036f
C4558 valid net82 0.060784f
C4559 net67 FILLER_0_8_24/a_36_472# 0.001252f
C4560 net57 FILLER_0_13_142/a_572_375# 0.011369f
C4561 net18 _417_/a_1308_423# 0.015651f
C4562 net20 _429_/a_2665_112# 0.062922f
C4563 FILLER_0_12_236/a_484_472# vss 0.002739f
C4564 FILLER_0_16_89/a_932_472# _131_ 0.008223f
C4565 net15 _160_ 0.046497f
C4566 FILLER_0_21_206/a_36_472# vss 0.004971f
C4567 net63 mask\[1\] 0.120872f
C4568 FILLER_0_21_125/a_484_472# _098_ 0.002964f
C4569 fanout66/a_36_113# net66 0.032757f
C4570 net82 FILLER_0_3_221/a_932_472# 0.004092f
C4571 _086_ _129_ 0.051553f
C4572 vss _416_/a_36_151# 0.044403f
C4573 output21/a_224_472# result[8] 0.149245f
C4574 FILLER_0_7_72/a_3172_472# _077_ 0.001923f
C4575 vdd net6 0.134918f
C4576 _137_ FILLER_0_17_104/a_1020_375# 0.001676f
C4577 net65 cal_itt\[1\] 0.049124f
C4578 mask\[2\] FILLER_0_16_154/a_124_375# 0.087247f
C4579 _110_ net71 0.004816f
C4580 net62 net78 0.001947f
C4581 _035_ _166_ 0.034749f
C4582 net68 _232_/a_67_603# 0.00184f
C4583 _094_ mask\[2\] 0.089828f
C4584 fanout82/a_36_113# output48/a_224_472# 0.009784f
C4585 output48/a_224_472# _425_/a_448_472# 0.001155f
C4586 FILLER_0_9_223/a_124_375# net4 0.061757f
C4587 _140_ FILLER_0_22_128/a_2364_375# 0.003037f
C4588 _131_ _136_ 1.42765f
C4589 _176_ FILLER_0_10_94/a_124_375# 0.009888f
C4590 _370_/a_692_472# net47 0.001021f
C4591 _119_ _129_ 0.055585f
C4592 FILLER_0_15_142/a_124_375# net74 0.005931f
C4593 net58 calibrate 0.205792f
C4594 output8/a_224_472# _000_ 0.182377f
C4595 net48 _123_ 0.153061f
C4596 _021_ _098_ 0.014179f
C4597 _432_/a_1308_423# _091_ 0.008903f
C4598 FILLER_0_15_282/a_484_472# net18 0.018113f
C4599 _337_/a_665_69# mask\[1\] 0.002125f
C4600 net74 _154_ 0.002976f
C4601 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_36_472# 0.001723f
C4602 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_572_375# 0.026339f
C4603 net65 sample 0.148853f
C4604 mask\[3\] _143_ 0.023322f
C4605 vss net40 0.898805f
C4606 FILLER_0_5_109/a_124_375# vdd 0.060786f
C4607 net23 _146_ 0.034955f
C4608 FILLER_0_21_28/a_1380_472# vdd 0.007073f
C4609 _169_ vss 0.037006f
C4610 _163_ vdd 0.418075f
C4611 net35 _436_/a_1308_423# 0.008773f
C4612 _057_ _311_/a_692_473# 0.002083f
C4613 FILLER_0_18_171/a_124_375# FILLER_0_19_171/a_124_375# 0.05841f
C4614 _032_ _370_/a_124_24# 0.007035f
C4615 net82 net9 0.004599f
C4616 net15 FILLER_0_5_54/a_1020_375# 0.015944f
C4617 net65 vss 0.471168f
C4618 _114_ _062_ 0.028432f
C4619 FILLER_0_22_128/a_2364_375# FILLER_0_21_150/a_36_472# 0.001543f
C4620 net52 FILLER_0_2_111/a_572_375# 0.00245f
C4621 cal_itt\[2\] FILLER_0_3_221/a_1020_375# 0.010951f
C4622 _372_/a_170_472# _070_ 0.024545f
C4623 _131_ _070_ 0.161861f
C4624 _069_ _090_ 1.067281f
C4625 fanout62/a_36_160# FILLER_0_11_282/a_124_375# 0.058702f
C4626 result[5] net62 0.041722f
C4627 cal_itt\[1\] net59 0.227495f
C4628 _115_ vdd 0.455713f
C4629 _093_ vss 2.002012f
C4630 net68 _453_/a_1000_472# 0.001816f
C4631 result[2] FILLER_0_15_282/a_124_375# 0.001114f
C4632 FILLER_0_18_2/a_1828_472# net17 0.008573f
C4633 cal_itt\[3\] net57 0.001586f
C4634 _256_/a_36_68# _128_ 0.001702f
C4635 FILLER_0_4_107/a_572_375# _157_ 0.001032f
C4636 _173_ _039_ 0.0326f
C4637 FILLER_0_21_133/a_124_375# net54 0.013027f
C4638 _415_/a_448_472# net64 0.02484f
C4639 net57 FILLER_0_16_154/a_1380_472# 0.041458f
C4640 FILLER_0_7_72/a_36_472# net52 0.014911f
C4641 FILLER_0_6_177/a_572_375# _163_ 0.001839f
C4642 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_36_472# 0.007947f
C4643 _415_/a_36_151# FILLER_0_11_282/a_124_375# 0.001822f
C4644 FILLER_0_20_107/a_36_472# net71 0.004375f
C4645 FILLER_0_17_72/a_2364_375# _131_ 0.006037f
C4646 _133_ _160_ 0.043549f
C4647 FILLER_0_4_49/a_484_472# vdd 0.003356f
C4648 FILLER_0_4_49/a_36_472# vss 0.001931f
C4649 net57 _081_ 0.023513f
C4650 net37 FILLER_0_5_148/a_484_472# 0.001212f
C4651 FILLER_0_11_109/a_36_472# _135_ 0.001891f
C4652 FILLER_0_19_195/a_124_375# FILLER_0_19_187/a_572_375# 0.012001f
C4653 net81 FILLER_0_15_212/a_1020_375# 0.006974f
C4654 net65 FILLER_0_2_171/a_124_375# 0.023202f
C4655 FILLER_0_5_72/a_932_472# net47 0.003953f
C4656 sample net59 0.001181f
C4657 FILLER_0_7_72/a_2812_375# vdd 0.02125f
C4658 mask\[4\] _069_ 0.001182f
C4659 _069_ net22 0.327999f
C4660 net80 FILLER_0_20_169/a_124_375# 0.054969f
C4661 FILLER_0_15_180/a_572_375# vss 0.010974f
C4662 FILLER_0_15_180/a_36_472# vdd 0.017678f
C4663 output45/a_224_472# net45 0.019483f
C4664 FILLER_0_24_290/a_36_472# FILLER_0_23_290/a_36_472# 0.05841f
C4665 net59 vss 1.191297f
C4666 _415_/a_2248_156# vdd 0.009114f
C4667 FILLER_0_20_177/a_36_472# _434_/a_36_151# 0.001723f
C4668 FILLER_0_20_177/a_1468_375# _434_/a_448_472# 0.008952f
C4669 _111_ FILLER_0_18_76/a_124_375# 0.002494f
C4670 _428_/a_796_472# _095_ 0.00117f
C4671 trim_val\[1\] trim_mask\[1\] 0.519723f
C4672 _340_/a_36_160# FILLER_0_20_169/a_36_472# 0.195478f
C4673 _155_ net50 0.012085f
C4674 _408_/a_244_524# net47 0.001066f
C4675 _000_ _253_/a_36_68# 0.005121f
C4676 net16 _174_ 0.022224f
C4677 output35/a_224_472# vss 0.01667f
C4678 net51 cal_count\[0\] 0.030963f
C4679 net74 _058_ 0.026905f
C4680 _430_/a_448_472# net36 0.011598f
C4681 FILLER_0_3_78/a_484_472# vss 0.005811f
C4682 net39 _444_/a_36_151# 0.14155f
C4683 _074_ FILLER_0_5_164/a_572_375# 0.001307f
C4684 net72 FILLER_0_21_28/a_1380_472# 0.048287f
C4685 _452_/a_836_156# net40 0.023204f
C4686 _095_ FILLER_0_15_72/a_572_375# 0.00352f
C4687 net16 _444_/a_2248_156# 0.065914f
C4688 _326_/a_36_160# _131_ 0.023688f
C4689 FILLER_0_11_142/a_36_472# net23 0.002015f
C4690 _432_/a_36_151# mask\[1\] 0.003001f
C4691 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_36_472# 0.026657f
C4692 _077_ _439_/a_2560_156# 0.012523f
C4693 net46 FILLER_0_21_28/a_124_375# 0.011995f
C4694 FILLER_0_4_107/a_932_472# vdd 0.00987f
C4695 net65 FILLER_0_2_165/a_124_375# 0.001177f
C4696 FILLER_0_2_171/a_124_375# net59 0.006603f
C4697 FILLER_0_8_24/a_572_375# net47 0.0353f
C4698 net67 _450_/a_1353_112# 0.025358f
C4699 FILLER_0_12_20/a_572_375# vdd 0.013384f
C4700 _149_ FILLER_0_20_107/a_124_375# 0.001244f
C4701 _086_ net57 0.126563f
C4702 _411_/a_36_151# net10 0.127193f
C4703 FILLER_0_15_212/a_36_472# net22 0.003143f
C4704 _435_/a_1000_472# vdd 0.032539f
C4705 FILLER_0_17_226/a_36_472# vss 0.007552f
C4706 net33 _146_ 0.306187f
C4707 FILLER_0_9_72/a_484_472# _439_/a_36_151# 0.001723f
C4708 FILLER_0_11_64/a_124_375# cal_count\[3\] 0.002495f
C4709 FILLER_0_4_144/a_484_472# _443_/a_36_151# 0.002841f
C4710 vdd FILLER_0_6_231/a_124_375# 0.024542f
C4711 _431_/a_1000_472# _136_ 0.024253f
C4712 _411_/a_36_151# FILLER_0_0_232/a_124_375# 0.059049f
C4713 output9/a_224_472# FILLER_0_1_266/a_484_472# 0.0323f
C4714 net41 trim_val\[1\] 0.001912f
C4715 _074_ _251_/a_1130_472# 0.00237f
C4716 _119_ net57 0.30462f
C4717 net55 FILLER_0_17_64/a_36_472# 0.034504f
C4718 _077_ _122_ 0.144611f
C4719 _164_ _382_/a_224_472# 0.011658f
C4720 FILLER_0_7_195/a_124_375# vdd 0.007788f
C4721 _128_ calibrate 0.039365f
C4722 _141_ net35 0.003655f
C4723 vss FILLER_0_21_60/a_484_472# 0.004134f
C4724 result[4] _417_/a_2560_156# 0.001076f
C4725 FILLER_0_19_171/a_932_472# _434_/a_36_151# 0.00271f
C4726 _451_/a_1040_527# _040_ 0.007154f
C4727 _126_ _136_ 0.086459f
C4728 net63 FILLER_0_18_177/a_1828_472# 0.047684f
C4729 _091_ _430_/a_1000_472# 0.025041f
C4730 _394_/a_728_93# vdd 0.006211f
C4731 net31 _199_/a_36_160# 0.007888f
C4732 _394_/a_1336_472# vss 0.040135f
C4733 _126_ net21 0.024842f
C4734 net48 _305_/a_36_159# 0.059079f
C4735 trim_mask\[4\] _160_ 0.244284f
C4736 FILLER_0_2_165/a_124_375# net59 0.00999f
C4737 FILLER_0_19_28/a_124_375# vdd 0.028695f
C4738 FILLER_0_16_57/a_572_375# FILLER_0_17_56/a_572_375# 0.026339f
C4739 _002_ net76 0.213703f
C4740 FILLER_0_10_78/a_932_472# FILLER_0_9_72/a_1468_375# 0.001543f
C4741 FILLER_0_18_177/a_2812_375# _202_/a_36_160# 0.026361f
C4742 _050_ FILLER_0_22_128/a_124_375# 0.002607f
C4743 output38/a_224_472# net66 0.148811f
C4744 FILLER_0_10_256/a_124_375# net28 0.034928f
C4745 FILLER_0_15_2/a_572_375# vdd 0.017581f
C4746 FILLER_0_15_2/a_124_375# vss 0.002713f
C4747 _428_/a_2560_156# net53 0.002265f
C4748 fanout71/a_36_113# FILLER_0_20_107/a_36_472# 0.001645f
C4749 FILLER_0_21_28/a_1380_472# _424_/a_36_151# 0.001723f
C4750 _314_/a_224_472# net23 0.001238f
C4751 trim_mask\[2\] net40 0.401672f
C4752 _069_ _076_ 0.033276f
C4753 _126_ _070_ 0.089475f
C4754 FILLER_0_19_195/a_36_472# vss 0.005146f
C4755 FILLER_0_13_80/a_124_375# vss 0.042254f
C4756 FILLER_0_13_80/a_36_472# vdd 0.087291f
C4757 FILLER_0_5_54/a_1380_472# net47 0.003924f
C4758 _095_ _406_/a_36_159# 0.131137f
C4759 net16 _166_ 0.146913f
C4760 _077_ _061_ 0.031458f
C4761 _016_ _428_/a_36_151# 0.001824f
C4762 net81 FILLER_0_15_235/a_124_375# 0.008139f
C4763 net82 FILLER_0_3_172/a_1380_472# 0.007879f
C4764 _449_/a_36_151# _043_ 0.001572f
C4765 FILLER_0_15_116/a_572_375# _136_ 0.001706f
C4766 output40/a_224_472# output41/a_224_472# 0.292611f
C4767 net4 FILLER_0_12_236/a_484_472# 0.014212f
C4768 _122_ _066_ 0.001217f
C4769 net20 _094_ 0.677838f
C4770 FILLER_0_10_256/a_124_375# FILLER_0_10_247/a_124_375# 0.002036f
C4771 net18 _418_/a_1308_423# 0.015651f
C4772 result[1] vss 0.311464f
C4773 FILLER_0_17_142/a_484_472# vdd 0.004902f
C4774 FILLER_0_17_142/a_36_472# vss 0.008239f
C4775 net17 _041_ 0.002779f
C4776 net62 net28 0.05491f
C4777 state\[1\] _121_ 0.006184f
C4778 _394_/a_2215_68# _095_ 0.001134f
C4779 net18 _419_/a_2665_112# 0.0371f
C4780 FILLER_0_18_2/a_484_472# vss 0.001228f
C4781 _016_ _114_ 0.041462f
C4782 _346_/a_49_472# vss 0.0031f
C4783 FILLER_0_9_28/a_484_472# net16 0.021584f
C4784 _086_ FILLER_0_10_107/a_572_375# 0.001179f
C4785 _004_ net19 0.112289f
C4786 _073_ vdd 0.258125f
C4787 _127_ _135_ 0.00622f
C4788 net55 FILLER_0_21_60/a_572_375# 0.041903f
C4789 FILLER_0_18_76/a_572_375# vss 0.007413f
C4790 FILLER_0_18_76/a_36_472# vdd 0.014249f
C4791 net52 _440_/a_448_472# 0.067294f
C4792 net81 _425_/a_2665_112# 0.010188f
C4793 _432_/a_448_472# _139_ 0.001772f
C4794 FILLER_0_13_100/a_36_472# _043_ 0.012726f
C4795 FILLER_0_18_107/a_484_472# FILLER_0_17_104/a_932_472# 0.026657f
C4796 _429_/a_2665_112# vss 0.012165f
C4797 net15 _012_ 0.043755f
C4798 _176_ _124_ 0.036117f
C4799 _423_/a_2248_156# vdd 0.013707f
C4800 _147_ net23 0.011375f
C4801 mask\[4\] FILLER_0_19_171/a_1020_375# 0.006236f
C4802 net57 net53 0.053565f
C4803 _129_ FILLER_0_11_135/a_36_472# 0.078373f
C4804 net69 _152_ 0.002532f
C4805 _443_/a_2248_156# trim_mask\[4\] 0.002315f
C4806 net82 _084_ 0.020793f
C4807 _122_ net37 3.870625f
C4808 net76 _078_ 0.029213f
C4809 FILLER_0_17_72/a_1020_375# _175_ 0.028592f
C4810 fanout69/a_36_113# _160_ 0.005933f
C4811 _321_/a_170_472# net23 0.025371f
C4812 net41 FILLER_0_21_28/a_124_375# 0.003254f
C4813 _074_ _082_ 0.069835f
C4814 FILLER_0_7_72/a_1468_375# net50 0.020186f
C4815 FILLER_0_12_20/a_484_472# FILLER_0_12_28/a_36_472# 0.013277f
C4816 FILLER_0_19_125/a_36_472# vss 0.001056f
C4817 net65 net4 0.614946f
C4818 mask\[8\] _214_/a_36_160# 0.001264f
C4819 net47 _450_/a_448_472# 0.012172f
C4820 _441_/a_2665_112# FILLER_0_3_78/a_572_375# 0.010688f
C4821 trim_mask\[2\] FILLER_0_3_78/a_484_472# 0.008122f
C4822 _013_ FILLER_0_17_56/a_572_375# 0.001047f
C4823 result[0] fanout65/a_36_113# 0.001816f
C4824 FILLER_0_22_128/a_1380_472# vdd 0.005746f
C4825 FILLER_0_22_128/a_932_472# vss 0.003452f
C4826 _128_ _125_ 0.017316f
C4827 _422_/a_796_472# _109_ 0.002086f
C4828 net38 FILLER_0_20_15/a_124_375# 0.012947f
C4829 net50 net16 0.015448f
C4830 _070_ FILLER_0_10_107/a_124_375# 0.009848f
C4831 _024_ _435_/a_1000_472# 0.002902f
C4832 trim_val\[0\] _453_/a_36_151# 0.001629f
C4833 result[6] _420_/a_1204_472# 0.002681f
C4834 _449_/a_2665_112# _172_ 0.003296f
C4835 net66 vdd 0.646189f
C4836 _128_ _315_/a_1657_68# 0.0013f
C4837 result[9] net61 0.014374f
C4838 _086_ _267_/a_672_472# 0.004515f
C4839 _452_/a_36_151# _041_ 0.013289f
C4840 ctln[8] trim_val\[3\] 0.007f
C4841 _053_ FILLER_0_6_47/a_484_472# 0.006301f
C4842 net49 net17 0.029142f
C4843 _415_/a_2560_156# vss 0.001286f
C4844 output20/a_224_472# vdd 0.09529f
C4845 FILLER_0_9_28/a_36_472# vss -0.001119f
C4846 _445_/a_1308_423# vdd 0.001478f
C4847 vss trim[3] 0.235724f
C4848 net68 net17 0.601273f
C4849 trim_val\[1\] _164_ 0.100504f
C4850 net68 _377_/a_36_472# 0.001305f
C4851 net75 _073_ 0.34505f
C4852 _029_ _365_/a_36_68# 0.013994f
C4853 _136_ _137_ 0.417639f
C4854 output35/a_224_472# mask\[7\] 0.004608f
C4855 FILLER_0_15_116/a_36_472# net53 0.005099f
C4856 net4 net59 0.102012f
C4857 mask\[5\] FILLER_0_18_177/a_1916_375# 0.002014f
C4858 _411_/a_2665_112# net8 0.036782f
C4859 FILLER_0_15_282/a_484_472# _417_/a_36_151# 0.059367f
C4860 FILLER_0_15_282/a_36_472# _417_/a_448_472# 0.011962f
C4861 FILLER_0_10_78/a_484_472# vss 0.005854f
C4862 trim_mask\[4\] _170_ 0.09738f
C4863 FILLER_0_10_78/a_1020_375# _389_/a_36_148# 0.001335f
C4864 net58 FILLER_0_9_270/a_572_375# 0.006256f
C4865 _425_/a_36_151# vdd 0.078723f
C4866 _072_ _375_/a_1388_497# 0.001138f
C4867 FILLER_0_10_78/a_1468_375# _308_/a_124_24# 0.001565f
C4868 FILLER_0_9_282/a_124_375# vdd 0.01273f
C4869 _104_ result[6] 0.096535f
C4870 _091_ FILLER_0_18_177/a_484_472# 0.004272f
C4871 vdd _167_ 0.012869f
C4872 mask\[7\] _435_/a_796_472# 0.009587f
C4873 net36 FILLER_0_15_228/a_36_472# 0.008225f
C4874 result[6] _421_/a_2665_112# 0.034452f
C4875 net60 net62 0.002144f
C4876 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_36_472# 0.086904f
C4877 vss FILLER_0_22_107/a_124_375# 0.002881f
C4878 vdd FILLER_0_22_107/a_572_375# 0.005745f
C4879 _092_ FILLER_0_18_209/a_572_375# 0.00609f
C4880 FILLER_0_15_212/a_1020_375# mask\[1\] 0.017527f
C4881 _444_/a_36_151# net42 0.006866f
C4882 _350_/a_49_472# _208_/a_36_160# 0.078981f
C4883 _147_ net33 0.001686f
C4884 output9/a_224_472# vss 0.007544f
C4885 _050_ _436_/a_36_151# 0.037103f
C4886 output37/a_224_472# fanout65/a_36_113# 0.013171f
C4887 _067_ vdd 0.853589f
C4888 _289_/a_36_472# _094_ 0.00922f
C4889 FILLER_0_16_57/a_124_375# _131_ 0.012982f
C4890 FILLER_0_18_107/a_3172_472# FILLER_0_17_133/a_124_375# 0.001543f
C4891 cal_itt\[2\] vdd 0.267121f
C4892 FILLER_0_17_282/a_124_375# net30 0.001288f
C4893 FILLER_0_7_59/a_36_472# fanout67/a_36_160# 0.013068f
C4894 FILLER_0_4_177/a_572_375# net22 0.006125f
C4895 net19 FILLER_0_23_274/a_124_375# 0.01233f
C4896 net55 _424_/a_2665_112# 0.056555f
C4897 net77 _007_ 0.002591f
C4898 FILLER_0_15_72/a_572_375# cal_count\[1\] 0.135344f
C4899 net1 vdd 0.63891f
C4900 _448_/a_2248_156# _443_/a_2248_156# 0.006556f
C4901 FILLER_0_14_99/a_124_375# vdd 0.040312f
C4902 _120_ vss 0.42505f
C4903 net54 vdd 0.877573f
C4904 _104_ mask\[4\] 0.001621f
C4905 _119_ _322_/a_124_24# 0.020461f
C4906 result[6] fanout61/a_36_113# 0.003917f
C4907 _189_/a_67_603# net62 0.001695f
C4908 net31 net33 0.002465f
C4909 FILLER_0_20_15/a_1468_375# vdd 0.009742f
C4910 FILLER_0_16_107/a_484_472# vss 0.004223f
C4911 ctln[6] _442_/a_448_472# 0.003039f
C4912 _232_/a_67_603# net47 0.014888f
C4913 _412_/a_36_151# vdd 0.080326f
C4914 FILLER_0_21_142/a_572_375# FILLER_0_22_128/a_2276_472# 0.001543f
C4915 net17 FILLER_0_20_15/a_932_472# 0.047256f
C4916 _115_ _315_/a_244_497# 0.00153f
C4917 _168_ _164_ 0.092012f
C4918 net79 FILLER_0_12_236/a_484_472# 0.009305f
C4919 _290_/a_224_472# _094_ 0.003006f
C4920 net75 _425_/a_36_151# 0.02868f
C4921 FILLER_0_8_127/a_124_375# _129_ 0.056784f
C4922 FILLER_0_4_177/a_124_375# _087_ 0.002288f
C4923 net79 _416_/a_36_151# 0.062626f
C4924 _090_ net22 0.032492f
C4925 _127_ _129_ 0.716384f
C4926 _273_/a_36_68# FILLER_0_10_214/a_36_472# 0.003036f
C4927 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1468_375# 0.086742f
C4928 FILLER_0_16_107/a_36_472# _451_/a_36_151# 0.059367f
C4929 _009_ _107_ 0.027726f
C4930 _432_/a_36_151# _097_ 0.003144f
C4931 net38 _444_/a_1288_156# 0.001147f
C4932 cal_count\[2\] _402_/a_244_567# 0.004411f
C4933 fanout80/a_36_113# vdd 0.033884f
C4934 net75 cal_itt\[2\] 0.143064f
C4935 _134_ FILLER_0_9_105/a_484_472# 0.011499f
C4936 _448_/a_2248_156# _170_ 0.00254f
C4937 _448_/a_1000_472# _037_ 0.03564f
C4938 _444_/a_796_472# net40 0.005776f
C4939 _062_ _310_/a_49_472# 0.020509f
C4940 _265_/a_916_472# _001_ 0.001719f
C4941 net72 _067_ 0.055817f
C4942 net63 _435_/a_1308_423# 0.003621f
C4943 FILLER_0_20_193/a_572_375# vdd 0.029393f
C4944 net34 _422_/a_2665_112# 0.006103f
C4945 output31/a_224_472# result[9] 0.082001f
C4946 net56 _136_ 0.462275f
C4947 _442_/a_36_151# net23 0.00157f
C4948 _078_ _083_ 0.01015f
C4949 fanout54/a_36_160# FILLER_0_19_155/a_36_472# 0.193804f
C4950 net21 _434_/a_2248_156# 0.001467f
C4951 net75 net1 0.098901f
C4952 _439_/a_2665_112# net14 0.004943f
C4953 _165_ trim_val\[0\] 0.164683f
C4954 FILLER_0_9_28/a_124_375# output42/a_224_472# 0.003337f
C4955 _093_ FILLER_0_19_134/a_36_472# 0.002415f
C4956 _441_/a_448_472# net49 0.001245f
C4957 FILLER_0_9_105/a_36_472# vdd 0.009746f
C4958 FILLER_0_9_105/a_572_375# vss 0.020145f
C4959 mask\[4\] net22 0.075713f
C4960 FILLER_0_5_198/a_124_375# net59 0.00174f
C4961 _308_/a_848_380# _114_ 0.005266f
C4962 FILLER_0_12_2/a_36_472# net67 0.013281f
C4963 _235_/a_67_603# net68 0.027525f
C4964 _181_ _179_ 0.011848f
C4965 FILLER_0_18_139/a_36_472# vss 0.007877f
C4966 FILLER_0_18_139/a_484_472# vdd 0.003106f
C4967 net75 _412_/a_36_151# 0.060039f
C4968 _009_ FILLER_0_23_274/a_124_375# 0.010723f
C4969 net49 _440_/a_1204_472# 0.006692f
C4970 _414_/a_2665_112# _074_ 0.004912f
C4971 output34/a_224_472# _103_ 0.027876f
C4972 FILLER_0_15_116/a_484_472# FILLER_0_14_107/a_1468_375# 0.001723f
C4973 _053_ _042_ 0.00242f
C4974 net64 FILLER_0_15_235/a_124_375# 0.025203f
C4975 _121_ vdd 0.106437f
C4976 net81 _136_ 0.021146f
C4977 net63 _019_ 0.004471f
C4978 FILLER_0_16_154/a_124_375# vss 0.004317f
C4979 FILLER_0_16_154/a_572_375# vdd 0.004706f
C4980 net81 net21 0.185411f
C4981 _032_ _031_ 0.013851f
C4982 _094_ vss 0.24519f
C4983 FILLER_0_15_235/a_124_375# mask\[1\] 0.013103f
C4984 net74 _172_ 0.006643f
C4985 _440_/a_2665_112# trim_mask\[1\] 0.007959f
C4986 _370_/a_848_380# vss 0.051599f
C4987 mask\[7\] FILLER_0_22_128/a_932_472# 0.017448f
C4988 trim[4] net47 0.009333f
C4989 _141_ _093_ 0.396041f
C4990 _432_/a_448_472# _098_ 0.032293f
C4991 net20 _043_ 0.094689f
C4992 FILLER_0_12_50/a_36_472# _453_/a_36_151# 0.001748f
C4993 FILLER_0_15_116/a_36_472# _451_/a_36_151# 0.096503f
C4994 _060_ net21 0.074356f
C4995 FILLER_0_16_73/a_484_472# _131_ 0.007761f
C4996 FILLER_0_7_104/a_124_375# vdd 0.031505f
C4997 _070_ _248_/a_36_68# 0.007095f
C4998 net63 FILLER_0_19_195/a_124_375# 0.017284f
C4999 net39 net49 0.158007f
C5000 net32 _419_/a_1308_423# 0.00191f
C5001 net2 net18 0.030437f
C5002 net55 FILLER_0_17_56/a_484_472# 0.023554f
C5003 _021_ _137_ 0.002807f
C5004 _021_ FILLER_0_18_171/a_124_375# 0.004621f
C5005 net73 FILLER_0_18_107/a_2364_375# 0.015484f
C5006 ctln[4] _411_/a_36_151# 0.0022f
C5007 _115_ FILLER_0_9_72/a_1380_472# 0.007262f
C5008 _153_ net14 0.260217f
C5009 _227_/a_36_160# vss 0.010455f
C5010 net68 FILLER_0_6_47/a_1828_472# 0.009096f
C5011 net38 _034_ 0.025823f
C5012 FILLER_0_4_185/a_36_472# net76 0.023698f
C5013 net82 calibrate 0.002345f
C5014 net15 ctln[8] 0.205163f
C5015 _239_/a_36_160# _065_ 0.032139f
C5016 _418_/a_1308_423# _417_/a_36_151# 0.001518f
C5017 FILLER_0_18_107/a_1020_375# vdd -0.008765f
C5018 _273_/a_36_68# _246_/a_36_68# 0.001168f
C5019 trim_mask\[1\] FILLER_0_6_47/a_2724_472# 0.003645f
C5020 net39 _445_/a_1204_472# 0.002681f
C5021 net52 FILLER_0_9_72/a_124_375# 0.029702f
C5022 _049_ FILLER_0_22_128/a_2812_375# 0.001905f
C5023 FILLER_0_12_124/a_36_472# net74 0.021369f
C5024 net54 FILLER_0_22_128/a_572_375# 0.048634f
C5025 _433_/a_1308_423# _145_ 0.026613f
C5026 FILLER_0_18_37/a_572_375# vdd 0.02259f
C5027 FILLER_0_18_37/a_124_375# vss 0.002958f
C5028 _412_/a_448_472# net18 0.049704f
C5029 _070_ _060_ 0.822179f
C5030 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_572_375# 0.086635f
C5031 FILLER_0_7_72/a_1380_472# _053_ 0.01339f
C5032 output42/a_224_472# net44 0.079084f
C5033 FILLER_0_12_220/a_1380_472# _060_ 0.01563f
C5034 _030_ _367_/a_36_68# 0.015584f
C5035 net37 _160_ 0.003563f
C5036 FILLER_0_11_64/a_124_375# _120_ 0.004514f
C5037 _446_/a_2665_112# vdd 0.044081f
C5038 _415_/a_1308_423# result[1] 0.00761f
C5039 ctln[4] _413_/a_448_472# 0.001072f
C5040 _421_/a_2665_112# _419_/a_2248_156# 0.001545f
C5041 state\[2\] FILLER_0_13_142/a_484_472# 0.004186f
C5042 net53 FILLER_0_13_142/a_1380_472# 0.041222f
C5043 cal net18 0.123815f
C5044 _415_/a_796_472# net27 0.004502f
C5045 FILLER_0_5_72/a_932_472# vdd 0.002735f
C5046 FILLER_0_5_72/a_484_472# vss 0.003738f
C5047 output14/a_224_472# _442_/a_2248_156# 0.001723f
C5048 net75 _411_/a_796_472# 0.006358f
C5049 net16 _054_ 0.044357f
C5050 _157_ _160_ 0.010231f
C5051 FILLER_0_4_144/a_572_375# _081_ 0.002236f
C5052 FILLER_0_4_144/a_124_375# _152_ 0.007333f
C5053 _065_ _036_ 0.031728f
C5054 _272_/a_36_472# vdd 0.058326f
C5055 _029_ _154_ 0.116532f
C5056 _128_ _069_ 0.018491f
C5057 _176_ _180_ 0.030701f
C5058 _076_ net22 0.03249f
C5059 result[6] _419_/a_2248_156# 0.002634f
C5060 FILLER_0_20_107/a_124_375# _098_ 0.01186f
C5061 FILLER_0_5_109/a_572_375# _163_ 0.003096f
C5062 output32/a_224_472# net30 0.001139f
C5063 _003_ _079_ 0.035497f
C5064 _089_ _088_ 0.009863f
C5065 result[8] _422_/a_36_151# 0.001488f
C5066 _032_ _371_/a_36_113# 0.030245f
C5067 FILLER_0_6_90/a_484_472# _163_ 0.011711f
C5068 _413_/a_36_151# FILLER_0_3_172/a_1468_375# 0.001252f
C5069 _067_ cal_count\[0\] 0.201595f
C5070 FILLER_0_2_93/a_36_472# net69 0.010977f
C5071 output9/a_224_472# net4 0.042449f
C5072 _324_/a_224_472# _129_ 0.009728f
C5073 FILLER_0_4_197/a_484_472# _088_ 0.014756f
C5074 FILLER_0_8_107/a_124_375# _219_/a_36_160# 0.002515f
C5075 _070_ _330_/a_224_472# 0.001096f
C5076 FILLER_0_18_177/a_1468_375# FILLER_0_20_177/a_1380_472# 0.0027f
C5077 _079_ net21 0.065561f
C5078 mask\[5\] vdd 0.79138f
C5079 _176_ _451_/a_2225_156# 0.030788f
C5080 net60 net33 0.008865f
C5081 _069_ FILLER_0_11_142/a_572_375# 0.020472f
C5082 FILLER_0_18_209/a_124_375# vss 0.004598f
C5083 FILLER_0_18_209/a_572_375# vdd 0.021356f
C5084 _040_ net14 0.069672f
C5085 _286_/a_224_472# vdd 0.00154f
C5086 FILLER_0_8_24/a_572_375# vdd 0.011353f
C5087 FILLER_0_7_72/a_572_375# vss 0.006884f
C5088 _256_/a_2124_68# _070_ 0.002444f
C5089 _184_ net17 0.007958f
C5090 net15 _449_/a_2248_156# 0.001705f
C5091 FILLER_0_18_107/a_36_472# mask\[9\] 0.005458f
C5092 _345_/a_36_160# _098_ 0.002041f
C5093 FILLER_0_12_220/a_124_375# vdd -0.008946f
C5094 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_36_472# 0.086905f
C5095 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2812_375# 0.001597f
C5096 net57 _071_ 0.12089f
C5097 FILLER_0_22_128/a_1380_472# _433_/a_36_151# 0.001973f
C5098 net23 _433_/a_2665_112# 0.015555f
C5099 mask\[3\] net36 0.002974f
C5100 net26 vdd 0.487733f
C5101 net78 net18 1.351707f
C5102 net31 _046_ 0.008368f
C5103 FILLER_0_4_107/a_572_375# _160_ 0.008945f
C5104 _426_/a_796_472# net64 0.006933f
C5105 net15 FILLER_0_17_72/a_36_472# 0.006905f
C5106 FILLER_0_11_124/a_124_375# vdd 0.016626f
C5107 _136_ _095_ 0.043768f
C5108 FILLER_0_23_274/a_36_472# vss 0.002346f
C5109 _053_ _169_ 0.014161f
C5110 output29/a_224_472# _416_/a_36_151# 0.07368f
C5111 output23/a_224_472# net23 0.122379f
C5112 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_36_472# 0.016748f
C5113 result[1] net79 0.25261f
C5114 net29 _006_ 0.135646f
C5115 net57 _386_/a_692_472# 0.00409f
C5116 _170_ _066_ 0.189122f
C5117 _063_ _166_ 0.025402f
C5118 output36/a_224_472# net30 0.083671f
C5119 _449_/a_1204_472# _038_ 0.005899f
C5120 FILLER_0_16_57/a_932_472# _176_ 0.010635f
C5121 FILLER_0_5_117/a_36_472# vss 0.001215f
C5122 result[5] net18 0.173673f
C5123 net65 FILLER_0_1_212/a_124_375# 0.005253f
C5124 FILLER_0_5_109/a_572_375# FILLER_0_4_107/a_932_472# 0.001684f
C5125 fanout70/a_36_113# net53 0.031633f
C5126 net73 net70 0.040702f
C5127 FILLER_0_7_59/a_124_375# net68 0.019553f
C5128 _104_ result[7] 0.475003f
C5129 _346_/a_49_472# _141_ 0.104653f
C5130 _012_ net71 0.004946f
C5131 net65 FILLER_0_2_177/a_36_472# 0.016652f
C5132 net27 vss 0.534444f
C5133 _093_ _397_/a_36_472# 0.001509f
C5134 FILLER_0_5_54/a_932_472# vss 0.003426f
C5135 FILLER_0_5_54/a_1380_472# vdd 0.008983f
C5136 cal_count\[2\] _452_/a_1353_112# 0.002558f
C5137 _133_ _068_ 0.002552f
C5138 _195_/a_67_603# vdd 0.022493f
C5139 net52 FILLER_0_3_78/a_36_472# 0.034084f
C5140 _053_ net59 0.145863f
C5141 _093_ FILLER_0_17_218/a_484_472# 0.004665f
C5142 net48 _074_ 1.192591f
C5143 _424_/a_36_151# FILLER_0_18_37/a_572_375# 0.002807f
C5144 output8/a_224_472# _080_ 0.001971f
C5145 net17 net47 2.009509f
C5146 FILLER_0_7_72/a_1380_472# _028_ 0.001777f
C5147 result[7] result[6] 0.119475f
C5148 net26 net72 0.868238f
C5149 FILLER_0_16_37/a_36_472# _184_ 0.001522f
C5150 net15 _440_/a_36_151# 0.016061f
C5151 _074_ _162_ 0.112872f
C5152 net54 _436_/a_448_472# 0.006129f
C5153 _414_/a_1288_156# cal_itt\[3\] 0.001354f
C5154 vdd net30 0.636147f
C5155 net62 output30/a_224_472# 0.074425f
C5156 net44 net6 0.005889f
C5157 _440_/a_2665_112# _164_ 0.067034f
C5158 FILLER_0_24_63/a_36_472# output26/a_224_472# 0.023414f
C5159 _431_/a_2248_156# vss 0.041929f
C5160 _151_ vss 0.050544f
C5161 net76 _263_/a_224_472# 0.00132f
C5162 _088_ FILLER_0_4_213/a_36_472# 0.01735f
C5163 _183_ _180_ 0.002621f
C5164 _285_/a_36_472# _196_/a_36_160# 0.004619f
C5165 net8 FILLER_0_0_266/a_124_375# 0.001181f
C5166 net54 _433_/a_36_151# 0.00661f
C5167 result[8] net21 0.166555f
C5168 FILLER_0_7_162/a_36_472# net57 0.015199f
C5169 _438_/a_448_472# net71 0.044454f
C5170 FILLER_0_2_177/a_36_472# net59 0.007582f
C5171 FILLER_0_10_28/a_124_375# net40 0.047331f
C5172 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_36_472# 0.012267f
C5173 FILLER_0_21_142/a_484_472# vss 0.034607f
C5174 mask\[3\] _432_/a_2248_156# 0.002775f
C5175 _315_/a_716_497# _120_ 0.001321f
C5176 _187_ _188_ 0.001453f
C5177 _413_/a_448_472# net21 0.052657f
C5178 FILLER_0_19_47/a_484_472# FILLER_0_18_37/a_1468_375# 0.001684f
C5179 _394_/a_1336_472# FILLER_0_15_72/a_124_375# 0.016876f
C5180 net58 output27/a_224_472# 0.121438f
C5181 _013_ _012_ 0.003113f
C5182 FILLER_0_9_223/a_484_472# _223_/a_36_160# 0.004695f
C5183 net81 valid 0.11798f
C5184 net73 _132_ 0.460325f
C5185 _292_/a_36_160# vss 0.009517f
C5186 net16 _217_/a_36_160# 0.00629f
C5187 net31 net18 0.114197f
C5188 _104_ _008_ 0.135471f
C5189 FILLER_0_9_28/a_3260_375# net68 0.009969f
C5190 FILLER_0_17_38/a_572_375# vss 0.007503f
C5191 FILLER_0_17_38/a_36_472# vdd 0.01637f
C5192 vss _450_/a_36_151# 0.02803f
C5193 vdd _450_/a_448_472# 0.011591f
C5194 _074_ net19 0.035973f
C5195 _098_ _433_/a_1000_472# 0.0184f
C5196 _136_ mask\[1\] 0.407932f
C5197 _255_/a_224_552# _090_ 0.001598f
C5198 net32 net19 0.65591f
C5199 net63 _202_/a_36_160# 0.004414f
C5200 mask\[1\] net21 0.023956f
C5201 _043_ vss 1.362912f
C5202 net16 _035_ 0.034977f
C5203 _115_ _171_ 0.033359f
C5204 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_484_472# 0.013277f
C5205 net47 _452_/a_36_151# 0.021978f
C5206 net41 _444_/a_448_472# 0.031876f
C5207 FILLER_0_17_200/a_572_375# FILLER_0_18_177/a_3172_472# 0.001597f
C5208 net74 _152_ 1.007413f
C5209 net26 _424_/a_36_151# 0.062638f
C5210 _038_ FILLER_0_11_78/a_484_472# 0.001782f
C5211 net32 mask\[6\] 0.003248f
C5212 _057_ cal_itt\[3\] 0.014849f
C5213 _065_ output15/a_224_472# 0.037721f
C5214 _267_/a_672_472# _071_ 0.00255f
C5215 _106_ output18/a_224_472# 0.005393f
C5216 net54 FILLER_0_19_134/a_124_375# 0.002681f
C5217 FILLER_0_13_65/a_36_472# vdd 0.005885f
C5218 _185_ vss 0.021437f
C5219 _448_/a_2665_112# net22 0.010428f
C5220 net64 FILLER_0_12_220/a_1380_472# 0.011079f
C5221 _434_/a_2560_156# mask\[6\] 0.010913f
C5222 FILLER_0_19_125/a_124_375# _022_ 0.055527f
C5223 FILLER_0_16_37/a_36_472# net47 0.008304f
C5224 output15/a_224_472# FILLER_0_0_96/a_36_472# 0.023414f
C5225 _058_ FILLER_0_9_105/a_124_375# 0.014234f
C5226 FILLER_0_21_28/a_2812_375# _012_ 0.016736f
C5227 net74 _318_/a_224_472# 0.001513f
C5228 ctlp[4] vdd 0.278868f
C5229 FILLER_0_5_164/a_36_472# _169_ 0.00284f
C5230 FILLER_0_5_164/a_572_375# _163_ 0.046852f
C5231 _422_/a_2248_156# net19 0.003451f
C5232 _175_ vss 0.162988f
C5233 net80 _340_/a_36_160# 0.004225f
C5234 _256_/a_1612_497# _068_ 0.002759f
C5235 _093_ FILLER_0_17_104/a_572_375# 0.01418f
C5236 output36/a_224_472# FILLER_0_14_263/a_36_472# 0.001711f
C5237 _115_ _176_ 1.300336f
C5238 net57 net55 0.001926f
C5239 _430_/a_1204_472# _069_ 0.001629f
C5240 net72 FILLER_0_17_38/a_36_472# 0.123542f
C5241 FILLER_0_5_117/a_124_375# _154_ 0.005866f
C5242 _261_/a_36_160# vss 0.05095f
C5243 _233_/a_36_160# FILLER_0_6_37/a_124_375# 0.001713f
C5244 _157_ _156_ 0.005264f
C5245 net50 net14 0.192231f
C5246 net36 FILLER_0_20_87/a_36_472# 0.074773f
C5247 _122_ _160_ 0.004488f
C5248 FILLER_0_10_107/a_484_472# vss 0.00298f
C5249 output35/a_224_472# ctlp[2] 0.001465f
C5250 net55 _027_ 0.002104f
C5251 _328_/a_36_113# _070_ 0.016264f
C5252 net74 _136_ 0.042043f
C5253 _086_ _057_ 0.82902f
C5254 trim_mask\[1\] FILLER_0_6_90/a_36_472# 0.001162f
C5255 _414_/a_448_472# vdd 0.013377f
C5256 mask\[4\] FILLER_0_18_177/a_932_472# 0.016924f
C5257 FILLER_0_17_200/a_484_472# _069_ 0.001396f
C5258 mask\[4\] _140_ 0.001697f
C5259 _075_ FILLER_0_5_206/a_36_472# 0.001503f
C5260 FILLER_0_20_177/a_484_472# vss 0.001256f
C5261 FILLER_0_20_177/a_932_472# vdd 0.035019f
C5262 _088_ FILLER_0_3_221/a_484_472# 0.002245f
C5263 net32 _009_ 0.003756f
C5264 _440_/a_1204_472# net47 0.006257f
C5265 net35 FILLER_0_22_86/a_572_375# 0.010986f
C5266 mask\[8\] FILLER_0_22_86/a_1020_375# 0.009431f
C5267 net52 _442_/a_448_472# 0.044149f
C5268 _232_/a_67_603# vdd 0.007565f
C5269 FILLER_0_17_200/a_36_472# _093_ 0.005101f
C5270 FILLER_0_13_65/a_36_472# net72 0.00272f
C5271 FILLER_0_14_263/a_124_375# vss 0.007923f
C5272 FILLER_0_14_263/a_36_472# vdd 0.02759f
C5273 FILLER_0_16_89/a_36_472# _451_/a_2225_156# 0.001329f
C5274 _045_ mask\[1\] 0.024178f
C5275 net50 _447_/a_2665_112# 0.015374f
C5276 _221_/a_36_160# net40 0.002952f
C5277 _096_ mask\[0\] 0.052773f
C5278 _069_ _429_/a_1000_472# 0.029501f
C5279 _411_/a_2560_156# ctln[1] 0.001413f
C5280 net52 _029_ 0.03261f
C5281 net74 _070_ 0.394108f
C5282 _321_/a_3126_472# _176_ 0.001932f
C5283 _069_ _395_/a_1492_488# 0.002565f
C5284 _004_ _415_/a_448_472# 0.044374f
C5285 net82 _443_/a_1204_472# 0.004056f
C5286 FILLER_0_3_142/a_36_472# _370_/a_848_380# 0.001207f
C5287 net65 _425_/a_2248_156# 0.003451f
C5288 _323_/a_36_113# _223_/a_36_160# 0.238626f
C5289 _095_ FILLER_0_14_107/a_484_472# 0.014431f
C5290 _083_ _263_/a_224_472# 0.003191f
C5291 net78 _109_ 0.001432f
C5292 FILLER_0_18_177/a_572_375# vdd 0.031241f
C5293 FILLER_0_18_177/a_124_375# vss 0.00364f
C5294 net57 net23 0.324262f
C5295 net44 FILLER_0_15_2/a_572_375# 0.041552f
C5296 ctln[5] _448_/a_796_472# 0.001484f
C5297 _192_/a_67_603# mask\[1\] 0.020097f
C5298 net39 net47 0.13057f
C5299 result[7] _419_/a_2248_156# 0.001916f
C5300 net58 ctln[1] 0.014147f
C5301 _131_ FILLER_0_17_56/a_124_375# 0.001609f
C5302 FILLER_0_2_127/a_36_472# vdd 0.08468f
C5303 FILLER_0_2_127/a_124_375# vss 0.008566f
C5304 _128_ _090_ 0.018296f
C5305 _178_ FILLER_0_14_50/a_36_472# 0.001492f
C5306 FILLER_0_7_59/a_572_375# net67 0.007538f
C5307 _071_ FILLER_0_13_142/a_1380_472# 0.001617f
C5308 FILLER_0_14_91/a_124_375# vdd -0.010114f
C5309 net27 net4 0.025834f
C5310 _255_/a_224_552# _076_ 0.081663f
C5311 net79 _094_ 0.301878f
C5312 _138_ vdd 0.090752f
C5313 net47 _039_ 0.042757f
C5314 vdd FILLER_0_10_94/a_36_472# 0.086035f
C5315 vss FILLER_0_10_94/a_572_375# 0.013232f
C5316 ctlp[5] _147_ 0.001406f
C5317 mask\[8\] _437_/a_2248_156# 0.004415f
C5318 _422_/a_2248_156# _009_ 0.061786f
C5319 FILLER_0_16_57/a_1468_375# net15 0.012909f
C5320 _095_ _451_/a_448_472# 0.002474f
C5321 _348_/a_49_472# vdd 0.038046f
C5322 _417_/a_448_472# _006_ 0.068545f
C5323 _430_/a_448_472# net80 0.00896f
C5324 FILLER_0_10_37/a_124_375# _173_ 0.00262f
C5325 _074_ FILLER_0_3_172/a_484_472# 0.001763f
C5326 FILLER_0_19_55/a_36_472# net36 0.001068f
C5327 _093_ FILLER_0_17_133/a_36_472# 0.010432f
C5328 _389_/a_36_148# _172_ 0.039684f
C5329 net13 _170_ 0.001668f
C5330 FILLER_0_19_171/a_1380_472# vss 0.004488f
C5331 _091_ FILLER_0_13_212/a_932_472# 0.008749f
C5332 FILLER_0_5_172/a_124_375# net22 0.002388f
C5333 comp FILLER_0_15_2/a_36_472# 0.001941f
C5334 _178_ cal_count\[3\] 0.002061f
C5335 FILLER_0_11_101/a_124_375# cal_count\[3\] 0.00419f
C5336 FILLER_0_21_142/a_484_472# mask\[7\] 0.001603f
C5337 FILLER_0_10_78/a_36_472# _453_/a_2665_112# 0.007491f
C5338 _176_ _394_/a_728_93# 0.002001f
C5339 _128_ net22 0.03249f
C5340 FILLER_0_18_177/a_1828_472# net21 0.001887f
C5341 _131_ _040_ 0.211618f
C5342 _438_/a_2248_156# vdd 0.024595f
C5343 output21/a_224_472# _107_ 0.086601f
C5344 _444_/a_36_151# net67 0.055072f
C5345 _373_/a_1254_68# _090_ 0.001326f
C5346 _131_ _125_ 0.013932f
C5347 result[9] _420_/a_2248_156# 0.046636f
C5348 FILLER_0_18_2/a_3260_375# FILLER_0_20_31/a_36_472# 0.001338f
C5349 _430_/a_36_151# FILLER_0_18_177/a_2276_472# 0.001793f
C5350 FILLER_0_4_177/a_36_472# net37 0.004017f
C5351 net60 net18 0.949607f
C5352 FILLER_0_17_72/a_3260_375# _451_/a_1040_527# 0.001117f
C5353 _083_ _265_/a_224_472# 0.003404f
C5354 FILLER_0_15_282/a_36_472# _006_ 0.003055f
C5355 trim[4] vdd 0.198218f
C5356 _413_/a_2665_112# cal_itt\[2\] 0.003007f
C5357 _301_/a_36_472# net35 0.051887f
C5358 _008_ _418_/a_448_472# 0.052899f
C5359 _137_ FILLER_0_19_155/a_572_375# 0.030256f
C5360 _074_ cal_itt\[0\] 0.076802f
C5361 _450_/a_836_156# _039_ 0.019042f
C5362 output36/a_224_472# _417_/a_2665_112# 0.008243f
C5363 _110_ _012_ 0.046196f
C5364 _432_/a_448_472# _137_ 0.008956f
C5365 _178_ net40 0.029542f
C5366 ctlp[3] _109_ 0.001371f
C5367 _449_/a_36_151# FILLER_0_13_72/a_484_472# 0.001723f
C5368 FILLER_0_12_136/a_124_375# vss 0.004063f
C5369 FILLER_0_12_136/a_572_375# vdd 0.016972f
C5370 _413_/a_2248_156# FILLER_0_1_212/a_36_472# 0.035805f
C5371 _402_/a_728_93# vdd 0.050988f
C5372 net62 _196_/a_36_160# 0.029171f
C5373 net27 _415_/a_1308_423# 0.02437f
C5374 _174_ _131_ 0.002314f
C5375 _410_/a_36_68# _187_ 0.038745f
C5376 trim_val\[4\] _443_/a_2560_156# 0.049334f
C5377 _448_/a_2560_156# trim_mask\[4\] 0.001306f
C5378 net53 _451_/a_3129_107# 0.002806f
C5379 net20 _418_/a_2248_156# 0.003507f
C5380 valid net64 0.022969f
C5381 _423_/a_448_472# _012_ 0.038928f
C5382 net41 FILLER_0_20_31/a_36_472# 0.030033f
C5383 _016_ fanout73/a_36_113# 0.001731f
C5384 net73 FILLER_0_19_111/a_124_375# 0.005778f
C5385 FILLER_0_17_104/a_36_472# net14 0.012286f
C5386 _031_ _369_/a_692_472# 0.00359f
C5387 ctln[6] _031_ 0.004486f
C5388 _086_ cal_count\[3\] 0.259095f
C5389 _069_ FILLER_0_15_205/a_124_375# 0.002728f
C5390 FILLER_0_3_172/a_2276_472# net22 0.012151f
C5391 net81 FILLER_0_10_256/a_36_472# 0.089055f
C5392 _427_/a_2248_156# _043_ 0.001148f
C5393 _384_/a_224_472# vss 0.004801f
C5394 _081_ _169_ 0.260462f
C5395 _417_/a_2665_112# vdd 0.03015f
C5396 net62 _417_/a_1000_472# 0.005762f
C5397 fanout57/a_36_113# net22 0.024465f
C5398 net57 trim_val\[4\] 0.295336f
C5399 result[7] FILLER_0_23_282/a_484_472# 0.013947f
C5400 FILLER_0_14_107/a_1020_375# FILLER_0_16_115/a_36_472# 0.001512f
C5401 _074_ FILLER_0_6_177/a_484_472# 0.002068f
C5402 FILLER_0_9_28/a_2276_472# net68 0.023299f
C5403 _069_ _098_ 0.029447f
C5404 _424_/a_1204_472# _012_ 0.003572f
C5405 _295_/a_244_68# _107_ 0.00123f
C5406 FILLER_0_18_2/a_124_375# vdd 0.008721f
C5407 _077_ _068_ 0.601166f
C5408 _130_ _428_/a_2248_156# 0.006602f
C5409 ctlp[3] _422_/a_448_472# 0.001441f
C5410 sample result[0] 0.081581f
C5411 FILLER_0_18_53/a_572_375# vdd 0.018416f
C5412 _128_ _076_ 0.04562f
C5413 net35 FILLER_0_22_177/a_36_472# 0.005721f
C5414 FILLER_0_22_86/a_484_472# net71 0.00583f
C5415 output38/a_224_472# net17 0.04454f
C5416 FILLER_0_3_172/a_1916_375# vdd -0.010166f
C5417 net44 _067_ 0.001203f
C5418 _136_ _097_ 0.002577f
C5419 result[0] vss 0.291352f
C5420 FILLER_0_21_206/a_124_375# net21 0.035287f
C5421 _052_ FILLER_0_21_28/a_1916_375# 0.002388f
C5422 _422_/a_2665_112# vss 0.006352f
C5423 _033_ vss 0.019158f
C5424 _067_ _171_ 0.007069f
C5425 FILLER_0_21_28/a_572_375# net17 0.001455f
C5426 cal_itt\[3\] net59 0.018616f
C5427 _438_/a_36_151# net14 0.008367f
C5428 FILLER_0_16_255/a_36_472# net19 0.001273f
C5429 trim_val\[4\] _037_ 0.258184f
C5430 FILLER_0_2_111/a_124_375# _157_ 0.028285f
C5431 net34 _050_ 0.004662f
C5432 _001_ cal_itt\[1\] 0.057933f
C5433 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_124_375# 0.012267f
C5434 _274_/a_2960_68# _070_ 0.001963f
C5435 FILLER_0_13_212/a_1020_375# _043_ 0.01418f
C5436 _093_ FILLER_0_18_107/a_36_472# 0.008683f
C5437 _087_ FILLER_0_3_172/a_1828_472# 0.027954f
C5438 _414_/a_36_151# _079_ 0.037562f
C5439 FILLER_0_11_142/a_572_375# _076_ 0.031784f
C5440 _102_ mask\[2\] 0.036292f
C5441 FILLER_0_12_2/a_572_375# vdd 0.022401f
C5442 _412_/a_2248_156# vdd 0.005671f
C5443 _030_ net49 0.046089f
C5444 _081_ net59 0.185504f
C5445 _098_ FILLER_0_15_212/a_36_472# 0.011079f
C5446 _126_ _125_ 0.032402f
C5447 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_36_472# 0.001963f
C5448 net69 _441_/a_2560_156# 0.002904f
C5449 FILLER_0_8_138/a_124_375# vdd 0.024547f
C5450 _087_ net37 0.23484f
C5451 _093_ FILLER_0_16_89/a_484_472# 0.001526f
C5452 _439_/a_36_151# _453_/a_2665_112# 0.001738f
C5453 _005_ _416_/a_36_151# 0.018752f
C5454 net15 FILLER_0_17_64/a_36_472# 0.015524f
C5455 fanout50/a_36_160# _164_ 0.08721f
C5456 output13/a_224_472# net23 0.00255f
C5457 _431_/a_448_472# _020_ 0.05255f
C5458 _036_ net66 0.04474f
C5459 net68 _030_ 0.007737f
C5460 FILLER_0_12_220/a_1380_472# FILLER_0_12_236/a_36_472# 0.013277f
C5461 net27 net79 0.059863f
C5462 FILLER_0_5_72/a_124_375# FILLER_0_5_54/a_1468_375# 0.005439f
C5463 FILLER_0_18_2/a_2724_472# net17 0.017841f
C5464 trimb[0] FILLER_0_20_2/a_124_375# 0.006864f
C5465 net50 _444_/a_2560_156# 0.001479f
C5466 _277_/a_36_160# vdd 0.115507f
C5467 FILLER_0_3_172/a_3172_472# net21 0.037958f
C5468 ctlp[8] vss 0.107975f
C5469 mask\[9\] FILLER_0_19_111/a_484_472# 0.041744f
C5470 _001_ vss 0.004381f
C5471 _187_ net41 0.002046f
C5472 _448_/a_36_151# net76 0.03831f
C5473 FILLER_0_22_86/a_1020_375# _026_ 0.001032f
C5474 output29/a_224_472# _094_ 0.006731f
C5475 net52 FILLER_0_5_72/a_36_472# 0.014911f
C5476 _176_ _067_ 0.046599f
C5477 net22 _435_/a_36_151# 0.001559f
C5478 FILLER_0_0_130/a_124_375# _442_/a_36_151# 0.059049f
C5479 output48/a_224_472# net76 0.069862f
C5480 mask\[0\] _429_/a_36_151# 0.026729f
C5481 output37/a_224_472# sample 0.015298f
C5482 _079_ _084_ 0.046584f
C5483 net35 FILLER_0_23_88/a_36_472# 0.00675f
C5484 FILLER_0_4_197/a_124_375# net76 0.00811f
C5485 _350_/a_49_472# vdd 0.026837f
C5486 net42 net47 0.237866f
C5487 net51 _450_/a_3129_107# 0.030082f
C5488 FILLER_0_2_111/a_484_472# vdd 0.005951f
C5489 _105_ _205_/a_36_160# 0.001167f
C5490 _062_ vss 0.58133f
C5491 _430_/a_36_151# _093_ 0.00184f
C5492 output37/a_224_472# vss 0.026983f
C5493 FILLER_0_20_177/a_124_375# _098_ 0.018701f
C5494 output32/a_224_472# _418_/a_2665_112# 0.011048f
C5495 _428_/a_1204_472# _131_ 0.012968f
C5496 net73 vdd 0.44835f
C5497 _036_ _167_ 0.003223f
C5498 _057_ _161_ 1.09228f
C5499 _105_ net19 0.049611f
C5500 FILLER_0_9_60/a_36_472# net51 0.059421f
C5501 net78 _418_/a_36_151# 0.003648f
C5502 _073_ _082_ 0.009987f
C5503 _068_ net37 0.006392f
C5504 _198_/a_67_603# mask\[2\] 0.005143f
C5505 _136_ FILLER_0_15_180/a_124_375# 0.002442f
C5506 net81 output28/a_224_472# 0.01335f
C5507 _016_ FILLER_0_12_136/a_484_472# 0.001516f
C5508 _149_ _437_/a_2560_156# 0.008064f
C5509 output17/a_224_472# net43 0.006661f
C5510 net17 vdd 2.139315f
C5511 _086_ _321_/a_2590_472# 0.001522f
C5512 FILLER_0_3_2/a_124_375# _446_/a_36_151# 0.023595f
C5513 net34 _435_/a_1204_472# 0.004285f
C5514 FILLER_0_17_56/a_484_472# FILLER_0_18_61/a_36_472# 0.026657f
C5515 _105_ mask\[6\] 0.029716f
C5516 net41 _445_/a_2248_156# 0.065247f
C5517 _093_ FILLER_0_17_72/a_1916_375# 0.017467f
C5518 FILLER_0_18_2/a_2724_472# _452_/a_36_151# 0.011733f
C5519 FILLER_0_10_78/a_36_472# vdd 0.001865f
C5520 FILLER_0_13_142/a_1380_472# net23 0.026285f
C5521 _031_ _154_ 0.037238f
C5522 net69 _153_ 0.003678f
C5523 net15 FILLER_0_21_60/a_572_375# 0.03167f
C5524 mask\[4\] FILLER_0_19_155/a_484_472# 0.024522f
C5525 net47 clkc 0.002956f
C5526 net79 _043_ 0.393702f
C5527 FILLER_0_8_107/a_36_472# vdd 0.117254f
C5528 net81 _429_/a_1308_423# 0.008913f
C5529 _441_/a_1308_423# _168_ 0.044302f
C5530 _430_/a_1204_472# net22 0.028536f
C5531 _053_ _372_/a_3126_472# 0.001056f
C5532 FILLER_0_7_72/a_572_375# _053_ 0.014569f
C5533 FILLER_0_13_65/a_124_375# _067_ 0.001283f
C5534 result[5] _418_/a_36_151# 0.009705f
C5535 FILLER_0_9_223/a_572_375# vdd 0.007158f
C5536 FILLER_0_14_50/a_36_472# FILLER_0_12_50/a_124_375# 0.0027f
C5537 ctln[1] FILLER_0_0_266/a_36_472# 0.011046f
C5538 _099_ _195_/a_67_603# 0.065049f
C5539 output24/a_224_472# _050_ 0.061723f
C5540 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_124_375# 0.012222f
C5541 cal_count\[3\] FILLER_0_11_78/a_124_375# 0.019818f
C5542 result[7] FILLER_0_24_290/a_36_472# 0.005185f
C5543 FILLER_0_9_28/a_124_375# FILLER_0_8_24/a_572_375# 0.05841f
C5544 _098_ FILLER_0_15_235/a_36_472# 0.093007f
C5545 FILLER_0_17_200/a_484_472# mask\[4\] 0.001701f
C5546 FILLER_0_4_144/a_484_472# vss 0.033414f
C5547 FILLER_0_17_200/a_484_472# net22 0.020589f
C5548 _099_ net30 0.05959f
C5549 FILLER_0_3_142/a_36_472# _261_/a_36_160# 0.001542f
C5550 net60 _109_ 0.021502f
C5551 _098_ _438_/a_36_151# 0.009083f
C5552 net63 FILLER_0_19_171/a_932_472# 0.00128f
C5553 cal_count\[3\] FILLER_0_12_50/a_124_375# 0.060164f
C5554 ctln[0] output40/a_224_472# 0.017541f
C5555 net76 FILLER_0_5_212/a_36_472# 0.00377f
C5556 _274_/a_3368_68# _069_ 0.001414f
C5557 FILLER_0_19_125/a_36_472# _022_ 0.013011f
C5558 _452_/a_36_151# vdd 0.109842f
C5559 _176_ _121_ 0.035608f
C5560 net55 _052_ 0.095046f
C5561 _136_ _019_ 0.049263f
C5562 _430_/a_2560_156# net36 0.00164f
C5563 _429_/a_1000_472# net22 0.007429f
C5564 output13/a_224_472# trim_val\[4\] 0.001014f
C5565 _053_ _220_/a_255_603# 0.001311f
C5566 _058_ FILLER_0_10_94/a_124_375# 0.001597f
C5567 FILLER_0_8_138/a_36_472# _059_ 0.02252f
C5568 _019_ net21 0.065941f
C5569 net72 net17 0.004503f
C5570 _041_ FILLER_0_18_37/a_1468_375# 0.001032f
C5571 net17 _452_/a_1040_527# 0.034254f
C5572 _143_ vdd 0.074199f
C5573 net35 _023_ 0.008361f
C5574 net60 _417_/a_36_151# 0.007446f
C5575 FILLER_0_17_72/a_1828_472# vss 0.001443f
C5576 FILLER_0_17_72/a_2276_472# vdd 0.001409f
C5577 _021_ _097_ 0.002219f
C5578 _228_/a_36_68# _060_ 0.016962f
C5579 _105_ _009_ 0.01731f
C5580 _425_/a_36_151# FILLER_0_8_247/a_36_472# 0.02628f
C5581 _425_/a_1308_423# FILLER_0_8_247/a_1020_375# 0.001064f
C5582 FILLER_0_21_206/a_36_472# _204_/a_67_603# 0.003123f
C5583 FILLER_0_7_72/a_3260_375# vss 0.053035f
C5584 _068_ FILLER_0_5_148/a_484_472# 0.016952f
C5585 FILLER_0_16_37/a_124_375# vss 0.021237f
C5586 FILLER_0_16_37/a_36_472# vdd 0.142203f
C5587 net38 output39/a_224_472# 0.036027f
C5588 net34 output19/a_224_472# 0.122464f
C5589 _053_ FILLER_0_5_54/a_932_472# 0.001578f
C5590 FILLER_0_9_223/a_484_472# state\[0\] 0.007034f
C5591 ctln[4] _413_/a_2248_156# 0.001253f
C5592 net60 _421_/a_2248_156# 0.036944f
C5593 FILLER_0_19_195/a_124_375# net21 0.039225f
C5594 _418_/a_2665_112# vdd 0.028061f
C5595 mask\[2\] FILLER_0_15_180/a_484_472# 0.00848f
C5596 net33 _434_/a_2665_112# 0.001043f
C5597 _422_/a_2665_112# mask\[7\] 0.028271f
C5598 _440_/a_2665_112# FILLER_0_4_91/a_124_375# 0.006271f
C5599 cal_itt\[2\] _082_ 0.032565f
C5600 net81 calibrate 0.047274f
C5601 net57 _428_/a_1000_472# 0.024803f
C5602 _091_ FILLER_0_15_212/a_484_472# 0.049391f
C5603 _450_/a_2225_156# net40 0.04513f
C5604 net20 _102_ 0.081029f
C5605 output7/a_224_472# trim[2] 0.008581f
C5606 output23/a_224_472# ctlp[5] 0.005152f
C5607 _426_/a_2665_112# calibrate 0.004837f
C5608 cal_count\[3\] FILLER_0_11_109/a_36_472# 0.00702f
C5609 _413_/a_1204_472# net82 0.00291f
C5610 net1 _082_ 0.033169f
C5611 _011_ vss 0.003987f
C5612 output9/a_224_472# fanout81/a_36_160# 0.012218f
C5613 FILLER_0_4_213/a_36_472# net59 0.044235f
C5614 _140_ FILLER_0_21_150/a_36_472# 0.015502f
C5615 _136_ FILLER_0_17_142/a_572_375# 0.001371f
C5616 cal_count\[3\] FILLER_0_11_135/a_36_472# 0.005101f
C5617 net82 net22 1.960347f
C5618 FILLER_0_12_28/a_124_375# vdd 0.040988f
C5619 _053_ _151_ 0.538643f
C5620 _402_/a_1948_68# cal_count\[1\] 0.037053f
C5621 _028_ FILLER_0_5_72/a_484_472# 0.003042f
C5622 _428_/a_1308_423# _043_ 0.024052f
C5623 _205_/a_36_160# _047_ 0.013528f
C5624 net18 output30/a_224_472# 0.08667f
C5625 _412_/a_36_151# _082_ 0.016538f
C5626 net15 _424_/a_2665_112# 0.046592f
C5627 FILLER_0_12_20/a_484_472# net47 0.020293f
C5628 output33/a_224_472# output19/a_224_472# 0.115114f
C5629 _070_ _389_/a_36_148# 0.010534f
C5630 net34 FILLER_0_22_128/a_1828_472# 0.005158f
C5631 _052_ _424_/a_796_472# 0.002115f
C5632 _083_ FILLER_0_3_221/a_572_375# 0.001072f
C5633 _098_ _434_/a_1000_472# 0.00725f
C5634 _441_/a_448_472# vdd 0.007984f
C5635 _441_/a_36_151# vss 0.015116f
C5636 _235_/a_67_603# vdd 0.026582f
C5637 FILLER_0_16_107/a_572_375# net36 0.001706f
C5638 net49 trim_mask\[3\] 0.03723f
C5639 _086_ _268_/a_245_68# 0.001044f
C5640 _449_/a_2560_156# net55 0.004835f
C5641 net72 _452_/a_36_151# 0.040035f
C5642 _442_/a_2248_156# trim_mask\[3\] 0.003039f
C5643 result[1] _005_ 0.001478f
C5644 net15 _447_/a_2560_156# 0.001586f
C5645 _155_ net14 0.10433f
C5646 mask\[3\] FILLER_0_18_177/a_1468_375# 0.002924f
C5647 _016_ vss 0.069165f
C5648 ctln[6] ctln[5] 0.017291f
C5649 output47/a_224_472# net40 0.002339f
C5650 FILLER_0_15_228/a_124_375# vdd 0.013701f
C5651 _161_ cal_count\[3\] 0.047389f
C5652 _057_ _071_ 0.139904f
C5653 _238_/a_67_603# vdd 0.004498f
C5654 net63 _434_/a_2560_156# 0.014333f
C5655 FILLER_0_11_101/a_124_375# _120_ 0.008016f
C5656 net55 FILLER_0_17_72/a_932_472# 0.024922f
C5657 _440_/a_1000_472# vss 0.031704f
C5658 FILLER_0_19_142/a_124_375# vdd 0.022448f
C5659 FILLER_0_4_107/a_1468_375# trim_mask\[4\] 0.00157f
C5660 comp cal_count\[2\] 0.015029f
C5661 FILLER_0_4_185/a_124_375# vdd 0.02924f
C5662 _112_ _425_/a_36_151# 0.032941f
C5663 _053_ FILLER_0_7_72/a_2364_375# 0.015932f
C5664 net68 net67 0.147318f
C5665 _439_/a_36_151# vdd 0.095368f
C5666 _104_ FILLER_0_17_226/a_124_375# 0.024833f
C5667 FILLER_0_16_37/a_36_472# net72 0.005134f
C5668 _044_ vss 0.038421f
C5669 _132_ _334_/a_36_160# 0.026495f
C5670 net70 net36 0.066607f
C5671 _432_/a_1000_472# _091_ 0.026097f
C5672 _443_/a_2248_156# _170_ 0.068179f
C5673 FILLER_0_7_72/a_572_375# _028_ 0.003837f
C5674 _061_ _113_ 0.012561f
C5675 net1 _265_/a_244_68# 0.023821f
C5676 FILLER_0_19_47/a_572_375# vss 0.055293f
C5677 FILLER_0_19_47/a_36_472# vdd 0.072773f
C5678 FILLER_0_15_142/a_572_375# net36 0.006382f
C5679 trim_val\[4\] FILLER_0_3_172/a_572_375# 0.001076f
C5680 _000_ _083_ 0.017601f
C5681 _131_ FILLER_0_17_104/a_36_472# 0.004125f
C5682 _426_/a_36_151# FILLER_0_8_247/a_124_375# 0.059049f
C5683 _275_/a_224_472# _069_ 0.004466f
C5684 _118_ _122_ 0.046796f
C5685 _008_ _006_ 0.02963f
C5686 net20 _198_/a_67_603# 0.013603f
C5687 FILLER_0_16_73/a_484_472# cal_count\[1\] 0.001135f
C5688 vss FILLER_0_16_115/a_36_472# 0.003243f
C5689 _308_/a_848_380# FILLER_0_7_72/a_2724_472# 0.001797f
C5690 FILLER_0_6_47/a_1380_472# vss 0.001431f
C5691 FILLER_0_6_47/a_1828_472# vdd 0.002735f
C5692 FILLER_0_9_72/a_36_472# _453_/a_2665_112# 0.001167f
C5693 output21/a_224_472# net32 0.017976f
C5694 _316_/a_124_24# vss 0.00516f
C5695 _316_/a_848_380# vdd 0.048727f
C5696 _140_ _149_ 0.0088f
C5697 _175_ FILLER_0_15_72/a_124_375# 0.009573f
C5698 FILLER_0_4_144/a_572_375# net23 0.019114f
C5699 net39 vdd 0.2282f
C5700 _112_ net1 0.001653f
C5701 _444_/a_2560_156# _054_ 0.003269f
C5702 _412_/a_36_151# _265_/a_244_68# 0.072351f
C5703 output35/a_224_472# _204_/a_67_603# 0.012678f
C5704 vdd _039_ 0.219985f
C5705 _413_/a_1308_423# net21 0.065716f
C5706 _062_ _311_/a_692_473# 0.008632f
C5707 input4/a_36_68# vss 0.058179f
C5708 FILLER_0_10_37/a_124_375# net68 0.012617f
C5709 FILLER_0_21_125/a_124_375# vdd -0.010326f
C5710 _087_ _122_ 0.007241f
C5711 FILLER_0_17_72/a_3260_375# net14 0.040606f
C5712 _144_ _348_/a_257_69# 0.001978f
C5713 _156_ _160_ 0.299745f
C5714 _162_ _163_ 0.011497f
C5715 _014_ _123_ 0.050082f
C5716 _418_/a_448_472# _007_ 0.050316f
C5717 ctln[1] net82 0.001141f
C5718 FILLER_0_21_142/a_124_375# _433_/a_2665_112# 0.004834f
C5719 FILLER_0_15_205/a_124_375# net22 0.049201f
C5720 net16 _063_ 0.038576f
C5721 FILLER_0_8_247/a_124_375# FILLER_0_8_239/a_124_375# 0.003732f
C5722 net29 result[2] 0.001786f
C5723 net54 FILLER_0_18_107/a_3260_375# 0.001619f
C5724 net70 FILLER_0_14_123/a_124_375# 0.032077f
C5725 FILLER_0_22_86/a_36_472# net14 0.003007f
C5726 _091_ FILLER_0_19_171/a_1468_375# 0.002731f
C5727 mask\[4\] _098_ 0.041526f
C5728 net34 _299_/a_36_472# 0.003396f
C5729 _098_ net22 0.157058f
C5730 _072_ _116_ 0.283323f
C5731 output14/a_224_472# vdd 0.054725f
C5732 state\[0\] _323_/a_36_113# 0.016796f
C5733 _448_/a_1000_472# net59 0.007647f
C5734 mask\[3\] net80 0.02972f
C5735 _061_ _118_ 0.268815f
C5736 FILLER_0_10_78/a_572_375# vss 0.004588f
C5737 _427_/a_448_472# vss 0.040679f
C5738 _427_/a_1308_423# vdd 0.002814f
C5739 net68 FILLER_0_8_37/a_572_375# 0.011704f
C5740 _397_/a_36_472# _175_ 0.004667f
C5741 _132_ net36 0.029615f
C5742 _289_/a_36_472# _102_ 0.046918f
C5743 _086_ _120_ 0.408014f
C5744 _432_/a_2665_112# _139_ 0.004089f
C5745 _433_/a_1288_156# _022_ 0.001147f
C5746 net28 _192_/a_255_603# 0.003166f
C5747 FILLER_0_2_93/a_484_472# FILLER_0_2_101/a_36_472# 0.013277f
C5748 FILLER_0_3_221/a_484_472# net59 0.001655f
C5749 _257_/a_36_472# vdd -0.001779f
C5750 FILLER_0_11_78/a_572_375# _389_/a_36_148# 0.021545f
C5751 _093_ FILLER_0_18_177/a_3260_375# 0.002695f
C5752 net75 _316_/a_848_380# 0.044673f
C5753 _401_/a_36_68# _180_ 0.051459f
C5754 net54 _354_/a_257_69# 0.001135f
C5755 net15 FILLER_0_17_56/a_484_472# 0.001758f
C5756 vss FILLER_0_8_156/a_572_375# 0.007969f
C5757 vdd FILLER_0_8_156/a_36_472# 0.002891f
C5758 _068_ _122_ 0.096251f
C5759 _002_ FILLER_0_3_172/a_3260_375# 0.001683f
C5760 _119_ _120_ 0.036534f
C5761 _437_/a_2560_156# net14 0.00349f
C5762 net44 _450_/a_448_472# 0.050752f
C5763 _127_ cal_count\[3\] 0.306114f
C5764 _413_/a_2248_156# net21 0.009186f
C5765 mask\[4\] _433_/a_2248_156# 0.001082f
C5766 result[8] FILLER_0_23_290/a_36_472# 0.001414f
C5767 _144_ _340_/a_36_160# 0.008886f
C5768 _028_ _151_ 0.020076f
C5769 _449_/a_448_472# _067_ 0.0432f
C5770 FILLER_0_22_177/a_1380_472# _435_/a_36_151# 0.001723f
C5771 _163_ FILLER_0_6_79/a_36_472# 0.001789f
C5772 _114_ FILLER_0_10_94/a_484_472# 0.011954f
C5773 _033_ _444_/a_796_472# 0.0099f
C5774 _165_ _444_/a_2248_156# 0.006027f
C5775 net36 _282_/a_36_160# 0.002754f
C5776 FILLER_0_12_136/a_1380_472# cal_count\[3\] 0.00383f
C5777 _068_ _311_/a_2180_473# 0.001454f
C5778 net76 FILLER_0_6_177/a_124_375# 0.00227f
C5779 FILLER_0_9_223/a_124_375# _246_/a_36_68# 0.005308f
C5780 net2 net37 0.05083f
C5781 FILLER_0_14_81/a_36_472# net55 0.015878f
C5782 net73 _433_/a_36_151# 0.004541f
C5783 _370_/a_124_24# _152_ 0.069015f
C5784 _370_/a_848_380# _081_ 0.035068f
C5785 output34/a_224_472# net32 0.027498f
C5786 FILLER_0_16_57/a_1020_375# FILLER_0_17_64/a_124_375# 0.026339f
C5787 mask\[5\] _434_/a_36_151# 0.00104f
C5788 cal_count\[3\] _373_/a_438_68# 0.003743f
C5789 net60 _418_/a_36_151# 0.016348f
C5790 net60 _419_/a_1204_472# 0.023544f
C5791 net61 _419_/a_2665_112# 0.022394f
C5792 net50 net69 0.634381f
C5793 net52 _031_ 0.633473f
C5794 _011_ mask\[7\] 0.043474f
C5795 FILLER_0_7_72/a_2364_375# _028_ 0.003884f
C5796 _061_ _068_ 1.857322f
C5797 _289_/a_36_472# _198_/a_67_603# 0.027695f
C5798 _443_/a_1204_472# net69 0.002642f
C5799 cal_count\[3\] _071_ 0.214649f
C5800 trimb[3] vdd 0.283005f
C5801 net27 _425_/a_2248_156# 0.027078f
C5802 FILLER_0_5_172/a_36_472# net37 0.013857f
C5803 FILLER_0_10_78/a_1380_472# _077_ 0.001548f
C5804 FILLER_0_18_177/a_3172_472# vss 0.002639f
C5805 FILLER_0_18_2/a_484_472# output47/a_224_472# 0.00175f
C5806 FILLER_0_12_124/a_124_375# _131_ 0.07304f
C5807 FILLER_0_7_59/a_124_375# vdd -0.006113f
C5808 _130_ _118_ 0.053869f
C5809 FILLER_0_14_99/a_36_472# FILLER_0_13_100/a_36_472# 0.026657f
C5810 FILLER_0_12_28/a_124_375# cal_count\[0\] 0.001414f
C5811 net35 net23 0.04007f
C5812 _106_ _291_/a_36_160# 0.054237f
C5813 net35 FILLER_0_22_128/a_1916_375# 0.014552f
C5814 _178_ _408_/a_56_524# 0.014421f
C5815 net21 _202_/a_36_160# 0.09166f
C5816 FILLER_0_4_49/a_484_472# FILLER_0_3_54/a_36_472# 0.026657f
C5817 net20 FILLER_0_6_231/a_572_375# 0.01215f
C5818 net38 cal_count\[3\] 0.002225f
C5819 _079_ FILLER_0_5_198/a_484_472# 0.008167f
C5820 _335_/a_257_69# _043_ 0.001043f
C5821 vss FILLER_0_13_72/a_484_472# 0.008682f
C5822 _002_ vdd 0.152662f
C5823 net64 calibrate 0.096329f
C5824 FILLER_0_16_57/a_1380_472# vss 0.011192f
C5825 trim_mask\[1\] FILLER_0_6_47/a_572_375# 0.007164f
C5826 FILLER_0_9_142/a_124_375# _120_ 0.04442f
C5827 _303_/a_36_472# vss 0.011549f
C5828 _102_ vss 0.068703f
C5829 _114_ FILLER_0_12_136/a_1020_375# 0.006974f
C5830 FILLER_0_15_116/a_36_472# FILLER_0_17_104/a_1468_375# 0.001512f
C5831 _070_ FILLER_0_9_105/a_124_375# 0.017687f
C5832 _308_/a_848_380# vss 0.043591f
C5833 FILLER_0_22_86/a_36_472# _098_ 0.182093f
C5834 FILLER_0_7_146/a_36_472# _062_ 0.011622f
C5835 _091_ _113_ 0.006236f
C5836 _444_/a_1308_423# net17 0.028709f
C5837 _421_/a_36_151# _419_/a_36_151# 0.561555f
C5838 output22/a_224_472# net22 0.032714f
C5839 ctlp[0] vdd 0.08832f
C5840 net55 _451_/a_3129_107# 0.098091f
C5841 _065_ trim_val\[2\] 0.002278f
C5842 _428_/a_2665_112# FILLER_0_13_142/a_36_472# 0.003706f
C5843 fanout79/a_36_160# vss 0.002268f
C5844 _013_ FILLER_0_17_64/a_36_472# 0.001991f
C5845 net36 state\[1\] 0.004105f
C5846 _065_ _447_/a_796_472# 0.007495f
C5847 _119_ _227_/a_36_160# 0.01123f
C5848 net41 FILLER_0_23_44/a_36_472# 0.001116f
C5849 _093_ FILLER_0_19_111/a_484_472# 0.001009f
C5850 _140_ FILLER_0_19_155/a_484_472# 0.004155f
C5851 _005_ _094_ 0.162984f
C5852 net38 net40 1.103743f
C5853 _025_ _352_/a_49_472# 0.003933f
C5854 _431_/a_36_151# _131_ 0.03645f
C5855 _446_/a_796_472# _035_ 0.013039f
C5856 net81 _015_ 0.002818f
C5857 _070_ _370_/a_124_24# 0.00219f
C5858 FILLER_0_4_123/a_36_472# vss 0.004542f
C5859 FILLER_0_9_28/a_3260_375# vdd 0.017581f
C5860 net35 _025_ 0.02169f
C5861 FILLER_0_14_181/a_36_472# _043_ 0.008613f
C5862 _015_ _426_/a_2665_112# 0.018623f
C5863 result[4] FILLER_0_17_282/a_124_375# 0.018106f
C5864 _174_ _095_ 0.977766f
C5865 output11/a_224_472# net65 0.001529f
C5866 _386_/a_692_472# _169_ 0.004014f
C5867 _386_/a_848_380# _163_ 0.026484f
C5868 _098_ _437_/a_2560_156# 0.001174f
C5869 _039_ cal_count\[0\] 0.219667f
C5870 _417_/a_36_151# output30/a_224_472# 0.004902f
C5871 net42 vdd 0.178782f
C5872 net65 FILLER_0_3_172/a_932_472# 0.002604f
C5873 FILLER_0_5_128/a_36_472# net47 0.008459f
C5874 FILLER_0_21_125/a_572_375# net54 0.024701f
C5875 input4/a_36_68# net4 0.004679f
C5876 FILLER_0_11_78/a_124_375# _120_ 0.014367f
C5877 net41 output7/a_224_472# 0.003942f
C5878 _359_/a_636_68# _062_ 0.001578f
C5879 FILLER_0_9_72/a_36_472# vdd 0.109576f
C5880 FILLER_0_9_72/a_1468_375# vss 0.013085f
C5881 result[9] net78 0.015761f
C5882 net27 _426_/a_1308_423# 0.00384f
C5883 FILLER_0_10_78/a_1468_375# _114_ 0.01836f
C5884 _171_ FILLER_0_10_94/a_36_472# 0.001514f
C5885 _172_ FILLER_0_10_94/a_124_375# 0.003341f
C5886 _451_/a_1040_527# net14 0.029964f
C5887 net55 FILLER_0_13_72/a_572_375# 0.005919f
C5888 net35 net33 1.594925f
C5889 _359_/a_36_488# vdd 0.083138f
C5890 _078_ vdd 0.181583f
C5891 FILLER_0_16_57/a_484_472# net55 0.001797f
C5892 _182_ vss 0.068928f
C5893 fanout51/a_36_113# FILLER_0_11_64/a_36_472# 0.001396f
C5894 _277_/a_36_160# _099_ 0.001628f
C5895 FILLER_0_12_50/a_124_375# _120_ 0.002753f
C5896 _198_/a_67_603# vss 0.003647f
C5897 output8/a_224_472# FILLER_0_3_221/a_1468_375# 0.032044f
C5898 net50 _165_ 0.056964f
C5899 _188_ vss 0.032923f
C5900 FILLER_0_6_90/a_36_472# FILLER_0_4_91/a_124_375# 0.001188f
C5901 net58 net82 0.022761f
C5902 net43 FILLER_0_20_15/a_124_375# 0.005925f
C5903 net57 FILLER_0_13_142/a_1468_375# 0.011369f
C5904 _320_/a_1120_472# _043_ 0.002242f
C5905 net18 _417_/a_1000_472# 0.056791f
C5906 net57 fanout53/a_36_160# 0.009946f
C5907 output46/a_224_472# net17 0.082914f
C5908 fanout66/a_36_113# _030_ 0.038252f
C5909 net26 FILLER_0_18_37/a_932_472# 0.002613f
C5910 net53 FILLER_0_16_154/a_124_375# 0.003458f
C5911 FILLER_0_15_282/a_572_375# output30/a_224_472# 0.029138f
C5912 net62 _416_/a_36_151# 0.054002f
C5913 vss _416_/a_1308_423# 0.001962f
C5914 output11/a_224_472# net59 0.002364f
C5915 result[5] result[9] 0.064058f
C5916 fanout67/a_36_160# vss 0.005344f
C5917 net67 FILLER_0_8_37/a_36_472# 0.001479f
C5918 vdd clkc 0.190259f
C5919 _408_/a_1336_472# _186_ 0.010089f
C5920 FILLER_0_13_142/a_572_375# _043_ 0.009328f
C5921 mask\[2\] FILLER_0_16_154/a_1020_375# 0.020485f
C5922 FILLER_0_15_142/a_124_375# _427_/a_36_151# 0.059049f
C5923 FILLER_0_14_91/a_124_375# _176_ 0.019567f
C5924 _431_/a_2665_112# FILLER_0_16_154/a_124_375# 0.006271f
C5925 trim[4] net44 0.188184f
C5926 _116_ state\[1\] 0.693219f
C5927 FILLER_0_12_124/a_124_375# _126_ 0.02249f
C5928 net48 _425_/a_36_151# 0.020568f
C5929 _176_ FILLER_0_10_94/a_36_472# 0.009089f
C5930 _140_ FILLER_0_22_128/a_3260_375# 0.003524f
C5931 fanout49/a_36_160# _160_ 0.009662f
C5932 mask\[0\] FILLER_0_15_212/a_1020_375# 0.001158f
C5933 FILLER_0_7_72/a_2276_472# vdd 0.004035f
C5934 _069_ _248_/a_36_68# 0.058746f
C5935 ctln[7] FILLER_0_0_96/a_36_472# 0.01317f
C5936 output8/a_224_472# net20 0.084627f
C5937 net34 output18/a_224_472# 0.17524f
C5938 _335_/a_49_472# _138_ 0.005957f
C5939 FILLER_0_11_109/a_36_472# _120_ 0.014554f
C5940 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_484_472# 0.001723f
C5941 net81 _069_ 0.034401f
C5942 vss trim[2] 0.026644f
C5943 trim_val\[0\] _220_/a_67_603# 0.005346f
C5944 _050_ vss 0.26237f
C5945 ctlp[1] FILLER_0_24_274/a_572_375# 0.002408f
C5946 FILLER_0_21_28/a_2276_472# vdd 0.002733f
C5947 FILLER_0_21_28/a_1828_472# vss -0.001894f
C5948 FILLER_0_6_90/a_124_375# vdd 0.020992f
C5949 FILLER_0_22_128/a_2812_375# _146_ 0.001336f
C5950 _178_ FILLER_0_17_38/a_572_375# 0.031538f
C5951 _057_ _311_/a_1660_473# 0.004637f
C5952 FILLER_0_11_135/a_36_472# _120_ 0.012562f
C5953 net35 _436_/a_1000_472# 0.009213f
C5954 _075_ _074_ 0.058521f
C5955 FILLER_0_5_109/a_124_375# _365_/a_36_68# 0.004633f
C5956 _443_/a_2665_112# net22 0.00621f
C5957 _163_ _365_/a_36_68# 0.004035f
C5958 _086_ FILLER_0_5_117/a_36_472# 0.042352f
C5959 FILLER_0_7_59/a_484_472# _439_/a_36_151# 0.001061f
C5960 FILLER_0_11_64/a_36_472# net51 0.009015f
C5961 _126_ FILLER_0_11_101/a_484_472# 0.001488f
C5962 cal_itt\[2\] FILLER_0_3_221/a_36_472# 0.003825f
C5963 net48 net1 0.006424f
C5964 _129_ _133_ 0.080636f
C5965 _372_/a_170_472# _076_ 0.049892f
C5966 _372_/a_2034_472# _133_ 0.001257f
C5967 _069_ _060_ 0.538161f
C5968 _126_ _090_ 0.003538f
C5969 _004_ _192_/a_67_603# 0.020219f
C5970 FILLER_0_11_282/a_124_375# vdd 0.026044f
C5971 _178_ _043_ 0.130207f
C5972 net25 _051_ 0.090798f
C5973 FILLER_0_7_104/a_932_472# _151_ 0.002092f
C5974 _233_/a_36_160# net40 0.001875f
C5975 FILLER_0_21_125/a_124_375# _433_/a_36_151# 0.059049f
C5976 FILLER_0_7_72/a_36_472# net50 0.011974f
C5977 net55 cal_count\[3\] 0.005157f
C5978 net67 net47 0.126281f
C5979 _253_/a_36_68# FILLER_0_3_221/a_1468_375# 0.014131f
C5980 _163_ FILLER_0_5_148/a_124_375# 0.001706f
C5981 FILLER_0_6_177/a_484_472# _163_ 0.002256f
C5982 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_124_375# 0.012222f
C5983 FILLER_0_8_24/a_484_472# FILLER_0_8_37/a_36_472# 0.001963f
C5984 _057_ _056_ 0.167928f
C5985 FILLER_0_17_72/a_3260_375# _131_ 0.004986f
C5986 _119_ FILLER_0_5_117/a_36_472# 0.002628f
C5987 trim_mask\[0\] FILLER_0_10_94/a_572_375# 0.003359f
C5988 output33/a_224_472# output18/a_224_472# 0.111946f
C5989 _068_ _160_ 0.003424f
C5990 _412_/a_36_151# net48 0.001091f
C5991 _106_ mask\[3\] 0.249479f
C5992 _053_ _062_ 0.185944f
C5993 _425_/a_36_151# net19 0.009499f
C5994 FILLER_0_19_142/a_124_375# FILLER_0_19_134/a_124_375# 0.003732f
C5995 _178_ _185_ 0.979797f
C5996 vdd FILLER_0_14_235/a_572_375# 0.006167f
C5997 vss FILLER_0_14_235/a_124_375# 0.002686f
C5998 FILLER_0_5_128/a_484_472# vss 0.004051f
C5999 net81 FILLER_0_15_212/a_36_472# 0.003945f
C6000 trim_mask\[1\] FILLER_0_6_79/a_124_375# 0.0042f
C6001 _093_ _199_/a_36_160# 0.05226f
C6002 FILLER_0_14_181/a_124_375# _138_ 0.001663f
C6003 net20 _223_/a_36_160# 0.066119f
C6004 FILLER_0_16_107/a_484_472# _451_/a_36_151# 0.027244f
C6005 net68 trim_val\[1\] 0.006974f
C6006 FILLER_0_15_180/a_484_472# vss 0.001207f
C6007 FILLER_0_5_206/a_124_375# net37 0.005485f
C6008 FILLER_0_18_2/a_124_375# net44 0.051228f
C6009 net66 FILLER_0_3_54/a_36_472# 0.008174f
C6010 _334_/a_36_160# vdd 0.041716f
C6011 output12/a_224_472# _037_ 0.00827f
C6012 FILLER_0_20_177/a_932_472# _434_/a_36_151# 0.001723f
C6013 _111_ FILLER_0_18_76/a_36_472# 0.006706f
C6014 FILLER_0_5_72/a_572_375# _440_/a_36_151# 0.035849f
C6015 _086_ _151_ 0.002442f
C6016 _164_ FILLER_0_6_47/a_572_375# 0.010099f
C6017 net79 _044_ 0.013636f
C6018 output21/a_224_472# _105_ 0.034631f
C6019 _149_ net14 0.102004f
C6020 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1380_472# 0.003468f
C6021 net1 net19 0.024768f
C6022 net67 FILLER_0_6_47/a_124_375# 0.005516f
C6023 net74 _125_ 0.071757f
C6024 FILLER_0_17_226/a_124_375# _008_ 0.006576f
C6025 _093_ FILLER_0_19_155/a_124_375# 0.001864f
C6026 _132_ FILLER_0_18_107/a_1916_375# 0.019011f
C6027 net55 net40 0.043962f
C6028 trim[1] _444_/a_36_151# 0.001391f
C6029 ctlp[7] vdd 0.481613f
C6030 _074_ FILLER_0_5_164/a_484_472# 0.003556f
C6031 _095_ FILLER_0_15_72/a_484_472# 0.002306f
C6032 output36/a_224_472# net36 0.009109f
C6033 output13/a_224_472# FILLER_0_0_130/a_124_375# 0.00363f
C6034 ctln[1] clk 0.551557f
C6035 net16 _444_/a_2560_156# 0.010829f
C6036 FILLER_0_9_28/a_124_375# net17 0.009179f
C6037 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_484_472# 0.026657f
C6038 FILLER_0_18_2/a_484_472# net38 0.003391f
C6039 mask\[0\] _335_/a_665_69# 0.001711f
C6040 FILLER_0_4_107/a_1380_472# vss 0.004455f
C6041 _307_/a_234_472# _085_ 0.001966f
C6042 _103_ net77 0.004691f
C6043 cal_count\[3\] net23 0.045417f
C6044 FILLER_0_8_24/a_484_472# net47 0.042018f
C6045 net67 _450_/a_836_156# 0.008805f
C6046 FILLER_0_12_2/a_572_375# net44 0.041552f
C6047 FILLER_0_12_20/a_484_472# vdd 0.003108f
C6048 _431_/a_36_151# FILLER_0_15_116/a_572_375# 0.001543f
C6049 _058_ FILLER_0_8_156/a_124_375# 0.006325f
C6050 FILLER_0_18_2/a_1828_472# _452_/a_1353_112# 0.001313f
C6051 _412_/a_36_151# net19 0.03393f
C6052 _435_/a_2248_156# vdd 0.00571f
C6053 FILLER_0_11_101/a_572_375# FILLER_0_10_107/a_36_472# 0.001684f
C6054 _049_ _146_ 0.042698f
C6055 _093_ net55 0.182194f
C6056 FILLER_0_18_2/a_1380_472# vss -0.001894f
C6057 _013_ _424_/a_2665_112# 0.001222f
C6058 cal_count\[1\] _040_ 0.019478f
C6059 FILLER_0_9_72/a_1380_472# _439_/a_36_151# 0.001723f
C6060 net75 _411_/a_448_472# 0.072712f
C6061 input1/a_36_113# net2 0.018839f
C6062 vss FILLER_0_6_231/a_572_375# 0.057794f
C6063 vdd FILLER_0_6_231/a_36_472# 0.014642f
C6064 net67 FILLER_0_9_60/a_124_375# 0.003083f
C6065 _122_ FILLER_0_5_172/a_36_472# 0.003007f
C6066 _434_/a_36_151# _348_/a_49_472# 0.017459f
C6067 _140_ _098_ 0.647503f
C6068 FILLER_0_20_87/a_124_375# vdd 0.008846f
C6069 _081_ _261_/a_36_160# 0.049069f
C6070 _126_ _038_ 0.031198f
C6071 net25 vdd 0.195306f
C6072 comp FILLER_0_12_2/a_36_472# 0.003875f
C6073 net63 FILLER_0_18_177/a_2724_472# 0.001857f
C6074 net49 _168_ 0.031157f
C6075 FILLER_0_20_193/a_572_375# _205_/a_36_160# 0.002828f
C6076 _440_/a_36_151# _160_ 0.002966f
C6077 _174_ net74 0.00916f
C6078 _394_/a_56_524# vss 0.003797f
C6079 fanout55/a_36_160# FILLER_0_13_80/a_36_472# 0.003699f
C6080 net36 vdd 0.939735f
C6081 FILLER_0_10_78/a_1020_375# _115_ 0.064761f
C6082 net26 FILLER_0_23_44/a_484_472# 0.003796f
C6083 _044_ _416_/a_2665_112# 0.01372f
C6084 FILLER_0_19_28/a_572_375# vss 0.002775f
C6085 FILLER_0_19_28/a_36_472# vdd 0.052986f
C6086 FILLER_0_16_57/a_36_472# FILLER_0_17_56/a_124_375# 0.001723f
C6087 _050_ FILLER_0_22_128/a_1020_375# 0.002647f
C6088 state\[1\] _225_/a_36_160# 0.0535f
C6089 FILLER_0_15_2/a_36_472# vss 0.002136f
C6090 net23 _169_ 0.00151f
C6091 cal input1/a_36_113# 0.025739f
C6092 net25 FILLER_0_23_60/a_36_472# 0.005618f
C6093 _098_ FILLER_0_21_150/a_36_472# 0.002964f
C6094 net16 _131_ 0.001308f
C6095 _053_ FILLER_0_7_72/a_3260_375# 0.071059f
C6096 FILLER_0_21_28/a_2276_472# _424_/a_36_151# 0.001723f
C6097 net80 _333_/a_36_160# 0.001594f
C6098 net76 _080_ 0.03728f
C6099 _127_ _120_ 0.198577f
C6100 _174_ cal_count\[1\] 0.081252f
C6101 FILLER_0_20_193/a_572_375# mask\[6\] 0.001262f
C6102 _093_ net23 0.042838f
C6103 _073_ cal_itt\[0\] 0.211566f
C6104 net64 FILLER_0_9_270/a_572_375# 0.017924f
C6105 _126_ _076_ 0.005517f
C6106 _140_ _433_/a_2248_156# 0.003337f
C6107 _015_ net64 1.212892f
C6108 _267_/a_36_472# _113_ 0.014178f
C6109 _285_/a_36_472# _094_ 0.045394f
C6110 net38 _445_/a_448_472# 0.023336f
C6111 net18 rstn 0.015842f
C6112 _016_ _428_/a_1308_423# 0.00107f
C6113 net81 FILLER_0_15_235/a_36_472# 0.001855f
C6114 net44 net17 0.046636f
C6115 net82 FILLER_0_3_172/a_2276_472# 0.007729f
C6116 net82 _386_/a_1084_68# 0.001068f
C6117 FILLER_0_15_116/a_484_472# _136_ 0.002712f
C6118 FILLER_0_4_107/a_484_472# _369_/a_36_68# 0.001049f
C6119 FILLER_0_4_107/a_1020_375# _158_ 0.003535f
C6120 _144_ _207_/a_67_603# 0.064623f
C6121 FILLER_0_1_98/a_124_375# vdd 0.036865f
C6122 fanout57/a_36_113# net82 0.017696f
C6123 net46 vss 0.110452f
C6124 FILLER_0_10_256/a_36_472# FILLER_0_10_247/a_36_472# 0.001963f
C6125 FILLER_0_4_185/a_36_472# vdd 0.122463f
C6126 net18 _418_/a_1000_472# 0.050485f
C6127 _413_/a_36_151# FILLER_0_4_197/a_36_472# 0.001512f
C6128 FILLER_0_5_54/a_1020_375# _440_/a_36_151# 0.059049f
C6129 output34/a_224_472# _105_ 0.007506f
C6130 net62 result[1] 0.061866f
C6131 _431_/a_2248_156# net53 0.003335f
C6132 net61 net78 1.588656f
C6133 FILLER_0_14_123/a_124_375# vdd 0.034436f
C6134 output19/a_224_472# vss 0.048948f
C6135 _431_/a_36_151# _137_ 0.011412f
C6136 FILLER_0_9_28/a_2276_472# vdd 0.003276f
C6137 FILLER_0_9_28/a_2364_375# _053_ 0.029866f
C6138 FILLER_0_21_150/a_124_375# _433_/a_2665_112# 0.029834f
C6139 _086_ _375_/a_960_497# 0.001454f
C6140 FILLER_0_21_206/a_36_472# net33 0.001447f
C6141 mask\[4\] FILLER_0_18_171/a_124_375# 0.008445f
C6142 mask\[4\] _137_ 0.086066f
C6143 net55 FILLER_0_21_60/a_484_472# 0.098472f
C6144 FILLER_0_19_55/a_124_375# vdd 0.035786f
C6145 _052_ FILLER_0_18_61/a_36_472# 0.001508f
C6146 FILLER_0_18_76/a_484_472# vss 0.005065f
C6147 _165_ _054_ 0.001337f
C6148 _056_ cal_count\[3\] 0.186969f
C6149 _050_ mask\[7\] 0.128172f
C6150 net40 _381_/a_36_472# 0.020876f
C6151 _410_/a_36_68# vss 0.02717f
C6152 output8/a_224_472# cal_itt\[1\] 0.003894f
C6153 FILLER_0_18_107/a_932_472# FILLER_0_17_104/a_1380_472# 0.026657f
C6154 net72 _394_/a_244_524# 0.001083f
C6155 net62 _429_/a_2665_112# 0.02887f
C6156 trim_mask\[1\] FILLER_0_4_91/a_484_472# 0.002806f
C6157 _423_/a_2665_112# vss 0.016881f
C6158 net54 FILLER_0_19_111/a_36_472# 0.003467f
C6159 mask\[4\] FILLER_0_19_171/a_36_472# 0.001776f
C6160 FILLER_0_2_101/a_124_375# net14 0.0239f
C6161 net57 state\[2\] 1.25275f
C6162 _050_ _148_ 0.002456f
C6163 _104_ _420_/a_2665_112# 0.053555f
C6164 _116_ vdd 0.399137f
C6165 _149_ _098_ 0.398643f
C6166 _106_ FILLER_0_17_218/a_124_375# 0.004655f
C6167 net41 FILLER_0_21_28/a_1020_375# 0.010649f
C6168 result[5] net61 0.092275f
C6169 FILLER_0_20_169/a_124_375# vss 0.017635f
C6170 FILLER_0_20_169/a_36_472# vdd 0.010522f
C6171 _239_/a_36_160# net17 0.014703f
C6172 net15 _453_/a_448_472# 0.040851f
C6173 _013_ FILLER_0_17_56/a_484_472# 0.002659f
C6174 _131_ FILLER_0_14_107/a_1380_472# 0.01797f
C6175 _392_/a_36_68# cal_count\[3\] 0.003072f
C6176 FILLER_0_22_128/a_2276_472# vdd 0.00565f
C6177 FILLER_0_22_128/a_1828_472# vss 0.009137f
C6178 net53 _043_ 0.053033f
C6179 result[4] vdd 0.205815f
C6180 _422_/a_1204_472# _109_ 0.001807f
C6181 FILLER_0_5_109/a_124_375# _154_ 0.058658f
C6182 net55 FILLER_0_13_80/a_124_375# 0.069951f
C6183 _432_/a_2248_156# vdd 0.02369f
C6184 _178_ _402_/a_1296_93# 0.062418f
C6185 _070_ FILLER_0_10_107/a_36_472# 0.013252f
C6186 output8/a_224_472# vss 0.076244f
C6187 _163_ _154_ 0.190662f
C6188 _030_ vdd 0.244909f
C6189 fanout49/a_36_160# _156_ 0.002871f
C6190 net57 trim_mask\[4\] 0.259381f
C6191 result[9] net60 0.251903f
C6192 _086_ _267_/a_1568_472# 0.002143f
C6193 _442_/a_1204_472# vdd 0.001128f
C6194 FILLER_0_6_79/a_124_375# _164_ 0.061565f
C6195 _053_ FILLER_0_6_47/a_1380_472# 0.004472f
C6196 FILLER_0_18_2/a_3260_375# vss 0.026159f
C6197 _069_ mask\[1\] 0.029447f
C6198 _036_ net17 0.153479f
C6199 trim_mask\[1\] vss 0.449335f
C6200 net47 _382_/a_224_472# 0.001795f
C6201 _424_/a_2248_156# FILLER_0_21_60/a_124_375# 0.001068f
C6202 FILLER_0_15_290/a_124_375# result[3] 0.020277f
C6203 _445_/a_2665_112# net17 0.006445f
C6204 _428_/a_1204_472# net74 0.009712f
C6205 mask\[5\] _205_/a_36_160# 0.003775f
C6206 output29/a_224_472# _044_ 0.087528f
C6207 net29 mask\[1\] 0.023266f
C6208 _421_/a_36_151# _010_ 0.015107f
C6209 _065_ net52 0.017184f
C6210 cal_itt\[2\] cal_itt\[0\] 0.011453f
C6211 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_36_472# 0.026657f
C6212 output37/a_224_472# _425_/a_2248_156# 0.00114f
C6213 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_124_375# 0.012222f
C6214 _308_/a_1084_68# net14 0.002892f
C6215 fanout55/a_36_160# _067_ 0.126784f
C6216 net55 FILLER_0_18_76/a_572_375# 0.002278f
C6217 net1 fanout58/a_36_160# 0.060243f
C6218 ctlp[3] net61 0.007397f
C6219 FILLER_0_3_54/a_124_375# _164_ 0.008654f
C6220 net58 FILLER_0_9_270/a_484_472# 0.061043f
C6221 output46/a_224_472# trimb[3] 0.050924f
C6222 fanout82/a_36_113# vss 0.023533f
C6223 _253_/a_36_68# cal_itt\[1\] 0.039692f
C6224 _425_/a_1308_423# vdd 0.021703f
C6225 net81 output27/a_224_472# 0.011872f
C6226 net20 FILLER_0_12_220/a_572_375# 0.007386f
C6227 fanout79/a_36_160# net79 0.011193f
C6228 net65 trim_val\[4\] 0.015549f
C6229 FILLER_0_9_282/a_36_472# vdd 0.106034f
C6230 FILLER_0_9_282/a_572_375# vss 0.058599f
C6231 FILLER_0_14_50/a_124_375# _174_ 0.033245f
C6232 mask\[7\] _435_/a_1204_472# 0.007888f
C6233 net70 FILLER_0_14_107/a_124_375# 0.029975f
C6234 vdd FILLER_0_22_107/a_484_472# 0.035591f
C6235 mask\[5\] mask\[6\] 0.140269f
C6236 vss FILLER_0_22_107/a_36_472# 0.001514f
C6237 _092_ FILLER_0_18_209/a_484_472# 0.006303f
C6238 _411_/a_1308_423# net65 0.004122f
C6239 FILLER_0_15_212/a_36_472# mask\[1\] 0.006865f
C6240 FILLER_0_7_72/a_3260_375# _028_ 0.003505f
C6241 _248_/a_36_68# _090_ 0.041161f
C6242 _292_/a_36_160# _204_/a_67_603# 0.003478f
C6243 _147_ _049_ 0.001131f
C6244 net73 FILLER_0_17_133/a_124_375# 0.022541f
C6245 _059_ net47 0.00606f
C6246 _070_ FILLER_0_10_94/a_124_375# 0.008294f
C6247 _223_/a_36_160# vss 0.007187f
C6248 _050_ _436_/a_1308_423# 0.022688f
C6249 output35/a_224_472# net33 0.170613f
C6250 net31 net61 0.053131f
C6251 _431_/a_36_151# net56 0.001371f
C6252 _371_/a_36_113# _152_ 0.001083f
C6253 cal_count\[3\] FILLER_0_12_196/a_124_375# 0.007717f
C6254 FILLER_0_16_57/a_1020_375# _131_ 0.012481f
C6255 FILLER_0_7_195/a_124_375# _055_ 0.001597f
C6256 _056_ net59 0.001756f
C6257 net41 vss 0.810444f
C6258 ctlp[2] _011_ 0.101324f
C6259 mask\[4\] net56 0.006006f
C6260 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_572_375# 0.086635f
C6261 FILLER_0_4_177/a_484_472# net22 0.006506f
C6262 FILLER_0_9_28/a_3172_472# vss 0.001977f
C6263 FILLER_0_15_72/a_484_472# cal_count\[1\] 0.013337f
C6264 _083_ _080_ 0.043927f
C6265 output25/a_224_472# _213_/a_67_603# 0.032497f
C6266 _117_ vdd 0.050188f
C6267 FILLER_0_4_107/a_36_472# _153_ 0.042459f
C6268 FILLER_0_4_107/a_932_472# _154_ 0.017867f
C6269 fanout72/a_36_113# _043_ 0.017862f
C6270 FILLER_0_14_99/a_36_472# vss 0.003598f
C6271 _253_/a_36_68# vss 0.002481f
C6272 net52 fanout51/a_36_113# 0.036773f
C6273 _346_/a_49_472# net23 0.022558f
C6274 FILLER_0_9_223/a_36_472# state\[0\] 0.002846f
C6275 _090_ _060_ 0.396493f
C6276 _345_/a_36_160# _145_ 0.001141f
C6277 trim_val\[4\] net59 0.062701f
C6278 _115_ _058_ 0.038308f
C6279 _248_/a_36_68# net22 0.002193f
C6280 FILLER_0_3_172/a_124_375# net22 0.01308f
C6281 _074_ _014_ 0.001557f
C6282 net81 net22 0.064261f
C6283 _115_ _315_/a_36_68# 0.001683f
C6284 net75 _425_/a_1308_423# 0.034219f
C6285 _077_ _129_ 0.08682f
C6286 _003_ _074_ 0.00476f
C6287 net79 _416_/a_1308_423# 0.030119f
C6288 net39 net44 0.0112f
C6289 FILLER_0_8_247/a_124_375# vss 0.002674f
C6290 _322_/a_848_380# _070_ 0.006182f
C6291 FILLER_0_8_247/a_572_375# vdd -0.007963f
C6292 output47/a_224_472# _185_ 0.001177f
C6293 mask\[0\] _136_ 0.025838f
C6294 _060_ net22 0.533421f
C6295 net76 FILLER_0_2_177/a_124_375# 0.00439f
C6296 FILLER_0_15_10/a_124_375# FILLER_0_15_2/a_572_375# 0.012001f
C6297 _421_/a_36_151# vdd -0.053849f
C6298 _132_ FILLER_0_14_107/a_124_375# 0.003315f
C6299 mask\[0\] net21 0.050431f
C6300 net44 _039_ 0.15647f
C6301 _074_ net21 0.186175f
C6302 mask\[9\] FILLER_0_20_98/a_36_472# 0.005917f
C6303 FILLER_0_14_107/a_36_472# _043_ 0.001661f
C6304 mask\[5\] _009_ 0.001095f
C6305 _225_/a_36_160# vdd 0.058272f
C6306 _448_/a_2248_156# _037_ 0.027079f
C6307 _444_/a_1204_472# net40 0.017496f
C6308 _308_/a_124_24# vdd 0.011014f
C6309 net63 _435_/a_1000_472# 0.002536f
C6310 net79 _283_/a_36_472# 0.010249f
C6311 FILLER_0_20_193/a_36_472# vss 0.001978f
C6312 FILLER_0_20_193/a_484_472# vdd 0.00749f
C6313 net19 net30 0.311153f
C6314 output19/a_224_472# mask\[7\] 0.001181f
C6315 _442_/a_36_151# net13 0.009343f
C6316 _118_ _113_ 0.005092f
C6317 _446_/a_36_151# net40 0.015376f
C6318 _081_ _001_ 0.012101f
C6319 FILLER_0_9_105/a_484_472# vss 0.004412f
C6320 _116_ _279_/a_244_68# 0.001752f
C6321 _415_/a_36_151# _426_/a_36_151# 0.002121f
C6322 net52 net51 0.091698f
C6323 _095_ FILLER_0_13_142/a_36_472# 0.001782f
C6324 net22 net12 0.032084f
C6325 FILLER_0_5_198/a_36_472# net59 0.059378f
C6326 _074_ _070_ 0.102481f
C6327 _139_ _098_ 0.026578f
C6328 cal_itt\[3\] _062_ 0.009718f
C6329 _004_ FILLER_0_10_256/a_36_472# 0.00402f
C6330 _414_/a_1000_472# _053_ 0.029433f
C6331 ctln[4] ctln[5] 0.031901f
C6332 _235_/a_67_603# _036_ 0.043345f
C6333 net55 _120_ 0.001054f
C6334 vss _433_/a_3041_156# 0.001287f
C6335 FILLER_0_18_139/a_932_472# vss 0.041568f
C6336 FILLER_0_18_139/a_1380_472# vdd 0.005855f
C6337 trim_val\[1\] net47 0.34878f
C6338 mask\[5\] FILLER_0_19_187/a_572_375# 0.005529f
C6339 net49 _440_/a_2665_112# 0.025303f
C6340 _064_ _445_/a_36_151# 0.03209f
C6341 _447_/a_36_151# net68 0.040925f
C6342 trim_mask\[2\] trim_mask\[1\] 0.002186f
C6343 net64 FILLER_0_15_235/a_36_472# 0.046292f
C6344 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_124_375# 0.026339f
C6345 FILLER_0_16_154/a_1020_375# vss 0.001453f
C6346 FILLER_0_16_154/a_1468_375# vdd 0.017574f
C6347 _322_/a_848_380# FILLER_0_9_142/a_36_472# 0.011591f
C6348 _431_/a_36_151# FILLER_0_18_107/a_2276_472# 0.002799f
C6349 FILLER_0_7_195/a_36_472# vss 0.002568f
C6350 net62 _094_ 0.04063f
C6351 FILLER_0_15_235/a_36_472# mask\[1\] 0.009316f
C6352 net75 _263_/a_224_472# 0.004396f
C6353 FILLER_0_7_104/a_932_472# _062_ 0.001184f
C6354 mask\[7\] FILLER_0_22_128/a_1828_472# 0.004503f
C6355 net75 FILLER_0_8_247/a_572_375# 0.003962f
C6356 _130_ _321_/a_170_472# 0.001018f
C6357 net16 _453_/a_36_151# 0.001634f
C6358 net38 FILLER_0_8_24/a_124_375# 0.001013f
C6359 FILLER_0_15_150/a_36_472# _136_ 0.002967f
C6360 _079_ net22 0.039221f
C6361 FILLER_0_7_104/a_1020_375# vdd 0.010571f
C6362 net31 output31/a_224_472# 0.002146f
C6363 trim_val\[2\] _167_ 0.011787f
C6364 _318_/a_224_472# _124_ 0.001288f
C6365 net73 FILLER_0_18_107/a_3260_375# 0.001629f
C6366 _431_/a_2560_156# net73 0.001018f
C6367 trimb[1] FILLER_0_18_2/a_1916_375# 0.001855f
C6368 output8/a_224_472# net4 0.015359f
C6369 trim[0] _034_ 0.044322f
C6370 net26 FILLER_0_21_28/a_1468_375# 0.041169f
C6371 FILLER_0_18_107/a_1916_375# vdd 0.018831f
C6372 trim_val\[1\] FILLER_0_6_47/a_124_375# 0.002577f
C6373 net39 _445_/a_2665_112# 0.002831f
C6374 _317_/a_36_113# FILLER_0_7_233/a_124_375# 0.03227f
C6375 net15 _052_ 0.001074f
C6376 net52 FILLER_0_9_72/a_1020_375# 0.00799f
C6377 trim_mask\[3\] vdd 0.233305f
C6378 _164_ vss 0.597051f
C6379 _207_/a_67_603# FILLER_0_22_128/a_3172_472# 0.005759f
C6380 _093_ _046_ 0.061989f
C6381 _432_/a_36_151# FILLER_0_15_180/a_36_472# 0.002018f
C6382 _120_ net23 0.147166f
C6383 _086_ _062_ 0.066419f
C6384 net54 FILLER_0_22_128/a_1468_375# 0.004731f
C6385 _433_/a_1000_472# _145_ 0.004227f
C6386 FILLER_0_18_37/a_1468_375# vdd 0.021186f
C6387 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_484_472# 0.013276f
C6388 net67 vdd 0.638702f
C6389 FILLER_0_16_89/a_572_375# vdd 0.005006f
C6390 FILLER_0_8_107/a_36_472# FILLER_0_7_104/a_484_472# 0.026657f
C6391 _292_/a_36_160# _201_/a_67_603# 0.003917f
C6392 ctln[2] FILLER_0_1_266/a_124_375# 0.047145f
C6393 _027_ net71 0.057875f
C6394 _131_ FILLER_0_17_64/a_124_375# 0.005913f
C6395 FILLER_0_3_204/a_36_472# _088_ 0.004381f
C6396 _317_/a_36_113# vdd 0.054289f
C6397 state\[2\] FILLER_0_13_142/a_1380_472# 0.019965f
C6398 FILLER_0_24_274/a_36_472# vdd 0.107635f
C6399 FILLER_0_24_274/a_1468_375# vss 0.060201f
C6400 _077_ net57 0.025864f
C6401 _072_ _247_/a_36_160# 0.005008f
C6402 cal net8 0.271166f
C6403 _098_ net14 0.061285f
C6404 FILLER_0_5_72/a_1380_472# vss 0.004538f
C6405 _178_ FILLER_0_16_37/a_124_375# 0.036901f
C6406 _119_ _062_ 0.080398f
C6407 FILLER_0_4_144/a_36_472# _152_ 0.008211f
C6408 FILLER_0_4_144/a_484_472# _081_ 0.001145f
C6409 calibrate _123_ 0.016296f
C6410 ctlp[4] mask\[6\] 0.003054f
C6411 _029_ _153_ 0.023421f
C6412 _077_ _219_/a_36_160# 0.01438f
C6413 _104_ result[8] 0.00201f
C6414 FILLER_0_17_161/a_124_375# _098_ 0.002013f
C6415 FILLER_0_9_28/a_124_375# net42 0.007403f
C6416 net61 net60 0.059237f
C6417 _390_/a_36_68# vss 0.002334f
C6418 _128_ _126_ 0.008298f
C6419 mask\[3\] FILLER_0_17_218/a_572_375# 0.015907f
C6420 _025_ FILLER_0_22_107/a_124_375# 0.001891f
C6421 _000_ FILLER_0_3_221/a_1020_375# 0.016709f
C6422 FILLER_0_10_28/a_36_472# net51 0.00703f
C6423 result[8] _422_/a_1308_423# 0.001356f
C6424 FILLER_0_10_37/a_124_375# vdd 0.048346f
C6425 _413_/a_36_151# FILLER_0_3_172/a_2364_375# 0.059049f
C6426 output22/a_224_472# _435_/a_36_151# 0.12978f
C6427 mask\[7\] _299_/a_36_472# 0.033949f
C6428 _187_ _173_ 0.03421f
C6429 net4 _223_/a_36_160# 0.020711f
C6430 _053_ fanout67/a_36_160# 0.05724f
C6431 _004_ output28/a_224_472# 0.024204f
C6432 cal_count\[2\] vss 0.361185f
C6433 _068_ _118_ 1.374452f
C6434 _070_ _124_ 0.114614f
C6435 _099_ FILLER_0_14_235/a_572_375# 0.013281f
C6436 _069_ FILLER_0_11_142/a_484_472# 0.005789f
C6437 FILLER_0_18_209/a_36_472# vss 0.005442f
C6438 FILLER_0_18_209/a_484_472# vdd 0.00367f
C6439 net18 _416_/a_36_151# 0.027435f
C6440 FILLER_0_8_24/a_36_472# vss 0.001239f
C6441 FILLER_0_8_24/a_484_472# vdd 0.009032f
C6442 _091_ FILLER_0_13_228/a_36_472# 0.001826f
C6443 FILLER_0_18_107/a_932_472# mask\[9\] 0.005296f
C6444 net15 mask\[9\] 0.128816f
C6445 FILLER_0_3_78/a_572_375# _160_ 0.003506f
C6446 output27/a_224_472# net64 0.04953f
C6447 net19 FILLER_0_14_263/a_36_472# 0.135429f
C6448 net52 _163_ 0.00157f
C6449 FILLER_0_12_220/a_572_375# vss 0.007775f
C6450 FILLER_0_12_220/a_1020_375# vdd -0.014642f
C6451 output13/a_224_472# _448_/a_2248_156# 0.009013f
C6452 net57 _066_ 0.069098f
C6453 ctlp[7] net24 0.078667f
C6454 net55 FILLER_0_18_37/a_124_375# 0.005899f
C6455 result[7] _420_/a_2665_112# 0.039448f
C6456 FILLER_0_4_107/a_1468_375# _160_ 0.028099f
C6457 net20 state\[0\] 0.396139f
C6458 net15 FILLER_0_17_72/a_932_472# 0.001122f
C6459 net75 _317_/a_36_113# 0.030797f
C6460 FILLER_0_17_72/a_124_375# vdd 0.0132f
C6461 _079_ _076_ 0.001575f
C6462 FILLER_0_8_37/a_572_375# vdd 0.013575f
C6463 FILLER_0_8_37/a_124_375# vss 0.00252f
C6464 _115_ net52 0.022268f
C6465 _091_ net31 0.001465f
C6466 _430_/a_448_472# mask\[2\] 0.045973f
C6467 FILLER_0_11_124/a_36_472# vss 0.002545f
C6468 net23 FILLER_0_16_154/a_124_375# 0.002689f
C6469 net47 FILLER_0_4_91/a_572_375# 0.008167f
C6470 result[8] net22 0.278936f
C6471 _370_/a_848_380# net23 0.001196f
C6472 net27 FILLER_0_10_256/a_124_375# 0.006216f
C6473 net38 _450_/a_36_151# 0.035458f
C6474 ctlp[4] _009_ 0.004522f
C6475 output18/a_224_472# vss 0.086897f
C6476 _449_/a_2665_112# _038_ 0.024406f
C6477 net65 net18 0.879399f
C6478 FILLER_0_21_142/a_124_375# net35 0.00123f
C6479 net80 FILLER_0_22_177/a_572_375# 0.005202f
C6480 trim[0] FILLER_0_3_2/a_124_375# 0.020708f
C6481 net16 _165_ 0.021744f
C6482 FILLER_0_15_59/a_124_375# vdd 0.017243f
C6483 _392_/a_244_472# _067_ 0.001893f
C6484 net38 _043_ 0.117134f
C6485 net57 net37 0.091923f
C6486 _227_/a_36_160# net23 0.055152f
C6487 net25 net24 0.031854f
C6488 FILLER_0_7_59/a_36_472# net68 0.050931f
C6489 _348_/a_49_472# mask\[6\] 0.005525f
C6490 net27 net62 0.008623f
C6491 mask\[1\] net22 0.029526f
C6492 net74 FILLER_0_13_142/a_36_472# 0.003568f
C6493 _392_/a_36_68# _120_ 0.001738f
C6494 _437_/a_36_151# vss 0.006865f
C6495 _437_/a_448_472# vdd 0.010432f
C6496 trim_mask\[2\] _164_ 1.859062f
C6497 FILLER_0_10_28/a_36_472# net6 0.038613f
C6498 output19/a_224_472# _295_/a_36_472# 0.003896f
C6499 _424_/a_448_472# FILLER_0_18_37/a_1020_375# 0.001674f
C6500 _105_ _422_/a_36_151# 0.030571f
C6501 trim_mask\[4\] FILLER_0_2_111/a_1020_375# 0.02806f
C6502 _098_ FILLER_0_15_205/a_124_375# 0.009558f
C6503 _328_/a_36_113# FILLER_0_11_101/a_484_472# 0.001826f
C6504 FILLER_0_12_124/a_124_375# net74 0.049113f
C6505 net36 _099_ 0.325141f
C6506 _238_/a_67_603# output15/a_224_472# 0.019027f
C6507 _447_/a_1308_423# _164_ 0.001422f
C6508 net18 net59 0.695067f
C6509 net15 _440_/a_1308_423# 0.015192f
C6510 output25/a_224_472# mask\[8\] 0.015742f
C6511 vdd result[3] 0.181788f
C6512 _360_/a_36_160# vss 0.028817f
C6513 _081_ _316_/a_124_24# 0.011421f
C6514 net44 clkc 0.184915f
C6515 trim_val\[2\] _446_/a_2665_112# 0.012621f
C6516 FILLER_0_6_177/a_124_375# net47 0.002925f
C6517 FILLER_0_4_99/a_36_472# _030_ 0.002699f
C6518 _411_/a_36_151# ctln[1] 0.018351f
C6519 _112_ _316_/a_848_380# 0.022235f
C6520 _305_/a_36_159# calibrate 0.003505f
C6521 output31/a_224_472# net60 0.216716f
C6522 _445_/a_2248_156# _444_/a_36_151# 0.001081f
C6523 _308_/a_848_380# trim_mask\[0\] 0.035693f
C6524 net54 _433_/a_1308_423# 0.004372f
C6525 FILLER_0_23_44/a_1020_375# vdd -0.014642f
C6526 fanout54/a_36_160# FILLER_0_18_139/a_1020_375# 0.031033f
C6527 _438_/a_796_472# net71 0.00514f
C6528 _077_ _453_/a_448_472# 0.057515f
C6529 _177_ vss 0.074896f
C6530 _446_/a_36_151# trim[3] 0.00699f
C6531 FILLER_0_7_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001723f
C6532 FILLER_0_5_72/a_124_375# _029_ 0.010208f
C6533 output23/a_224_472# _049_ 0.001034f
C6534 FILLER_0_20_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001543f
C6535 _091_ _429_/a_1204_472# 0.024554f
C6536 _394_/a_728_93# FILLER_0_15_72/a_572_375# 0.02852f
C6537 net72 FILLER_0_15_59/a_124_375# 0.022905f
C6538 _131_ net14 0.037705f
C6539 _132_ _134_ 0.029512f
C6540 net58 net81 0.375649f
C6541 FILLER_0_23_60/a_124_375# FILLER_0_23_44/a_1468_375# 0.012001f
C6542 net15 net35 0.01797f
C6543 net63 FILLER_0_20_193/a_572_375# 0.015818f
C6544 FILLER_0_17_38/a_484_472# vss 0.001229f
C6545 vdd _450_/a_1040_527# 0.005529f
C6546 _074_ net9 0.002862f
C6547 _098_ _433_/a_2248_156# 0.034774f
C6548 net17 _450_/a_3129_107# 0.004255f
C6549 net73 _020_ 0.057454f
C6550 FILLER_0_16_73/a_124_375# FILLER_0_17_72/a_124_375# 0.026339f
C6551 net62 _043_ 0.00426f
C6552 net47 _452_/a_1353_112# 0.003681f
C6553 FILLER_0_16_107/a_124_375# _136_ 0.00661f
C6554 mask\[9\] _437_/a_2665_112# 0.014146f
C6555 net26 _424_/a_1308_423# 0.001179f
C6556 net19 _417_/a_2665_112# 0.042961f
C6557 _136_ FILLER_0_16_115/a_124_375# 0.006372f
C6558 FILLER_0_4_144/a_572_375# trim_mask\[4\] 0.014071f
C6559 net34 _207_/a_67_603# 0.008585f
C6560 input3/a_36_113# cal_count\[2\] 0.00555f
C6561 _005_ _044_ 0.50767f
C6562 _015_ FILLER_0_10_247/a_36_472# 0.007508f
C6563 _382_/a_224_472# vdd 0.001663f
C6564 _058_ FILLER_0_9_105/a_36_472# 0.011426f
C6565 fanout75/a_36_113# net59 0.00817f
C6566 _093_ FILLER_0_18_61/a_36_472# 0.004039f
C6567 net16 _095_ 0.042842f
C6568 FILLER_0_19_171/a_1380_472# FILLER_0_19_187/a_36_472# 0.013277f
C6569 FILLER_0_5_164/a_484_472# _163_ 0.029894f
C6570 FILLER_0_10_37/a_124_375# cal_count\[0\] 0.016543f
C6571 FILLER_0_7_72/a_3172_472# _219_/a_36_160# 0.035111f
C6572 FILLER_0_12_136/a_124_375# _127_ 0.004013f
C6573 _093_ FILLER_0_17_104/a_1468_375# 0.010965f
C6574 _448_/a_36_151# vdd 0.133302f
C6575 net57 en_co_clk 0.195533f
C6576 _315_/a_36_68# _121_ 0.031617f
C6577 FILLER_0_5_117/a_124_375# _153_ 0.079379f
C6578 FILLER_0_5_128/a_572_375# _152_ 0.00813f
C6579 result[1] net18 0.056799f
C6580 FILLER_0_24_63/a_36_472# vss 0.008178f
C6581 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_36_472# 0.026657f
C6582 net55 FILLER_0_17_38/a_572_375# 0.007646f
C6583 FILLER_0_14_107/a_124_375# vdd 0.013327f
C6584 _059_ vdd 0.161836f
C6585 output48/a_224_472# vdd 0.038342f
C6586 _161_ _062_ 0.046903f
C6587 FILLER_0_22_177/a_124_375# vdd 0.001293f
C6588 FILLER_0_4_197/a_124_375# vdd 0.011327f
C6589 net4 FILLER_0_12_220/a_572_375# 0.019052f
C6590 FILLER_0_3_221/a_124_375# vss 0.034009f
C6591 FILLER_0_7_104/a_124_375# _058_ 0.006125f
C6592 net36 FILLER_0_15_212/a_124_375# 0.004391f
C6593 FILLER_0_9_28/a_572_375# net40 0.001406f
C6594 _016_ net53 0.180698f
C6595 _075_ FILLER_0_7_195/a_124_375# 0.008178f
C6596 net55 _043_ 0.053191f
C6597 mask\[5\] _343_/a_49_472# 0.002228f
C6598 FILLER_0_17_200/a_572_375# mask\[3\] 0.013879f
C6599 _414_/a_1000_472# cal_itt\[3\] 0.08528f
C6600 net74 _038_ 0.055774f
C6601 _375_/a_36_68# vdd 0.010344f
C6602 net5 vdd 0.516129f
C6603 _144_ _208_/a_36_160# 0.00717f
C6604 mask\[4\] FILLER_0_18_177/a_1828_472# 0.014226f
C6605 FILLER_0_18_107/a_1916_375# _433_/a_36_151# 0.002709f
C6606 _443_/a_1456_156# net23 0.001009f
C6607 FILLER_0_5_54/a_572_375# _029_ 0.00494f
C6608 _293_/a_36_472# net31 0.005692f
C6609 FILLER_0_20_177/a_1380_472# vss 0.004504f
C6610 FILLER_0_18_100/a_124_375# _438_/a_2665_112# 0.010688f
C6611 net34 _108_ 0.297364f
C6612 FILLER_0_16_255/a_36_472# _045_ 0.001653f
C6613 FILLER_0_4_197/a_932_472# net76 0.003693f
C6614 fanout50/a_36_160# net49 0.030626f
C6615 _440_/a_2665_112# net47 0.014066f
C6616 _414_/a_1000_472# _081_ 0.006091f
C6617 _119_ FILLER_0_8_156/a_572_375# 0.01739f
C6618 net35 FILLER_0_22_86/a_1468_375# 0.010438f
C6619 mask\[8\] FILLER_0_22_86/a_36_472# 0.012471f
C6620 net52 _442_/a_796_472# 0.004871f
C6621 _093_ FILLER_0_17_200/a_124_375# 0.00419f
C6622 net57 _395_/a_1044_488# 0.002526f
C6623 FILLER_0_21_142/a_484_472# net23 0.005353f
C6624 net62 FILLER_0_14_263/a_124_375# 0.037111f
C6625 FILLER_0_21_142/a_484_472# FILLER_0_22_128/a_1916_375# 0.001543f
C6626 FILLER_0_18_2/a_3172_472# net55 0.00602f
C6627 net78 _420_/a_2248_156# 0.001534f
C6628 net50 _029_ 0.025102f
C6629 _429_/a_448_472# _043_ 0.003615f
C6630 state\[0\] vss 0.126943f
C6631 _095_ FILLER_0_14_107/a_1380_472# 0.011439f
C6632 _000_ vdd 0.215988f
C6633 _126_ net14 0.238336f
C6634 FILLER_0_18_177/a_1468_375# vdd 0.024167f
C6635 net55 _175_ 0.142124f
C6636 _128_ _426_/a_2665_112# 0.025626f
C6637 _072_ _311_/a_66_473# 0.031716f
C6638 _350_/a_49_472# mask\[6\] 0.033488f
C6639 net44 FILLER_0_15_2/a_484_472# 0.047161f
C6640 FILLER_0_2_101/a_36_472# _156_ 0.001487f
C6641 net82 FILLER_0_3_212/a_36_472# 0.011542f
C6642 _431_/a_448_472# _136_ 0.064724f
C6643 ctln[5] _448_/a_1204_472# 0.005186f
C6644 _308_/a_124_24# FILLER_0_9_72/a_1380_472# 0.003595f
C6645 _070_ FILLER_0_8_156/a_124_375# 0.004329f
C6646 mask\[5\] net63 0.112147f
C6647 _131_ FILLER_0_17_56/a_36_472# 0.001491f
C6648 _136_ _451_/a_2225_156# 0.01289f
C6649 _053_ trim_mask\[1\] 0.110786f
C6650 _128_ _060_ 0.022833f
C6651 FILLER_0_7_59/a_484_472# net67 0.03109f
C6652 FILLER_0_14_91/a_572_375# vss 0.054783f
C6653 FILLER_0_14_91/a_36_472# vdd 0.08739f
C6654 net75 output48/a_224_472# 0.070114f
C6655 vss FILLER_0_10_94/a_484_472# 0.001244f
C6656 net15 FILLER_0_13_72/a_572_375# 0.003021f
C6657 mask\[8\] _437_/a_2560_156# 0.001171f
C6658 _422_/a_2560_156# _009_ 0.002551f
C6659 net23 _043_ 0.042095f
C6660 _453_/a_2248_156# vdd 0.010767f
C6661 FILLER_0_16_57/a_484_472# net15 0.008573f
C6662 _415_/a_2560_156# net18 0.010318f
C6663 _095_ _451_/a_1040_527# 0.002316f
C6664 net69 FILLER_0_3_78/a_124_375# 0.004201f
C6665 _417_/a_796_472# _006_ 0.014427f
C6666 _072_ _374_/a_244_472# 0.001816f
C6667 _012_ FILLER_0_21_60/a_572_375# 0.011991f
C6668 _230_/a_652_68# _062_ 0.001144f
C6669 _141_ FILLER_0_16_154/a_1020_375# 0.003441f
C6670 mask\[3\] FILLER_0_16_154/a_484_472# 0.002067f
C6671 result[7] result[8] 0.201281f
C6672 _414_/a_36_151# _074_ 0.070632f
C6673 _178_ _182_ 0.067534f
C6674 _429_/a_2665_112# FILLER_0_15_212/a_1468_375# 0.010688f
C6675 net69 FILLER_0_2_101/a_124_375# 0.015032f
C6676 result[8] FILLER_0_23_282/a_484_472# 0.001908f
C6677 _414_/a_1000_472# _089_ 0.001754f
C6678 FILLER_0_20_2/a_124_375# vss 0.002737f
C6679 FILLER_0_20_2/a_572_375# vdd 0.010844f
C6680 FILLER_0_4_123/a_124_375# _152_ 0.039668f
C6681 FILLER_0_11_101/a_36_472# cal_count\[3\] 0.005101f
C6682 FILLER_0_5_212/a_36_472# vdd 0.107657f
C6683 FILLER_0_5_212/a_124_375# vss 0.006344f
C6684 _176_ net36 0.336675f
C6685 FILLER_0_18_177/a_2724_472# net21 0.048803f
C6686 _438_/a_2560_156# vdd 0.001166f
C6687 _438_/a_2665_112# vss 0.001389f
C6688 net53 _427_/a_448_472# 0.047356f
C6689 _444_/a_1308_423# net67 0.021684f
C6690 _373_/a_1458_68# _113_ 0.001257f
C6691 trim_val\[1\] vdd 0.173304f
C6692 result[9] _420_/a_2560_156# 0.002295f
C6693 FILLER_0_1_266/a_572_375# vdd 0.030477f
C6694 trim_mask\[1\] FILLER_0_5_88/a_36_472# 0.038642f
C6695 mask\[5\] output21/a_224_472# 0.009585f
C6696 _139_ _137_ 0.093639f
C6697 FILLER_0_8_127/a_124_375# _062_ 0.046401f
C6698 net3 _190_/a_36_160# 0.013324f
C6699 _430_/a_36_151# FILLER_0_18_177/a_3172_472# 0.001512f
C6700 net7 net40 0.025164f
C6701 net57 _122_ 0.034045f
C6702 _127_ _062_ 0.020537f
C6703 net16 ctln[9] 0.07797f
C6704 net75 _000_ 0.096899f
C6705 output9/a_224_472# net18 0.114757f
C6706 net38 _033_ 0.03598f
C6707 output19/a_224_472# ctlp[2] 0.04607f
C6708 _091_ _273_/a_36_68# 0.00155f
C6709 _413_/a_36_151# net76 0.084453f
C6710 _074_ _084_ 0.110937f
C6711 _450_/a_3129_107# _039_ 0.012762f
C6712 _308_/a_692_472# trim_mask\[0\] 0.004377f
C6713 _057_ state\[2\] 0.054838f
C6714 fanout57/a_36_113# FILLER_0_3_172/a_124_375# 0.006548f
C6715 net80 vdd 1.045288f
C6716 _261_/a_36_160# net23 0.005015f
C6717 _130_ _129_ 0.021732f
C6718 _402_/a_728_93# _401_/a_36_68# 0.002178f
C6719 _087_ FILLER_0_5_172/a_36_472# 0.00443f
C6720 FILLER_0_21_206/a_124_375# net22 0.05301f
C6721 _413_/a_1000_472# _002_ 0.006249f
C6722 _276_/a_36_160# _291_/a_36_160# 0.239422f
C6723 _024_ FILLER_0_22_177/a_124_375# 0.005166f
C6724 _340_/a_36_160# vss 0.029871f
C6725 trimb[1] _452_/a_2225_156# 0.004072f
C6726 FILLER_0_12_136/a_1468_375# vdd 0.026145f
C6727 FILLER_0_12_136/a_1020_375# vss 0.018233f
C6728 _144_ FILLER_0_18_107/a_2364_375# 0.002388f
C6729 net21 _047_ 0.048701f
C6730 net15 cal_count\[3\] 0.045013f
C6731 _182_ FILLER_0_18_37/a_1380_472# 0.004074f
C6732 net53 _451_/a_2449_156# 0.015332f
C6733 net57 _061_ 0.127011f
C6734 net58 net64 0.590523f
C6735 _423_/a_796_472# _012_ 0.015809f
C6736 _013_ _052_ 0.284735f
C6737 net19 _418_/a_2665_112# 0.040822f
C6738 FILLER_0_17_104/a_932_472# net14 0.002113f
C6739 net73 FILLER_0_19_111/a_36_472# 0.001412f
C6740 net69 _158_ 0.033459f
C6741 mask\[9\] net71 0.344312f
C6742 _159_ vss 0.102545f
C6743 _116_ _176_ 0.067051f
C6744 _105_ _204_/a_255_603# 0.002146f
C6745 _008_ net64 0.001427f
C6746 _429_/a_36_151# _138_ 0.002064f
C6747 FILLER_0_3_172/a_3172_472# net22 0.010714f
C6748 _306_/a_36_68# _116_ 0.00183f
C6749 net79 FILLER_0_12_220/a_572_375# 0.010889f
C6750 _168_ vdd 0.083621f
C6751 _152_ _163_ 0.05157f
C6752 output26/a_224_472# vdd 0.047141f
C6753 FILLER_0_17_72/a_932_472# net71 0.001418f
C6754 net62 _417_/a_2248_156# 0.005537f
C6755 _412_/a_2248_156# fanout58/a_36_160# 0.005856f
C6756 _424_/a_2665_112# _012_ 0.01024f
C6757 _092_ _106_ 0.140596f
C6758 FILLER_0_4_123/a_124_375# _070_ 0.001677f
C6759 net48 _316_/a_848_380# 0.026413f
C6760 ctln[2] net76 0.001008f
C6761 net16 cal_count\[1\] 0.007291f
C6762 net41 FILLER_0_10_28/a_124_375# 0.003909f
C6763 FILLER_0_18_53/a_36_472# vss 0.001471f
C6764 FILLER_0_18_53/a_484_472# vdd 0.002358f
C6765 _430_/a_2248_156# _091_ 0.053571f
C6766 FILLER_0_17_161/a_124_375# _137_ 0.016092f
C6767 FILLER_0_18_76/a_124_375# _438_/a_36_151# 0.001252f
C6768 FILLER_0_10_78/a_1468_375# vss 0.054053f
C6769 net35 FILLER_0_22_177/a_932_472# 0.00643f
C6770 FILLER_0_22_86/a_1380_472# net71 0.011277f
C6771 output26/a_224_472# FILLER_0_23_60/a_36_472# 0.003292f
C6772 _247_/a_36_160# vdd 0.060423f
C6773 net20 FILLER_0_15_228/a_36_472# 0.020589f
C6774 FILLER_0_8_263/a_124_375# FILLER_0_8_247/a_1468_375# 0.012001f
C6775 cal_count\[3\] _186_ 0.012453f
C6776 FILLER_0_21_28/a_124_375# vdd 0.014155f
C6777 _028_ trim_mask\[1\] 0.148182f
C6778 net69 net14 0.056927f
C6779 FILLER_0_3_172/a_2812_375# vdd -0.012025f
C6780 _052_ FILLER_0_21_28/a_2812_375# 0.002388f
C6781 _067_ _172_ 0.010195f
C6782 FILLER_0_5_128/a_484_472# _081_ 0.00169f
C6783 net4 FILLER_0_3_221/a_124_375# 0.015788f
C6784 _132_ _436_/a_36_151# 0.00162f
C6785 _438_/a_1308_423# net14 0.005201f
C6786 output12/a_224_472# net59 0.015069f
C6787 FILLER_0_3_204/a_36_472# net65 0.001777f
C6788 _076_ _269_/a_36_472# 0.001618f
C6789 FILLER_0_13_212/a_36_472# _043_ 0.011752f
C6790 _093_ FILLER_0_18_107/a_932_472# 0.008683f
C6791 FILLER_0_2_93/a_484_472# FILLER_0_0_96/a_124_375# 0.001338f
C6792 _131_ _372_/a_170_472# 0.002967f
C6793 _093_ net15 0.145303f
C6794 _079_ FILLER_0_3_172/a_2276_472# 0.00261f
C6795 _412_/a_2560_156# net1 0.005618f
C6796 FILLER_0_12_2/a_36_472# vss 0.003757f
C6797 FILLER_0_8_263/a_124_375# _426_/a_36_151# 0.001252f
C6798 _444_/a_448_472# net47 0.030563f
C6799 _098_ FILLER_0_15_212/a_932_472# 0.011837f
C6800 _094_ net18 0.468109f
C6801 _363_/a_36_68# _151_ 0.020916f
C6802 _013_ mask\[9\] 0.011224f
C6803 _233_/a_36_160# _033_ 0.017573f
C6804 _063_ _165_ 0.021839f
C6805 _005_ _416_/a_1308_423# 0.020096f
C6806 FILLER_0_16_255/a_36_472# _287_/a_36_472# 0.004546f
C6807 output13/a_224_472# net13 0.058196f
C6808 _053_ FILLER_0_7_104/a_572_375# 0.005239f
C6809 _129_ _160_ 0.001631f
C6810 _430_/a_448_472# vss 0.003371f
C6811 _036_ _030_ 0.430683f
C6812 vdd FILLER_0_4_91/a_572_375# 0.019853f
C6813 output27/a_224_472# FILLER_0_9_290/a_36_472# 0.001711f
C6814 _447_/a_2665_112# net69 0.002067f
C6815 FILLER_0_4_99/a_124_375# net47 0.001409f
C6816 trimb[0] FILLER_0_20_2/a_36_472# 0.005458f
C6817 net82 net69 0.005307f
C6818 _445_/a_2248_156# net49 0.029744f
C6819 result[8] FILLER_0_24_290/a_36_472# 0.004676f
C6820 net19 _316_/a_848_380# 0.00558f
C6821 net81 _139_ 0.001762f
C6822 ctlp[2] _299_/a_36_472# 0.012937f
C6823 _267_/a_1792_472# _055_ 0.003058f
C6824 state\[0\] net4 0.13193f
C6825 mask\[8\] _140_ 0.003375f
C6826 ctln[5] FILLER_0_1_192/a_124_375# 0.001391f
C6827 _160_ _034_ 0.00905f
C6828 _053_ _164_ 0.058788f
C6829 FILLER_0_22_86/a_932_472# _149_ 0.001205f
C6830 FILLER_0_22_86/a_36_472# _026_ 0.001503f
C6831 FILLER_0_7_162/a_36_472# _062_ 0.016683f
C6832 net52 FILLER_0_5_72/a_932_472# 0.008749f
C6833 trimb[2] net43 0.011999f
C6834 mask\[3\] mask\[2\] 0.077703f
C6835 _432_/a_796_472# net80 0.007731f
C6836 FILLER_0_3_204/a_36_472# net59 0.001606f
C6837 _432_/a_1308_423# _093_ 0.016365f
C6838 net20 _291_/a_36_160# 0.002375f
C6839 net80 _024_ 0.064854f
C6840 mask\[0\] _429_/a_1308_423# 0.019225f
C6841 net55 FILLER_0_18_53/a_124_375# 0.011674f
C6842 net72 FILLER_0_18_53/a_484_472# 0.001067f
C6843 _256_/a_716_497# calibrate 0.001066f
C6844 net51 _450_/a_2449_156# 0.008215f
C6845 FILLER_0_2_111/a_932_472# vss -0.001894f
C6846 FILLER_0_2_111/a_1380_472# vdd 0.002688f
C6847 _321_/a_170_472# _118_ 0.034852f
C6848 _134_ vdd 0.482157f
C6849 _016_ _127_ 0.01898f
C6850 _070_ _163_ 1.884485f
C6851 _043_ FILLER_0_12_196/a_124_375# 0.003935f
C6852 FILLER_0_20_177/a_1020_375# _098_ 0.013949f
C6853 _428_/a_2665_112# _131_ 0.006081f
C6854 _128_ net64 0.291788f
C6855 fanout71/a_36_113# mask\[9\] 0.044939f
C6856 _103_ _418_/a_448_472# 0.002678f
C6857 state\[2\] cal_count\[3\] 0.005312f
C6858 ctlp[4] output21/a_224_472# 0.052556f
C6859 fanout62/a_36_160# vss 0.01343f
C6860 _115_ _070_ 0.890903f
C6861 _136_ FILLER_0_15_180/a_36_472# 0.006924f
C6862 FILLER_0_5_88/a_36_472# _164_ 0.011718f
C6863 net35 net71 0.042275f
C6864 FILLER_0_5_128/a_124_375# net74 0.013683f
C6865 FILLER_0_5_206/a_36_472# net22 0.049294f
C6866 _412_/a_2665_112# vdd 0.014403f
C6867 net63 FILLER_0_20_177/a_932_472# 0.004375f
C6868 fanout49/a_36_160# FILLER_0_3_78/a_572_375# 0.00805f
C6869 _078_ FILLER_0_4_213/a_572_375# 0.02957f
C6870 _086_ _321_/a_3662_472# 0.002598f
C6871 _414_/a_2248_156# FILLER_0_5_212/a_36_472# 0.035805f
C6872 _415_/a_36_151# vss 0.003124f
C6873 net34 _435_/a_2665_112# 0.009214f
C6874 output34/a_224_472# net30 0.002189f
C6875 net41 _445_/a_2560_156# 0.002221f
C6876 _093_ FILLER_0_17_72/a_2812_375# 0.019521f
C6877 _315_/a_244_497# _059_ 0.00101f
C6878 net56 FILLER_0_17_161/a_124_375# 0.001108f
C6879 FILLER_0_23_60/a_124_375# vdd 0.031398f
C6880 _031_ _153_ 0.009316f
C6881 FILLER_0_6_177/a_124_375# vdd 0.017329f
C6882 net15 FILLER_0_21_60/a_484_472# 0.001552f
C6883 _428_/a_36_151# FILLER_0_13_100/a_124_375# 0.023595f
C6884 net20 net76 0.021613f
C6885 FILLER_0_5_72/a_1380_472# FILLER_0_5_88/a_36_472# 0.013277f
C6886 mask\[4\] _145_ 0.340415f
C6887 net81 _429_/a_1000_472# 0.011018f
C6888 net64 FILLER_0_12_236/a_124_375# 0.043517f
C6889 net63 FILLER_0_18_177/a_572_375# 0.004407f
C6890 mask\[4\] FILLER_0_19_195/a_124_375# 0.006236f
C6891 _441_/a_1000_472# _168_ 0.036305f
C6892 FILLER_0_9_28/a_1380_472# _054_ 0.004017f
C6893 FILLER_0_24_96/a_36_472# ctlp[7] 0.001551f
C6894 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_36_472# 0.002296f
C6895 net15 _394_/a_1336_472# 0.01144f
C6896 FILLER_0_18_171/a_124_375# _098_ 0.032114f
C6897 _137_ _098_ 0.07262f
C6898 _411_/a_1000_472# _000_ 0.023042f
C6899 _431_/a_2560_156# net36 0.001858f
C6900 net27 FILLER_0_9_270/a_124_375# 0.079454f
C6901 _114_ _072_ 0.078148f
C6902 _444_/a_2665_112# FILLER_0_6_37/a_124_375# 0.005477f
C6903 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_36_472# 0.086742f
C6904 cal_count\[3\] FILLER_0_11_78/a_36_472# 0.031399f
C6905 _098_ FILLER_0_19_171/a_36_472# 0.021559f
C6906 net20 _108_ 0.125627f
C6907 FILLER_0_16_89/a_36_472# net36 0.010907f
C6908 net60 _420_/a_2248_156# 0.035104f
C6909 _428_/a_36_151# net70 0.040167f
C6910 _115_ FILLER_0_9_142/a_36_472# 0.00336f
C6911 _091_ net57 0.006076f
C6912 net50 _220_/a_67_603# 0.005566f
C6913 mask\[8\] _149_ 0.0498f
C6914 _074_ calibrate 0.046632f
C6915 _144_ _132_ 0.185339f
C6916 _098_ _438_/a_1308_423# 0.004124f
C6917 _126_ _131_ 0.626666f
C6918 net7 trim[3] 0.044017f
C6919 _188_ FILLER_0_12_50/a_124_375# 0.00157f
C6920 _326_/a_36_160# _115_ 0.051266f
C6921 FILLER_0_2_111/a_572_375# _158_ 0.031641f
C6922 FILLER_0_7_195/a_124_375# net21 0.007906f
C6923 net54 FILLER_0_20_98/a_124_375# 0.001639f
C6924 net82 FILLER_0_3_172/a_124_375# 0.011418f
C6925 FILLER_0_0_266/a_124_375# rstn 0.073089f
C6926 FILLER_0_24_96/a_36_472# net25 0.040228f
C6927 _452_/a_1353_112# vdd 0.008539f
C6928 net81 net82 0.063498f
C6929 net44 net67 0.08001f
C6930 output20/a_224_472# _422_/a_36_151# 0.053592f
C6931 _260_/a_36_68# FILLER_0_3_221/a_1380_472# 0.001652f
C6932 _080_ FILLER_0_3_221/a_1020_375# 0.001414f
C6933 _058_ FILLER_0_10_94/a_36_472# 0.009346f
C6934 net52 FILLER_0_5_54/a_1380_472# 0.00179f
C6935 net17 _452_/a_1293_527# 0.001011f
C6936 _128_ net74 0.121254f
C6937 trim_mask\[4\] _169_ 0.042442f
C6938 FILLER_0_9_223/a_124_375# _077_ 0.008762f
C6939 FILLER_0_17_72/a_3172_472# vdd 0.002712f
C6940 FILLER_0_7_146/a_124_375# _059_ 0.029514f
C6941 _028_ FILLER_0_7_104/a_572_375# 0.003664f
C6942 trim_mask\[2\] FILLER_0_4_91/a_124_375# 0.003591f
C6943 output38/a_224_472# trim[1] 0.003114f
C6944 _077_ _057_ 0.584179f
C6945 FILLER_0_21_142/a_572_375# vss 0.097474f
C6946 net60 _421_/a_2560_156# 0.001951f
C6947 FILLER_0_15_116/a_572_375# _131_ 0.051323f
C6948 _440_/a_2665_112# FILLER_0_4_91/a_36_472# 0.007491f
C6949 _028_ _164_ 0.019799f
C6950 _038_ _389_/a_36_148# 0.003749f
C6951 net27 net18 0.092379f
C6952 net57 _428_/a_2248_156# 0.022587f
C6953 _091_ FILLER_0_15_212/a_1380_472# 0.002787f
C6954 result[7] _103_ 0.298427f
C6955 _115_ FILLER_0_11_78/a_572_375# 0.034089f
C6956 net43 net40 0.018193f
C6957 output44/a_224_472# net40 0.006489f
C6958 _062_ net23 0.061239f
C6959 net31 _419_/a_2665_112# 0.004446f
C6960 _106_ vdd 0.232973f
C6961 _132_ _428_/a_36_151# 0.013691f
C6962 fanout59/a_36_160# net59 0.021522f
C6963 FILLER_0_6_37/a_124_375# _160_ 0.04948f
C6964 FILLER_0_17_72/a_1468_375# net36 0.047507f
C6965 FILLER_0_12_28/a_36_472# vss 0.003004f
C6966 _359_/a_244_68# _059_ 0.002986f
C6967 _028_ FILLER_0_5_72/a_1380_472# 0.002164f
C6968 FILLER_0_6_239/a_124_375# net37 0.001989f
C6969 _428_/a_1000_472# _043_ 0.020031f
C6970 FILLER_0_22_128/a_124_375# vdd 0.013058f
C6971 trim_mask\[4\] net59 0.012971f
C6972 _144_ FILLER_0_21_133/a_124_375# 0.001885f
C6973 _322_/a_848_380# _125_ 0.013667f
C6974 net25 FILLER_0_22_86/a_124_375# 0.004298f
C6975 ctln[5] FILLER_0_0_198/a_124_375# 0.002726f
C6976 _132_ _114_ 0.08562f
C6977 net41 _178_ 0.019945f
C6978 net34 FILLER_0_22_128/a_2724_472# 0.004465f
C6979 _052_ _424_/a_1204_472# 0.002681f
C6980 _098_ _434_/a_2248_156# 0.016991f
C6981 net80 _337_/a_49_472# 0.015686f
C6982 _441_/a_1308_423# vss 0.016854f
C6983 net57 _443_/a_2248_156# 0.001117f
C6984 FILLER_0_13_212/a_484_472# mask\[0\] 0.001794f
C6985 _399_/a_224_472# _182_ 0.002729f
C6986 FILLER_0_13_206/a_124_375# vdd 0.034528f
C6987 mask\[3\] FILLER_0_18_177/a_2364_375# 0.002935f
C6988 trim_val\[2\] net17 0.019133f
C6989 _447_/a_36_151# vdd 0.067176f
C6990 trimb[0] vdd 0.10929f
C6991 net20 mask\[3\] 0.047107f
C6992 FILLER_0_15_228/a_36_472# vss 0.006585f
C6993 _187_ _408_/a_1936_472# 0.017573f
C6994 FILLER_0_11_101/a_36_472# _120_ 0.007656f
C6995 _213_/a_67_603# _098_ 0.018092f
C6996 net55 FILLER_0_17_72/a_1828_472# 0.001217f
C6997 _440_/a_2248_156# vss 0.010006f
C6998 _440_/a_2665_112# vdd -0.002297f
C6999 _110_ mask\[9\] 0.00319f
C7000 FILLER_0_19_142/a_36_472# vss 0.011026f
C7001 _439_/a_448_472# vss 0.036535f
C7002 _439_/a_1308_423# vdd 0.002368f
C7003 net81 FILLER_0_15_205/a_124_375# 0.015134f
C7004 FILLER_0_8_138/a_124_375# _313_/a_67_603# 0.00744f
C7005 vdd FILLER_0_13_290/a_36_472# 0.027484f
C7006 vss FILLER_0_13_290/a_124_375# 0.031844f
C7007 net4 _264_/a_224_472# 0.001408f
C7008 mask\[7\] _350_/a_257_69# 0.001135f
C7009 net62 _044_ 0.101165f
C7010 _095_ net14 0.043065f
C7011 _073_ _070_ 0.001892f
C7012 fanout56/a_36_113# vdd 0.078814f
C7013 _077_ _042_ 0.045685f
C7014 net81 _098_ 0.029506f
C7015 _443_/a_2560_156# _170_ 0.00758f
C7016 _443_/a_2248_156# _037_ 0.005717f
C7017 net76 FILLER_0_5_181/a_36_472# 0.014784f
C7018 _412_/a_448_472# net2 0.033994f
C7019 _035_ _445_/a_36_151# 0.002276f
C7020 FILLER_0_19_47/a_484_472# vss 0.001338f
C7021 _008_ _103_ 0.092504f
C7022 _131_ FILLER_0_17_104/a_932_472# 0.002988f
C7023 net20 _083_ 0.230786f
C7024 _426_/a_36_151# FILLER_0_8_247/a_1020_375# 0.059049f
C7025 _020_ _334_/a_36_160# 0.028435f
C7026 FILLER_0_18_2/a_36_472# vss 0.001872f
C7027 FILLER_0_6_47/a_2276_472# vss 0.004086f
C7028 FILLER_0_6_47/a_2724_472# vdd 0.002467f
C7029 net56 FILLER_0_18_139/a_572_375# 0.005919f
C7030 _175_ FILLER_0_15_72/a_36_472# 0.006746f
C7031 FILLER_0_4_144/a_484_472# net23 0.01239f
C7032 trim[1] vdd 0.089624f
C7033 _428_/a_36_151# FILLER_0_14_107/a_572_375# 0.001597f
C7034 _155_ _029_ 0.174512f
C7035 cal net2 0.081236f
C7036 net57 _170_ 0.057355f
C7037 en vdd 0.282941f
C7038 _425_/a_36_151# _014_ 0.12681f
C7039 FILLER_0_10_78/a_932_472# vdd 0.005517f
C7040 _139_ mask\[1\] 0.017315f
C7041 mask\[5\] FILLER_0_19_171/a_124_375# 0.002206f
C7042 _118_ _311_/a_3220_473# 0.001133f
C7043 FILLER_0_21_142/a_36_472# net54 0.02217f
C7044 _063_ FILLER_0_6_47/a_36_472# 0.007244f
C7045 mask\[9\] FILLER_0_20_107/a_36_472# 0.006047f
C7046 _291_/a_36_160# vss 0.012222f
C7047 _150_ _027_ 0.006689f
C7048 _418_/a_796_472# _007_ 0.012286f
C7049 _311_/a_66_473# vdd 0.106886f
C7050 _398_/a_36_113# _178_ 0.004282f
C7051 net3 _095_ 0.002383f
C7052 _111_ _303_/a_244_68# 0.001153f
C7053 FILLER_0_9_223/a_572_375# _055_ 0.022619f
C7054 _207_/a_67_603# vss 0.00837f
C7055 net15 _120_ 0.028275f
C7056 FILLER_0_11_101/a_572_375# FILLER_0_9_105/a_36_472# 0.0027f
C7057 _091_ FILLER_0_19_171/a_484_472# 0.013944f
C7058 _367_/a_36_68# vss 0.001589f
C7059 FILLER_0_22_86/a_932_472# net14 0.020589f
C7060 _056_ _062_ 0.320621f
C7061 FILLER_0_7_72/a_1380_472# _077_ 0.001315f
C7062 _072_ _085_ 0.408915f
C7063 net76 cal_itt\[1\] 0.027781f
C7064 net34 _208_/a_36_160# 0.002666f
C7065 output46/a_224_472# FILLER_0_20_2/a_572_375# 0.03228f
C7066 _448_/a_2248_156# net59 0.005684f
C7067 FILLER_0_24_274/a_484_472# _420_/a_36_151# 0.002841f
C7068 _176_ FILLER_0_15_59/a_124_375# 0.007169f
C7069 _170_ _037_ 0.05171f
C7070 _427_/a_796_472# vss 0.001131f
C7071 _077_ FILLER_0_9_72/a_572_375# 0.008103f
C7072 net68 FILLER_0_8_37/a_484_472# 0.002696f
C7073 _136_ _067_ 0.051914f
C7074 _141_ _340_/a_36_160# 0.00584f
C7075 FILLER_0_8_138/a_124_375# _058_ 0.009863f
C7076 FILLER_0_7_162/a_36_472# FILLER_0_8_156/a_572_375# 0.001543f
C7077 _432_/a_2665_112# _019_ 0.002852f
C7078 _331_/a_448_472# _134_ 0.001126f
C7079 FILLER_0_11_78/a_484_472# _389_/a_36_148# 0.001043f
C7080 FILLER_0_19_47/a_572_375# net55 0.003447f
C7081 fanout72/a_36_113# _394_/a_56_524# 0.002775f
C7082 mask\[4\] _202_/a_36_160# 0.007912f
C7083 _020_ net36 0.001995f
C7084 _448_/a_36_151# FILLER_0_2_177/a_572_375# 0.001597f
C7085 _136_ FILLER_0_14_99/a_124_375# 0.007209f
C7086 net22 _202_/a_36_160# 0.052766f
C7087 net47 FILLER_0_5_164/a_124_375# 0.011983f
C7088 _077_ cal_count\[3\] 0.176576f
C7089 vss FILLER_0_8_156/a_484_472# 0.004078f
C7090 net76 vss 0.436111f
C7091 net44 _450_/a_1040_527# 0.002267f
C7092 FILLER_0_7_162/a_124_375# _074_ 0.007213f
C7093 FILLER_0_7_195/a_36_472# cal_itt\[3\] 0.070665f
C7094 mask\[4\] FILLER_0_18_139/a_1468_375# 0.023004f
C7095 _128_ FILLER_0_12_236/a_36_472# 0.001043f
C7096 net7 _446_/a_2248_156# 0.001166f
C7097 _070_ _067_ 0.001869f
C7098 _449_/a_796_472# _067_ 0.004874f
C7099 FILLER_0_12_220/a_932_472# _223_/a_36_160# 0.001323f
C7100 _114_ state\[1\] 0.087216f
C7101 FILLER_0_13_212/a_124_375# vdd 0.010978f
C7102 net52 FILLER_0_2_127/a_36_472# 0.001964f
C7103 mask\[3\] _289_/a_36_472# 0.02347f
C7104 _033_ _444_/a_1204_472# 0.002294f
C7105 _110_ net35 0.053239f
C7106 _436_/a_36_151# vdd 0.078019f
C7107 net27 FILLER_0_15_235/a_572_375# 0.001554f
C7108 _053_ FILLER_0_7_72/a_1828_472# 0.013271f
C7109 _068_ _311_/a_3220_473# 0.004371f
C7110 _430_/a_796_472# net63 0.002914f
C7111 _149_ _026_ 0.243704f
C7112 _235_/a_255_603# trim_mask\[2\] 0.001488f
C7113 _235_/a_67_603# trim_val\[2\] 0.00747f
C7114 FILLER_0_11_142/a_124_375# cal_count\[3\] 0.010782f
C7115 output47/a_224_472# FILLER_0_15_2/a_36_472# 0.035046f
C7116 _108_ vss 0.160825f
C7117 _370_/a_692_472# _152_ 0.005908f
C7118 _370_/a_1152_472# _081_ 0.001901f
C7119 _125_ _124_ 0.085897f
C7120 _409_/a_245_68# cal_count\[3\] 0.001164f
C7121 _133_ _120_ 0.003762f
C7122 _413_/a_448_472# net82 0.004927f
C7123 _054_ _220_/a_67_603# 0.004333f
C7124 cal_count\[3\] _373_/a_1060_68# 0.00165f
C7125 output35/a_224_472# _048_ 0.009509f
C7126 net60 _418_/a_1308_423# 0.016365f
C7127 _173_ vss 0.063821f
C7128 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_124_375# 0.003228f
C7129 net34 _210_/a_67_603# 0.01049f
C7130 _093_ net71 0.133323f
C7131 _445_/a_2248_156# net47 0.028909f
C7132 net60 _419_/a_2665_112# 0.059916f
C7133 net58 FILLER_0_9_290/a_36_472# 0.005553f
C7134 _095_ _098_ 0.057687f
C7135 _343_/a_49_472# _143_ 0.00918f
C7136 FILLER_0_7_72/a_2724_472# FILLER_0_6_90/a_572_375# 0.001684f
C7137 fanout80/a_36_113# _136_ 0.006151f
C7138 _104_ _107_ 0.021508f
C7139 ctln[6] output14/a_224_472# 0.007421f
C7140 _431_/a_1000_472# _137_ 0.010168f
C7141 fanout80/a_36_113# net21 0.021603f
C7142 mask\[8\] net14 0.040566f
C7143 net57 _267_/a_36_472# 0.032037f
C7144 FILLER_0_19_47/a_36_472# _424_/a_1308_423# 0.010224f
C7145 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_572_375# 0.086635f
C7146 FILLER_0_20_193/a_572_375# net21 0.002103f
C7147 FILLER_0_7_59/a_36_472# vdd 0.016778f
C7148 FILLER_0_7_59/a_572_375# vss 0.017487f
C7149 _147_ _146_ 0.001164f
C7150 FILLER_0_8_107/a_36_472# _058_ 0.015262f
C7151 net54 FILLER_0_22_86/a_1020_375# 0.001597f
C7152 _053_ FILLER_0_5_212/a_124_375# 0.048501f
C7153 FILLER_0_8_239/a_36_472# _317_/a_36_113# 0.00191f
C7154 net35 FILLER_0_22_128/a_2812_375# 0.010399f
C7155 FILLER_0_1_204/a_36_472# vdd 0.009339f
C7156 FILLER_0_1_204/a_124_375# vss 0.018397f
C7157 _328_/a_36_113# net14 0.002272f
C7158 net20 FILLER_0_6_231/a_484_472# 0.017025f
C7159 net68 FILLER_0_6_47/a_572_375# 0.007672f
C7160 _075_ _414_/a_448_472# 0.020304f
C7161 FILLER_0_9_223/a_484_472# vdd 0.004285f
C7162 output46/a_224_472# FILLER_0_21_28/a_124_375# 0.003337f
C7163 _092_ FILLER_0_17_218/a_572_375# 0.006125f
C7164 _103_ _006_ 0.00205f
C7165 _178_ cal_count\[2\] 0.119443f
C7166 _104_ FILLER_0_23_274/a_124_375# 0.002159f
C7167 _136_ FILLER_0_16_154/a_572_375# 0.003842f
C7168 trim_mask\[1\] FILLER_0_6_47/a_1468_375# 0.007169f
C7169 output15/a_224_472# trim_mask\[3\] 0.024718f
C7170 _435_/a_2248_156# mask\[6\] 0.001778f
C7171 net53 FILLER_0_14_99/a_36_472# 0.004153f
C7172 _086_ FILLER_0_7_104/a_572_375# 0.003137f
C7173 _114_ FILLER_0_12_136/a_36_472# 0.003953f
C7174 _080_ vdd 0.123811f
C7175 _070_ FILLER_0_9_105/a_36_472# 0.023853f
C7176 _274_/a_2552_68# vss 0.003123f
C7177 _333_/a_36_160# mask\[2\] 0.022517f
C7178 FILLER_0_14_123/a_124_375# FILLER_0_14_107/a_1468_375# 0.012001f
C7179 _444_/a_36_151# vss 0.003795f
C7180 _444_/a_448_472# vdd 0.03285f
C7181 FILLER_0_22_86/a_932_472# _098_ 0.001442f
C7182 _093_ _013_ 0.064462f
C7183 FILLER_0_7_72/a_124_375# FILLER_0_7_59/a_572_375# 0.003228f
C7184 net74 net14 0.034568f
C7185 trim_mask\[2\] _367_/a_36_68# 0.001302f
C7186 _444_/a_1000_472# net17 0.02064f
C7187 net54 _437_/a_2248_156# 0.046559f
C7188 _027_ _438_/a_448_472# 0.053901f
C7189 _066_ _169_ 0.222791f
C7190 net36 net19 0.031858f
C7191 _427_/a_448_472# net23 0.014853f
C7192 FILLER_0_8_138/a_36_472# vss 0.008189f
C7193 _065_ _064_ 0.007356f
C7194 FILLER_0_4_99/a_124_375# vdd 0.029154f
C7195 net25 FILLER_0_23_88/a_124_375# 0.010782f
C7196 output34/a_224_472# _277_/a_36_160# 0.014508f
C7197 fanout62/a_36_160# net79 0.011515f
C7198 _065_ _447_/a_1204_472# 0.017675f
C7199 _070_ _121_ 0.285424f
C7200 trim[0] net40 0.005988f
C7201 _083_ cal_itt\[1\] 0.046464f
C7202 result[5] net78 0.020038f
C7203 output13/a_224_472# _170_ 0.024999f
C7204 _415_/a_36_151# net79 0.001156f
C7205 mask\[3\] vss 0.664467f
C7206 FILLER_0_6_239/a_124_375# _122_ 0.01772f
C7207 FILLER_0_9_28/a_1380_472# net16 0.005297f
C7208 FILLER_0_2_93/a_124_375# _030_ 0.001641f
C7209 FILLER_0_8_2/a_124_375# net40 0.002839f
C7210 _414_/a_36_151# _163_ 0.001186f
C7211 _386_/a_1152_472# _163_ 0.004076f
C7212 FILLER_0_12_50/a_36_472# _067_ 0.011087f
C7213 _417_/a_1308_423# output30/a_224_472# 0.001434f
C7214 net82 net74 0.007059f
C7215 _116_ _162_ 0.00156f
C7216 FILLER_0_21_125/a_484_472# net54 0.022347f
C7217 net41 _450_/a_2225_156# 0.024042f
C7218 FILLER_0_11_78/a_36_472# _120_ 0.014169f
C7219 FILLER_0_9_72/a_484_472# vss 0.008087f
C7220 FILLER_0_9_72/a_932_472# vdd 0.00604f
C7221 _131_ _330_/a_224_472# 0.001186f
C7222 net27 _426_/a_1000_472# 0.002971f
C7223 mask\[1\] FILLER_0_15_205/a_124_375# 0.007883f
C7224 _169_ net37 0.03934f
C7225 net64 _098_ 0.281888f
C7226 _272_/a_36_472# _003_ 0.001634f
C7227 _129_ _118_ 0.213736f
C7228 _436_/a_448_472# FILLER_0_22_128/a_124_375# 0.006782f
C7229 net65 net37 0.008382f
C7230 _066_ net59 0.002935f
C7231 net55 FILLER_0_13_72/a_484_472# 0.004375f
C7232 net35 _049_ 0.022439f
C7233 _083_ vss 0.0284f
C7234 net48 _251_/a_244_472# 0.001259f
C7235 _144_ vdd 0.40911f
C7236 _094_ _418_/a_36_151# 0.041823f
C7237 FILLER_0_16_57/a_1380_472# net55 0.002219f
C7238 _098_ mask\[1\] 1.476748f
C7239 _069_ mask\[0\] 0.040599f
C7240 FILLER_0_1_192/a_36_472# net59 0.082738f
C7241 output8/a_224_472# FILLER_0_3_221/a_484_472# 0.001699f
C7242 _390_/a_692_472# _136_ 0.004782f
C7243 net44 FILLER_0_20_2/a_572_375# 0.002597f
C7244 _073_ net9 0.005417f
C7245 _028_ FILLER_0_7_72/a_1828_472# 0.001777f
C7246 FILLER_0_6_90/a_484_472# FILLER_0_4_91/a_572_375# 0.00108f
C7247 net57 FILLER_0_13_142/a_484_472# 0.011685f
C7248 _320_/a_1792_472# _043_ 0.002235f
C7249 net18 _417_/a_2248_156# 0.001601f
C7250 FILLER_0_20_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001543f
C7251 FILLER_0_15_282/a_484_472# output30/a_224_472# 0.001711f
C7252 FILLER_0_15_282/a_124_375# net30 0.00123f
C7253 net62 _416_/a_1308_423# 0.002665f
C7254 vss _416_/a_1000_472# 0.001784f
C7255 ctlp[6] output23/a_224_472# 0.024575f
C7256 FILLER_0_16_89/a_124_375# FILLER_0_17_72/a_1916_375# 0.026339f
C7257 mask\[2\] FILLER_0_16_154/a_36_472# 0.312123f
C7258 FILLER_0_13_142/a_1468_375# _043_ 0.009636f
C7259 FILLER_0_14_91/a_36_472# _176_ 0.076419f
C7260 mask\[8\] _098_ 0.096999f
C7261 output14/a_224_472# ctln[7] 0.076006f
C7262 result[0] net18 0.085445f
C7263 _085_ state\[1\] 0.182697f
C7264 mask\[5\] net21 0.212814f
C7265 net37 net59 0.03883f
C7266 _086_ FILLER_0_11_124/a_36_472# 0.010729f
C7267 _095_ _405_/a_67_603# 0.012596f
C7268 net62 _283_/a_36_472# 0.002309f
C7269 result[4] net19 0.015095f
C7270 net76 net4 0.024291f
C7271 _323_/a_36_113# vdd 0.009958f
C7272 _111_ net36 0.102444f
C7273 FILLER_0_18_76/a_572_375# net71 0.006025f
C7274 _430_/a_36_151# FILLER_0_18_209/a_36_472# 0.002841f
C7275 _131_ _095_ 0.043211f
C7276 _432_/a_36_151# _143_ 0.001486f
C7277 FILLER_0_18_2/a_1380_472# net38 0.029747f
C7278 FILLER_0_16_107/a_124_375# _040_ 0.008721f
C7279 mask\[7\] _108_ 0.785154f
C7280 net57 _113_ 0.012056f
C7281 ctlp[1] FILLER_0_24_274/a_1468_375# 0.01305f
C7282 FILLER_0_21_28/a_2724_472# vss -0.001553f
C7283 net36 _280_/a_224_472# 0.001012f
C7284 FILLER_0_6_90/a_36_472# vdd 0.00366f
C7285 FILLER_0_6_90/a_572_375# vss 0.006421f
C7286 FILLER_0_16_73/a_36_472# _131_ 0.008223f
C7287 net35 _436_/a_2248_156# 0.014499f
C7288 output31/a_224_472# FILLER_0_16_255/a_124_375# 0.001274f
C7289 _428_/a_36_151# vdd 0.131612f
C7290 _415_/a_1204_472# _004_ 0.002391f
C7291 trim_mask\[4\] _370_/a_848_380# 0.027744f
C7292 net15 FILLER_0_5_54/a_932_472# 0.008904f
C7293 net52 FILLER_0_2_111/a_484_472# 0.061249f
C7294 valid net1 0.00347f
C7295 cal_itt\[2\] FILLER_0_3_221/a_932_472# 0.016327f
C7296 FILLER_0_14_99/a_36_472# FILLER_0_14_107/a_36_472# 0.002296f
C7297 _411_/a_2248_156# vdd 0.006283f
C7298 _372_/a_2590_472# _076_ 0.002268f
C7299 _129_ _068_ 0.104827f
C7300 FILLER_0_11_282/a_36_472# vss 0.007114f
C7301 net55 _182_ 0.012838f
C7302 FILLER_0_16_89/a_124_375# net53 0.001032f
C7303 FILLER_0_12_220/a_124_375# _070_ 0.007554f
C7304 FILLER_0_4_107/a_484_472# _157_ 0.027364f
C7305 _114_ vdd 1.30767f
C7306 _163_ FILLER_0_5_148/a_36_472# 0.002454f
C7307 en_co_clk cal_count\[3\] 0.001359f
C7308 _414_/a_36_151# FILLER_0_7_195/a_124_375# 0.059049f
C7309 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_36_472# 0.086742f
C7310 fanout50/a_36_160# vdd 0.009536f
C7311 _057_ _061_ 0.030546f
C7312 FILLER_0_17_72/a_484_472# _131_ 0.002672f
C7313 trim_mask\[0\] FILLER_0_10_94/a_484_472# 0.015575f
C7314 _412_/a_36_151# valid 0.009757f
C7315 vdd FILLER_0_14_235/a_484_472# 0.010228f
C7316 vss FILLER_0_14_235/a_36_472# 0.001602f
C7317 _425_/a_1308_423# net19 0.058462f
C7318 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_36_472# 0.002296f
C7319 net62 FILLER_0_14_235/a_124_375# 0.015659f
C7320 net81 FILLER_0_15_212/a_932_472# 0.003953f
C7321 _443_/a_36_151# vdd 0.175472f
C7322 _142_ _132_ 0.006253f
C7323 output47/a_224_472# _398_/a_36_113# 0.001605f
C7324 FILLER_0_24_130/a_36_472# net54 0.06125f
C7325 FILLER_0_4_197/a_36_472# _270_/a_36_472# 0.004546f
C7326 output48/a_224_472# _082_ 0.002393f
C7327 output37/a_224_472# net18 0.046654f
C7328 FILLER_0_10_78/a_36_472# net52 0.014225f
C7329 _414_/a_1308_423# _053_ 0.029387f
C7330 _430_/a_2560_156# mask\[2\] 0.010268f
C7331 _428_/a_2665_112# _095_ 0.001471f
C7332 _445_/a_2665_112# trim_val\[1\] 0.015206f
C7333 net57 _118_ 0.036179f
C7334 _072_ FILLER_0_12_220/a_36_472# 0.01861f
C7335 _088_ FILLER_0_3_212/a_124_375# 0.0042f
C7336 net79 FILLER_0_13_290/a_124_375# 0.043673f
C7337 net68 FILLER_0_3_54/a_124_375# 0.022559f
C7338 _026_ net14 0.010792f
C7339 _147_ _435_/a_448_472# 0.001008f
C7340 _093_ FILLER_0_19_155/a_36_472# 0.001737f
C7341 _116_ _373_/a_244_68# 0.001213f
C7342 _132_ FILLER_0_18_107/a_2812_375# 0.002706f
C7343 net39 _444_/a_1000_472# 0.001323f
C7344 _432_/a_2560_156# vdd 0.003219f
C7345 FILLER_0_2_177/a_124_375# vdd 0.019296f
C7346 net75 _411_/a_2248_156# 0.032114f
C7347 _096_ _116_ 0.020685f
C7348 _103_ _007_ 0.002514f
C7349 net15 _043_ 0.042278f
C7350 FILLER_0_12_2/a_484_472# net44 0.046864f
C7351 _058_ FILLER_0_8_156/a_36_472# 0.011885f
C7352 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001597f
C7353 FILLER_0_17_218/a_572_375# vdd 0.019414f
C7354 FILLER_0_17_218/a_124_375# vss 0.012673f
C7355 net71 FILLER_0_22_107/a_124_375# 0.018295f
C7356 _412_/a_36_151# net9 0.005212f
C7357 _435_/a_2560_156# vdd 0.001372f
C7358 _435_/a_2665_112# vss 0.002665f
C7359 FILLER_0_10_78/a_484_472# _077_ 0.002486f
C7360 output18/a_224_472# ctlp[1] 0.039734f
C7361 FILLER_0_18_61/a_124_375# FILLER_0_18_53/a_572_375# 0.012001f
C7362 FILLER_0_9_72/a_1468_375# _439_/a_2248_156# 0.001901f
C7363 FILLER_0_8_263/a_124_375# vss 0.007944f
C7364 FILLER_0_8_263/a_36_472# vdd 0.092694f
C7365 vss FILLER_0_6_231/a_484_472# 0.005629f
C7366 FILLER_0_20_31/a_36_472# vdd 0.097195f
C7367 FILLER_0_20_31/a_124_375# vss 0.049142f
C7368 _093_ _110_ 0.08348f
C7369 net56 _137_ 0.0313f
C7370 trimb[0] output46/a_224_472# 0.048191f
C7371 net20 _421_/a_448_472# 0.015767f
C7372 FILLER_0_21_286/a_124_375# vdd 0.026138f
C7373 FILLER_0_4_197/a_1380_472# net22 0.012286f
C7374 net76 FILLER_0_5_198/a_124_375# 0.006974f
C7375 FILLER_0_20_87/a_36_472# vss 0.006244f
C7376 _406_/a_36_159# net17 0.053547f
C7377 net70 FILLER_0_13_100/a_36_472# 0.00585f
C7378 _421_/a_36_151# net19 0.016842f
C7379 _132_ _354_/a_49_472# 0.034372f
C7380 result[4] fanout78/a_36_113# 0.001531f
C7381 _451_/a_2225_156# _040_ 0.015815f
C7382 cal_itt\[3\] _375_/a_1612_497# 0.003901f
C7383 net16 _408_/a_728_93# 0.107634f
C7384 result[7] FILLER_0_24_274/a_124_375# 0.006125f
C7385 FILLER_0_20_193/a_484_472# _205_/a_36_160# 0.001684f
C7386 _440_/a_1308_423# _160_ 0.002554f
C7387 _211_/a_36_160# net14 0.005761f
C7388 net15 _175_ 0.052586f
C7389 _394_/a_718_524# vss 0.002666f
C7390 FILLER_0_7_195/a_36_472# _161_ 0.015074f
C7391 net58 _004_ 0.00116f
C7392 output48/a_224_472# _112_ 0.027383f
C7393 _036_ _168_ 0.01699f
C7394 FILLER_0_2_93/a_124_375# trim_mask\[3\] 0.003033f
C7395 FILLER_0_19_28/a_484_472# vss 0.001207f
C7396 FILLER_0_16_57/a_484_472# FILLER_0_17_56/a_572_375# 0.001723f
C7397 _050_ net23 0.003752f
C7398 net57 _068_ 0.029812f
C7399 _186_ _043_ 0.045082f
C7400 mask\[4\] FILLER_0_20_177/a_36_472# 0.001215f
C7401 _077_ _120_ 0.205715f
C7402 output8/a_224_472# output11/a_224_472# 0.003437f
C7403 FILLER_0_21_28/a_3172_472# _424_/a_36_151# 0.001723f
C7404 FILLER_0_10_28/a_36_472# net17 0.012954f
C7405 mask\[5\] _021_ 0.001088f
C7406 _174_ _180_ 0.102241f
C7407 net4 _083_ 0.135165f
C7408 _073_ _084_ 0.048469f
C7409 net64 FILLER_0_9_270/a_484_472# 0.017924f
C7410 _186_ _185_ 0.007962f
C7411 trim[0] trim[3] 0.012429f
C7412 net34 FILLER_0_22_177/a_572_375# 0.006974f
C7413 _195_/a_67_603# _045_ 0.004028f
C7414 net82 FILLER_0_3_172/a_3172_472# 0.007677f
C7415 _139_ _019_ 0.094494f
C7416 net75 FILLER_0_8_263/a_36_472# 0.020293f
C7417 _150_ mask\[9\] 0.162185f
C7418 net80 _434_/a_36_151# 0.067037f
C7419 _041_ vss 0.012963f
C7420 FILLER_0_5_128/a_124_375# _370_/a_124_24# 0.023285f
C7421 ctlp[4] net21 0.04068f
C7422 FILLER_0_18_2/a_1380_472# net55 0.007469f
C7423 net48 _317_/a_36_113# 0.018494f
C7424 FILLER_0_11_142/a_124_375# _120_ 0.036088f
C7425 FILLER_0_15_116/a_572_375# _095_ 0.00152f
C7426 net60 net78 0.030634f
C7427 net52 _441_/a_448_472# 0.04874f
C7428 net72 FILLER_0_20_31/a_36_472# 0.002751f
C7429 output47/a_224_472# cal_count\[2\] 0.080405f
C7430 FILLER_0_24_96/a_124_375# net35 0.001886f
C7431 fanout63/a_36_160# FILLER_0_15_228/a_36_472# 0.014197f
C7432 FILLER_0_5_109/a_484_472# vss 0.00212f
C7433 _115_ _439_/a_2665_112# 0.003617f
C7434 comp vdd 0.108153f
C7435 _238_/a_67_603# net52 0.006325f
C7436 result[7] FILLER_0_23_274/a_124_375# 0.017938f
C7437 net52 _440_/a_1204_472# 0.003916f
C7438 _176_ _134_ 0.035146f
C7439 _061_ cal_count\[3\] 0.003415f
C7440 net74 _372_/a_170_472# 0.079123f
C7441 _187_ vdd 0.194575f
C7442 _131_ net74 0.227843f
C7443 net52 _439_/a_36_151# 0.01388f
C7444 _122_ _169_ 0.014463f
C7445 calibrate _163_ 0.026892f
C7446 _414_/a_448_472# _003_ 0.023209f
C7447 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_36_472# 0.002296f
C7448 mask\[4\] FILLER_0_19_171/a_932_472# 0.004669f
C7449 net41 net38 0.059214f
C7450 _050_ _025_ 0.033887f
C7451 _085_ vdd 0.227153f
C7452 _106_ FILLER_0_17_218/a_36_472# 0.002777f
C7453 FILLER_0_5_164/a_124_375# vdd 0.00419f
C7454 _026_ _098_ 0.197713f
C7455 net55 FILLER_0_19_28/a_572_375# 0.002115f
C7456 _010_ _420_/a_36_151# 0.001838f
C7457 _421_/a_36_151# _009_ 0.00246f
C7458 _414_/a_448_472# net21 0.040301f
C7459 result[5] net60 0.16275f
C7460 FILLER_0_5_212/a_124_375# _081_ 0.01149f
C7461 FILLER_0_18_107/a_2276_472# _137_ 0.001752f
C7462 state\[0\] _274_/a_1164_497# 0.002914f
C7463 _098_ FILLER_0_21_206/a_124_375# 0.001882f
C7464 _104_ net32 0.342568f
C7465 _131_ cal_count\[1\] 0.001497f
C7466 net69 FILLER_0_2_111/a_572_375# 0.015789f
C7467 state\[2\] _043_ 0.028842f
C7468 FILLER_0_22_128/a_3172_472# vdd 0.003395f
C7469 FILLER_0_22_128/a_2724_472# vss 0.005195f
C7470 _108_ _295_/a_36_472# 0.014558f
C7471 _098_ _097_ 0.034041f
C7472 net32 _421_/a_2665_112# 0.019532f
C7473 net38 FILLER_0_20_15/a_36_472# 0.070475f
C7474 _018_ vdd 0.048119f
C7475 FILLER_0_5_109/a_124_375# _153_ 0.040726f
C7476 _163_ _153_ 0.243815f
C7477 FILLER_0_8_107/a_124_375# FILLER_0_9_105/a_484_472# 0.001684f
C7478 _133_ FILLER_0_10_107/a_484_472# 0.001798f
C7479 net18 _044_ 0.174456f
C7480 net49 vss 0.689397f
C7481 _251_/a_468_472# vss 0.001679f
C7482 _442_/a_2665_112# vdd 0.056153f
C7483 _452_/a_836_156# _041_ 0.001052f
C7484 _053_ FILLER_0_6_47/a_2276_472# 0.004472f
C7485 _096_ _225_/a_36_160# 0.004807f
C7486 net68 vss 0.635359f
C7487 FILLER_0_14_50/a_36_472# _181_ 0.001514f
C7488 _093_ fanout54/a_36_160# 0.003506f
C7489 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_572_375# 0.001597f
C7490 _144_ _433_/a_36_151# 0.086558f
C7491 _122_ net59 0.041453f
C7492 net32 result[6] 0.048987f
C7493 net29 FILLER_0_16_255/a_36_472# 0.086886f
C7494 _445_/a_2248_156# vdd 0.018573f
C7495 _440_/a_2665_112# FILLER_0_5_88/a_124_375# 0.02132f
C7496 FILLER_0_14_91/a_124_375# _136_ 0.013064f
C7497 net24 _436_/a_36_151# 0.075327f
C7498 _424_/a_2665_112# FILLER_0_21_60/a_572_375# 0.001077f
C7499 _136_ _138_ 0.186242f
C7500 _428_/a_2665_112# net74 0.048822f
C7501 _048_ FILLER_0_18_209/a_124_375# 0.001615f
C7502 _065_ net50 0.123581f
C7503 output14/a_224_472# net52 0.02346f
C7504 cal_itt\[2\] _084_ 0.061303f
C7505 _077_ _227_/a_36_160# 0.012587f
C7506 mask\[5\] FILLER_0_18_177/a_36_472# 0.001063f
C7507 _138_ net21 0.003242f
C7508 _282_/a_36_160# mask\[2\] 0.023533f
C7509 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_36_472# 0.086742f
C7510 _104_ _422_/a_2248_156# 0.041703f
C7511 net55 FILLER_0_18_76/a_484_472# 0.003745f
C7512 _322_/a_124_24# _118_ 0.04952f
C7513 net1 _084_ 0.008356f
C7514 net16 FILLER_0_17_38/a_124_375# 0.046435f
C7515 FILLER_0_16_241/a_124_375# _198_/a_67_603# 0.002082f
C7516 net55 _423_/a_2665_112# 0.002379f
C7517 _425_/a_1000_472# vdd 0.019072f
C7518 state\[0\] FILLER_0_12_220/a_932_472# 0.001003f
C7519 mask\[9\] _012_ 0.008145f
C7520 net20 FILLER_0_12_220/a_1468_375# 0.016974f
C7521 mask\[0\] net22 0.054097f
C7522 FILLER_0_9_282/a_484_472# vss 0.00561f
C7523 net38 _398_/a_36_113# 0.061273f
C7524 _074_ net22 0.079421f
C7525 mask\[7\] _435_/a_2665_112# 0.030393f
C7526 net70 FILLER_0_14_107/a_1020_375# 0.011157f
C7527 FILLER_0_7_72/a_484_472# vss 0.003793f
C7528 net32 net22 0.042885f
C7529 _130_ cal_count\[3\] 0.037708f
C7530 FILLER_0_15_212/a_932_472# mask\[1\] 0.014799f
C7531 _248_/a_36_68# _060_ 0.004581f
C7532 _070_ FILLER_0_10_94/a_36_472# 0.001866f
C7533 _274_/a_2124_68# net4 0.00137f
C7534 _050_ _436_/a_1000_472# 0.02064f
C7535 _159_ _081_ 0.003646f
C7536 net31 net60 0.012623f
C7537 FILLER_0_16_57/a_36_472# _131_ 0.00864f
C7538 _328_/a_36_113# _126_ 0.023932f
C7539 fanout73/a_36_113# net70 0.00238f
C7540 net81 _060_ 0.019654f
C7541 _420_/a_36_151# vdd 0.137919f
C7542 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_484_472# 0.013277f
C7543 _291_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C7544 FILLER_0_7_195/a_124_375# calibrate 0.00576f
C7545 fanout65/a_36_113# vdd 0.10473f
C7546 _333_/a_36_160# vss 0.030799f
C7547 _189_/a_67_603# FILLER_0_13_228/a_36_472# 0.005759f
C7548 _320_/a_224_472# vdd 0.001757f
C7549 trimb[0] net44 0.00246f
C7550 mask\[3\] _141_ 0.361692f
C7551 _098_ FILLER_0_15_180/a_124_375# 0.019007f
C7552 _208_/a_36_160# vss 0.012188f
C7553 net20 _419_/a_36_151# 0.001225f
C7554 _415_/a_1000_472# result[1] 0.005365f
C7555 FILLER_0_18_2/a_3260_375# net55 0.004262f
C7556 _053_ net76 0.022571f
C7557 FILLER_0_20_15/a_1380_472# vdd 0.007068f
C7558 net41 _233_/a_36_160# 0.053625f
C7559 mask\[9\] _438_/a_448_472# 0.046823f
C7560 _093_ FILLER_0_18_139/a_124_375# 0.008393f
C7561 net16 FILLER_0_6_37/a_36_472# 0.013074f
C7562 _115_ _125_ 0.049021f
C7563 FILLER_0_3_172/a_1020_375# net22 0.013048f
C7564 _126_ net74 1.001749f
C7565 FILLER_0_9_28/a_484_472# net51 0.001023f
C7566 FILLER_0_18_171/a_36_472# _143_ 0.005167f
C7567 FILLER_0_17_72/a_1380_472# _438_/a_36_151# 0.001221f
C7568 FILLER_0_17_200/a_572_375# vdd 0.006861f
C7569 net75 _425_/a_1000_472# 0.038919f
C7570 FILLER_0_15_142/a_124_375# net36 0.006533f
C7571 net79 _416_/a_1000_472# 0.024811f
C7572 _322_/a_848_380# _076_ 0.006699f
C7573 FILLER_0_8_247/a_1468_375# vdd 0.011086f
C7574 FILLER_0_18_2/a_2276_472# net47 0.001369f
C7575 net76 FILLER_0_2_177/a_36_472# 0.003526f
C7576 FILLER_0_14_91/a_572_375# net53 0.063988f
C7577 _421_/a_448_472# vss -0.001027f
C7578 _421_/a_1308_423# vdd 0.021664f
C7579 _132_ FILLER_0_14_107/a_1020_375# 0.029702f
C7580 net23 FILLER_0_22_128/a_1828_472# 0.003857f
C7581 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1380_472# 0.013276f
C7582 result[9] _094_ 0.03984f
C7583 _028_ _439_/a_448_472# 0.017606f
C7584 _239_/a_36_160# _447_/a_36_151# 0.137659f
C7585 FILLER_0_14_107/a_932_472# _043_ 0.0017f
C7586 _415_/a_448_472# FILLER_0_11_282/a_124_375# 0.008952f
C7587 _448_/a_2560_156# _037_ 0.011661f
C7588 _127_ FILLER_0_11_124/a_36_472# 0.001641f
C7589 net63 _435_/a_2248_156# 0.045342f
C7590 _426_/a_36_151# vdd 0.086652f
C7591 _427_/a_2665_112# net36 0.009904f
C7592 _029_ net14 0.042032f
C7593 net41 net55 0.033821f
C7594 _446_/a_1308_423# net40 0.038281f
C7595 _198_/a_67_603# _046_ 0.007349f
C7596 net75 _253_/a_1100_68# 0.001047f
C7597 _441_/a_2248_156# _030_ 0.003495f
C7598 _310_/a_49_472# vdd 0.043164f
C7599 trim_mask\[2\] net49 0.041781f
C7600 _064_ net66 0.304028f
C7601 _053_ FILLER_0_7_59/a_572_375# 0.014569f
C7602 net56 _095_ 0.004847f
C7603 _095_ FILLER_0_13_142/a_932_472# 0.001782f
C7604 _074_ _076_ 0.03553f
C7605 _210_/a_67_603# vss 0.038142f
C7606 _019_ _098_ 0.010193f
C7607 _137_ mask\[1\] 0.782055f
C7608 _028_ FILLER_0_6_47/a_2276_472# 0.002066f
C7609 en_co_clk _120_ 0.008507f
C7610 trim_mask\[2\] net68 0.099597f
C7611 _116_ _055_ 0.72331f
C7612 _287_/a_36_472# net30 0.005402f
C7613 _257_/a_36_472# _075_ 0.005709f
C7614 _292_/a_36_160# _048_ 0.008475f
C7615 mask\[5\] FILLER_0_19_187/a_484_472# 0.007596f
C7616 FILLER_0_3_142/a_124_375# _443_/a_36_151# 0.059049f
C7617 FILLER_0_15_235/a_124_375# FILLER_0_15_228/a_124_375# 0.002868f
C7618 net66 output41/a_224_472# 0.015427f
C7619 _064_ _445_/a_1308_423# 0.01485f
C7620 _447_/a_1308_423# net68 0.006686f
C7621 _447_/a_36_151# _036_ 0.007244f
C7622 _187_ cal_count\[0\] 0.645851f
C7623 net79 FILLER_0_11_282/a_36_472# 0.004358f
C7624 FILLER_0_1_98/a_124_375# ctln[7] 0.004533f
C7625 net35 _012_ 0.007543f
C7626 FILLER_0_16_154/a_484_472# vdd 0.001006f
C7627 FILLER_0_16_154/a_36_472# vss 0.005098f
C7628 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_36_472# 0.001723f
C7629 _414_/a_1308_423# cal_itt\[3\] 0.044184f
C7630 FILLER_0_8_239/a_124_375# vdd 0.035205f
C7631 output19/a_224_472# net33 0.126671f
C7632 net63 net36 0.010544f
C7633 _431_/a_36_151# FILLER_0_18_107/a_3172_472# 0.00271f
C7634 _413_/a_1308_423# net82 0.003079f
C7635 _098_ _145_ 0.007514f
C7636 FILLER_0_1_212/a_124_375# FILLER_0_1_204/a_124_375# 0.003732f
C7637 _142_ vdd 0.090938f
C7638 FILLER_0_10_78/a_932_472# _176_ 0.0109f
C7639 mask\[7\] FILLER_0_22_128/a_2724_472# 0.001055f
C7640 net38 cal_count\[2\] 0.047195f
C7641 net75 FILLER_0_8_247/a_1468_375# 0.047331f
C7642 _414_/a_1308_423# _081_ 0.003429f
C7643 ctlp[9] net26 0.02213f
C7644 result[9] FILLER_0_24_274/a_572_375# 0.003576f
C7645 net38 FILLER_0_8_24/a_36_472# 0.015829f
C7646 result[4] fanout60/a_36_160# 0.027276f
C7647 _276_/a_36_160# _092_ 0.06772f
C7648 mask\[3\] fanout63/a_36_160# 0.002585f
C7649 FILLER_0_7_104/a_36_472# vdd 0.096343f
C7650 FILLER_0_7_104/a_1468_375# vss 0.003442f
C7651 _011_ _109_ 0.055905f
C7652 net32 _419_/a_2248_156# 0.034827f
C7653 output48/a_224_472# net48 0.001786f
C7654 FILLER_0_12_136/a_124_375# state\[2\] 0.001029f
C7655 FILLER_0_12_136/a_1020_375# net53 0.002709f
C7656 net73 FILLER_0_18_107/a_484_472# 0.0052f
C7657 net75 _426_/a_36_151# 0.070626f
C7658 _114_ FILLER_0_9_72/a_1380_472# 0.001043f
C7659 output32/a_224_472# _419_/a_448_472# 0.010723f
C7660 net26 FILLER_0_21_28/a_2364_375# 0.003691f
C7661 FILLER_0_18_107/a_2812_375# vdd 0.004212f
C7662 net40 _160_ 0.152292f
C7663 net52 FILLER_0_9_72/a_36_472# 0.014911f
C7664 net20 _282_/a_36_160# 0.016884f
C7665 _433_/a_2248_156# _145_ 0.009108f
C7666 FILLER_0_18_139/a_572_375# _145_ 0.00346f
C7667 _098_ FILLER_0_18_76/a_124_375# 0.001831f
C7668 FILLER_0_18_37/a_484_472# vdd 0.008381f
C7669 FILLER_0_18_37/a_36_472# vss 0.003026f
C7670 net34 vdd 1.161282f
C7671 net54 FILLER_0_20_107/a_124_375# 0.072539f
C7672 _091_ _093_ 0.035503f
C7673 FILLER_0_16_89/a_1468_375# vdd 0.038266f
C7674 _375_/a_36_68# _162_ 0.011065f
C7675 _375_/a_1612_497# _161_ 0.003325f
C7676 FILLER_0_8_138/a_124_375# _070_ 0.002997f
C7677 ctln[2] FILLER_0_1_266/a_36_472# 0.052489f
C7678 _030_ _154_ 0.004803f
C7679 _010_ _419_/a_448_472# 0.003295f
C7680 _377_/a_36_472# trim_val\[0\] 0.135527f
C7681 _069_ _047_ 0.001975f
C7682 _425_/a_36_151# calibrate 0.071513f
C7683 _087_ _088_ 0.001219f
C7684 _413_/a_2248_156# net82 0.009308f
C7685 net75 _265_/a_916_472# 0.001686f
C7686 _381_/a_244_68# _167_ 0.001153f
C7687 ctlp[2] _108_ 0.034027f
C7688 net73 _136_ 0.050578f
C7689 _077_ FILLER_0_7_72/a_2364_375# 0.002969f
C7690 _053_ _359_/a_1044_488# 0.001474f
C7691 FILLER_0_4_49/a_36_472# _160_ 0.00202f
C7692 _394_/a_728_93# _174_ 0.012471f
C7693 FILLER_0_4_197/a_932_472# vdd 0.003395f
C7694 _011_ _422_/a_448_472# 0.044695f
C7695 _354_/a_49_472# vdd -0.001073f
C7696 ctln[5] net22 0.072969f
C7697 _430_/a_2560_156# vss 0.002924f
C7698 mask\[3\] FILLER_0_17_218/a_484_472# 0.017442f
C7699 output48/a_224_472# net19 0.054227f
C7700 result[9] FILLER_0_23_274/a_36_472# 0.0064f
C7701 net20 FILLER_0_3_221/a_1020_375# 0.025371f
C7702 _057_ _267_/a_36_472# 0.038568f
C7703 net74 net69 0.143604f
C7704 _055_ _117_ 0.242156f
C7705 result[8] _422_/a_1000_472# 0.001104f
C7706 net10 _411_/a_448_472# 0.010544f
C7707 output33/a_224_472# vdd -0.031734f
C7708 _411_/a_1204_472# ctln[1] 0.031348f
C7709 FILLER_0_10_37/a_36_472# vss 0.003659f
C7710 _413_/a_36_151# FILLER_0_3_172/a_3260_375# 0.059049f
C7711 output22/a_224_472# _435_/a_1308_423# 0.005111f
C7712 _133_ _062_ 1.210949f
C7713 mask\[7\] _208_/a_36_160# 0.105845f
C7714 FILLER_0_22_177/a_124_375# mask\[6\] 0.002672f
C7715 _430_/a_2665_112# mask\[3\] 0.002697f
C7716 net63 _432_/a_2248_156# 0.047337f
C7717 _430_/a_796_472# net21 0.015066f
C7718 net47 _386_/a_124_24# 0.024696f
C7719 _321_/a_170_472# _129_ 0.024601f
C7720 _122_ _120_ 0.143427f
C7721 _184_ vss 0.068129f
C7722 _176_ _451_/a_3081_151# 0.001255f
C7723 _379_/a_36_472# _160_ 0.023459f
C7724 net27 net37 0.003648f
C7725 output26/a_224_472# FILLER_0_23_44/a_484_472# 0.0323f
C7726 _099_ FILLER_0_14_235/a_484_472# 0.00281f
C7727 output8/a_224_472# _411_/a_1308_423# 0.005111f
C7728 _101_ vss 0.05721f
C7729 net18 _416_/a_1308_423# 0.021956f
C7730 FILLER_0_9_28/a_1916_375# _054_ 0.005889f
C7731 _449_/a_36_151# vdd 0.09324f
C7732 FILLER_0_3_78/a_484_472# _160_ 0.004988f
C7733 _395_/a_36_488# _121_ 0.009689f
C7734 net50 _163_ 0.068547f
C7735 FILLER_0_12_220/a_36_472# vdd 0.027911f
C7736 FILLER_0_12_220/a_1468_375# vss 0.057853f
C7737 net81 net64 0.455159f
C7738 _311_/a_1212_473# _117_ 0.001673f
C7739 net55 FILLER_0_18_37/a_1020_375# 0.005661f
C7740 FILLER_0_4_107/a_484_472# _160_ 0.008194f
C7741 _028_ FILLER_0_7_59/a_572_375# 0.00133f
C7742 _426_/a_2665_112# net64 0.01548f
C7743 FILLER_0_17_72/a_572_375# vss 0.008057f
C7744 FILLER_0_17_72/a_1020_375# vdd 0.002541f
C7745 net2 input5/a_36_113# 0.007518f
C7746 input2/a_36_113# net5 0.001761f
C7747 FILLER_0_8_37/a_484_472# vdd 0.009603f
C7748 net81 mask\[1\] 2.509493f
C7749 _115_ net50 0.008628f
C7750 net47 FILLER_0_4_91/a_484_472# 0.007531f
C7751 _132_ FILLER_0_19_111/a_572_375# 0.01675f
C7752 _072_ FILLER_0_7_233/a_36_472# 0.00241f
C7753 _053_ FILLER_0_6_90/a_572_375# 0.073688f
C7754 net64 _060_ 0.05104f
C7755 net65 FILLER_0_3_212/a_124_375# 0.003807f
C7756 result[7] net32 0.103491f
C7757 FILLER_0_8_107/a_36_472# _070_ 0.001287f
C7758 mask\[8\] _213_/a_67_603# 0.039626f
C7759 FILLER_0_9_28/a_1828_472# vss 0.001663f
C7760 _092_ net20 0.001458f
C7761 FILLER_0_13_100/a_36_472# vdd 0.021826f
C7762 FILLER_0_13_100/a_124_375# vss 0.00513f
C7763 FILLER_0_16_107/a_572_375# vss 0.055104f
C7764 net38 _450_/a_1353_112# 0.02208f
C7765 _165_ FILLER_0_6_47/a_36_472# 0.077573f
C7766 _419_/a_36_151# vss -0.00139f
C7767 _419_/a_448_472# vdd 0.022174f
C7768 _256_/a_3368_68# net22 0.001285f
C7769 _072_ vss 0.439154f
C7770 ctln[5] net11 0.004569f
C7771 en_co_clk _390_/a_244_472# 0.001238f
C7772 net65 net8 0.203388f
C7773 FILLER_0_15_59/a_572_375# vss 0.018573f
C7774 FILLER_0_15_59/a_36_472# vdd 0.031071f
C7775 FILLER_0_7_72/a_2812_375# net50 0.006598f
C7776 FILLER_0_9_223/a_36_472# vdd 0.030289f
C7777 FILLER_0_18_107/a_124_375# net14 0.005202f
C7778 mask\[5\] FILLER_0_19_155/a_572_375# 0.007026f
C7779 _075_ _078_ 0.001896f
C7780 _017_ _134_ 0.017998f
C7781 fanout66/a_36_113# FILLER_0_3_54/a_124_375# 0.002853f
C7782 FILLER_0_17_72/a_2276_472# _136_ 0.055635f
C7783 net82 _370_/a_124_24# 0.001011f
C7784 _210_/a_67_603# mask\[7\] 0.039004f
C7785 output24/a_224_472# vdd 0.08781f
C7786 FILLER_0_5_88/a_124_375# FILLER_0_6_90/a_36_472# 0.001543f
C7787 FILLER_0_5_117/a_124_375# _158_ 0.001068f
C7788 output42/a_224_472# _054_ 0.013225f
C7789 _443_/a_2248_156# net59 0.002471f
C7790 net70 vss 0.175272f
C7791 _413_/a_36_151# vdd 0.130213f
C7792 _115_ _069_ 0.022355f
C7793 _104_ _105_ 0.931514f
C7794 net55 cal_count\[2\] 0.022989f
C7795 cal_count\[2\] _452_/a_3129_107# 0.008853f
C7796 _255_/a_224_552# _074_ 0.005907f
C7797 FILLER_0_15_142/a_572_375# vss 0.095176f
C7798 net15 _441_/a_36_151# 0.01821f
C7799 net59 FILLER_0_3_212/a_124_375# 0.057221f
C7800 net47 vss 0.919407f
C7801 mask\[2\] vdd 0.433058f
C7802 _093_ _150_ 0.406318f
C7803 _441_/a_2665_112# _164_ 0.021931f
C7804 net58 _074_ 0.004651f
C7805 output37/a_224_472# fanout59/a_36_160# 0.021845f
C7806 net34 _024_ 0.009705f
C7807 _193_/a_36_160# result[3] 0.002218f
C7808 net47 _365_/a_692_472# 0.002051f
C7809 _449_/a_36_151# net72 0.039436f
C7810 _431_/a_36_151# FILLER_0_16_115/a_124_375# 0.035117f
C7811 FILLER_0_4_213/a_124_375# vdd 0.009037f
C7812 FILLER_0_7_72/a_1916_375# vdd 0.015888f
C7813 net8 net59 0.062623f
C7814 net15 _440_/a_1000_472# 0.056791f
C7815 _427_/a_2665_112# _225_/a_36_160# 0.001394f
C7816 FILLER_0_4_107/a_572_375# _151_ 0.00162f
C7817 trimb[1] FILLER_0_18_2/a_2364_375# 0.001523f
C7818 _440_/a_3041_156# _164_ 0.001221f
C7819 _105_ result[6] 0.001477f
C7820 _064_ _446_/a_2665_112# 0.039211f
C7821 _446_/a_448_472# net66 0.017696f
C7822 FILLER_0_6_177/a_36_472# net47 0.011891f
C7823 _058_ _117_ 0.003932f
C7824 net32 _297_/a_36_472# 0.001843f
C7825 _112_ _316_/a_1152_472# 0.001449f
C7826 _126_ FILLER_0_15_180/a_124_375# 0.001238f
C7827 _341_/a_49_472# _137_ 0.059288f
C7828 _445_/a_2665_112# _444_/a_448_472# 0.001178f
C7829 net54 _433_/a_1000_472# 0.0025f
C7830 net25 _214_/a_36_160# 0.019894f
C7831 FILLER_0_23_44/a_36_472# vdd 0.01833f
C7832 FILLER_0_23_44/a_1468_375# vss 0.055902f
C7833 _077_ _453_/a_796_472# 0.003409f
C7834 _122_ _227_/a_36_160# 0.005128f
C7835 fanout81/a_36_160# net76 0.001905f
C7836 FILLER_0_17_38/a_572_375# _179_ 0.002825f
C7837 FILLER_0_5_72/a_1020_375# _029_ 0.010208f
C7838 net15 FILLER_0_6_47/a_1380_472# 0.00464f
C7839 FILLER_0_6_47/a_572_375# vdd 0.003158f
C7840 _308_/a_1152_472# trim_mask\[0\] 0.004076f
C7841 net80 mask\[6\] 0.080689f
C7842 _091_ _429_/a_2665_112# 0.002597f
C7843 net72 FILLER_0_15_59/a_36_472# 0.049812f
C7844 _256_/a_716_497# _128_ 0.001035f
C7845 _170_ net59 0.002301f
C7846 net26 _423_/a_36_151# 0.067024f
C7847 _164_ _381_/a_36_472# 0.007224f
C7848 _098_ _202_/a_36_160# 0.006831f
C7849 net63 FILLER_0_20_193/a_484_472# 0.015851f
C7850 FILLER_0_24_63/a_124_375# ctlp[8] 0.005758f
C7851 mask\[4\] _105_ 0.025209f
C7852 _105_ net22 0.01308f
C7853 _276_/a_36_160# vdd 0.010213f
C7854 _174_ _067_ 0.002678f
C7855 output7/a_224_472# vdd 0.086699f
C7856 FILLER_0_17_200/a_36_472# mask\[3\] 0.27914f
C7857 ctln[2] vdd 0.245598f
C7858 _132_ vss 0.492496f
C7859 _098_ _433_/a_2560_156# 0.004273f
C7860 _130_ _120_ 0.014675f
C7861 _057_ _113_ 0.339862f
C7862 FILLER_0_7_104/a_124_375# _153_ 0.001205f
C7863 FILLER_0_7_104/a_1020_375# _154_ 0.005051f
C7864 net17 _450_/a_2449_156# 0.05017f
C7865 output32/a_224_472# net20 0.050019f
C7866 _256_/a_3368_68# _076_ 0.001183f
C7867 FILLER_0_18_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001684f
C7868 _095_ mask\[1\] 0.001297f
C7869 FILLER_0_9_60/a_124_375# vss 0.003217f
C7870 FILLER_0_9_60/a_572_375# vdd 0.031403f
C7871 net47 _452_/a_836_156# 0.002075f
C7872 _137_ _097_ 0.001654f
C7873 cal_itt\[3\] net76 0.017174f
C7874 _114_ _171_ 0.203692f
C7875 _093_ _293_/a_36_472# 0.004121f
C7876 FILLER_0_15_290/a_124_375# vss 0.032056f
C7877 FILLER_0_15_290/a_36_472# vdd 0.092839f
C7878 net26 _424_/a_1000_472# 0.003207f
C7879 net41 _446_/a_36_151# 0.143017f
C7880 FILLER_0_4_144/a_484_472# trim_mask\[4\] 0.015778f
C7881 net58 _415_/a_2665_112# 0.005219f
C7882 FILLER_0_18_2/a_1916_375# net17 0.013121f
C7883 _226_/a_1044_68# net21 0.001903f
C7884 ctln[7] trim_mask\[3\] 0.059414f
C7885 net66 _166_ 0.011066f
C7886 FILLER_0_8_127/a_36_472# vss 0.004344f
C7887 _081_ FILLER_0_8_156/a_484_472# 0.001772f
C7888 net76 _081_ 0.706096f
C7889 _322_/a_848_380# _128_ 0.012288f
C7890 _300_/a_224_472# _011_ 0.007508f
C7891 FILLER_0_4_197/a_572_375# _088_ 0.013597f
C7892 net20 _010_ 0.016197f
C7893 _216_/a_67_603# net36 0.028132f
C7894 ctln[8] FILLER_0_0_96/a_124_375# 0.002726f
C7895 FILLER_0_1_98/a_124_375# net52 0.001167f
C7896 _028_ FILLER_0_6_90/a_572_375# 0.015802f
C7897 FILLER_0_11_109/a_124_375# _134_ 0.027704f
C7898 _432_/a_1000_472# _093_ 0.007509f
C7899 _320_/a_36_472# net79 0.029189f
C7900 _282_/a_36_160# vss 0.005221f
C7901 net55 _177_ 0.327874f
C7902 fanout58/a_36_160# net5 0.003758f
C7903 _093_ FILLER_0_17_104/a_484_472# 0.014431f
C7904 _093_ _012_ 0.141641f
C7905 result[9] FILLER_0_14_263/a_124_375# 0.003706f
C7906 _057_ _118_ 0.055726f
C7907 FILLER_0_17_282/a_124_375# vss 0.024404f
C7908 FILLER_0_17_282/a_36_472# vdd 0.107351f
C7909 _074_ FILLER_0_5_172/a_124_375# 0.068565f
C7910 _448_/a_1308_423# vdd 0.006042f
C7911 FILLER_0_14_81/a_124_375# _095_ 0.009791f
C7912 _114_ _176_ 0.147182f
C7913 _114_ _306_/a_36_68# 0.032258f
C7914 cal_count\[2\] FILLER_0_15_10/a_36_472# 0.015502f
C7915 net55 FILLER_0_17_38/a_484_472# 0.013624f
C7916 FILLER_0_14_107/a_1020_375# vdd 0.008956f
C7917 _063_ FILLER_0_6_37/a_36_472# 0.014315f
C7918 _415_/a_1000_472# net27 0.017938f
C7919 _126_ _389_/a_36_148# 0.007813f
C7920 FILLER_0_21_133/a_124_375# vss 0.015693f
C7921 FILLER_0_22_177/a_1020_375# vdd 0.001695f
C7922 _270_/a_36_472# net76 0.009569f
C7923 _284_/a_224_472# _094_ 0.001731f
C7924 _341_/a_49_472# net56 0.018486f
C7925 net66 FILLER_0_5_54/a_572_375# 0.002203f
C7926 _423_/a_36_151# FILLER_0_23_44/a_124_375# 0.059049f
C7927 FILLER_0_3_221/a_1020_375# vss 0.003948f
C7928 FILLER_0_3_221/a_1468_375# vdd 0.008815f
C7929 _086_ net76 0.049988f
C7930 net36 FILLER_0_15_212/a_1020_375# 0.004863f
C7931 _016_ state\[2\] 0.002937f
C7932 en_co_clk _043_ 0.041355f
C7933 fanout73/a_36_113# vdd 0.048166f
C7934 output31/a_224_472# _094_ 0.004668f
C7935 mask\[4\] FILLER_0_18_177/a_2724_472# 0.014625f
C7936 FILLER_0_18_177/a_2724_472# net22 0.004297f
C7937 _059_ FILLER_0_5_148/a_124_375# 0.007657f
C7938 _021_ _143_ 0.007778f
C7939 _089_ net76 0.017609f
C7940 fanout66/a_36_113# vss 0.014789f
C7941 FILLER_0_19_55/a_124_375# _216_/a_67_603# 0.003017f
C7942 FILLER_0_3_204/a_124_375# FILLER_0_3_172/a_3260_375# 0.012001f
C7943 FILLER_0_5_54/a_124_375# trim_mask\[1\] 0.024065f
C7944 FILLER_0_5_54/a_1468_375# _029_ 0.008339f
C7945 _304_/a_224_472# _111_ 0.003461f
C7946 _093_ _438_/a_448_472# 0.0106f
C7947 net74 _095_ 0.04188f
C7948 net52 _030_ 0.035783f
C7949 net50 net66 0.016385f
C7950 _119_ FILLER_0_8_156/a_484_472# 0.00979f
C7951 net35 FILLER_0_22_86/a_484_472# 0.008347f
C7952 mask\[8\] FILLER_0_22_86/a_932_472# 0.012284f
C7953 _137_ FILLER_0_15_180/a_124_375# 0.003108f
C7954 net52 _442_/a_1204_472# 0.005558f
C7955 FILLER_0_4_197/a_484_472# net76 0.003719f
C7956 net20 FILLER_0_7_233/a_124_375# 0.017217f
C7957 _144_ _434_/a_36_151# 0.004055f
C7958 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_124_375# 0.003732f
C7959 _162_ FILLER_0_6_177/a_124_375# 0.031168f
C7960 _072_ net4 0.097916f
C7961 _150_ FILLER_0_18_76/a_572_375# 0.008337f
C7962 _449_/a_2665_112# net74 0.001185f
C7963 _257_/a_36_472# _070_ 0.002295f
C7964 _307_/a_672_472# _096_ 0.001367f
C7965 _095_ cal_count\[1\] 0.853949f
C7966 FILLER_0_18_177/a_2364_375# vdd 0.020562f
C7967 net64 mask\[1\] 0.038611f
C7968 _363_/a_36_68# FILLER_0_7_104/a_572_375# 0.002308f
C7969 net20 vdd 2.14128f
C7970 FILLER_0_9_223/a_124_375# _068_ 0.010485f
C7971 _350_/a_665_69# mask\[6\] 0.001069f
C7972 _339_/a_36_160# vdd 0.01226f
C7973 _053_ net68 0.239882f
C7974 output18/a_224_472# net33 0.135766f
C7975 FILLER_0_18_2/a_2276_472# vdd 0.004679f
C7976 net32 _006_ 0.0012f
C7977 _070_ FILLER_0_8_156/a_36_472# 0.001338f
C7978 _076_ FILLER_0_8_156/a_124_375# 0.0062f
C7979 _354_/a_49_472# _433_/a_36_151# 0.001715f
C7980 _013_ FILLER_0_18_53/a_124_375# 0.015996f
C7981 FILLER_0_7_59/a_124_375# trim_val\[0\] 0.002169f
C7982 FILLER_0_14_91/a_484_472# vss 0.003257f
C7983 _119_ _319_/a_672_472# 0.00488f
C7984 _057_ _068_ 0.393271f
C7985 state\[1\] vss 0.294171f
C7986 net15 FILLER_0_13_72/a_484_472# 0.002925f
C7987 _453_/a_2665_112# vss 0.037567f
C7988 _092_ vss 0.346097f
C7989 FILLER_0_16_57/a_1380_472# net15 0.017841f
C7990 net69 FILLER_0_3_78/a_36_472# 0.002068f
C7991 _417_/a_1204_472# _006_ 0.014354f
C7992 _432_/a_36_151# FILLER_0_16_154/a_1468_375# 0.001107f
C7993 _012_ FILLER_0_21_60/a_484_472# 0.01517f
C7994 mask\[4\] _047_ 0.080091f
C7995 net22 _047_ 0.132529f
C7996 _141_ FILLER_0_16_154/a_36_472# 0.00126f
C7997 fanout60/a_36_160# result[3] 0.00188f
C7998 _031_ FILLER_0_2_101/a_124_375# 0.00179f
C7999 _002_ _270_/a_244_68# 0.001153f
C8000 FILLER_0_6_79/a_124_375# vdd 0.015119f
C8001 FILLER_0_20_2/a_484_472# vdd 0.001049f
C8002 cal_count\[3\] _113_ 0.093684f
C8003 _079_ _260_/a_244_472# 0.00325f
C8004 _053_ FILLER_0_7_72/a_484_472# 0.00887f
C8005 _070_ _319_/a_234_472# 0.004015f
C8006 state\[2\] _427_/a_448_472# 0.00237f
C8007 net53 _427_/a_796_472# 0.001983f
C8008 _444_/a_1000_472# net67 0.025169f
C8009 FILLER_0_12_236/a_36_472# _060_ 0.014046f
C8010 FILLER_0_1_266/a_484_472# vdd 0.003622f
C8011 comp net44 0.079931f
C8012 _077_ _062_ 0.037598f
C8013 FILLER_0_3_204/a_124_375# vdd 0.023302f
C8014 FILLER_0_3_54/a_124_375# vdd 0.029897f
C8015 _114_ FILLER_0_13_142/a_124_375# 0.00191f
C8016 output9/a_224_472# net8 0.020421f
C8017 _002_ net21 0.056631f
C8018 net75 net20 0.092951f
C8019 _083_ _081_ 0.03934f
C8020 FILLER_0_7_72/a_2724_472# vdd 0.007669f
C8021 _359_/a_36_488# _152_ 0.032195f
C8022 _128_ _124_ 0.111918f
C8023 _008_ _418_/a_1204_472# 0.002933f
C8024 _450_/a_2449_156# _039_ 0.013285f
C8025 _132_ _148_ 0.002873f
C8026 net36 FILLER_0_15_235/a_124_375# 0.007232f
C8027 FILLER_0_18_2/a_2276_472# _452_/a_1040_527# 0.008652f
C8028 _402_/a_1296_93# _179_ 0.001692f
C8029 result[9] _417_/a_2248_156# 0.046399f
C8030 _238_/a_67_603# FILLER_0_2_93/a_36_472# 0.002778f
C8031 _119_ FILLER_0_8_138/a_36_472# 0.003894f
C8032 output24/a_224_472# _436_/a_448_472# 0.009204f
C8033 FILLER_0_12_136/a_484_472# vdd 0.005304f
C8034 FILLER_0_12_136/a_36_472# vss 0.003185f
C8035 FILLER_0_10_214/a_124_375# _247_/a_36_160# 0.005732f
C8036 _065_ net16 0.068602f
C8037 cal_count\[3\] _118_ 0.009058f
C8038 FILLER_0_17_142/a_572_375# _137_ 0.006974f
C8039 FILLER_0_4_197/a_1380_472# net82 0.003084f
C8040 FILLER_0_9_28/a_1916_375# net16 0.001431f
C8041 _423_/a_1204_472# _012_ 0.003181f
C8042 trim_mask\[2\] fanout66/a_36_113# 0.015961f
C8043 net79 _101_ 0.014383f
C8044 _031_ _158_ 0.015116f
C8045 _085_ _176_ 0.024708f
C8046 _430_/a_36_151# mask\[3\] 0.005848f
C8047 _337_/a_49_472# mask\[2\] 0.00188f
C8048 _415_/a_2248_156# output27/a_224_472# 0.001506f
C8049 output32/a_224_472# vss -0.003023f
C8050 FILLER_0_19_111/a_572_375# vdd -0.008314f
C8051 net2 rstn 0.002598f
C8052 _163_ net22 0.005017f
C8053 _306_/a_36_68# _085_ 0.00755f
C8054 net79 FILLER_0_12_220/a_1468_375# 0.012754f
C8055 _415_/a_796_472# vdd 0.001842f
C8056 FILLER_0_14_50/a_124_375# _095_ 0.052375f
C8057 FILLER_0_19_187/a_124_375# vdd 0.030349f
C8058 _289_/a_36_472# vdd 0.006886f
C8059 net62 _417_/a_2560_156# 0.003361f
C8060 _446_/a_2248_156# _160_ 0.002464f
C8061 _256_/a_2960_68# _076_ 0.001292f
C8062 net14 FILLER_0_10_94/a_124_375# 0.007086f
C8063 FILLER_0_21_133/a_124_375# mask\[7\] 0.00145f
C8064 mask\[7\] FILLER_0_22_177/a_572_375# 0.001315f
C8065 _328_/a_36_113# net74 0.002214f
C8066 _132_ _332_/a_36_472# 0.055537f
C8067 net16 _180_ 0.00101f
C8068 _051_ vss 0.050185f
C8069 _010_ vss 0.064717f
C8070 FILLER_0_2_93/a_572_375# _367_/a_36_68# 0.001069f
C8071 FILLER_0_5_181/a_124_375# vss 0.011456f
C8072 FILLER_0_5_181/a_36_472# vdd 0.081434f
C8073 _062_ net37 0.082701f
C8074 FILLER_0_21_28/a_1020_375# vdd 0.04353f
C8075 _031_ net14 0.00913f
C8076 FILLER_0_3_172/a_36_472# vdd 0.006145f
C8077 FILLER_0_3_172/a_3260_375# vss 0.054783f
C8078 _386_/a_124_24# vdd 0.014293f
C8079 output37/a_224_472# net37 0.011407f
C8080 FILLER_0_16_241/a_36_472# net30 0.001025f
C8081 _438_/a_1000_472# net14 0.003275f
C8082 net4 FILLER_0_3_221/a_1020_375# 0.006974f
C8083 FILLER_0_2_111/a_36_472# _157_ 0.104961f
C8084 FILLER_0_5_54/a_124_375# _164_ 0.004076f
C8085 FILLER_0_14_81/a_124_375# cal_count\[1\] 0.070473f
C8086 _359_/a_36_488# _070_ 0.028563f
C8087 FILLER_0_13_212/a_932_472# _043_ 0.014431f
C8088 _093_ FILLER_0_18_107/a_1828_472# 0.001872f
C8089 FILLER_0_18_100/a_124_375# vdd 0.044014f
C8090 _095_ _097_ 0.030222f
C8091 _385_/a_36_68# vss 0.002408f
C8092 _088_ FILLER_0_3_172/a_2724_472# 0.005827f
C8093 _059_ _313_/a_67_603# 0.061666f
C8094 _449_/a_2248_156# cal_count\[3\] 0.002041f
C8095 net28 _196_/a_36_160# 0.060575f
C8096 output15/a_224_472# fanout50/a_36_160# 0.003531f
C8097 _005_ _416_/a_1000_472# 0.027013f
C8098 net52 trim_mask\[3\] 0.666362f
C8099 _442_/a_448_472# net69 0.004308f
C8100 _053_ FILLER_0_7_104/a_1468_375# 0.001492f
C8101 net56 _145_ 0.009307f
C8102 vdd FILLER_0_4_91/a_484_472# 0.007304f
C8103 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1468_375# 0.016748f
C8104 _069_ _121_ 0.137961f
C8105 _155_ _163_ 0.296236f
C8106 output36/a_224_472# vss -0.002521f
C8107 _445_/a_2560_156# net49 0.001208f
C8108 _105_ _297_/a_36_472# 0.03208f
C8109 net81 _019_ 0.004079f
C8110 FILLER_0_9_28/a_2364_375# _077_ 0.00397f
C8111 cal_itt\[1\] vdd 0.410279f
C8112 _412_/a_2665_112# fanout58/a_36_160# 0.001221f
C8113 FILLER_0_22_86/a_932_472# _026_ 0.001587f
C8114 net56 FILLER_0_17_142/a_572_375# 0.014948f
C8115 net16 net51 0.035455f
C8116 mask\[0\] _429_/a_1000_472# 0.020553f
C8117 FILLER_0_4_107/a_484_472# FILLER_0_2_111/a_124_375# 0.001404f
C8118 _415_/a_36_151# FILLER_0_10_256/a_124_375# 0.035117f
C8119 net4 state\[1\] 0.010195f
C8120 net55 FILLER_0_18_53/a_36_472# 0.00953f
C8121 FILLER_0_7_233/a_36_472# vdd 0.016804f
C8122 FILLER_0_7_233/a_124_375# vss 0.003952f
C8123 _181_ _185_ 0.061846f
C8124 net38 _452_/a_448_472# 0.016895f
C8125 _321_/a_2590_472# _118_ 0.002396f
C8126 net35 _146_ 0.096468f
C8127 FILLER_0_12_136/a_1020_375# net23 0.005919f
C8128 sample vdd 0.154389f
C8129 net72 FILLER_0_21_28/a_1020_375# 0.040811f
C8130 _076_ _163_ 0.030003f
C8131 FILLER_0_20_177/a_36_472# _098_ 0.015061f
C8132 FILLER_0_5_117/a_36_472# _160_ 0.005314f
C8133 FILLER_0_4_123/a_36_472# trim_mask\[4\] 0.003692f
C8134 input2/a_36_113# en 0.002108f
C8135 fanout62/a_36_160# net62 0.02201f
C8136 vdd vss 15.42941f
C8137 _091_ net27 0.023019f
C8138 _115_ _076_ 0.051404f
C8139 _207_/a_255_603# mask\[6\] 0.003114f
C8140 _136_ _334_/a_36_160# 0.005574f
C8141 _058_ _059_ 0.990213f
C8142 output24/a_224_472# net24 0.005559f
C8143 fanout49/a_36_160# FILLER_0_3_78/a_484_472# 0.003699f
C8144 _078_ FILLER_0_4_213/a_484_472# 0.003702f
C8145 net50 FILLER_0_8_24/a_572_375# 0.001597f
C8146 _415_/a_36_151# net62 0.00514f
C8147 FILLER_0_18_100/a_36_472# FILLER_0_17_72/a_3172_472# 0.05841f
C8148 _427_/a_2248_156# state\[1\] 0.001849f
C8149 net47 _380_/a_224_472# 0.001405f
C8150 FILLER_0_9_28/a_572_375# net41 0.025588f
C8151 net58 _412_/a_1308_423# 0.037719f
C8152 _093_ FILLER_0_17_72/a_36_472# 0.001971f
C8153 FILLER_0_13_65/a_36_472# _174_ 0.011724f
C8154 FILLER_0_23_60/a_36_472# vss 0.006794f
C8155 FILLER_0_5_128/a_484_472# _133_ 0.037369f
C8156 FILLER_0_6_177/a_36_472# vdd 0.109918f
C8157 FILLER_0_6_177/a_572_375# vss 0.008666f
C8158 _074_ net82 0.123449f
C8159 net81 _429_/a_2248_156# 0.017036f
C8160 net64 FILLER_0_12_236/a_36_472# 0.052381f
C8161 FILLER_0_2_171/a_124_375# vdd 0.042659f
C8162 net75 cal_itt\[1\] 0.704169f
C8163 net74 FILLER_0_13_72/a_124_375# 0.014594f
C8164 net63 FILLER_0_18_177/a_1468_375# 0.020059f
C8165 FILLER_0_15_290/a_124_375# net79 0.051113f
C8166 net81 FILLER_0_10_247/a_36_472# 0.015109f
C8167 net15 _394_/a_56_524# 0.006099f
C8168 FILLER_0_7_72/a_124_375# vdd 0.01526f
C8169 _068_ net59 0.001388f
C8170 net27 FILLER_0_9_270/a_36_472# 0.041681f
C8171 _144_ FILLER_0_21_125/a_572_375# 0.003787f
C8172 net20 FILLER_0_13_212/a_572_375# 0.002085f
C8173 _099_ mask\[2\] 0.776725f
C8174 _097_ mask\[1\] 0.001232f
C8175 FILLER_0_21_142/a_124_375# FILLER_0_22_128/a_1828_472# 0.001543f
C8176 _435_/a_2248_156# net21 0.012406f
C8177 FILLER_0_19_47/a_572_375# _013_ 0.012993f
C8178 _053_ FILLER_0_8_37/a_36_472# 0.001011f
C8179 _098_ FILLER_0_19_171/a_932_472# 0.003573f
C8180 FILLER_0_16_255/a_36_472# _006_ 0.006621f
C8181 _088_ FILLER_0_5_206/a_124_375# 0.001374f
C8182 _079_ FILLER_0_5_206/a_36_472# 0.008243f
C8183 FILLER_0_16_89/a_932_472# net36 0.001709f
C8184 net60 _420_/a_2560_156# 0.001358f
C8185 _428_/a_36_151# _017_ 0.021229f
C8186 FILLER_0_21_28/a_1020_375# _424_/a_36_151# 0.001252f
C8187 FILLER_0_15_72/a_124_375# FILLER_0_15_59/a_572_375# 0.003228f
C8188 FILLER_0_16_57/a_36_472# cal_count\[1\] 0.002116f
C8189 result[9] _418_/a_2248_156# 0.043716f
C8190 mask\[8\] _026_ 0.001638f
C8191 _077_ FILLER_0_10_78/a_572_375# 0.001886f
C8192 _098_ _438_/a_1000_472# 0.001492f
C8193 _104_ output20/a_224_472# 0.019295f
C8194 _343_/a_49_472# net80 0.001646f
C8195 net75 vss 0.662689f
C8196 _114_ _017_ 0.071595f
C8197 net82 FILLER_0_3_172/a_1020_375# 0.010679f
C8198 _053_ _072_ 0.001774f
C8199 net72 vss 0.472104f
C8200 FILLER_0_2_165/a_124_375# vdd 0.020315f
C8201 _452_/a_836_156# vdd 0.002533f
C8202 output20/a_224_472# _422_/a_1308_423# 0.005632f
C8203 FILLER_0_18_139/a_1468_375# _137_ 0.004111f
C8204 _136_ net36 1.151311f
C8205 FILLER_0_4_123/a_36_472# fanout69/a_36_113# 0.007864f
C8206 FILLER_0_16_37/a_124_375# _179_ 0.005434f
C8207 _091_ _043_ 0.041409f
C8208 net36 net21 0.034415f
C8209 _369_/a_244_472# vdd 0.001255f
C8210 _070_ FILLER_0_6_231/a_36_472# 0.001096f
C8211 _076_ FILLER_0_6_231/a_124_375# 0.001382f
C8212 net17 _452_/a_2225_156# 0.001943f
C8213 _450_/a_1697_156# net6 0.00236f
C8214 _041_ FILLER_0_18_37/a_1380_472# 0.003776f
C8215 _299_/a_36_472# _109_ 0.030751f
C8216 output18/a_224_472# net18 0.01698f
C8217 trim_mask\[2\] FILLER_0_4_91/a_36_472# 0.003327f
C8218 _077_ FILLER_0_8_156/a_572_375# 0.007238f
C8219 _432_/a_1204_472# _091_ 0.00563f
C8220 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_124_375# 0.007947f
C8221 _274_/a_36_68# net20 0.021022f
C8222 _114_ _250_/a_36_68# 0.017773f
C8223 _053_ net47 0.011652f
C8224 output27/a_224_472# FILLER_0_9_282/a_124_375# 0.029138f
C8225 FILLER_0_15_116/a_484_472# _131_ 0.042796f
C8226 net15 _423_/a_2665_112# 0.061217f
C8227 _350_/a_257_69# net23 0.003052f
C8228 net63 net80 0.337396f
C8229 net7 net41 0.243942f
C8230 net57 _428_/a_2560_156# 0.010877f
C8231 FILLER_0_14_50/a_124_375# cal_count\[1\] 0.023752f
C8232 net61 _422_/a_2665_112# 0.023601f
C8233 _356_/a_36_472# net36 0.004539f
C8234 _115_ FILLER_0_11_78/a_484_472# 0.003641f
C8235 _423_/a_36_151# net17 0.002865f
C8236 _443_/a_36_151# _032_ 0.0737f
C8237 net69 _370_/a_124_24# 0.001491f
C8238 _316_/a_124_24# net37 0.011141f
C8239 _413_/a_2560_156# vss 0.001097f
C8240 _132_ _428_/a_1308_423# 0.027389f
C8241 FILLER_0_17_72/a_2364_375# net36 0.005483f
C8242 FILLER_0_16_73/a_124_375# vss 0.026383f
C8243 _413_/a_36_151# FILLER_0_2_177/a_572_375# 0.073306f
C8244 mask\[1\] FILLER_0_15_180/a_124_375# 0.004011f
C8245 FILLER_0_8_138/a_124_375# calibrate 0.013177f
C8246 _428_/a_2248_156# _043_ 0.011841f
C8247 FILLER_0_22_128/a_572_375# vss 0.00243f
C8248 FILLER_0_22_128/a_1020_375# vdd 0.002503f
C8249 FILLER_0_1_98/a_36_472# vdd 0.009937f
C8250 _449_/a_2248_156# FILLER_0_13_80/a_124_375# 0.001068f
C8251 _024_ vss 0.132549f
C8252 trimb[2] output17/a_224_472# 0.008375f
C8253 _424_/a_36_151# vss 0.030774f
C8254 _424_/a_448_472# vdd 0.014219f
C8255 _052_ _424_/a_2665_112# 0.003027f
C8256 _083_ FILLER_0_3_221/a_484_472# 0.02695f
C8257 _098_ _434_/a_2560_156# 0.003888f
C8258 _441_/a_1000_472# vss 0.01858f
C8259 trim_mask\[2\] vdd 0.376424f
C8260 FILLER_0_5_88/a_36_472# net47 0.003953f
C8261 FILLER_0_11_64/a_124_375# vdd 0.045435f
C8262 mask\[5\] FILLER_0_20_177/a_124_375# 0.013531f
C8263 net29 _195_/a_67_603# 0.048817f
C8264 FILLER_0_13_212/a_1380_472# mask\[0\] 0.002361f
C8265 net55 _452_/a_448_472# 0.05323f
C8266 _053_ FILLER_0_6_47/a_124_375# 0.002541f
C8267 FILLER_0_13_206/a_36_472# vss 0.003985f
C8268 _447_/a_1308_423# vdd 0.004739f
C8269 _193_/a_36_160# FILLER_0_13_290/a_36_472# 0.004828f
C8270 _064_ net17 0.108825f
C8271 net79 state\[1\] 0.005861f
C8272 net62 FILLER_0_15_228/a_36_472# 0.002128f
C8273 trim_val\[3\] _164_ 0.018411f
C8274 ctln[1] _073_ 0.001457f
C8275 net15 trim_mask\[1\] 0.042093f
C8276 net73 _345_/a_36_160# 0.032139f
C8277 _440_/a_2560_156# vss 0.002793f
C8278 _116_ net21 0.036746f
C8279 FILLER_0_4_107/a_1380_472# trim_mask\[4\] 0.011766f
C8280 net29 net30 0.053996f
C8281 _035_ net66 1.624557f
C8282 _112_ _425_/a_1000_472# 0.001973f
C8283 _439_/a_796_472# vss 0.003859f
C8284 _367_/a_244_472# _157_ 0.002529f
C8285 fanout58/a_36_160# en 0.00568f
C8286 input3/a_36_113# vdd 0.117445f
C8287 net31 FILLER_0_16_255/a_124_375# 0.029277f
C8288 net62 FILLER_0_13_290/a_124_375# 0.032026f
C8289 net17 output41/a_224_472# 0.030456f
C8290 _073_ _076_ 0.011358f
C8291 _279_/a_652_68# vdd 0.001562f
C8292 _181_ _402_/a_1296_93# 0.040412f
C8293 _142_ FILLER_0_17_133/a_124_375# 0.022066f
C8294 _122_ _062_ 0.190871f
C8295 net76 FILLER_0_3_172/a_932_472# 0.005391f
C8296 net36 _045_ 0.091033f
C8297 _426_/a_36_151# FILLER_0_8_247/a_36_472# 0.001723f
C8298 _432_/a_2248_156# net21 0.002329f
C8299 fanout63/a_36_160# _282_/a_36_160# 0.23939f
C8300 _130_ FILLER_0_12_136/a_124_375# 0.010514f
C8301 _255_/a_224_552# _163_ 0.002169f
C8302 _114_ FILLER_0_11_109/a_124_375# 0.009676f
C8303 _116_ _070_ 0.166494f
C8304 mask\[7\] vdd 1.098711f
C8305 FILLER_0_4_197/a_572_375# net59 0.001512f
C8306 FILLER_0_6_47/a_3172_472# vss 0.014726f
C8307 _077_ _308_/a_848_380# 0.010515f
C8308 net56 FILLER_0_18_139/a_1468_375# 0.065206f
C8309 _091_ FILLER_0_18_177/a_124_375# 0.010316f
C8310 _316_/a_1084_68# vdd 0.001166f
C8311 mask\[4\] net54 0.009909f
C8312 _148_ vdd 0.01565f
C8313 _276_/a_36_160# FILLER_0_17_218/a_36_472# 0.035111f
C8314 fanout64/a_36_160# fanout65/a_36_113# 0.001627f
C8315 vss cal_count\[0\] 0.160743f
C8316 net35 _435_/a_448_472# 0.007865f
C8317 net4 vdd 1.218939f
C8318 net25 FILLER_0_23_44/a_1380_472# 0.0014f
C8319 _019_ mask\[1\] 0.007797f
C8320 mask\[5\] FILLER_0_19_171/a_1020_375# 0.007169f
C8321 _144_ mask\[6\] 0.230129f
C8322 _414_/a_2248_156# vss 0.00384f
C8323 _035_ _167_ 0.01574f
C8324 net72 _424_/a_448_472# 0.011745f
C8325 net10 _000_ 0.001954f
C8326 mask\[9\] _424_/a_2665_112# 0.015491f
C8327 _118_ _120_ 0.339442f
C8328 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_124_375# 0.009654f
C8329 output31/a_224_472# _417_/a_2248_156# 0.024448f
C8330 _091_ FILLER_0_19_171/a_1380_472# 0.001044f
C8331 net53 FILLER_0_14_123/a_36_472# 0.062713f
C8332 _061_ _062_ 0.344031f
C8333 _000_ FILLER_0_0_232/a_124_375# 0.001391f
C8334 net20 _099_ 0.011124f
C8335 FILLER_0_9_223/a_572_375# calibrate 0.002082f
C8336 output46/a_224_472# FILLER_0_20_2/a_484_472# 0.001699f
C8337 _432_/a_36_151# net80 0.035794f
C8338 _448_/a_2560_156# net59 0.007516f
C8339 _176_ FILLER_0_15_59/a_36_472# 0.00622f
C8340 FILLER_0_5_128/a_36_472# _152_ 0.013822f
C8341 FILLER_0_21_142/a_572_375# net23 0.007884f
C8342 net81 _100_ 0.24831f
C8343 _427_/a_2248_156# vdd -0.002315f
C8344 _427_/a_1204_472# vss 0.0041f
C8345 FILLER_0_5_128/a_124_375# _163_ 0.009765f
C8346 _374_/a_36_68# vss 0.047832f
C8347 _077_ FILLER_0_9_72/a_1468_375# 0.008273f
C8348 _291_/a_36_160# _199_/a_36_160# 0.005575f
C8349 net58 _415_/a_2248_156# 0.001869f
C8350 _038_ _067_ 0.503045f
C8351 FILLER_0_8_138/a_124_375# _125_ 0.001589f
C8352 FILLER_0_4_152/a_36_472# _386_/a_124_24# 0.004755f
C8353 net81 _004_ 0.993594f
C8354 _376_/a_36_160# trim_mask\[1\] 0.003111f
C8355 FILLER_0_8_24/a_572_375# _054_ 0.004858f
C8356 FILLER_0_19_47/a_484_472# net55 0.061087f
C8357 net75 _316_/a_1084_68# 0.001531f
C8358 FILLER_0_13_65/a_124_375# _449_/a_36_151# 0.059049f
C8359 _322_/a_124_24# _129_ 0.017754f
C8360 net41 _186_ 0.054661f
C8361 _429_/a_36_151# FILLER_0_13_206/a_124_375# 0.001597f
C8362 _448_/a_448_472# FILLER_0_2_177/a_36_472# 0.001927f
C8363 _448_/a_36_151# FILLER_0_2_177/a_484_472# 0.059367f
C8364 _411_/a_2248_156# net19 0.001197f
C8365 net47 FILLER_0_5_164/a_36_472# 0.046908f
C8366 _077_ _188_ 0.1656f
C8367 _117_ net21 0.016722f
C8368 FILLER_0_18_2/a_36_472# _452_/a_3129_107# 0.035307f
C8369 _332_/a_36_472# vdd 0.017097f
C8370 cal_itt\[2\] ctln[1] 0.053339f
C8371 net38 _444_/a_36_151# 0.009033f
C8372 net75 net4 0.031823f
C8373 FILLER_0_10_247/a_36_472# net64 0.059367f
C8374 ctln[1] net1 0.003756f
C8375 _449_/a_1204_472# _067_ 0.014354f
C8376 _077_ fanout67/a_36_160# 0.017322f
C8377 _411_/a_1000_472# vss 0.002964f
C8378 FILLER_0_13_212/a_1020_375# vdd -0.014642f
C8379 FILLER_0_13_212/a_572_375# vss 0.007991f
C8380 net46 net43 0.215092f
C8381 _081_ _265_/a_468_472# 0.005156f
C8382 _033_ _444_/a_2665_112# 0.004024f
C8383 net46 output44/a_224_472# 0.003211f
C8384 net65 net2 0.035908f
C8385 _436_/a_1308_423# vdd 0.005258f
C8386 _415_/a_1308_423# vdd 0.004258f
C8387 output45/a_224_472# net17 0.092967f
C8388 _058_ _134_ 0.034211f
C8389 _070_ _117_ 0.080445f
C8390 _050_ net71 0.033192f
C8391 FILLER_0_24_130/a_36_472# ctlp[7] 0.012298f
C8392 _013_ _182_ 0.001681f
C8393 _235_/a_67_603# _064_ 0.003796f
C8394 net52 _453_/a_2248_156# 0.011419f
C8395 FILLER_0_11_142/a_36_472# cal_count\[3\] 0.008454f
C8396 FILLER_0_16_57/a_932_472# FILLER_0_17_64/a_124_375# 0.001723f
C8397 _068_ _120_ 0.447243f
C8398 _447_/a_2248_156# _441_/a_36_151# 0.035837f
C8399 trim_mask\[2\] _447_/a_448_472# 0.002533f
C8400 trim_val\[2\] _447_/a_36_151# 0.022122f
C8401 FILLER_0_18_107/a_2364_375# _022_ 0.001902f
C8402 FILLER_0_16_107/a_124_375# net14 0.004684f
C8403 vss _433_/a_36_151# 0.00618f
C8404 vdd _433_/a_448_472# 0.003821f
C8405 net60 _418_/a_1000_472# 0.007557f
C8406 _413_/a_2665_112# net20 0.015855f
C8407 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_36_472# 0.007947f
C8408 _445_/a_2560_156# net47 0.014069f
C8409 _337_/a_257_69# vdd 0.002972f
C8410 _369_/a_36_68# _367_/a_36_68# 0.038188f
C8411 _187_ _450_/a_3129_107# 0.00126f
C8412 _412_/a_448_472# net65 0.043862f
C8413 _315_/a_244_497# vss 0.008724f
C8414 FILLER_0_5_172/a_124_375# _163_ 0.006403f
C8415 _132_ FILLER_0_17_104/a_572_375# 0.003857f
C8416 net57 _267_/a_672_472# 0.004637f
C8417 _440_/a_448_472# _029_ 0.043511f
C8418 _352_/a_49_472# FILLER_0_22_128/a_36_472# 0.063744f
C8419 mask\[7\] FILLER_0_22_128/a_572_375# 0.01909f
C8420 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_484_472# 0.013276f
C8421 FILLER_0_20_193/a_484_472# net21 0.00371f
C8422 net65 cal 0.023638f
C8423 FILLER_0_5_198/a_124_375# vdd 0.010749f
C8424 net47 _221_/a_36_160# 0.012197f
C8425 mask\[7\] _024_ 0.122185f
C8426 _384_/a_224_472# _160_ 0.00324f
C8427 FILLER_0_4_152/a_36_472# vss 0.009467f
C8428 FILLER_0_7_59/a_484_472# vss 0.005804f
C8429 net2 net59 0.334636f
C8430 _115_ _128_ 0.263909f
C8431 FILLER_0_10_78/a_124_375# _115_ 0.001718f
C8432 net35 FILLER_0_22_128/a_36_472# 0.00784f
C8433 FILLER_0_5_128/a_36_472# _070_ 0.036f
C8434 _118_ _227_/a_36_160# 0.017547f
C8435 _064_ net39 0.558387f
C8436 net36 _451_/a_448_472# 0.042223f
C8437 net16 net66 0.030521f
C8438 _274_/a_36_68# vss 0.052669f
C8439 FILLER_0_20_98/a_36_472# _437_/a_36_151# 0.001723f
C8440 FILLER_0_8_263/a_36_472# net19 0.047387f
C8441 net68 FILLER_0_6_47/a_1468_375# 0.022624f
C8442 _092_ FILLER_0_17_218/a_484_472# 0.007838f
C8443 _065_ net14 0.005438f
C8444 _178_ _184_ 0.436202f
C8445 _308_/a_124_24# _070_ 0.001465f
C8446 _013_ FILLER_0_21_28/a_1828_472# 0.003978f
C8447 _136_ FILLER_0_16_154/a_1468_375# 0.0028f
C8448 trim_mask\[1\] FILLER_0_6_47/a_2364_375# 0.007169f
C8449 net15 _164_ 0.026132f
C8450 fanout52/a_36_160# _386_/a_124_24# 0.004695f
C8451 _412_/a_448_472# net59 0.001462f
C8452 FILLER_0_3_142/a_36_472# vdd 0.10948f
C8453 FILLER_0_3_142/a_124_375# vss 0.008128f
C8454 net23 _207_/a_67_603# 0.002734f
C8455 _411_/a_2560_156# _073_ 0.002649f
C8456 output10/a_224_472# _411_/a_2248_156# 0.019736f
C8457 cal_count\[3\] _314_/a_224_472# 0.002143f
C8458 _289_/a_36_472# _099_ 0.035055f
C8459 _086_ FILLER_0_7_104/a_1468_375# 0.065371f
C8460 _114_ FILLER_0_12_136/a_932_472# 0.003953f
C8461 vdd FILLER_0_19_134/a_36_472# 0.092128f
C8462 vss FILLER_0_19_134/a_124_375# 0.021427f
C8463 FILLER_0_0_96/a_36_472# net14 0.009584f
C8464 _412_/a_2560_156# net5 0.007446f
C8465 _033_ _160_ 0.020281f
C8466 _092_ _430_/a_2665_112# 0.004778f
C8467 FILLER_0_12_220/a_124_375# _090_ 0.001521f
C8468 cal net59 0.297816f
C8469 _155_ FILLER_0_7_104/a_124_375# 0.007925f
C8470 _027_ _438_/a_796_472# 0.031292f
C8471 _150_ _438_/a_1204_472# 0.003696f
C8472 ctlp[1] _421_/a_448_472# 0.011026f
C8473 net54 _437_/a_2560_156# 0.009745f
C8474 net58 _073_ 0.057725f
C8475 FILLER_0_4_99/a_36_472# vss 0.002273f
C8476 net67 trim_val\[0\] 0.382079f
C8477 _119_ FILLER_0_7_104/a_1468_375# 0.022368f
C8478 _446_/a_448_472# net17 0.026011f
C8479 net79 vdd 1.283563f
C8480 _431_/a_2248_156# FILLER_0_15_142/a_484_472# 0.016128f
C8481 FILLER_0_4_99/a_124_375# _365_/a_36_68# 0.001918f
C8482 FILLER_0_7_146/a_36_472# vdd 0.072981f
C8483 FILLER_0_7_146/a_124_375# vss 0.050543f
C8484 _096_ _114_ 0.066848f
C8485 _065_ _447_/a_2665_112# 0.034757f
C8486 _316_/a_124_24# _122_ 0.040082f
C8487 _316_/a_848_380# calibrate 0.012121f
C8488 _076_ _121_ 0.013717f
C8489 mask\[5\] mask\[4\] 0.176881f
C8490 mask\[5\] net22 0.04021f
C8491 _233_/a_36_160# _444_/a_36_151# 0.032942f
C8492 mask\[4\] FILLER_0_18_209/a_572_375# 0.032112f
C8493 trim[0] trim[2] 0.002289f
C8494 net16 _167_ 0.001124f
C8495 net22 FILLER_0_18_209/a_572_375# 0.005202f
C8496 _165_ _220_/a_67_603# 0.004199f
C8497 _317_/a_36_113# _014_ 0.037134f
C8498 output13/a_224_472# _037_ 0.019694f
C8499 _322_/a_848_380# _126_ 0.002519f
C8500 net63 _106_ 0.034574f
C8501 _141_ vdd 0.439746f
C8502 FILLER_0_21_28/a_36_472# net40 0.032105f
C8503 net16 _067_ 0.039705f
C8504 net52 _168_ 0.726039f
C8505 _055_ _311_/a_66_473# 0.040326f
C8506 FILLER_0_18_2/a_1828_472# net38 0.006713f
C8507 FILLER_0_16_89/a_572_375# _136_ 0.069752f
C8508 _417_/a_448_472# net30 0.042386f
C8509 net65 FILLER_0_3_172/a_2724_472# 0.001777f
C8510 _097_ FILLER_0_15_180/a_124_375# 0.007065f
C8511 vdd _295_/a_36_472# 0.0083f
C8512 _182_ _179_ 0.109377f
C8513 FILLER_0_16_37/a_124_375# _181_ 0.001198f
C8514 FILLER_0_9_72/a_1380_472# vss 0.007254f
C8515 net27 _426_/a_2248_156# 0.002303f
C8516 _068_ _227_/a_36_160# 0.053563f
C8517 _131_ _124_ 0.002448f
C8518 _104_ net30 0.001375f
C8519 cal_itt\[3\] _072_ 2.019868f
C8520 input1/a_36_113# input4/a_36_68# 0.015796f
C8521 _077_ _308_/a_692_472# 0.002268f
C8522 net48 _251_/a_906_472# 0.001362f
C8523 _094_ _418_/a_1308_423# 0.029276f
C8524 _126_ mask\[0\] 0.067513f
C8525 _062_ _160_ 0.001024f
C8526 _178_ net47 0.09023f
C8527 output8/a_224_472# FILLER_0_3_221/a_1380_472# 0.001699f
C8528 net44 FILLER_0_20_2/a_484_472# 0.039736f
C8529 output46/a_224_472# vss 0.00432f
C8530 net43 FILLER_0_20_15/a_36_472# 0.002803f
C8531 net57 FILLER_0_13_142/a_1380_472# 0.011768f
C8532 output44/a_224_472# FILLER_0_20_15/a_36_472# 0.0323f
C8533 output31/a_224_472# _418_/a_2248_156# 0.023576f
C8534 fanout52/a_36_160# vss 0.010082f
C8535 net26 _217_/a_36_160# 0.021067f
C8536 _303_/a_36_472# _110_ 0.001606f
C8537 vdd _380_/a_224_472# 0.001733f
C8538 _376_/a_36_160# _164_ 0.004503f
C8539 _207_/a_67_603# net33 0.005153f
C8540 FILLER_0_20_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001543f
C8541 FILLER_0_15_282/a_36_472# net30 0.001692f
C8542 FILLER_0_15_282/a_124_375# result[3] 0.004601f
C8543 vdd _416_/a_2665_112# 0.027256f
C8544 net53 FILLER_0_16_154/a_36_472# 0.006261f
C8545 net62 _416_/a_1000_472# 0.002399f
C8546 net24 vss 0.172755f
C8547 FILLER_0_21_286/a_124_375# _009_ 0.001024f
C8548 trimb[1] FILLER_0_18_2/a_1020_375# 0.01376f
C8549 cal_itt\[3\] net47 0.00247f
C8550 FILLER_0_16_89/a_572_375# FILLER_0_17_72/a_2364_375# 0.026339f
C8551 _408_/a_728_93# _095_ 0.040366f
C8552 mask\[2\] FILLER_0_16_154/a_932_472# 0.021665f
C8553 calibrate FILLER_0_8_156/a_36_472# 0.001283f
C8554 _122_ FILLER_0_8_156/a_572_375# 0.002572f
C8555 FILLER_0_13_142/a_484_472# _043_ 0.011974f
C8556 _431_/a_2665_112# FILLER_0_16_154/a_36_472# 0.007491f
C8557 _411_/a_2248_156# cal_itt\[0\] 0.006897f
C8558 _053_ _385_/a_36_68# 0.018437f
C8559 net29 _417_/a_2665_112# 0.002977f
C8560 _376_/a_36_160# FILLER_0_5_72/a_1380_472# 0.035111f
C8561 _081_ net47 1.302193f
C8562 net58 FILLER_0_9_282/a_124_375# 0.021949f
C8563 _186_ cal_count\[2\] 0.001605f
C8564 _099_ vss 0.255039f
C8565 FILLER_0_18_76/a_484_472# net71 0.004649f
C8566 net64 _100_ 0.001674f
C8567 FILLER_0_5_109/a_572_375# vss 0.055343f
C8568 FILLER_0_17_104/a_36_472# _438_/a_2248_156# 0.001731f
C8569 ctlp[1] FILLER_0_24_274/a_484_472# 0.001875f
C8570 net58 cal_itt\[2\] 0.003431f
C8571 FILLER_0_6_90/a_484_472# vss 0.00243f
C8572 _086_ _072_ 0.220767f
C8573 _100_ mask\[1\] 0.002229f
C8574 _428_/a_1308_423# vdd 0.004352f
C8575 net35 _436_/a_2560_156# 0.003198f
C8576 _101_ _005_ 0.003946f
C8577 _130_ _016_ 0.114514f
C8578 _004_ net64 0.001495f
C8579 mask\[7\] _433_/a_36_151# 0.001832f
C8580 trim_mask\[4\] _370_/a_1152_472# 0.001449f
C8581 _105_ _098_ 0.055065f
C8582 net58 net1 0.626432f
C8583 net52 FILLER_0_2_111/a_1380_472# 0.050754f
C8584 _372_/a_3126_472# _068_ 0.005304f
C8585 _004_ mask\[1\] 0.052788f
C8586 net62 FILLER_0_11_282/a_36_472# 0.00149f
C8587 _077_ _410_/a_36_68# 0.020334f
C8588 result[8] FILLER_0_24_274/a_124_375# 0.00726f
C8589 _061_ FILLER_0_8_156/a_572_375# 0.023346f
C8590 _119_ _072_ 0.189217f
C8591 _043_ _113_ 0.048005f
C8592 _132_ _022_ 0.001404f
C8593 net37 FILLER_0_6_231/a_572_375# 0.001989f
C8594 FILLER_0_15_72/a_124_375# vdd 0.020511f
C8595 _093_ net31 0.274432f
C8596 fanout63/a_36_160# vdd 0.020165f
C8597 FILLER_0_17_72/a_1380_472# _131_ 0.006873f
C8598 net58 _412_/a_36_151# 0.010226f
C8599 net75 _416_/a_2665_112# 0.001785f
C8600 output43/a_224_472# net17 0.083607f
C8601 net69 _031_ 0.450281f
C8602 FILLER_0_22_177/a_124_375# _434_/a_1308_423# 0.001064f
C8603 net33 _108_ 0.001901f
C8604 net50 net17 0.010654f
C8605 _425_/a_1000_472# net19 0.020388f
C8606 net62 FILLER_0_14_235/a_36_472# 0.00534f
C8607 _443_/a_1308_423# vdd 0.00203f
C8608 _443_/a_448_472# vss 0.030448f
C8609 FILLER_0_14_99/a_124_375# _451_/a_1040_527# 0.010005f
C8610 output36/a_224_472# output29/a_224_472# 0.007726f
C8611 _093_ FILLER_0_21_60/a_572_375# 0.011177f
C8612 FILLER_0_9_223/a_484_472# _055_ 0.026026f
C8613 FILLER_0_13_206/a_36_472# net79 0.00402f
C8614 _053_ vdd 1.467835f
C8615 _327_/a_36_472# _114_ 0.019746f
C8616 output34/a_224_472# _106_ 0.01606f
C8617 _142_ _020_ 0.010094f
C8618 FILLER_0_5_72/a_484_472# _440_/a_36_151# 0.001723f
C8619 result[8] _107_ 0.041984f
C8620 _413_/a_2665_112# vss 0.012213f
C8621 fanout62/a_36_160# net18 0.008106f
C8622 net19 _420_/a_36_151# 0.016882f
C8623 _036_ FILLER_0_3_54/a_124_375# 0.010221f
C8624 _274_/a_36_68# net4 0.037848f
C8625 net80 FILLER_0_19_171/a_124_375# 0.024758f
C8626 FILLER_0_1_212/a_124_375# vdd 0.020159f
C8627 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_124_375# 0.012001f
C8628 _126_ _124_ 0.012466f
C8629 _053_ FILLER_0_6_177/a_572_375# 0.01663f
C8630 net54 _140_ 1.37516f
C8631 _308_/a_1084_68# _115_ 0.001451f
C8632 _415_/a_36_151# net18 0.015992f
C8633 net16 FILLER_0_18_37/a_572_375# 0.03477f
C8634 ctln[4] _000_ 0.002823f
C8635 net55 FILLER_0_21_28/a_2724_472# 0.049771f
C8636 _397_/a_36_472# vdd 0.094023f
C8637 mask\[3\] _294_/a_224_472# 0.00233f
C8638 _320_/a_1120_472# state\[1\] 0.001998f
C8639 FILLER_0_2_177/a_572_375# vss 0.008507f
C8640 FILLER_0_2_177/a_36_472# vdd 0.110255f
C8641 mask\[0\] _137_ 0.009052f
C8642 output9/a_224_472# net2 0.003405f
C8643 _096_ _085_ 0.0099f
C8644 FILLER_0_18_171/a_36_472# net80 0.041571f
C8645 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1380_472# 0.026657f
C8646 net16 _446_/a_2665_112# 0.045966f
C8647 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001597f
C8648 FILLER_0_17_218/a_36_472# vss 0.006061f
C8649 FILLER_0_17_218/a_484_472# vdd 0.004777f
C8650 FILLER_0_18_2/a_1828_472# net55 0.011802f
C8651 FILLER_0_5_88/a_36_472# vdd 0.090268f
C8652 FILLER_0_5_88/a_124_375# vss 0.015423f
C8653 net71 FILLER_0_22_107/a_36_472# 0.034505f
C8654 output29/a_224_472# vdd 0.103437f
C8655 FILLER_0_5_206/a_124_375# net59 0.008027f
C8656 ctlp[4] net22 0.257841f
C8657 net74 _370_/a_124_24# 0.083426f
C8658 ctlp[1] _419_/a_36_151# 0.015335f
C8659 _086_ _132_ 0.014693f
C8660 trim[4] _054_ 0.005511f
C8661 output28/a_224_472# FILLER_0_11_282/a_124_375# 0.002977f
C8662 _093_ FILLER_0_17_142/a_124_375# 0.009328f
C8663 _441_/a_36_151# _160_ 0.030777f
C8664 _360_/a_36_160# _133_ 0.001878f
C8665 net54 FILLER_0_21_150/a_36_472# 0.005439f
C8666 _430_/a_2665_112# vdd 0.021353f
C8667 _412_/a_448_472# output9/a_224_472# 0.001025f
C8668 FILLER_0_21_286/a_572_375# vss 0.031895f
C8669 FILLER_0_21_286/a_36_472# vdd 0.008714f
C8670 net76 FILLER_0_5_198/a_36_472# 0.003987f
C8671 FILLER_0_21_28/a_2276_472# _423_/a_36_151# 0.013806f
C8672 _421_/a_1308_423# net19 0.055838f
C8673 _152_ _059_ 0.038141f
C8674 output45/a_224_472# trimb[3] 0.076387f
C8675 net69 _371_/a_36_113# 0.016091f
C8676 result[7] FILLER_0_24_274/a_1020_375# 0.006125f
C8677 FILLER_0_15_212/a_124_375# vss 0.005813f
C8678 FILLER_0_15_212/a_572_375# vdd -0.014642f
C8679 output9/a_224_472# cal 0.011495f
C8680 FILLER_0_5_164/a_124_375# _386_/a_848_380# 0.014613f
C8681 _394_/a_1936_472# vss 0.006085f
C8682 FILLER_0_4_144/a_572_375# net57 0.001254f
C8683 _163_ net14 0.040169f
C8684 FILLER_0_16_107/a_124_375# _131_ 0.016011f
C8685 _426_/a_36_151# net19 0.04851f
C8686 _131_ FILLER_0_16_115/a_124_375# 0.016715f
C8687 FILLER_0_2_93/a_36_472# trim_mask\[3\] 0.003417f
C8688 FILLER_0_9_28/a_3172_472# _077_ 0.011059f
C8689 FILLER_0_7_72/a_572_375# FILLER_0_6_47/a_3260_375# 0.026339f
C8690 FILLER_0_5_164/a_36_472# _385_/a_36_68# 0.001674f
C8691 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_124_375# 0.012222f
C8692 _414_/a_448_472# net22 0.047364f
C8693 FILLER_0_10_28/a_124_375# vdd 0.039012f
C8694 net16 FILLER_0_8_24/a_572_375# 0.002225f
C8695 _115_ net14 0.037635f
C8696 net38 net49 0.117427f
C8697 net70 net53 1.170795f
C8698 _119_ FILLER_0_8_127/a_36_472# 0.053962f
C8699 FILLER_0_15_142/a_572_375# net53 0.021481f
C8700 _093_ FILLER_0_17_161/a_36_472# 0.006224f
C8701 net16 net26 0.273031f
C8702 output39/a_224_472# _034_ 0.002236f
C8703 net44 vss 0.477283f
C8704 FILLER_0_7_72/a_2276_472# _439_/a_2665_112# 0.001167f
C8705 net34 FILLER_0_22_177/a_1468_375# 0.006974f
C8706 _420_/a_36_151# _009_ 0.018171f
C8707 _093_ _424_/a_2665_112# 0.001854f
C8708 _171_ vss 0.004501f
C8709 _016_ _428_/a_2248_156# 0.048889f
C8710 net20 FILLER_0_8_239/a_36_472# 0.004483f
C8711 _098_ _047_ 0.062495f
C8712 net82 _163_ 0.00269f
C8713 _027_ mask\[9\] 0.050723f
C8714 _288_/a_224_472# _102_ 0.002528f
C8715 net80 _434_/a_1308_423# 0.006837f
C8716 FILLER_0_7_72/a_2812_375# net14 0.025092f
C8717 FILLER_0_4_107/a_932_472# _158_ 0.029116f
C8718 mask\[4\] FILLER_0_18_177/a_572_375# 0.015941f
C8719 FILLER_0_5_54/a_932_472# _440_/a_36_151# 0.001723f
C8720 FILLER_0_11_142/a_36_472# _120_ 0.040786f
C8721 output45/a_224_472# ctlp[0] 0.007867f
C8722 net32 _420_/a_2665_112# 0.002753f
C8723 FILLER_0_15_116/a_484_472# _095_ 0.001069f
C8724 net54 _149_ 0.212511f
C8725 net50 _441_/a_448_472# 0.074088f
C8726 FILLER_0_13_212/a_572_375# net79 0.009626f
C8727 ctlp[2] vdd 0.617599f
C8728 FILLER_0_12_136/a_572_375# FILLER_0_13_142/a_36_472# 0.001684f
C8729 FILLER_0_16_89/a_572_375# _451_/a_448_472# 0.001597f
C8730 _131_ _427_/a_36_151# 0.0012f
C8731 _096_ _320_/a_224_472# 0.001285f
C8732 _238_/a_67_603# net50 0.002229f
C8733 mask\[4\] _348_/a_49_472# 0.001241f
C8734 net52 _440_/a_2665_112# 0.005084f
C8735 _028_ vdd 0.626868f
C8736 net52 _439_/a_1308_423# 0.033366f
C8737 net50 _439_/a_36_151# 0.009774f
C8738 FILLER_0_4_197/a_124_375# net21 0.018398f
C8739 FILLER_0_17_104/a_572_375# vdd 0.03661f
C8740 ctln[3] vdd 0.167569f
C8741 fanout82/a_36_113# net37 0.046126f
C8742 _425_/a_448_472# net37 0.002755f
C8743 _077_ FILLER_0_9_105/a_484_472# 0.002951f
C8744 _176_ vss 0.761803f
C8745 FILLER_0_5_164/a_36_472# vdd 0.004144f
C8746 FILLER_0_5_164/a_572_375# vss 0.055055f
C8747 net55 FILLER_0_19_28/a_484_472# 0.001426f
C8748 _239_/a_36_160# vss 0.001596f
C8749 _114_ _055_ 0.071738f
C8750 net45 net26 0.002978f
C8751 _321_/a_786_69# net23 0.001073f
C8752 _306_/a_36_68# vss 0.008326f
C8753 _132_ net53 0.035348f
C8754 net34 net19 0.039959f
C8755 net47 _450_/a_2225_156# 0.057106f
C8756 cal_count\[3\] _135_ 0.039115f
C8757 _068_ _261_/a_36_160# 0.008557f
C8758 _070_ _059_ 0.041498f
C8759 _131_ _180_ 0.016104f
C8760 _031_ FILLER_0_2_111/a_572_375# 0.023633f
C8761 net69 FILLER_0_2_111/a_1468_375# 0.021524f
C8762 net52 FILLER_0_6_47/a_2724_472# 0.011079f
C8763 net81 mask\[0\] 0.320022f
C8764 net18 FILLER_0_13_290/a_124_375# 0.007717f
C8765 net34 mask\[6\] 0.231853f
C8766 _128_ _121_ 0.051501f
C8767 _251_/a_1130_472# vss 0.001211f
C8768 FILLER_0_10_78/a_932_472# net52 0.00207f
C8769 _086_ state\[1\] 0.043298f
C8770 net55 _041_ 0.972122f
C8771 _431_/a_448_472# _131_ 0.006194f
C8772 FILLER_0_10_78/a_1380_472# _120_ 0.003228f
C8773 _274_/a_36_68# net79 0.009814f
C8774 _053_ FILLER_0_6_47/a_3172_472# 0.001777f
C8775 mask\[3\] FILLER_0_16_241/a_124_375# 0.006824f
C8776 _036_ vss 0.161195f
C8777 FILLER_0_18_107/a_1468_375# net71 0.001292f
C8778 _131_ _451_/a_2225_156# 0.008232f
C8779 mask\[0\] _060_ 0.002039f
C8780 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_1020_375# 0.001597f
C8781 _144_ _433_/a_1308_423# 0.027969f
C8782 _428_/a_2665_112# _427_/a_36_151# 0.028591f
C8783 _445_/a_2560_156# vdd 0.002586f
C8784 _445_/a_2665_112# vss 0.004455f
C8785 FILLER_0_17_200/a_36_472# vdd 0.001039f
C8786 FILLER_0_14_91/a_36_472# _136_ 0.008573f
C8787 _163_ FILLER_0_5_136/a_124_375# 0.009765f
C8788 trim_mask\[0\] vdd 0.154098f
C8789 output33/a_224_472# net19 0.12997f
C8790 _233_/a_36_160# net49 0.035342f
C8791 output47/a_224_472# net47 0.023797f
C8792 input5/a_36_113# rstn 0.019149f
C8793 FILLER_0_11_142/a_572_375# _121_ 0.003107f
C8794 _414_/a_2248_156# _053_ 0.013478f
C8795 _421_/a_1000_472# _010_ 0.01379f
C8796 _181_ _182_ 0.02735f
C8797 FILLER_0_19_55/a_36_472# net55 0.062683f
C8798 mask\[5\] _140_ 0.103728f
C8799 _104_ _422_/a_2560_156# 0.003223f
C8800 FILLER_0_18_2/a_1468_375# _452_/a_448_472# 0.001597f
C8801 net75 ctln[3] 0.066513f
C8802 _322_/a_692_472# _118_ 0.002849f
C8803 net16 FILLER_0_17_38/a_36_472# 0.014381f
C8804 FILLER_0_15_150/a_36_472# net56 0.011741f
C8805 _221_/a_36_160# vdd 0.073414f
C8806 FILLER_0_13_65/a_124_375# vss 0.030194f
C8807 FILLER_0_14_181/a_36_472# vdd 0.027265f
C8808 FILLER_0_14_181/a_124_375# vss 0.009291f
C8809 _253_/a_1528_68# cal_itt\[1\] 0.002251f
C8810 _072_ _161_ 0.048567f
C8811 _425_/a_2248_156# vdd 0.010067f
C8812 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_36_472# 0.086635f
C8813 net20 FILLER_0_12_220/a_484_472# 0.001758f
C8814 _430_/a_36_151# _092_ 0.002363f
C8815 net17 _054_ 0.034759f
C8816 _017_ FILLER_0_14_107/a_1020_375# 0.001363f
C8817 net70 FILLER_0_14_107/a_36_472# 0.054561f
C8818 FILLER_0_12_2/a_124_375# _450_/a_36_151# 0.001543f
C8819 _110_ _423_/a_2665_112# 0.001668f
C8820 FILLER_0_24_290/a_124_375# FILLER_0_24_274/a_1468_375# 0.012001f
C8821 _122_ FILLER_0_6_231/a_572_375# 0.016091f
C8822 _050_ _436_/a_2248_156# 0.023725f
C8823 _449_/a_1308_423# _453_/a_2665_112# 0.001066f
C8824 FILLER_0_16_57/a_932_472# _131_ 0.007885f
C8825 net78 _094_ 0.050187f
C8826 FILLER_0_17_133/a_36_472# vdd 0.097394f
C8827 FILLER_0_17_133/a_124_375# vss 0.015434f
C8828 _420_/a_1308_423# vdd 0.00284f
C8829 _420_/a_448_472# vss 0.007371f
C8830 _321_/a_170_472# _120_ 0.040613f
C8831 _063_ _167_ 0.002201f
C8832 net70 _451_/a_36_151# 0.04524f
C8833 cal_itt\[1\] _082_ 0.921465f
C8834 _320_/a_1120_472# vdd 0.001676f
C8835 net3 FILLER_0_15_2/a_572_375# 0.004377f
C8836 net34 _009_ 0.325819f
C8837 _098_ FILLER_0_15_180/a_36_472# 0.101593f
C8838 net20 _419_/a_1308_423# 0.022245f
C8839 net33 _435_/a_2665_112# 0.005831f
C8840 _013_ FILLER_0_18_37/a_1020_375# 0.023067f
C8841 net19 _419_/a_448_472# 0.037199f
C8842 net80 _136_ 0.034194f
C8843 net44 input3/a_36_113# 0.016865f
C8844 _093_ FILLER_0_18_139/a_1020_375# 0.003529f
C8845 mask\[9\] _438_/a_796_472# 0.004751f
C8846 _236_/a_36_160# output39/a_224_472# 0.042231f
C8847 _395_/a_36_488# _116_ 0.033784f
C8848 net80 net21 0.016911f
C8849 _079_ _074_ 0.025058f
C8850 FILLER_0_3_172/a_1916_375# net22 0.00941f
C8851 _114_ _058_ 0.013316f
C8852 _434_/a_36_151# vss 0.006401f
C8853 _434_/a_448_472# vdd 0.020387f
C8854 _008_ net30 1.112351f
C8855 FILLER_0_13_142/a_572_375# vdd 0.017472f
C8856 FILLER_0_13_142/a_124_375# vss 0.009543f
C8857 net76 net18 0.002264f
C8858 _132_ FILLER_0_11_109/a_36_472# 0.005748f
C8859 result[4] net77 0.003336f
C8860 FILLER_0_9_28/a_2724_472# _077_ 0.006001f
C8861 _429_/a_36_151# _018_ 0.118135f
C8862 result[5] _094_ 0.065897f
C8863 _183_ vss 0.009822f
C8864 _057_ net57 0.873864f
C8865 _081_ _385_/a_36_68# 0.006303f
C8866 mask\[3\] _046_ 0.018595f
C8867 _082_ vss 0.053349f
C8868 _073_ net82 0.028504f
C8869 net79 _416_/a_2248_156# 0.026136f
C8870 output43/a_224_472# trimb[3] 0.070044f
C8871 FILLER_0_8_247/a_36_472# vss 0.003706f
C8872 FILLER_0_8_247/a_484_472# vdd 0.005485f
C8873 FILLER_0_14_91/a_484_472# net53 0.00544f
C8874 _421_/a_1000_472# vdd 0.006281f
C8875 _432_/a_2560_156# net63 0.00227f
C8876 net53 state\[1\] 0.00554f
C8877 fanout77/a_36_113# vss 0.004099f
C8878 _132_ FILLER_0_14_107/a_36_472# 0.002187f
C8879 cal_count\[3\] _408_/a_1336_472# 0.010351f
C8880 net23 FILLER_0_22_128/a_2724_472# 0.054521f
C8881 FILLER_0_4_197/a_1020_375# vss 0.001981f
C8882 _116_ _228_/a_36_68# 0.013091f
C8883 FILLER_0_4_123/a_36_472# _160_ 0.050308f
C8884 mask\[0\] _095_ 0.006711f
C8885 fanout81/a_36_160# vdd 0.095319f
C8886 _412_/a_2560_156# en 0.049213f
C8887 net50 FILLER_0_7_59/a_124_375# 0.002292f
C8888 _028_ _439_/a_796_472# 0.013039f
C8889 net63 FILLER_0_17_218/a_572_375# 0.006355f
C8890 FILLER_0_11_101/a_572_375# _134_ 0.0024f
C8891 _062_ _113_ 0.020368f
C8892 net63 _435_/a_2560_156# 0.023868f
C8893 _265_/a_244_68# cal_itt\[1\] 0.024108f
C8894 _426_/a_1308_423# vdd 0.008509f
C8895 net79 _099_ 0.010543f
C8896 _446_/a_1000_472# net40 0.0368f
C8897 _178_ vdd 0.440802f
C8898 _086_ FILLER_0_5_181/a_124_375# 0.006872f
C8899 net61 output19/a_224_472# 0.077658f
C8900 FILLER_0_11_101/a_124_375# vdd 0.024363f
C8901 net75 _253_/a_1732_68# 0.001047f
C8902 _129_ cal_count\[3\] 0.005967f
C8903 _132_ _451_/a_36_151# 0.007777f
C8904 _441_/a_2665_112# net49 0.062459f
C8905 _053_ FILLER_0_7_59/a_484_472# 0.013665f
C8906 _028_ FILLER_0_6_47/a_3172_472# 0.015585f
C8907 trim_val\[3\] _441_/a_1308_423# 0.001312f
C8908 trim_mask\[2\] _036_ 0.466145f
C8909 _085_ _055_ 0.240451f
C8910 vdd _022_ 0.082842f
C8911 net71 _437_/a_36_151# 0.055761f
C8912 _064_ _445_/a_1000_472# 0.015908f
C8913 _431_/a_36_151# net73 0.015086f
C8914 _447_/a_1000_472# net68 0.006223f
C8915 _447_/a_1308_423# _036_ 0.003079f
C8916 _116_ calibrate 0.018482f
C8917 cal_itt\[3\] vdd 0.571239f
C8918 _247_/a_36_160# net21 0.002254f
C8919 fanout80/a_36_113# _139_ 0.009968f
C8920 FILLER_0_16_154/a_932_472# vss 0.001652f
C8921 FILLER_0_16_154/a_1380_472# vdd 0.001901f
C8922 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3260_375# 0.001597f
C8923 FILLER_0_3_172/a_2812_375# net21 0.015743f
C8924 FILLER_0_8_239/a_36_472# vss 0.003115f
C8925 _265_/a_244_68# vss 0.009604f
C8926 _408_/a_1336_472# net40 0.020063f
C8927 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_36_472# 0.002296f
C8928 _257_/a_244_68# _053_ 0.001138f
C8929 ctln[2] net19 0.073057f
C8930 _081_ vdd 0.729534f
C8931 net75 FILLER_0_8_247/a_484_472# 0.003007f
C8932 fanout75/a_36_113# net76 0.040306f
C8933 net31 _094_ 0.203395f
C8934 sample fanout64/a_36_160# 0.007266f
C8935 _112_ vss 0.145781f
C8936 _118_ _062_ 0.029651f
C8937 cal_itt\[3\] FILLER_0_6_177/a_572_375# 0.00225f
C8938 _189_/a_67_603# _429_/a_2665_112# 0.015187f
C8939 FILLER_0_7_104/a_932_472# vdd 0.020291f
C8940 _070_ _247_/a_36_160# 0.0169f
C8941 net32 _419_/a_2560_156# 0.029586f
C8942 net36 _040_ 0.429029f
C8943 output48/a_224_472# valid 0.046397f
C8944 fanout64/a_36_160# vss 0.007097f
C8945 FILLER_0_12_136/a_1020_375# state\[2\] 0.001952f
C8946 FILLER_0_14_99/a_124_375# net14 0.04852f
C8947 net73 FILLER_0_18_107/a_1380_472# 0.039646f
C8948 _053_ FILLER_0_7_146/a_124_375# 0.005844f
C8949 net82 _425_/a_36_151# 0.002959f
C8950 FILLER_0_15_150/a_36_472# _095_ 0.001526f
C8951 net75 _426_/a_1308_423# 0.002552f
C8952 net68 _381_/a_36_472# 0.003421f
C8953 _081_ FILLER_0_6_177/a_572_375# 0.007285f
C8954 net54 net14 0.121719f
C8955 _072_ _071_ 0.296543f
C8956 FILLER_0_18_107/a_3260_375# vss 0.056926f
C8957 FILLER_0_18_107/a_36_472# vdd 0.116746f
C8958 output15/a_224_472# vss 0.067969f
C8959 FILLER_0_19_195/a_124_375# _202_/a_36_160# 0.005489f
C8960 FILLER_0_20_2/a_124_375# net43 0.001563f
C8961 _431_/a_2560_156# vss 0.004767f
C8962 net40 _034_ 0.04333f
C8963 valid net5 0.044555f
C8964 net52 FILLER_0_9_72/a_932_472# 0.008749f
C8965 net23 _208_/a_36_160# 0.112626f
C8966 _115_ _131_ 0.410424f
C8967 result[8] net32 0.024881f
C8968 FILLER_0_14_107/a_572_375# _451_/a_36_151# 0.02627f
C8969 net27 FILLER_0_12_236/a_572_375# 0.083731f
C8970 _178_ net72 0.007093f
C8971 FILLER_0_18_139/a_1468_375# _145_ 0.002318f
C8972 _433_/a_2560_156# _145_ 0.007651f
C8973 FILLER_0_18_37/a_1380_472# vdd 0.004422f
C8974 FILLER_0_16_241/a_36_472# net36 0.001988f
C8975 FILLER_0_16_89/a_36_472# vss 0.001289f
C8976 _270_/a_36_472# vdd 0.09815f
C8977 cal_itt\[2\] net82 0.663246f
C8978 FILLER_0_8_138/a_124_375# _076_ 0.031436f
C8979 FILLER_0_5_109/a_36_472# net47 0.005565f
C8980 _421_/a_36_151# net77 0.028951f
C8981 _030_ _153_ 0.026157f
C8982 FILLER_0_9_28/a_1916_375# _453_/a_36_151# 0.001543f
C8983 _010_ _419_/a_796_472# 0.001613f
C8984 ctlp[1] _010_ 0.002794f
C8985 net82 net1 0.029512f
C8986 _086_ vdd 1.212255f
C8987 FILLER_0_24_274/a_1380_472# vss 0.005744f
C8988 _425_/a_448_472# _122_ 0.002863f
C8989 _425_/a_1308_423# calibrate 0.022697f
C8990 fanout82/a_36_113# _122_ 0.007118f
C8991 net39 _054_ 0.049797f
C8992 mask\[0\] net64 0.45093f
C8993 _065_ net69 0.051511f
C8994 ctln[7] _442_/a_2665_112# 0.01075f
C8995 _035_ net17 0.021052f
C8996 _089_ vdd 0.087336f
C8997 FILLER_0_16_57/a_1468_375# _175_ 0.001654f
C8998 net10 _411_/a_2248_156# 0.002419f
C8999 mask\[0\] mask\[1\] 0.01742f
C9000 net75 _081_ 0.060976f
C9001 net20 net48 0.035427f
C9002 _011_ _422_/a_796_472# 0.009261f
C9003 ctln[5] net12 0.41364f
C9004 _416_/a_36_151# output30/a_224_472# 0.012025f
C9005 _411_/a_1000_472# ctln[3] 0.00283f
C9006 _132_ _127_ 0.112364f
C9007 FILLER_0_5_128/a_484_472# _160_ 0.003335f
C9008 _412_/a_36_151# net82 0.064296f
C9009 _119_ vdd 0.38257f
C9010 FILLER_0_4_197/a_484_472# vdd 0.002749f
C9011 _086_ FILLER_0_6_177/a_572_375# 0.012909f
C9012 _091_ FILLER_0_15_180/a_484_472# 0.001757f
C9013 _000_ FILLER_0_3_221/a_932_472# 0.008308f
C9014 FILLER_0_24_96/a_36_472# vss 0.003218f
C9015 net79 FILLER_0_21_286/a_572_375# 0.001476f
C9016 _021_ net80 0.254353f
C9017 cal_count\[2\] _179_ 0.404284f
C9018 trim_mask\[4\] _159_ 0.049552f
C9019 net38 net47 0.352245f
C9020 net28 _094_ 0.007842f
C9021 net16 _402_/a_728_93# 0.040925f
C9022 FILLER_0_4_185/a_124_375# FILLER_0_4_177/a_572_375# 0.012001f
C9023 _006_ net30 0.284414f
C9024 mask\[4\] _143_ 0.352305f
C9025 _072_ FILLER_0_10_214/a_36_472# 0.015199f
C9026 _430_/a_36_151# vdd 0.112575f
C9027 output14/a_224_472# FILLER_0_0_130/a_36_472# 0.023414f
C9028 net57 cal_count\[3\] 0.02848f
C9029 FILLER_0_7_72/a_2276_472# net50 0.030391f
C9030 _068_ _062_ 0.089152f
C9031 _070_ _134_ 0.087767f
C9032 net47 _386_/a_692_472# 0.003299f
C9033 FILLER_0_22_177/a_1020_375# mask\[6\] 0.002657f
C9034 _155_ FILLER_0_8_107/a_36_472# 0.002068f
C9035 _321_/a_2590_472# _129_ 0.005391f
C9036 output10/a_224_472# ctln[2] 0.024524f
C9037 _161_ state\[1\] 0.002512f
C9038 output26/a_224_472# FILLER_0_23_44/a_1380_472# 0.0323f
C9039 _005_ vdd 0.506158f
C9040 net62 _101_ 0.023932f
C9041 net18 _416_/a_1000_472# 0.046085f
C9042 _431_/a_448_472# _137_ 0.008493f
C9043 _449_/a_1308_423# vdd 0.002584f
C9044 _449_/a_448_472# vss 0.032274f
C9045 _210_/a_67_603# net23 0.005398f
C9046 net50 FILLER_0_6_90/a_124_375# 0.041764f
C9047 _395_/a_1492_488# _121_ 0.002537f
C9048 _412_/a_1204_472# net65 0.001629f
C9049 FILLER_0_12_220/a_484_472# vss 0.006724f
C9050 FILLER_0_12_220/a_932_472# vdd 0.003359f
C9051 _431_/a_796_472# net70 0.001754f
C9052 _052_ mask\[9\] 0.007224f
C9053 net55 FILLER_0_18_37/a_36_472# 0.006084f
C9054 FILLER_0_4_107/a_1380_472# _160_ 0.020979f
C9055 _322_/a_848_380# net74 0.00168f
C9056 _450_/a_36_151# output6/a_224_472# 0.134892f
C9057 _414_/a_2665_112# vss 0.010021f
C9058 net35 _434_/a_2665_112# 0.024254f
C9059 FILLER_0_17_72/a_1916_375# vdd 0.002595f
C9060 FILLER_0_17_72/a_1468_375# vss 0.003461f
C9061 FILLER_0_5_109/a_484_472# _363_/a_36_68# 0.001709f
C9062 _308_/a_124_24# _439_/a_2665_112# 0.002245f
C9063 _105_ _420_/a_2665_112# 0.001159f
C9064 _132_ FILLER_0_19_111/a_484_472# 0.004619f
C9065 _004_ FILLER_0_10_247/a_36_472# 0.001551f
C9066 net23 FILLER_0_16_154/a_36_472# 0.035678f
C9067 net20 net19 0.384932f
C9068 _053_ FILLER_0_6_90/a_484_472# 0.011443f
C9069 output29/a_224_472# _416_/a_2248_156# 0.024448f
C9070 result[2] _416_/a_448_472# 0.003015f
C9071 FILLER_0_8_247/a_572_375# calibrate 0.008498f
C9072 fanout50/a_36_160# net52 0.037383f
C9073 _401_/a_36_68# FILLER_0_15_59/a_36_472# 0.019798f
C9074 net35 _213_/a_255_603# 0.001597f
C9075 _301_/a_36_472# _051_ 0.001277f
C9076 FILLER_0_22_86/a_572_375# vdd 0.017472f
C9077 FILLER_0_22_86/a_124_375# vss 0.00285f
C9078 net4 _082_ 0.004529f
C9079 FILLER_0_4_197/a_1468_375# vss 0.057762f
C9080 net38 _450_/a_836_156# 0.0039f
C9081 _116_ FILLER_0_12_196/a_36_472# 0.010951f
C9082 FILLER_0_9_223/a_572_375# _076_ 0.034523f
C9083 _415_/a_2665_112# net64 0.074373f
C9084 net52 _443_/a_36_151# 0.020518f
C9085 ctlp[1] vdd 0.942436f
C9086 _303_/a_36_472# _012_ 0.001735f
C9087 net57 _169_ 0.033365f
C9088 _140_ _348_/a_49_472# 0.023816f
C9089 en_co_clk _390_/a_36_68# 0.086301f
C9090 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_36_472# 0.026657f
C9091 net80 FILLER_0_22_177/a_484_472# 0.005297f
C9092 FILLER_0_16_107/a_36_472# _093_ 0.001526f
C9093 FILLER_0_15_59/a_484_472# vss 0.007866f
C9094 mask\[5\] FILLER_0_19_155/a_484_472# 0.043011f
C9095 _412_/a_1204_472# net59 0.001824f
C9096 _055_ _310_/a_49_472# 0.00384f
C9097 net18 FILLER_0_11_282/a_36_472# 0.048657f
C9098 _326_/a_36_160# _134_ 0.003299f
C9099 FILLER_0_9_142/a_124_375# vdd 0.015952f
C9100 FILLER_0_17_72/a_3172_472# _136_ 0.002925f
C9101 _453_/a_448_472# _042_ 0.053209f
C9102 _453_/a_36_151# net51 0.012537f
C9103 _053_ _414_/a_796_472# 0.008213f
C9104 fanout75/a_36_113# _083_ 0.002133f
C9105 net54 _098_ 0.116416f
C9106 net74 _371_/a_36_113# 0.027966f
C9107 fanout69/a_36_113# _159_ 0.005623f
C9108 FILLER_0_4_185/a_124_375# net22 0.004776f
C9109 _178_ cal_count\[0\] 0.011488f
C9110 net53 vdd 0.78288f
C9111 _017_ vss 0.022624f
C9112 _135_ _120_ 0.017522f
C9113 net34 FILLER_0_22_128/a_1468_375# 0.003214f
C9114 net15 _441_/a_1308_423# 0.009697f
C9115 _072_ _246_/a_36_68# 0.064797f
C9116 _093_ _027_ 0.047164f
C9117 _016_ _118_ 0.001549f
C9118 _431_/a_2665_112# vdd 0.015335f
C9119 FILLER_0_4_177/a_124_375# net76 0.003962f
C9120 FILLER_0_4_213/a_36_472# vdd 0.087733f
C9121 FILLER_0_4_213/a_572_375# vss 0.017689f
C9122 _064_ net67 0.006691f
C9123 _109_ _108_ 0.001806f
C9124 net54 _436_/a_2665_112# 0.042428f
C9125 net60 _094_ 0.579872f
C9126 net55 FILLER_0_17_72/a_572_375# 0.023585f
C9127 _446_/a_796_472# net66 0.002296f
C9128 net15 _439_/a_448_472# 0.038829f
C9129 net47 FILLER_0_5_148/a_572_375# 0.062581f
C9130 _233_/a_36_160# net47 0.054273f
C9131 _414_/a_2248_156# cal_itt\[3\] 0.032294f
C9132 net4 FILLER_0_8_239/a_36_472# 0.008503f
C9133 _032_ vss 0.02257f
C9134 net27 FILLER_0_9_290/a_124_375# 0.002657f
C9135 _250_/a_36_68# vss 0.005108f
C9136 net63 FILLER_0_17_200/a_572_375# 0.007512f
C9137 _112_ _316_/a_1084_68# 0.005773f
C9138 _236_/a_36_160# net40 0.035082f
C9139 net41 _181_ 0.043679f
C9140 net54 _433_/a_2248_156# 0.04755f
C9141 _077_ FILLER_0_10_94/a_484_472# 0.001548f
C9142 net54 FILLER_0_18_139/a_572_375# 0.00217f
C9143 _077_ _453_/a_1204_472# 0.011124f
C9144 fanout80/a_36_113# _098_ 0.011559f
C9145 _414_/a_2248_156# _081_ 0.002027f
C9146 _446_/a_1000_472# trim[3] 0.001257f
C9147 _431_/a_448_472# net56 0.001464f
C9148 FILLER_0_21_125/a_36_472# vdd 0.007233f
C9149 FILLER_0_21_125/a_572_375# vss 0.054783f
C9150 FILLER_0_11_78/a_124_375# vdd -0.011022f
C9151 FILLER_0_20_193/a_572_375# _098_ 0.078973f
C9152 FILLER_0_5_72/a_36_472# _029_ 0.007282f
C9153 FILLER_0_5_72/a_572_375# trim_mask\[1\] 0.010714f
C9154 net20 _009_ 0.026064f
C9155 net15 FILLER_0_6_47/a_2276_472# 0.049487f
C9156 FILLER_0_6_47/a_1468_375# vdd -0.014642f
C9157 _037_ net59 0.799647f
C9158 output16/a_224_472# vdd 0.006151f
C9159 cal_itt\[3\] _374_/a_36_68# 0.001569f
C9160 _321_/a_3126_472# _126_ 0.002939f
C9161 _321_/a_358_69# _069_ 0.001124f
C9162 _301_/a_36_472# vdd 0.013061f
C9163 FILLER_0_12_50/a_124_375# vdd 0.039185f
C9164 vdd _450_/a_2225_156# 0.020301f
C9165 net16 net17 0.034209f
C9166 _091_ FILLER_0_20_169/a_124_375# 0.003958f
C9167 FILLER_0_13_228/a_36_472# _043_ 0.02119f
C9168 _292_/a_36_160# net31 0.010041f
C9169 mask\[3\] FILLER_0_17_200/a_124_375# 0.01841f
C9170 FILLER_0_7_104/a_1020_375# _153_ 0.026997f
C9171 _317_/a_36_113# calibrate 0.011799f
C9172 fanout56/a_36_113# _136_ 0.002316f
C9173 cal_count\[3\] _453_/a_448_472# 0.001494f
C9174 _422_/a_448_472# _108_ 0.03293f
C9175 net58 _412_/a_2248_156# 0.010702f
C9176 FILLER_0_17_133/a_36_472# FILLER_0_19_134/a_124_375# 0.001188f
C9177 ctln[4] FILLER_0_1_204/a_36_472# 0.006408f
C9178 FILLER_0_18_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001684f
C9179 _115_ FILLER_0_10_107/a_124_375# 0.011098f
C9180 net55 net47 0.049398f
C9181 _098_ FILLER_0_16_154/a_572_375# 0.001791f
C9182 _370_/a_848_380# FILLER_0_5_136/a_36_472# 0.001177f
C9183 FILLER_0_9_60/a_484_472# vdd 0.005181f
C9184 FILLER_0_9_60/a_36_472# vss 0.001327f
C9185 _449_/a_36_151# FILLER_0_11_64/a_36_472# 0.046516f
C9186 _204_/a_67_603# vdd 0.039556f
C9187 _020_ vss 0.008954f
C9188 fanout72/a_36_113# vdd -0.002193f
C9189 _415_/a_796_472# net19 0.001468f
C9190 _114_ _172_ 0.045798f
C9191 net62 FILLER_0_15_290/a_124_375# 0.034614f
C9192 _412_/a_1000_472# net65 0.00929f
C9193 output12/a_224_472# net76 0.00803f
C9194 state\[1\] _071_ 0.196063f
C9195 net41 _446_/a_1308_423# 0.056251f
C9196 _412_/a_1308_423# net81 0.006961f
C9197 _110_ _437_/a_36_151# 0.00125f
C9198 net74 FILLER_0_2_111/a_1468_375# 0.003854f
C9199 FILLER_0_23_282/a_124_375# vdd -0.003896f
C9200 net42 _054_ 0.006314f
C9201 _028_ FILLER_0_6_90/a_484_472# 0.01566f
C9202 output47/a_224_472# vdd 0.028666f
C9203 FILLER_0_12_124/a_36_472# _428_/a_36_151# 0.001723f
C9204 FILLER_0_21_28/a_1828_472# _012_ 0.021162f
C9205 net74 _124_ 0.180235f
C9206 _072_ net23 0.006278f
C9207 _069_ net36 0.032818f
C9208 _178_ _407_/a_36_472# 0.001699f
C9209 _445_/a_448_472# _034_ 0.03826f
C9210 _433_/a_36_151# _022_ 0.017789f
C9211 trim_mask\[1\] _160_ 0.051511f
C9212 net27 FILLER_0_10_247/a_124_375# 0.015466f
C9213 FILLER_0_18_2/a_932_472# net38 0.020589f
C9214 FILLER_0_11_109/a_124_375# vss 0.006764f
C9215 FILLER_0_11_109/a_36_472# vdd 0.109453f
C9216 FILLER_0_12_136/a_36_472# _127_ 0.023927f
C9217 FILLER_0_16_57/a_124_375# FILLER_0_18_53/a_484_472# 0.001512f
C9218 _076_ _226_/a_1044_68# 0.0023f
C9219 _093_ FILLER_0_17_104/a_1380_472# 0.014431f
C9220 FILLER_0_2_93/a_572_375# vdd 0.022073f
C9221 net29 net36 0.370099f
C9222 net48 FILLER_0_7_233/a_36_472# 0.01015f
C9223 input5/a_36_113# net59 0.257143f
C9224 FILLER_0_12_124/a_36_472# _114_ 0.003953f
C9225 _086_ _374_/a_36_68# 0.009872f
C9226 _311_/a_66_473# net21 0.02018f
C9227 FILLER_0_11_135/a_36_472# vdd 0.091206f
C9228 FILLER_0_11_135/a_124_375# vss 0.02843f
C9229 net45 net17 0.192181f
C9230 _448_/a_1000_472# vdd 0.004267f
C9231 _412_/a_1000_472# net59 0.00147f
C9232 FILLER_0_14_107/a_36_472# vdd 0.114495f
C9233 net38 FILLER_0_20_2/a_36_472# 0.002204f
C9234 FILLER_0_14_107/a_1468_375# vss 0.055167f
C9235 net72 FILLER_0_12_50/a_124_375# 0.011077f
C9236 FILLER_0_15_142/a_572_375# net23 0.006327f
C9237 net23 net47 0.090948f
C9238 net48 vss 0.161385f
C9239 FILLER_0_22_177/a_1468_375# vss 0.028064f
C9240 FILLER_0_22_177/a_36_472# vdd 0.111906f
C9241 output44/a_224_472# _452_/a_448_472# 0.004683f
C9242 _119_ _374_/a_36_68# 0.001756f
C9243 net4 FILLER_0_12_220/a_484_472# 0.022264f
C9244 net34 net63 0.050865f
C9245 mask\[3\] fanout53/a_36_160# 0.001205f
C9246 _091_ _223_/a_36_160# 0.001976f
C9247 _423_/a_36_151# FILLER_0_23_44/a_1020_375# 0.059049f
C9248 _086_ _331_/a_448_472# 0.004356f
C9249 FILLER_0_3_221/a_36_472# vss 0.046345f
C9250 FILLER_0_3_221/a_484_472# vdd 0.002974f
C9251 FILLER_0_7_104/a_36_472# _058_ 0.006613f
C9252 net36 FILLER_0_15_212/a_36_472# 0.005396f
C9253 net16 FILLER_0_16_37/a_36_472# 0.015199f
C9254 _162_ vss 0.08357f
C9255 _161_ vdd 0.262564f
C9256 _427_/a_36_151# _095_ 0.029048f
C9257 net68 FILLER_0_5_54/a_124_375# 0.018458f
C9258 _399_/a_224_472# vdd 0.001593f
C9259 fanout72/a_36_113# net72 0.02315f
C9260 net19 cal_itt\[1\] 0.044717f
C9261 net41 _160_ 0.006523f
C9262 _059_ FILLER_0_5_148/a_36_472# 0.010977f
C9263 _129_ _120_ 0.017802f
C9264 _451_/a_36_151# vdd 0.088651f
C9265 FILLER_0_5_212/a_124_375# net37 0.005414f
C9266 FILLER_0_5_54/a_1020_375# trim_mask\[1\] 0.010745f
C9267 FILLER_0_9_223/a_36_472# _055_ 0.014713f
C9268 _093_ _438_/a_796_472# 0.001924f
C9269 net50 _030_ 0.073046f
C9270 _441_/a_36_151# _440_/a_36_151# 0.003983f
C9271 net61 output18/a_224_472# 0.059062f
C9272 mask\[0\] FILLER_0_12_236/a_36_472# 0.002801f
C9273 net35 FILLER_0_22_86/a_1380_472# 0.00813f
C9274 net52 _442_/a_2665_112# 0.031179f
C9275 _137_ FILLER_0_15_180/a_36_472# 0.004437f
C9276 _140_ _350_/a_49_472# 0.028997f
C9277 _413_/a_1204_472# _002_ 0.003057f
C9278 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_36_472# 0.009654f
C9279 FILLER_0_16_89/a_572_375# _040_ 0.004252f
C9280 _162_ FILLER_0_6_177/a_36_472# 0.001723f
C9281 _161_ FILLER_0_6_177/a_572_375# 0.004064f
C9282 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_124_375# 0.001597f
C9283 _285_/a_36_472# vdd 0.073338f
C9284 trim[4] FILLER_0_8_2/a_36_472# 0.019134f
C9285 _027_ FILLER_0_18_76/a_572_375# 0.08501f
C9286 _150_ FILLER_0_18_76/a_484_472# 0.003548f
C9287 _002_ net22 0.038848f
C9288 FILLER_0_15_150/a_124_375# net56 0.011873f
C9289 mask\[5\] _098_ 1.316993f
C9290 _205_/a_36_160# vss 0.003612f
C9291 net16 FILLER_0_12_28/a_124_375# 0.002225f
C9292 _069_ _116_ 0.390834f
C9293 _098_ FILLER_0_18_209/a_572_375# 0.001352f
C9294 net2 _001_ 0.081616f
C9295 _258_/a_36_160# _079_ 0.026618f
C9296 _095_ _180_ 0.013383f
C9297 FILLER_0_18_177/a_3260_375# vdd 0.003399f
C9298 net15 FILLER_0_7_59/a_572_375# 0.033245f
C9299 FILLER_0_21_206/a_36_472# _434_/a_2665_112# 0.00243f
C9300 net32 _103_ 0.038496f
C9301 _063_ _232_/a_67_603# 0.005404f
C9302 net19 vss 1.140787f
C9303 output8/a_224_472# net8 0.034396f
C9304 FILLER_0_9_28/a_932_472# net68 0.003603f
C9305 _076_ FILLER_0_8_156/a_36_472# 0.006989f
C9306 _068_ FILLER_0_8_156/a_572_375# 0.00185f
C9307 _013_ FILLER_0_18_53/a_36_472# 0.013138f
C9308 net16 _235_/a_67_603# 0.038585f
C9309 FILLER_0_7_59/a_36_472# trim_val\[0\] 0.003014f
C9310 FILLER_0_23_88/a_36_472# vdd 0.002576f
C9311 FILLER_0_23_88/a_124_375# vss 0.014165f
C9312 output16/a_224_472# _447_/a_448_472# 0.003175f
C9313 output13/a_224_472# net59 0.007733f
C9314 _412_/a_448_472# _001_ 0.01124f
C9315 output26/a_224_472# ctlp[9] 0.034572f
C9316 _095_ _451_/a_2225_156# 0.001102f
C9317 _440_/a_36_151# FILLER_0_6_47/a_1380_472# 0.001512f
C9318 mask\[6\] vss 0.348967f
C9319 _417_/a_2665_112# _006_ 0.023025f
C9320 _072_ _056_ 0.061377f
C9321 _173_ _186_ 0.002111f
C9322 _439_/a_36_151# FILLER_0_6_47/a_2812_375# 0.001512f
C9323 FILLER_0_1_266/a_124_375# FILLER_0_0_266/a_124_375# 0.05841f
C9324 net4 FILLER_0_4_213/a_572_375# 0.001015f
C9325 _105_ result[8] 0.011678f
C9326 input2/a_36_113# vss 0.055539f
C9327 _430_/a_36_151# _337_/a_49_472# 0.023882f
C9328 _189_/a_67_603# net27 0.008028f
C9329 FILLER_0_6_79/a_36_472# vss 0.008693f
C9330 FILLER_0_16_73/a_572_375# vss 0.030752f
C9331 _444_/a_2665_112# _164_ 0.015644f
C9332 _399_/a_224_472# net72 0.002538f
C9333 _088_ _260_/a_36_68# 0.003476f
C9334 _412_/a_448_472# output37/a_224_472# 0.001155f
C9335 net53 _427_/a_1204_472# 0.004293f
C9336 _444_/a_2248_156# net67 0.028782f
C9337 net16 FILLER_0_19_47/a_36_472# 0.009509f
C9338 _015_ FILLER_0_8_247/a_572_375# 0.00706f
C9339 _181_ cal_count\[2\] 0.375819f
C9340 FILLER_0_1_204/a_36_472# net21 0.076466f
C9341 FILLER_0_5_72/a_572_375# _164_ 0.005919f
C9342 _139_ _138_ 0.00256f
C9343 output38/a_224_472# net38 0.018882f
C9344 vdd _201_/a_67_603# 0.031337f
C9345 net35 _352_/a_49_472# 0.02594f
C9346 mask\[8\] _352_/a_257_69# 0.003259f
C9347 _114_ FILLER_0_13_142/a_1020_375# 0.001964f
C9348 FILLER_0_3_54/a_36_472# vss 0.002818f
C9349 FILLER_0_8_127/a_124_375# vdd 0.019587f
C9350 net16 _039_ 0.031852f
C9351 _095_ FILLER_0_13_72/a_36_472# 0.00819f
C9352 FILLER_0_18_2/a_2364_375# net17 0.048345f
C9353 _017_ _332_/a_36_472# 0.033837f
C9354 _008_ _418_/a_2665_112# 0.010862f
C9355 trim_mask\[2\] FILLER_0_2_93/a_124_375# 0.046032f
C9356 _127_ vdd 0.155954f
C9357 FILLER_0_12_50/a_124_375# cal_count\[0\] 0.002359f
C9358 net36 FILLER_0_15_235/a_36_472# 0.00664f
C9359 net65 FILLER_0_3_172/a_572_375# 0.008318f
C9360 _259_/a_455_68# net20 0.001427f
C9361 FILLER_0_7_104/a_124_375# _131_ 0.001291f
C9362 trim_val\[4\] net47 0.003977f
C9363 net36 _438_/a_36_151# 0.076525f
C9364 result[9] _417_/a_2560_156# 0.00263f
C9365 _143_ _140_ 0.00806f
C9366 _389_/a_36_148# FILLER_0_10_94/a_124_375# 0.004673f
C9367 _024_ FILLER_0_22_177/a_36_472# 0.003242f
C9368 _274_/a_36_68# FILLER_0_12_220/a_932_472# 0.001237f
C9369 net63 mask\[2\] 0.553545f
C9370 FILLER_0_18_2/a_932_472# net55 0.012117f
C9371 net57 _120_ 0.012391f
C9372 FILLER_0_8_107/a_124_375# vdd 0.049132f
C9373 FILLER_0_12_136/a_932_472# vss 0.008682f
C9374 FILLER_0_12_136/a_1380_472# vdd 0.006419f
C9375 _069_ _117_ 0.041311f
C9376 _065_ ctln[9] 0.123393f
C9377 _130_ FILLER_0_11_124/a_36_472# 0.003572f
C9378 FILLER_0_17_142/a_484_472# _137_ 0.003953f
C9379 output10/a_224_472# vss 0.014205f
C9380 _009_ vss 0.105833f
C9381 net34 output34/a_224_472# 0.031833f
C9382 _437_/a_2248_156# _436_/a_36_151# 0.001837f
C9383 FILLER_0_9_28/a_1468_375# net68 0.013121f
C9384 _009_ _298_/a_224_472# 0.002441f
C9385 _111_ vss 0.233815f
C9386 net20 _429_/a_36_151# 0.002103f
C9387 _308_/a_124_24# net50 0.02221f
C9388 _423_/a_2665_112# _012_ 0.014394f
C9389 FILLER_0_5_109/a_36_472# vdd 0.042799f
C9390 _114_ FILLER_0_11_101/a_572_375# 0.051108f
C9391 FILLER_0_9_223/a_572_375# _128_ 0.006559f
C9392 _189_/a_67_603# _043_ 0.005635f
C9393 _164_ _160_ 1.863027f
C9394 FILLER_0_21_286/a_484_472# _420_/a_36_151# 0.027236f
C9395 _096_ vss 0.126096f
C9396 _071_ vdd 0.074299f
C9397 FILLER_0_19_111/a_484_472# vdd 0.009246f
C9398 net79 FILLER_0_12_220/a_484_472# 0.005464f
C9399 _023_ vdd 0.062542f
C9400 FILLER_0_19_187/a_36_472# vdd 0.09884f
C9401 FILLER_0_19_187/a_572_375# vss 0.055266f
C9402 fanout60/a_36_160# FILLER_0_17_282/a_36_472# 0.002647f
C9403 fanout78/a_36_113# vss 0.031944f
C9404 net44 _221_/a_36_160# 0.013363f
C9405 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_124_375# 0.012001f
C9406 net14 FILLER_0_10_94/a_36_472# 0.003391f
C9407 calibrate _059_ 0.506928f
C9408 mask\[7\] FILLER_0_22_177/a_1468_375# 0.001315f
C9409 _174_ FILLER_0_15_59/a_124_375# 0.00622f
C9410 output48/a_224_472# calibrate 0.003223f
C9411 ctlp[3] _422_/a_2665_112# 0.001024f
C9412 _414_/a_796_472# cal_itt\[3\] 0.019699f
C9413 _432_/a_448_472# net80 0.045963f
C9414 net38 vdd 0.906502f
C9415 state\[1\] net23 0.075055f
C9416 output11/a_224_472# vdd 0.01016f
C9417 FILLER_0_15_150/a_124_375# _095_ 0.003939f
C9418 valid en 0.026142f
C9419 _375_/a_36_68# calibrate 0.048799f
C9420 net48 net4 0.099614f
C9421 FILLER_0_21_28/a_1916_375# vdd -0.009753f
C9422 FILLER_0_21_125/a_36_472# _433_/a_36_151# 0.001723f
C9423 FILLER_0_3_172/a_932_472# vdd 0.009887f
C9424 _386_/a_848_380# vss 0.012638f
C9425 _442_/a_36_151# FILLER_0_2_127/a_124_375# 0.001597f
C9426 _414_/a_796_472# _081_ 0.003538f
C9427 net17 output40/a_224_472# 0.00187f
C9428 _443_/a_36_151# _152_ 0.002345f
C9429 _427_/a_36_151# net74 0.04306f
C9430 net4 FILLER_0_3_221/a_36_472# 0.010517f
C9431 _438_/a_2248_156# net14 0.045909f
C9432 fanout58/a_36_160# cal_itt\[1\] 0.010654f
C9433 cal_itt\[1\] cal_itt\[0\] 0.055355f
C9434 _076_ _078_ 0.012626f
C9435 _359_/a_1044_488# _133_ 0.001894f
C9436 _359_/a_1492_488# _070_ 0.0043f
C9437 _359_/a_36_488# _076_ 0.005184f
C9438 _093_ FILLER_0_18_107/a_2724_472# 0.00308f
C9439 FILLER_0_18_100/a_36_472# vss 0.002412f
C9440 trim_mask\[1\] _156_ 0.007519f
C9441 _431_/a_36_151# _334_/a_36_160# 0.032942f
C9442 FILLER_0_22_177/a_572_375# net33 0.013337f
C9443 FILLER_0_6_177/a_484_472# FILLER_0_5_181/a_36_472# 0.05841f
C9444 FILLER_0_15_142/a_124_375# fanout73/a_36_113# 0.00146f
C9445 _444_/a_1204_472# net47 0.007847f
C9446 _091_ FILLER_0_12_220/a_572_375# 0.003075f
C9447 net69 net66 0.09789f
C9448 _120_ FILLER_0_10_107/a_572_375# 0.002214f
C9449 FILLER_0_20_107/a_36_472# _438_/a_2665_112# 0.035266f
C9450 FILLER_0_10_214/a_36_472# vdd 0.026621f
C9451 FILLER_0_10_214/a_124_375# vss 0.013034f
C9452 net20 _055_ 0.203142f
C9453 _372_/a_358_69# _160_ 0.001562f
C9454 _005_ _416_/a_2248_156# 0.036714f
C9455 trim_val\[3\] net49 0.009336f
C9456 net50 trim_mask\[3\] 0.001654f
C9457 _442_/a_448_472# _031_ 0.019293f
C9458 _053_ FILLER_0_7_104/a_484_472# 0.005353f
C9459 _131_ FILLER_0_11_124/a_124_375# 0.008946f
C9460 result[0] FILLER_0_9_290/a_124_375# 0.030628f
C9461 FILLER_0_14_81/a_36_472# _451_/a_3129_107# 0.001557f
C9462 ctlp[7] output25/a_224_472# 0.002088f
C9463 output36/a_224_472# net62 0.317201f
C9464 mask\[7\] net19 0.003605f
C9465 _261_/a_36_160# FILLER_0_5_136/a_36_472# 0.00304f
C9466 net50 net67 0.518421f
C9467 fanout58/a_36_160# vss 0.039959f
C9468 cal_itt\[0\] vss 0.11965f
C9469 FILLER_0_21_125/a_124_375# _140_ 0.031374f
C9470 FILLER_0_10_256/a_124_375# vdd 0.041848f
C9471 _005_ _099_ 0.001603f
C9472 trim_mask\[2\] FILLER_0_3_54/a_36_472# 0.004063f
C9473 _432_/a_36_151# mask\[2\] 0.031341f
C9474 net4 net19 0.050898f
C9475 net56 FILLER_0_17_142/a_484_472# 0.008895f
C9476 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_572_375# 0.086635f
C9477 mask\[7\] mask\[6\] 0.227476f
C9478 fanout55/a_36_160# vss 0.005203f
C9479 net22 _435_/a_2248_156# 0.003453f
C9480 _114_ _136_ 0.003405f
C9481 mask\[0\] _429_/a_2248_156# 0.016246f
C9482 net75 output11/a_224_472# 0.015211f
C9483 FILLER_0_4_107/a_932_472# FILLER_0_2_111/a_572_375# 0.001512f
C9484 _088_ net59 0.270902f
C9485 FILLER_0_7_162/a_36_472# vdd 0.026981f
C9486 _114_ net21 0.022033f
C9487 _089_ _414_/a_796_472# 0.001426f
C9488 net63 FILLER_0_22_177/a_1020_375# 0.003419f
C9489 net38 _452_/a_1040_527# 0.002024f
C9490 cal_count\[1\] _180_ 0.300952f
C9491 _415_/a_2665_112# FILLER_0_9_290/a_36_472# 0.007376f
C9492 FILLER_0_5_128/a_572_375# net74 0.050735f
C9493 _193_/a_36_160# vss 0.035228f
C9494 FILLER_0_20_177/a_932_472# _098_ 0.008366f
C9495 net58 _412_/a_796_472# 0.001182f
C9496 output25/a_224_472# net25 0.179738f
C9497 FILLER_0_5_212/a_124_375# _122_ 0.001352f
C9498 _077_ _439_/a_448_472# 0.052962f
C9499 _103_ _418_/a_1204_472# 0.00582f
C9500 net2 input4/a_36_68# 0.031809f
C9501 output26/a_224_472# _423_/a_36_151# 0.011936f
C9502 net62 vdd 1.53102f
C9503 _431_/a_36_151# net36 0.006618f
C9504 _411_/a_448_472# ctln[1] 0.039538f
C9505 _365_/a_36_68# vss 0.029516f
C9506 _115_ _449_/a_2665_112# 0.00947f
C9507 FILLER_0_16_241/a_124_375# _282_/a_36_160# 0.005398f
C9508 FILLER_0_16_89/a_36_472# _397_/a_36_472# 0.004546f
C9509 FILLER_0_9_105/a_124_375# FILLER_0_10_107/a_36_472# 0.001543f
C9510 FILLER_0_11_101/a_124_375# _171_ 0.00105f
C9511 cal_count\[1\] _451_/a_2225_156# 0.006336f
C9512 FILLER_0_14_107/a_124_375# _040_ 0.001861f
C9513 net45 trimb[3] 0.001109f
C9514 _093_ mask\[9\] 0.460108f
C9515 net36 net22 0.034258f
C9516 _114_ _070_ 0.507391f
C9517 _011_ net78 0.002956f
C9518 FILLER_0_20_193/a_124_375# FILLER_0_20_177/a_1468_375# 0.012222f
C9519 net50 FILLER_0_8_24/a_484_472# 0.059367f
C9520 FILLER_0_18_2/a_2724_472# net55 0.007511f
C9521 _056_ state\[1\] 0.219625f
C9522 FILLER_0_9_28/a_932_472# FILLER_0_10_37/a_36_472# 0.026657f
C9523 _093_ FILLER_0_17_72/a_932_472# 0.004367f
C9524 vss FILLER_0_5_148/a_124_375# 0.018465f
C9525 vdd FILLER_0_5_148/a_572_375# -0.009701f
C9526 _233_/a_36_160# vdd 0.064615f
C9527 _024_ _023_ 0.005966f
C9528 result[4] _417_/a_448_472# 0.003485f
C9529 _199_/a_36_160# vdd 0.036579f
C9530 net81 _429_/a_2560_156# 0.003888f
C9531 _432_/a_2560_156# _136_ 0.001178f
C9532 FILLER_0_2_171/a_36_472# vss 0.002909f
C9533 net74 FILLER_0_13_72/a_36_472# 0.007448f
C9534 _246_/a_36_68# vdd 0.047419f
C9535 net63 FILLER_0_18_177/a_2364_375# 0.009893f
C9536 net63 net20 0.045207f
C9537 net75 FILLER_0_10_256/a_124_375# 0.027258f
C9538 net15 _394_/a_718_524# 0.027444f
C9539 _360_/a_36_160# _160_ 0.052885f
C9540 result[5] _418_/a_2248_156# 0.001309f
C9541 cal input4/a_36_68# 0.054357f
C9542 _144_ FILLER_0_21_125/a_484_472# 0.001616f
C9543 net20 FILLER_0_13_212/a_1468_375# 0.009573f
C9544 _098_ _348_/a_49_472# 0.011096f
C9545 ctlp[6] _050_ 0.100418f
C9546 FILLER_0_19_47/a_484_472# _013_ 0.009677f
C9547 _053_ _414_/a_2665_112# 0.032254f
C9548 mask\[7\] _009_ 0.078131f
C9549 _408_/a_1336_472# _043_ 0.023648f
C9550 FILLER_0_4_185/a_36_472# net22 0.006506f
C9551 _431_/a_36_151# FILLER_0_14_123/a_124_375# 0.002807f
C9552 _415_/a_1308_423# net19 0.001498f
C9553 _428_/a_1308_423# _017_ 0.005962f
C9554 _428_/a_448_472# net53 0.001959f
C9555 _116_ _090_ 0.122467f
C9556 FILLER_0_21_28/a_1916_375# _424_/a_36_151# 0.059049f
C9557 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_572_375# 0.007947f
C9558 FILLER_0_19_155/a_124_375# vdd 0.019233f
C9559 FILLER_0_18_107/a_3172_472# _145_ 0.002415f
C9560 _069_ FILLER_0_18_209/a_484_472# 0.013944f
C9561 FILLER_0_16_57/a_932_472# cal_count\[1\] 0.002217f
C9562 net7 net68 0.032489f
C9563 net45 ctlp[0] 0.001134f
C9564 net59 rstn 0.039664f
C9565 _074_ _123_ 0.157299f
C9566 _098_ _438_/a_2248_156# 0.002798f
C9567 _247_/a_36_160# _228_/a_36_68# 0.001919f
C9568 FILLER_0_2_111/a_484_472# _158_ 0.003604f
C9569 FILLER_0_5_54/a_124_375# net47 0.012889f
C9570 net82 FILLER_0_3_172/a_1916_375# 0.010202f
C9571 net55 vdd 1.248648f
C9572 FILLER_0_2_165/a_36_472# vss 0.001099f
C9573 _452_/a_3129_107# vdd 0.016611f
C9574 _080_ FILLER_0_3_221/a_932_472# 0.003217f
C9575 _397_/a_36_472# FILLER_0_17_72/a_1468_375# 0.001295f
C9576 FILLER_0_4_123/a_124_375# net74 0.002449f
C9577 _126_ FILLER_0_11_124/a_124_375# 0.038971f
C9578 _185_ _405_/a_255_603# 0.002565f
C9579 _369_/a_36_68# vdd 0.042534f
C9580 _076_ FILLER_0_6_231/a_36_472# 0.005517f
C9581 ctlp[4] output22/a_224_472# 0.008275f
C9582 ctln[6] vss 0.45431f
C9583 _267_/a_224_472# _121_ 0.0029f
C9584 _394_/a_728_93# _095_ 0.035417f
C9585 _302_/a_224_472# vss 0.005149f
C9586 net18 _419_/a_36_151# 0.021491f
C9587 _137_ FILLER_0_16_154/a_572_375# 0.010132f
C9588 _116_ net22 0.122052f
C9589 _028_ FILLER_0_7_104/a_484_472# 0.00499f
C9590 _077_ FILLER_0_8_156/a_484_472# 0.006446f
C9591 FILLER_0_7_72/a_1916_375# net52 0.001608f
C9592 FILLER_0_12_2/a_572_375# net3 0.001872f
C9593 cal_itt\[3\] _251_/a_1130_472# 0.001099f
C9594 _256_/a_2552_68# _072_ 0.001213f
C9595 _046_ _282_/a_36_160# 0.005584f
C9596 output39/a_224_472# net40 0.087367f
C9597 net81 _425_/a_36_151# 0.014663f
C9598 output27/a_224_472# FILLER_0_9_282/a_36_472# 0.001711f
C9599 _429_/a_36_151# vss 0.026298f
C9600 _429_/a_448_472# vdd 0.008822f
C9601 FILLER_0_10_78/a_1020_375# vss 0.002352f
C9602 _079_ _073_ 0.234533f
C9603 net39 FILLER_0_8_2/a_36_472# 0.010296f
C9604 FILLER_0_14_50/a_124_375# _180_ 0.022435f
C9605 FILLER_0_7_72/a_932_472# net52 0.008749f
C9606 net56 net54 0.018493f
C9607 _095_ FILLER_0_13_80/a_36_472# 0.004187f
C9608 _053_ FILLER_0_4_213/a_572_375# 0.003451f
C9609 state\[1\] FILLER_0_12_196/a_124_375# 0.063785f
C9610 _132_ _428_/a_1000_472# 0.027767f
C9611 _415_/a_2248_156# net64 0.051575f
C9612 _413_/a_36_151# FILLER_0_2_177/a_484_472# 0.006095f
C9613 _093_ net35 0.00127f
C9614 FILLER_0_16_89/a_484_472# _176_ 0.004026f
C9615 mask\[1\] FILLER_0_15_180/a_36_472# 0.001145f
C9616 _077_ _319_/a_672_472# 0.001602f
C9617 ctlp[1] FILLER_0_21_286/a_572_375# 0.026009f
C9618 _423_/a_36_151# FILLER_0_23_60/a_124_375# 0.005577f
C9619 net23 vdd 1.576398f
C9620 _428_/a_2560_156# _043_ 0.009909f
C9621 FILLER_0_22_128/a_1468_375# vss 0.006619f
C9622 _057_ cal_count\[3\] 0.416063f
C9623 net25 FILLER_0_22_86/a_36_472# 0.001265f
C9624 net81 net1 0.03613f
C9625 FILLER_0_18_2/a_572_375# net38 0.007477f
C9626 _086_ _176_ 0.837546f
C9627 _396_/a_224_472# _177_ 0.001254f
C9628 FILLER_0_23_290/a_124_375# vdd 0.030435f
C9629 _424_/a_796_472# vdd 0.001951f
C9630 _083_ FILLER_0_3_221/a_1380_472# 0.00181f
C9631 net79 net19 0.03862f
C9632 net15 net49 0.057277f
C9633 _441_/a_2665_112# vdd 0.012404f
C9634 _441_/a_2248_156# vss 0.005663f
C9635 trim_val\[2\] vss 0.027243f
C9636 FILLER_0_11_64/a_36_472# vss 0.006069f
C9637 mask\[5\] FILLER_0_20_177/a_1020_375# 0.013294f
C9638 FILLER_0_8_107/a_36_472# net14 0.001596f
C9639 net72 net55 0.233515f
C9640 net55 _452_/a_1040_527# 0.021721f
C9641 _053_ FILLER_0_6_47/a_1020_375# 0.015621f
C9642 net15 net68 0.205016f
C9643 mask\[3\] FILLER_0_18_177/a_484_472# 0.005654f
C9644 _447_/a_1000_472# vdd 0.003392f
C9645 _117_ _090_ 0.041465f
C9646 _412_/a_36_151# net81 0.014094f
C9647 fanout74/a_36_113# vdd 0.099021f
C9648 net76 FILLER_0_1_192/a_36_472# 0.003817f
C9649 net63 FILLER_0_19_187/a_124_375# 0.012282f
C9650 result[2] net30 0.019568f
C9651 _439_/a_1204_472# vss 0.006567f
C9652 _367_/a_36_68# _157_ 0.013352f
C9653 net74 _163_ 0.042013f
C9654 net4 cal_itt\[0\] 0.054266f
C9655 FILLER_0_17_56/a_124_375# FILLER_0_18_53/a_484_472# 0.001597f
C9656 _094_ _196_/a_36_160# 0.001668f
C9657 _153_ FILLER_0_4_91/a_572_375# 0.001735f
C9658 net3 net17 0.045911f
C9659 _177_ _150_ 0.002507f
C9660 _136_ _018_ 0.002892f
C9661 _141_ mask\[6\] 0.009844f
C9662 mask\[9\] FILLER_0_18_76/a_572_375# 0.006158f
C9663 output35/a_224_472# net35 0.007217f
C9664 output34/a_224_472# net20 0.023142f
C9665 _115_ net74 0.033145f
C9666 _018_ net21 0.077174f
C9667 net76 FILLER_0_3_172/a_1828_472# 0.051851f
C9668 _426_/a_36_151# FILLER_0_8_247/a_932_472# 0.001723f
C9669 _055_ vss 0.365503f
C9670 mask\[0\] _100_ 0.005921f
C9671 fanout49/a_36_160# trim_mask\[1\] 0.00358f
C9672 _116_ _076_ 0.008283f
C9673 _085_ _070_ 0.058787f
C9674 _091_ state\[0\] 0.012343f
C9675 FILLER_0_17_72/a_484_472# FILLER_0_18_76/a_36_472# 0.05841f
C9676 mask\[5\] _137_ 0.002972f
C9677 _091_ FILLER_0_18_177/a_1020_375# 0.002226f
C9678 net56 FILLER_0_18_139/a_484_472# 0.004375f
C9679 vdd _381_/a_36_472# 0.014305f
C9680 _428_/a_36_151# FILLER_0_14_107/a_484_472# 0.059367f
C9681 result[6] _421_/a_36_151# 0.032036f
C9682 fanout80/a_36_113# net81 0.097873f
C9683 net57 _043_ 1.955053f
C9684 net76 net37 0.549565f
C9685 fanout60/a_36_160# vss 0.035381f
C9686 net67 _054_ 0.391592f
C9687 _025_ vdd 0.259346f
C9688 net56 FILLER_0_16_154/a_572_375# 0.002321f
C9689 FILLER_0_16_73/a_124_375# net55 0.007695f
C9690 _074_ _305_/a_36_159# 0.012602f
C9691 FILLER_0_8_138/a_36_472# _077_ 0.005953f
C9692 _371_/a_36_113# _370_/a_124_24# 0.008354f
C9693 mask\[5\] FILLER_0_19_171/a_36_472# 0.002923f
C9694 _411_/a_36_151# _073_ 0.00135f
C9695 FILLER_0_15_10/a_36_472# vdd 0.086171f
C9696 FILLER_0_15_10/a_124_375# vss 0.002173f
C9697 _245_/a_672_472# net17 0.00121f
C9698 net19 _416_/a_2665_112# 0.059453f
C9699 cal_count\[3\] _042_ 0.001716f
C9700 net55 _424_/a_36_151# 0.007344f
C9701 net39 _063_ 0.004732f
C9702 FILLER_0_15_142/a_124_375# vss 0.009207f
C9703 _311_/a_1660_473# vdd 0.001435f
C9704 _285_/a_36_472# _099_ 0.040922f
C9705 net20 net10 0.02842f
C9706 _251_/a_906_472# _070_ 0.002124f
C9707 cal_itt\[2\] _079_ 0.017071f
C9708 net33 vdd 0.42212f
C9709 _431_/a_1308_423# vdd 0.002397f
C9710 _154_ vss 0.200253f
C9711 _313_/a_67_603# vss 0.016047f
C9712 net24 FILLER_0_23_88/a_36_472# 0.006289f
C9713 _081_ _082_ 0.008298f
C9714 _343_/a_49_472# vss 0.002581f
C9715 ctln[7] vss 0.132613f
C9716 _079_ net1 0.099822f
C9717 _062_ FILLER_0_5_136/a_36_472# 0.001404f
C9718 net18 FILLER_0_17_282/a_124_375# 0.048177f
C9719 _053_ net48 0.003159f
C9720 _077_ FILLER_0_9_72/a_484_472# 0.004472f
C9721 _427_/a_2665_112# vss 0.01229f
C9722 _056_ vdd 0.423512f
C9723 result[9] _108_ 0.015443f
C9724 result[4] _418_/a_448_472# 0.004918f
C9725 FILLER_0_3_221/a_124_375# FILLER_0_3_212/a_124_375# 0.002036f
C9726 mask\[4\] FILLER_0_20_193/a_484_472# 0.001215f
C9727 trim_val\[1\] _166_ 0.06773f
C9728 FILLER_0_10_28/a_124_375# _450_/a_3129_107# 0.010735f
C9729 net73 _098_ 0.004745f
C9730 net28 _044_ 0.481924f
C9731 _053_ _162_ 0.00209f
C9732 _176_ net53 0.083005f
C9733 FILLER_0_8_24/a_484_472# _054_ 0.009315f
C9734 FILLER_0_14_81/a_124_375# _394_/a_728_93# 0.004587f
C9735 _095_ _067_ 0.00784f
C9736 FILLER_0_14_263/a_124_375# output30/a_224_472# 0.011584f
C9737 _096_ net79 0.015605f
C9738 _322_/a_692_472# _129_ 0.004891f
C9739 _002_ FILLER_0_3_172/a_2276_472# 0.030358f
C9740 trim_val\[4\] vdd 0.245329f
C9741 _069_ _059_ 0.002034f
C9742 _392_/a_36_68# vdd 0.036386f
C9743 net38 _444_/a_1308_423# 0.007915f
C9744 FILLER_0_14_50/a_36_472# cal_count\[3\] 0.005814f
C9745 _024_ net23 0.001994f
C9746 fanout78/a_36_113# net79 0.029496f
C9747 mask\[4\] FILLER_0_18_139/a_1380_472# 0.003851f
C9748 FILLER_0_8_37/a_572_375# _054_ 0.137749f
C9749 FILLER_0_14_99/a_124_375# _095_ 0.012128f
C9750 net63 vss 0.566021f
C9751 _238_/a_67_603# net14 0.004718f
C9752 _449_/a_2665_112# _067_ 0.03661f
C9753 output38/a_224_472# _446_/a_36_151# 0.117966f
C9754 net34 _422_/a_36_151# 0.032272f
C9755 FILLER_0_13_212/a_1468_375# vss 0.062822f
C9756 FILLER_0_13_212/a_36_472# vdd 0.105926f
C9757 net62 FILLER_0_13_212/a_572_375# 0.001597f
C9758 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_124_375# 0.001597f
C9759 net32 _107_ 0.003155f
C9760 _081_ _265_/a_244_68# 0.03338f
C9761 _012_ FILLER_0_23_44/a_572_375# 0.002827f
C9762 _436_/a_1000_472# vdd 0.006522f
C9763 output20/a_224_472# result[8] 0.038114f
C9764 _125_ _134_ 0.00437f
C9765 trim_mask\[2\] trim_val\[2\] 0.21814f
C9766 FILLER_0_17_200/a_572_375# net21 0.011557f
C9767 _064_ _447_/a_36_151# 0.004185f
C9768 mask\[5\] _434_/a_2248_156# 0.003462f
C9769 vss _433_/a_1308_423# 0.002695f
C9770 _112_ _081_ 0.037903f
C9771 _176_ FILLER_0_11_78/a_124_375# 0.004803f
C9772 _438_/a_448_472# _437_/a_36_151# 0.00198f
C9773 net60 _418_/a_2248_156# 0.045472f
C9774 _058_ vss 0.19427f
C9775 output47/a_224_472# net44 0.077292f
C9776 net66 _440_/a_448_472# 0.023934f
C9777 net60 _419_/a_3041_156# 0.001022f
C9778 net52 FILLER_0_6_79/a_124_375# 0.010099f
C9779 FILLER_0_18_2/a_572_375# _452_/a_3129_107# 0.001073f
C9780 _431_/a_1288_156# net73 0.001033f
C9781 net20 FILLER_0_1_212/a_36_472# 0.013846f
C9782 mask\[8\] _423_/a_2248_156# 0.001648f
C9783 _315_/a_36_68# vss 0.02467f
C9784 _394_/a_728_93# cal_count\[1\] 0.057049f
C9785 net60 _011_ 0.003094f
C9786 result[2] FILLER_0_14_263/a_36_472# 0.001134f
C9787 net74 FILLER_0_13_80/a_36_472# 0.00679f
C9788 _132_ FILLER_0_17_104/a_1468_375# 0.051996f
C9789 output21/a_224_472# vss 0.082781f
C9790 net50 trim_val\[1\] 0.002079f
C9791 ctlp[1] _420_/a_448_472# 0.038053f
C9792 _440_/a_796_472# _029_ 0.009261f
C9793 _159_ _160_ 0.021804f
C9794 mask\[7\] FILLER_0_22_128/a_1468_375# 0.0178f
C9795 FILLER_0_16_241/a_124_375# vdd 0.035603f
C9796 FILLER_0_5_198/a_36_472# vdd 0.088893f
C9797 FILLER_0_5_198/a_572_375# vss 0.055087f
C9798 _260_/a_36_68# net59 0.004346f
C9799 _053_ FILLER_0_6_79/a_36_472# 0.001777f
C9800 net54 FILLER_0_22_86/a_932_472# 0.047897f
C9801 _254_/a_244_472# _074_ 0.002716f
C9802 net35 FILLER_0_22_128/a_932_472# 0.007806f
C9803 _126_ _138_ 0.003253f
C9804 output29/a_224_472# net19 0.09445f
C9805 _064_ trim[1] 0.166575f
C9806 net36 _451_/a_1040_527# 0.00974f
C9807 FILLER_0_12_220/a_124_375# _248_/a_36_68# 0.005308f
C9808 cal_count\[1\] FILLER_0_13_80/a_36_472# 0.001559f
C9809 output46/a_224_472# net38 0.003296f
C9810 _411_/a_1308_423# net75 0.028281f
C9811 _367_/a_692_472# net14 0.00423f
C9812 vdd FILLER_0_12_196/a_124_375# 0.015159f
C9813 _363_/a_36_68# vdd 0.04306f
C9814 cal_count\[3\] net40 0.080767f
C9815 net82 _316_/a_848_380# 0.087022f
C9816 net64 FILLER_0_9_282/a_124_375# 0.046477f
C9817 output14/a_224_472# net14 0.018674f
C9818 _136_ FILLER_0_16_154/a_484_472# 0.007583f
C9819 output39/a_224_472# _445_/a_448_472# 0.009352f
C9820 trim_mask\[1\] FILLER_0_6_47/a_3260_375# 0.003764f
C9821 FILLER_0_1_266/a_124_375# net8 0.012703f
C9822 net20 FILLER_0_15_212/a_1020_375# 0.001629f
C9823 _024_ net33 0.001047f
C9824 _070_ _310_/a_49_472# 0.00564f
C9825 _052_ FILLER_0_18_37/a_124_375# 0.03242f
C9826 _444_/a_1204_472# vdd 0.001086f
C9827 net31 _102_ 0.060034f
C9828 net79 _193_/a_36_160# 0.010228f
C9829 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_124_375# 0.003732f
C9830 FILLER_0_10_78/a_932_472# _439_/a_2665_112# 0.001182f
C9831 _176_ FILLER_0_11_109/a_36_472# 0.002951f
C9832 _446_/a_36_151# vdd 0.06703f
C9833 _421_/a_36_151# _419_/a_2248_156# 0.001203f
C9834 ctlp[1] _421_/a_796_472# 0.001754f
C9835 ctlp[1] fanout77/a_36_113# 0.012793f
C9836 net53 FILLER_0_13_142/a_124_375# 0.001599f
C9837 _430_/a_448_472# _091_ 0.065306f
C9838 _316_/a_692_472# _122_ 0.002929f
C9839 _316_/a_1152_472# calibrate 0.001604f
C9840 fanout54/a_36_160# FILLER_0_19_142/a_36_472# 0.002647f
C9841 mask\[4\] FILLER_0_18_209/a_484_472# 0.021522f
C9842 _255_/a_224_552# _116_ 0.027303f
C9843 net4 _055_ 0.216844f
C9844 net22 FILLER_0_18_209/a_484_472# 0.005297f
C9845 FILLER_0_4_91/a_124_375# _160_ 0.009765f
C9846 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1468_375# 0.086635f
C9847 FILLER_0_11_101/a_36_472# FILLER_0_13_100/a_124_375# 0.001436f
C9848 _432_/a_36_151# vss 0.003647f
C9849 _372_/a_1602_69# _152_ 0.00262f
C9850 _414_/a_2665_112# cal_itt\[3\] 0.02392f
C9851 FILLER_0_6_239/a_36_472# _123_ 0.004433f
C9852 FILLER_0_20_87/a_36_472# net71 0.003995f
C9853 mask\[8\] FILLER_0_22_107/a_572_375# 0.030641f
C9854 net35 FILLER_0_22_107/a_124_375# 0.010439f
C9855 net50 _168_ 0.306226f
C9856 _272_/a_36_472# _079_ 0.0237f
C9857 FILLER_0_12_136/a_124_375# net57 0.001727f
C9858 _055_ _311_/a_692_473# 0.003127f
C9859 _417_/a_448_472# result[3] 0.003109f
C9860 FILLER_0_16_89/a_1468_375# _136_ 0.005791f
C9861 _245_/a_672_472# _039_ 0.001025f
C9862 FILLER_0_13_65/a_124_375# fanout72/a_36_113# 0.005467f
C9863 net34 net21 0.036237f
C9864 FILLER_0_7_104/a_1468_375# _133_ 0.003206f
C9865 _097_ FILLER_0_15_180/a_36_472# 0.005242f
C9866 _414_/a_2665_112# _081_ 0.00247f
C9867 _129_ _062_ 0.20212f
C9868 FILLER_0_13_80/a_124_375# FILLER_0_13_72/a_572_375# 0.012001f
C9869 FILLER_0_12_136/a_572_375# _126_ 0.01289f
C9870 _098_ FILLER_0_15_228/a_124_375# 0.080662f
C9871 net27 _426_/a_2560_156# 0.004199f
C9872 _176_ _451_/a_36_151# 0.003176f
C9873 net81 _195_/a_67_603# 0.002322f
C9874 net73 _131_ 0.022043f
C9875 output35/a_224_472# FILLER_0_21_206/a_36_472# 0.0323f
C9876 output34/a_224_472# vss 0.011966f
C9877 _405_/a_67_603# net17 0.014714f
C9878 ctlp[2] net19 0.017506f
C9879 _094_ _418_/a_1000_472# 0.053462f
C9880 net54 mask\[8\] 0.162104f
C9881 FILLER_0_18_107/a_572_375# mask\[9\] 0.005368f
C9882 _046_ vdd 0.041841f
C9883 _430_/a_1308_423# vdd 0.00218f
C9884 output32/a_224_472# net18 0.022521f
C9885 net52 _386_/a_124_24# 0.001051f
C9886 cal_count\[3\] FILLER_0_12_20/a_124_375# 0.008038f
C9887 _008_ result[4] 0.134001f
C9888 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_36_472# 0.003468f
C9889 output45/a_224_472# trimb[0] 0.003753f
C9890 FILLER_0_4_197/a_932_472# net21 0.00663f
C9891 output44/a_224_472# FILLER_0_20_15/a_932_472# 0.0323f
C9892 FILLER_0_11_124/a_36_472# _118_ 0.002798f
C9893 net15 FILLER_0_17_72/a_572_375# 0.003021f
C9894 fanout80/a_36_113# mask\[1\] 0.020046f
C9895 _207_/a_67_603# _049_ 0.003205f
C9896 ctln[3] net19 0.003077f
C9897 net62 _416_/a_2248_156# 0.043158f
C9898 _420_/a_36_151# FILLER_0_23_282/a_572_375# 0.059049f
C9899 FILLER_0_21_286/a_36_472# _009_ 0.003266f
C9900 _414_/a_2248_156# _056_ 0.001452f
C9901 FILLER_0_16_89/a_36_472# FILLER_0_17_72/a_1916_375# 0.001723f
C9902 FILLER_0_16_89/a_1020_375# FILLER_0_17_72/a_2812_375# 0.026339f
C9903 FILLER_0_20_169/a_36_472# _140_ 0.023696f
C9904 _149_ FILLER_0_20_87/a_124_375# 0.004191f
C9905 net74 _067_ 0.674895f
C9906 _413_/a_2665_112# output11/a_224_472# 0.001492f
C9907 _122_ FILLER_0_8_156/a_484_472# 0.007378f
C9908 FILLER_0_13_142/a_1380_472# _043_ 0.011974f
C9909 net76 _122_ 0.028025f
C9910 _056_ _311_/a_254_473# 0.005937f
C9911 net10 vss 0.324553f
C9912 net65 net59 0.790496f
C9913 _411_/a_2248_156# _084_ 0.002258f
C9914 net50 FILLER_0_4_91/a_572_375# 0.007234f
C9915 FILLER_0_4_152/a_36_472# net23 0.047194f
C9916 net28 fanout79/a_36_160# 0.036675f
C9917 net63 mask\[7\] 0.069252f
C9918 FILLER_0_21_125/a_124_375# _098_ 0.006462f
C9919 _140_ FILLER_0_22_128/a_2276_472# 0.002954f
C9920 FILLER_0_18_139/a_572_375# FILLER_0_19_142/a_124_375# 0.026339f
C9921 net58 FILLER_0_9_282/a_36_472# 0.062389f
C9922 _186_ _184_ 0.047995f
C9923 net15 FILLER_0_15_59/a_572_375# 0.033245f
C9924 net62 _099_ 0.062012f
C9925 FILLER_0_0_232/a_36_472# vdd 0.050082f
C9926 FILLER_0_0_232/a_124_375# vss 0.019863f
C9927 _028_ FILLER_0_6_79/a_36_472# 0.016281f
C9928 _069_ _247_/a_36_160# 0.046764f
C9929 _137_ _138_ 0.045916f
C9930 FILLER_0_9_270/a_124_375# vdd 0.013312f
C9931 _392_/a_36_68# cal_count\[0\] 0.038691f
C9932 _339_/a_36_160# FILLER_0_19_171/a_124_375# 0.006021f
C9933 FILLER_0_16_255/a_124_375# _094_ 0.004398f
C9934 net20 FILLER_0_15_235/a_124_375# 0.001278f
C9935 _144_ FILLER_0_19_155/a_572_375# 0.003611f
C9936 _374_/a_36_68# _056_ 0.011052f
C9937 ctlp[1] FILLER_0_24_274/a_1380_472# 0.008573f
C9938 FILLER_0_21_125/a_572_375# _022_ 0.006025f
C9939 _025_ _436_/a_448_472# 0.044246f
C9940 FILLER_0_3_142/a_124_375# net23 0.25251f
C9941 _428_/a_1000_472# vdd 0.005345f
C9942 _431_/a_2560_156# net53 0.002265f
C9943 _429_/a_36_151# net79 0.02414f
C9944 net69 FILLER_0_2_127/a_36_472# 0.019383f
C9945 net61 _108_ 0.030767f
C9946 trim_mask\[4\] _370_/a_1084_68# 0.005157f
C9947 FILLER_0_5_54/a_124_375# vdd 0.007387f
C9948 net80 FILLER_0_20_177/a_124_375# 0.001198f
C9949 net55 _404_/a_36_472# 0.001746f
C9950 FILLER_0_10_247/a_124_375# fanout79/a_36_160# 0.010334f
C9951 net15 net47 0.035839f
C9952 valid fanout65/a_36_113# 0.001646f
C9953 FILLER_0_22_128/a_2724_472# FILLER_0_21_150/a_124_375# 0.001543f
C9954 output36/a_224_472# net18 0.010751f
C9955 _214_/a_36_160# vss 0.007045f
C9956 _136_ FILLER_0_13_100/a_36_472# 0.005029f
C9957 net36 _006_ 0.001331f
C9958 FILLER_0_16_89/a_36_472# net53 0.004701f
C9959 FILLER_0_12_220/a_36_472# _070_ 0.087648f
C9960 FILLER_0_17_226/a_36_472# _093_ 0.004282f
C9961 result[8] FILLER_0_24_274/a_1020_375# 0.00726f
C9962 fanout76/a_36_160# vss 0.028897f
C9963 _061_ FILLER_0_8_156/a_484_472# 0.00255f
C9964 output21/a_224_472# mask\[7\] 0.032297f
C9965 FILLER_0_15_290/a_124_375# FILLER_0_15_282/a_572_375# 0.012001f
C9966 _002_ net82 0.034599f
C9967 net37 FILLER_0_6_231/a_484_472# 0.004323f
C9968 FILLER_0_17_282/a_124_375# _417_/a_36_151# 0.059049f
C9969 FILLER_0_15_72/a_572_375# vss 0.007579f
C9970 FILLER_0_15_72/a_36_472# vdd 0.108844f
C9971 fanout74/a_36_113# FILLER_0_3_142/a_124_375# 0.002073f
C9972 _013_ _041_ 0.00271f
C9973 net52 vss 1.608047f
C9974 FILLER_0_17_72/a_2276_472# _131_ 0.004125f
C9975 FILLER_0_7_146/a_124_375# net23 0.00129f
C9976 _074_ _375_/a_692_497# 0.004556f
C9977 _440_/a_36_151# _164_ 0.003699f
C9978 _196_/a_36_160# FILLER_0_14_263/a_124_375# 0.005732f
C9979 ctlp[2] _009_ 0.220631f
C9980 _425_/a_2248_156# net19 0.010557f
C9981 _128_ _116_ 0.069335f
C9982 _127_ _176_ 0.319517f
C9983 _443_/a_796_472# vss 0.001654f
C9984 _093_ FILLER_0_21_60/a_484_472# 0.001396f
C9985 _033_ FILLER_0_6_37/a_124_375# 0.018812f
C9986 net15 FILLER_0_23_44/a_1468_375# 0.001307f
C9987 result[1] _416_/a_36_151# 0.007739f
C9988 mask\[4\] _343_/a_257_69# 0.001786f
C9989 _431_/a_1000_472# net73 0.035816f
C9990 _413_/a_36_151# net21 0.012223f
C9991 net57 _062_ 0.067654f
C9992 _053_ _365_/a_36_68# 0.001572f
C9993 FILLER_0_9_28/a_932_472# vdd 0.04397f
C9994 FILLER_0_19_55/a_36_472# _013_ 0.005889f
C9995 _136_ mask\[2\] 1.822289f
C9996 net75 FILLER_0_0_232/a_36_472# 0.001514f
C9997 output10/a_224_472# ctln[3] 0.064347f
C9998 _086_ _250_/a_36_68# 0.001132f
C9999 net38 net44 0.523774f
C10000 mask\[2\] net21 0.033368f
C10001 FILLER_0_9_223/a_36_472# _070_ 0.006158f
C10002 _077_ _251_/a_468_472# 0.002497f
C10003 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_124_375# 0.003228f
C10004 net18 vdd 1.496006f
C10005 net19 _420_/a_1308_423# 0.010051f
C10006 mask\[5\] result[8] 0.003797f
C10007 fanout82/a_36_113# net2 0.008681f
C10008 FILLER_0_9_28/a_1380_472# net51 0.002012f
C10009 FILLER_0_1_212/a_36_472# vss 0.00858f
C10010 FILLER_0_7_72/a_124_375# net52 0.029774f
C10011 _067_ FILLER_0_13_72/a_124_375# 0.001782f
C10012 net60 _102_ 0.008212f
C10013 _077_ net68 0.003823f
C10014 _216_/a_67_603# vss 0.012211f
C10015 _053_ FILLER_0_6_177/a_484_472# 0.015994f
C10016 trim_val\[0\] FILLER_0_6_47/a_572_375# 0.03235f
C10017 _132_ FILLER_0_18_107/a_932_472# 0.001369f
C10018 output29/a_224_472# _193_/a_36_160# 0.006363f
C10019 net16 FILLER_0_18_37/a_1468_375# 0.002269f
C10020 net16 net67 0.038448f
C10021 ctln[4] net20 0.00225f
C10022 output27/a_224_472# net5 0.008663f
C10023 _320_/a_1792_472# state\[1\] 0.001901f
C10024 net46 FILLER_0_21_28/a_36_472# 0.051176f
C10025 fanout52/a_36_160# net23 0.009496f
C10026 net15 FILLER_0_9_60/a_124_375# 0.003602f
C10027 _115_ _389_/a_36_148# 0.029505f
C10028 _176_ _071_ 0.002542f
C10029 net74 _370_/a_692_472# 0.005066f
C10030 _120_ _042_ 0.031451f
C10031 ctlp[1] _419_/a_1308_423# 0.00678f
C10032 fanout60/a_36_160# net79 0.069956f
C10033 _096_ _335_/a_257_69# 0.001084f
C10034 net17 _190_/a_36_160# 0.04702f
C10035 _306_/a_36_68# _071_ 0.054312f
C10036 _016_ _129_ 0.002216f
C10037 _387_/a_36_113# vss 0.047621f
C10038 net82 _078_ 0.00197f
C10039 _093_ FILLER_0_17_142/a_36_472# 0.011974f
C10040 state\[1\] FILLER_0_13_142/a_1468_375# 0.010245f
C10041 _406_/a_36_159# vss 0.002509f
C10042 net52 FILLER_0_2_165/a_124_375# 0.002214f
C10043 _448_/a_36_151# net22 0.027581f
C10044 FILLER_0_7_72/a_2276_472# net14 0.004375f
C10045 _434_/a_448_472# mask\[6\] 0.060756f
C10046 net20 _421_/a_1204_472# 0.019627f
C10047 net62 FILLER_0_21_286/a_572_375# 0.003744f
C10048 FILLER_0_21_286/a_484_472# vss 0.008522f
C10049 FILLER_0_2_171/a_36_472# FILLER_0_2_177/a_36_472# 0.003468f
C10050 _077_ FILLER_0_7_72/a_484_472# 0.001332f
C10051 _144_ _345_/a_36_160# 0.00465f
C10052 _256_/a_1164_497# net20 0.001462f
C10053 _421_/a_1000_472# net19 0.03394f
C10054 result[4] _006_ 0.271278f
C10055 _412_/a_2560_156# cal_itt\[1\] 0.00454f
C10056 cal_itt\[3\] _162_ 0.141474f
C10057 FILLER_0_10_37/a_124_375# net16 0.010358f
C10058 _072_ state\[2\] 0.002629f
C10059 net20 _422_/a_36_151# 0.083307f
C10060 result[7] FILLER_0_24_274/a_36_472# 0.006454f
C10061 FILLER_0_15_212/a_1020_375# vss 0.035883f
C10062 FILLER_0_15_212/a_1468_375# vdd 0.010445f
C10063 FILLER_0_4_99/a_124_375# _153_ 0.030839f
C10064 net48 _081_ 0.137029f
C10065 _093_ FILLER_0_18_76/a_572_375# 0.025143f
C10066 FILLER_0_4_197/a_124_375# net22 0.00145f
C10067 FILLER_0_6_90/a_124_375# net14 0.005361f
C10068 state\[0\] _426_/a_2248_156# 0.001198f
C10069 FILLER_0_22_86/a_484_472# _437_/a_36_151# 0.013806f
C10070 FILLER_0_5_164/a_36_472# _386_/a_848_380# 0.001177f
C10071 FILLER_0_7_146/a_36_472# _313_/a_67_603# 0.002287f
C10072 _095_ _450_/a_448_472# 0.001393f
C10073 FILLER_0_4_144/a_484_472# net57 0.003724f
C10074 _363_/a_692_472# _028_ 0.001416f
C10075 FILLER_0_10_78/a_484_472# cal_count\[3\] 0.001112f
C10076 net81 _138_ 0.006815f
C10077 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_36_472# 0.086743f
C10078 FILLER_0_10_28/a_36_472# vss 0.001102f
C10079 _075_ vss 0.046342f
C10080 _050_ FILLER_0_22_128/a_36_472# 0.001098f
C10081 _128_ _117_ 0.045015f
C10082 _343_/a_49_472# _141_ 0.04106f
C10083 _114_ _395_/a_36_488# 0.005314f
C10084 _449_/a_36_151# FILLER_0_12_50/a_36_472# 0.003462f
C10085 fanout75/a_36_113# vdd 0.028614f
C10086 _096_ FILLER_0_14_181/a_36_472# 0.028078f
C10087 FILLER_0_9_28/a_1468_375# vdd 0.009854f
C10088 _086_ FILLER_0_11_135/a_124_375# 0.008238f
C10089 net16 FILLER_0_8_37/a_572_375# 0.004285f
C10090 _172_ vss 0.054608f
C10091 FILLER_0_13_65/a_36_472# _095_ 0.003171f
C10092 net34 FILLER_0_22_177/a_484_472# 0.003953f
C10093 _420_/a_1308_423# _009_ 0.014359f
C10094 _016_ _428_/a_2560_156# 0.003934f
C10095 _445_/a_448_472# net40 0.044285f
C10096 FILLER_0_9_28/a_36_472# net40 0.020589f
C10097 _105_ _107_ 0.020727f
C10098 net40 trim[3] 0.084824f
C10099 ctln[3] cal_itt\[0\] 0.002081f
C10100 net80 _434_/a_1000_472# 0.01421f
C10101 _139_ net36 0.024268f
C10102 _029_ _163_ 0.007545f
C10103 mask\[4\] FILLER_0_18_177/a_1468_375# 0.01587f
C10104 FILLER_0_1_98/a_36_472# net52 0.005688f
C10105 net15 fanout66/a_36_113# 0.024302f
C10106 _443_/a_448_472# net23 0.038188f
C10107 net54 _026_ 0.006401f
C10108 net50 _441_/a_796_472# 0.010626f
C10109 net52 trim_mask\[2\] 0.036196f
C10110 FILLER_0_8_127/a_36_472# _133_ 0.004423f
C10111 cal_count\[3\] _120_ 4.687877f
C10112 _442_/a_2248_156# _157_ 0.002731f
C10113 FILLER_0_13_212/a_1468_375# net79 0.009597f
C10114 output43/a_224_472# trimb[0] 0.043402f
C10115 FILLER_0_4_49/a_572_375# net66 0.074393f
C10116 FILLER_0_5_109/a_484_472# FILLER_0_4_107/a_572_375# 0.001684f
C10117 FILLER_0_12_136/a_1020_375# FILLER_0_13_142/a_484_472# 0.001684f
C10118 trim_mask\[4\] net47 0.264421f
C10119 _086_ _162_ 0.107276f
C10120 _195_/a_67_603# mask\[1\] 0.016836f
C10121 _367_/a_36_68# _160_ 0.013113f
C10122 _096_ _320_/a_1120_472# 0.004315f
C10123 FILLER_0_18_61/a_36_472# vdd 0.08828f
C10124 FILLER_0_18_61/a_124_375# vss 0.021307f
C10125 _114_ _439_/a_2665_112# 0.011015f
C10126 net50 _440_/a_2665_112# 0.009767f
C10127 _202_/a_36_160# _047_ 0.02265f
C10128 net52 _439_/a_1000_472# 0.03537f
C10129 net50 _439_/a_1308_423# 0.008832f
C10130 FILLER_0_12_124/a_36_472# vss 0.001443f
C10131 FILLER_0_4_49/a_124_375# trim_mask\[1\] 0.006676f
C10132 _106_ _069_ 0.006716f
C10133 FILLER_0_17_104/a_1468_375# vdd 0.022331f
C10134 fanout73/a_36_113# _136_ 0.002661f
C10135 _044_ output30/a_224_472# 0.00717f
C10136 _119_ _162_ 0.036701f
C10137 FILLER_0_5_164/a_484_472# vss 0.003257f
C10138 net73 _137_ 0.047989f
C10139 _434_/a_36_151# _023_ 0.035162f
C10140 FILLER_0_17_72/a_932_472# _175_ 0.003281f
C10141 FILLER_0_5_212/a_36_472# net22 0.0015f
C10142 output9/a_224_472# net65 0.095296f
C10143 net75 fanout75/a_36_113# 0.035159f
C10144 net74 FILLER_0_11_124/a_124_375# 0.047331f
C10145 FILLER_0_19_187/a_36_472# _434_/a_36_151# 0.002398f
C10146 FILLER_0_21_286/a_124_375# net77 0.00301f
C10147 _016_ net57 0.028276f
C10148 ctln[1] FILLER_0_3_221/a_572_375# 0.001554f
C10149 _030_ FILLER_0_3_78/a_124_375# 0.010439f
C10150 net20 _014_ 0.008597f
C10151 net15 _453_/a_2665_112# 0.011775f
C10152 net69 FILLER_0_2_111/a_484_472# 0.010567f
C10153 _031_ FILLER_0_2_111/a_1468_375# 0.013595f
C10154 _076_ _059_ 1.03702f
C10155 fanout52/a_36_160# trim_val\[4\] 0.019286f
C10156 ctln[1] net5 0.050549f
C10157 _341_/a_49_472# FILLER_0_16_154/a_572_375# 0.001643f
C10158 net55 net44 0.018961f
C10159 FILLER_0_9_28/a_1916_375# _220_/a_67_603# 0.014522f
C10160 net44 _452_/a_3129_107# 0.067848f
C10161 _429_/a_36_151# FILLER_0_15_212/a_572_375# 0.059049f
C10162 fanout76/a_36_160# net4 0.002206f
C10163 net54 _211_/a_36_160# 0.001244f
C10164 _069_ FILLER_0_13_206/a_124_375# 0.009695f
C10165 FILLER_0_19_171/a_572_375# vdd 0.022516f
C10166 FILLER_0_20_15/a_1020_375# net40 0.005742f
C10167 _442_/a_3041_156# vdd 0.001178f
C10168 FILLER_0_4_123/a_124_375# _370_/a_124_24# 0.007188f
C10169 _114_ _311_/a_1920_473# 0.005579f
C10170 ctlp[5] vdd 0.293399f
C10171 FILLER_0_15_235/a_124_375# vss 0.001993f
C10172 FILLER_0_15_235/a_572_375# vdd -0.005887f
C10173 trim_val\[3\] vdd 0.211478f
C10174 FILLER_0_18_177/a_2364_375# net21 0.018463f
C10175 _415_/a_448_472# net79 0.001602f
C10176 net36 net14 0.037175f
C10177 _144_ _433_/a_1000_472# 0.029564f
C10178 FILLER_0_18_171/a_36_472# vss 0.0032f
C10179 FILLER_0_9_28/a_572_375# vdd 0.023246f
C10180 mask\[4\] net80 0.034957f
C10181 ctlp[4] result[8] 0.151286f
C10182 FILLER_0_17_200/a_124_375# vdd -0.010938f
C10183 _307_/a_234_472# _113_ 0.007518f
C10184 ctln[1] _000_ 0.223573f
C10185 output9/a_224_472# net59 0.051763f
C10186 mask\[5\] FILLER_0_18_177/a_1828_472# 0.001038f
C10187 FILLER_0_14_91/a_124_375# _095_ 0.01418f
C10188 _432_/a_2248_156# _139_ 0.002904f
C10189 _424_/a_2248_156# net36 0.017101f
C10190 FILLER_0_0_130/a_124_375# vdd 0.012493f
C10191 net20 _070_ 0.075448f
C10192 _425_/a_2560_156# vdd 0.001827f
C10193 _425_/a_2665_112# vss 0.002983f
C10194 _005_ net19 0.033451f
C10195 _253_/a_1100_68# _084_ 0.001651f
C10196 _053_ _154_ 0.41707f
C10197 FILLER_0_8_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001597f
C10198 net20 FILLER_0_12_220/a_1380_472# 0.029747f
C10199 net55 _176_ 0.300149f
C10200 net53 FILLER_0_14_107/a_1468_375# 0.001642f
C10201 net70 FILLER_0_14_107/a_932_472# 0.008396f
C10202 FILLER_0_20_98/a_124_375# vss 0.013019f
C10203 FILLER_0_20_98/a_36_472# vdd 0.095266f
C10204 FILLER_0_17_72/a_3172_472# FILLER_0_17_104/a_36_472# 0.013277f
C10205 FILLER_0_1_98/a_124_375# net14 0.049552f
C10206 FILLER_0_5_128/a_484_472# FILLER_0_5_136/a_36_472# 0.013276f
C10207 FILLER_0_8_263/a_36_472# calibrate 0.006968f
C10208 _122_ FILLER_0_6_231/a_484_472# 0.017477f
C10209 _123_ FILLER_0_6_231/a_124_375# 0.001259f
C10210 _247_/a_36_160# _090_ 0.010285f
C10211 _190_/a_36_160# _039_ 0.003926f
C10212 _050_ _436_/a_2560_156# 0.01099f
C10213 _420_/a_796_472# vss 0.001659f
C10214 result[9] _421_/a_448_472# 0.015264f
C10215 FILLER_0_3_204/a_124_375# net21 0.010054f
C10216 _143_ _137_ 0.009932f
C10217 FILLER_0_18_171/a_124_375# _143_ 0.005331f
C10218 net63 fanout63/a_36_160# 0.011149f
C10219 trim_val\[4\] _443_/a_448_472# 0.038063f
C10220 FILLER_0_14_81/a_36_472# _043_ 0.001714f
C10221 FILLER_0_24_130/a_36_472# output24/a_224_472# 0.023414f
C10222 net70 _451_/a_1353_112# 0.00194f
C10223 _115_ FILLER_0_9_105/a_124_375# 0.002316f
C10224 _320_/a_1792_472# vdd 0.001113f
C10225 net3 FILLER_0_15_2/a_484_472# 0.002224f
C10226 _109_ vdd 0.059259f
C10227 _432_/a_36_151# _141_ 0.008193f
C10228 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_36_472# 0.026657f
C10229 ctln[1] FILLER_0_1_266/a_572_375# 0.004319f
C10230 FILLER_0_9_290/a_124_375# FILLER_0_9_282/a_572_375# 0.012001f
C10231 net20 _419_/a_1000_472# 0.022734f
C10232 FILLER_0_16_241/a_124_375# _099_ 0.040547f
C10233 ctlp[1] net19 0.029153f
C10234 _130_ _327_/a_244_68# 0.00117f
C10235 ctln[4] vss 0.244634f
C10236 _093_ FILLER_0_18_139/a_36_472# 0.008761f
C10237 output23/a_224_472# _050_ 0.014495f
C10238 mask\[9\] _438_/a_1204_472# 0.03521f
C10239 _395_/a_36_488# _085_ 0.020572f
C10240 _247_/a_36_160# net22 0.048614f
C10241 FILLER_0_22_86/a_124_375# FILLER_0_23_88/a_36_472# 0.001684f
C10242 FILLER_0_3_172/a_2812_375# net22 0.013048f
C10243 FILLER_0_4_177/a_124_375# vdd 0.021637f
C10244 FILLER_0_13_142/a_1468_375# vdd 0.028002f
C10245 fanout53/a_36_160# vdd 0.016868f
C10246 FILLER_0_13_142/a_1020_375# vss 0.005307f
C10247 net57 FILLER_0_8_156/a_572_375# 0.014948f
C10248 _415_/a_2560_156# result[1] 0.002282f
C10249 FILLER_0_21_133/a_36_472# vdd 0.092168f
C10250 _417_/a_36_151# vdd 0.140703f
C10251 FILLER_0_10_256/a_36_472# _426_/a_36_151# 0.059238f
C10252 _093_ _094_ 0.003586f
C10253 _176_ net23 0.036283f
C10254 FILLER_0_16_57/a_124_375# FILLER_0_15_59/a_36_472# 0.001543f
C10255 FILLER_0_14_81/a_36_472# _175_ 0.076977f
C10256 net7 vdd 0.321735f
C10257 net79 _416_/a_2560_156# 0.013576f
C10258 FILLER_0_8_247/a_1380_472# vdd 0.036604f
C10259 _091_ mask\[3\] 0.044304f
C10260 _052_ FILLER_0_18_53/a_124_375# 0.001585f
C10261 _421_/a_2248_156# vdd 0.035239f
C10262 state\[2\] state\[1\] 0.229832f
C10263 _030_ net14 0.079892f
C10264 _053_ _058_ 0.075418f
C10265 _132_ FILLER_0_14_107/a_932_472# 0.014911f
C10266 cal_count\[3\] _408_/a_56_524# 0.001685f
C10267 FILLER_0_21_142/a_124_375# vdd 0.020936f
C10268 FILLER_0_13_65/a_36_472# net74 0.014937f
C10269 _057_ _043_ 0.02152f
C10270 _069_ FILLER_0_13_212/a_124_375# 0.070185f
C10271 net50 FILLER_0_7_59/a_36_472# 0.01018f
C10272 _422_/a_36_151# vss 0.014056f
C10273 _422_/a_448_472# vdd 0.032865f
C10274 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3260_375# 0.086635f
C10275 _378_/a_224_472# vdd 0.002263f
C10276 _067_ _389_/a_36_148# 0.002789f
C10277 net63 FILLER_0_17_218/a_484_472# 0.002672f
C10278 net44 FILLER_0_15_10/a_36_472# 0.012286f
C10279 _426_/a_1000_472# vdd 0.007031f
C10280 FILLER_0_18_100/a_36_472# FILLER_0_18_107/a_36_472# 0.002764f
C10281 _093_ FILLER_0_18_107/a_572_375# 0.008393f
C10282 _359_/a_36_488# _131_ 0.006398f
C10283 _232_/a_67_603# FILLER_0_6_47/a_36_472# 0.010206f
C10284 _165_ _377_/a_36_472# 0.025689f
C10285 _098_ FILLER_0_20_87/a_124_375# 0.019333f
C10286 FILLER_0_15_282/a_124_375# vss 0.004893f
C10287 _287_/a_36_472# mask\[2\] 0.00492f
C10288 FILLER_0_15_282/a_572_375# vdd 0.002928f
C10289 _446_/a_2248_156# net40 0.037373f
C10290 net54 _145_ 0.087336f
C10291 net36 FILLER_0_15_205/a_124_375# 0.004337f
C10292 _081_ cal_itt\[0\] 0.036569f
C10293 FILLER_0_11_101/a_572_375# vss 0.055325f
C10294 FILLER_0_11_101/a_36_472# vdd 0.093852f
C10295 mask\[5\] FILLER_0_21_206/a_124_375# 0.011644f
C10296 net25 _098_ 0.001267f
C10297 ctlp[5] _024_ 0.022549f
C10298 FILLER_0_19_47/a_484_472# _012_ 0.001667f
C10299 net63 _430_/a_2665_112# 0.075661f
C10300 net69 _441_/a_448_472# 0.028545f
C10301 _077_ _072_ 0.178678f
C10302 FILLER_0_13_65/a_36_472# cal_count\[1\] 0.016393f
C10303 _138_ mask\[1\] 0.085445f
C10304 net36 _098_ 3.387566f
C10305 net52 FILLER_0_3_142/a_36_472# 0.001122f
C10306 _003_ FILLER_0_5_181/a_36_472# 0.003545f
C10307 _447_/a_2665_112# _030_ 0.001226f
C10308 FILLER_0_4_49/a_124_375# _164_ 0.017213f
C10309 net71 _437_/a_1308_423# 0.023981f
C10310 _445_/a_36_151# net66 0.058093f
C10311 _363_/a_692_472# _086_ 0.001353f
C10312 net63 FILLER_0_15_212/a_572_375# 0.001597f
C10313 _447_/a_1000_472# _036_ 0.002902f
C10314 net66 _029_ 0.056971f
C10315 _064_ _445_/a_2248_156# 0.013127f
C10316 fanout80/a_36_113# _019_ 0.003644f
C10317 output12/a_224_472# vdd 0.106635f
C10318 FILLER_0_9_223/a_572_375# _426_/a_2665_112# 0.005202f
C10319 _408_/a_56_524# net40 0.001367f
C10320 _420_/a_36_151# net77 0.023469f
C10321 FILLER_0_18_100/a_124_375# _136_ 0.002528f
C10322 FILLER_0_5_117/a_124_375# _163_ 0.003096f
C10323 _127_ _017_ 0.005836f
C10324 ctlp[1] _009_ 0.085933f
C10325 net55 _183_ 0.024948f
C10326 _152_ vss 0.140215f
C10327 ctln[2] net9 0.022757f
C10328 net75 FILLER_0_8_247/a_1380_472# 0.020589f
C10329 result[9] FILLER_0_24_274/a_484_472# 0.003507f
C10330 _046_ _099_ 0.005245f
C10331 _028_ _154_ 0.174927f
C10332 _155_ FILLER_0_4_91/a_572_375# 0.004038f
C10333 _116_ _311_/a_2700_473# 0.001555f
C10334 FILLER_0_8_24/a_124_375# net40 0.002431f
C10335 _175_ _451_/a_3129_107# 0.021546f
C10336 FILLER_0_7_104/a_1380_472# vss 0.003236f
C10337 net58 output48/a_224_472# 0.065357f
C10338 FILLER_0_21_142/a_36_472# vss 0.009084f
C10339 FILLER_0_3_78/a_572_375# _164_ 0.055492f
C10340 FILLER_0_20_193/a_124_375# FILLER_0_19_195/a_36_472# 0.001543f
C10341 net73 FILLER_0_18_107/a_2276_472# 0.016723f
C10342 output32/a_224_472# _418_/a_36_151# 0.07368f
C10343 _081_ FILLER_0_5_148/a_124_375# 0.021583f
C10344 net75 _426_/a_1000_472# 0.002727f
C10345 _036_ _381_/a_36_472# 0.023012f
C10346 _367_/a_36_68# _156_ 0.096366f
C10347 _081_ FILLER_0_6_177/a_484_472# 0.010037f
C10348 _255_/a_224_552# _375_/a_36_68# 0.00229f
C10349 _043_ FILLER_0_13_72/a_572_375# 0.013294f
C10350 _093_ FILLER_0_18_209/a_124_375# 0.00333f
C10351 FILLER_0_2_101/a_124_375# trim_mask\[3\] 0.033692f
C10352 _074_ _312_/a_672_472# 0.005399f
C10353 FILLER_0_18_107/a_932_472# vdd 0.009633f
C10354 _308_/a_848_380# _219_/a_36_160# 0.001045f
C10355 net15 vdd 2.073988f
C10356 _420_/a_36_151# FILLER_0_23_290/a_36_472# 0.001723f
C10357 net58 net5 0.387314f
C10358 _014_ FILLER_0_7_233/a_36_472# 0.002089f
C10359 net19 FILLER_0_23_282/a_124_375# 0.001668f
C10360 _208_/a_36_160# FILLER_0_22_128/a_2812_375# 0.026361f
C10361 FILLER_0_3_204/a_36_472# vdd 0.092654f
C10362 net16 trim_val\[1\] 0.164715f
C10363 net27 FILLER_0_12_236/a_484_472# 0.042937f
C10364 _149_ _437_/a_448_472# 0.009274f
C10365 net54 FILLER_0_22_128/a_484_472# 0.055436f
C10366 FILLER_0_18_139/a_484_472# _145_ 0.002415f
C10367 _132_ net71 0.099427f
C10368 trim_val\[0\] vss 0.11063f
C10369 FILLER_0_19_55/a_124_375# FILLER_0_17_56/a_36_472# 0.001338f
C10370 FILLER_0_16_89/a_1380_472# vdd 0.010554f
C10371 _014_ vss 0.034646f
C10372 FILLER_0_12_124/a_36_472# _332_/a_36_472# 0.004546f
C10373 net15 FILLER_0_23_60/a_36_472# 0.004561f
C10374 FILLER_0_13_142/a_124_375# net23 0.003962f
C10375 net74 FILLER_0_2_127/a_36_472# 0.001261f
C10376 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_572_375# 0.001597f
C10377 _425_/a_796_472# _122_ 0.001701f
C10378 _425_/a_36_151# _123_ 0.006319f
C10379 _425_/a_1000_472# calibrate 0.027245f
C10380 _104_ _106_ 0.17237f
C10381 _323_/a_36_113# _015_ 0.003795f
C10382 net47 _066_ 0.096823f
C10383 FILLER_0_20_169/a_36_472# _098_ 0.007354f
C10384 FILLER_0_17_72/a_124_375# FILLER_0_17_64/a_124_375# 0.003732f
C10385 _003_ vss 0.095366f
C10386 net58 _000_ 0.00389f
C10387 _063_ net67 0.039144f
C10388 _011_ _422_/a_1204_472# 0.002176f
C10389 _136_ vss 0.947188f
C10390 _432_/a_1308_423# vdd 0.029938f
C10391 net73 _095_ 0.003688f
C10392 _086_ FILLER_0_6_177/a_484_472# 0.017841f
C10393 _308_/a_124_24# net14 0.005016f
C10394 _057_ _267_/a_1568_472# 0.002083f
C10395 net21 vss 1.123312f
C10396 net20 FILLER_0_3_221/a_932_472# 0.054476f
C10397 _077_ FILLER_0_9_60/a_124_375# 0.051389f
C10398 FILLER_0_10_78/a_484_472# _120_ 0.004669f
C10399 _432_/a_2665_112# net80 0.041304f
C10400 _186_ vdd 0.074983f
C10401 net56 FILLER_0_19_142/a_124_375# 0.003154f
C10402 _103_ net30 0.013544f
C10403 _250_/a_36_68# _071_ 0.199512f
C10404 _070_ FILLER_0_7_233/a_36_472# 0.07194f
C10405 _005_ _193_/a_36_160# 0.009892f
C10406 _006_ result[3] 0.016909f
C10407 _028_ _058_ 0.041158f
C10408 _229_/a_224_472# net22 0.007346f
C10409 _095_ net17 0.172789f
C10410 FILLER_0_22_177/a_36_472# mask\[6\] 0.006882f
C10411 _077_ FILLER_0_8_127/a_36_472# 0.003023f
C10412 FILLER_0_13_228/a_124_375# FILLER_0_12_220/a_1020_375# 0.05841f
C10413 net18 _416_/a_2248_156# 0.002106f
C10414 net47 net37 0.057409f
C10415 _133_ vdd 0.27652f
C10416 net15 net72 0.157843f
C10417 _070_ vss 1.363355f
C10418 _449_/a_796_472# vss 0.00143f
C10419 net81 FILLER_0_15_228/a_124_375# 0.006974f
C10420 FILLER_0_6_239/a_36_472# _074_ 0.004715f
C10421 net50 FILLER_0_6_90/a_36_472# 0.049285f
C10422 FILLER_0_12_220/a_1380_472# vss 0.006172f
C10423 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2724_472# 0.026657f
C10424 cal_count\[3\] _043_ 0.721078f
C10425 FILLER_0_18_177/a_3260_375# _205_/a_36_160# 0.001313f
C10426 _091_ FILLER_0_17_218/a_124_375# 0.013726f
C10427 cal_itt\[2\] _413_/a_2248_156# 0.002527f
C10428 net63 FILLER_0_17_200/a_36_472# 0.005648f
C10429 net55 FILLER_0_18_37/a_932_472# 0.00769f
C10430 _426_/a_3041_156# net64 0.001046f
C10431 _450_/a_1353_112# output6/a_224_472# 0.008732f
C10432 FILLER_0_17_72/a_2812_375# vdd 0.005986f
C10433 _376_/a_36_160# vdd -0.006711f
C10434 mask\[4\] _106_ 0.091207f
C10435 net10 FILLER_0_1_212/a_124_375# 0.002314f
C10436 _208_/a_36_160# _049_ 0.04568f
C10437 _009_ FILLER_0_23_282/a_124_375# 0.012402f
C10438 _127_ FILLER_0_11_135/a_124_375# 0.040456f
C10439 FILLER_0_8_247/a_1468_375# calibrate 0.006404f
C10440 fanout50/a_36_160# net50 0.052685f
C10441 _187_ _174_ 0.001321f
C10442 FILLER_0_22_86/a_1468_375# vdd 0.035441f
C10443 _105_ net32 2.08459f
C10444 net33 _434_/a_36_151# 0.002776f
C10445 _418_/a_36_151# vdd 0.155643f
C10446 _422_/a_36_151# mask\[7\] 0.043316f
C10447 net52 _443_/a_1308_423# 0.02003f
C10448 _131_ net36 0.068899f
C10449 output39/a_224_472# _033_ 0.045759f
C10450 _058_ trim_mask\[0\] 0.076069f
C10451 _426_/a_36_151# calibrate 0.004525f
C10452 _300_/a_224_472# vdd 0.001344f
C10453 net31 output18/a_224_472# 0.04975f
C10454 FILLER_0_13_206/a_124_375# net22 0.024537f
C10455 _053_ net52 0.042556f
C10456 trim_mask\[3\] net14 0.142743f
C10457 _256_/a_1164_497# net4 0.004729f
C10458 _132_ fanout71/a_36_113# 0.055078f
C10459 mask\[5\] _145_ 0.012075f
C10460 FILLER_0_16_73/a_124_375# net15 0.005202f
C10461 mask\[5\] FILLER_0_19_195/a_124_375# 0.007169f
C10462 FILLER_0_9_142/a_36_472# vss 0.004305f
C10463 _095_ _452_/a_36_151# 0.002974f
C10464 _453_/a_796_472# _042_ 0.005463f
C10465 _453_/a_1308_423# net51 0.001804f
C10466 _043_ net40 0.031043f
C10467 _402_/a_728_93# cal_count\[1\] 0.057043f
C10468 FILLER_0_16_89/a_572_375# net14 0.00106f
C10469 state\[2\] vdd 0.392508f
C10470 _326_/a_36_160# vss 0.002357f
C10471 FILLER_0_4_107/a_572_375# net47 0.006041f
C10472 cal_itt\[3\] _055_ 0.007428f
C10473 _114_ _069_ 0.029875f
C10474 net34 FILLER_0_22_128/a_2364_375# 0.009656f
C10475 net15 _441_/a_1000_472# 0.025912f
C10476 _178_ FILLER_0_15_10/a_124_375# 0.002355f
C10477 _045_ vss 0.032891f
C10478 _437_/a_2665_112# vdd 0.050182f
C10479 _185_ net40 0.048742f
C10480 _449_/a_1000_472# net72 0.001247f
C10481 _449_/a_448_472# net55 0.004439f
C10482 _420_/a_2248_156# _108_ 0.021735f
C10483 net15 _447_/a_448_472# 0.001766f
C10484 FILLER_0_8_239/a_124_375# calibrate 0.008393f
C10485 FILLER_0_4_177/a_36_472# net76 0.003007f
C10486 FILLER_0_18_2/a_3172_472# net40 0.046864f
C10487 FILLER_0_4_213/a_484_472# vss 0.007857f
C10488 fanout59/a_36_160# vdd 0.02169f
C10489 net63 _434_/a_448_472# 0.008139f
C10490 FILLER_0_7_72/a_36_472# _439_/a_36_151# 0.013806f
C10491 net55 FILLER_0_17_72/a_1468_375# 0.014449f
C10492 ctlp[8] net35 0.001859f
C10493 _020_ _431_/a_796_472# 0.012284f
C10494 _131_ FILLER_0_14_123/a_124_375# 0.016964f
C10495 _446_/a_1204_472# net66 0.001885f
C10496 _305_/a_36_159# _425_/a_36_151# 0.001404f
C10497 net15 _439_/a_796_472# 0.001822f
C10498 net47 FILLER_0_5_148/a_484_472# 0.009741f
C10499 _192_/a_67_603# vss 0.007021f
C10500 trim_mask\[4\] vdd 0.20602f
C10501 net80 _140_ 0.188514f
C10502 _096_ _161_ 0.00104f
C10503 FILLER_0_5_72/a_572_375# net49 0.001158f
C10504 _062_ _226_/a_276_68# 0.001286f
C10505 _273_/a_36_68# _223_/a_36_160# 0.002786f
C10506 net54 _433_/a_2560_156# 0.014333f
C10507 FILLER_0_23_44/a_1380_472# vss 0.003905f
C10508 _077_ _453_/a_2665_112# 0.002824f
C10509 en_co_clk FILLER_0_13_100/a_124_375# 0.002325f
C10510 FILLER_0_19_47/a_572_375# _052_ 0.020156f
C10511 FILLER_0_21_125/a_484_472# vss 0.002399f
C10512 FILLER_0_11_78/a_36_472# vdd -0.001328f
C10513 FILLER_0_11_78/a_572_375# vss 0.004808f
C10514 FILLER_0_20_193/a_484_472# _098_ 0.012457f
C10515 FILLER_0_5_109/a_484_472# _160_ 0.001598f
C10516 FILLER_0_5_72/a_932_472# _029_ 0.007801f
C10517 FILLER_0_5_72/a_1468_375# trim_mask\[1\] 0.017105f
C10518 FILLER_0_6_47/a_2364_375# vdd 0.015888f
C10519 FILLER_0_6_47/a_1916_375# vss 0.005279f
C10520 FILLER_0_21_133/a_36_472# _433_/a_36_151# 0.001723f
C10521 net26 _423_/a_1000_472# 0.001338f
C10522 FILLER_0_24_130/a_124_375# net54 0.001269f
C10523 _305_/a_36_159# net1 0.013619f
C10524 _444_/a_448_472# _054_ 0.017318f
C10525 _411_/a_2665_112# vdd 0.026095f
C10526 FILLER_0_18_171/a_36_472# _141_ 0.002037f
C10527 FILLER_0_12_50/a_36_472# vss 0.0027f
C10528 _412_/a_796_472# net81 0.038712f
C10529 net43 vdd 0.210686f
C10530 _086_ _055_ 0.113385f
C10531 output44/a_224_472# vdd 0.043902f
C10532 FILLER_0_17_218/a_572_375# _069_ 0.001464f
C10533 FILLER_0_7_104/a_932_472# _154_ 0.002023f
C10534 _422_/a_796_472# _108_ 0.007356f
C10535 _021_ vss 0.142648f
C10536 _115_ FILLER_0_10_107/a_36_472# 0.016715f
C10537 _098_ FILLER_0_16_154/a_1468_375# 0.009042f
C10538 net10 ctln[3] 0.873575f
C10539 _419_/a_448_472# net77 0.007659f
C10540 net27 result[1] 0.187252f
C10541 net54 FILLER_0_18_107/a_124_375# 0.001636f
C10542 _431_/a_1000_472# net36 0.001771f
C10543 _075_ _053_ 0.634359f
C10544 net41 _446_/a_1000_472# 0.01097f
C10545 ctln[3] FILLER_0_0_232/a_124_375# 0.012394f
C10546 net49 _160_ 1.243817f
C10547 mask\[7\] net21 0.050718f
C10548 FILLER_0_23_282/a_36_472# vdd 0.106034f
C10549 FILLER_0_23_282/a_572_375# vss 0.058599f
C10550 _322_/a_1084_68# _128_ 0.002629f
C10551 _023_ mask\[6\] 0.077441f
C10552 FILLER_0_11_101/a_124_375# _058_ 0.002209f
C10553 FILLER_0_24_63/a_124_375# vdd 0.029514f
C10554 valid cal_itt\[1\] 0.011576f
C10555 FILLER_0_21_28/a_2724_472# _012_ 0.020109f
C10556 net68 _160_ 0.072339f
C10557 _075_ _414_/a_2560_156# 0.026328f
C10558 net73 net74 0.016949f
C10559 _086_ _154_ 0.102849f
C10560 _320_/a_1568_472# net79 0.001157f
C10561 trimb[4] net17 0.004628f
C10562 _445_/a_796_472# _034_ 0.009261f
C10563 _433_/a_1308_423# _022_ 0.015376f
C10564 fanout69/a_36_113# vdd 0.00378f
C10565 _408_/a_728_93# _067_ 0.006262f
C10566 FILLER_0_12_136/a_932_472# _127_ 0.002804f
C10567 FILLER_0_2_93/a_484_472# vdd 0.005163f
C10568 _057_ _062_ 0.062063f
C10569 cal_itt\[3\] _058_ 0.002207f
C10570 net41 _408_/a_1336_472# 0.063099f
C10571 _411_/a_2665_112# net75 0.005223f
C10572 _119_ _154_ 0.01697f
C10573 _119_ _313_/a_67_603# 0.015457f
C10574 _437_/a_448_472# net14 0.090442f
C10575 _448_/a_2248_156# vdd 0.008296f
C10576 valid sample 0.103192f
C10577 _028_ net52 0.150861f
C10578 _099_ FILLER_0_15_235/a_572_375# 0.001327f
C10579 _178_ _278_/a_36_160# 0.269109f
C10580 _176_ FILLER_0_15_72/a_36_472# 0.002101f
C10581 FILLER_0_14_107/a_484_472# vss -0.001894f
C10582 FILLER_0_14_107/a_932_472# vdd 0.006908f
C10583 _051_ net71 0.001617f
C10584 _115_ FILLER_0_10_94/a_124_375# 0.010311f
C10585 net4 _070_ 0.169392f
C10586 valid vss 0.308766f
C10587 FILLER_0_22_177/a_484_472# vss -0.001894f
C10588 FILLER_0_22_177/a_932_472# vdd 0.029547f
C10589 _087_ net76 0.529571f
C10590 _043_ FILLER_0_13_80/a_124_375# 0.013485f
C10591 FILLER_0_22_177/a_124_375# _435_/a_36_151# 0.059049f
C10592 net58 _412_/a_2665_112# 0.006815f
C10593 net4 FILLER_0_12_220/a_1380_472# 0.016375f
C10594 net66 FILLER_0_5_54/a_484_472# 0.001863f
C10595 _423_/a_36_151# FILLER_0_23_44/a_36_472# 0.001723f
C10596 FILLER_0_12_136/a_124_375# cal_count\[3\] 0.005006f
C10597 FILLER_0_3_221/a_932_472# vss 0.002881f
C10598 FILLER_0_3_221/a_1380_472# vdd 0.003819f
C10599 FILLER_0_7_104/a_932_472# _058_ 0.002096f
C10600 _394_/a_1336_472# _175_ 0.002792f
C10601 net36 FILLER_0_15_212/a_932_472# 0.008239f
C10602 _076_ _311_/a_66_473# 0.003077f
C10603 FILLER_0_15_116/a_572_375# net36 0.007321f
C10604 _427_/a_1308_423# _095_ 0.022677f
C10605 net68 FILLER_0_5_54/a_1020_375# 0.00648f
C10606 _415_/a_2560_156# net27 0.008433f
C10607 net41 _034_ 0.026084f
C10608 net9 cal_itt\[1\] 0.028339f
C10609 _081_ FILLER_0_5_198/a_572_375# 0.001285f
C10610 _091_ _333_/a_36_160# 0.031262f
C10611 _451_/a_1353_112# vdd 0.009693f
C10612 _250_/a_36_68# net23 0.002628f
C10613 _032_ net23 0.019676f
C10614 FILLER_0_5_54/a_36_472# trim_mask\[1\] 0.101342f
C10615 FILLER_0_5_54/a_1380_472# _029_ 0.01027f
C10616 FILLER_0_10_256/a_124_375# net19 0.002884f
C10617 FILLER_0_24_130/a_36_472# vss 0.001687f
C10618 _441_/a_36_151# _440_/a_1308_423# 0.001736f
C10619 net61 _419_/a_36_151# 0.019141f
C10620 net60 output18/a_224_472# 0.001518f
C10621 net79 FILLER_0_15_282/a_124_375# 0.001058f
C10622 FILLER_0_9_270/a_484_472# FILLER_0_9_282/a_36_472# 0.002296f
C10623 _137_ _334_/a_36_160# 0.015722f
C10624 FILLER_0_16_89/a_1468_375# _040_ 0.004985f
C10625 _374_/a_244_472# _076_ 0.001567f
C10626 _161_ FILLER_0_6_177/a_484_472# 0.001723f
C10627 _128_ _247_/a_36_160# 0.00163f
C10628 _027_ FILLER_0_18_76/a_484_472# 0.00705f
C10629 mask\[1\] FILLER_0_15_228/a_124_375# 0.013558f
C10630 _048_ vdd 0.270091f
C10631 _086_ _058_ 0.054155f
C10632 _429_/a_2665_112# _043_ 0.007641f
C10633 fanout74/a_36_113# _032_ 0.012909f
C10634 _069_ _085_ 0.032519f
C10635 FILLER_0_18_177/a_484_472# vdd 0.006177f
C10636 FILLER_0_18_177/a_36_472# vss 0.002187f
C10637 net15 FILLER_0_7_59/a_484_472# 0.015199f
C10638 _430_/a_36_151# net63 0.026607f
C10639 _115_ _322_/a_848_380# 0.011372f
C10640 _086_ _315_/a_36_68# 0.003329f
C10641 net9 vss 0.086497f
C10642 _122_ net47 0.030693f
C10643 net62 net19 0.352148f
C10644 _119_ _058_ 0.692466f
C10645 _069_ _018_ 0.002777f
C10646 _245_/a_234_472# net47 0.00188f
C10647 _136_ _337_/a_257_69# 0.002933f
C10648 net16 _447_/a_36_151# 0.133348f
C10649 FILLER_0_15_142/a_124_375# net53 0.033224f
C10650 FILLER_0_16_57/a_572_375# vdd 0.004039f
C10651 FILLER_0_16_57/a_124_375# vss 0.001678f
C10652 _440_/a_36_151# FILLER_0_6_47/a_2276_472# 0.001512f
C10653 FILLER_0_9_142/a_124_375# _313_/a_67_603# 0.029786f
C10654 _072_ _061_ 0.448032f
C10655 mask\[5\] _202_/a_36_160# 0.00164f
C10656 FILLER_0_3_2/a_36_472# net66 0.011419f
C10657 fanout68/a_36_113# _441_/a_36_151# 0.138322f
C10658 _074_ _163_ 0.446493f
C10659 FILLER_0_11_124/a_36_472# _135_ 0.110114f
C10660 FILLER_0_21_150/a_124_375# vdd 0.020581f
C10661 _002_ _079_ 0.051048f
C10662 FILLER_0_18_177/a_1468_375# _139_ 0.001359f
C10663 FILLER_0_5_198/a_124_375# net21 0.029659f
C10664 FILLER_0_21_125/a_484_472# mask\[7\] 0.003404f
C10665 net71 vdd 0.775031f
C10666 _444_/a_2560_156# net67 0.012781f
C10667 net53 _427_/a_2665_112# 0.042564f
C10668 _181_ _184_ 0.022711f
C10669 FILLER_0_1_204/a_36_472# net11 0.014707f
C10670 output38/a_224_472# trim[0] 0.026911f
C10671 FILLER_0_5_72/a_1468_375# _164_ 0.040819f
C10672 _019_ _138_ 0.003734f
C10673 _066_ _385_/a_36_68# 0.001405f
C10674 net36 _137_ 0.048198f
C10675 FILLER_0_12_2/a_36_472# output6/a_224_472# 0.00108f
C10676 _339_/a_36_160# FILLER_0_19_155/a_572_375# 0.003589f
C10677 trimb[1] FILLER_0_19_28/a_124_375# 0.00285f
C10678 FILLER_0_12_124/a_124_375# _428_/a_36_151# 0.058722f
C10679 FILLER_0_24_290/a_124_375# vdd 0.026739f
C10680 mask\[4\] _144_ 0.268823f
C10681 FILLER_0_6_239/a_124_375# _316_/a_124_24# 0.003524f
C10682 FILLER_0_20_87/a_36_472# _438_/a_448_472# 0.004782f
C10683 _077_ vdd 1.61568f
C10684 _015_ _426_/a_36_151# 0.01243f
C10685 _063_ trim_val\[1\] 0.038045f
C10686 FILLER_0_2_93/a_124_375# _441_/a_2665_112# 0.006271f
C10687 trim_mask\[2\] FILLER_0_2_93/a_36_472# 0.281054f
C10688 _033_ net40 0.298492f
C10689 _098_ _437_/a_448_472# 0.050691f
C10690 output32/a_224_472# result[9] 0.047198f
C10691 FILLER_0_5_212/a_124_375# FILLER_0_5_206/a_124_375# 0.005439f
C10692 FILLER_0_12_124/a_124_375# _114_ 0.006974f
C10693 FILLER_0_7_104/a_1020_375# _131_ 0.016404f
C10694 net65 result[0] 0.011634f
C10695 FILLER_0_5_181/a_124_375# net37 0.005396f
C10696 net80 _435_/a_36_151# 0.035259f
C10697 net36 _438_/a_1308_423# 0.012976f
C10698 _106_ _008_ 0.034748f
C10699 _277_/a_36_160# _103_ 0.032112f
C10700 FILLER_0_9_223/a_484_472# _076_ 0.001736f
C10701 _389_/a_36_148# FILLER_0_10_94/a_36_472# 0.001723f
C10702 net79 _136_ 0.00111f
C10703 cal_count\[3\] _062_ 0.004405f
C10704 fanout81/a_36_160# fanout76/a_36_160# 0.01081f
C10705 FILLER_0_16_57/a_572_375# net72 0.012909f
C10706 net79 net21 0.645949f
C10707 _385_/a_36_68# net37 0.047762f
C10708 _449_/a_36_151# _174_ 0.002252f
C10709 FILLER_0_19_55/a_36_472# _012_ 0.001667f
C10710 _256_/a_36_68# net20 0.02797f
C10711 FILLER_0_11_142/a_124_375# vdd 0.010672f
C10712 ctln[4] FILLER_0_1_212/a_124_375# 0.008197f
C10713 _327_/a_36_472# _127_ 0.002934f
C10714 result[9] _010_ 0.121471f
C10715 _303_/a_36_472# mask\[9\] 0.013976f
C10716 _076_ _080_ 0.005433f
C10717 _131_ FILLER_0_18_37/a_1468_375# 0.001151f
C10718 output48/a_224_472# net82 0.048965f
C10719 _015_ FILLER_0_8_239/a_124_375# 0.007342f
C10720 _013_ vdd 0.372605f
C10721 output44/a_224_472# FILLER_0_18_2/a_572_375# 0.001296f
C10722 net20 _429_/a_1308_423# 0.001186f
C10723 FILLER_0_16_89/a_572_375# _131_ 0.012481f
C10724 net81 FILLER_0_14_235/a_572_375# 0.029643f
C10725 _079_ _078_ 0.03338f
C10726 FILLER_0_9_142/a_124_375# _315_/a_36_68# 0.028077f
C10727 FILLER_0_9_28/a_2276_472# _453_/a_36_151# 0.059367f
C10728 _114_ FILLER_0_11_101/a_484_472# 0.025975f
C10729 FILLER_0_16_73/a_572_375# net55 0.015207f
C10730 _114_ _090_ 0.001909f
C10731 FILLER_0_3_78/a_124_375# _168_ 0.009374f
C10732 _431_/a_1308_423# _020_ 0.001997f
C10733 net82 FILLER_0_3_221/a_572_375# 0.005424f
C10734 net80 _139_ 0.178583f
C10735 FILLER_0_5_109/a_36_472# _365_/a_36_68# 0.07596f
C10736 FILLER_0_7_72/a_572_375# FILLER_0_5_72/a_484_472# 0.001512f
C10737 _074_ FILLER_0_6_231/a_124_375# 0.006087f
C10738 _444_/a_2248_156# FILLER_0_8_37/a_484_472# 0.013656f
C10739 net79 _070_ 0.009715f
C10740 FILLER_0_7_146/a_124_375# _133_ 0.001577f
C10741 FILLER_0_17_200/a_572_375# _069_ 0.011239f
C10742 _066_ vdd 0.14893f
C10743 net79 FILLER_0_12_220/a_1380_472# 0.010583f
C10744 fanout77/a_36_113# net18 0.060158f
C10745 FILLER_0_19_187/a_484_472# vss 0.004504f
C10746 ctlp[9] vss 0.013018f
C10747 net62 fanout78/a_36_113# 0.014177f
C10748 FILLER_0_7_195/a_124_375# _074_ 0.019559f
C10749 FILLER_0_1_192/a_124_375# vss 0.049811f
C10750 FILLER_0_1_192/a_36_472# vdd 0.011806f
C10751 _140_ FILLER_0_22_128/a_124_375# 0.011452f
C10752 FILLER_0_18_2/a_2364_375# _452_/a_1353_112# 0.001068f
C10753 FILLER_0_16_241/a_36_472# mask\[2\] 0.025337f
C10754 output36/a_224_472# result[9] 0.059164f
C10755 mask\[5\] _107_ 0.01249f
C10756 _430_/a_2560_156# _091_ 0.047345f
C10757 trim[0] vdd 0.125774f
C10758 _161_ _055_ 0.078364f
C10759 FILLER_0_16_73/a_484_472# vss 0.007212f
C10760 net65 output37/a_224_472# 0.096416f
C10761 FILLER_0_9_28/a_2364_375# _042_ 0.001216f
C10762 _405_/a_255_603# cal_count\[2\] 0.001576f
C10763 net58 en 0.029072f
C10764 _000_ net82 0.032846f
C10765 _432_/a_2248_156# _137_ 0.001775f
C10766 net23 mask\[6\] 0.025699f
C10767 FILLER_0_21_28/a_2812_375# vdd -0.014642f
C10768 fanout71/a_36_113# vdd 0.028178f
C10769 FILLER_0_3_172/a_1828_472# vdd 0.0083f
C10770 _414_/a_36_151# vss 0.002101f
C10771 _255_/a_224_552# _311_/a_66_473# 0.002588f
C10772 _442_/a_448_472# FILLER_0_2_127/a_36_472# 0.008634f
C10773 FILLER_0_4_197/a_572_375# net76 0.006026f
C10774 FILLER_0_8_2/a_124_375# vdd 0.016103f
C10775 _427_/a_1308_423# net74 0.005627f
C10776 _413_/a_448_472# _002_ 0.044695f
C10777 net4 FILLER_0_3_221/a_932_472# 0.002116f
C10778 _438_/a_2560_156# net14 0.049389f
C10779 _115_ _124_ 0.045023f
C10780 FILLER_0_5_54/a_36_472# _164_ 0.003923f
C10781 output27/a_224_472# FILLER_0_8_263/a_36_472# 0.002002f
C10782 cal_itt\[1\] _084_ 0.495918f
C10783 net56 net36 0.772486f
C10784 FILLER_0_4_152/a_36_472# trim_mask\[4\] 0.011746f
C10785 _069_ _310_/a_49_472# 0.023925f
C10786 _001_ net59 0.001439f
C10787 net37 vdd 0.544653f
C10788 FILLER_0_22_177/a_1468_375# net33 0.017455f
C10789 _053_ _152_ 0.032961f
C10790 net25 _213_/a_67_603# 0.027452f
C10791 net57 FILLER_0_16_154/a_1020_375# 0.001902f
C10792 _161_ _311_/a_1212_473# 0.004138f
C10793 _111_ net55 0.002855f
C10794 _013_ net72 0.006579f
C10795 _157_ vdd 0.419501f
C10796 net69 _030_ 0.49547f
C10797 FILLER_0_17_72/a_124_375# _131_ 0.006224f
C10798 _005_ _416_/a_2560_156# 0.004273f
C10799 _442_/a_796_472# _031_ 0.013039f
C10800 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1380_472# 0.003468f
C10801 net48 _056_ 0.001581f
C10802 _178_ _406_/a_36_159# 0.007052f
C10803 net20 calibrate 0.044792f
C10804 result[9] vdd 0.597071f
C10805 FILLER_0_5_72/a_572_375# net47 0.006974f
C10806 result[6] FILLER_0_21_286/a_124_375# 0.019179f
C10807 FILLER_0_3_142/a_124_375# trim_mask\[4\] 0.002514f
C10808 output37/a_224_472# net59 0.001014f
C10809 net81 net36 0.030215f
C10810 fanout75/a_36_113# _082_ 0.016843f
C10811 output34/a_224_472# ctlp[1] 0.00277f
C10812 _162_ _056_ 0.018616f
C10813 FILLER_0_2_177/a_124_375# net22 0.001318f
C10814 _084_ vss 0.082779f
C10815 FILLER_0_10_256/a_36_472# vss 0.001792f
C10816 _074_ _073_ 0.040339f
C10817 net80 FILLER_0_17_161/a_124_375# 0.021914f
C10818 net4 net9 0.008183f
C10819 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_484_472# 0.013276f
C10820 _053_ trim_val\[0\] 0.446477f
C10821 net22 _435_/a_2560_156# 0.002281f
C10822 mask\[0\] _429_/a_2560_156# 0.010913f
C10823 _091_ _072_ 0.162027f
C10824 net79 _192_/a_67_603# 0.017688f
C10825 FILLER_0_4_107/a_1380_472# FILLER_0_2_111/a_1020_375# 0.001512f
C10826 FILLER_0_0_266/a_124_375# vdd 0.006328f
C10827 _321_/a_3126_472# _124_ 0.001072f
C10828 net24 FILLER_0_22_86/a_1468_375# 0.008075f
C10829 FILLER_0_12_136/a_932_472# net23 0.004375f
C10830 _179_ vdd 0.049022f
C10831 net62 _193_/a_36_160# 0.00227f
C10832 _411_/a_2248_156# ctln[1] 0.013381f
C10833 net19 net33 0.254336f
C10834 ctln[4] ctln[3] 0.073214f
C10835 net16 _444_/a_448_472# 0.038803f
C10836 _053_ _003_ 0.021223f
C10837 _077_ _439_/a_796_472# 0.007471f
C10838 FILLER_0_4_107/a_124_375# vss 0.00322f
C10839 FILLER_0_4_107/a_572_375# vdd 0.034678f
C10840 net75 net37 0.07785f
C10841 _103_ _418_/a_2665_112# 0.0066f
C10842 _009_ FILLER_0_23_290/a_124_375# 0.002666f
C10843 result[0] result[1] 0.06045f
C10844 _075_ cal_itt\[3\] 0.731221f
C10845 _207_/a_67_603# _146_ 0.026192f
C10846 net33 mask\[6\] 0.881813f
C10847 FILLER_0_9_105/a_572_375# FILLER_0_10_107/a_484_472# 0.001543f
C10848 _013_ _424_/a_36_151# 0.012928f
C10849 _053_ net21 0.036284f
C10850 FILLER_0_9_72/a_124_375# _439_/a_36_151# 0.059049f
C10851 _114_ _076_ 0.088609f
C10852 ctlp[2] _422_/a_36_151# 0.068086f
C10853 net67 _190_/a_36_160# 0.023989f
C10854 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1468_375# 0.086742f
C10855 FILLER_0_3_54/a_36_472# _381_/a_36_472# 0.010679f
C10856 net47 _160_ 0.2966f
C10857 _016_ cal_count\[3\] 0.004588f
C10858 _061_ state\[1\] 0.02716f
C10859 _093_ FILLER_0_17_72/a_1828_472# 0.053526f
C10860 net57 _390_/a_36_68# 0.001112f
C10861 _075_ _081_ 0.001195f
C10862 FILLER_0_9_28/a_1916_375# net51 0.001008f
C10863 vss FILLER_0_5_148/a_36_472# 0.029152f
C10864 output31/a_224_472# FILLER_0_17_282/a_124_375# 0.002977f
C10865 net7 _239_/a_36_160# 0.068281f
C10866 _161_ _058_ 0.101968f
C10867 _116_ _248_/a_36_68# 0.007314f
C10868 net50 FILLER_0_8_37/a_484_472# 0.003311f
C10869 _077_ cal_count\[0\] 0.018501f
C10870 _053_ _070_ 2.345795f
C10871 net15 _394_/a_1936_472# 0.001592f
C10872 fanout52/a_36_160# trim_mask\[4\] 0.014356f
C10873 _021_ _141_ 0.047816f
C10874 _230_/a_244_68# _056_ 0.001844f
C10875 net20 FILLER_0_13_212/a_484_472# 0.001273f
C10876 _447_/a_2665_112# _168_ 0.001107f
C10877 _192_/a_67_603# _416_/a_2665_112# 0.012638f
C10878 _044_ _416_/a_36_151# 0.032206f
C10879 net55 fanout55/a_36_160# 0.028425f
C10880 _052_ FILLER_0_19_28/a_572_375# 0.011078f
C10881 _140_ _436_/a_36_151# 0.031519f
C10882 FILLER_0_7_72/a_3172_472# vdd 0.003913f
C10883 _408_/a_56_524# _043_ 0.10151f
C10884 net73 _145_ 0.009144f
C10885 _430_/a_796_472# _019_ 0.006511f
C10886 _428_/a_1000_472# _017_ 0.012268f
C10887 _345_/a_36_160# FILLER_0_19_111/a_572_375# 0.132282f
C10888 _085_ _090_ 0.001012f
C10889 _116_ _060_ 0.020653f
C10890 FILLER_0_21_28/a_2812_375# _424_/a_36_151# 0.059049f
C10891 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_484_472# 0.001963f
C10892 FILLER_0_19_155/a_572_375# vss 0.004538f
C10893 fanout51/a_36_113# net51 0.013081f
C10894 net72 _179_ 0.083699f
C10895 net76 net2 0.039533f
C10896 FILLER_0_5_54/a_1020_375# net47 0.005159f
C10897 output46/a_224_472# net43 0.10562f
C10898 net14 FILLER_0_4_91/a_572_375# 0.047331f
C10899 _408_/a_56_524# _185_ 0.002484f
C10900 output46/a_224_472# output44/a_224_472# 0.005749f
C10901 _071_ _055_ 0.002641f
C10902 _077_ _374_/a_36_68# 0.012411f
C10903 FILLER_0_0_198/a_124_375# vss 0.017602f
C10904 FILLER_0_0_198/a_36_472# vdd 0.052226f
C10905 net82 FILLER_0_3_172/a_2812_375# 0.010439f
C10906 en_co_clk vdd 0.245319f
C10907 cal_itt\[3\] FILLER_0_5_164/a_484_472# 0.001518f
C10908 _273_/a_36_68# state\[0\] 0.012187f
C10909 cal_itt\[2\] _074_ 0.082824f
C10910 output28/a_224_472# vss -0.0033f
C10911 _412_/a_448_472# net76 0.026446f
C10912 _110_ vdd 0.041979f
C10913 net20 FILLER_0_16_241/a_36_472# 0.001528f
C10914 net18 _419_/a_1308_423# 0.013637f
C10915 _137_ FILLER_0_16_154/a_1468_375# 0.014214f
C10916 _074_ net1 0.128466f
C10917 net64 FILLER_0_11_282/a_124_375# 0.023042f
C10918 _081_ FILLER_0_5_164/a_484_472# 0.001105f
C10919 _095_ net36 0.127549f
C10920 net71 _436_/a_448_472# 0.005274f
C10921 ctlp[4] _107_ 0.080312f
C10922 FILLER_0_5_109/a_36_472# _154_ 0.070958f
C10923 _415_/a_36_151# net28 0.001195f
C10924 net80 _098_ 1.289178f
C10925 FILLER_0_10_78/a_572_375# cal_count\[3\] 0.002314f
C10926 FILLER_0_7_72/a_1916_375# net50 0.059471f
C10927 _256_/a_36_68# vss 0.055568f
C10928 FILLER_0_15_150/a_124_375# _427_/a_36_151# 0.001822f
C10929 mask\[4\] FILLER_0_22_128/a_3172_472# 0.001484f
C10930 _122_ FILLER_0_5_181/a_124_375# 0.001352f
C10931 net81 _425_/a_1308_423# 0.004202f
C10932 _050_ _352_/a_49_472# 0.005393f
C10933 _134_ net14 0.001303f
C10934 net71 _433_/a_36_151# 0.014126f
C10935 _359_/a_36_488# net74 0.037211f
C10936 net77 vss 0.327705f
C10937 _018_ net22 0.141743f
C10938 net64 FILLER_0_14_235/a_572_375# 0.008689f
C10939 _429_/a_1308_423# vss 0.008906f
C10940 _423_/a_36_151# vss 0.012999f
C10941 _423_/a_448_472# vdd 0.01351f
C10942 _056_ _373_/a_244_68# 0.00229f
C10943 FILLER_0_7_72/a_932_472# net50 0.074005f
C10944 net35 _050_ 0.28822f
C10945 net15 _176_ 0.038396f
C10946 _093_ FILLER_0_16_115/a_36_472# 0.001526f
C10947 net38 FILLER_0_15_10/a_124_375# 0.047331f
C10948 _122_ _385_/a_36_68# 0.003549f
C10949 _096_ _056_ 0.001946f
C10950 FILLER_0_18_2/a_2812_375# net17 0.012909f
C10951 FILLER_0_17_72/a_484_472# net36 0.001629f
C10952 FILLER_0_10_214/a_36_472# _055_ 0.027657f
C10953 net52 FILLER_0_11_78/a_124_375# 0.006273f
C10954 FILLER_0_8_127/a_124_375# _058_ 0.007791f
C10955 _372_/a_170_472# _059_ 0.033956f
C10956 ctlp[1] FILLER_0_21_286/a_484_472# 0.045536f
C10957 net13 vdd 0.264116f
C10958 output27/a_224_472# fanout65/a_36_113# 0.011564f
C10959 FILLER_0_22_128/a_2812_375# vdd 0.003766f
C10960 FILLER_0_22_128/a_2364_375# vss 0.017496f
C10961 _069_ mask\[2\] 0.032781f
C10962 FILLER_0_20_107/a_124_375# vss 0.002749f
C10963 FILLER_0_20_107/a_36_472# vdd 0.117841f
C10964 _095_ FILLER_0_14_123/a_124_375# 0.014486f
C10965 _415_/a_1000_472# vdd 0.002497f
C10966 FILLER_0_23_290/a_36_472# vss 0.0074f
C10967 _424_/a_1204_472# vdd 0.001573f
C10968 fanout80/a_36_113# mask\[0\] 0.002212f
C10969 result[6] _420_/a_36_151# 0.011901f
C10970 _441_/a_2560_156# vss 0.001374f
C10971 _064_ vss 0.228443f
C10972 mask\[5\] FILLER_0_20_177/a_36_472# 0.017871f
C10973 net29 mask\[2\] 0.122202f
C10974 output29/a_224_472# _045_ 0.002303f
C10975 output15/a_224_472# trim_val\[3\] 0.042209f
C10976 net69 trim_mask\[3\] 0.017779f
C10977 net15 _036_ 0.036489f
C10978 _053_ FILLER_0_6_47/a_1916_375# 0.008103f
C10979 _228_/a_36_68# vss 0.031389f
C10980 mask\[3\] FILLER_0_18_177/a_1380_472# 0.005654f
C10981 _447_/a_2248_156# vdd 0.009094f
C10982 net47 _170_ 0.010131f
C10983 _117_ _060_ 0.149558f
C10984 net23 FILLER_0_5_148/a_124_375# 0.01836f
C10985 FILLER_0_8_107/a_124_375# _058_ 0.01823f
C10986 _320_/a_36_472# _113_ 0.030365f
C10987 _077_ FILLER_0_7_59/a_484_472# 0.001371f
C10988 vss output41/a_224_472# -0.007739f
C10989 net63 FILLER_0_19_187/a_36_472# 0.006753f
C10990 result[2] result[3] 0.09741f
C10991 _439_/a_2665_112# vss 0.003954f
C10992 _104_ _421_/a_1308_423# 0.001621f
C10993 net4 _084_ 0.029194f
C10994 _445_/a_36_151# net17 0.009838f
C10995 _345_/a_36_160# vss 0.003697f
C10996 FILLER_0_17_56/a_36_472# FILLER_0_18_53/a_484_472# 0.026657f
C10997 FILLER_0_15_116/a_124_375# net70 0.02416f
C10998 fanout49/a_36_160# net49 0.032999f
C10999 fanout66/a_36_113# _160_ 0.015681f
C11000 input4/a_36_68# net59 0.003625f
C11001 _181_ _402_/a_718_527# 0.00461f
C11002 calibrate FILLER_0_7_233/a_36_472# 0.013262f
C11003 mask\[2\] FILLER_0_15_212/a_36_472# 0.001181f
C11004 FILLER_0_9_223/a_484_472# _128_ 0.005152f
C11005 mask\[9\] FILLER_0_18_76/a_484_472# 0.002672f
C11006 sample calibrate 0.001861f
C11007 trim_val\[4\] FILLER_0_3_172/a_484_472# 0.002633f
C11008 FILLER_0_10_37/a_124_375# _453_/a_36_151# 0.017882f
C11009 FILLER_0_13_65/a_124_375# net15 0.048002f
C11010 trim_val\[4\] _386_/a_848_380# 0.007605f
C11011 output42/a_224_472# net6 0.010571f
C11012 net78 _108_ 0.056528f
C11013 mask\[9\] _423_/a_2665_112# 0.001735f
C11014 _144_ _140_ 0.415736f
C11015 FILLER_0_18_2/a_2812_375# _452_/a_36_151# 0.001597f
C11016 _130_ FILLER_0_12_136/a_36_472# 0.082451f
C11017 FILLER_0_17_72/a_932_472# FILLER_0_18_76/a_484_472# 0.05841f
C11018 net56 FILLER_0_18_139/a_1380_472# 0.048069f
C11019 calibrate vss 1.140031f
C11020 _122_ vdd 0.379907f
C11021 _428_/a_448_472# FILLER_0_14_107/a_932_472# 0.007f
C11022 result[6] _421_/a_1308_423# 0.023269f
C11023 FILLER_0_9_28/a_2724_472# _453_/a_448_472# 0.008036f
C11024 net61 vdd 0.46584f
C11025 fanout60/a_36_160# net62 0.049222f
C11026 net64 net36 0.037523f
C11027 fanout53/a_36_160# FILLER_0_16_154/a_932_472# 0.001426f
C11028 net52 FILLER_0_2_93/a_572_375# 0.007787f
C11029 _147_ _207_/a_67_603# 0.001123f
C11030 net58 _411_/a_2248_156# 0.014884f
C11031 _255_/a_224_552# _114_ 0.005131f
C11032 FILLER_0_17_200/a_36_472# net21 0.036768f
C11033 mask\[5\] FILLER_0_19_171/a_932_472# 0.007596f
C11034 FILLER_0_17_72/a_3172_472# net14 0.046864f
C11035 net36 mask\[1\] 0.28584f
C11036 net41 _052_ 0.001927f
C11037 _188_ _042_ 0.015684f
C11038 output32/a_224_472# output31/a_224_472# 0.00289f
C11039 _092_ _091_ 0.028594f
C11040 net55 _424_/a_1308_423# 0.00168f
C11041 FILLER_0_6_239/a_124_375# FILLER_0_6_231/a_572_375# 0.012001f
C11042 FILLER_0_17_200/a_572_375# net22 0.047331f
C11043 input1/a_36_113# vdd 0.099655f
C11044 _246_/a_36_68# _055_ 0.028938f
C11045 _311_/a_2180_473# vdd 0.001974f
C11046 fanout71/a_36_113# _433_/a_36_151# 0.138322f
C11047 ctln[6] net23 0.003826f
C11048 _096_ FILLER_0_12_196/a_124_375# 0.002309f
C11049 FILLER_0_19_142/a_124_375# _145_ 0.009109f
C11050 FILLER_0_5_128/a_572_375# _163_ 0.007391f
C11051 _049_ vdd 0.199608f
C11052 net31 _291_/a_36_160# 0.005683f
C11053 net5 clk 0.042578f
C11054 _153_ vss 0.256017f
C11055 fanout54/a_36_160# vdd 0.008482f
C11056 _310_/a_49_472# _090_ 0.059827f
C11057 _153_ _365_/a_692_472# 0.002377f
C11058 mask\[8\] net25 0.035648f
C11059 net51 net6 0.142515f
C11060 net20 _015_ 0.005917f
C11061 _070_ trim_mask\[0\] 0.006144f
C11062 _072_ _267_/a_36_472# 0.024239f
C11063 net17 FILLER_0_20_15/a_572_375# 0.018398f
C11064 _077_ FILLER_0_9_72/a_1380_472# 0.006408f
C11065 net80 output22/a_224_472# 0.00955f
C11066 _132_ FILLER_0_15_116/a_124_375# 0.047331f
C11067 _061_ vdd 0.295557f
C11068 net38 _278_/a_36_160# 0.010587f
C11069 net15 _183_ 0.007353f
C11070 FILLER_0_10_78/a_124_375# FILLER_0_9_72/a_932_472# 0.001543f
C11071 _175_ _043_ 0.001037f
C11072 net24 net71 0.015101f
C11073 _093_ FILLER_0_18_177/a_3172_472# 0.003708f
C11074 net75 _122_ 0.052177f
C11075 _429_/a_2248_156# FILLER_0_15_228/a_124_375# 0.030666f
C11076 net47 _156_ 0.040298f
C11077 FILLER_0_17_56/a_572_375# vdd 0.003489f
C11078 FILLER_0_17_56/a_124_375# vss 0.00143f
C11079 _002_ FILLER_0_3_172/a_3172_472# 0.002313f
C11080 net23 FILLER_0_22_128/a_1468_375# 0.001866f
C11081 _104_ net34 0.293336f
C11082 _079_ _263_/a_224_472# 0.002505f
C11083 output44/a_224_472# net44 0.051347f
C11084 net38 _444_/a_1000_472# 0.027886f
C11085 FILLER_0_8_37/a_484_472# _054_ 0.022621f
C11086 net34 _421_/a_2665_112# 0.001056f
C11087 _214_/a_36_160# FILLER_0_23_88/a_36_472# 0.006647f
C11088 ctlp[3] _108_ 0.009437f
C11089 output45/a_224_472# vss 0.00543f
C11090 output31/a_224_472# output36/a_224_472# 0.00289f
C11091 _269_/a_36_472# _078_ 0.033601f
C11092 FILLER_0_13_212/a_484_472# vss 0.002397f
C11093 net62 FILLER_0_13_212/a_1468_375# 0.003327f
C11094 _093_ _303_/a_36_472# 0.096502f
C11095 _142_ _431_/a_36_151# 0.030496f
C11096 _165_ net67 0.045827f
C11097 net58 FILLER_0_8_263/a_36_472# 0.059769f
C11098 _144_ _149_ 0.032178f
C11099 _012_ FILLER_0_23_44/a_1468_375# 0.002827f
C11100 _093_ _102_ 0.008937f
C11101 _436_/a_2248_156# vdd 0.011151f
C11102 _288_/a_224_472# vdd 0.002071f
C11103 mask\[5\] net32 0.304094f
C11104 net74 net36 0.012494f
C11105 _081_ _152_ 0.172002f
C11106 net34 result[6] 0.072393f
C11107 cal_count\[3\] _188_ 0.048745f
C11108 _040_ vss 0.216709f
C11109 vss _433_/a_1000_472# 0.002059f
C11110 net76 FILLER_0_5_206/a_124_375# 0.006974f
C11111 _176_ FILLER_0_11_78/a_36_472# 0.003603f
C11112 _125_ vss 0.149512f
C11113 _187_ net16 0.161791f
C11114 FILLER_0_22_86/a_1380_472# FILLER_0_22_107/a_36_472# 0.001963f
C11115 net60 _418_/a_2560_156# 0.020147f
C11116 FILLER_0_18_139/a_124_375# vdd 0.023256f
C11117 net66 _440_/a_796_472# 0.002718f
C11118 net49 _440_/a_36_151# 0.021133f
C11119 _256_/a_36_68# net4 0.017783f
C11120 _432_/a_2248_156# mask\[1\] 0.002293f
C11121 net50 FILLER_0_6_79/a_124_375# 0.004402f
C11122 _323_/a_36_113# _128_ 0.014377f
C11123 _104_ output33/a_224_472# 0.032929f
C11124 _369_/a_36_68# _154_ 0.042308f
C11125 FILLER_0_7_146/a_124_375# net37 0.005315f
C11126 net19 net18 0.028285f
C11127 net35 _423_/a_2665_112# 0.019085f
C11128 output33/a_224_472# _421_/a_2665_112# 0.010726f
C11129 net36 cal_count\[1\] 0.011481f
C11130 net68 _440_/a_36_151# 0.080854f
C11131 FILLER_0_5_54/a_124_375# FILLER_0_3_54/a_36_472# 0.001512f
C11132 _132_ FILLER_0_17_104/a_484_472# 0.002737f
C11133 _181_ vdd 0.209604f
C11134 FILLER_0_8_107/a_36_472# FILLER_0_9_105/a_124_375# 0.001684f
C11135 ctlp[1] _420_/a_796_472# 0.001468f
C11136 mask\[7\] FILLER_0_22_128/a_2364_375# 0.003632f
C11137 _095_ _225_/a_36_160# 0.001084f
C11138 FILLER_0_16_241/a_36_472# vss 0.004432f
C11139 FILLER_0_5_198/a_484_472# vss 0.001338f
C11140 output31/a_224_472# vdd 0.083516f
C11141 net34 net22 0.031404f
C11142 _062_ _227_/a_36_160# 0.015411f
C11143 net34 mask\[4\] 0.001774f
C11144 net35 FILLER_0_22_128/a_1828_472# 0.016187f
C11145 output33/a_224_472# result[6] 0.035032f
C11146 net50 FILLER_0_3_54/a_124_375# 0.00189f
C11147 _130_ vdd 0.046379f
C11148 trim_val\[2\] _381_/a_36_472# 0.005253f
C11149 _174_ _401_/a_244_472# 0.001957f
C11150 FILLER_0_7_72/a_2724_472# net50 0.007192f
C11151 _114_ _128_ 0.047516f
C11152 _343_/a_257_69# _137_ 0.003494f
C11153 net72 FILLER_0_17_56/a_572_375# 0.004473f
C11154 _003_ cal_itt\[3\] 0.054183f
C11155 net73 FILLER_0_18_107/a_124_375# 0.003742f
C11156 trim_val\[4\] FILLER_0_2_165/a_36_472# 0.007765f
C11157 vss FILLER_0_12_196/a_36_472# 0.003551f
C11158 output15/a_224_472# net15 0.028578f
C11159 net64 FILLER_0_9_282/a_36_472# 0.031302f
C11160 FILLER_0_15_142/a_124_375# net23 0.002212f
C11161 _136_ FILLER_0_16_154/a_1380_472# 0.006517f
C11162 trim_mask\[1\] FILLER_0_6_47/a_484_472# 0.022211f
C11163 _174_ vss 0.188373f
C11164 net39 _445_/a_36_151# 0.006056f
C11165 FILLER_0_1_266/a_36_472# net8 0.0138f
C11166 cal_itt\[3\] net21 0.175781f
C11167 _003_ _081_ 0.041822f
C11168 net16 _445_/a_2248_156# 0.003321f
C11169 _093_ _198_/a_67_603# 0.004447f
C11170 _086_ FILLER_0_7_104/a_1380_472# 0.034829f
C11171 FILLER_0_4_197/a_932_472# net22 0.0473f
C11172 FILLER_0_11_101/a_124_375# _070_ 0.052406f
C11173 _052_ FILLER_0_18_37/a_1020_375# 0.001287f
C11174 FILLER_0_1_98/a_36_472# _153_ 0.001463f
C11175 _444_/a_2248_156# vss 0.001329f
C11176 _444_/a_2665_112# vdd 0.029351f
C11177 _086_ _318_/a_224_472# 0.007024f
C11178 FILLER_0_12_220/a_36_472# _090_ 0.023446f
C11179 _081_ net21 0.030964f
C11180 net10 output11/a_224_472# 0.095679f
C11181 _155_ FILLER_0_7_104/a_36_472# 0.005042f
C11182 trim_mask\[2\] _153_ 0.007934f
C11183 fanout77/a_36_113# _418_/a_36_151# 0.001082f
C11184 _446_/a_1308_423# vdd 0.002346f
C11185 _421_/a_448_472# _419_/a_2665_112# 0.002393f
C11186 ctlp[1] _421_/a_1204_472# 0.003759f
C11187 _427_/a_2665_112# net23 0.032729f
C11188 _065_ net66 0.003956f
C11189 state\[2\] FILLER_0_13_142/a_124_375# 0.010494f
C11190 net53 FILLER_0_13_142/a_1020_375# 0.001597f
C11191 _119_ FILLER_0_7_104/a_1380_472# 0.002603f
C11192 FILLER_0_5_72/a_572_375# vdd -0.00211f
C11193 FILLER_0_5_72/a_124_375# vss 0.041166f
C11194 FILLER_0_17_226/a_124_375# _106_ 0.061857f
C11195 output14/a_224_472# _442_/a_448_472# 0.008149f
C11196 _446_/a_1204_472# net17 0.003628f
C11197 output11/a_224_472# FILLER_0_0_232/a_124_375# 0.00515f
C11198 _316_/a_848_380# _123_ 0.0018f
C11199 FILLER_0_7_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001723f
C11200 _076_ FILLER_0_8_239/a_124_375# 0.007237f
C11201 net32 net30 0.004658f
C11202 _143_ FILLER_0_18_139/a_1468_375# 0.001097f
C11203 FILLER_0_4_91/a_36_472# _160_ 0.007864f
C11204 net72 _181_ 0.004503f
C11205 _070_ _081_ 0.00804f
C11206 net4 calibrate 0.04302f
C11207 mask\[8\] FILLER_0_22_107/a_484_472# 0.024416f
C11208 net35 FILLER_0_22_107/a_36_472# 0.007196f
C11209 FILLER_0_7_162/a_124_375# vss 0.018732f
C11210 FILLER_0_5_109/a_124_375# _163_ 0.002658f
C11211 _414_/a_2248_156# _122_ 0.002838f
C11212 _104_ mask\[2\] 0.002737f
C11213 _404_/a_36_472# _179_ 0.00141f
C11214 FILLER_0_21_142/a_572_375# _433_/a_2665_112# 0.001092f
C11215 _417_/a_1204_472# net30 0.001496f
C11216 FILLER_0_16_89/a_484_472# _136_ 0.032722f
C11217 _417_/a_796_472# result[3] 0.001206f
C11218 net27 result[0] 0.106157f
C11219 FILLER_0_9_223/a_36_472# _090_ 0.001057f
C11220 output9/a_224_472# input4/a_36_68# 0.009732f
C11221 trim_val\[3\] FILLER_0_2_93/a_124_375# 0.001032f
C11222 _258_/a_36_160# _073_ 0.079254f
C11223 _408_/a_728_93# net17 0.005494f
C11224 _270_/a_36_472# net21 0.001606f
C11225 _131_ _134_ 0.887647f
C11226 FILLER_0_12_136/a_1468_375# _126_ 0.012732f
C11227 _089_ _003_ 0.014763f
C11228 FILLER_0_16_107/a_484_472# FILLER_0_16_115/a_36_472# 0.013276f
C11229 _436_/a_2248_156# FILLER_0_22_128/a_572_375# 0.006739f
C11230 _436_/a_2665_112# FILLER_0_22_128/a_124_375# 0.004834f
C11231 _092_ _293_/a_36_472# 0.004828f
C11232 _056_ _055_ 0.155993f
C11233 net15 _449_/a_448_472# 0.040076f
C11234 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_572_375# 0.086635f
C11235 _094_ _418_/a_2248_156# 0.028557f
C11236 fanout56/a_36_113# _098_ 0.019463f
C11237 _089_ net21 0.006605f
C11238 _091_ vdd 1.011371f
C11239 _058_ net23 0.075446f
C11240 result[7] _420_/a_36_151# 0.006868f
C11241 fanout78/a_36_113# net18 0.001419f
C11242 _307_/a_672_472# _126_ 0.00121f
C11243 FILLER_0_4_197/a_484_472# net21 0.046864f
C11244 _185_ _402_/a_1296_93# 0.001714f
C11245 vss _166_ 0.011302f
C11246 vdd _160_ 0.606139f
C11247 _315_/a_36_68# net23 0.030384f
C11248 _086_ _070_ 0.123033f
C11249 net62 _416_/a_2560_156# 0.010748f
C11250 _420_/a_36_151# FILLER_0_23_282/a_484_472# 0.001723f
C11251 _414_/a_36_151# _053_ 0.035994f
C11252 output34/a_224_472# _199_/a_36_160# 0.003531f
C11253 _430_/a_36_151# _136_ 0.02044f
C11254 _141_ FILLER_0_19_155/a_572_375# 0.033271f
C11255 FILLER_0_16_89/a_1468_375# FILLER_0_17_72/a_3260_375# 0.026339f
C11256 FILLER_0_16_89/a_484_472# FILLER_0_17_72/a_2364_375# 0.001723f
C11257 _410_/a_36_68# _042_ 0.041079f
C11258 _408_/a_2215_68# _186_ 0.001205f
C11259 _026_ FILLER_0_20_87/a_124_375# 0.031902f
C11260 _430_/a_36_151# net21 0.019114f
C11261 _072_ _118_ 0.120452f
C11262 FILLER_0_10_78/a_572_375# _120_ 0.006134f
C11263 net50 FILLER_0_4_91/a_484_472# 0.008749f
C11264 FILLER_0_24_96/a_124_375# vdd 0.029269f
C11265 output28/a_224_472# net79 0.04262f
C11266 valid _425_/a_2248_156# 0.00154f
C11267 _140_ FILLER_0_22_128/a_3172_472# 0.005458f
C11268 _119_ _070_ 1.949038f
C11269 _449_/a_36_151# _038_ 0.019666f
C11270 _432_/a_2248_156# FILLER_0_18_177/a_1828_472# 0.035805f
C11271 mask\[2\] net22 0.034216f
C11272 net15 FILLER_0_15_59/a_484_472# 0.015199f
C11273 FILLER_0_16_57/a_572_375# _176_ 0.006422f
C11274 _267_/a_36_472# state\[1\] 0.001647f
C11275 ctlp[7] _211_/a_36_160# 0.003488f
C11276 FILLER_0_9_270/a_36_472# vdd 0.008742f
C11277 FILLER_0_9_270/a_572_375# vss 0.017196f
C11278 _015_ vss 0.090048f
C11279 ctlp[4] net32 0.001413f
C11280 FILLER_0_17_72/a_1916_375# _136_ 0.009573f
C11281 net20 FILLER_0_15_235/a_36_472# 0.002227f
C11282 _144_ FILLER_0_19_155/a_484_472# 0.006137f
C11283 _374_/a_36_68# _061_ 0.026111f
C11284 net36 _097_ 0.022089f
C11285 FILLER_0_22_128/a_2724_472# _146_ 0.002471f
C11286 _025_ _436_/a_796_472# 0.026852f
C11287 FILLER_0_21_125/a_484_472# _022_ 0.004649f
C11288 result[7] _421_/a_1308_423# 0.022204f
C11289 net79 net77 0.431572f
C11290 _428_/a_2248_156# vdd 0.006977f
C11291 _031_ FILLER_0_2_127/a_36_472# 0.016207f
C11292 _120_ FILLER_0_8_156/a_572_375# 0.030218f
C11293 FILLER_0_5_54/a_572_375# vss 0.002617f
C11294 FILLER_0_5_54/a_1020_375# vdd -0.014642f
C11295 FILLER_0_4_99/a_124_375# net14 0.003714f
C11296 net63 net33 0.048496f
C11297 FILLER_0_16_73/a_36_472# FILLER_0_17_72/a_124_375# 0.001723f
C11298 FILLER_0_16_89/a_932_472# net53 0.012534f
C11299 FILLER_0_12_220/a_932_472# _070_ 0.001282f
C11300 result[8] FILLER_0_24_274/a_36_472# 0.005458f
C11301 output43/a_224_472# vss -0.005182f
C11302 _413_/a_1308_423# _002_ 0.002178f
C11303 _326_/a_36_160# _086_ 0.063565f
C11304 FILLER_0_15_72/a_484_472# vss 0.010761f
C11305 FILLER_0_7_72/a_1020_375# vdd 0.004039f
C11306 FILLER_0_12_124/a_36_472# _127_ 0.01468f
C11307 FILLER_0_7_195/a_124_375# _163_ 0.001308f
C11308 net50 vss 1.178736f
C11309 FILLER_0_17_72/a_3172_472# _131_ 0.003717f
C11310 _074_ _375_/a_1388_497# 0.005488f
C11311 _077_ _176_ 0.00497f
C11312 FILLER_0_5_128/a_36_472# net74 0.01163f
C11313 _281_/a_234_472# _098_ 0.003724f
C11314 _414_/a_448_472# _074_ 0.008725f
C11315 _181_ cal_count\[0\] 0.001114f
C11316 _443_/a_1204_472# vss 0.005425f
C11317 _443_/a_2248_156# vdd 0.010579f
C11318 _128_ _085_ 0.004532f
C11319 _276_/a_36_160# mask\[4\] 0.025336f
C11320 _412_/a_1308_423# net1 0.022273f
C11321 FILLER_0_19_28/a_572_375# net40 0.00139f
C11322 mask\[3\] FILLER_0_17_161/a_36_472# 0.13873f
C11323 vdd FILLER_0_3_212/a_124_375# 0.025095f
C11324 net53 _136_ 0.099584f
C11325 _326_/a_36_160# _119_ 0.003944f
C11326 FILLER_0_4_197/a_36_472# _088_ 0.067725f
C11327 output28/a_224_472# _416_/a_2665_112# 0.008243f
C11328 result[1] _416_/a_1308_423# 0.002597f
C11329 net18 _193_/a_36_160# 0.114176f
C11330 net80 _137_ 0.260786f
C11331 FILLER_0_18_171/a_124_375# net80 0.024341f
C11332 net58 FILLER_0_8_247/a_1468_375# 0.001669f
C11333 _430_/a_1308_423# _429_/a_36_151# 0.001722f
C11334 _072_ _068_ 0.185471f
C11335 _410_/a_36_68# cal_count\[3\] 0.001096f
C11336 FILLER_0_5_72/a_1468_375# _440_/a_2248_156# 0.030666f
C11337 FILLER_0_5_72/a_1020_375# _440_/a_2665_112# 0.010688f
C11338 output21/a_224_472# net33 0.001166f
C11339 _431_/a_2665_112# _136_ 0.035394f
C11340 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_36_472# 0.086635f
C11341 FILLER_0_9_223/a_36_472# _076_ 0.00146f
C11342 _056_ _058_ 0.988919f
C11343 net8 vdd 0.593788f
C11344 _164_ FILLER_0_6_47/a_484_472# 0.012286f
C11345 net19 _420_/a_1000_472# 0.006558f
C11346 net81 output48/a_224_472# 0.040059f
C11347 net80 FILLER_0_19_171/a_36_472# 0.040915f
C11348 FILLER_0_7_72/a_124_375# net50 0.009304f
C11349 net44 FILLER_0_8_2/a_124_375# 0.083677f
C11350 net19 _109_ 0.005991f
C11351 net67 FILLER_0_6_47/a_36_472# 0.004607f
C11352 net58 _426_/a_36_151# 0.002612f
C11353 _052_ FILLER_0_17_38/a_484_472# 0.001368f
C11354 _132_ FILLER_0_18_107/a_1828_472# 0.045833f
C11355 net16 FILLER_0_18_37/a_484_472# 0.054878f
C11356 _144_ FILLER_0_22_128/a_3260_375# 0.006444f
C11357 _069_ vss 0.323941f
C11358 net46 net40 0.254778f
C11359 _308_/a_1084_68# _114_ 0.00178f
C11360 mask\[0\] _138_ 0.22533f
C11361 net81 net5 0.006276f
C11362 _432_/a_796_472# _091_ 0.018082f
C11363 _068_ net47 0.001491f
C11364 _150_ vdd 0.05295f
C11365 _363_/a_36_68# _154_ 0.149319f
C11366 net36 FILLER_0_15_180/a_124_375# 0.004275f
C11367 FILLER_0_7_146/a_36_472# calibrate 0.060587f
C11368 net29 vss 0.259409f
C11369 ctlp[1] _419_/a_1000_472# 0.005263f
C11370 _121_ FILLER_0_8_156/a_124_375# 0.033427f
C11371 _170_ vdd 0.18848f
C11372 net52 net55 0.016401f
C11373 _104_ net20 0.482229f
C11374 _005_ _192_/a_67_603# 0.013886f
C11375 _448_/a_36_151# net12 0.133216f
C11376 _448_/a_1308_423# net22 0.045644f
C11377 _434_/a_796_472# mask\[6\] 0.004416f
C11378 trimb[1] FILLER_0_18_2/a_124_375# 0.01352f
C11379 _432_/a_2560_156# _139_ 0.002737f
C11380 _421_/a_2248_156# net19 0.016721f
C11381 result[7] FILLER_0_24_274/a_932_472# 0.006454f
C11382 FILLER_0_15_212/a_36_472# vss 0.002853f
C11383 _093_ FILLER_0_18_76/a_484_472# 0.024853f
C11384 FILLER_0_15_116/a_124_375# vdd 0.012886f
C11385 FILLER_0_6_90/a_36_472# net14 0.002705f
C11386 fanout81/a_36_160# net9 0.002274f
C11387 _422_/a_448_472# net19 0.003382f
C11388 net69 _168_ 0.035976f
C11389 _428_/a_36_151# net14 0.004485f
C11390 net75 net8 0.553872f
C11391 net20 result[6] 0.026511f
C11392 FILLER_0_5_164/a_572_375# net37 0.014025f
C11393 FILLER_0_19_47/a_124_375# net26 0.008432f
C11394 ctln[1] ctln[2] 0.047127f
C11395 _050_ FILLER_0_22_128/a_932_472# 0.001098f
C11396 _114_ net14 0.127764f
C11397 _134_ FILLER_0_10_107/a_124_375# 0.009573f
C11398 net55 _216_/a_67_603# 0.071821f
C11399 _429_/a_2665_112# FILLER_0_14_235/a_124_375# 0.006271f
C11400 FILLER_0_17_38/a_124_375# _452_/a_36_151# 0.006111f
C11401 _407_/a_36_472# _181_ 0.035594f
C11402 state\[1\] _113_ 0.107642f
C11403 FILLER_0_18_2/a_3260_375# net40 0.035372f
C11404 _397_/a_244_68# net55 0.001173f
C11405 output8/a_224_472# net65 0.084944f
C11406 net16 FILLER_0_8_37/a_484_472# 0.004272f
C11407 net34 FILLER_0_22_177/a_1380_472# 0.003953f
C11408 _420_/a_1000_472# _009_ 0.019219f
C11409 output35/a_224_472# output19/a_224_472# 0.015892f
C11410 net41 cal_count\[3\] 0.028902f
C11411 trim[2] trim[3] 0.056575f
C11412 net52 net23 0.093434f
C11413 output48/a_224_472# _079_ 0.003556f
C11414 _293_/a_36_472# vdd 0.087136f
C11415 _019_ net36 0.309649f
C11416 _009_ _109_ 0.006736f
C11417 mask\[4\] FILLER_0_18_177/a_2364_375# 0.01602f
C11418 FILLER_0_4_197/a_124_375# _079_ 0.004772f
C11419 mask\[5\] _105_ 0.706158f
C11420 mask\[4\] _339_/a_36_160# 0.003234f
C11421 _443_/a_796_472# net23 0.002306f
C11422 _443_/a_448_472# net13 0.002263f
C11423 FILLER_0_20_177/a_572_375# vdd -0.001627f
C11424 FILLER_0_20_177/a_124_375# vss 0.002674f
C11425 _088_ FILLER_0_3_221/a_124_375# 0.002378f
C11426 _250_/a_36_68# state\[2\] 0.038165f
C11427 output28/a_224_472# output29/a_224_472# 0.00289f
C11428 net34 _297_/a_36_472# 0.005603f
C11429 _067_ net6 0.015232f
C11430 net50 _441_/a_1204_472# 0.006986f
C11431 net52 _441_/a_2665_112# 0.004975f
C11432 net50 trim_mask\[2\] 0.267074f
C11433 _440_/a_36_151# net47 0.013626f
C11434 _188_ _120_ 0.046757f
C11435 FILLER_0_13_212/a_484_472# net79 0.00402f
C11436 FILLER_0_4_49/a_484_472# net66 0.015555f
C11437 FILLER_0_4_49/a_124_375# net49 0.005427f
C11438 net55 _406_/a_36_159# 0.001219f
C11439 FILLER_0_12_136/a_1468_375# FILLER_0_13_142/a_932_472# 0.001684f
C11440 fanout50/a_36_160# _447_/a_2665_112# 0.002885f
C11441 _432_/a_1000_472# vdd 0.010431f
C11442 FILLER_0_16_89/a_484_472# _451_/a_448_472# 0.059367f
C11443 _096_ _320_/a_1792_472# 0.001419f
C11444 net52 fanout74/a_36_113# 0.001514f
C11445 FILLER_0_4_49/a_124_375# net68 0.008422f
C11446 FILLER_0_16_255/a_36_472# net30 0.00209f
C11447 _102_ _094_ 0.727442f
C11448 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_36_472# 0.086635f
C11449 net74 _372_/a_786_69# 0.00149f
C11450 net82 _443_/a_36_151# 0.03565f
C11451 _003_ _161_ 0.004981f
C11452 net50 _439_/a_1000_472# 0.005154f
C11453 net52 _439_/a_2248_156# 0.00258f
C11454 _070_ FILLER_0_11_109/a_36_472# 0.001091f
C11455 FILLER_0_17_104/a_36_472# vss 0.002744f
C11456 FILLER_0_17_104/a_484_472# vdd 0.020339f
C11457 net81 net80 0.006516f
C11458 _095_ FILLER_0_14_107/a_124_375# 0.01418f
C11459 output8/a_224_472# net59 0.00398f
C11460 _015_ net4 0.003985f
C11461 _012_ vdd 0.261844f
C11462 net65 FILLER_0_9_282/a_572_375# 0.001388f
C11463 _050_ FILLER_0_22_107/a_124_375# 0.002634f
C11464 _425_/a_1204_472# net37 0.001403f
C11465 _144_ _098_ 1.252524f
C11466 _013_ _183_ 0.00176f
C11467 FILLER_0_4_144/a_124_375# _059_ 0.031451f
C11468 _161_ net21 0.011799f
C11469 result[7] _419_/a_448_472# 0.021809f
C11470 _032_ trim_mask\[4\] 0.010578f
C11471 vdd _156_ 0.178622f
C11472 _010_ _420_/a_2248_156# 0.047408f
C11473 _131_ _331_/a_244_472# 0.002331f
C11474 net41 net40 2.687418f
C11475 _136_ _451_/a_36_151# 0.043941f
C11476 net41 FILLER_0_21_28/a_932_472# 0.014034f
C11477 net34 _140_ 0.033459f
C11478 _000_ _079_ 0.032884f
C11479 _365_/a_244_472# _156_ 0.003847f
C11480 _053_ _439_/a_2665_112# 0.006037f
C11481 _267_/a_36_472# vdd 0.005477f
C11482 fanout79/a_36_160# _094_ 0.008308f
C11483 FILLER_0_21_286/a_36_472# net77 0.001557f
C11484 _422_/a_448_472# _009_ 0.018984f
C11485 ctlp[1] FILLER_0_23_282/a_572_375# 0.009848f
C11486 mask\[8\] _437_/a_448_472# 0.008198f
C11487 ctln[1] FILLER_0_3_221/a_1468_375# 0.001235f
C11488 _030_ FILLER_0_3_78/a_36_472# 0.007376f
C11489 net49 FILLER_0_3_78/a_572_375# 0.066078f
C11490 _012_ FILLER_0_23_60/a_36_472# 0.001572f
C11491 _031_ FILLER_0_2_111/a_484_472# 0.027347f
C11492 net69 FILLER_0_2_111/a_1380_472# 0.021896f
C11493 net63 _430_/a_1308_423# 0.01125f
C11494 trimb[1] net17 0.084269f
C11495 en clk 0.067072f
C11496 FILLER_0_3_204/a_124_375# net22 0.031438f
C11497 _379_/a_36_472# trim_mask\[1\] 0.003592f
C11498 net44 _452_/a_2449_156# 0.0059f
C11499 _178_ _402_/a_1948_68# 0.00815f
C11500 _126_ FILLER_0_13_206/a_124_375# 0.002746f
C11501 net36 FILLER_0_18_76/a_124_375# 0.001741f
C11502 ctln[0] output7/a_224_472# 0.081823f
C11503 ctln[4] output11/a_224_472# 0.072677f
C11504 net23 _387_/a_36_113# 0.031688f
C11505 _077_ FILLER_0_8_239/a_36_472# 0.001289f
C11506 FILLER_0_19_171/a_1468_375# vdd 0.064097f
C11507 en_co_clk _171_ 0.003472f
C11508 _091_ FILLER_0_13_212/a_572_375# 0.022882f
C11509 _161_ _070_ 0.027757f
C11510 FILLER_0_16_73/a_572_375# net15 0.002076f
C11511 net82 FILLER_0_2_177/a_124_375# 0.003837f
C11512 _140_ _354_/a_49_472# 0.004731f
C11513 _114_ _311_/a_2700_473# 0.005178f
C11514 _016_ _043_ 0.030341f
C11515 FILLER_0_15_235/a_484_472# vdd 0.006f
C11516 FILLER_0_15_235/a_36_472# vss 0.003138f
C11517 net62 FILLER_0_15_235/a_124_375# 0.001315f
C11518 _053_ calibrate 0.081635f
C11519 net78 _421_/a_448_472# 0.025808f
C11520 FILLER_0_17_282/a_36_472# _418_/a_448_472# 0.011962f
C11521 FILLER_0_18_177/a_3260_375# net21 0.005704f
C11522 _144_ _433_/a_2248_156# 0.021805f
C11523 _438_/a_448_472# vdd 0.009409f
C11524 _438_/a_36_151# vss 0.014203f
C11525 FILLER_0_18_2/a_2812_375# FILLER_0_19_28/a_36_472# 0.001684f
C11526 FILLER_0_4_177/a_124_375# _386_/a_848_380# 0.001277f
C11527 FILLER_0_21_286/a_484_472# FILLER_0_23_290/a_124_375# 0.001404f
C11528 result[2] FILLER_0_13_290/a_36_472# 0.016496f
C11529 _079_ FILLER_0_5_212/a_36_472# 0.005671f
C11530 fanout60/a_36_160# net18 0.004124f
C11531 net20 ctln[1] 0.135151f
C11532 _091_ _337_/a_49_472# 0.014992f
C11533 net55 FILLER_0_18_61/a_124_375# 0.040701f
C11534 cal_count\[1\] FILLER_0_15_59/a_124_375# 0.010034f
C11535 FILLER_0_14_91/a_36_472# _095_ 0.014431f
C11536 _189_/a_67_603# FILLER_0_14_235/a_36_472# 0.002778f
C11537 FILLER_0_0_130/a_36_472# vss 0.00351f
C11538 FILLER_0_14_81/a_36_472# _177_ 0.004294f
C11539 FILLER_0_15_142/a_36_472# vdd 0.106034f
C11540 _063_ _445_/a_2248_156# 0.008121f
C11541 _054_ vss 0.176655f
C11542 net20 _076_ 0.228128f
C11543 net72 _012_ 0.002382f
C11544 FILLER_0_15_212/a_1380_472# FILLER_0_15_228/a_36_472# 0.013277f
C11545 _053_ _153_ 0.015583f
C11546 _008_ _419_/a_448_472# 0.01758f
C11547 en_co_clk _176_ 0.099475f
C11548 _017_ FILLER_0_14_107/a_932_472# 0.001941f
C11549 _069_ net4 0.07542f
C11550 _067_ FILLER_0_12_20/a_572_375# 0.01186f
C11551 _147_ _208_/a_36_160# 0.006056f
C11552 fanout69/a_36_113# _032_ 0.003681f
C11553 _247_/a_36_160# _060_ 0.055366f
C11554 _412_/a_1204_472# net76 0.020975f
C11555 _274_/a_36_68# _091_ 0.025773f
C11556 net52 trim_val\[4\] 0.21532f
C11557 mask\[4\] FILLER_0_19_187/a_124_375# 0.006236f
C11558 _420_/a_2248_156# vdd 0.00331f
C11559 FILLER_0_15_142/a_484_472# vdd 0.001097f
C11560 _094_ _283_/a_36_472# 0.004373f
C11561 net15 _111_ 0.049514f
C11562 net53 _451_/a_448_472# 0.026909f
C11563 net70 _451_/a_836_156# 0.006451f
C11564 _115_ FILLER_0_9_105/a_36_472# 0.004013f
C11565 _411_/a_36_151# _000_ 0.023297f
C11566 output48/a_224_472# net64 0.002845f
C11567 _430_/a_2248_156# mask\[3\] 0.004211f
C11568 _008_ mask\[2\] 0.003475f
C11569 ctln[1] FILLER_0_1_266/a_484_472# 0.002068f
C11570 _414_/a_36_151# cal_itt\[3\] 0.049033f
C11571 _013_ FILLER_0_18_37/a_932_472# 0.010651f
C11572 FILLER_0_8_138/a_36_472# _129_ 0.055537f
C11573 mask\[9\] _438_/a_2665_112# 0.040085f
C11574 _183_ _179_ 0.017086f
C11575 net64 net5 0.098088f
C11576 _376_/a_36_160# FILLER_0_6_79/a_36_472# 0.003913f
C11577 FILLER_0_3_172/a_36_472# net22 0.012287f
C11578 _434_/a_1204_472# vdd 0.005382f
C11579 _427_/a_448_472# _043_ 0.002896f
C11580 _414_/a_36_151# _081_ 0.016708f
C11581 FILLER_0_4_177/a_36_472# vdd 0.114788f
C11582 FILLER_0_4_177/a_572_375# vss 0.054783f
C11583 FILLER_0_13_142/a_36_472# vss 0.005768f
C11584 net57 FILLER_0_8_156/a_484_472# 0.008895f
C11585 fanout66/a_36_113# _440_/a_36_151# 0.017895f
C11586 _417_/a_448_472# vss 0.005289f
C11587 _417_/a_1308_423# vdd 0.002263f
C11588 _285_/a_36_472# _045_ 0.00269f
C11589 FILLER_0_4_99/a_36_472# _160_ 0.006222f
C11590 _149_ _354_/a_49_472# 0.017453f
C11591 _424_/a_36_151# _012_ 0.005964f
C11592 FILLER_0_16_57/a_572_375# FILLER_0_15_59/a_484_472# 0.001543f
C11593 FILLER_0_8_127/a_124_375# _070_ 0.003265f
C11594 cal_count\[3\] _390_/a_36_68# 0.003074f
C11595 FILLER_0_12_124/a_124_375# vss 0.012672f
C11596 _411_/a_1000_472# net8 0.007241f
C11597 sample output27/a_224_472# 0.006116f
C11598 _127_ _070_ 0.031272f
C11599 _104_ vss 0.564464f
C11600 _112_ net37 0.070289f
C11601 FILLER_0_17_226/a_124_375# FILLER_0_17_218/a_572_375# 0.012001f
C11602 _177_ _451_/a_3129_107# 0.043731f
C11603 _044_ FILLER_0_14_263/a_124_375# 0.001047f
C11604 _421_/a_2665_112# vss 0.002792f
C11605 _421_/a_2560_156# vdd 0.001862f
C11606 FILLER_0_22_86/a_124_375# net71 0.002239f
C11607 _104_ _298_/a_224_472# 0.001731f
C11608 ctln[6] FILLER_0_0_130/a_124_375# 0.026786f
C11609 net58 ctln[2] 0.025352f
C11610 ctlp[4] _105_ 0.002221f
C11611 cal_count\[3\] _408_/a_718_524# 0.005968f
C11612 comp net3 0.05248f
C11613 _442_/a_2665_112# net14 0.011563f
C11614 _164_ net40 0.048933f
C11615 _414_/a_2665_112# _077_ 0.001675f
C11616 output27/a_224_472# vss 0.027374f
C11617 _422_/a_796_472# vdd 0.003546f
C11618 trim_val\[4\] _387_/a_36_113# 0.005339f
C11619 net76 _037_ 0.010891f
C11620 FILLER_0_8_107/a_124_375# _070_ 0.003069f
C11621 _426_/a_2248_156# vdd 0.003943f
C11622 FILLER_0_12_136/a_484_472# _076_ 0.001683f
C11623 output34/a_224_472# _046_ 0.006059f
C11624 _087_ FILLER_0_5_181/a_124_375# 0.068f
C11625 cal_count\[3\] cal_count\[2\] 0.005307f
C11626 _414_/a_1456_156# cal_itt\[3\] 0.001134f
C11627 _359_/a_1044_488# _129_ 0.001111f
C11628 _088_ FILLER_0_3_172/a_2364_375# 0.002377f
C11629 result[6] vss 0.310169f
C11630 FILLER_0_15_282/a_36_472# vss 0.004616f
C11631 net62 FILLER_0_15_282/a_124_375# 0.012711f
C11632 _446_/a_2560_156# net40 0.012204f
C11633 _081_ _084_ 0.016804f
C11634 FILLER_0_11_101/a_484_472# vss 0.003923f
C11635 _075_ _056_ 0.001957f
C11636 _086_ _414_/a_36_151# 0.002687f
C11637 _090_ vss 0.267577f
C11638 _113_ vdd 0.774039f
C11639 net69 _441_/a_796_472# 0.002057f
C11640 fanout61/a_36_113# vss 0.05514f
C11641 _093_ FILLER_0_16_89/a_124_375# 0.004086f
C11642 trim_val\[3\] _441_/a_2248_156# 0.027464f
C11643 FILLER_0_4_49/a_36_472# _164_ 0.033727f
C11644 _414_/a_36_151# _089_ 0.039611f
C11645 net71 _437_/a_1000_472# 0.014459f
C11646 _447_/a_36_151# net69 0.001216f
C11647 FILLER_0_9_223/a_36_472# _128_ 0.00702f
C11648 _064_ _445_/a_2560_156# 0.005361f
C11649 cal_count\[3\] FILLER_0_11_124/a_36_472# 0.00702f
C11650 ctlp[7] FILLER_0_24_130/a_124_375# 0.002726f
C11651 cal_itt\[2\] _073_ 0.202415f
C11652 _070_ _071_ 0.001757f
C11653 _122_ FILLER_0_5_164/a_572_375# 0.001352f
C11654 net74 _059_ 0.004133f
C11655 net46 FILLER_0_20_15/a_1020_375# 0.0302f
C11656 _127_ FILLER_0_9_142/a_36_472# 0.004721f
C11657 output25/a_224_472# vss 0.080847f
C11658 _431_/a_36_151# vss 0.00849f
C11659 _411_/a_2665_112# net19 0.00934f
C11660 _408_/a_718_524# net40 0.011463f
C11661 _415_/a_448_472# net18 0.057688f
C11662 mask\[4\] vss 0.426009f
C11663 FILLER_0_5_172/a_36_472# net47 0.0015f
C11664 net22 vss 1.28233f
C11665 _330_/a_224_472# _134_ 0.007508f
C11666 fanout49/a_36_160# FILLER_0_4_91/a_36_472# 0.001461f
C11667 _300_/a_224_472# _009_ 0.001405f
C11668 cal_count\[2\] net40 0.313209f
C11669 _439_/a_2665_112# trim_mask\[0\] 0.020363f
C11670 _410_/a_36_68# _120_ 0.073688f
C11671 _379_/a_36_472# _164_ 0.026812f
C11672 _028_ _153_ 0.008011f
C11673 _431_/a_796_472# _136_ 0.009889f
C11674 FILLER_0_2_111/a_124_375# vdd 0.024756f
C11675 net66 _167_ 0.016569f
C11676 result[7] net20 0.134149f
C11677 FILLER_0_4_152/a_36_472# _170_ 0.005476f
C11678 FILLER_0_24_96/a_124_375# net24 0.040364f
C11679 FILLER_0_3_78/a_484_472# _164_ 0.05311f
C11680 FILLER_0_20_193/a_484_472# FILLER_0_19_195/a_124_375# 0.001543f
C11681 net73 FILLER_0_18_107/a_3172_472# 0.00533f
C11682 _428_/a_36_151# _131_ 0.00821f
C11683 _081_ FILLER_0_5_148/a_36_472# 0.020403f
C11684 _118_ vdd 0.292155f
C11685 _043_ FILLER_0_13_72/a_484_472# 0.016114f
C11686 _093_ FILLER_0_18_209/a_36_472# 0.007068f
C11687 FILLER_0_4_107/a_36_472# trim_mask\[3\] 0.00152f
C11688 _412_/a_1000_472# net76 0.024114f
C11689 FILLER_0_18_107/a_1828_472# vdd 0.004446f
C11690 ctln[8] vdd 0.125219f
C11691 net26 FILLER_0_21_28/a_1380_472# 0.035291f
C11692 fanout78/a_36_113# _418_/a_36_151# 0.030244f
C11693 FILLER_0_2_171/a_124_375# net22 0.009924f
C11694 trim_val\[1\] FILLER_0_6_47/a_36_472# 0.00351f
C11695 FILLER_0_5_109/a_572_375# _160_ 0.004207f
C11696 net78 _419_/a_36_151# 0.007437f
C11697 _016_ FILLER_0_12_136/a_124_375# 0.008914f
C11698 FILLER_0_14_107/a_484_472# _451_/a_36_151# 0.001723f
C11699 net80 mask\[1\] 0.015535f
C11700 _026_ _437_/a_448_472# 0.026072f
C11701 net10 FILLER_0_0_232/a_36_472# 0.016287f
C11702 net54 FILLER_0_22_128/a_1380_472# 0.008765f
C11703 FILLER_0_18_139/a_1380_472# _145_ 0.002077f
C11704 _114_ _131_ 0.036548f
C11705 _053_ FILLER_0_7_162/a_124_375# 0.007494f
C11706 net34 _435_/a_36_151# 0.011954f
C11707 _087_ vdd 0.281159f
C11708 FILLER_0_9_223/a_124_375# state\[0\] 0.002912f
C11709 FILLER_0_13_65/a_36_472# FILLER_0_13_72/a_36_472# 0.002765f
C11710 FILLER_0_10_214/a_36_472# _070_ 0.014734f
C11711 net41 _445_/a_448_472# 0.002211f
C11712 _069_ net79 0.045808f
C11713 net41 trim[3] 0.005906f
C11714 _035_ vss 0.105648f
C11715 FILLER_0_13_142/a_1020_375# net23 0.047331f
C11716 _425_/a_2248_156# calibrate 0.022237f
C11717 fanout49/a_36_160# vdd 0.099887f
C11718 net47 output6/a_224_472# 0.070584f
C11719 output14/a_224_472# _031_ 0.001077f
C11720 _413_/a_796_472# _002_ 0.009261f
C11721 _018_ FILLER_0_15_205/a_124_375# 0.002309f
C11722 trim_val\[4\] FILLER_0_5_164/a_484_472# 0.00172f
C11723 _155_ vss 0.13648f
C11724 FILLER_0_16_57/a_1380_472# _175_ 0.002834f
C11725 net27 _283_/a_36_472# 0.023243f
C11726 _038_ vss 0.373776f
C11727 result[5] _419_/a_36_151# 0.006539f
C11728 output34/a_224_472# net18 0.126175f
C11729 FILLER_0_2_165/a_124_375# net22 0.206491f
C11730 net11 vss 0.057193f
C11731 _077_ FILLER_0_9_60/a_36_472# 0.038809f
C11732 FILLER_0_16_255/a_36_472# _417_/a_2665_112# 0.003221f
C11733 _413_/a_36_151# FILLER_0_3_172/a_2276_472# 0.001723f
C11734 _236_/a_36_160# _444_/a_36_151# 0.034413f
C11735 _324_/a_224_472# _070_ 0.00142f
C11736 net20 _008_ 0.153014f
C11737 FILLER_0_17_38/a_572_375# _182_ 0.035561f
C11738 FILLER_0_17_104/a_572_375# _040_ 0.001228f
C11739 ctln[7] FILLER_0_0_130/a_124_375# 0.002726f
C11740 output10/a_224_472# _411_/a_2665_112# 0.008469f
C11741 ctln[1] vss 0.27233f
C11742 net56 fanout56/a_36_113# 0.015924f
C11743 FILLER_0_22_177/a_932_472# mask\[6\] 0.006573f
C11744 result[9] _419_/a_1308_423# 0.012036f
C11745 ctlp[9] FILLER_0_23_44/a_932_472# 0.001195f
C11746 _114_ _428_/a_2665_112# 0.002329f
C11747 net54 FILLER_0_22_107/a_572_375# 0.002239f
C11748 _068_ vdd 0.793549f
C11749 _076_ vss 1.132839f
C11750 _449_/a_2248_156# vdd -0.001225f
C11751 _449_/a_1204_472# vss 0.006048f
C11752 _205_/a_36_160# _048_ 0.040317f
C11753 _093_ _437_/a_36_151# 0.056554f
C11754 _091_ FILLER_0_17_218/a_36_472# 0.066133f
C11755 trim_mask\[4\] _386_/a_848_380# 0.001657f
C11756 _450_/a_448_472# net6 0.041113f
C11757 fanout60/a_36_160# _417_/a_36_151# 0.062739f
C11758 net63 FILLER_0_17_200/a_124_375# 0.008905f
C11759 net27 FILLER_0_14_235/a_124_375# 0.002299f
C11760 FILLER_0_17_72/a_3260_375# vss 0.052993f
C11761 FILLER_0_17_72/a_36_472# vdd 0.111688f
C11762 FILLER_0_4_49/a_124_375# net47 0.006524f
C11763 _339_/a_36_160# _140_ 0.025058f
C11764 fanout52/a_36_160# _170_ 0.024724f
C11765 _104_ mask\[7\] 0.069172f
C11766 _009_ FILLER_0_23_282/a_36_472# 0.005974f
C11767 FILLER_0_8_247/a_484_472# calibrate 0.009318f
C11768 _412_/a_36_151# net1 0.020184f
C11769 _152_ net23 0.001895f
C11770 _070_ _246_/a_36_68# 0.056186f
C11771 net60 _421_/a_448_472# 0.052759f
C11772 FILLER_0_22_86/a_36_472# vss 0.002319f
C11773 net61 fanout77/a_36_113# 0.080943f
C11774 _077_ net48 0.142015f
C11775 _418_/a_448_472# vss 0.005772f
C11776 _418_/a_1308_423# vdd 0.002258f
C11777 _093_ _177_ 0.001194f
C11778 _422_/a_1308_423# mask\[7\] 0.045368f
C11779 net52 _443_/a_1000_472# 0.016322f
C11780 _419_/a_2665_112# vdd 0.030085f
C11781 _091_ FILLER_0_15_212/a_124_375# 0.025529f
C11782 cal_count\[2\] FILLER_0_15_2/a_124_375# 0.033559f
C11783 output7/a_224_472# output40/a_224_472# 0.038066f
C11784 _426_/a_1308_423# calibrate 0.001708f
C11785 FILLER_0_21_142/a_36_472# net23 0.001629f
C11786 fanout58/a_36_160# fanout59/a_36_160# 0.001216f
C11787 _077_ _162_ 0.013298f
C11788 FILLER_0_11_142/a_124_375# FILLER_0_11_135/a_124_375# 0.004426f
C11789 _053_ net50 0.711279f
C11790 net81 en 0.071123f
C11791 _257_/a_36_472# _074_ 0.011352f
C11792 _126_ _428_/a_36_151# 0.032026f
C11793 fanout74/a_36_113# _152_ 0.017267f
C11794 fanout76/a_36_160# net18 0.003319f
C11795 _453_/a_1204_472# _042_ 0.002408f
C11796 FILLER_0_18_2/a_1916_375# net38 0.006403f
C11797 fanout53/a_36_160# _427_/a_2665_112# 0.00285f
C11798 output42/a_224_472# trim[4] 0.017153f
C11799 _402_/a_728_93# _180_ 0.008035f
C11800 ctlp[6] vdd 0.207209f
C11801 FILLER_0_16_89/a_1468_375# net14 0.022582f
C11802 FILLER_0_4_107/a_1468_375# net47 0.012534f
C11803 _086_ _395_/a_36_488# 0.00825f
C11804 _114_ _126_ 3.341247f
C11805 net4 _090_ 0.06324f
C11806 net34 FILLER_0_22_128/a_3260_375# 0.006974f
C11807 FILLER_0_4_99/a_36_472# _156_ 0.0255f
C11808 net15 FILLER_0_11_64/a_36_472# 0.020589f
C11809 net62 _045_ 0.029263f
C11810 cal_itt\[3\] calibrate 1.141592f
C11811 _413_/a_2665_112# FILLER_0_3_212/a_124_375# 0.001077f
C11812 _429_/a_448_472# net21 0.014792f
C11813 ctln[0] vss 0.125714f
C11814 FILLER_0_17_282/a_36_472# _006_ 0.002964f
C11815 mask\[7\] net22 0.275179f
C11816 FILLER_0_17_56/a_572_375# _183_ 0.002605f
C11817 net50 FILLER_0_5_88/a_36_472# 0.00867f
C11818 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_124_375# 0.004426f
C11819 _440_/a_36_151# vdd 0.117768f
C11820 net20 _128_ 0.041f
C11821 _411_/a_2665_112# cal_itt\[0\] 0.010667f
C11822 _446_/a_2665_112# net66 0.00195f
C11823 net80 FILLER_0_18_177/a_1828_472# 0.00195f
C11824 trim_mask\[2\] _035_ 0.004455f
C11825 _112_ _122_ 0.120159f
C11826 FILLER_0_5_72/a_1468_375# net49 0.001276f
C11827 _062_ _226_/a_860_68# 0.001842f
C11828 _136_ net23 0.031512f
C11829 net4 net22 0.036966f
C11830 _443_/a_448_472# _170_ 0.056211f
C11831 _139_ mask\[2\] 0.035793f
C11832 net76 FILLER_0_3_172/a_572_375# 0.003315f
C11833 FILLER_0_7_72/a_1468_375# vss 0.003253f
C11834 FILLER_0_19_47/a_484_472# _052_ 0.01589f
C11835 FILLER_0_11_78/a_484_472# vss 0.004063f
C11836 ctln[2] FILLER_0_0_266/a_36_472# 0.049163f
C11837 FILLER_0_5_72/a_484_472# trim_mask\[1\] 0.012321f
C11838 output23/a_224_472# _208_/a_36_160# 0.014541f
C11839 FILLER_0_6_47/a_2812_375# vss 0.035758f
C11840 FILLER_0_6_47/a_3260_375# vdd 0.003435f
C11841 _343_/a_665_69# _141_ 0.002451f
C11842 FILLER_0_4_197/a_932_472# net82 0.001826f
C11843 _444_/a_796_472# _054_ 0.001838f
C11844 net16 vss 0.679042f
C11845 _070_ net23 0.047632f
C11846 net48 net37 0.081653f
C11847 _414_/a_36_151# _161_ 0.033054f
C11848 FILLER_0_12_2/a_124_375# vdd 0.0247f
C11849 _432_/a_2665_112# vss 0.002577f
C11850 _317_/a_36_113# _123_ 0.037893f
C11851 _086_ calibrate 0.041755f
C11852 _188_ _453_/a_796_472# 0.00103f
C11853 FILLER_0_21_286/a_484_472# net18 0.001956f
C11854 _422_/a_1204_472# _108_ 0.015401f
C11855 ctlp[1] net77 0.716304f
C11856 net41 FILLER_0_18_37/a_124_375# 0.004639f
C11857 _419_/a_796_472# net77 0.001053f
C11858 net20 _006_ 0.014721f
C11859 _114_ FILLER_0_10_107/a_124_375# 0.004825f
C11860 fanout56/a_36_113# _095_ 0.004331f
C11861 output29/a_224_472# net29 0.038602f
C11862 FILLER_0_4_197/a_572_375# vdd 0.002455f
C11863 result[7] vss 0.49466f
C11864 FILLER_0_13_100/a_36_472# net14 0.046864f
C11865 net41 _446_/a_2248_156# 0.016492f
C11866 _072_ _395_/a_244_68# 0.001406f
C11867 FILLER_0_7_72/a_124_375# FILLER_0_6_47/a_2812_375# 0.026339f
C11868 result[7] _298_/a_224_472# 0.007724f
C11869 net73 _427_/a_36_151# 0.006328f
C11870 _119_ calibrate 0.062309f
C11871 net49 _034_ 0.031359f
C11872 FILLER_0_23_282/a_484_472# vss 0.005378f
C11873 _065_ net17 0.035195f
C11874 _111_ net71 0.002668f
C11875 net58 cal_itt\[1\] 0.79493f
C11876 trim_mask\[4\] FILLER_0_2_165/a_36_472# 0.265591f
C11877 _036_ _160_ 0.034434f
C11878 _086_ _153_ 0.017325f
C11879 _445_/a_1204_472# _034_ 0.003057f
C11880 _433_/a_1000_472# _022_ 0.05526f
C11881 _062_ FILLER_0_8_156/a_572_375# 0.002944f
C11882 ctlp[1] FILLER_0_23_290/a_36_472# 0.038596f
C11883 FILLER_0_3_221/a_124_375# net59 0.008996f
C11884 net45 vss 0.028798f
C11885 _118_ _331_/a_448_472# 0.001166f
C11886 _412_/a_2560_156# net18 0.015371f
C11887 net55 FILLER_0_11_78/a_572_375# 0.002321f
C11888 output23/a_224_472# _210_/a_67_603# 0.021084f
C11889 FILLER_0_9_142/a_36_472# net23 0.001099f
C11890 net19 net37 0.030961f
C11891 _431_/a_1308_423# _136_ 0.027758f
C11892 ctln[1] net4 0.009703f
C11893 _119_ _153_ 0.001741f
C11894 net58 sample 0.006906f
C11895 _448_/a_2665_112# vss 0.009029f
C11896 _028_ net50 0.087995f
C11897 net33 net21 0.052426f
C11898 _099_ FILLER_0_15_235/a_484_472# 0.002657f
C11899 _255_/a_224_552# vss 0.001019f
C11900 FILLER_0_9_223/a_484_472# _426_/a_2665_112# 0.004209f
C11901 net79 _417_/a_448_472# 0.028398f
C11902 FILLER_0_14_107/a_1380_472# vss 0.001338f
C11903 FILLER_0_17_161/a_124_375# mask\[2\] 0.00227f
C11904 net4 _076_ 1.140706f
C11905 _115_ FILLER_0_10_94/a_36_472# 0.014605f
C11906 net58 vss 0.589419f
C11907 _106_ net64 0.001587f
C11908 _414_/a_2665_112# _122_ 0.007441f
C11909 FILLER_0_22_177/a_1380_472# vss 0.001502f
C11910 trim[4] net6 0.002404f
C11911 _114_ _267_/a_224_472# 0.001264f
C11912 _088_ net76 0.214494f
C11913 FILLER_0_12_136/a_932_472# FILLER_0_11_142/a_124_375# 0.001543f
C11914 FILLER_0_22_177/a_1020_375# _435_/a_36_151# 0.059049f
C11915 FILLER_0_9_223/a_484_472# _060_ 0.001529f
C11916 FILLER_0_12_136/a_1020_375# cal_count\[3\] 0.002916f
C11917 _178_ _174_ 0.012157f
C11918 _423_/a_36_151# FILLER_0_23_44/a_932_472# 0.001723f
C11919 result[9] net19 0.540761f
C11920 _056_ net21 0.484506f
C11921 _431_/a_448_472# net73 0.050964f
C11922 _106_ mask\[1\] 0.005728f
C11923 _068_ _311_/a_254_473# 0.002606f
C11924 FILLER_0_15_116/a_484_472# net36 0.009319f
C11925 _427_/a_1000_472# _095_ 0.021594f
C11926 _413_/a_36_151# net82 0.00601f
C11927 _297_/a_36_472# vss 0.003601f
C11928 net68 FILLER_0_5_54/a_36_472# 0.012107f
C11929 _008_ vss 0.355468f
C11930 _074_ _078_ 0.003088f
C11931 _396_/a_224_472# _176_ 0.008359f
C11932 _354_/a_49_472# _098_ 0.009677f
C11933 FILLER_0_18_2/a_1916_375# net55 0.008235f
C11934 _133_ _154_ 0.0133f
C11935 _133_ _313_/a_67_603# 0.002974f
C11936 FILLER_0_18_139/a_124_375# FILLER_0_18_107/a_3260_375# 0.012552f
C11937 _451_/a_836_156# vdd 0.003786f
C11938 net65 FILLER_0_1_266/a_124_375# 0.002654f
C11939 FILLER_0_5_54/a_932_472# trim_mask\[1\] 0.016187f
C11940 fanout60/a_36_160# _418_/a_36_151# 0.029017f
C11941 _111_ _013_ 0.024203f
C11942 _189_/a_67_603# FILLER_0_12_220/a_1468_375# 0.029786f
C11943 _093_ _438_/a_2665_112# 0.003293f
C11944 _118_ _315_/a_244_497# 0.003007f
C11945 net60 _419_/a_36_151# 0.016173f
C11946 net61 _419_/a_1308_423# 0.00793f
C11947 output42/a_224_472# net17 0.047757f
C11948 _095_ _281_/a_234_472# 0.001467f
C11949 FILLER_0_3_172/a_36_472# FILLER_0_5_172/a_124_375# 0.0027f
C11950 FILLER_0_16_89/a_484_472# _040_ 0.009871f
C11951 net52 trim_val\[3\] 0.082691f
C11952 net82 FILLER_0_4_213/a_124_375# 0.00123f
C11953 _056_ _070_ 0.045548f
C11954 comp _190_/a_36_160# 0.001891f
C11955 FILLER_0_11_124/a_36_472# _120_ 0.014712f
C11956 output47/a_224_472# _452_/a_2225_156# 0.012077f
C11957 _443_/a_36_151# net69 0.069715f
C11958 FILLER_0_9_142/a_124_375# calibrate 0.001505f
C11959 net20 FILLER_0_13_228/a_124_375# 0.047331f
C11960 fanout61/a_36_113# net79 0.001865f
C11961 _086_ _125_ 0.490983f
C11962 net50 trim_mask\[0\] 0.002835f
C11963 _126_ _085_ 0.02154f
C11964 net27 FILLER_0_9_282/a_572_375# 0.002809f
C11965 FILLER_0_18_177/a_1380_472# vdd 0.005692f
C11966 FILLER_0_18_177/a_932_472# vss -0.001894f
C11967 _072_ _311_/a_3220_473# 0.001995f
C11968 output34/a_224_472# _421_/a_2248_156# 0.001144f
C11969 _140_ vss 0.53195f
C11970 _402_/a_56_567# net40 0.033835f
C11971 FILLER_0_5_212/a_124_375# net59 0.045135f
C11972 net52 FILLER_0_0_130/a_124_375# 0.004055f
C11973 net16 trim_mask\[2\] 0.002527f
C11974 mask\[5\] FILLER_0_20_193/a_572_375# 0.036451f
C11975 _119_ _125_ 0.11554f
C11976 output32/a_224_472# net78 0.002901f
C11977 _126_ _018_ 0.001243f
C11978 net79 net22 0.042486f
C11979 ctln[4] FILLER_0_0_232/a_36_472# 0.012298f
C11980 net16 _447_/a_1308_423# 0.001178f
C11981 ctln[9] _447_/a_36_151# 0.010503f
C11982 FILLER_0_16_57/a_1020_375# vss 0.004487f
C11983 FILLER_0_16_57/a_1468_375# vdd 0.020146f
C11984 _440_/a_36_151# FILLER_0_6_47/a_3172_472# 0.001653f
C11985 _146_ vdd 0.031209f
C11986 net17 net51 0.026974f
C11987 _092_ net31 0.04309f
C11988 FILLER_0_21_150/a_36_472# vss 0.012815f
C11989 ctln[2] net82 0.005498f
C11990 _053_ _054_ 0.015389f
C11991 net2 vdd 0.434557f
C11992 en net64 0.01789f
C11993 mask\[4\] _141_ 0.948091f
C11994 _256_/a_1612_497# _055_ 0.001438f
C11995 FILLER_0_5_198/a_36_472# net21 0.014911f
C11996 _066_ _386_/a_848_380# 0.00416f
C11997 output17/a_224_472# vdd 0.026649f
C11998 _065_ _441_/a_448_472# 0.001973f
C11999 _079_ _080_ 0.022852f
C12000 _065_ _235_/a_67_603# 0.004135f
C12001 _133_ _058_ 0.092697f
C12002 state\[2\] _427_/a_2665_112# 0.007007f
C12003 _425_/a_2665_112# net18 0.003301f
C12004 FILLER_0_23_290/a_124_375# FILLER_0_23_282/a_572_375# 0.012001f
C12005 result[9] _009_ 0.19745f
C12006 FILLER_0_5_72/a_484_472# _164_ 0.003769f
C12007 _015_ FILLER_0_8_247/a_484_472# 0.005458f
C12008 output32/a_224_472# result[5] 0.047325f
C12009 _068_ _315_/a_244_497# 0.004768f
C12010 FILLER_0_12_2/a_572_375# net6 0.058881f
C12011 _339_/a_36_160# FILLER_0_19_155/a_484_472# 0.00304f
C12012 trimb[1] FILLER_0_19_28/a_36_472# 0.01233f
C12013 mask\[0\] FILLER_0_14_235/a_572_375# 0.002003f
C12014 _238_/a_67_603# _065_ 0.005075f
C12015 _412_/a_448_472# vdd 0.011f
C12016 net21 FILLER_0_12_196/a_124_375# 0.005374f
C12017 net47 FILLER_0_5_136/a_36_472# 0.006139f
C12018 _016_ _427_/a_448_472# 0.016416f
C12019 trim_mask\[4\] _154_ 0.014658f
C12020 FILLER_0_24_290/a_36_472# vss 0.007621f
C12021 FILLER_0_5_172/a_36_472# vdd 0.092294f
C12022 FILLER_0_5_172/a_124_375# vss 0.028247f
C12023 _015_ _426_/a_1308_423# 0.029444f
C12024 FILLER_0_2_93/a_36_472# _441_/a_2665_112# 0.007491f
C12025 cal vdd 0.318671f
C12026 _128_ vss 0.859962f
C12027 _098_ mask\[2\] 0.06158f
C12028 FILLER_0_10_78/a_124_375# vss 0.006775f
C12029 _098_ _437_/a_796_472# 0.0049f
C12030 _067_ _450_/a_448_472# 0.003113f
C12031 net65 FILLER_0_3_172/a_2364_375# 0.003745f
C12032 fanout57/a_36_113# FILLER_0_3_172/a_36_472# 0.19419f
C12033 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_36_472# 0.003468f
C12034 result[5] _010_ 0.00244f
C12035 output10/a_224_472# FILLER_0_0_266/a_124_375# 0.00515f
C12036 FILLER_0_7_104/a_1468_375# _129_ 0.001165f
C12037 FILLER_0_7_104/a_36_472# _131_ 0.002019f
C12038 _323_/a_36_113# _060_ 0.002584f
C12039 net36 _438_/a_1000_472# 0.072117f
C12040 net57 _333_/a_36_160# 0.008292f
C12041 _104_ fanout63/a_36_160# 0.007014f
C12042 _386_/a_848_380# net37 0.006086f
C12043 net35 _207_/a_67_603# 0.005045f
C12044 net41 _043_ 0.03188f
C12045 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_36_472# 0.002296f
C12046 _126_ _320_/a_224_472# 0.003754f
C12047 FILLER_0_11_142/a_36_472# vdd 0.110248f
C12048 FILLER_0_11_142/a_572_375# vss 0.052505f
C12049 _149_ vss 0.005314f
C12050 FILLER_0_5_109/a_36_472# FILLER_0_4_107/a_124_375# 0.001684f
C12051 net53 _040_ 0.035628f
C12052 FILLER_0_14_99/a_36_472# _043_ 0.001242f
C12053 FILLER_0_16_89/a_1468_375# _131_ 0.016581f
C12054 net81 FILLER_0_14_235/a_484_472# 0.015266f
C12055 _088_ _083_ 0.007169f
C12056 FILLER_0_12_236/a_124_375# vss 0.001024f
C12057 FILLER_0_12_236/a_572_375# vdd 0.024713f
C12058 _119_ FILLER_0_7_162/a_124_375# 0.059009f
C12059 _114_ _060_ 0.003352f
C12060 net63 _430_/a_1000_472# 0.016386f
C12061 FILLER_0_3_78/a_36_472# _168_ 0.063262f
C12062 _161_ _228_/a_36_68# 0.055774f
C12063 net41 _185_ 0.029318f
C12064 net82 FILLER_0_3_221/a_1468_375# 0.009095f
C12065 net26 FILLER_0_18_37/a_572_375# 0.00109f
C12066 net80 _019_ 0.265857f
C12067 fanout62/a_36_160# _416_/a_36_151# 0.016215f
C12068 _074_ FILLER_0_6_231/a_36_472# 0.004325f
C12069 net41 FILLER_0_18_2/a_3172_472# 0.00982f
C12070 vdd output6/a_224_472# 0.009312f
C12071 _232_/a_67_603# net66 0.001758f
C12072 FILLER_0_7_146/a_36_472# _076_ 0.001843f
C12073 FILLER_0_7_146/a_124_375# _068_ 0.033245f
C12074 _187_ _453_/a_36_151# 0.001829f
C12075 net65 _264_/a_224_472# 0.001866f
C12076 net17 net6 0.063494f
C12077 net60 FILLER_0_17_282/a_124_375# 0.039003f
C12078 _035_ _380_/a_224_472# 0.001921f
C12079 _085_ _267_/a_224_472# 0.002907f
C12080 _176_ _267_/a_36_472# 0.001681f
C12081 net78 vdd 0.265913f
C12082 _006_ vss 0.111492f
C12083 _408_/a_1336_472# _184_ 0.003286f
C12084 _431_/a_2248_156# FILLER_0_18_139/a_932_472# 0.001148f
C12085 net48 _122_ 0.110769f
C12086 FILLER_0_6_239/a_124_375# net76 0.001286f
C12087 _392_/a_36_68# FILLER_0_12_50/a_36_472# 0.002811f
C12088 _132_ _135_ 0.345161f
C12089 _430_/a_1308_423# net21 0.008506f
C12090 _415_/a_1000_472# net19 0.001125f
C12091 FILLER_0_15_282/a_124_375# net18 0.048284f
C12092 FILLER_0_16_73/a_124_375# FILLER_0_16_57/a_1468_375# 0.012222f
C12093 vss output40/a_224_472# 0.002459f
C12094 net58 net4 0.858616f
C12095 mask\[7\] _297_/a_36_472# 0.003196f
C12096 _161_ calibrate 0.044443f
C12097 FILLER_0_21_28/a_3260_375# vss 0.054959f
C12098 FILLER_0_21_28/a_36_472# vdd 0.090954f
C12099 net20 net82 0.026007f
C12100 FILLER_0_3_172/a_2724_472# vdd 0.006405f
C12101 net79 _418_/a_448_472# 0.034736f
C12102 mask\[8\] _436_/a_36_151# 0.032521f
C12103 FILLER_0_8_2/a_36_472# vss 0.004429f
C12104 _427_/a_1000_472# net74 0.009646f
C12105 fanout57/a_36_113# vss 0.046378f
C12106 FILLER_0_21_28/a_1380_472# net17 0.001709f
C12107 output42/a_224_472# net39 0.027208f
C12108 net81 FILLER_0_8_263/a_36_472# 0.007373f
C12109 result[5] vdd 0.142481f
C12110 _398_/a_36_113# _043_ 0.005985f
C12111 FILLER_0_22_177/a_484_472# net33 0.013149f
C12112 _232_/a_67_603# _167_ 0.014152f
C12113 _053_ net22 0.039386f
C12114 net68 _453_/a_448_472# 0.01245f
C12115 output42/a_224_472# _039_ 0.001254f
C12116 _391_/a_245_68# cal_count\[0\] 0.001201f
C12117 net15 FILLER_0_15_72/a_572_375# 0.002741f
C12118 _077_ FILLER_0_10_78/a_1020_375# 0.001131f
C12119 net15 net52 0.166073f
C12120 _091_ FILLER_0_12_220/a_484_472# 0.001453f
C12121 FILLER_0_17_72/a_1020_375# _131_ 0.005847f
C12122 _439_/a_36_151# net51 0.00711f
C12123 FILLER_0_17_64/a_36_472# vdd 0.094397f
C12124 FILLER_0_17_64/a_124_375# vss 0.022351f
C12125 FILLER_0_4_49/a_124_375# vdd 0.008637f
C12126 FILLER_0_7_72/a_2724_472# net14 0.012436f
C12127 _414_/a_2560_156# net22 0.00603f
C12128 _127_ _395_/a_36_488# 0.00519f
C12129 _140_ mask\[7\] 0.064343f
C12130 FILLER_0_10_78/a_36_472# _115_ 0.002611f
C12131 _111_ _110_ 0.00195f
C12132 FILLER_0_5_72/a_1468_375# net47 0.005049f
C12133 result[6] FILLER_0_21_286/a_36_472# 0.015369f
C12134 net61 net19 0.132027f
C12135 _140_ _148_ 0.011699f
C12136 FILLER_0_2_177/a_36_472# net22 0.002517f
C12137 _162_ _061_ 0.001665f
C12138 mask\[4\] FILLER_0_17_218/a_484_472# 0.001232f
C12139 _428_/a_36_151# _095_ 0.006658f
C12140 FILLER_0_20_177/a_572_375# _434_/a_36_151# 0.059049f
C12141 _401_/a_36_68# _179_ 0.007074f
C12142 FILLER_0_3_204/a_124_375# net82 0.014222f
C12143 _077_ FILLER_0_11_64/a_36_472# 0.076102f
C12144 FILLER_0_15_150/a_36_472# net36 0.012318f
C12145 _147_ vdd 0.09215f
C12146 FILLER_0_0_266/a_36_472# vss 0.003738f
C12147 net51 _039_ 0.398642f
C12148 net15 _216_/a_67_603# 0.060076f
C12149 net63 FILLER_0_22_177/a_932_472# 0.060639f
C12150 ctlp[3] vdd 0.251098f
C12151 net38 _452_/a_2225_156# 0.034415f
C12152 output11/a_224_472# FILLER_0_0_198/a_124_375# 0.00363f
C12153 FILLER_0_16_73/a_484_472# net55 0.004188f
C12154 FILLER_0_3_78/a_572_375# vdd 0.014442f
C12155 FILLER_0_3_78/a_124_375# vss 0.004739f
C12156 _114_ _095_ 0.001338f
C12157 output39/a_224_472# _444_/a_36_151# 0.062717f
C12158 FILLER_0_8_37/a_572_375# _220_/a_67_603# 0.00744f
C12159 _452_/a_448_472# net40 0.047031f
C12160 _321_/a_170_472# vdd 0.060585f
C12161 FILLER_0_13_228/a_36_472# vdd 0.085375f
C12162 FILLER_0_13_228/a_124_375# vss 0.007465f
C12163 FILLER_0_2_101/a_36_472# vdd 0.099518f
C12164 FILLER_0_2_101/a_124_375# vss 0.04897f
C12165 FILLER_0_4_107/a_1468_375# vdd 0.023541f
C12166 _155_ _053_ 0.122798f
C12167 _077_ _439_/a_1204_472# 0.016471f
C12168 _104_ ctlp[2] 1.420577f
C12169 fanout57/a_36_113# FILLER_0_2_165/a_124_375# 0.008057f
C12170 _395_/a_36_488# _071_ 0.00276f
C12171 _435_/a_448_472# vdd 0.029967f
C12172 trimb[1] FILLER_0_20_15/a_484_472# 0.001292f
C12173 FILLER_0_12_20/a_572_375# net17 0.041149f
C12174 fanout72/a_36_113# _174_ 0.026207f
C12175 _013_ _424_/a_1308_423# 0.007751f
C12176 FILLER_0_9_72/a_1020_375# _439_/a_36_151# 0.059049f
C12177 _259_/a_455_68# net37 0.0023f
C12178 net31 vdd 0.542738f
C12179 output19/a_224_472# _422_/a_2665_112# 0.024396f
C12180 input1/a_36_113# input2/a_36_113# 0.029417f
C12181 _086_ _069_ 0.580351f
C12182 _077_ _055_ 0.083808f
C12183 _221_/a_36_160# _054_ 0.02124f
C12184 net47 _034_ 0.052602f
C12185 _093_ FILLER_0_17_72/a_2724_472# 0.02416f
C12186 net20 _098_ 0.087341f
C12187 FILLER_0_17_226/a_124_375# net20 0.001895f
C12188 net72 FILLER_0_17_64/a_36_472# 0.001145f
C12189 result[6] ctlp[2] 0.001324f
C12190 _063_ vss 0.157186f
C12191 FILLER_0_21_28/a_1916_375# _423_/a_36_151# 0.001597f
C12192 _369_/a_692_472# _157_ 0.0025f
C12193 _127_ calibrate 0.004656f
C12194 fanout49/a_36_160# FILLER_0_5_88/a_124_375# 0.001154f
C12195 vdd FILLER_0_21_60/a_572_375# 0.022291f
C12196 vss FILLER_0_21_60/a_124_375# 0.003723f
C12197 FILLER_0_1_212/a_124_375# net11 0.029766f
C12198 _130_ FILLER_0_11_135/a_124_375# 0.001198f
C12199 net54 _438_/a_2248_156# 0.014423f
C12200 _451_/a_36_151# _040_ 0.018648f
C12201 net52 _376_/a_36_160# 0.00267f
C12202 FILLER_0_9_290/a_124_375# vdd 0.028723f
C12203 _119_ _069_ 0.00226f
C12204 net63 FILLER_0_18_177/a_484_472# 0.061539f
C12205 _053_ _076_ 0.108358f
C12206 FILLER_0_5_206/a_124_375# vdd 0.038311f
C12207 _139_ vss 0.052996f
C12208 _128_ net4 0.039671f
C12209 net20 FILLER_0_13_212/a_1380_472# 0.006746f
C12210 FILLER_0_12_28/a_36_472# net40 0.020589f
C12211 net26 FILLER_0_23_44/a_124_375# 0.007775f
C12212 FILLER_0_13_290/a_124_375# _416_/a_36_151# 0.026277f
C12213 en_co_clk fanout55/a_36_160# 0.041263f
C12214 _052_ FILLER_0_19_28/a_484_472# 0.003325f
C12215 _430_/a_36_151# _069_ 0.026308f
C12216 FILLER_0_18_100/a_124_375# net14 0.04037f
C12217 fanout56/a_36_113# _097_ 0.062226f
C12218 fanout80/a_36_113# _138_ 0.002489f
C12219 _408_/a_718_524# _043_ 0.003719f
C12220 net38 _064_ 0.02996f
C12221 FILLER_0_19_28/a_124_375# net17 0.007234f
C12222 _288_/a_224_472# net19 0.002252f
C12223 _077_ _313_/a_67_603# 0.007446f
C12224 net61 _009_ 0.042703f
C12225 _345_/a_36_160# FILLER_0_19_111/a_484_472# 0.007907f
C12226 FILLER_0_19_155/a_484_472# vss 0.004002f
C12227 _144_ mask\[8\] 0.131592f
C12228 net81 _018_ 0.081888f
C12229 _149_ _148_ 0.001124f
C12230 _306_/a_36_68# _113_ 0.010109f
C12231 net41 _402_/a_1296_93# 0.001707f
C12232 _323_/a_36_113# net64 0.06154f
C12233 FILLER_0_5_117/a_36_472# _360_/a_36_160# 0.003913f
C12234 FILLER_0_5_54/a_36_472# net47 0.00679f
C12235 net14 FILLER_0_4_91/a_484_472# 0.020589f
C12236 net16 _380_/a_224_472# 0.008718f
C12237 net29 _005_ 0.020239f
C12238 net82 FILLER_0_3_172/a_36_472# 0.007612f
C12239 net4 FILLER_0_12_236/a_124_375# 0.001558f
C12240 net73 FILLER_0_17_142/a_484_472# 0.001122f
C12241 output32/a_224_472# net60 0.191561f
C12242 _185_ cal_count\[2\] 0.205002f
C12243 _033_ trim_mask\[1\] 0.001251f
C12244 _173_ _042_ 0.002294f
C12245 FILLER_0_17_142/a_124_375# vdd 0.020936f
C12246 _158_ vss 0.007784f
C12247 fanout62/a_36_160# result[1] 0.036633f
C12248 net62 output28/a_224_472# 0.206137f
C12249 net28 vdd 0.489756f
C12250 _039_ net6 0.104745f
C12251 net57 FILLER_0_13_100/a_124_375# 0.012636f
C12252 FILLER_0_17_72/a_1468_375# _150_ 0.001076f
C12253 net61 fanout78/a_36_113# 0.056484f
C12254 net18 _419_/a_1000_472# 0.008295f
C12255 _137_ FILLER_0_16_154/a_484_472# 0.00631f
C12256 _411_/a_2665_112# net10 0.007912f
C12257 FILLER_0_8_127/a_36_472# _129_ 0.060819f
C12258 net57 _072_ 0.108982f
C12259 FILLER_0_17_200/a_484_472# vss 0.003134f
C12260 _093_ FILLER_0_19_142/a_36_472# 0.002415f
C12261 _292_/a_36_160# output18/a_224_472# 0.009736f
C12262 output31/a_224_472# net19 0.072666f
C12263 _142_ _137_ 1.401722f
C12264 FILLER_0_5_109/a_36_472# _153_ 0.034328f
C12265 _415_/a_36_151# result[1] 0.012965f
C12266 mask\[5\] ctlp[4] 0.001643f
C12267 net15 FILLER_0_18_61/a_124_375# 0.001179f
C12268 mask\[9\] FILLER_0_20_87/a_36_472# 0.00596f
C12269 FILLER_0_19_55/a_36_472# _052_ 0.019665f
C12270 net60 _010_ 0.108311f
C12271 result[0] FILLER_0_9_282/a_572_375# 0.042859f
C12272 _007_ vss 0.017377f
C12273 net62 net77 0.122747f
C12274 net64 FILLER_0_14_235/a_484_472# 0.012355f
C12275 _429_/a_1000_472# vss 0.006901f
C12276 _176_ _118_ 0.392531f
C12277 _423_/a_1308_423# vss 0.001726f
C12278 _423_/a_796_472# vdd 0.001494f
C12279 net52 trim_mask\[4\] 0.034276f
C12280 net57 net70 0.012088f
C12281 FILLER_0_10_247/a_124_375# vdd 0.040502f
C12282 _024_ _147_ 0.006801f
C12283 net82 cal_itt\[1\] 0.396149f
C12284 vss net14 1.003274f
C12285 FILLER_0_19_28/a_124_375# _452_/a_36_151# 0.002709f
C12286 net57 net47 0.279638f
C12287 fanout51/a_36_113# FILLER_0_9_72/a_36_472# 0.001391f
C12288 FILLER_0_17_72/a_1380_472# net36 0.021039f
C12289 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_124_375# 0.012001f
C12290 net52 FILLER_0_11_78/a_36_472# 0.005678f
C12291 net41 _033_ 0.033812f
C12292 FILLER_0_8_127/a_124_375# _125_ 0.003105f
C12293 mask\[4\] FILLER_0_17_200/a_36_472# 0.001242f
C12294 trim_mask\[2\] FILLER_0_3_78/a_124_375# 0.010185f
C12295 _372_/a_2590_472# _059_ 0.002974f
C12296 _077_ _058_ 3.018054f
C12297 FILLER_0_17_161/a_124_375# vss 0.00824f
C12298 FILLER_0_17_161/a_36_472# vdd 0.006972f
C12299 net52 FILLER_0_6_47/a_2364_375# 0.002577f
C12300 FILLER_0_22_128/a_36_472# vdd 0.004601f
C12301 FILLER_0_22_128/a_3260_375# vss 0.006346f
C12302 _297_/a_36_472# _295_/a_36_472# 0.004259f
C12303 _281_/a_234_472# _097_ 0.004169f
C12304 _328_/a_36_113# _428_/a_36_151# 0.030244f
C12305 net32 _421_/a_36_151# 0.008275f
C12306 ctln[2] clk 0.004558f
C12307 _127_ _125_ 0.053419f
C12308 _422_/a_36_151# _109_ 0.036674f
C12309 output42/a_224_472# net42 0.117956f
C12310 _155_ _028_ 0.049284f
C12311 _424_/a_2665_112# vdd 0.013636f
C12312 _424_/a_2248_156# vss 0.004855f
C12313 _024_ _435_/a_448_472# 0.039244f
C12314 result[6] _420_/a_1308_423# 0.008756f
C12315 FILLER_0_7_72/a_1468_375# _053_ 0.014569f
C12316 _093_ _291_/a_36_160# 0.017281f
C12317 mask\[5\] FILLER_0_20_177/a_932_472# 0.016114f
C12318 _442_/a_36_151# vdd 0.102701f
C12319 net55 _452_/a_2225_156# 0.022788f
C12320 net66 net17 0.023639f
C12321 _031_ trim_mask\[3\] 0.016747f
C12322 _053_ FILLER_0_6_47/a_2812_375# 0.003818f
C12323 mask\[3\] FILLER_0_18_177/a_2276_472# 0.01204f
C12324 _447_/a_2665_112# vss 0.012813f
C12325 _412_/a_2248_156# net1 0.044934f
C12326 _328_/a_36_113# _114_ 0.058671f
C12327 net23 FILLER_0_5_148/a_36_472# 0.011079f
C12328 _320_/a_1120_472# _090_ 0.001215f
C12329 _187_ _095_ 0.00765f
C12330 _141_ _140_ 0.131685f
C12331 net82 vss 0.550252f
C12332 _414_/a_36_151# _056_ 0.00356f
C12333 _154_ _157_ 0.447829f
C12334 FILLER_0_15_290/a_124_375# output30/a_224_472# 0.02894f
C12335 _258_/a_36_160# _078_ 0.006096f
C12336 FILLER_0_8_263/a_36_472# net64 0.00399f
C12337 net3 vss 0.02666f
C12338 _445_/a_1308_423# net17 0.002172f
C12339 FILLER_0_15_116/a_36_472# net70 0.051129f
C12340 _428_/a_36_151# net74 0.020444f
C12341 ctln[1] ctln[3] 0.926618f
C12342 _431_/a_36_151# FILLER_0_17_133/a_36_472# 0.001723f
C12343 fanout82/a_36_113# output37/a_224_472# 0.023409f
C12344 FILLER_0_7_162/a_36_472# calibrate 0.014431f
C12345 mask\[5\] FILLER_0_18_177/a_572_375# 0.002653f
C12346 _430_/a_2248_156# _092_ 0.003124f
C12347 FILLER_0_16_107/a_36_472# _132_ 0.001538f
C12348 FILLER_0_9_28/a_3260_375# net51 0.001597f
C12349 _422_/a_36_151# _421_/a_2248_156# 0.001189f
C12350 _132_ net57 0.029479f
C12351 _074_ _265_/a_224_472# 0.001223f
C12352 output42/a_224_472# clkc 0.004924f
C12353 net55 _423_/a_36_151# 0.001124f
C12354 _114_ net74 0.559239f
C12355 net82 FILLER_0_2_171/a_124_375# 0.003818f
C12356 _141_ FILLER_0_21_150/a_36_472# 0.002773f
C12357 net65 net76 0.14935f
C12358 output12/a_224_472# ctln[4] 0.041517f
C12359 _449_/a_2248_156# _176_ 0.013753f
C12360 mask\[7\] _435_/a_36_151# 0.037736f
C12361 result[6] _421_/a_1000_472# 0.024206f
C12362 net60 vdd 0.575502f
C12363 net81 _426_/a_36_151# 0.060652f
C12364 FILLER_0_13_228/a_124_375# net4 0.002641f
C12365 FILLER_0_16_255/a_36_472# net36 0.034335f
C12366 mask\[5\] _348_/a_49_472# 0.025962f
C12367 net50 FILLER_0_2_93/a_572_375# 0.00275f
C12368 net52 FILLER_0_2_93/a_484_472# 0.009006f
C12369 FILLER_0_12_20/a_572_375# _039_ 0.005679f
C12370 _211_/a_36_160# _436_/a_36_151# 0.068534f
C12371 net74 _443_/a_36_151# 0.003682f
C12372 _059_ _242_/a_36_160# 0.001942f
C12373 net35 _435_/a_2665_112# 0.007912f
C12374 _449_/a_36_151# _453_/a_36_151# 0.007757f
C12375 _142_ net56 0.028797f
C12376 net52 _448_/a_2248_156# 0.002555f
C12377 FILLER_0_17_200/a_124_375# net21 0.048656f
C12378 _067_ net17 0.17227f
C12379 net55 _424_/a_1000_472# 0.001357f
C12380 _269_/a_36_472# _080_ 0.003981f
C12381 _083_ _260_/a_36_68# 0.047191f
C12382 ctln[6] net13 0.065837f
C12383 FILLER_0_17_226/a_36_472# _291_/a_36_160# 0.035111f
C12384 FILLER_0_4_107/a_572_375# _154_ 0.052251f
C12385 FILLER_0_16_107/a_124_375# net36 0.001706f
C12386 net36 FILLER_0_16_115/a_124_375# 0.001706f
C12387 _310_/a_49_472# _060_ 0.001122f
C12388 _189_/a_67_603# vdd 0.01494f
C12389 FILLER_0_21_133/a_36_472# FILLER_0_21_142/a_36_472# 0.001963f
C12390 FILLER_0_20_15/a_124_375# vdd 0.006513f
C12391 net76 net59 3.439686f
C12392 _426_/a_2665_112# FILLER_0_8_239/a_124_375# 0.010736f
C12393 net17 FILLER_0_20_15/a_1468_375# 0.010099f
C12394 _132_ FILLER_0_15_116/a_36_472# 0.020589f
C12395 _074_ _317_/a_36_113# 0.003383f
C12396 net16 FILLER_0_10_28/a_124_375# 0.002225f
C12397 FILLER_0_15_205/a_124_375# vss 0.026372f
C12398 FILLER_0_15_205/a_36_472# vdd 0.010089f
C12399 FILLER_0_5_136/a_124_375# vss 0.053395f
C12400 FILLER_0_5_136/a_36_472# vdd 0.092379f
C12401 FILLER_0_23_290/a_124_375# net77 0.001783f
C12402 net79 FILLER_0_12_236/a_124_375# 0.010367f
C12403 valid net18 0.03851f
C12404 FILLER_0_5_198/a_572_375# net37 0.009149f
C12405 FILLER_0_14_263/a_36_472# net30 0.003972f
C12406 FILLER_0_1_98/a_36_472# net14 0.023583f
C12407 _098_ vss 0.958032f
C12408 FILLER_0_17_226/a_124_375# vss 0.025007f
C12409 FILLER_0_3_54/a_36_472# _160_ 0.00702f
C12410 trim_mask\[2\] net14 0.060278f
C12411 _135_ vdd 0.018662f
C12412 FILLER_0_17_56/a_36_472# vss 0.00167f
C12413 FILLER_0_17_56/a_484_472# vdd 0.002789f
C12414 net23 FILLER_0_22_128/a_2364_375# 0.018463f
C12415 net79 _006_ 0.050445f
C12416 _137_ mask\[2\] 0.440828f
C12417 cal_count\[2\] _402_/a_1296_93# 0.022009f
C12418 net44 FILLER_0_12_2/a_124_375# 0.01836f
C12419 _101_ _196_/a_36_160# 0.009836f
C12420 _134_ FILLER_0_9_105/a_124_375# 0.005919f
C12421 cal_count\[3\] FILLER_0_9_72/a_484_472# 0.004129f
C12422 _448_/a_448_472# _037_ 0.044085f
C12423 _033_ _164_ 0.007117f
C12424 _444_/a_36_151# net40 0.032012f
C12425 cal_itt\[3\] net22 0.134309f
C12426 fanout53/a_36_160# _136_ 0.001471f
C12427 FILLER_0_13_212/a_1380_472# vss 0.010223f
C12428 net62 FILLER_0_13_212/a_484_472# 0.059367f
C12429 _069_ _161_ 0.017831f
C12430 _012_ FILLER_0_23_44/a_484_472# 0.001572f
C12431 _436_/a_2665_112# vss 0.007905f
C12432 _441_/a_448_472# net66 0.023761f
C12433 FILLER_0_7_72/a_1468_375# _028_ 0.003785f
C12434 net42 net6 0.166896f
C12435 _081_ net22 0.103561f
C12436 net73 FILLER_0_18_139/a_484_472# 0.00131f
C12437 _028_ FILLER_0_6_47/a_2812_375# 0.023189f
C12438 FILLER_0_7_195/a_36_472# _062_ 0.0045f
C12439 vss _433_/a_2248_156# 0.034403f
C12440 vdd _433_/a_2665_112# 0.002569f
C12441 _181_ _401_/a_36_68# 0.010647f
C12442 FILLER_0_18_139/a_1020_375# vdd 0.001285f
C12443 FILLER_0_18_139/a_572_375# vss 0.009977f
C12444 net41 FILLER_0_16_37/a_124_375# 0.008195f
C12445 FILLER_0_1_204/a_124_375# net59 0.00999f
C12446 _018_ mask\[1\] 0.001206f
C12447 net49 _440_/a_1308_423# 0.022006f
C12448 net19 net8 0.056454f
C12449 _369_/a_36_68# _153_ 0.008048f
C12450 _065_ FILLER_0_1_98/a_124_375# 0.001136f
C12451 _086_ _090_ 0.065807f
C12452 _132_ FILLER_0_17_104/a_1380_472# 0.02114f
C12453 output23/a_224_472# vdd 0.033718f
C12454 _273_/a_36_68# vdd 0.041825f
C12455 net57 state\[1\] 0.154183f
C12456 mask\[7\] FILLER_0_22_128/a_3260_375# 0.00186f
C12457 calibrate net23 0.032259f
C12458 mask\[3\] _093_ 2.443356f
C12459 _427_/a_36_151# FILLER_0_14_123/a_124_375# 0.023595f
C12460 _067_ FILLER_0_12_28/a_124_375# 0.012779f
C12461 _431_/a_448_472# net36 0.010914f
C12462 net35 FILLER_0_22_128/a_2724_472# 0.012359f
C12463 net6 clkc 0.036083f
C12464 _270_/a_36_472# net22 0.002857f
C12465 input3/a_36_113# net3 0.015124f
C12466 output39/a_224_472# net49 0.039256f
C12467 _011_ _299_/a_36_472# 0.004407f
C12468 net36 _451_/a_2225_156# 0.044144f
C12469 net55 FILLER_0_17_56/a_124_375# 0.014472f
C12470 net72 FILLER_0_17_56/a_484_472# 0.003359f
C12471 FILLER_0_12_220/a_36_472# _248_/a_36_68# 0.006596f
C12472 _256_/a_36_68# _056_ 0.008305f
C12473 _077_ net52 0.047585f
C12474 net73 FILLER_0_18_107/a_1020_375# 0.04487f
C12475 _086_ net22 0.00117f
C12476 net68 FILLER_0_6_47/a_484_472# 0.005391f
C12477 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_36_472# 0.009654f
C12478 output46/a_224_472# FILLER_0_21_28/a_36_472# 0.010684f
C12479 output38/a_224_472# _034_ 0.039873f
C12480 output15/a_224_472# ctln[8] 0.079231f
C12481 trim_mask\[1\] FILLER_0_6_47/a_1380_472# 0.006166f
C12482 trim[1] _445_/a_36_151# 0.008362f
C12483 net39 _445_/a_1308_423# 0.008252f
C12484 _363_/a_244_472# vdd 0.002075f
C12485 FILLER_0_7_72/a_3172_472# _058_ 0.001085f
C12486 _383_/a_36_472# vdd -0.002154f
C12487 _414_/a_1204_472# net21 0.007637f
C12488 FILLER_0_11_101/a_36_472# _070_ 0.033113f
C12489 net82 net4 1.982825f
C12490 _327_/a_36_472# _130_ 0.001474f
C12491 FILLER_0_4_197/a_484_472# net22 0.007955f
C12492 fanout68/a_36_113# net68 0.027807f
C12493 _104_ ctlp[1] 0.076863f
C12494 FILLER_0_13_228/a_124_375# net79 0.008554f
C12495 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_36_472# 0.009654f
C12496 _432_/a_2665_112# FILLER_0_17_200/a_36_472# 0.007491f
C12497 _446_/a_1000_472# vdd 0.001598f
C12498 ctlp[1] _421_/a_2665_112# 0.008695f
C12499 net55 _040_ 0.107198f
C12500 _065_ _030_ 0.001499f
C12501 fanout65/a_36_113# net64 0.002858f
C12502 state\[2\] FILLER_0_13_142/a_1020_375# 0.007311f
C12503 net53 FILLER_0_13_142/a_36_472# 0.059367f
C12504 _425_/a_36_151# _316_/a_848_380# 0.035903f
C12505 _091_ FILLER_0_10_214/a_124_375# 0.006331f
C12506 FILLER_0_5_72/a_1020_375# vss 0.004157f
C12507 FILLER_0_5_72/a_1468_375# vdd 0.001826f
C12508 _430_/a_36_151# net22 0.005321f
C12509 _446_/a_2665_112# net17 0.00149f
C12510 cal_itt\[3\] _076_ 0.002726f
C12511 _114_ _097_ 0.004412f
C12512 net56 mask\[2\] 0.090254f
C12513 net54 FILLER_0_19_142/a_124_375# 0.056556f
C12514 net58 ctln[3] 0.00479f
C12515 fanout60/a_36_160# net61 0.001167f
C12516 FILLER_0_13_212/a_36_472# _429_/a_1308_423# 0.009119f
C12517 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1380_472# 0.013276f
C12518 _083_ net59 0.408831f
C12519 _127_ _069_ 0.048146f
C12520 _056_ _228_/a_36_68# 0.043669f
C12521 result[6] ctlp[1] 0.677825f
C12522 _430_/a_2248_156# vdd 0.008989f
C12523 _076_ _081_ 0.010091f
C12524 _133_ _152_ 0.124374f
C12525 net52 _066_ 0.022601f
C12526 FILLER_0_17_226/a_36_472# mask\[3\] 0.011509f
C12527 FILLER_0_3_204/a_36_472# net21 0.01535f
C12528 output10/a_224_472# net8 0.010088f
C12529 FILLER_0_6_90/a_124_375# _163_ 0.013948f
C12530 _408_/a_1336_472# vdd 0.040992f
C12531 fanout61/a_36_113# ctlp[1] 0.019606f
C12532 _417_/a_2665_112# net30 0.015638f
C12533 FILLER_0_16_89/a_1380_472# _136_ 0.009079f
C12534 _067_ _039_ 0.221585f
C12535 FILLER_0_7_104/a_1380_472# _133_ 0.004838f
C12536 trim_val\[3\] FILLER_0_2_93/a_36_472# 0.015653f
C12537 FILLER_0_12_136/a_484_472# _126_ 0.014541f
C12538 trim_val\[1\] FILLER_0_6_37/a_36_472# 0.011347f
C12539 _405_/a_67_603# vss 0.008564f
C12540 _405_/a_255_603# vdd 0.001044f
C12541 net81 mask\[2\] 0.002083f
C12542 net64 FILLER_0_8_247/a_1468_375# 0.002559f
C12543 _013_ _216_/a_67_603# 0.006454f
C12544 FILLER_0_8_127/a_36_472# _322_/a_124_24# 0.00171f
C12545 _436_/a_2665_112# FILLER_0_22_128/a_1020_375# 0.029834f
C12546 _372_/a_170_472# vss 0.027819f
C12547 net15 _449_/a_796_472# 0.006722f
C12548 _129_ vdd 0.314544f
C12549 _061_ _055_ 0.853642f
C12550 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_484_472# 0.013276f
C12551 _094_ _418_/a_2560_156# 0.011088f
C12552 _131_ vss 0.549133f
C12553 FILLER_0_8_24/a_572_375# net17 0.007101f
C12554 FILLER_0_21_125/a_124_375# net54 0.008377f
C12555 _056_ calibrate 0.00931f
C12556 FILLER_0_22_128/a_36_472# _433_/a_36_151# 0.001653f
C12557 _426_/a_36_151# net64 0.022056f
C12558 FILLER_0_20_177/a_572_375# mask\[6\] 0.001158f
C12559 _274_/a_3368_68# vss 0.001714f
C12560 vdd _034_ 0.424437f
C12561 FILLER_0_10_256/a_124_375# _015_ 0.001151f
C12562 _185_ _402_/a_56_567# 0.107713f
C12563 net26 net17 0.132516f
C12564 _086_ _076_ 0.79237f
C12565 _075_ _077_ 0.004518f
C12566 _431_/a_36_151# net53 0.001579f
C12567 _141_ FILLER_0_19_155/a_484_472# 0.015625f
C12568 FILLER_0_16_89/a_932_472# FILLER_0_17_72/a_2812_375# 0.001723f
C12569 net52 _157_ 0.005889f
C12570 net58 _425_/a_2248_156# 0.051603f
C12571 FILLER_0_18_139/a_484_472# FILLER_0_19_142/a_124_375# 0.001723f
C12572 output36/a_224_472# output30/a_224_472# 0.003578f
C12573 _119_ _076_ 0.083673f
C12574 _415_/a_2248_156# FILLER_0_11_282/a_124_375# 0.001221f
C12575 _449_/a_1308_423# _038_ 0.021006f
C12576 output9/a_224_472# net76 0.002042f
C12577 FILLER_0_16_57/a_1468_375# _176_ 0.006445f
C12578 FILLER_0_18_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001684f
C12579 FILLER_0_15_150/a_124_375# net36 0.005687f
C12580 _277_/a_36_160# net30 0.014059f
C12581 _339_/a_36_160# FILLER_0_19_171/a_36_472# 0.195478f
C12582 net57 _385_/a_36_68# 0.03315f
C12583 mask\[7\] _436_/a_2665_112# 0.004274f
C12584 net81 ctln[2] 0.003762f
C12585 _449_/a_36_151# _095_ 0.003412f
C12586 net31 _099_ 0.01086f
C12587 FILLER_0_17_72/a_2812_375# _136_ 0.017702f
C12588 fanout70/a_36_113# net70 0.073707f
C12589 net16 _178_ 0.30147f
C12590 _144_ _145_ 0.671767f
C12591 _025_ _436_/a_1204_472# 0.01349f
C12592 result[7] _421_/a_1000_472# 0.015328f
C12593 net79 _007_ 0.096772f
C12594 _428_/a_2665_112# vss 0.005991f
C12595 net27 fanout62/a_36_160# 0.005558f
C12596 trim_mask\[4\] _152_ 0.224909f
C12597 FILLER_0_5_54/a_36_472# vdd 0.006056f
C12598 FILLER_0_5_54/a_1468_375# vss 0.053407f
C12599 net34 result[8] 0.076645f
C12600 trimb[1] FILLER_0_20_2/a_572_375# 0.003431f
C12601 _058_ _122_ 0.040376f
C12602 FILLER_0_20_31/a_124_375# net40 0.011967f
C12603 _070_ _133_ 0.436976f
C12604 _093_ FILLER_0_17_218/a_124_375# 0.003338f
C12605 _441_/a_36_151# _164_ 0.008955f
C12606 clk vss 0.210484f
C12607 mask\[5\] _143_ 0.032539f
C12608 _412_/a_796_472# net1 0.002922f
C12609 net68 _042_ 0.037716f
C12610 net27 _415_/a_36_151# 0.019856f
C12611 _413_/a_36_151# _079_ 0.0017f
C12612 FILLER_0_10_214/a_36_472# _069_ 0.085701f
C12613 result[8] FILLER_0_24_274/a_932_472# 0.005458f
C12614 cal_itt\[0\] net8 0.026229f
C12615 FILLER_0_21_28/a_3172_472# FILLER_0_21_60/a_36_472# 0.013276f
C12616 _095_ FILLER_0_13_100/a_36_472# 0.003036f
C12617 net82 FILLER_0_3_142/a_36_472# 0.0172f
C12618 _414_/a_2665_112# _068_ 0.002324f
C12619 FILLER_0_16_37/a_124_375# cal_count\[2\] 0.008393f
C12620 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_572_375# 0.086635f
C12621 _074_ _375_/a_36_68# 0.003157f
C12622 vdd output30/a_224_472# 0.068123f
C12623 _327_/a_36_472# _428_/a_2248_156# 0.001757f
C12624 net44 output6/a_224_472# 0.078248f
C12625 _064_ _446_/a_36_151# 0.006723f
C12626 _235_/a_67_603# _446_/a_2665_112# 0.017036f
C12627 _122_ FILLER_0_5_198/a_572_375# 0.001352f
C12628 _443_/a_2665_112# vss 0.007913f
C12629 _073_ _078_ 0.098575f
C12630 FILLER_0_19_28/a_484_472# net40 0.020293f
C12631 _141_ FILLER_0_17_161/a_124_375# 0.040332f
C12632 vss FILLER_0_3_212/a_36_472# 0.00838f
C12633 _173_ _120_ 0.004205f
C12634 _141_ FILLER_0_22_128/a_3260_375# 0.003544f
C12635 result[1] _416_/a_1000_472# 0.001529f
C12636 net28 _416_/a_2248_156# 0.001082f
C12637 _446_/a_36_151# output41/a_224_472# 0.135198f
C12638 _448_/a_448_472# FILLER_0_3_172/a_572_375# 0.00123f
C12639 _448_/a_36_151# FILLER_0_3_172/a_1020_375# 0.001512f
C12640 net17 FILLER_0_23_44/a_124_375# 0.007634f
C12641 _013_ FILLER_0_18_61/a_124_375# 0.016976f
C12642 _410_/a_36_68# _188_ 0.007731f
C12643 FILLER_0_16_107/a_36_472# vdd 0.110244f
C12644 net20 _420_/a_2665_112# 0.030202f
C12645 net15 FILLER_0_6_47/a_1916_375# 0.029774f
C12646 FILLER_0_11_101/a_484_472# FILLER_0_11_109/a_36_472# 0.013276f
C12647 _431_/a_1000_472# vss 0.002491f
C12648 net69 FILLER_0_3_54/a_124_375# 0.004245f
C12649 net22 _204_/a_67_603# 0.006495f
C12650 _091_ _429_/a_36_151# 0.006557f
C12651 _061_ _058_ 0.02828f
C12652 net19 _420_/a_2248_156# 0.058662f
C12653 _075_ net37 0.001054f
C12654 _275_/a_224_472# vss 0.001498f
C12655 net57 vdd 1.260693f
C12656 _000_ _074_ 0.003542f
C12657 net58 fanout81/a_36_160# 0.013959f
C12658 FILLER_0_4_185/a_124_375# _272_/a_36_472# 0.001781f
C12659 _076_ FILLER_0_9_142/a_124_375# 0.001774f
C12660 output35/a_224_472# _435_/a_2665_112# 0.008469f
C12661 FILLER_0_4_144/a_572_375# net47 0.011686f
C12662 _132_ FILLER_0_18_107/a_2724_472# 0.002229f
C12663 net16 FILLER_0_18_37/a_1380_472# 0.002932f
C12664 _041_ net40 0.082688f
C12665 _219_/a_36_160# vdd 0.013125f
C12666 _098_ _433_/a_448_472# 0.027678f
C12667 _126_ vss 0.399848f
C12668 net62 _069_ 0.010033f
C12669 FILLER_0_3_2/a_124_375# vdd 0.021963f
C12670 net17 _450_/a_448_472# 0.017832f
C12671 _430_/a_1000_472# net21 0.053061f
C12672 _140_ _434_/a_448_472# 0.00128f
C12673 _027_ vdd 0.146607f
C12674 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2724_472# 0.026657f
C12675 _363_/a_36_68# _153_ 0.008003f
C12676 net36 FILLER_0_15_180/a_36_472# 0.007275f
C12677 net62 net29 0.082455f
C12678 result[2] vss 0.327009f
C12679 _159_ FILLER_0_2_127/a_124_375# 0.020951f
C12680 ctlp[1] _419_/a_2248_156# 0.028734f
C12681 _114_ _389_/a_36_148# 0.009465f
C12682 _037_ vdd 0.158731f
C12683 _255_/a_224_552# cal_itt\[3\] 0.003266f
C12684 _161_ _090_ 0.207838f
C12685 result[1] FILLER_0_11_282/a_36_472# 0.01775f
C12686 _056_ FILLER_0_12_196/a_36_472# 0.039555f
C12687 state\[1\] FILLER_0_13_142/a_1380_472# 0.006475f
C12688 _065_ trim_mask\[3\] 0.020092f
C12689 trim_val\[2\] _160_ 0.051804f
C12690 _448_/a_1000_472# net22 0.011389f
C12691 _323_/a_36_113# FILLER_0_10_247/a_36_472# 0.00136f
C12692 _434_/a_36_151# _146_ 0.003818f
C12693 _434_/a_1204_472# mask\[6\] 0.006692f
C12694 mask\[8\] _354_/a_49_472# 0.105272f
C12695 output22/a_224_472# mask\[7\] 0.05527f
C12696 FILLER_0_21_28/a_1468_375# _012_ 0.00351f
C12697 FILLER_0_0_96/a_36_472# trim_mask\[3\] 0.005343f
C12698 _443_/a_2665_112# FILLER_0_2_165/a_124_375# 0.006271f
C12699 _421_/a_2560_156# net19 0.006572f
C12700 FILLER_0_8_138/a_36_472# _120_ 0.006759f
C12701 net20 net81 0.036173f
C12702 FILLER_0_15_212/a_1380_472# vdd 0.003213f
C12703 FILLER_0_15_212/a_932_472# vss 0.019114f
C12704 FILLER_0_15_116/a_36_472# vdd 0.013454f
C12705 vdd FILLER_0_6_37/a_124_375# 0.041381f
C12706 net20 _426_/a_2665_112# 0.018602f
C12707 _236_/a_36_160# vdd 0.023428f
C12708 _411_/a_448_472# _073_ 0.004279f
C12709 FILLER_0_10_78/a_1380_472# _176_ 0.009351f
C12710 FILLER_0_5_164/a_484_472# net37 0.013857f
C12711 output34/a_224_472# net61 0.008309f
C12712 net2 _082_ 0.034094f
C12713 _091_ _055_ 0.003332f
C12714 net20 _060_ 0.0426f
C12715 FILLER_0_19_47/a_36_472# net26 0.050805f
C12716 _430_/a_36_151# _432_/a_2665_112# 0.030053f
C12717 _134_ FILLER_0_10_107/a_36_472# 0.006746f
C12718 net49 net40 0.093233f
C12719 output28/a_224_472# net18 0.015144f
C12720 _429_/a_2665_112# FILLER_0_14_235/a_36_472# 0.007491f
C12721 FILLER_0_17_38/a_36_472# _452_/a_36_151# 0.096503f
C12722 _140_ _022_ 0.001997f
C12723 _132_ mask\[9\] 0.203851f
C12724 net68 net40 0.036106f
C12725 _162_ _118_ 0.005444f
C12726 _120_ FILLER_0_9_72/a_484_472# 0.001645f
C12727 FILLER_0_10_107/a_124_375# vss 0.003015f
C12728 FILLER_0_10_107/a_572_375# vdd 0.043678f
C12729 _420_/a_2248_156# _009_ 0.00681f
C12730 _412_/a_448_472# _082_ 0.022743f
C12731 _445_/a_1204_472# net40 0.003916f
C12732 net52 net13 0.018118f
C12733 _086_ _255_/a_224_552# 0.073601f
C12734 input5/a_36_113# vdd 0.026855f
C12735 mask\[4\] FILLER_0_18_177/a_3260_375# 0.013881f
C12736 FILLER_0_18_177/a_3260_375# net22 0.049279f
C12737 _053_ net14 0.713784f
C12738 net18 net77 0.378783f
C12739 _412_/a_1000_472# vdd 0.002008f
C12740 _443_/a_1204_472# net23 0.026261f
C12741 _141_ _098_ 0.0697f
C12742 FILLER_0_20_177/a_1468_375# vdd 0.016422f
C12743 net50 _441_/a_2665_112# 0.056602f
C12744 net64 mask\[2\] 0.046428f
C12745 _440_/a_1308_423# net47 0.009738f
C12746 FILLER_0_12_124/a_124_375# _127_ 0.003767f
C12747 _301_/a_36_472# FILLER_0_22_86/a_36_472# 0.010679f
C12748 FILLER_0_4_49/a_36_472# net49 0.010951f
C12749 net38 _054_ 0.640545f
C12750 FILLER_0_13_212/a_1380_472# net79 0.006824f
C12751 ctln[3] FILLER_0_0_266/a_36_472# 0.012298f
C12752 output46/a_224_472# FILLER_0_20_15/a_124_375# 0.029497f
C12753 mask\[2\] mask\[1\] 0.059794f
C12754 ctln[6] _170_ 0.005146f
C12755 calibrate FILLER_0_9_270/a_124_375# 0.002292f
C12756 _154_ _160_ 0.395185f
C12757 output42/a_224_472# net67 0.05585f
C12758 FILLER_0_11_142/a_36_472# FILLER_0_13_142/a_124_375# 0.0027f
C12759 _069_ _429_/a_448_472# 0.035108f
C12760 _411_/a_1204_472# _000_ 0.002575f
C12761 FILLER_0_4_49/a_36_472# net68 0.00894f
C12762 net78 _420_/a_448_472# 0.001091f
C12763 net82 _443_/a_1308_423# 0.006706f
C12764 net50 _439_/a_2248_156# 0.007461f
C12765 _321_/a_170_472# _176_ 0.059301f
C12766 _449_/a_36_151# net74 0.032989f
C12767 _073_ FILLER_0_6_231/a_36_472# 0.001898f
C12768 FILLER_0_17_104/a_1380_472# vdd 0.010877f
C12769 _095_ FILLER_0_14_107/a_1020_375# 0.014156f
C12770 _050_ FILLER_0_22_107/a_36_472# 0.001098f
C12771 _425_/a_2665_112# net37 0.008519f
C12772 ctln[5] _448_/a_36_151# 0.009209f
C12773 result[7] ctlp[1] 0.07619f
C12774 _131_ _332_/a_36_472# 0.006825f
C12775 _010_ _420_/a_2560_156# 0.070902f
C12776 _136_ _451_/a_1353_112# 0.058703f
C12777 _069_ net23 0.418375f
C12778 _365_/a_36_68# _156_ 0.027744f
C12779 fanout73/a_36_113# _095_ 0.003989f
C12780 net20 _079_ 0.177911f
C12781 _137_ vss 0.343959f
C12782 FILLER_0_18_171/a_124_375# vss 0.048769f
C12783 _422_/a_796_472# _009_ 0.001178f
C12784 ctlp[1] FILLER_0_23_282/a_484_472# 0.007608f
C12785 net49 FILLER_0_3_78/a_484_472# 0.048729f
C12786 _453_/a_448_472# vdd 0.010005f
C12787 _453_/a_36_151# vss 0.007105f
C12788 _031_ FILLER_0_2_111/a_1380_472# 0.01562f
C12789 FILLER_0_16_57/a_124_375# net15 0.001594f
C12790 net48 _068_ 0.054333f
C12791 mask\[4\] _201_/a_67_603# 0.029139f
C12792 net22 _201_/a_67_603# 0.004491f
C12793 net63 _091_ 0.767908f
C12794 net25 _423_/a_2248_156# 0.005535f
C12795 _429_/a_36_151# FILLER_0_15_212/a_484_472# 0.001723f
C12796 net74 FILLER_0_13_100/a_36_472# 0.003924f
C12797 net36 FILLER_0_18_76/a_36_472# 0.001728f
C12798 net13 _387_/a_36_113# 0.00189f
C12799 _076_ FILLER_0_3_221/a_484_472# 0.001225f
C12800 net67 net51 0.010753f
C12801 en_co_clk _172_ 0.025699f
C12802 FILLER_0_19_171/a_484_472# vdd 0.009225f
C12803 FILLER_0_19_171/a_36_472# vss 0.001338f
C12804 FILLER_0_20_15/a_932_472# net40 0.002705f
C12805 mask\[3\] _094_ 0.00554f
C12806 _142_ _341_/a_49_472# 0.011026f
C12807 _091_ FILLER_0_13_212/a_1468_375# 0.003576f
C12808 _161_ _076_ 0.042123f
C12809 net69 vss 0.34555f
C12810 net82 FILLER_0_2_177/a_36_472# 0.001777f
C12811 _432_/a_1308_423# FILLER_0_18_177/a_36_472# 0.009119f
C12812 fanout77/a_36_113# net78 0.019286f
C12813 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_484_472# 0.026657f
C12814 _144_ _433_/a_2560_156# 0.01064f
C12815 output36/a_224_472# _196_/a_36_160# 0.001309f
C12816 FILLER_0_4_177/a_36_472# _386_/a_848_380# 0.007646f
C12817 _415_/a_796_472# net81 0.002008f
C12818 output13/a_224_472# vdd 0.045929f
C12819 _057_ _072_ 0.048392f
C12820 calibrate net18 0.014127f
C12821 _096_ _113_ 0.650985f
C12822 cal_count\[1\] FILLER_0_15_59/a_36_472# 0.00544f
C12823 _180_ FILLER_0_15_59/a_124_375# 0.009926f
C12824 output16/a_224_472# net16 0.054603f
C12825 FILLER_0_18_177/a_3172_472# FILLER_0_18_209/a_36_472# 0.013276f
C12826 net16 _450_/a_2225_156# 0.001015f
C12827 output7/a_224_472# ctln[9] 0.001987f
C12828 FILLER_0_5_128/a_36_472# _163_ 0.009857f
C12829 FILLER_0_10_37/a_124_375# net51 0.006198f
C12830 _322_/a_124_24# vdd 0.01572f
C12831 _450_/a_448_472# _039_ 0.047559f
C12832 _008_ ctlp[1] 0.002566f
C12833 _008_ _419_/a_796_472# 0.013039f
C12834 net53 FILLER_0_14_107/a_1380_472# 0.059367f
C12835 _302_/a_224_472# _012_ 0.002675f
C12836 fanout63/a_36_160# _098_ 0.003627f
C12837 _086_ FILLER_0_5_172/a_124_375# 0.007355f
C12838 FILLER_0_17_226/a_124_375# fanout63/a_36_160# 0.008215f
C12839 _067_ FILLER_0_12_20/a_484_472# 0.011046f
C12840 _449_/a_36_151# FILLER_0_13_72/a_124_375# 0.059049f
C12841 output12/a_224_472# FILLER_0_1_192/a_124_375# 0.032639f
C12842 _196_/a_36_160# vdd 0.106963f
C12843 _086_ _128_ 0.085571f
C12844 _115_ _308_/a_124_24# 0.039354f
C12845 output44/a_224_472# FILLER_0_18_2/a_1916_375# 0.032639f
C12846 mask\[4\] FILLER_0_19_187/a_36_472# 0.004669f
C12847 _420_/a_2560_156# vdd 0.001652f
C12848 _420_/a_2665_112# vss 0.001749f
C12849 _432_/a_448_472# FILLER_0_19_171/a_572_375# 0.00184f
C12850 result[9] _421_/a_1204_472# 0.014964f
C12851 ctlp[7] net54 0.004355f
C12852 net61 FILLER_0_21_286/a_484_472# 0.001829f
C12853 _147_ _434_/a_36_151# 0.001817f
C12854 net53 _451_/a_1040_527# 0.023651f
C12855 net57 _374_/a_36_68# 0.001052f
C12856 valid fanout59/a_36_160# 0.029107f
C12857 _411_/a_36_151# net20 0.011179f
C12858 _308_/a_1084_68# trim_mask\[0\] 0.001592f
C12859 _028_ net14 0.066292f
C12860 _077_ net21 0.032627f
C12861 net19 _419_/a_2665_112# 0.00276f
C12862 FILLER_0_17_104/a_572_375# net14 0.004285f
C12863 _069_ _056_ 0.035189f
C12864 net69 _369_/a_244_472# 0.002456f
C12865 _086_ FILLER_0_11_142/a_572_375# 0.011726f
C12866 FILLER_0_10_214/a_36_472# _090_ 0.011963f
C12867 FILLER_0_18_209/a_484_472# _047_ 0.002188f
C12868 net81 cal_itt\[1\] 0.387207f
C12869 FILLER_0_22_86/a_484_472# FILLER_0_23_88/a_124_375# 0.001684f
C12870 result[9] FILLER_0_15_282/a_124_375# 0.001233f
C12871 FILLER_0_3_172/a_932_472# net22 0.012284f
C12872 FILLER_0_9_28/a_1828_472# _042_ 0.001809f
C12873 _434_/a_2665_112# vdd 0.030225f
C12874 _075_ _122_ 0.030339f
C12875 FILLER_0_13_142/a_1380_472# vdd 0.001977f
C12876 FILLER_0_13_142/a_932_472# vss 0.005192f
C12877 FILLER_0_4_177/a_484_472# vss 0.002399f
C12878 net20 result[8] 0.014571f
C12879 net56 vss 0.367812f
C12880 result[7] FILLER_0_23_282/a_124_375# 0.016009f
C12881 _417_/a_796_472# vss 0.001608f
C12882 net62 _417_/a_448_472# 0.011318f
C12883 _074_ FILLER_0_6_177/a_124_375# 0.003608f
C12884 net67 net6 0.345681f
C12885 _424_/a_1308_423# _012_ 0.007041f
C12886 _415_/a_448_472# FILLER_0_9_270/a_36_472# 0.012285f
C12887 _077_ _070_ 0.29321f
C12888 net41 FILLER_0_19_28/a_572_375# 0.040551f
C12889 _126_ _332_/a_36_472# 0.009299f
C12890 _213_/a_67_603# vss 0.019344f
C12891 FILLER_0_5_109/a_36_472# _155_ 0.001872f
C12892 _127_ _076_ 0.137964f
C12893 _091_ _432_/a_36_151# 0.054497f
C12894 _177_ _451_/a_2449_156# 0.002085f
C12895 FILLER_0_16_73/a_484_472# net15 0.001946f
C12896 net35 FILLER_0_22_177/a_572_375# 0.007797f
C12897 _248_/a_36_68# vss 0.027935f
C12898 net54 net36 0.005827f
C12899 FILLER_0_10_214/a_36_472# net22 0.001634f
C12900 cal_count\[3\] _408_/a_1936_472# 0.007046f
C12901 FILLER_0_3_172/a_572_375# vdd 0.007121f
C12902 _422_/a_1204_472# vdd 0.001062f
C12903 cal_count\[2\] _182_ 0.044348f
C12904 net20 net64 0.374636f
C12905 _069_ FILLER_0_13_212/a_36_472# 0.047013f
C12906 net81 vss 0.766885f
C12907 _165_ vss 0.048027f
C12908 _399_/a_224_472# net16 0.003817f
C12909 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001597f
C12910 _426_/a_2665_112# vss 0.006288f
C12911 FILLER_0_11_64/a_124_375# _453_/a_36_151# 0.005577f
C12912 FILLER_0_12_136/a_1380_472# _076_ 0.001809f
C12913 FILLER_0_19_125/a_124_375# _132_ 0.009167f
C12914 net38 _035_ 0.02987f
C12915 net20 mask\[1\] 0.09671f
C12916 _088_ FILLER_0_3_172/a_3260_375# 0.002239f
C12917 net62 FILLER_0_15_282/a_36_472# 0.013655f
C12918 trim_mask\[0\] net14 0.499565f
C12919 result[6] net62 0.005382f
C12920 _104_ _199_/a_36_160# 0.095519f
C12921 ctlp[1] FILLER_0_24_290/a_36_472# 0.037615f
C12922 _060_ vss 0.318005f
C12923 net41 net46 0.061224f
C12924 net66 _030_ 0.087608f
C12925 _098_ FILLER_0_15_212/a_572_375# 0.009099f
C12926 FILLER_0_1_192/a_36_472# net21 0.016033f
C12927 FILLER_0_17_142/a_124_375# FILLER_0_17_133/a_124_375# 0.003228f
C12928 net69 _441_/a_1204_472# 0.014374f
C12929 trim_mask\[2\] net69 0.051795f
C12930 fanout61/a_36_113# net62 0.031315f
C12931 _093_ FILLER_0_16_89/a_1020_375# 0.004133f
C12932 FILLER_0_21_125/a_36_472# _140_ 0.101284f
C12933 FILLER_0_3_172/a_124_375# FILLER_0_2_171/a_124_375# 0.026339f
C12934 _089_ FILLER_0_3_172/a_2276_472# 0.001522f
C12935 FILLER_0_16_37/a_36_472# _402_/a_728_93# 0.0108f
C12936 _321_/a_358_69# _121_ 0.00135f
C12937 net71 _437_/a_2248_156# 0.025557f
C12938 ctln[4] FILLER_0_0_198/a_36_472# 0.02582f
C12939 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_124_375# 0.026339f
C12940 _445_/a_448_472# net49 0.00122f
C12941 net63 FILLER_0_15_212/a_484_472# 0.059367f
C12942 FILLER_0_4_152/a_36_472# net57 0.015332f
C12943 output11/a_224_472# net11 0.003448f
C12944 _122_ FILLER_0_5_164/a_484_472# 0.002997f
C12945 _267_/a_36_472# _055_ 0.035376f
C12946 _128_ FILLER_0_9_142/a_124_375# 0.004439f
C12947 fanout80/a_36_113# net36 0.007625f
C12948 _003_ net37 0.046745f
C12949 mask\[9\] FILLER_0_19_111/a_124_375# 0.031474f
C12950 _326_/a_36_160# _077_ 0.00419f
C12951 _253_/a_244_68# _073_ 0.002878f
C12952 net52 FILLER_0_5_72/a_572_375# 0.024148f
C12953 _246_/a_36_68# _090_ 0.001712f
C12954 net12 vss 0.043754f
C12955 _341_/a_49_472# mask\[2\] 0.026222f
C12956 ctln[1] output11/a_224_472# 0.004299f
C12957 _059_ FILLER_0_8_156/a_124_375# 0.00593f
C12958 fanout73/a_36_113# net74 0.04136f
C12959 net37 net21 0.03272f
C12960 _072_ cal_count\[3\] 0.028346f
C12961 _184_ net40 0.122833f
C12962 _079_ cal_itt\[1\] 0.012324f
C12963 net57 FILLER_0_3_142/a_124_375# 0.003738f
C12964 _124_ _134_ 0.002508f
C12965 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_124_375# 0.007947f
C12966 FILLER_0_2_111/a_1020_375# vdd 0.007918f
C12967 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3260_375# 0.086635f
C12968 _372_/a_786_69# _163_ 0.001179f
C12969 FILLER_0_18_2/a_2812_375# FILLER_0_20_15/a_1380_472# 0.001338f
C12970 _360_/a_36_160# FILLER_0_4_123/a_36_472# 0.001165f
C12971 fanout70/a_36_113# vdd 0.015969f
C12972 _428_/a_1308_423# _131_ 0.037599f
C12973 _154_ _156_ 0.019471f
C12974 _255_/a_224_552# _161_ 0.025424f
C12975 FILLER_0_7_72/a_36_472# vss 0.033878f
C12976 net26 FILLER_0_21_28/a_2276_472# 0.001561f
C12977 FILLER_0_18_107/a_2724_472# vdd 0.004677f
C12978 _103_ _419_/a_448_472# 0.001207f
C12979 _418_/a_2665_112# _417_/a_2665_112# 0.00131f
C12980 _070_ net37 0.036662f
C12981 _052_ vdd 0.264744f
C12982 net78 _419_/a_1308_423# 0.018598f
C12983 _016_ FILLER_0_12_136/a_1020_375# 0.001659f
C12984 net63 FILLER_0_20_177/a_572_375# 0.00281f
C12985 _149_ _437_/a_1204_472# 0.024276f
C12986 _026_ _437_/a_796_472# 0.008884f
C12987 cal_count\[3\] net47 0.043032f
C12988 net28 _426_/a_448_472# 0.00154f
C12989 net41 FILLER_0_18_2/a_3260_375# 0.042057f
C12990 net34 _435_/a_1308_423# 0.008652f
C12991 _088_ vdd 0.140259f
C12992 _079_ vss 0.124667f
C12993 _093_ FILLER_0_17_72/a_572_375# 0.005609f
C12994 _126_ net79 0.085443f
C12995 mask\[0\] FILLER_0_13_206/a_124_375# 0.005989f
C12996 FILLER_0_10_78/a_124_375# FILLER_0_11_78/a_124_375# 0.05841f
C12997 trim[4] net39 0.004535f
C12998 FILLER_0_13_142/a_36_472# net23 0.003007f
C12999 _425_/a_2560_156# calibrate 0.010842f
C13000 mask\[4\] FILLER_0_19_155/a_124_375# 0.043876f
C13001 net68 _120_ 0.001304f
C13002 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_124_375# 0.012001f
C13003 result[2] net79 0.077934f
C13004 _077_ FILLER_0_12_50/a_36_472# 0.177624f
C13005 output12/a_224_472# FILLER_0_0_198/a_124_375# 0.00515f
C13006 net52 _160_ 0.133292f
C13007 _103_ mask\[2\] 0.002168f
C13008 _053_ _372_/a_170_472# 0.05895f
C13009 _053_ _131_ 0.086215f
C13010 FILLER_0_16_107/a_572_375# _093_ 0.002827f
C13011 FILLER_0_21_125/a_36_472# _149_ 0.008849f
C13012 _057_ state\[1\] 0.284428f
C13013 _449_/a_2248_156# fanout55/a_36_160# 0.027388f
C13014 net7 _064_ 0.001538f
C13015 _142_ FILLER_0_17_142/a_572_375# 0.012321f
C13016 _095_ vss 1.465527f
C13017 _413_/a_36_151# FILLER_0_3_172/a_3172_472# 0.001723f
C13018 FILLER_0_11_101/a_124_375# net14 0.011983f
C13019 FILLER_0_18_107/a_2812_375# _145_ 0.030158f
C13020 FILLER_0_17_38/a_484_472# _182_ 0.00527f
C13021 net47 net40 0.635497f
C13022 FILLER_0_4_144/a_124_375# vss 0.017638f
C13023 FILLER_0_4_144/a_572_375# vdd -0.013698f
C13024 net57 fanout52/a_36_160# 0.122432f
C13025 net47 _169_ 0.528536f
C13026 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_124_375# 0.003732f
C13027 FILLER_0_16_73/a_36_472# vss 0.035175f
C13028 result[9] _419_/a_1000_472# 0.012469f
C13029 _397_/a_36_472# _131_ 0.012338f
C13030 net27 FILLER_0_11_282/a_36_472# 0.001526f
C13031 net63 FILLER_0_19_171/a_1468_375# 0.006671f
C13032 _093_ net70 0.001888f
C13033 _430_/a_1308_423# _069_ 0.024499f
C13034 net7 output41/a_224_472# 0.019483f
C13035 _132_ cal_count\[3\] 0.193553f
C13036 net54 FILLER_0_22_107/a_484_472# 0.005897f
C13037 _104_ _294_/a_224_472# 0.003008f
C13038 result[6] FILLER_0_23_290/a_124_375# 0.001492f
C13039 _449_/a_2665_112# vss 0.007395f
C13040 net72 _052_ 0.138281f
C13041 net55 _217_/a_36_160# 0.001311f
C13042 fanout81/a_36_160# net82 0.027351f
C13043 FILLER_0_9_28/a_1468_375# _444_/a_2248_156# 0.001074f
C13044 mask\[9\] vdd 0.940144f
C13045 _429_/a_448_472# net22 0.054866f
C13046 cal_itt\[2\] _253_/a_244_68# 0.001073f
C13047 net10 net8 0.003331f
C13048 _337_/a_257_69# _137_ 0.001822f
C13049 net17 _452_/a_36_151# 0.041497f
C13050 _431_/a_2560_156# FILLER_0_17_142/a_124_375# 0.001178f
C13051 _450_/a_448_472# clkc 0.003011f
C13052 _450_/a_1040_527# net6 0.019715f
C13053 FILLER_0_19_47/a_572_375# FILLER_0_18_53/a_36_472# 0.001684f
C13054 net27 FILLER_0_14_235/a_36_472# 0.003401f
C13055 FILLER_0_17_72/a_484_472# vss 0.005334f
C13056 FILLER_0_4_49/a_36_472# net47 0.002964f
C13057 FILLER_0_14_181/a_36_472# _098_ 0.004669f
C13058 _425_/a_36_151# FILLER_0_8_247/a_572_375# 0.001597f
C13059 FILLER_0_12_136/a_572_375# _427_/a_1308_423# 0.001238f
C13060 vdd rstn 0.160093f
C13061 _068_ FILLER_0_5_148/a_124_375# 0.003986f
C13062 _430_/a_36_151# _139_ 0.012035f
C13063 net18 FILLER_0_9_270/a_572_375# 0.005977f
C13064 FILLER_0_8_247/a_1380_472# calibrate 0.008605f
C13065 output38/a_224_472# output39/a_224_472# 0.002978f
C13066 FILLER_0_7_72/a_1020_375# net52 0.00799f
C13067 _178_ net3 0.257606f
C13068 mask\[4\] net23 0.111873f
C13069 net35 _051_ 0.019252f
C13070 net60 _421_/a_796_472# 0.002046f
C13071 FILLER_0_22_86/a_1380_472# vdd 0.008224f
C13072 FILLER_0_22_86/a_932_472# vss -0.001553f
C13073 _422_/a_1000_472# mask\[7\] 0.039617f
C13074 _418_/a_796_472# vss 0.00145f
C13075 net15 _423_/a_36_151# 0.003422f
C13076 net52 _443_/a_2248_156# 0.045316f
C13077 _411_/a_36_151# vss 0.035447f
C13078 net57 _428_/a_448_472# 0.032029f
C13079 _091_ FILLER_0_15_212/a_1020_375# 0.00799f
C13080 net55 _038_ 0.05656f
C13081 en_co_clk _136_ 0.034892f
C13082 net61 _422_/a_36_151# 0.003736f
C13083 cal_count\[2\] FILLER_0_15_2/a_36_472# 0.037661f
C13084 _426_/a_1000_472# calibrate 0.002865f
C13085 net4 _248_/a_36_68# 0.054512f
C13086 FILLER_0_18_107/a_36_472# net14 0.005297f
C13087 _065_ _168_ 0.020406f
C13088 _162_ FILLER_0_5_172/a_36_472# 0.001501f
C13089 net20 _260_/a_244_472# 0.001593f
C13090 _379_/a_36_472# net47 0.016584f
C13091 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_124_375# 0.012267f
C13092 _055_ _113_ 0.153988f
C13093 _128_ _161_ 0.027657f
C13094 net81 net4 0.003327f
C13095 FILLER_0_16_241/a_36_472# FILLER_0_15_235/a_572_375# 0.001543f
C13096 FILLER_0_9_28/a_2812_375# _077_ 0.006629f
C13097 _104_ net33 0.037008f
C13098 net2 net19 0.031976f
C13099 _453_/a_2248_156# net51 0.05329f
C13100 FILLER_0_24_63/a_124_375# ctlp[9] 0.002726f
C13101 result[8] vss 0.235206f
C13102 _426_/a_2665_112# net4 0.011288f
C13103 _402_/a_2172_497# cal_count\[1\] 0.008211f
C13104 _421_/a_2665_112# net33 0.007127f
C13105 _028_ FILLER_0_5_72/a_1020_375# 0.00123f
C13106 mask\[6\] _146_ 0.181681f
C13107 FILLER_0_12_2/a_572_375# _039_ 0.005407f
C13108 net17 FILLER_0_12_28/a_124_375# 0.009108f
C13109 _093_ _132_ 0.105039f
C13110 FILLER_0_4_107/a_484_472# net47 0.001975f
C13111 _308_/a_848_380# FILLER_0_10_94/a_484_472# 0.019491f
C13112 _086_ _395_/a_1492_488# 0.001769f
C13113 FILLER_0_12_20/a_124_375# net47 0.047331f
C13114 _052_ _424_/a_36_151# 0.010844f
C13115 net4 _060_ 0.327437f
C13116 output34/a_224_472# _293_/a_36_472# 0.001888f
C13117 _098_ _434_/a_448_472# 0.015893f
C13118 net57 _443_/a_448_472# 0.001956f
C13119 net27 FILLER_0_8_263/a_124_375# 0.016669f
C13120 FILLER_0_17_200/a_484_472# _430_/a_36_151# 0.001723f
C13121 sample net64 0.209777f
C13122 _412_/a_448_472# net19 0.001526f
C13123 mask\[3\] FILLER_0_18_177/a_124_375# 0.002924f
C13124 _235_/a_67_603# net17 0.018056f
C13125 FILLER_0_8_239/a_124_375# _123_ 0.001286f
C13126 result[6] net33 0.363421f
C13127 _187_ _408_/a_728_93# 0.002598f
C13128 input2/a_36_113# net2 0.015844f
C13129 FILLER_0_16_255/a_124_375# vdd 0.029925f
C13130 net64 vss 0.636644f
C13131 _440_/a_1308_423# vdd 0.00218f
C13132 _440_/a_448_472# vss 0.032037f
C13133 _446_/a_2248_156# net49 0.006196f
C13134 trim_mask\[1\] _164_ 0.195956f
C13135 mask\[1\] vss 0.46268f
C13136 fanout49/a_36_160# _441_/a_2248_156# 0.027388f
C13137 net52 _170_ 0.378738f
C13138 _141_ _137_ 0.40175f
C13139 _118_ _055_ 0.042556f
C13140 _056_ _090_ 0.177189f
C13141 net1 _265_/a_224_472# 0.005504f
C13142 _019_ mask\[2\] 0.155325f
C13143 _131_ FILLER_0_17_104/a_572_375# 0.003214f
C13144 net76 FILLER_0_3_172/a_1468_375# 0.039469f
C13145 net36 _195_/a_67_603# 0.034361f
C13146 FILLER_0_10_78/a_36_472# _439_/a_36_151# 0.00271f
C13147 _141_ FILLER_0_19_171/a_36_472# 0.001292f
C13148 mask\[5\] FILLER_0_20_169/a_36_472# 0.016469f
C13149 FILLER_0_5_72/a_1380_472# trim_mask\[1\] 0.01221f
C13150 net65 _448_/a_448_472# 0.001006f
C13151 _352_/a_49_472# vdd 0.077542f
C13152 FILLER_0_6_47/a_36_472# vss 0.002433f
C13153 FILLER_0_6_47/a_484_472# vdd 0.005065f
C13154 _176_ _129_ 0.036112f
C13155 output39/a_224_472# vdd 0.022593f
C13156 net33 net22 0.066751f
C13157 _059_ _163_ 0.038651f
C13158 ctln[9] vss 0.167242f
C13159 net20 FILLER_0_12_236/a_36_472# 0.003143f
C13160 FILLER_0_12_20/a_484_472# _450_/a_448_472# 0.04564f
C13161 net39 net17 0.099429f
C13162 output18/a_224_472# output19/a_224_472# 0.00124f
C13163 mask\[8\] vss 0.378558f
C13164 net35 vdd 1.0365f
C13165 _425_/a_36_151# _317_/a_36_113# 0.002361f
C13166 FILLER_0_6_239/a_124_375# vdd 0.031271f
C13167 _076_ net23 0.105196f
C13168 valid net37 0.051518f
C13169 cal_count\[3\] state\[1\] 0.236393f
C13170 _098_ _022_ 0.013131f
C13171 FILLER_0_2_111/a_124_375# _154_ 0.004032f
C13172 net65 FILLER_0_3_221/a_1020_375# 0.001641f
C13173 net17 _039_ 0.079171f
C13174 _056_ net22 0.075673f
C13175 _014_ _122_ 0.001529f
C13176 fanout68/a_36_113# vdd 0.012621f
C13177 _422_/a_2665_112# _108_ 0.023365f
C13178 _418_/a_36_151# net77 0.019316f
C13179 net67 _067_ 0.151887f
C13180 FILLER_0_5_109/a_484_472# FILLER_0_5_117/a_36_472# 0.013276f
C13181 _140_ _023_ 0.079452f
C13182 net20 _103_ 0.261438f
C13183 FILLER_0_16_57/a_1468_375# _111_ 0.001371f
C13184 _098_ FILLER_0_16_154/a_1380_472# 0.00417f
C13185 _118_ _313_/a_67_603# 0.001793f
C13186 _328_/a_36_113# vss 0.044028f
C13187 _079_ net4 0.023763f
C13188 _081_ FILLER_0_5_136/a_124_375# 0.025819f
C13189 net16 _233_/a_36_160# 0.01152f
C13190 FILLER_0_14_81/a_124_375# vss 0.03341f
C13191 FILLER_0_14_81/a_36_472# vdd 0.00958f
C13192 _114_ FILLER_0_10_107/a_36_472# 0.00263f
C13193 output29/a_224_472# result[2] 0.058798f
C13194 _003_ _122_ 0.033778f
C13195 FILLER_0_22_86/a_572_375# net14 0.009573f
C13196 _091_ FILLER_0_19_171/a_124_375# 0.028992f
C13197 net78 net19 0.507249f
C13198 net41 _446_/a_2560_156# 0.005695f
C13199 ctln[7] ctln[8] 0.004643f
C13200 _448_/a_448_472# net59 0.050956f
C13201 trim[4] net42 0.016428f
C13202 trim_val\[4\] net22 0.144267f
C13203 _127_ _128_ 0.257374f
C13204 _122_ net21 0.026632f
C13205 _387_/a_36_113# _170_ 0.017801f
C13206 _086_ _311_/a_2700_473# 0.00176f
C13207 FILLER_0_18_171/a_36_472# _091_ 0.00395f
C13208 FILLER_0_0_96/a_124_375# vdd 0.034959f
C13209 trimb[4] vss 0.039934f
C13210 FILLER_0_13_212/a_36_472# net22 0.002402f
C13211 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_124_375# 0.012001f
C13212 _062_ FILLER_0_8_156/a_484_472# 0.006123f
C13213 net74 vss 0.589483f
C13214 _321_/a_170_472# FILLER_0_11_135/a_124_375# 0.001153f
C13215 output37/a_224_472# net76 0.004028f
C13216 net53 net14 0.04525f
C13217 _068_ _055_ 0.443477f
C13218 FILLER_0_9_223/a_124_375# vdd 0.006153f
C13219 net55 FILLER_0_11_78/a_484_472# 0.038269f
C13220 _242_/a_36_160# FILLER_0_5_164/a_124_375# 0.005705f
C13221 result[5] net19 0.003542f
C13222 net15 FILLER_0_17_56/a_124_375# 0.001854f
C13223 _133_ calibrate 0.0188f
C13224 _070_ _122_ 0.153373f
C13225 _002_ FILLER_0_3_172/a_1916_375# 0.047331f
C13226 _437_/a_1204_472# net14 0.004949f
C13227 net79 _417_/a_796_472# 0.001042f
C13228 net68 _220_/a_255_603# 0.001908f
C13229 _057_ vdd 0.801978f
C13230 net16 net55 0.035875f
C13231 net75 FILLER_0_6_239/a_124_375# 0.013962f
C13232 FILLER_0_7_104/a_36_472# FILLER_0_9_105/a_124_375# 0.001188f
C13233 net41 cal_count\[2\] 0.079279f
C13234 FILLER_0_17_38/a_572_375# _041_ 0.021754f
C13235 cal_count\[1\] vss 0.307993f
C13236 FILLER_0_4_123/a_36_472# _159_ 0.004956f
C13237 _092_ _093_ 0.287983f
C13238 trim[4] clkc 0.005f
C13239 FILLER_0_12_136/a_1380_472# FILLER_0_11_142/a_572_375# 0.001543f
C13240 _114_ FILLER_0_10_94/a_124_375# 0.040691f
C13241 _141_ net56 0.012364f
C13242 _033_ _444_/a_36_151# 0.014843f
C13243 FILLER_0_12_136/a_36_472# cal_count\[3\] 0.006102f
C13244 _061_ net21 0.049282f
C13245 FILLER_0_19_125/a_124_375# vdd 0.032954f
C13246 _068_ _311_/a_1212_473# 0.002835f
C13247 net79 _248_/a_36_68# 0.018243f
C13248 _427_/a_2248_156# _095_ 0.022479f
C13249 net68 FILLER_0_5_54/a_932_472# 0.013043f
C13250 _058_ _118_ 0.001451f
C13251 _068_ _313_/a_67_603# 0.012208f
C13252 FILLER_0_18_2/a_2364_375# net38 0.001683f
C13253 result[4] net30 0.298966f
C13254 net81 net79 0.178225f
C13255 _451_/a_3129_107# vdd 0.008569f
C13256 net65 FILLER_0_1_266/a_36_472# 0.003529f
C13257 FILLER_0_9_28/a_36_472# net47 0.006712f
C13258 _445_/a_448_472# net47 0.005429f
C13259 _118_ _315_/a_36_68# 0.005792f
C13260 FILLER_0_14_123/a_36_472# _043_ 0.001782f
C13261 _420_/a_36_151# FILLER_0_23_274/a_124_375# 0.059049f
C13262 net61 _419_/a_1000_472# 0.017712f
C13263 net60 _419_/a_1308_423# 0.029697f
C13264 _216_/a_67_603# _012_ 0.001014f
C13265 net57 _176_ 0.192223f
C13266 FILLER_0_16_89/a_1380_472# _040_ 0.008446f
C13267 net50 trim_val\[3\] 0.111824f
C13268 net82 FILLER_0_4_213/a_36_472# 0.003042f
C13269 _056_ _076_ 0.938912f
C13270 _061_ _070_ 0.02813f
C13271 net79 _060_ 0.019511f
C13272 _443_/a_1308_423# net69 0.004128f
C13273 _443_/a_36_151# _031_ 0.014344f
C13274 _032_ _442_/a_36_151# 0.005632f
C13275 net57 _306_/a_36_68# 0.042596f
C13276 FILLER_0_18_2/a_3172_472# _041_ 0.001503f
C13277 FILLER_0_9_28/a_572_375# net50 0.002807f
C13278 result[8] mask\[7\] 0.110637f
C13279 net78 _009_ 0.02395f
C13280 _008_ _199_/a_36_160# 0.002015f
C13281 net2 fanout58/a_36_160# 0.010424f
C13282 net27 FILLER_0_9_282/a_484_472# 0.006955f
C13283 FILLER_0_18_177/a_1828_472# vss -0.001107f
C13284 FILLER_0_18_177/a_2276_472# vdd 0.005211f
C13285 trimb[3] net17 0.005798f
C13286 _147_ mask\[6\] 0.103475f
C13287 FILLER_0_12_28/a_124_375# _039_ 0.004669f
C13288 _132_ FILLER_0_19_125/a_36_472# 0.008568f
C13289 _104_ _046_ 0.035267f
C13290 FILLER_0_9_28/a_1828_472# _120_ 0.00108f
C13291 _044_ FILLER_0_13_290/a_124_375# 0.001855f
C13292 net35 FILLER_0_22_128/a_572_375# 0.010439f
C13293 _411_/a_1308_423# ctln[1] 0.037098f
C13294 trimb[2] vdd 0.084666f
C13295 net35 _024_ 0.001335f
C13296 _079_ FILLER_0_5_198/a_124_375# 0.013896f
C13297 mask\[5\] FILLER_0_20_193/a_484_472# 0.02147f
C13298 net31 net19 0.023019f
C13299 _128_ FILLER_0_10_214/a_36_472# 0.00186f
C13300 vdd FILLER_0_13_72/a_572_375# -0.001166f
C13301 vss FILLER_0_13_72/a_124_375# 0.043492f
C13302 _042_ vdd 0.261947f
C13303 _398_/a_36_113# cal_count\[2\] 0.004895f
C13304 _178_ _405_/a_67_603# 0.02427f
C13305 output16/a_224_472# _447_/a_2665_112# 0.005471f
C13306 net16 _447_/a_1000_472# 0.003207f
C13307 FILLER_0_16_57/a_484_472# vdd 0.005894f
C13308 FILLER_0_16_57/a_36_472# vss 0.003789f
C13309 net15 _174_ 0.090215f
C13310 _106_ _105_ 0.038327f
C13311 fanout78/a_36_113# net78 0.004202f
C13312 output15/a_224_472# _383_/a_36_472# 0.001154f
C13313 _260_/a_36_68# vdd 0.011119f
C13314 FILLER_0_8_138/a_36_472# _062_ 0.001109f
C13315 cal fanout58/a_36_160# 0.047586f
C13316 net4 net64 0.060449f
C13317 FILLER_0_22_86/a_572_375# _098_ 0.001139f
C13318 result[7] FILLER_0_23_290/a_124_375# 0.018455f
C13319 FILLER_0_16_107/a_484_472# net70 0.002732f
C13320 ctlp[1] _098_ 0.0012f
C13321 net54 _437_/a_448_472# 0.004418f
C13322 _133_ _125_ 0.014858f
C13323 _068_ _058_ 0.092852f
C13324 _444_/a_2665_112# trim_val\[0\] 0.007249f
C13325 FILLER_0_2_93/a_572_375# net14 0.044606f
C13326 net15 FILLER_0_5_72/a_124_375# 0.006403f
C13327 _155_ _363_/a_36_68# 0.013915f
C13328 FILLER_0_5_72/a_1380_472# _164_ 0.049427f
C13329 ctlp[0] net17 0.006778f
C13330 net66 _382_/a_224_472# 0.001902f
C13331 _065_ _447_/a_36_151# 0.043351f
C13332 _068_ _315_/a_36_68# 0.003516f
C13333 _093_ FILLER_0_19_111/a_124_375# 0.00186f
C13334 FILLER_0_12_2/a_484_472# net6 0.005586f
C13335 FILLER_0_24_63/a_36_472# _423_/a_2665_112# 0.001873f
C13336 _101_ _094_ 0.304499f
C13337 mask\[0\] FILLER_0_14_235/a_484_472# 0.004688f
C13338 _083_ _001_ 0.002625f
C13339 output38/a_224_472# net40 0.072234f
C13340 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_572_375# 0.086635f
C13341 FILLER_0_18_177/a_1916_375# FILLER_0_19_195/a_36_472# 0.001684f
C13342 output27/a_224_472# FILLER_0_9_270/a_124_375# 0.001274f
C13343 mask\[8\] mask\[7\] 0.021731f
C13344 result[5] fanout78/a_36_113# 0.018989f
C13345 _126_ FILLER_0_14_181/a_36_472# 0.008653f
C13346 _446_/a_36_151# _035_ 0.012914f
C13347 _016_ _427_/a_796_472# 0.001666f
C13348 _341_/a_49_472# vss 0.003485f
C13349 FILLER_0_21_28/a_572_375# net40 0.001406f
C13350 _430_/a_1308_423# net22 0.035518f
C13351 mask\[8\] _148_ 0.356546f
C13352 _015_ _426_/a_1000_472# 0.033582f
C13353 _017_ _135_ 0.094281f
C13354 _443_/a_36_151# _371_/a_36_113# 0.001252f
C13355 _176_ FILLER_0_10_107/a_572_375# 0.012296f
C13356 _098_ _437_/a_1204_472# 0.005729f
C13357 _067_ _450_/a_1040_527# 0.007414f
C13358 FILLER_0_14_50/a_124_375# vss 0.002412f
C13359 FILLER_0_14_50/a_36_472# vdd 0.081414f
C13360 net65 FILLER_0_3_172/a_3260_375# 0.002696f
C13361 output47/a_224_472# net3 0.002186f
C13362 trimb[4] input3/a_36_113# 0.001221f
C13363 FILLER_0_7_104/a_932_472# _131_ 0.011713f
C13364 _402_/a_1948_68# _179_ 0.005403f
C13365 FILLER_0_9_72/a_124_375# vss 0.047932f
C13366 FILLER_0_9_72/a_572_375# vdd -0.014642f
C13367 net80 _435_/a_1000_472# 0.001079f
C13368 ctlp[3] _009_ 0.018168f
C13369 _152_ _160_ 0.286108f
C13370 _011_ _108_ 0.036521f
C13371 net17 net42 0.056318f
C13372 net34 _107_ 0.017589f
C13373 _451_/a_36_151# net14 0.037503f
C13374 net28 net19 0.115252f
C13375 FILLER_0_18_2/a_2724_472# net40 0.011079f
C13376 _000_ _073_ 0.222349f
C13377 _269_/a_36_472# vss 0.014227f
C13378 FILLER_0_16_57/a_1020_375# net55 0.003303f
C13379 FILLER_0_16_57/a_484_472# net72 0.017841f
C13380 FILLER_0_11_142/a_484_472# vss 0.033416f
C13381 output8/a_224_472# FILLER_0_3_221/a_124_375# 0.03228f
C13382 _026_ vss 0.005992f
C13383 _132_ _120_ 0.034714f
C13384 cal_count\[3\] vdd 1.020669f
C13385 _320_/a_36_472# _043_ 0.019162f
C13386 _131_ FILLER_0_18_37/a_1380_472# 0.035078f
C13387 _128_ _246_/a_36_68# 0.01024f
C13388 net57 FILLER_0_13_142/a_124_375# 0.011369f
C13389 net18 _417_/a_448_472# 0.03772f
C13390 FILLER_0_16_107/a_484_472# _132_ 0.005391f
C13391 net20 _429_/a_2248_156# 0.027661f
C13392 FILLER_0_16_89/a_484_472# _131_ 0.01075f
C13393 FILLER_0_12_236/a_36_472# vss 0.001526f
C13394 FILLER_0_12_236/a_484_472# vdd 0.00923f
C13395 FILLER_0_21_206/a_36_472# vdd 0.00971f
C13396 FILLER_0_21_206/a_124_375# vss 0.05074f
C13397 FILLER_0_21_125/a_36_472# _098_ 0.002923f
C13398 net82 FILLER_0_3_221/a_484_472# 0.013492f
C13399 _086_ _131_ 0.886615f
C13400 vdd _416_/a_36_151# 0.142481f
C13401 _097_ vss 0.00839f
C13402 _104_ net18 0.039321f
C13403 output24/a_224_472# FILLER_0_24_130/a_124_375# 0.00515f
C13404 _053_ _165_ 0.123461f
C13405 _103_ vss 0.098913f
C13406 _415_/a_36_151# _416_/a_1308_423# 0.00119f
C13407 _301_/a_36_472# _098_ 0.010091f
C13408 output27/a_224_472# net18 0.058296f
C13409 net62 _006_ 0.136418f
C13410 _140_ net23 0.06742f
C13411 output48/a_224_472# _425_/a_36_151# 0.004037f
C13412 FILLER_0_18_2/a_2364_375# net55 0.005899f
C13413 _119_ _372_/a_170_472# 0.003159f
C13414 FILLER_0_9_28/a_1468_375# _054_ 0.005381f
C13415 FILLER_0_23_88/a_36_472# net14 0.003077f
C13416 _370_/a_848_380# net47 0.004223f
C13417 _119_ _131_ 0.073868f
C13418 net16 _392_/a_36_68# 0.002191f
C13419 FILLER_0_4_152/a_124_375# _386_/a_124_24# 0.010472f
C13420 _091_ _136_ 0.075998f
C13421 result[6] net18 0.026875f
C13422 FILLER_0_15_282/a_36_472# net18 0.036858f
C13423 _098_ _204_/a_67_603# 0.00539f
C13424 _091_ net21 0.030022f
C13425 output45/a_224_472# net43 0.024629f
C13426 vdd net40 1.984115f
C13427 FILLER_0_21_28/a_932_472# vdd 0.04815f
C13428 _211_/a_36_160# vss 0.002041f
C13429 FILLER_0_3_172/a_3172_472# vss 0.003689f
C13430 _115_ _134_ 0.051655f
C13431 fanout61/a_36_113# net18 0.001668f
C13432 _169_ vdd 0.055642f
C13433 _057_ _311_/a_254_473# 0.002364f
C13434 net35 _436_/a_448_472# 0.012374f
C13435 net15 FILLER_0_5_54/a_572_375# 0.002259f
C13436 net65 vdd 1.430654f
C13437 net23 FILLER_0_21_150/a_36_472# 0.016375f
C13438 net52 FILLER_0_2_111/a_124_375# 0.00483f
C13439 output48/a_224_472# net1 0.006536f
C13440 _126_ FILLER_0_11_101/a_124_375# 0.011403f
C13441 cal_itt\[2\] FILLER_0_3_221/a_572_375# 0.060779f
C13442 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_124_375# 0.003732f
C13443 _256_/a_36_68# _077_ 0.027906f
C13444 _093_ vdd 1.439861f
C13445 FILLER_0_22_177/a_1380_472# net33 0.016037f
C13446 net68 _453_/a_796_472# 0.001516f
C13447 FILLER_0_4_107/a_124_375# _157_ 0.001427f
C13448 _091_ _070_ 0.162632f
C13449 net57 FILLER_0_16_154/a_932_472# 0.003453f
C13450 FILLER_0_16_107/a_484_472# FILLER_0_14_107/a_572_375# 0.001404f
C13451 net72 cal_count\[3\] 0.059493f
C13452 net15 FILLER_0_15_72/a_484_472# 0.002925f
C13453 ctln[8] net52 0.005231f
C13454 net15 net50 0.177988f
C13455 net1 net5 0.266194f
C13456 FILLER_0_6_177/a_124_375# _163_ 0.025831f
C13457 FILLER_0_20_107/a_124_375# net71 0.03452f
C13458 _255_/a_224_552# _056_ 0.033615f
C13459 FILLER_0_17_72/a_1916_375# _131_ 0.006589f
C13460 FILLER_0_4_185/a_124_375# _002_ 0.013895f
C13461 _412_/a_36_151# output48/a_224_472# 0.229574f
C13462 _070_ _160_ 0.065914f
C13463 FILLER_0_4_49/a_36_472# vdd 0.090733f
C13464 FILLER_0_4_49/a_572_375# vss 0.008729f
C13465 net74 _332_/a_36_472# 0.003752f
C13466 net33 _297_/a_36_472# 0.00521f
C13467 FILLER_0_11_109/a_124_375# _135_ 0.009057f
C13468 net20 _123_ 0.034801f
C13469 ctlp[2] _420_/a_2665_112# 0.01544f
C13470 net81 FILLER_0_15_212/a_572_375# 0.006974f
C13471 FILLER_0_5_72/a_484_472# net47 0.00169f
C13472 FILLER_0_7_72/a_36_472# _053_ 0.01287f
C13473 state\[0\] _223_/a_36_160# 0.070065f
C13474 net73 _334_/a_36_160# 0.003275f
C13475 net60 net19 0.102311f
C13476 ctln[1] FILLER_0_0_232/a_36_472# 0.005158f
C13477 _448_/a_2665_112# trim_val\[4\] 0.004707f
C13478 output34/a_224_472# _419_/a_2665_112# 0.010731f
C13479 FILLER_0_15_180/a_572_375# vdd 0.068901f
C13480 _128_ net23 0.041791f
C13481 cal_itt\[2\] _000_ 0.042235f
C13482 net59 vdd 2.180407f
C13483 net79 net64 0.049663f
C13484 _428_/a_1308_423# _095_ 0.001504f
C13485 FILLER_0_20_177/a_1468_375# _434_/a_36_151# 0.001822f
C13486 _340_/a_36_160# FILLER_0_20_169/a_124_375# 0.005494f
C13487 _345_/a_36_160# net71 0.002396f
C13488 FILLER_0_16_89/a_124_375# _177_ 0.008257f
C13489 _379_/a_36_472# vdd 0.004183f
C13490 _053_ _079_ 0.007118f
C13491 FILLER_0_14_91/a_36_472# _067_ 0.004194f
C13492 _408_/a_56_524# net47 0.040511f
C13493 net79 mask\[1\] 0.029512f
C13494 output35/a_224_472# vdd 0.064053f
C13495 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_572_375# 0.026339f
C13496 _042_ cal_count\[0\] 0.006265f
C13497 FILLER_0_4_152/a_124_375# vss 0.019426f
C13498 _413_/a_2248_156# net20 0.002515f
C13499 _140_ net33 0.026401f
C13500 net24 FILLER_0_22_86/a_1380_472# 0.003096f
C13501 FILLER_0_17_133/a_36_472# _137_ 0.001963f
C13502 FILLER_0_3_78/a_36_472# vss 0.004461f
C13503 net72 net40 0.001815f
C13504 FILLER_0_8_37/a_484_472# _220_/a_67_603# 0.005759f
C13505 _452_/a_1040_527# net40 0.007832f
C13506 net75 net65 0.135447f
C13507 _095_ FILLER_0_15_72/a_124_375# 0.001474f
C13508 net55 FILLER_0_21_28/a_3260_375# 0.006399f
C13509 net72 FILLER_0_21_28/a_932_472# 0.015756f
C13510 FILLER_0_9_28/a_572_375# _054_ 0.002983f
C13511 net53 _131_ 0.059223f
C13512 FILLER_0_11_142/a_572_375# net23 0.010863f
C13513 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_36_472# 0.086635f
C13514 FILLER_0_4_107/a_36_472# vss 0.002634f
C13515 FILLER_0_4_107/a_484_472# vdd 0.03151f
C13516 _077_ _439_/a_2665_112# 0.035688f
C13517 FILLER_0_8_24/a_124_375# net47 0.025599f
C13518 net67 _450_/a_448_472# 0.068692f
C13519 FILLER_0_12_20/a_124_375# vdd 0.017452f
C13520 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_124_375# 0.001597f
C13521 _435_/a_796_472# vdd 0.003478f
C13522 FILLER_0_17_226/a_36_472# vdd 0.087587f
C13523 mask\[0\] _018_ 0.328328f
C13524 _120_ _453_/a_2665_112# 0.002925f
C13525 FILLER_0_12_20/a_484_472# net17 0.05005f
C13526 _013_ _424_/a_1000_472# 0.037585f
C13527 FILLER_0_19_55/a_36_472# FILLER_0_18_53/a_124_375# 0.001684f
C13528 _254_/a_448_472# _072_ 0.002611f
C13529 FILLER_0_9_72/a_36_472# _439_/a_36_151# 0.001723f
C13530 FILLER_0_4_144/a_36_472# _443_/a_36_151# 0.00271f
C13531 _086_ _126_ 0.063495f
C13532 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1380_472# 0.013276f
C13533 output9/a_224_472# FILLER_0_1_266/a_36_472# 0.001007f
C13534 _094_ FILLER_0_17_282/a_124_375# 0.001151f
C13535 _074_ _251_/a_906_472# 0.002887f
C13536 _077_ calibrate 0.055446f
C13537 FILLER_0_19_125/a_124_375# _433_/a_36_151# 0.001597f
C13538 net55 FILLER_0_17_64/a_124_375# 0.020021f
C13539 vdd FILLER_0_21_60/a_484_472# 0.005181f
C13540 vss FILLER_0_21_60/a_36_472# 0.001384f
C13541 FILLER_0_19_171/a_484_472# _434_/a_36_151# 0.002841f
C13542 _451_/a_1353_112# _040_ 0.005265f
C13543 net50 _376_/a_36_160# 0.018407f
C13544 net63 FILLER_0_18_177/a_1380_472# 0.070445f
C13545 net73 net36 0.073334f
C13546 FILLER_0_9_290/a_36_472# vss 0.011755f
C13547 net75 net59 0.06935f
C13548 FILLER_0_18_2/a_3172_472# FILLER_0_18_37/a_36_472# 0.002765f
C13549 ctln[1] net18 0.004646f
C13550 FILLER_0_3_142/a_36_472# net74 0.001098f
C13551 FILLER_0_5_206/a_36_472# vss 0.003493f
C13552 _394_/a_1336_472# vdd 0.003226f
C13553 _019_ vss 0.10954f
C13554 _150_ _136_ 0.039815f
C13555 net42 _039_ 0.001096f
C13556 net26 FILLER_0_23_44/a_1020_375# 0.001646f
C13557 _413_/a_2560_156# net65 0.011101f
C13558 _144_ _352_/a_257_69# 0.001662f
C13559 _233_/a_36_160# _063_ 0.002771f
C13560 FILLER_0_5_117/a_36_472# net47 0.005919f
C13561 FILLER_0_15_2/a_124_375# vdd 0.010829f
C13562 trim[0] _064_ 0.014422f
C13563 fanout71/a_36_113# FILLER_0_20_107/a_124_375# 0.002853f
C13564 FILLER_0_19_28/a_36_472# net17 0.009277f
C13565 _430_/a_796_472# net36 0.00117f
C13566 _428_/a_2665_112# net53 0.002379f
C13567 net60 _009_ 0.006086f
C13568 _308_/a_124_24# FILLER_0_10_94/a_36_472# 0.001811f
C13569 vss _145_ 0.399701f
C13570 net4 _269_/a_36_472# 0.033296f
C13571 FILLER_0_19_195/a_124_375# vss 0.020433f
C13572 FILLER_0_19_195/a_36_472# vdd 0.094409f
C13573 _432_/a_796_472# _093_ 0.002586f
C13574 _256_/a_2552_68# _076_ 0.00144f
C13575 net41 _402_/a_56_567# 0.021641f
C13576 FILLER_0_13_80/a_124_375# vdd 0.018971f
C13577 _033_ net49 0.003904f
C13578 cal_count\[3\] cal_count\[0\] 0.098735f
C13579 FILLER_0_5_54/a_932_472# net47 0.006386f
C13580 trim[0] output41/a_224_472# 0.018464f
C13581 _389_/a_36_148# vss 0.001935f
C13582 result[2] _005_ 0.060821f
C13583 _411_/a_796_472# _000_ 0.044697f
C13584 net82 FILLER_0_3_172/a_932_472# 0.007986f
C13585 _098_ _201_/a_67_603# 0.005932f
C13586 _128_ _056_ 0.026612f
C13587 net4 FILLER_0_12_236/a_36_472# 0.016315f
C13588 net38 net3 0.103189f
C13589 _150_ _356_/a_36_472# 0.007271f
C13590 FILLER_0_12_220/a_1468_375# _043_ 0.002509f
C13591 _021_ _091_ 0.016024f
C13592 net35 net24 0.01339f
C13593 FILLER_0_18_2/a_1380_472# _452_/a_448_472# 0.059367f
C13594 _185_ _184_ 0.047803f
C13595 net18 _418_/a_448_472# 0.026048f
C13596 result[7] _046_ 0.003397f
C13597 FILLER_0_17_142/a_572_375# vss 0.049716f
C13598 FILLER_0_17_142/a_36_472# vdd 0.108843f
C13599 result[1] vdd 0.221634f
C13600 _039_ clkc 0.003104f
C13601 FILLER_0_17_72/a_2364_375# _150_ 0.001083f
C13602 FILLER_0_18_2/a_484_472# vdd 0.003495f
C13603 net18 _419_/a_2248_156# 0.014287f
C13604 _137_ FILLER_0_16_154/a_1380_472# 0.005667f
C13605 _413_/a_2560_156# net59 0.016463f
C13606 _346_/a_49_472# vdd -0.002208f
C13607 _253_/a_1100_68# _074_ 0.001563f
C13608 _431_/a_2248_156# FILLER_0_15_142/a_572_375# 0.001374f
C13609 _232_/a_255_603# _164_ 0.001274f
C13610 fanout63/a_36_160# net64 0.016132f
C13611 net55 FILLER_0_21_60/a_124_375# 0.015315f
C13612 _258_/a_36_160# _080_ 0.261387f
C13613 FILLER_0_7_72/a_36_472# _028_ 0.020625f
C13614 FILLER_0_18_76/a_124_375# vss 0.006877f
C13615 FILLER_0_18_76/a_572_375# vdd -0.009037f
C13616 net52 _440_/a_36_151# 0.01571f
C13617 net81 _425_/a_2248_156# 0.058229f
C13618 FILLER_0_13_100/a_124_375# _043_ 0.010818f
C13619 result[0] FILLER_0_9_282/a_484_472# 0.018647f
C13620 fanout63/a_36_160# mask\[1\] 0.009907f
C13621 net30 result[3] 0.002746f
C13622 _429_/a_2248_156# vss 0.040729f
C13623 _429_/a_2665_112# vdd 0.010552f
C13624 trim_mask\[1\] FILLER_0_4_91/a_124_375# 0.006803f
C13625 net38 _245_/a_672_472# 0.006341f
C13626 fanout80/a_36_113# net80 0.004615f
C13627 net57 _017_ 0.045694f
C13628 mask\[4\] FILLER_0_19_171/a_572_375# 0.006277f
C13629 FILLER_0_10_247/a_36_472# vss 0.002828f
C13630 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_36_472# 0.026657f
C13631 _129_ FILLER_0_11_135/a_124_375# 0.009882f
C13632 calibrate net37 0.101109f
C13633 ctlp[5] net22 0.001542f
C13634 _075_ _068_ 0.006297f
C13635 _132_ _428_/a_1456_156# 0.001009f
C13636 _104_ _109_ 0.029532f
C13637 trimb[3] ctlp[0] 0.384753f
C13638 result[5] fanout60/a_36_160# 0.001585f
C13639 _069_ state\[2\] 0.023375f
C13640 FILLER_0_17_72/a_2276_472# net36 0.004399f
C13641 FILLER_0_19_125/a_36_472# vdd 0.003414f
C13642 _421_/a_2665_112# _109_ 0.002029f
C13643 net47 _450_/a_36_151# 0.029201f
C13644 _441_/a_2248_156# FILLER_0_3_78/a_572_375# 0.001068f
C13645 _423_/a_2248_156# FILLER_0_23_60/a_124_375# 0.001901f
C13646 _013_ FILLER_0_17_56/a_124_375# 0.001047f
C13647 trim_mask\[2\] FILLER_0_3_78/a_36_472# 0.005209f
C13648 _077_ _125_ 0.017422f
C13649 net52 FILLER_0_6_47/a_3260_375# 0.040612f
C13650 _415_/a_1204_472# net18 0.001828f
C13651 FILLER_0_22_128/a_932_472# vdd 0.004405f
C13652 FILLER_0_22_128/a_484_472# vss 0.002338f
C13653 net20 FILLER_0_24_274/a_124_375# 0.002751f
C13654 FILLER_0_17_200/a_124_375# net22 0.003602f
C13655 net70 _043_ 0.045182f
C13656 _115_ FILLER_0_10_78/a_932_472# 0.013773f
C13657 net32 _421_/a_1308_423# 0.005394f
C13658 output43/a_224_472# net43 0.11662f
C13659 _424_/a_2560_156# vss 0.001554f
C13660 _043_ net47 0.043824f
C13661 _024_ _435_/a_796_472# 0.006511f
C13662 result[6] _420_/a_1000_472# 0.007761f
C13663 net57 _250_/a_36_68# 0.001141f
C13664 FILLER_0_21_28/a_124_375# FILLER_0_20_15/a_1468_375# 0.026339f
C13665 _098_ _023_ 0.004191f
C13666 _086_ _267_/a_224_472# 0.004041f
C13667 _442_/a_1308_423# vdd 0.00782f
C13668 _442_/a_448_472# vss 0.001428f
C13669 _008_ _046_ 0.067769f
C13670 _430_/a_1000_472# _069_ 0.00929f
C13671 _445_/a_36_151# vss 0.009726f
C13672 _445_/a_448_472# vdd 0.007946f
C13673 FILLER_0_9_28/a_36_472# vdd 0.086674f
C13674 _185_ net47 0.185634f
C13675 _029_ vss 0.11129f
C13676 vdd trim[3] 0.147228f
C13677 FILLER_0_9_28/a_932_472# net16 0.017841f
C13678 _369_/a_36_68# _158_ 0.042315f
C13679 _029_ _365_/a_692_472# 0.001426f
C13680 _153_ _157_ 0.050552f
C13681 _428_/a_1308_423# net74 0.0098f
C13682 FILLER_0_15_116/a_572_375# net53 0.012526f
C13683 _181_ _402_/a_1948_68# 0.001223f
C13684 _065_ fanout50/a_36_160# 0.022932f
C13685 _123_ FILLER_0_7_233/a_36_472# 0.002812f
C13686 mask\[5\] FILLER_0_18_177/a_1468_375# 0.002726f
C13687 FILLER_0_10_78/a_484_472# vdd 0.004673f
C13688 _414_/a_2248_156# net59 0.004437f
C13689 _104_ _422_/a_448_472# 0.001955f
C13690 _446_/a_2665_112# trim_val\[1\] 0.001275f
C13691 mask\[3\] _102_ 0.142836f
C13692 trim_val\[4\] _386_/a_1084_68# 0.002659f
C13693 _430_/a_2665_112# mask\[1\] 0.004574f
C13694 _072_ _375_/a_960_497# 0.001322f
C13695 fanout57/a_36_113# trim_val\[4\] 0.078297f
C13696 _274_/a_244_497# net27 0.010334f
C13697 fanout81/a_36_160# net81 0.025745f
C13698 _123_ vss 0.016878f
C13699 _091_ FILLER_0_18_177/a_36_472# 0.012695f
C13700 trim[4] net67 0.06366f
C13701 mask\[7\] _435_/a_1308_423# 0.028235f
C13702 net36 FILLER_0_15_228/a_124_375# 0.00167f
C13703 result[6] _421_/a_2248_156# 0.031832f
C13704 net81 _426_/a_1308_423# 0.002332f
C13705 vdd FILLER_0_22_107/a_124_375# 0.029828f
C13706 FILLER_0_12_20/a_484_472# _039_ 0.006288f
C13707 _070_ _267_/a_36_472# 0.002617f
C13708 FILLER_0_15_212/a_572_375# mask\[1\] 0.012463f
C13709 net50 FILLER_0_2_93/a_484_472# 0.002377f
C13710 result[7] net18 0.098317f
C13711 output32/a_224_472# _094_ 0.005545f
C13712 _411_/a_1000_472# net65 0.001916f
C13713 output9/a_224_472# vdd 0.102412f
C13714 _261_/a_36_160# net47 0.010976f
C13715 _132_ _043_ 0.038747f
C13716 FILLER_0_4_177/a_124_375# net22 0.006125f
C13717 _274_/a_36_68# FILLER_0_12_236/a_484_472# 0.001237f
C13718 _053_ net74 0.09773f
C13719 FILLER_0_15_72/a_124_375# cal_count\[1\] 0.00816f
C13720 net55 _424_/a_2248_156# 0.057967f
C13721 _415_/a_796_472# _004_ 0.005395f
C13722 FILLER_0_4_107/a_1468_375# _154_ 0.005202f
C13723 FILLER_0_4_107/a_572_375# _153_ 0.010165f
C13724 result[8] ctlp[2] 0.068359f
C13725 _341_/a_49_472# _141_ 0.006222f
C13726 FILLER_0_15_142/a_36_472# _136_ 0.003745f
C13727 _411_/a_36_151# ctln[3] 0.004014f
C13728 _412_/a_2665_112# net1 0.063655f
C13729 _413_/a_2248_156# vss 0.004157f
C13730 _120_ vdd 0.750809f
C13731 FILLER_0_20_15/a_1020_375# vdd 0.005198f
C13732 FILLER_0_16_107/a_484_472# vdd 0.02929f
C13733 ctln[6] _442_/a_36_151# 0.007031f
C13734 FILLER_0_18_107/a_572_375# FILLER_0_19_111/a_124_375# 0.058411f
C13735 FILLER_0_14_181/a_36_472# _095_ 0.071989f
C13736 net34 net32 0.330134f
C13737 net17 FILLER_0_20_15/a_484_472# 0.011079f
C13738 _126_ FILLER_0_11_109/a_36_472# 0.00136f
C13739 net79 FILLER_0_12_236/a_36_472# 0.009225f
C13740 net58 net18 0.091503f
C13741 _126_ FILLER_0_11_135/a_36_472# 0.002321f
C13742 mask\[3\] _198_/a_67_603# 0.024102f
C13743 FILLER_0_14_81/a_36_472# _394_/a_1936_472# 0.010394f
C13744 mask\[5\] net80 0.036014f
C13745 FILLER_0_5_198/a_484_472# net37 0.009858f
C13746 _127_ _131_ 0.470047f
C13747 FILLER_0_9_28/a_1468_375# net16 0.005202f
C13748 _273_/a_36_68# FILLER_0_10_214/a_124_375# 0.003707f
C13749 net53 _137_ 0.008376f
C13750 _441_/a_2665_112# net14 0.00104f
C13751 net23 FILLER_0_22_128/a_3260_375# 0.012171f
C13752 _008_ net18 0.113775f
C13753 output36/a_224_472# _094_ 0.001477f
C13754 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_36_472# 0.086635f
C13755 cal_count\[2\] _402_/a_56_567# 0.07745f
C13756 _448_/a_796_472# _037_ 0.009263f
C13757 _134_ FILLER_0_9_105/a_36_472# 0.004375f
C13758 output33/a_224_472# net32 0.018183f
C13759 _431_/a_2665_112# _137_ 0.010924f
C13760 _444_/a_1308_423# net40 0.043396f
C13761 net63 _435_/a_448_472# 0.009878f
C13762 trim[0] _446_/a_448_472# 0.007307f
C13763 FILLER_0_8_107/a_124_375# _131_ 0.001624f
C13764 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_124_375# 0.004426f
C13765 FILLER_0_20_193/a_124_375# vdd 0.009092f
C13766 net34 _422_/a_2248_156# 0.005617f
C13767 net62 FILLER_0_13_212/a_1380_472# 0.059367f
C13768 output12/a_224_472# net22 0.002662f
C13769 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_572_375# 0.086635f
C13770 FILLER_0_4_197/a_1020_375# _088_ 0.013641f
C13771 _439_/a_2248_156# net14 0.001279f
C13772 net41 _452_/a_448_472# 0.052165f
C13773 FILLER_0_9_28/a_2364_375# net68 0.019969f
C13774 _012_ FILLER_0_23_44/a_1380_472# 0.001572f
C13775 _093_ FILLER_0_19_134/a_124_375# 0.003473f
C13776 FILLER_0_9_105/a_572_375# vdd 0.074717f
C13777 _441_/a_448_472# _030_ 0.038429f
C13778 _441_/a_36_151# net49 0.010951f
C13779 net82 net23 0.18994f
C13780 vss _202_/a_36_160# 0.010418f
C13781 _335_/a_257_69# mask\[1\] 0.001543f
C13782 FILLER_0_12_2/a_572_375# net67 0.007509f
C13783 net68 _441_/a_36_151# 0.031891f
C13784 fanout76/a_36_160# net2 0.023033f
C13785 output21/a_224_472# ctlp[3] 0.021951f
C13786 vss _433_/a_2560_156# 0.003477f
C13787 net61 net77 0.986569f
C13788 FILLER_0_18_139/a_1468_375# vss 0.009191f
C13789 FILLER_0_18_139/a_36_472# vdd 0.089771f
C13790 net49 _440_/a_1000_472# 0.020434f
C13791 net9 net8 0.027272f
C13792 FILLER_0_16_154/a_124_375# vdd 0.00439f
C13793 fanout74/a_36_113# net82 0.018392f
C13794 net68 _440_/a_1000_472# 0.002604f
C13795 _094_ vdd 0.717159f
C13796 _100_ vss 0.020176f
C13797 FILLER_0_24_130/a_124_375# vss 0.018125f
C13798 _127_ _428_/a_2665_112# 0.001162f
C13799 net72 _403_/a_224_472# 0.002276f
C13800 _440_/a_2248_156# trim_mask\[1\] 0.004408f
C13801 _370_/a_848_380# vdd -0.001256f
C13802 _370_/a_124_24# vss 0.005764f
C13803 cal_itt\[3\] _079_ 0.015743f
C13804 FILLER_0_11_109/a_36_472# FILLER_0_10_107/a_124_375# 0.001684f
C13805 mask\[7\] FILLER_0_22_128/a_484_472# 0.010605f
C13806 output26/a_224_472# net26 0.047008f
C13807 FILLER_0_3_204/a_36_472# net22 0.036788f
C13808 _430_/a_36_151# net81 0.017255f
C13809 FILLER_0_7_162/a_124_375# net37 0.011644f
C13810 _004_ vss 0.115789f
C13811 _305_/a_36_159# vss 0.003366f
C13812 _178_ _095_ 0.839141f
C13813 trim[1] net66 0.007756f
C13814 _079_ _081_ 1.441057f
C13815 net32 _419_/a_448_472# 0.011757f
C13816 _174_ _179_ 0.003183f
C13817 net81 _005_ 0.003646f
C13818 net55 FILLER_0_17_56/a_36_472# 0.019193f
C13819 _077_ net50 0.312283f
C13820 FILLER_0_14_91/a_484_472# _043_ 0.00134f
C13821 _115_ FILLER_0_9_72/a_932_472# 0.001837f
C13822 net73 FILLER_0_18_107/a_1916_375# 0.014643f
C13823 state\[1\] _043_ 0.1587f
C13824 net68 FILLER_0_6_47/a_1380_472# 0.049638f
C13825 _227_/a_36_160# vdd 0.007828f
C13826 output46/a_224_472# net40 0.002542f
C13827 FILLER_0_18_107/a_572_375# vdd 0.00419f
C13828 FILLER_0_18_107/a_124_375# vss 0.003425f
C13829 FILLER_0_14_181/a_36_472# mask\[1\] 0.006352f
C13830 trim_mask\[1\] FILLER_0_6_47/a_2276_472# 0.006166f
C13831 net39 _445_/a_1000_472# 0.007782f
C13832 _429_/a_36_151# FILLER_0_15_205/a_36_472# 0.001723f
C13833 FILLER_0_9_28/a_572_375# net16 0.042681f
C13834 net33 FILLER_0_22_128/a_3260_375# 0.001178f
C13835 _010_ FILLER_0_23_274/a_36_472# 0.008718f
C13836 output12/a_224_472# net11 0.009336f
C13837 net29 _287_/a_244_68# 0.001262f
C13838 net54 FILLER_0_22_128/a_124_375# 0.032013f
C13839 _433_/a_448_472# _145_ 0.045046f
C13840 FILLER_0_18_37/a_124_375# vdd 0.024546f
C13841 FILLER_0_5_206/a_124_375# FILLER_0_5_198/a_572_375# 0.012001f
C13842 _070_ _113_ 0.01052f
C13843 _052_ FILLER_0_18_37/a_932_472# 0.002749f
C13844 fanout68/a_36_113# _036_ 0.007847f
C13845 FILLER_0_12_220/a_932_472# _060_ 0.002471f
C13846 _030_ _367_/a_692_472# 0.002082f
C13847 _446_/a_2248_156# vdd 0.059236f
C13848 net67 net17 0.04175f
C13849 _421_/a_2248_156# _419_/a_2248_156# 0.001364f
C13850 _427_/a_3041_156# net23 0.001305f
C13851 _377_/a_36_472# net67 0.005639f
C13852 FILLER_0_24_274/a_124_375# vss 0.002674f
C13853 _432_/a_2665_112# FILLER_0_17_200/a_124_375# 0.006271f
C13854 state\[2\] FILLER_0_13_142/a_36_472# 0.022678f
C13855 FILLER_0_11_282/a_36_472# _416_/a_1308_423# 0.001295f
C13856 net56 net53 0.053535f
C13857 net53 FILLER_0_13_142/a_932_472# 0.059367f
C13858 FILLER_0_5_72/a_36_472# vss 0.031034f
C13859 FILLER_0_5_72/a_484_472# vdd 0.002735f
C13860 _303_/a_36_472# FILLER_0_20_87/a_36_472# 0.005725f
C13861 ctln[7] _442_/a_36_151# 0.007057f
C13862 net3 FILLER_0_15_10/a_36_472# 0.002825f
C13863 _270_/a_36_472# _079_ 0.036715f
C13864 FILLER_0_4_144/a_124_375# _081_ 0.004558f
C13865 calibrate _122_ 0.074949f
C13866 output19/a_224_472# _108_ 0.005075f
C13867 FILLER_0_7_72/a_2276_472# FILLER_0_6_90/a_124_375# 0.001684f
C13868 FILLER_0_8_127/a_124_375# _126_ 0.001799f
C13869 _143_ FILLER_0_18_139/a_1380_472# 0.002226f
C13870 _057_ _176_ 0.001304f
C13871 _431_/a_2665_112# net56 0.048214f
C13872 fanout60/a_36_160# net60 0.019034f
C13873 _098_ net23 0.036637f
C13874 _118_ net21 0.007371f
C13875 net15 _038_ 0.078028f
C13876 _127_ _126_ 0.398279f
C13877 _068_ _152_ 0.006744f
C13878 _057_ _306_/a_36_68# 0.019072f
C13879 _143_ FILLER_0_16_154/a_1468_375# 0.002033f
C13880 _093_ _099_ 0.001725f
C13881 _089_ _079_ 0.126206f
C13882 _003_ _087_ 0.054908f
C13883 fanout61/a_36_113# _418_/a_36_151# 0.001442f
C13884 FILLER_0_6_90/a_36_472# _163_ 0.016147f
C13885 _408_/a_56_524# vdd 0.003158f
C13886 _408_/a_728_93# vss 0.001345f
C13887 FILLER_0_5_117/a_124_375# vss 0.001764f
C13888 FILLER_0_2_93/a_572_375# net69 0.015032f
C13889 _410_/a_36_68# _173_ 0.009636f
C13890 vss _107_ 0.186994f
C13891 net7 ctln[0] 0.001209f
C13892 _242_/a_36_160# _386_/a_124_24# 0.031797f
C13893 FILLER_0_12_136/a_1380_472# _126_ 0.014722f
C13894 FILLER_0_19_134/a_36_472# _145_ 0.080913f
C13895 _033_ net47 0.056436f
C13896 _176_ _451_/a_3129_107# 0.021559f
C13897 FILLER_0_7_72/a_124_375# FILLER_0_5_72/a_36_472# 0.001512f
C13898 _069_ FILLER_0_11_142/a_124_375# 0.030279f
C13899 _070_ _118_ 0.302298f
C13900 FILLER_0_18_209/a_124_375# vdd 0.023676f
C13901 net1 en 0.068102f
C13902 net82 trim_val\[4\] 0.511271f
C13903 FILLER_0_7_72/a_572_375# vdd 0.004039f
C13904 FILLER_0_8_24/a_124_375# vdd 0.01166f
C13905 net57 _280_/a_224_472# 0.001032f
C13906 _372_/a_2590_472# vss 0.00106f
C13907 net15 _449_/a_1204_472# 0.01349f
C13908 _096_ net57 0.05086f
C13909 _120_ cal_count\[0\] 0.014209f
C13910 FILLER_0_19_125/a_36_472# _433_/a_36_151# 0.059367f
C13911 output34/a_224_472# net31 0.165772f
C13912 FILLER_0_8_24/a_484_472# net17 0.010321f
C13913 FILLER_0_4_185/a_36_472# _002_ 0.004231f
C13914 net23 _433_/a_2248_156# 0.005588f
C13915 _114_ _115_ 0.148291f
C13916 FILLER_0_22_128/a_932_472# _433_/a_36_151# 0.002841f
C13917 net72 FILLER_0_18_37/a_124_375# 0.05632f
C13918 FILLER_0_4_107/a_124_375# _160_ 0.005906f
C13919 _078_ FILLER_0_6_231/a_36_472# 0.013046f
C13920 _426_/a_1308_423# net64 0.021119f
C13921 FILLER_0_20_177/a_1468_375# mask\[6\] 0.001162f
C13922 net18 _006_ 0.082256f
C13923 input2/a_36_113# input5/a_36_113# 0.01088f
C13924 _185_ _402_/a_718_527# 0.001973f
C13925 _126_ _071_ 0.090032f
C13926 FILLER_0_23_274/a_36_472# vdd 0.010289f
C13927 FILLER_0_23_274/a_124_375# vss 0.017196f
C13928 _072_ _062_ 0.025795f
C13929 output23/a_224_472# FILLER_0_22_128/a_1468_375# 0.00242f
C13930 FILLER_0_16_89/a_1380_472# FILLER_0_17_72/a_3260_375# 0.001723f
C13931 net7 net16 0.033509f
C13932 _141_ _145_ 0.094128f
C13933 _187_ net51 0.04894f
C13934 FILLER_0_16_37/a_124_375# FILLER_0_18_37/a_36_472# 0.001512f
C13935 _073_ _080_ 0.455535f
C13936 net58 _425_/a_2560_156# 0.004835f
C13937 _033_ FILLER_0_6_47/a_124_375# 0.002521f
C13938 FILLER_0_5_148/a_36_472# _160_ 0.001025f
C13939 net57 _386_/a_848_380# 0.041622f
C13940 FILLER_0_9_28/a_124_375# net40 0.047331f
C13941 _449_/a_1000_472# _038_ 0.021492f
C13942 _413_/a_2665_112# net65 0.033675f
C13943 FILLER_0_16_57/a_484_472# _176_ 0.013507f
C13944 _232_/a_67_603# trim_val\[1\] 0.009588f
C13945 net16 _378_/a_224_472# 0.001007f
C13946 _220_/a_67_603# vss 0.001485f
C13947 _068_ net21 0.030836f
C13948 FILLER_0_18_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001684f
C13949 FILLER_0_5_117/a_36_472# vdd 0.092171f
C13950 _256_/a_716_497# net20 0.007413f
C13951 FILLER_0_9_142/a_36_472# _118_ 0.01533f
C13952 FILLER_0_4_197/a_1468_375# _088_ 0.012367f
C13953 net38 _190_/a_36_160# 0.062343f
C13954 _141_ FILLER_0_17_142/a_572_375# 0.029028f
C13955 ctlp[5] _140_ 0.002123f
C13956 _436_/a_36_151# FILLER_0_22_107/a_572_375# 0.059049f
C13957 net65 FILLER_0_2_177/a_572_375# 0.017058f
C13958 net27 vdd 0.88294f
C13959 trim_mask\[4\] net22 0.027368f
C13960 FILLER_0_7_59/a_572_375# trim_mask\[1\] 0.001548f
C13961 _331_/a_448_472# _120_ 0.001496f
C13962 _430_/a_1000_472# net22 0.032221f
C13963 FILLER_0_5_54/a_932_472# vdd 0.003166f
C13964 FILLER_0_5_54/a_484_472# vss 0.001929f
C13965 trimb[1] FILLER_0_20_2/a_484_472# 0.003628f
C13966 cal_count\[2\] _452_/a_448_472# 0.003314f
C13967 net74 FILLER_0_13_142/a_572_375# 0.001412f
C13968 _242_/a_36_160# vss 0.032884f
C13969 _133_ _076_ 0.11688f
C13970 _070_ _068_ 1.019801f
C13971 _093_ FILLER_0_17_218/a_36_472# 0.006994f
C13972 _441_/a_1308_423# _164_ 0.001807f
C13973 FILLER_0_10_28/a_36_472# output6/a_224_472# 0.010475f
C13974 net55 _131_ 0.314732f
C13975 _182_ _041_ 0.08834f
C13976 _193_/a_36_160# output30/a_224_472# 0.018f
C13977 _432_/a_448_472# _091_ 0.050539f
C13978 cal_count\[3\] _171_ 0.00961f
C13979 _273_/a_36_68# _055_ 0.081216f
C13980 net52 FILLER_0_2_101/a_36_472# 0.00749f
C13981 _084_ net8 0.001821f
C13982 ctlp[3] _296_/a_224_472# 0.005335f
C13983 _413_/a_2665_112# net59 0.066623f
C13984 _238_/a_67_603# trim_mask\[3\] 0.028437f
C13985 net54 _436_/a_36_151# 0.004179f
C13986 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_484_472# 0.013276f
C13987 _440_/a_2248_156# _164_ 0.054298f
C13988 _064_ _446_/a_1308_423# 0.001728f
C13989 _122_ FILLER_0_5_198/a_484_472# 0.002999f
C13990 FILLER_0_6_239/a_124_375# FILLER_0_8_239/a_36_472# 0.001512f
C13991 _431_/a_2248_156# vdd 0.00968f
C13992 _151_ vdd 0.157764f
C13993 net57 fanout55/a_36_160# 0.017476f
C13994 net63 FILLER_0_15_205/a_36_472# 0.047903f
C13995 _088_ FILLER_0_4_213/a_572_375# 0.022684f
C13996 result[9] net29 0.001272f
C13997 _432_/a_36_151# FILLER_0_17_161/a_36_472# 0.004847f
C13998 FILLER_0_2_177/a_572_375# net59 0.005397f
C13999 net67 _439_/a_36_151# 0.136402f
C14000 _438_/a_36_151# net71 0.053065f
C14001 _274_/a_1164_497# net64 0.002049f
C14002 result[1] _416_/a_2248_156# 0.001888f
C14003 _332_/a_244_68# _135_ 0.001325f
C14004 FILLER_0_21_142/a_484_472# vdd 0.004917f
C14005 net80 _138_ 0.002053f
C14006 net58 FILLER_0_8_247/a_1380_472# 0.0597f
C14007 _315_/a_244_497# _120_ 0.006419f
C14008 output22/a_224_472# net23 0.008048f
C14009 _008_ _417_/a_36_151# 0.001136f
C14010 net53 _095_ 0.431214f
C14011 net15 FILLER_0_6_47/a_2812_375# 0.002944f
C14012 net19 _196_/a_36_160# 0.027835f
C14013 FILLER_0_20_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001543f
C14014 _091_ _429_/a_1308_423# 0.031247f
C14015 net19 _420_/a_2560_156# 0.010978f
C14016 net44 net40 0.003336f
C14017 FILLER_0_16_107/a_124_375# FILLER_0_16_89/a_1468_375# 0.005439f
C14018 net20 mask\[0\] 0.103301f
C14019 net20 _074_ 0.038279f
C14020 _176_ cal_count\[3\] 0.067683f
C14021 _068_ FILLER_0_9_142/a_36_472# 0.009073f
C14022 _292_/a_36_160# vdd 0.01694f
C14023 FILLER_0_24_63/a_124_375# output25/a_224_472# 0.007304f
C14024 FILLER_0_17_38/a_572_375# vdd 0.01525f
C14025 vdd _450_/a_36_151# 0.08588f
C14026 net20 net32 0.006161f
C14027 FILLER_0_4_144/a_484_472# net47 0.008338f
C14028 net67 FILLER_0_6_47/a_1828_472# 0.001175f
C14029 net75 net27 0.037524f
C14030 _306_/a_36_68# cal_count\[3\] 0.007663f
C14031 net39 net67 0.049482f
C14032 FILLER_0_7_72/a_2364_375# vdd 0.018287f
C14033 _372_/a_170_472# net23 0.025555f
C14034 _098_ _433_/a_796_472# 0.002825f
C14035 _057_ _310_/a_741_69# 0.001002f
C14036 _178_ cal_count\[1\] 0.470244f
C14037 FILLER_0_7_72/a_3172_472# net50 0.001428f
C14038 FILLER_0_3_2/a_36_472# vss 0.004076f
C14039 fanout70/a_36_113# _020_ 0.001266f
C14040 net67 _039_ 0.302826f
C14041 cal_itt\[2\] _080_ 0.062471f
C14042 _043_ vdd 0.827689f
C14043 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3172_472# 0.026657f
C14044 FILLER_0_8_138/a_124_375# _059_ 0.007966f
C14045 net41 _444_/a_36_151# 0.013142f
C14046 FILLER_0_8_127/a_36_472# _062_ 0.01783f
C14047 FILLER_0_21_133/a_36_472# _140_ 0.008378f
C14048 net62 result[2] 0.311075f
C14049 net74 _081_ 0.093806f
C14050 ctlp[1] _419_/a_2560_156# 0.002551f
C14051 _038_ FILLER_0_11_78/a_36_472# 0.001782f
C14052 net64 _005_ 0.006192f
C14053 _161_ _060_ 0.042838f
C14054 _412_/a_2248_156# net5 0.048919f
C14055 FILLER_0_18_2/a_1020_375# net38 0.047331f
C14056 _432_/a_1204_472# vdd 0.004019f
C14057 output14/a_224_472# trim_mask\[3\] 0.001155f
C14058 ctlp[7] net25 0.003141f
C14059 _185_ vdd 0.325358f
C14060 _448_/a_2248_156# net22 0.07925f
C14061 _064_ _160_ 0.006705f
C14062 _005_ mask\[1\] 0.246517f
C14063 _434_/a_2665_112# mask\[6\] 0.026286f
C14064 FILLER_0_16_37/a_124_375# net47 0.002638f
C14065 output15/a_224_472# FILLER_0_0_96/a_124_375# 0.00515f
C14066 result[8] ctlp[1] 0.049662f
C14067 trim_mask\[4\] _076_ 0.001824f
C14068 net34 _105_ 0.784678f
C14069 FILLER_0_21_28/a_2364_375# _012_ 0.017669f
C14070 FILLER_0_18_2/a_3172_472# vdd 0.011201f
C14071 _411_/a_2248_156# _073_ 0.003809f
C14072 FILLER_0_21_142/a_124_375# _140_ 0.016087f
C14073 FILLER_0_24_96/a_36_472# net35 0.002526f
C14074 net16 _186_ 0.225785f
C14075 mask\[7\] _107_ 0.13732f
C14076 _239_/a_36_160# net40 0.010925f
C14077 FILLER_0_15_116/a_484_472# vss 0.003923f
C14078 net68 fanout67/a_36_160# 0.02648f
C14079 FILLER_0_18_2/a_36_472# cal_count\[2\] 0.001929f
C14080 _175_ vdd 0.147794f
C14081 vss FILLER_0_6_37/a_36_472# 0.006755f
C14082 FILLER_0_5_164/a_124_375# _163_ 0.048663f
C14083 _256_/a_1612_497# _076_ 0.001111f
C14084 _093_ FILLER_0_17_104/a_124_375# 0.01418f
C14085 _411_/a_2665_112# ctln[1] 0.004748f
C14086 output36/a_224_472# FILLER_0_14_263/a_124_375# 0.029138f
C14087 _004_ _415_/a_1308_423# 0.002098f
C14088 FILLER_0_4_197/a_572_375# net21 0.041173f
C14089 net57 FILLER_0_2_165/a_36_472# 0.001562f
C14090 FILLER_0_7_72/a_1468_375# _376_/a_36_160# 0.02985f
C14091 FILLER_0_4_197/a_1380_472# vss 0.007979f
C14092 _086_ net74 0.058077f
C14093 fanout72/a_36_113# _095_ 0.001842f
C14094 _149_ FILLER_0_20_98/a_36_472# 0.067283f
C14095 net72 FILLER_0_17_38/a_572_375# 0.010272f
C14096 _261_/a_36_160# vdd 0.0109f
C14097 net36 FILLER_0_20_87/a_124_375# 0.005853f
C14098 output33/a_224_472# _105_ 0.099107f
C14099 _036_ net40 0.599505f
C14100 _120_ FILLER_0_9_72/a_1380_472# 0.001723f
C14101 FILLER_0_10_107/a_36_472# vss 0.003894f
C14102 FILLER_0_10_107/a_484_472# vdd 0.034172f
C14103 _130_ _125_ 0.002745f
C14104 _431_/a_796_472# _137_ 0.002195f
C14105 _420_/a_2560_156# _009_ 0.001487f
C14106 net72 _043_ 0.05655f
C14107 _375_/a_960_497# vdd 0.004471f
C14108 output47/a_224_472# _095_ 0.012266f
C14109 _119_ net74 0.02813f
C14110 net22 _048_ 0.268142f
C14111 net24 FILLER_0_22_107/a_124_375# 0.001023f
C14112 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_36_472# 0.086635f
C14113 trim_mask\[1\] FILLER_0_6_90/a_572_375# 0.001263f
C14114 mask\[4\] FILLER_0_18_177/a_484_472# 0.016924f
C14115 _144_ net54 0.095482f
C14116 net18 _007_ 0.060872f
C14117 _075_ FILLER_0_5_206/a_124_375# 0.001024f
C14118 FILLER_0_20_177/a_484_472# vdd 0.010805f
C14119 FILLER_0_20_177/a_36_472# vss 0.003944f
C14120 _440_/a_1000_472# net47 0.011283f
C14121 net35 FILLER_0_22_86/a_124_375# 0.01209f
C14122 mask\[8\] FILLER_0_22_86/a_572_375# 0.013048f
C14123 _335_/a_49_472# FILLER_0_15_180/a_572_375# 0.001126f
C14124 net52 _442_/a_36_151# 0.029373f
C14125 output46/a_224_472# FILLER_0_20_15/a_1020_375# 0.001274f
C14126 FILLER_0_14_263/a_124_375# vdd 0.026205f
C14127 net50 _447_/a_2248_156# 0.007602f
C14128 ctln[6] _037_ 0.031407f
C14129 calibrate FILLER_0_9_270/a_36_472# 0.00119f
C14130 _153_ _160_ 0.304792f
C14131 FILLER_0_11_142/a_484_472# FILLER_0_13_142/a_572_375# 0.0027f
C14132 net63 _430_/a_2248_156# 0.051057f
C14133 _174_ _181_ 0.079407f
C14134 _069_ _429_/a_796_472# 0.003099f
C14135 FILLER_0_8_2/a_124_375# _054_ 0.001055f
C14136 net70 FILLER_0_16_115/a_36_472# 0.003407f
C14137 FILLER_0_2_111/a_1380_472# FILLER_0_2_127/a_36_472# 0.013276f
C14138 net82 _443_/a_1000_472# 0.008161f
C14139 net50 _439_/a_2560_156# 0.006321f
C14140 _321_/a_2590_472# _176_ 0.001932f
C14141 _069_ _395_/a_1044_488# 0.002244f
C14142 _291_/a_36_160# output18/a_224_472# 0.001175f
C14143 _095_ FILLER_0_14_107/a_36_472# 0.011439f
C14144 FILLER_0_18_177/a_124_375# vdd 0.033102f
C14145 state\[1\] _062_ 0.001179f
C14146 net44 FILLER_0_15_2/a_124_375# 0.017852f
C14147 FILLER_0_4_107/a_124_375# _156_ 0.00268f
C14148 ctln[5] _448_/a_1308_423# 0.004061f
C14149 result[7] _419_/a_1204_472# 0.018181f
C14150 _126_ net23 0.030487f
C14151 FILLER_0_2_127/a_124_375# vdd 0.013496f
C14152 FILLER_0_7_59/a_124_375# net67 0.036499f
C14153 trimb[1] vss 0.048527f
C14154 net79 _100_ 0.170973f
C14155 _141_ FILLER_0_18_139/a_1468_375# 0.005239f
C14156 vdd FILLER_0_10_94/a_572_375# 0.02784f
C14157 _422_/a_1204_472# _009_ 0.009783f
C14158 _453_/a_1308_423# vss 0.003012f
C14159 FILLER_0_16_57/a_1020_375# net15 0.048731f
C14160 _095_ _451_/a_36_151# 0.008311f
C14161 _074_ FILLER_0_5_181/a_36_472# 0.002385f
C14162 _417_/a_36_151# _006_ 0.015561f
C14163 mask\[3\] FILLER_0_16_154/a_1020_375# 0.001996f
C14164 _050_ _208_/a_36_160# 0.001038f
C14165 _004_ net79 0.27387f
C14166 _093_ FILLER_0_17_133/a_124_375# 0.009649f
C14167 FILLER_0_19_171/a_932_472# vss 0.001256f
C14168 FILLER_0_19_171/a_1380_472# vdd 0.03086f
C14169 _091_ FILLER_0_13_212/a_484_472# 0.04953f
C14170 FILLER_0_14_181/a_36_472# FILLER_0_15_180/a_124_375# 0.001723f
C14171 _031_ vss 0.18315f
C14172 FILLER_0_18_2/a_484_472# net44 0.047503f
C14173 _077_ net22 0.049592f
C14174 FILLER_0_13_206/a_36_472# _043_ 0.011439f
C14175 net78 _421_/a_1204_472# 0.006482f
C14176 ctlp[5] _435_/a_36_151# 0.003815f
C14177 _438_/a_1000_472# vss 0.001536f
C14178 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_932_472# 0.026657f
C14179 _129_ _058_ 0.050726f
C14180 _373_/a_1060_68# _090_ 0.002234f
C14181 FILLER_0_16_73/a_124_375# _175_ 0.005727f
C14182 _029_ FILLER_0_5_88/a_36_472# 0.007596f
C14183 net57 _055_ 0.008619f
C14184 net78 _422_/a_36_151# 0.023285f
C14185 net7 output40/a_224_472# 0.006944f
C14186 net53 net74 0.164124f
C14187 output16/a_224_472# ctln[9] 0.08624f
C14188 FILLER_0_15_282/a_572_375# _006_ 0.001054f
C14189 _132_ FILLER_0_16_115/a_36_472# 0.015199f
C14190 _180_ FILLER_0_15_59/a_36_472# 0.087308f
C14191 FILLER_0_18_2/a_1020_375# net55 0.003942f
C14192 _069_ _122_ 0.002164f
C14193 _301_/a_36_472# mask\[8\] 0.016751f
C14194 _137_ FILLER_0_19_155/a_124_375# 0.00129f
C14195 _008_ _418_/a_36_151# 0.016984f
C14196 _074_ cal_itt\[1\] 0.120296f
C14197 _322_/a_848_380# vss 0.026127f
C14198 _450_/a_1040_527# _039_ 0.015478f
C14199 output36/a_224_472# _417_/a_2248_156# 0.023576f
C14200 FILLER_0_18_2/a_3260_375# FILLER_0_19_28/a_484_472# 0.001684f
C14201 _162_ _312_/a_234_472# 0.003812f
C14202 net67 net42 0.101108f
C14203 _043_ cal_count\[0\] 0.019077f
C14204 _074_ FILLER_0_7_233/a_36_472# 0.001341f
C14205 _449_/a_36_151# FILLER_0_13_72/a_36_472# 0.001723f
C14206 FILLER_0_12_136/a_124_375# vdd 0.004378f
C14207 _004_ _416_/a_2665_112# 0.002631f
C14208 _402_/a_1296_93# vdd 0.017239f
C14209 _104_ result[9] 0.169685f
C14210 _050_ _210_/a_67_603# 0.006444f
C14211 FILLER_0_4_197/a_36_472# net76 0.003914f
C14212 _321_/a_1602_69# _120_ 0.00262f
C14213 ctlp[8] _051_ 0.010337f
C14214 trim_val\[4\] _443_/a_2665_112# 0.018733f
C14215 ctlp[6] FILLER_0_24_130/a_36_472# 0.005932f
C14216 _094_ _099_ 0.193065f
C14217 net57 _427_/a_2665_112# 0.016685f
C14218 _185_ cal_count\[0\] 0.008096f
C14219 mask\[0\] vss 0.694674f
C14220 _423_/a_36_151# _012_ 0.021631f
C14221 _013_ _217_/a_36_160# 0.001614f
C14222 _082_ net59 0.004251f
C14223 _074_ vss 0.404343f
C14224 _057_ _250_/a_36_68# 0.014333f
C14225 net41 FILLER_0_20_31/a_124_375# 0.049106f
C14226 net32 vss 0.824307f
C14227 fanout66/a_36_113# _441_/a_36_151# 0.032681f
C14228 FILLER_0_18_2/a_3260_375# _041_ 0.001024f
C14229 _069_ _061_ 0.024151f
C14230 _031_ _369_/a_244_472# 0.002741f
C14231 net69 _369_/a_36_68# 0.008024f
C14232 _086_ FILLER_0_11_142/a_484_472# 0.008338f
C14233 FILLER_0_10_214/a_36_472# _060_ 0.001378f
C14234 result[6] result[9] 0.026511f
C14235 FILLER_0_4_197/a_1020_375# net59 0.008989f
C14236 result[9] FILLER_0_15_282/a_36_472# 0.003213f
C14237 FILLER_0_3_172/a_1828_472# net22 0.009883f
C14238 net81 FILLER_0_10_256/a_124_375# 0.026113f
C14239 input2/a_36_113# rstn 0.002202f
C14240 net45 net43 0.131763f
C14241 result[7] FILLER_0_23_282/a_36_472# 0.014869f
C14242 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1468_375# 0.086635f
C14243 _417_/a_2248_156# vdd 0.004032f
C14244 _074_ FILLER_0_6_177/a_36_472# 0.045576f
C14245 net67 clkc 0.102244f
C14246 _114_ _121_ 0.002513f
C14247 net22 net37 0.03068f
C14248 ctln[6] output13/a_224_472# 0.080817f
C14249 output26/a_224_472# net17 0.004277f
C14250 _424_/a_1000_472# _012_ 0.00675f
C14251 _077_ _076_ 1.895143f
C14252 _328_/a_36_113# FILLER_0_11_109/a_36_472# 0.0161f
C14253 ctlp[3] _422_/a_36_151# 0.002627f
C14254 net41 FILLER_0_19_28/a_484_472# 0.047447f
C14255 fanout72/a_36_113# net74 0.02894f
C14256 FILLER_0_18_53/a_124_375# vdd 0.022f
C14257 net58 _411_/a_2665_112# 0.018133f
C14258 _274_/a_36_68# net27 0.027359f
C14259 net35 FILLER_0_22_177/a_1468_375# 0.048182f
C14260 _137_ net23 0.031218f
C14261 net65 fanout64/a_36_160# 0.214347f
C14262 FILLER_0_22_86/a_36_472# net71 0.005766f
C14263 net62 _248_/a_36_68# 0.002178f
C14264 output47/a_224_472# trimb[4] 0.044883f
C14265 _285_/a_36_472# mask\[1\] 0.036335f
C14266 FILLER_0_3_172/a_1468_375# vdd 0.045181f
C14267 _052_ FILLER_0_21_28/a_1468_375# 0.001757f
C14268 result[0] vdd 0.193436f
C14269 mask\[5\] _144_ 0.38642f
C14270 _422_/a_2248_156# vss 0.001755f
C14271 _422_/a_2665_112# vdd 0.008306f
C14272 net81 net62 0.245647f
C14273 trim_val\[3\] net14 0.01035f
C14274 _033_ vdd 0.509957f
C14275 FILLER_0_21_28/a_124_375# net17 0.005751f
C14276 net80 _143_ 0.023487f
C14277 FILLER_0_16_255/a_124_375# net19 0.008033f
C14278 trim[0] _035_ 0.171633f
C14279 net57 _058_ 0.028536f
C14280 FILLER_0_13_212/a_572_375# _043_ 0.01418f
C14281 _093_ FILLER_0_18_107/a_3260_375# 0.008393f
C14282 net69 net23 0.064573f
C14283 _265_/a_244_68# net59 0.001147f
C14284 _414_/a_36_151# _087_ 0.010359f
C14285 net41 _041_ 0.076779f
C14286 net57 _315_/a_36_68# 0.0036f
C14287 _098_ FILLER_0_15_212/a_1468_375# 0.008327f
C14288 _449_/a_448_472# cal_count\[3\] 0.007511f
C14289 _219_/a_36_160# _058_ 0.014194f
C14290 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_124_375# 0.007947f
C14291 FILLER_0_15_150/a_36_472# vss 0.00975f
C14292 FILLER_0_10_78/a_484_472# _176_ 0.001731f
C14293 net69 _441_/a_2665_112# 0.014995f
C14294 _111_ mask\[9\] 0.127919f
C14295 _120_ _171_ 0.414533f
C14296 net56 FILLER_0_19_155/a_124_375# 0.006762f
C14297 _093_ FILLER_0_16_89/a_36_472# 0.001338f
C14298 _063_ _378_/a_224_472# 0.002323f
C14299 _439_/a_36_151# _453_/a_2248_156# 0.001082f
C14300 net15 FILLER_0_17_64/a_124_375# 0.047331f
C14301 _112_ net59 0.002846f
C14302 net71 _437_/a_2560_156# 0.037081f
C14303 _415_/a_2665_112# vss 0.015461f
C14304 output10/a_224_472# rstn 0.001656f
C14305 fanout74/a_36_113# net69 0.006779f
C14306 net49 trim_mask\[1\] 0.003402f
C14307 _447_/a_2665_112# trim_val\[3\] 0.002721f
C14308 net50 _444_/a_2665_112# 0.023342f
C14309 _187_ _067_ 0.035532f
C14310 net38 _095_ 0.032393f
C14311 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3172_472# 0.026657f
C14312 FILLER_0_0_130/a_36_472# net13 0.002757f
C14313 fanout73/a_36_113# _427_/a_36_151# 0.032681f
C14314 FILLER_0_3_172/a_2724_472# net21 0.009426f
C14315 _166_ _160_ 0.492224f
C14316 ctlp[8] vdd 0.115254f
C14317 FILLER_0_20_98/a_36_472# net14 0.024154f
C14318 mask\[9\] FILLER_0_19_111/a_36_472# 0.285112f
C14319 _001_ vdd 0.122898f
C14320 net68 trim_mask\[1\] 0.054055f
C14321 net20 FILLER_0_6_239/a_36_472# 0.005138f
C14322 _101_ _283_/a_36_472# 0.002471f
C14323 FILLER_0_4_123/a_36_472# net47 0.012399f
C14324 _059_ FILLER_0_8_156/a_36_472# 0.18373f
C14325 net35 FILLER_0_23_88/a_124_375# 0.009071f
C14326 _126_ FILLER_0_12_196/a_124_375# 0.001392f
C14327 _407_/a_36_472# _185_ 0.009281f
C14328 net35 mask\[6\] 0.041818f
C14329 FILLER_0_2_111/a_36_472# vdd 0.033758f
C14330 FILLER_0_2_111/a_1468_375# vss 0.055168f
C14331 _413_/a_1000_472# net65 0.02866f
C14332 _062_ vdd 0.393862f
C14333 output37/a_224_472# vdd 0.082206f
C14334 _176_ _120_ 0.169846f
C14335 _411_/a_1204_472# vss 0.001746f
C14336 output32/a_224_472# _418_/a_2248_156# 0.024448f
C14337 _428_/a_1000_472# _131_ 0.035998f
C14338 _153_ _156_ 0.539362f
C14339 _124_ vss 0.110847f
C14340 _256_/a_716_497# net4 0.001936f
C14341 FILLER_0_18_107/a_3172_472# vss 0.006614f
C14342 _431_/a_1308_423# _137_ 0.008805f
C14343 FILLER_0_9_60/a_572_375# net51 0.002279f
C14344 _017_ cal_count\[3\] 0.003939f
C14345 _076_ net37 0.072179f
C14346 net41 net49 0.392356f
C14347 net78 _419_/a_1000_472# 0.040603f
C14348 FILLER_0_18_100/a_36_472# mask\[9\] 0.005719f
C14349 _016_ FILLER_0_12_136/a_36_472# 0.016227f
C14350 net63 FILLER_0_20_177/a_1468_375# 0.018435f
C14351 FILLER_0_15_150/a_124_375# mask\[2\] 0.002588f
C14352 FILLER_0_5_206/a_36_472# _081_ 0.014328f
C14353 _149_ _437_/a_2665_112# 0.020763f
C14354 _026_ _437_/a_1204_472# 0.022954f
C14355 _022_ _145_ 0.199016f
C14356 net41 net68 0.009755f
C14357 _086_ _321_/a_2034_472# 0.001815f
C14358 net34 _435_/a_1000_472# 0.007444f
C14359 FILLER_0_9_28/a_3172_472# net68 0.007929f
C14360 FILLER_0_8_107/a_36_472# _134_ 0.005632f
C14361 _093_ FILLER_0_17_72/a_1468_375# 0.005785f
C14362 _432_/a_36_151# net57 0.00484f
C14363 trim[4] trim[1] 0.001879f
C14364 net56 net23 0.930833f
C14365 FILLER_0_13_142/a_932_472# net23 0.020589f
C14366 _411_/a_36_151# output11/a_224_472# 0.095813f
C14367 mask\[4\] FILLER_0_19_155/a_36_472# 0.047448f
C14368 FILLER_0_18_2/a_2364_375# output44/a_224_472# 0.032639f
C14369 net81 _429_/a_448_472# 0.018517f
C14370 net75 _001_ 0.056236f
C14371 _413_/a_1000_472# net59 0.018099f
C14372 FILLER_0_5_109/a_572_375# FILLER_0_5_117/a_36_472# 0.086635f
C14373 net50 _160_ 0.048787f
C14374 _250_/a_36_68# cal_count\[3\] 0.004136f
C14375 _441_/a_448_472# _168_ 0.033059f
C14376 _053_ _372_/a_2590_472# 0.001932f
C14377 ctln[1] FILLER_0_0_266/a_124_375# 0.01186f
C14378 result[7] FILLER_0_24_290/a_124_375# 0.005026f
C14379 _098_ FILLER_0_19_171/a_572_375# 0.001946f
C14380 _142_ FILLER_0_17_142/a_484_472# 0.01467f
C14381 FILLER_0_16_89/a_572_375# net36 0.003629f
C14382 _414_/a_2665_112# net59 0.010265f
C14383 FILLER_0_11_101/a_36_472# net14 0.04522f
C14384 _098_ FILLER_0_15_235/a_572_375# 0.001343f
C14385 FILLER_0_4_144/a_36_472# vss 0.008308f
C14386 FILLER_0_4_144/a_484_472# vdd 0.004027f
C14387 FILLER_0_4_197/a_124_375# _002_ 0.001406f
C14388 net16 _013_ 0.060401f
C14389 net32 mask\[7\] 0.01969f
C14390 ctln[5] vss 0.132862f
C14391 net76 FILLER_0_5_212/a_124_375# 0.004635f
C14392 _258_/a_36_160# net20 0.041584f
C14393 valid net2 0.062523f
C14394 _091_ _069_ 0.741596f
C14395 FILLER_0_4_197/a_1468_375# net59 0.050218f
C14396 _074_ net4 0.088616f
C14397 _085_ _121_ 0.027373f
C14398 FILLER_0_8_127/a_124_375# net74 0.026604f
C14399 _429_/a_796_472# net22 0.020124f
C14400 _053_ _220_/a_67_603# 0.065611f
C14401 FILLER_0_4_144/a_572_375# FILLER_0_5_148/a_124_375# 0.05841f
C14402 FILLER_0_1_98/a_124_375# trim_mask\[3\] 0.058544f
C14403 net17 _452_/a_1353_112# 0.038603f
C14404 _450_/a_1040_527# clkc 0.001412f
C14405 _127_ net74 0.0588f
C14406 FILLER_0_17_72/a_1828_472# vdd 0.001969f
C14407 FILLER_0_17_72/a_1380_472# vss 0.003698f
C14408 _228_/a_36_68# _113_ 0.021898f
C14409 fanout57/a_36_113# trim_mask\[4\] 0.002404f
C14410 FILLER_0_21_206/a_124_375# _204_/a_67_603# 0.003591f
C14411 _068_ FILLER_0_5_148/a_36_472# 0.003015f
C14412 FILLER_0_7_72/a_3260_375# vdd 0.008342f
C14413 _430_/a_36_151# _019_ 0.019296f
C14414 FILLER_0_16_37/a_124_375# vdd 0.038329f
C14415 FILLER_0_5_128/a_484_472# net47 0.009309f
C14416 net18 FILLER_0_9_270/a_484_472# 0.004375f
C14417 FILLER_0_7_72/a_1020_375# net50 0.014749f
C14418 fanout67/a_36_160# FILLER_0_9_60/a_124_375# 0.02985f
C14419 _077_ _255_/a_224_552# 0.025141f
C14420 _104_ net61 1.149805f
C14421 _053_ FILLER_0_5_54/a_484_472# 0.001135f
C14422 _098_ FILLER_0_20_98/a_36_472# 0.0127f
C14423 net61 _421_/a_2665_112# 0.001339f
C14424 net60 _421_/a_1204_472# 0.021679f
C14425 _418_/a_2248_156# vdd 0.00423f
C14426 net15 _423_/a_1308_423# 0.001999f
C14427 _422_/a_2248_156# mask\[7\] 0.015008f
C14428 _449_/a_36_151# _394_/a_728_93# 0.002727f
C14429 net52 _443_/a_2560_156# 0.020855f
C14430 _426_/a_36_151# _425_/a_36_151# 0.006252f
C14431 cal valid 0.06045f
C14432 net57 _428_/a_796_472# 0.003017f
C14433 _091_ FILLER_0_15_212/a_36_472# 0.007355f
C14434 en_co_clk _038_ 0.014475f
C14435 net61 _422_/a_1308_423# 0.002171f
C14436 net60 _422_/a_36_151# 0.008119f
C14437 _450_/a_3129_107# net40 0.034729f
C14438 _426_/a_2248_156# calibrate 0.004597f
C14439 cal_count\[3\] FILLER_0_11_109/a_124_375# 0.004618f
C14440 FILLER_0_0_198/a_36_472# net11 0.056269f
C14441 _011_ vdd 0.182751f
C14442 FILLER_0_7_72/a_2364_375# FILLER_0_6_90/a_484_472# 0.001684f
C14443 _140_ FILLER_0_21_150/a_124_375# 0.019084f
C14444 _136_ FILLER_0_17_142/a_124_375# 0.001315f
C14445 clk net18 0.003519f
C14446 FILLER_0_4_213/a_572_375# net59 0.061684f
C14447 net55 _095_ 0.055644f
C14448 cal_count\[3\] FILLER_0_11_135/a_124_375# 0.004365f
C14449 _453_/a_2560_156# net51 0.013556f
C14450 result[6] net61 0.120359f
C14451 net2 net9 0.001033f
C14452 _402_/a_2172_497# _180_ 0.001094f
C14453 FILLER_0_9_28/a_2364_375# vdd 0.004562f
C14454 FILLER_0_16_89/a_1380_472# net14 0.049391f
C14455 _428_/a_448_472# _043_ 0.063478f
C14456 FILLER_0_12_2/a_484_472# _039_ 0.003082f
C14457 _140_ net71 0.005182f
C14458 FILLER_0_16_73/a_36_472# net55 0.002576f
C14459 net57 net52 0.016136f
C14460 net61 fanout61/a_36_113# 0.023179f
C14461 FILLER_0_4_107/a_1380_472# net47 0.008874f
C14462 net15 _424_/a_2248_156# 0.00415f
C14463 FILLER_0_12_20/a_36_472# net47 0.020589f
C14464 cal_count\[2\] _041_ 0.02197f
C14465 _412_/a_2248_156# en 0.022108f
C14466 _052_ _424_/a_1308_423# 0.008633f
C14467 net34 FILLER_0_22_128/a_1380_472# 0.001011f
C14468 _403_/a_224_472# _183_ 0.007508f
C14469 _441_/a_36_151# vdd 0.098562f
C14470 _098_ _434_/a_796_472# 0.001383f
C14471 net49 _164_ 0.428468f
C14472 _449_/a_2665_112# net55 0.057694f
C14473 FILLER_0_21_133/a_36_472# _098_ 0.002964f
C14474 trimb[4] net38 0.124219f
C14475 _057_ _096_ 0.001547f
C14476 _093_ _020_ 0.015474f
C14477 net15 _447_/a_2665_112# 0.063341f
C14478 _394_/a_56_524# FILLER_0_15_59/a_572_375# 0.003413f
C14479 mask\[3\] FILLER_0_18_177/a_1020_375# 0.002924f
C14480 _016_ vdd 0.114288f
C14481 net68 _164_ 0.189377f
C14482 FILLER_0_16_255/a_36_472# vss 0.00184f
C14483 net63 _434_/a_2665_112# 0.120476f
C14484 net62 net64 0.078454f
C14485 _122_ net22 0.024638f
C14486 _447_/a_36_151# net17 0.001448f
C14487 _440_/a_796_472# vss 0.001285f
C14488 net55 FILLER_0_17_72/a_484_472# 0.019636f
C14489 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_36_472# 0.012267f
C14490 FILLER_0_3_204/a_36_472# net82 0.008268f
C14491 _081_ _123_ 0.007811f
C14492 trimb[0] net17 0.006176f
C14493 _044_ vdd 0.406979f
C14494 fanout62/a_36_160# FILLER_0_13_290/a_124_375# 0.001138f
C14495 FILLER_0_16_37/a_124_375# net72 0.013591f
C14496 net62 mask\[1\] 0.227329f
C14497 net52 _037_ 0.103749f
C14498 FILLER_0_20_87/a_36_472# _437_/a_36_151# 0.001723f
C14499 FILLER_0_5_72/a_1380_472# net49 0.002057f
C14500 _256_/a_36_68# _068_ 0.029112f
C14501 FILLER_0_21_142/a_124_375# _098_ 0.006558f
C14502 _036_ _446_/a_2248_156# 0.001763f
C14503 result[7] result[9] 1.21288f
C14504 _443_/a_1204_472# _170_ 0.002808f
C14505 _056_ _060_ 0.085489f
C14506 _061_ _090_ 0.00832f
C14507 net1 _265_/a_916_472# 0.002088f
C14508 FILLER_0_16_107/a_124_375# vss 0.002683f
C14509 trim_val\[4\] FILLER_0_3_172/a_124_375# 0.002076f
C14510 FILLER_0_19_47/a_572_375# vdd 0.019566f
C14511 FILLER_0_19_47/a_124_375# vss 0.002211f
C14512 _131_ FILLER_0_17_104/a_1468_375# 0.006022f
C14513 net16 _179_ 0.007397f
C14514 _095_ net23 0.053365f
C14515 vss FILLER_0_16_115/a_124_375# 0.006358f
C14516 vdd FILLER_0_16_115/a_36_472# 0.093403f
C14517 _395_/a_244_68# _070_ 0.001481f
C14518 FILLER_0_6_47/a_1380_472# vdd 0.002735f
C14519 FILLER_0_9_72/a_36_472# _453_/a_2248_156# 0.013656f
C14520 FILLER_0_4_144/a_124_375# net23 0.011315f
C14521 _316_/a_124_24# vdd 0.033047f
C14522 result[2] net18 0.086474f
C14523 _444_/a_2665_112# _054_ 0.003576f
C14524 ctlp[5] output22/a_224_472# 0.024131f
C14525 input4/a_36_68# vdd 0.09828f
C14526 FILLER_0_6_239/a_36_472# vss 0.003177f
C14527 net58 net37 0.15273f
C14528 FILLER_0_17_72/a_2812_375# net14 0.018463f
C14529 _144_ _348_/a_49_472# 0.037768f
C14530 _061_ net22 0.123662f
C14531 _418_/a_36_151# _007_ 0.007397f
C14532 net41 FILLER_0_18_37/a_36_472# 0.007459f
C14533 _152_ FILLER_0_5_136/a_36_472# 0.049485f
C14534 FILLER_0_9_28/a_2724_472# net68 0.010755f
C14535 net53 FILLER_0_17_142/a_572_375# 0.023771f
C14536 output31/a_224_472# _417_/a_448_472# 0.008149f
C14537 _367_/a_244_472# vdd 0.001113f
C14538 FILLER_0_21_206/a_36_472# mask\[6\] 0.015735f
C14539 FILLER_0_22_86/a_1468_375# net14 0.024975f
C14540 _091_ FILLER_0_19_171/a_1020_375# 0.005708f
C14541 FILLER_0_5_212/a_36_472# _078_ 0.002235f
C14542 _374_/a_36_68# _062_ 0.004248f
C14543 net28 _045_ 0.05144f
C14544 _065_ vss 0.230397f
C14545 fanout77/a_36_113# _094_ 0.002244f
C14546 _431_/a_2665_112# FILLER_0_17_142/a_572_375# 0.001092f
C14547 _324_/a_224_472# net74 0.001704f
C14548 _077_ _128_ 0.005311f
C14549 _105_ vss 0.485198f
C14550 _448_/a_796_472# net59 0.004855f
C14551 FILLER_0_10_78/a_124_375# _077_ 0.001886f
C14552 FILLER_0_10_78/a_572_375# vdd -0.014642f
C14553 _149_ net71 0.827628f
C14554 net34 net54 0.003682f
C14555 _387_/a_36_113# _037_ 0.003577f
C14556 _427_/a_36_151# vss 0.019281f
C14557 FILLER_0_0_96/a_36_472# vss 0.00344f
C14558 net68 FILLER_0_8_37/a_124_375# 0.004818f
C14559 net48 net59 0.015963f
C14560 _008_ result[9] 0.048497f
C14561 mask\[0\] net79 0.243338f
C14562 trim_mask\[4\] _158_ 0.022724f
C14563 net28 _192_/a_67_603# 0.119061f
C14564 FILLER_0_3_221/a_36_472# net59 0.075858f
C14565 net65 net19 0.044106f
C14566 net15 _098_ 0.003965f
C14567 _093_ FILLER_0_18_177/a_2812_375# 0.001989f
C14568 net75 _316_/a_124_24# 0.003078f
C14569 output35/a_224_472# FILLER_0_22_177/a_1468_375# 0.018187f
C14570 _401_/a_244_472# _180_ 0.001689f
C14571 _242_/a_36_160# FILLER_0_5_164/a_36_472# 0.193804f
C14572 _127_ FILLER_0_11_142/a_484_472# 0.001177f
C14573 _095_ FILLER_0_15_10/a_36_472# 0.00335f
C14574 _068_ calibrate 0.110297f
C14575 _076_ _122_ 0.097035f
C14576 net54 _354_/a_49_472# 0.002169f
C14577 vss FILLER_0_8_156/a_124_375# 0.001766f
C14578 vdd FILLER_0_8_156/a_572_375# 0.014611f
C14579 _002_ FILLER_0_3_172/a_2812_375# 0.006403f
C14580 net44 _450_/a_36_151# 0.026203f
C14581 _437_/a_2665_112# net14 0.002936f
C14582 _411_/a_448_472# _000_ 0.073053f
C14583 FILLER_0_7_104/a_484_472# FILLER_0_9_105/a_572_375# 0.001188f
C14584 net41 _184_ 0.065857f
C14585 _412_/a_1308_423# cal_itt\[1\] 0.009991f
C14586 FILLER_0_17_38/a_484_472# _041_ 0.009607f
C14587 _180_ vss 0.106022f
C14588 ctln[1] input1/a_36_113# 0.004419f
C14589 _449_/a_36_151# _067_ 0.031377f
C14590 net50 _156_ 0.020099f
C14591 fanout51/a_36_113# vss 0.0844f
C14592 _113_ FILLER_0_12_196/a_36_472# 0.002495f
C14593 FILLER_0_22_177/a_932_472# _435_/a_36_151# 0.001723f
C14594 _114_ FILLER_0_10_94/a_36_472# 0.08191f
C14595 net32 _295_/a_36_472# 0.002637f
C14596 _033_ _444_/a_1308_423# 0.002877f
C14597 FILLER_0_12_136/a_932_472# cal_count\[3\] 0.007247f
C14598 _068_ _311_/a_1920_473# 0.001498f
C14599 _394_/a_1936_472# _175_ 0.017848f
C14600 _443_/a_36_151# FILLER_0_2_127/a_36_472# 0.006095f
C14601 _427_/a_2560_156# _095_ 0.009888f
C14602 FILLER_0_15_205/a_36_472# net21 0.007503f
C14603 _370_/a_124_24# _081_ 0.015048f
C14604 FILLER_0_14_81/a_124_375# net55 0.038949f
C14605 _431_/a_448_472# vss 0.005583f
C14606 _125_ _118_ 0.239695f
C14607 result[4] result[3] 0.089939f
C14608 _235_/a_67_603# _447_/a_36_151# 0.038675f
C14609 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3260_375# 0.086905f
C14610 _451_/a_2225_156# vss 0.003848f
C14611 net19 net59 0.0206f
C14612 _305_/a_36_159# _081_ 0.039192f
C14613 output42/a_224_472# vss 0.00418f
C14614 cal_count\[3\] _373_/a_244_68# 0.002341f
C14615 output35/a_224_472# _205_/a_36_160# 0.002043f
C14616 net61 _418_/a_448_472# 0.001253f
C14617 trim_mask\[1\] net47 0.306848f
C14618 FILLER_0_5_128/a_572_375# vss 0.057605f
C14619 FILLER_0_3_54/a_36_472# net40 0.069702f
C14620 net60 _419_/a_1000_472# 0.028992f
C14621 net61 _419_/a_2248_156# 0.022159f
C14622 _258_/a_36_160# vss 0.005039f
C14623 _096_ cal_count\[3\] 0.016393f
C14624 _061_ _076_ 0.024289f
C14625 trimb[4] net55 0.01379f
C14626 trimb[4] _452_/a_3129_107# 0.004943f
C14627 _443_/a_1000_472# net69 0.008276f
C14628 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_36_472# 0.026657f
C14629 _070_ FILLER_0_5_136/a_36_472# 0.029293f
C14630 output13/a_224_472# net52 0.018089f
C14631 FILLER_0_5_172/a_124_375# net37 0.014083f
C14632 net82 trim_mask\[4\] 0.21475f
C14633 net55 net74 0.048927f
C14634 FILLER_0_18_177/a_3172_472# vdd 0.002358f
C14635 FILLER_0_14_99/a_124_375# FILLER_0_13_100/a_36_472# 0.001597f
C14636 output35/a_224_472# mask\[6\] 0.069819f
C14637 _176_ _043_ 0.04106f
C14638 net35 FILLER_0_22_128/a_1468_375# 0.015932f
C14639 _414_/a_1000_472# vdd 0.002568f
C14640 _069_ _267_/a_36_472# 0.003607f
C14641 net20 FILLER_0_6_231/a_124_375# 0.060499f
C14642 _306_/a_36_68# _043_ 0.001086f
C14643 _079_ FILLER_0_5_198/a_36_472# 0.012251f
C14644 _088_ FILLER_0_5_198/a_572_375# 0.001374f
C14645 _335_/a_49_472# _043_ 0.00367f
C14646 fanout71/a_36_113# _149_ 0.001315f
C14647 vss FILLER_0_13_72/a_36_472# 0.034188f
C14648 net51 vss 0.21065f
C14649 net55 cal_count\[1\] 0.204733f
C14650 FILLER_0_16_57/a_932_472# vss 0.003388f
C14651 FILLER_0_16_57/a_1380_472# vdd 0.005673f
C14652 trim_mask\[1\] FILLER_0_6_47/a_124_375# 0.005902f
C14653 result[8] net33 0.474056f
C14654 net41 net47 0.19549f
C14655 mask\[5\] _346_/a_257_69# 0.001764f
C14656 _303_/a_36_472# vdd 0.015964f
C14657 output24/a_224_472# net54 0.177947f
C14658 _102_ vdd 0.211559f
C14659 _114_ FILLER_0_12_136/a_572_375# 0.006974f
C14660 _308_/a_848_380# vdd 0.013895f
C14661 _093_ _111_ 0.555171f
C14662 FILLER_0_7_146/a_124_375# _062_ 0.028312f
C14663 _176_ _175_ 0.054439f
C14664 _091_ _090_ 0.117348f
C14665 _150_ _438_/a_36_151# 0.032532f
C14666 _444_/a_448_472# net17 0.022222f
C14667 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_124_375# 0.026339f
C14668 _065_ trim_mask\[2\] 0.002792f
C14669 FILLER_0_2_93/a_484_472# net14 0.019214f
C14670 fanout79/a_36_160# vdd 0.099877f
C14671 _065_ _447_/a_1308_423# 0.024822f
C14672 net74 net23 0.0064f
C14673 vss _047_ 0.070755f
C14674 net39 trim[1] 0.115976f
C14675 _005_ _100_ 0.004305f
C14676 _073_ FILLER_0_3_221/a_1468_375# 0.006377f
C14677 _148_ _352_/a_257_69# 0.001417f
C14678 trim[0] output40/a_224_472# 0.005306f
C14679 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_484_472# 0.013276f
C14680 output13/a_224_472# _387_/a_36_113# 0.020974f
C14681 _446_/a_1308_423# _035_ 0.002639f
C14682 net81 FILLER_0_9_270/a_124_375# 0.014206f
C14683 _127_ _321_/a_2034_472# 0.003159f
C14684 _273_/a_36_68# _070_ 0.013247f
C14685 _372_/a_2034_472# _152_ 0.00171f
C14686 _129_ _152_ 0.041257f
C14687 _004_ _005_ 0.004158f
C14688 FILLER_0_4_123/a_36_472# vdd 0.091386f
C14689 FILLER_0_4_123/a_124_375# vss 0.009712f
C14690 FILLER_0_13_65/a_124_375# _043_ 0.013045f
C14691 FILLER_0_14_181/a_124_375# _043_ 0.008393f
C14692 mask\[8\] _025_ 0.036686f
C14693 _053_ _074_ 0.503728f
C14694 _015_ _426_/a_2248_156# 0.021465f
C14695 mask\[4\] _091_ 0.071954f
C14696 _176_ FILLER_0_10_107/a_484_472# 0.009571f
C14697 _091_ net22 0.031921f
C14698 _386_/a_848_380# _169_ 0.001355f
C14699 _386_/a_124_24# _163_ 0.001234f
C14700 _144_ _350_/a_49_472# 0.033348f
C14701 _098_ _437_/a_2665_112# 0.003567f
C14702 fanout74/a_36_113# net74 0.007425f
C14703 net65 FILLER_0_3_172/a_484_472# 0.003678f
C14704 net65 _386_/a_848_380# 0.00123f
C14705 _096_ FILLER_0_15_180/a_572_375# 0.001972f
C14706 FILLER_0_9_72/a_1468_375# vdd 0.026475f
C14707 FILLER_0_9_72/a_1020_375# vss 0.005622f
C14708 result[9] _006_ 0.05748f
C14709 net27 _426_/a_448_472# 0.023676f
C14710 _414_/a_2560_156# _074_ 0.001344f
C14711 _144_ net73 0.003657f
C14712 result[1] net19 0.084617f
C14713 _451_/a_1353_112# net14 0.041814f
C14714 _256_/a_244_497# calibrate 0.002421f
C14715 result[7] net61 0.021122f
C14716 net55 FILLER_0_13_72/a_124_375# 0.00281f
C14717 _105_ mask\[7\] 0.486236f
C14718 FILLER_0_24_96/a_124_375# output25/a_224_472# 0.002633f
C14719 net15 _131_ 0.037758f
C14720 _086_ FILLER_0_5_117/a_124_375# 0.003725f
C14721 _182_ vdd 0.161134f
C14722 fanout51/a_36_113# FILLER_0_11_64/a_124_375# 0.002335f
C14723 mask\[5\] net34 0.041303f
C14724 FILLER_0_7_195/a_36_472# _072_ 0.008357f
C14725 _198_/a_67_603# vdd 0.015843f
C14726 net20 _073_ 0.437482f
C14727 _120_ _450_/a_3129_107# 0.001598f
C14728 _093_ FILLER_0_18_100/a_36_472# 0.077197f
C14729 output8/a_224_472# FILLER_0_3_221/a_1020_375# 0.03228f
C14730 FILLER_0_15_150/a_124_375# vss 0.01957f
C14731 _173_ FILLER_0_12_28/a_36_472# 0.001633f
C14732 _193_/a_36_160# _416_/a_36_151# 0.065269f
C14733 _188_ vdd 0.022839f
C14734 net67 FILLER_0_8_24/a_484_472# 0.001065f
C14735 net57 FILLER_0_13_142/a_1020_375# 0.009442f
C14736 net18 _417_/a_796_472# 0.006722f
C14737 net20 _429_/a_2560_156# 0.002069f
C14738 FILLER_0_16_89/a_1380_472# _131_ 0.004201f
C14739 FILLER_0_9_223/a_124_375# _055_ 0.014525f
C14740 net82 FILLER_0_3_221/a_1380_472# 0.008049f
C14741 _119_ FILLER_0_5_117/a_124_375# 0.002747f
C14742 FILLER_0_15_282/a_124_375# output30/a_224_472# 0.029138f
C14743 vdd _416_/a_1308_423# 0.002623f
C14744 vss _416_/a_448_472# 0.004806f
C14745 net80 net36 0.036729f
C14746 fanout67/a_36_160# vdd 0.018829f
C14747 vss net6 0.096009f
C14748 _137_ FILLER_0_17_104/a_1468_375# 0.002679f
C14749 net65 cal_itt\[0\] 0.07564f
C14750 _057_ _055_ 0.290639f
C14751 mask\[2\] FILLER_0_16_154/a_572_375# 0.026605f
C14752 FILLER_0_13_142/a_124_375# _043_ 0.009328f
C14753 _035_ _160_ 0.120469f
C14754 net81 net18 0.102876f
C14755 _176_ FILLER_0_10_94/a_572_375# 0.011743f
C14756 _140_ FILLER_0_22_128/a_2812_375# 0.003154f
C14757 mask\[5\] output33/a_224_472# 0.0238f
C14758 _081_ _242_/a_36_160# 0.025059f
C14759 mask\[0\] FILLER_0_15_212/a_572_375# 0.001158f
C14760 _283_/a_36_472# vdd 0.092097f
C14761 ctln[7] FILLER_0_0_96/a_124_375# 0.025944f
C14762 trimb[0] trimb[3] 0.549457f
C14763 net63 net35 0.126544f
C14764 FILLER_0_11_109/a_124_375# _120_ 0.016902f
C14765 cal_count\[2\] _184_ 0.033241f
C14766 _018_ _138_ 0.008093f
C14767 vdd trim[2] 0.166648f
C14768 FILLER_0_21_28/a_1828_472# vdd 0.004227f
C14769 FILLER_0_21_28/a_1380_472# vss 0.001688f
C14770 _050_ vdd 0.484554f
C14771 net20 output20/a_224_472# 0.024692f
C14772 _163_ vss 0.638066f
C14773 _057_ _311_/a_1212_473# 0.004869f
C14774 FILLER_0_11_135/a_124_375# _120_ 0.017316f
C14775 net35 _436_/a_796_472# 0.002146f
C14776 mask\[8\] _436_/a_1000_472# 0.001091f
C14777 _008_ net61 0.004059f
C14778 _443_/a_2248_156# net22 0.001984f
C14779 net15 FILLER_0_5_54/a_1468_375# 0.039975f
C14780 FILLER_0_10_37/a_36_472# FILLER_0_8_37/a_124_375# 0.001512f
C14781 net71 net14 0.147175f
C14782 FILLER_0_11_64/a_124_375# net51 0.027848f
C14783 _126_ FILLER_0_11_101/a_36_472# 0.062336f
C14784 net52 FILLER_0_2_111/a_1020_375# 0.00245f
C14785 cal_itt\[2\] FILLER_0_3_221/a_1468_375# 0.016021f
C14786 _372_/a_170_472# _133_ 0.031518f
C14787 _069_ _113_ 0.027402f
C14788 fanout58/a_36_160# net59 0.048057f
C14789 _131_ _133_ 0.20118f
C14790 _129_ _070_ 0.056776f
C14791 fanout62/a_36_160# FILLER_0_11_282/a_36_472# 0.005262f
C14792 net72 _182_ 0.044895f
C14793 net47 _164_ 0.118311f
C14794 _115_ vss 0.372063f
C14795 result[2] FILLER_0_15_282/a_572_375# 0.0011f
C14796 FILLER_0_2_101/a_124_375# _157_ 0.002818f
C14797 FILLER_0_6_177/a_36_472# _163_ 0.025039f
C14798 ctln[8] net50 0.0032f
C14799 _144_ _143_ 0.001774f
C14800 FILLER_0_17_72/a_2812_375# _131_ 0.006589f
C14801 net16 _181_ 0.48682f
C14802 _076_ _160_ 0.006506f
C14803 FILLER_0_4_49/a_484_472# vss 0.002751f
C14804 _077_ net14 0.03359f
C14805 vdd FILLER_0_14_235/a_124_375# -0.011193f
C14806 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_572_375# 0.086635f
C14807 net81 FILLER_0_15_212/a_1468_375# 0.006906f
C14808 net65 FILLER_0_2_171/a_36_472# 0.023858f
C14809 FILLER_0_5_72/a_1380_472# net47 0.003924f
C14810 _341_/a_49_472# net23 0.031763f
C14811 FILLER_0_21_28/a_124_375# FILLER_0_19_28/a_36_472# 0.001512f
C14812 net80 FILLER_0_20_169/a_36_472# 0.024142f
C14813 FILLER_0_3_204/a_36_472# FILLER_0_3_212/a_36_472# 0.002296f
C14814 FILLER_0_15_180/a_484_472# vdd 0.037927f
C14815 FILLER_0_15_180/a_36_472# vss 0.00138f
C14816 net32 ctlp[2] 0.097138f
C14817 output9/a_224_472# net19 0.070689f
C14818 cal_itt\[2\] net20 0.715447f
C14819 _415_/a_2248_156# vss 0.00818f
C14820 net66 FILLER_0_3_54/a_124_375# 0.038548f
C14821 net50 fanout49/a_36_160# 0.059373f
C14822 _428_/a_1000_472# _095_ 0.001101f
C14823 FILLER_0_5_72/a_124_375# _440_/a_36_151# 0.059049f
C14824 FILLER_0_20_177/a_484_472# _434_/a_36_151# 0.001723f
C14825 _164_ FILLER_0_6_47/a_124_375# 0.069738f
C14826 net80 _432_/a_2248_156# 0.059406f
C14827 _000_ _253_/a_244_68# 0.001243f
C14828 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_484_472# 0.001723f
C14829 _069_ _118_ 0.010986f
C14830 _140_ _049_ 0.003069f
C14831 _052_ _216_/a_67_603# 0.006658f
C14832 net2 calibrate 0.003482f
C14833 net39 _444_/a_448_472# 0.002089f
C14834 _132_ FILLER_0_18_107/a_1468_375# 0.089207f
C14835 net16 _444_/a_2665_112# 0.011295f
C14836 _321_/a_3662_472# vdd 0.001229f
C14837 cal_count\[2\] net47 0.274891f
C14838 FILLER_0_7_233/a_36_472# FILLER_0_6_231/a_124_375# 0.001684f
C14839 FILLER_0_11_142/a_484_472# net23 0.006988f
C14840 FILLER_0_14_91/a_484_472# FILLER_0_14_99/a_36_472# 0.013276f
C14841 FILLER_0_4_107/a_1380_472# vdd 0.007022f
C14842 FILLER_0_2_171/a_36_472# net59 0.066486f
C14843 FILLER_0_8_24/a_36_472# net47 0.097212f
C14844 net67 _450_/a_1040_527# 0.032098f
C14845 FILLER_0_12_20/a_572_375# vss 0.054934f
C14846 FILLER_0_12_20/a_36_472# vdd 0.068477f
C14847 net78 net77 0.252376f
C14848 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_36_472# 0.026657f
C14849 FILLER_0_18_2/a_1828_472# _452_/a_448_472# 0.005748f
C14850 _435_/a_1204_472# vdd 0.013805f
C14851 FILLER_0_4_152/a_124_375# FILLER_0_5_148/a_572_375# 0.05841f
C14852 _057_ _058_ 0.098076f
C14853 FILLER_0_19_55/a_124_375# FILLER_0_18_53/a_484_472# 0.001684f
C14854 _013_ _424_/a_2248_156# 0.001828f
C14855 FILLER_0_9_72/a_932_472# _439_/a_36_151# 0.001723f
C14856 FILLER_0_16_107/a_36_472# _136_ 0.011469f
C14857 FILLER_0_11_64/a_36_472# cal_count\[3\] 0.0081f
C14858 vss FILLER_0_6_231/a_124_375# 0.00353f
C14859 vdd FILLER_0_6_231/a_572_375# 0.018694f
C14860 ctlp[2] _422_/a_2248_156# 0.001328f
C14861 _098_ _048_ 0.092201f
C14862 _411_/a_36_151# FILLER_0_0_232/a_36_472# 0.001723f
C14863 _093_ _302_/a_224_472# 0.011376f
C14864 fanout53/a_36_160# _137_ 0.001852f
C14865 _122_ FILLER_0_5_172/a_124_375# 0.001352f
C14866 net57 _136_ 0.168299f
C14867 _415_/a_36_151# FILLER_0_8_263/a_124_375# 0.001619f
C14868 FILLER_0_7_195/a_124_375# vss 0.006314f
C14869 _158_ _157_ 0.001663f
C14870 FILLER_0_4_197/a_1380_472# _081_ 0.001345f
C14871 _128_ _122_ 0.019207f
C14872 FILLER_0_19_171/a_1380_472# _434_/a_36_151# 0.00271f
C14873 _451_/a_836_156# _040_ 0.016371f
C14874 net63 FILLER_0_18_177/a_2276_472# 0.012025f
C14875 _030_ _168_ 0.015729f
C14876 ctln[1] net8 0.678616f
C14877 _394_/a_56_524# vdd 0.010692f
C14878 _394_/a_728_93# vss 0.024106f
C14879 _408_/a_728_93# _450_/a_2225_156# 0.00128f
C14880 result[5] net77 0.142532f
C14881 FILLER_0_20_193/a_36_472# FILLER_0_18_177/a_1916_375# 0.0027f
C14882 fanout55/a_36_160# FILLER_0_13_80/a_124_375# 0.00805f
C14883 _036_ _384_/a_224_472# 0.001921f
C14884 net26 FILLER_0_23_44/a_36_472# 0.013977f
C14885 FILLER_0_2_165/a_36_472# net59 0.067972f
C14886 net82 _066_ 0.029681f
C14887 mask\[4\] _293_/a_36_472# 0.023203f
C14888 _044_ _416_/a_2248_156# 0.005198f
C14889 FILLER_0_19_28/a_572_375# vdd 0.034691f
C14890 cal_count\[3\] _055_ 0.039546f
C14891 FILLER_0_18_177/a_3260_375# _202_/a_36_160# 0.001948f
C14892 _050_ FILLER_0_22_128/a_572_375# 0.002607f
C14893 net57 _070_ 0.202843f
C14894 FILLER_0_10_256/a_36_472# net28 0.00136f
C14895 _098_ FILLER_0_21_150/a_124_375# 0.006526f
C14896 net25 FILLER_0_23_60/a_124_375# 0.004431f
C14897 _276_/a_36_160# FILLER_0_18_209/a_572_375# 0.004736f
C14898 FILLER_0_15_2/a_572_375# vss 0.055203f
C14899 FILLER_0_15_2/a_36_472# vdd 0.104741f
C14900 mask\[0\] FILLER_0_14_181/a_36_472# 0.001234f
C14901 output23/a_224_472# FILLER_0_24_130/a_36_472# 0.001994f
C14902 ctln[6] net59 0.001267f
C14903 _428_/a_2665_112# state\[2\] 0.001746f
C14904 _008_ output31/a_224_472# 0.051074f
C14905 FILLER_0_21_28/a_1828_472# _424_/a_36_151# 0.001723f
C14906 trim_val\[2\] net40 0.06019f
C14907 _216_/a_67_603# mask\[9\] 0.003086f
C14908 _157_ net14 0.026868f
C14909 _144_ FILLER_0_21_125/a_124_375# 0.009117f
C14910 _073_ cal_itt\[1\] 0.058541f
C14911 _098_ net71 1.076897f
C14912 net64 FILLER_0_9_270/a_124_375# 0.013532f
C14913 _069_ _068_ 0.003779f
C14914 net41 _402_/a_718_527# 0.019628f
C14915 _267_/a_36_472# _090_ 0.001109f
C14916 FILLER_0_13_80/a_36_472# vss 0.009445f
C14917 net38 _445_/a_36_151# 0.112205f
C14918 net16 _160_ 0.354736f
C14919 _016_ _428_/a_448_472# 0.00347f
C14920 net81 FILLER_0_15_235/a_572_375# 0.009675f
C14921 _105_ _295_/a_36_472# 0.031356f
C14922 _195_/a_67_603# mask\[2\] 0.003161f
C14923 net82 FILLER_0_3_172/a_1828_472# 0.004472f
C14924 _079_ fanout75/a_36_113# 0.059598f
C14925 FILLER_0_15_116/a_36_472# _136_ 0.003818f
C14926 _128_ _061_ 0.76584f
C14927 _432_/a_2665_112# _091_ 0.002978f
C14928 FILLER_0_10_78/a_572_375# FILLER_0_9_72/a_1380_472# 0.001543f
C14929 net75 FILLER_0_6_231/a_572_375# 0.002577f
C14930 FILLER_0_4_107/a_36_472# _369_/a_36_68# 0.001709f
C14931 net46 vdd 0.255965f
C14932 net18 _418_/a_796_472# 0.003044f
C14933 _094_ net19 0.06304f
C14934 FILLER_0_17_142/a_484_472# vss 0.030872f
C14935 FILLER_0_5_54/a_572_375# _440_/a_36_151# 0.026916f
C14936 output45/a_224_472# output17/a_224_472# 0.071473f
C14937 fanout66/a_36_113# _164_ 0.010496f
C14938 net82 net37 0.037195f
C14939 net18 _419_/a_2560_156# 0.008155f
C14940 _360_/a_36_160# net47 0.011731f
C14941 _053_ _312_/a_672_472# 0.001065f
C14942 mask\[2\] net30 0.089173f
C14943 output19/a_224_472# vdd 0.063651f
C14944 FILLER_0_13_65/a_36_472# _449_/a_36_151# 0.001723f
C14945 FILLER_0_21_206/a_124_375# net33 0.001579f
C14946 _086_ _375_/a_692_497# 0.002565f
C14947 _073_ vss 0.216342f
C14948 net55 FILLER_0_21_60/a_36_472# 0.06794f
C14949 _052_ FILLER_0_18_61/a_124_375# 0.006877f
C14950 _411_/a_1204_472# ctln[3] 0.00185f
C14951 FILLER_0_18_76/a_36_472# vss 0.007456f
C14952 FILLER_0_15_150/a_124_375# _427_/a_2248_156# 0.001221f
C14953 net52 _440_/a_1308_423# 0.047012f
C14954 net81 _425_/a_2560_156# 0.022037f
C14955 _410_/a_36_68# vdd 0.039824f
C14956 comp net17 0.02802f
C14957 _321_/a_170_472# _395_/a_36_488# 0.007047f
C14958 _429_/a_2560_156# vss 0.005255f
C14959 net62 _429_/a_2248_156# 0.012262f
C14960 trim_mask\[1\] FILLER_0_4_91/a_36_472# 0.26171f
C14961 net72 _394_/a_56_524# 0.066156f
C14962 _423_/a_2248_156# vss 0.010039f
C14963 _423_/a_2665_112# vdd 0.022696f
C14964 FILLER_0_23_282/a_124_375# FILLER_0_23_274/a_124_375# 0.003732f
C14965 FILLER_0_19_155/a_124_375# _145_ 0.006057f
C14966 net41 output38/a_224_472# 0.017358f
C14967 FILLER_0_4_152/a_124_375# net23 0.039975f
C14968 _104_ _420_/a_2248_156# 0.027923f
C14969 net72 FILLER_0_19_28/a_572_375# 0.010026f
C14970 _443_/a_2665_112# trim_mask\[4\] 0.013708f
C14971 net76 _083_ 0.002446f
C14972 net41 FILLER_0_21_28/a_572_375# 0.054443f
C14973 FILLER_0_20_169/a_124_375# vdd 0.03036f
C14974 _126_ state\[2\] 0.030985f
C14975 net35 _214_/a_36_160# 0.0116f
C14976 fanout53/a_36_160# net56 0.196684f
C14977 net47 _450_/a_1353_112# 0.018879f
C14978 net15 _453_/a_36_151# 0.009841f
C14979 _013_ FILLER_0_17_56/a_36_472# 0.002659f
C14980 FILLER_0_22_128/a_1828_472# vdd 0.005724f
C14981 FILLER_0_22_128/a_1380_472# vss 0.007305f
C14982 net64 net18 1.557441f
C14983 _017_ _043_ 0.02569f
C14984 net32 _421_/a_1000_472# 0.002275f
C14985 _422_/a_1000_472# _109_ 0.003473f
C14986 _070_ FILLER_0_10_107/a_572_375# 0.003959f
C14987 result[6] _420_/a_2248_156# 0.003418f
C14988 output8/a_224_472# vdd 0.023187f
C14989 net66 vss 0.265973f
C14990 net15 net69 0.034091f
C14991 _086_ _267_/a_1120_472# 0.004245f
C14992 _442_/a_1000_472# vdd 0.003088f
C14993 net80 FILLER_0_16_154/a_1468_375# 0.013593f
C14994 _452_/a_448_472# _041_ 0.007f
C14995 _155_ _156_ 0.037229f
C14996 _053_ FILLER_0_6_47/a_932_472# 0.011457f
C14997 _183_ FILLER_0_18_53/a_124_375# 0.001032f
C14998 FILLER_0_18_2/a_3260_375# vdd 0.046682f
C14999 _343_/a_49_472# _093_ 0.001926f
C15000 output20/a_224_472# vss -0.004787f
C15001 trim_mask\[1\] vdd 0.241393f
C15002 output9/a_224_472# cal_itt\[0\] 0.008307f
C15003 output28/a_224_472# net28 0.048681f
C15004 _432_/a_1308_423# _137_ 0.002078f
C15005 _445_/a_2248_156# net17 0.06175f
C15006 FILLER_0_7_72/a_3172_472# net14 0.046751f
C15007 _428_/a_1000_472# net74 0.00735f
C15008 FILLER_0_15_116/a_484_472# net53 0.002804f
C15009 cal_itt\[2\] cal_itt\[1\] 0.057194f
C15010 mask\[5\] FILLER_0_18_177/a_2364_375# 0.002726f
C15011 fanout71/a_36_113# _098_ 0.012725f
C15012 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001597f
C15013 FILLER_0_15_282/a_36_472# _417_/a_1308_423# 0.001295f
C15014 mask\[5\] _339_/a_36_160# 0.007734f
C15015 net55 FILLER_0_18_76/a_124_375# 0.001706f
C15016 cal_itt\[3\] _074_ 0.584958f
C15017 _288_/a_224_472# _006_ 0.001278f
C15018 net1 cal_itt\[1\] 0.229522f
C15019 _425_/a_36_151# vss 0.00158f
C15020 fanout82/a_36_113# vdd 0.083174f
C15021 _425_/a_448_472# vdd 0.029071f
C15022 _072_ _375_/a_1612_497# 0.002646f
C15023 FILLER_0_18_2/a_2812_375# net55 0.007169f
C15024 net20 FILLER_0_12_220/a_124_375# 0.003161f
C15025 _021_ net57 0.00736f
C15026 FILLER_0_9_282/a_572_375# vdd 0.002928f
C15027 FILLER_0_9_282/a_124_375# vss 0.00451f
C15028 _091_ FILLER_0_18_177/a_932_472# 0.002113f
C15029 net23 _145_ 0.035734f
C15030 vss _167_ 0.043544f
C15031 _074_ _081_ 0.070546f
C15032 mask\[7\] _435_/a_1000_472# 0.024725f
C15033 _378_/a_224_472# _165_ 0.00481f
C15034 result[6] _421_/a_2560_156# 0.006943f
C15035 _091_ _140_ 0.006511f
C15036 FILLER_0_5_128/a_124_375# _160_ 0.001157f
C15037 vdd FILLER_0_22_107/a_36_472# 0.114332f
C15038 vss FILLER_0_22_107/a_572_375# 0.001944f
C15039 FILLER_0_15_212/a_1468_375# mask\[1\] 0.045287f
C15040 _412_/a_36_151# cal_itt\[1\] 0.025078f
C15041 _444_/a_448_472# net42 0.002526f
C15042 cal_count\[3\] _278_/a_36_160# 0.008398f
C15043 _050_ _436_/a_448_472# 0.064832f
C15044 _223_/a_36_160# vdd 0.018653f
C15045 _067_ vss 0.20904f
C15046 net63 _093_ 0.109689f
C15047 _176_ FILLER_0_17_72/a_1828_472# 0.001028f
C15048 FILLER_0_16_57/a_572_375# _131_ 0.015859f
C15049 cal_itt\[2\] vss 0.249871f
C15050 net41 vdd 1.983262f
C15051 output8/a_224_472# net75 0.044765f
C15052 fanout78/a_36_113# _094_ 0.01312f
C15053 FILLER_0_17_282/a_36_472# net30 0.001189f
C15054 FILLER_0_17_64/a_124_375# FILLER_0_17_56/a_572_375# 0.012001f
C15055 fanout56/a_36_113# net36 0.021321f
C15056 FILLER_0_4_177/a_36_472# net22 0.006506f
C15057 FILLER_0_4_197/a_1380_472# FILLER_0_4_213/a_36_472# 0.013277f
C15058 net19 FILLER_0_23_274/a_36_472# 0.075097f
C15059 FILLER_0_15_72/a_36_472# cal_count\[1\] 0.006408f
C15060 _259_/a_271_68# net4 0.003663f
C15061 net55 _424_/a_2560_156# 0.003707f
C15062 _078_ _080_ 0.030094f
C15063 net4 FILLER_0_6_231/a_124_375# 0.002212f
C15064 _001_ _082_ 0.46787f
C15065 net1 vss 0.161208f
C15066 _299_/a_36_472# vdd 0.098451f
C15067 FILLER_0_4_107/a_484_472# _154_ 0.040595f
C15068 output31/a_224_472# _006_ 0.090006f
C15069 state\[0\] _072_ 0.030642f
C15070 _341_/a_665_69# _141_ 0.001064f
C15071 FILLER_0_14_99/a_36_472# vdd 0.095251f
C15072 FILLER_0_14_99/a_124_375# vss 0.017196f
C15073 _253_/a_36_68# vdd 0.016219f
C15074 _090_ _113_ 0.263235f
C15075 net54 vss 0.715177f
C15076 FILLER_0_20_15/a_1468_375# vss 0.055156f
C15077 FILLER_0_20_15/a_36_472# vdd 0.086947f
C15078 _411_/a_2560_156# net8 0.013106f
C15079 FILLER_0_18_107/a_1020_375# FILLER_0_19_111/a_572_375# 0.05841f
C15080 _232_/a_255_603# net47 0.001241f
C15081 _412_/a_36_151# vss 0.003515f
C15082 net17 FILLER_0_20_15/a_1380_472# 0.012286f
C15083 FILLER_0_15_72/a_572_375# _451_/a_3129_107# 0.007026f
C15084 _092_ output18/a_224_472# 0.002205f
C15085 _168_ trim_mask\[3\] 0.007154f
C15086 _086_ _074_ 0.186795f
C15087 net58 net8 0.175026f
C15088 net75 _425_/a_448_472# 0.038993f
C15089 _077_ _131_ 0.03465f
C15090 net27 net19 0.036883f
C15091 net63 output35/a_224_472# 0.148302f
C15092 _102_ _099_ 0.151018f
C15093 FILLER_0_4_177/a_572_375# _087_ 0.006527f
C15094 net79 _416_/a_448_472# 0.078357f
C15095 FILLER_0_20_107/a_36_472# net14 0.002543f
C15096 _322_/a_124_24# _070_ 0.033355f
C15097 _119_ _074_ 0.153267f
C15098 _091_ _128_ 0.003717f
C15099 _116_ FILLER_0_13_206/a_124_375# 0.003926f
C15100 mask\[9\] FILLER_0_20_98/a_124_375# 0.003444f
C15101 _404_/a_36_472# _182_ 0.036415f
C15102 cal_count\[2\] _402_/a_718_527# 0.004645f
C15103 net20 net30 0.033149f
C15104 ctlp[7] _436_/a_36_151# 0.002655f
C15105 fanout80/a_36_113# vss 0.003526f
C15106 _448_/a_2665_112# _170_ 0.002715f
C15107 _448_/a_1204_472# _037_ 0.008883f
C15108 _444_/a_1000_472# net40 0.038229f
C15109 _265_/a_244_68# _001_ 0.008874f
C15110 FILLER_0_17_226/a_36_472# net63 0.001822f
C15111 FILLER_0_20_193/a_572_375# vss 0.005887f
C15112 FILLER_0_20_193/a_36_472# vdd 0.091886f
C15113 output12/a_224_472# net12 0.007193f
C15114 _118_ _090_ 0.005469f
C15115 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_484_472# 0.013276f
C15116 net21 _434_/a_2665_112# 0.004945f
C15117 net41 net72 0.319547f
C15118 _398_/a_36_113# vdd 0.030449f
C15119 FILLER_0_15_72/a_124_375# FILLER_0_13_72/a_36_472# 0.001418f
C15120 net75 _253_/a_36_68# 0.047906f
C15121 FILLER_0_9_105/a_36_472# vss 0.002744f
C15122 FILLER_0_9_105/a_484_472# vdd 0.03152f
C15123 _441_/a_796_472# _030_ 0.024278f
C15124 trim_mask\[2\] net66 0.036211f
C15125 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_572_375# 0.026339f
C15126 _032_ FILLER_0_2_127/a_124_375# 0.002221f
C15127 _013_ _131_ 0.001178f
C15128 fanout53/a_36_160# _095_ 0.007436f
C15129 _321_/a_170_472# _125_ 0.008492f
C15130 FILLER_0_5_198/a_572_375# net59 0.00183f
C15131 _112_ _001_ 0.002527f
C15132 _004_ FILLER_0_10_256/a_124_375# 0.006989f
C15133 output21/a_224_472# output35/a_224_472# 0.001374f
C15134 FILLER_0_12_2/a_484_472# net67 0.006435f
C15135 _036_ _441_/a_36_151# 0.005754f
C15136 FILLER_0_18_139/a_932_472# vdd 0.002904f
C15137 FILLER_0_18_139/a_484_472# vss 0.006719f
C15138 net60 net77 0.046792f
C15139 _073_ net4 0.076114f
C15140 _009_ FILLER_0_23_274/a_36_472# 0.005531f
C15141 _292_/a_36_160# _205_/a_36_160# 0.105676f
C15142 mask\[5\] FILLER_0_19_187/a_124_375# 0.007169f
C15143 net49 _440_/a_2248_156# 0.025137f
C15144 _410_/a_36_68# cal_count\[0\] 0.007618f
C15145 _187_ _039_ 0.228074f
C15146 _142_ net73 0.090025f
C15147 net64 FILLER_0_15_235/a_572_375# 0.007219f
C15148 FILLER_0_16_154/a_1020_375# vdd 0.004279f
C15149 FILLER_0_16_154/a_572_375# vss 0.003976f
C15150 _121_ vss 0.082882f
C15151 FILLER_0_18_2/a_1020_375# output44/a_224_472# 0.032639f
C15152 _411_/a_796_472# vss 0.00159f
C15153 _322_/a_848_380# FILLER_0_9_142/a_124_375# 0.001721f
C15154 _431_/a_36_151# FILLER_0_18_107/a_1828_472# 0.001221f
C15155 FILLER_0_7_195/a_36_472# vdd 0.04565f
C15156 _103_ _046_ 0.010317f
C15157 trim_mask\[4\] net69 0.185121f
C15158 net62 _100_ 0.006742f
C15159 FILLER_0_15_235/a_572_375# mask\[1\] 0.013718f
C15160 _326_/a_36_160# _322_/a_124_24# 0.004397f
C15161 FILLER_0_11_109/a_124_375# FILLER_0_10_107/a_484_472# 0.001684f
C15162 mask\[7\] FILLER_0_22_128/a_1380_472# 0.015814f
C15163 _105_ ctlp[2] 0.223601f
C15164 _432_/a_36_151# _093_ 0.018324f
C15165 net75 FILLER_0_8_247/a_124_375# 0.002085f
C15166 _198_/a_67_603# _099_ 0.0109f
C15167 output37/a_224_472# fanout64/a_36_160# 0.017421f
C15168 _004_ net62 0.001201f
C15169 _116_ _311_/a_66_473# 0.001527f
C15170 FILLER_0_10_78/a_1020_375# _120_ 0.003403f
C15171 net32 ctlp[1] 0.032275f
C15172 _087_ net22 0.028009f
C15173 FILLER_0_7_104/a_572_375# vdd 0.038253f
C15174 net63 FILLER_0_19_195/a_36_472# 0.030832f
C15175 trim_mask\[2\] _167_ 0.027204f
C15176 net34 _350_/a_49_472# 0.008001f
C15177 net73 FILLER_0_18_107/a_2812_375# 0.018753f
C15178 FILLER_0_7_72/a_1380_472# net52 0.003507f
C15179 _110_ _098_ 0.09704f
C15180 output20/a_224_472# mask\[7\] 0.024731f
C15181 net82 _122_ 0.001375f
C15182 net41 _424_/a_36_151# 0.00413f
C15183 _426_/a_2248_156# _076_ 0.015189f
C15184 FILLER_0_18_107/a_1468_375# vdd 0.004726f
C15185 FILLER_0_10_78/a_572_375# _176_ 0.005927f
C15186 output34/a_224_472# _093_ 0.012298f
C15187 _402_/a_56_567# net47 0.026503f
C15188 _196_/a_36_160# _045_ 0.036714f
C15189 trim_mask\[1\] FILLER_0_6_47/a_3172_472# 0.004605f
C15190 net39 _445_/a_2248_156# 0.003571f
C15191 net52 FILLER_0_9_72/a_572_375# 0.022582f
C15192 _164_ vdd 0.711488f
C15193 _049_ FILLER_0_22_128/a_3260_375# 0.16381f
C15194 net54 FILLER_0_22_128/a_1020_375# 0.010068f
C15195 FILLER_0_18_37/a_1020_375# vdd 0.020683f
C15196 net24 _050_ 0.049889f
C15197 FILLER_0_16_89/a_124_375# vdd 0.01011f
C15198 _086_ _124_ 0.063099f
C15199 _283_/a_36_472# _099_ 0.004667f
C15200 FILLER_0_11_64/a_36_472# _120_ 0.011673f
C15201 _446_/a_2560_156# vdd 0.003959f
C15202 _446_/a_2665_112# vss 0.001781f
C15203 _421_/a_2665_112# _419_/a_2665_112# 0.002588f
C15204 FILLER_0_24_274/a_1020_375# vss 0.003553f
C15205 net52 cal_count\[3\] 0.348542f
C15206 state\[2\] FILLER_0_13_142/a_932_472# 0.004118f
C15207 _159_ net47 0.01358f
C15208 FILLER_0_5_72/a_932_472# vss 0.003084f
C15209 FILLER_0_5_72/a_1380_472# vdd 0.001438f
C15210 output14/a_224_472# _442_/a_2665_112# 0.009771f
C15211 FILLER_0_4_144/a_36_472# _081_ 0.003547f
C15212 fanout70/a_36_113# _136_ 0.002788f
C15213 _063_ _444_/a_2665_112# 0.001996f
C15214 _390_/a_36_68# vdd 0.012472f
C15215 mask\[3\] FILLER_0_17_218/a_124_375# 0.016168f
C15216 _068_ net22 0.088209f
C15217 result[6] _419_/a_2665_112# 0.001225f
C15218 _148_ FILLER_0_22_107/a_572_375# 0.00652f
C15219 FILLER_0_20_107/a_36_472# _098_ 0.011046f
C15220 FILLER_0_10_28/a_124_375# net51 0.00979f
C15221 fanout69/a_36_113# net69 0.040451f
C15222 net15 _095_ 0.056214f
C15223 result[8] _422_/a_448_472# 0.002989f
C15224 FILLER_0_16_73/a_572_375# _175_ 0.138524f
C15225 _408_/a_718_524# vdd 0.002635f
C15226 _289_/a_36_472# net30 0.009623f
C15227 _413_/a_36_151# FILLER_0_3_172/a_1916_375# 0.059049f
C15228 FILLER_0_2_93/a_484_472# net69 0.0127f
C15229 _443_/a_2665_112# _066_ 0.001654f
C15230 _131_ _179_ 0.034602f
C15231 _088_ net21 0.053843f
C15232 net41 cal_count\[0\] 0.001014f
C15233 FILLER_0_16_73/a_36_472# net15 0.005297f
C15234 cal_itt\[2\] net4 0.333682f
C15235 net54 mask\[7\] 0.262465f
C15236 mask\[5\] vss 0.528441f
C15237 _076_ _118_ 0.06281f
C15238 cal_count\[2\] vdd 0.932907f
C15239 _176_ _451_/a_2449_156# 0.038547f
C15240 net64 FILLER_0_8_247/a_1380_472# 0.001021f
C15241 FILLER_0_18_209/a_572_375# vss 0.007545f
C15242 FILLER_0_18_209/a_36_472# vdd 0.089327f
C15243 net1 net4 0.03357f
C15244 FILLER_0_8_24/a_572_375# vss 0.012859f
C15245 FILLER_0_8_24/a_36_472# vdd 0.007423f
C15246 net54 _148_ 0.098648f
C15247 _091_ FILLER_0_13_228/a_124_375# 0.001657f
C15248 FILLER_0_18_107/a_484_472# mask\[9\] 0.001955f
C15249 FILLER_0_15_150/a_36_472# net53 0.016925f
C15250 FILLER_0_3_78/a_124_375# _160_ 0.003276f
C15251 net65 fanout76/a_36_160# 0.018025f
C15252 FILLER_0_19_47/a_572_375# _183_ 0.001186f
C15253 net19 FILLER_0_14_263/a_124_375# 0.032085f
C15254 FILLER_0_12_220/a_572_375# vdd -0.014642f
C15255 FILLER_0_12_220/a_124_375# vss 0.040895f
C15256 _415_/a_448_472# result[1] 0.005209f
C15257 _311_/a_66_473# _117_ 0.001055f
C15258 _103_ net18 0.11279f
C15259 FILLER_0_18_139/a_1468_375# net23 0.04546f
C15260 FILLER_0_2_101/a_124_375# _160_ 0.001047f
C15261 FILLER_0_4_107/a_1020_375# _160_ 0.015684f
C15262 _426_/a_1000_472# net64 0.008796f
C15263 net26 vss 0.263774f
C15264 result[7] _420_/a_2248_156# 0.034866f
C15265 net15 FILLER_0_17_72/a_484_472# 0.002925f
C15266 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_124_375# 0.026339f
C15267 _431_/a_2665_112# FILLER_0_15_150/a_36_472# 0.035266f
C15268 FILLER_0_8_37/a_124_375# vdd 0.029725f
C15269 net47 FILLER_0_4_91/a_124_375# 0.009482f
C15270 FILLER_0_11_124/a_36_472# vdd 0.005222f
C15271 FILLER_0_11_124/a_124_375# vss 0.017354f
C15272 _096_ _043_ 0.842762f
C15273 net32 _204_/a_67_603# 0.037639f
C15274 output29/a_224_472# _416_/a_448_472# 0.008149f
C15275 _053_ _163_ 0.763235f
C15276 FILLER_0_8_247/a_36_472# _316_/a_124_24# 0.001386f
C15277 _313_/a_67_603# _120_ 0.005873f
C15278 output23/a_224_472# FILLER_0_22_128/a_2364_375# 0.002439f
C15279 net7 ctln[9] 0.005103f
C15280 output12/a_224_472# _413_/a_448_472# 0.001495f
C15281 _186_ _095_ 0.042856f
C15282 _028_ net51 0.002321f
C15283 output18/a_224_472# vdd -0.01545f
C15284 _063_ _160_ 0.091185f
C15285 _449_/a_2248_156# _038_ 0.016483f
C15286 net80 FILLER_0_22_177/a_124_375# 0.013214f
C15287 FILLER_0_16_57/a_1380_472# _176_ 0.01346f
C15288 _136_ mask\[9\] 0.015204f
C15289 FILLER_0_18_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001684f
C15290 _091_ _139_ 0.05535f
C15291 net65 FILLER_0_1_212/a_36_472# 0.004414f
C15292 _141_ FILLER_0_17_142/a_484_472# 0.004527f
C15293 FILLER_0_7_59/a_572_375# net68 0.005738f
C15294 _069_ _314_/a_224_472# 0.003461f
C15295 _436_/a_36_151# FILLER_0_22_107/a_484_472# 0.001723f
C15296 net65 FILLER_0_2_177/a_484_472# 0.01675f
C15297 output42/a_224_472# _221_/a_36_160# 0.017421f
C15298 FILLER_0_5_88/a_36_472# _163_ 0.006541f
C15299 FILLER_0_17_200/a_36_472# FILLER_0_18_177/a_2724_472# 0.026657f
C15300 FILLER_0_7_72/a_2812_375# _053_ 0.016329f
C15301 net72 cal_count\[2\] 0.073818f
C15302 FILLER_0_5_54/a_1380_472# vss 0.007301f
C15303 FILLER_0_8_107/a_124_375# FILLER_0_10_107/a_36_472# 0.0027f
C15304 cal_count\[2\] _452_/a_1040_527# 0.002003f
C15305 _430_/a_1204_472# _091_ 0.007301f
C15306 net52 FILLER_0_3_78/a_484_472# 0.003143f
C15307 _076_ _068_ 0.35956f
C15308 _195_/a_67_603# vss 0.002638f
C15309 _437_/a_36_151# vdd 0.115376f
C15310 FILLER_0_10_28/a_124_375# net6 0.007948f
C15311 cal_count\[3\] _172_ 0.03048f
C15312 _356_/a_36_472# mask\[9\] 0.047632f
C15313 _444_/a_36_151# net49 0.007102f
C15314 _430_/a_796_472# mask\[2\] 0.006305f
C15315 net15 _440_/a_448_472# 0.036624f
C15316 net54 _436_/a_1308_423# 0.002665f
C15317 net46 output46/a_224_472# 0.008691f
C15318 _074_ _161_ 0.191658f
C15319 vss net30 0.17209f
C15320 _360_/a_36_160# vdd 0.006439f
C15321 _440_/a_2560_156# _164_ 0.003934f
C15322 FILLER_0_4_197/a_36_472# vdd 0.042721f
C15323 FILLER_0_1_212/a_36_472# net59 0.002567f
C15324 _242_/a_36_160# FILLER_0_5_148/a_572_375# 0.00805f
C15325 _119_ _312_/a_672_472# 0.00145f
C15326 _112_ _316_/a_124_24# 0.032665f
C15327 _088_ FILLER_0_4_213/a_484_472# 0.018066f
C15328 result[9] result[2] 0.001669f
C15329 _151_ _365_/a_36_68# 0.001944f
C15330 net41 _407_/a_36_472# 0.003257f
C15331 _158_ _160_ 0.018681f
C15332 net54 _433_/a_448_472# 0.008777f
C15333 fanout54/a_36_160# _433_/a_2248_156# 0.012122f
C15334 _058_ _120_ 0.008566f
C15335 FILLER_0_23_44/a_572_375# vdd -0.011314f
C15336 FILLER_0_2_177/a_484_472# net59 0.007829f
C15337 _077_ _453_/a_36_151# 0.042928f
C15338 FILLER_0_10_28/a_36_472# net40 0.020589f
C15339 FILLER_0_16_107/a_124_375# FILLER_0_18_107/a_36_472# 0.001512f
C15340 _177_ vdd 0.111636f
C15341 _315_/a_36_68# _120_ 0.00572f
C15342 net17 FILLER_0_23_44/a_36_472# 0.071244f
C15343 state\[2\] _095_ 0.001426f
C15344 FILLER_0_12_124/a_36_472# cal_count\[3\] 0.004109f
C15345 FILLER_0_21_142/a_36_472# net35 0.003079f
C15346 fanout55/a_36_160# _043_ 0.019538f
C15347 _176_ _182_ 0.008217f
C15348 _091_ _429_/a_1000_472# 0.029742f
C15349 FILLER_0_20_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001543f
C15350 FILLER_0_19_47/a_124_375# FILLER_0_18_37/a_1380_472# 0.001684f
C15351 FILLER_0_4_197/a_572_375# net22 0.016547f
C15352 _164_ FILLER_0_6_47/a_3172_472# 0.001058f
C15353 net15 ctln[9] 0.01475f
C15354 _321_/a_170_472# _069_ 0.025551f
C15355 net15 mask\[8\] 0.02403f
C15356 net63 FILLER_0_20_193/a_124_375# 0.075841f
C15357 FILLER_0_17_38/a_484_472# vdd 0.009211f
C15358 trim_val\[0\] FILLER_0_6_47/a_484_472# 0.001215f
C15359 vss _450_/a_448_472# -0.001661f
C15360 _098_ _433_/a_1204_472# 0.014374f
C15361 net14 _160_ 0.034023f
C15362 _178_ _180_ 0.004668f
C15363 output7/a_224_472# net17 0.001164f
C15364 _313_/a_67_603# _227_/a_36_160# 0.032438f
C15365 _125_ _135_ 0.001926f
C15366 net47 _452_/a_448_472# 0.005335f
C15367 net41 _444_/a_1308_423# 0.015841f
C15368 net26 _424_/a_448_472# 0.063966f
C15369 FILLER_0_4_144/a_124_375# trim_mask\[4\] 0.014395f
C15370 net31 net29 0.009564f
C15371 _274_/a_1612_497# net20 0.002057f
C15372 _075_ net59 0.01129f
C15373 net54 FILLER_0_19_134/a_36_472# 0.061344f
C15374 _448_/a_2560_156# net22 0.00766f
C15375 _064_ _034_ 1.397143f
C15376 FILLER_0_13_65/a_36_472# vss 0.007545f
C15377 _322_/a_848_380# _127_ 0.018892f
C15378 _015_ FILLER_0_10_247/a_124_375# 0.001261f
C15379 _058_ FILLER_0_9_105/a_572_375# 0.003832f
C15380 net48 _001_ 0.006122f
C15381 _028_ _163_ 0.199021f
C15382 FILLER_0_21_28/a_3260_375# _012_ 0.016427f
C15383 net35 net21 0.001845f
C15384 _093_ FILLER_0_18_61/a_124_375# 0.031062f
C15385 trimb[1] net38 0.161478f
C15386 net15 net74 0.05717f
C15387 ctlp[4] vss 0.102044f
C15388 mask\[5\] mask\[7\] 0.014384f
C15389 FILLER_0_5_164/a_36_472# _163_ 0.001777f
C15390 _422_/a_2665_112# net19 0.006987f
C15391 _093_ FILLER_0_17_104/a_1020_375# 0.01418f
C15392 _438_/a_2665_112# FILLER_0_19_111/a_124_375# 0.006271f
C15393 _372_/a_170_472# _122_ 0.018399f
C15394 _129_ calibrate 0.04134f
C15395 _255_/a_224_552# _118_ 0.002405f
C15396 _114_ _116_ 0.038641f
C15397 net15 cal_count\[1\] 0.089855f
C15398 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001597f
C15399 net55 FILLER_0_17_38/a_124_375# 0.003236f
C15400 net72 FILLER_0_17_38/a_484_472# 0.00547f
C15401 FILLER_0_5_128/a_572_375# _081_ 0.023853f
C15402 net23 _242_/a_36_160# 0.007466f
C15403 FILLER_0_24_63/a_36_472# vdd 0.055524f
C15404 _233_/a_36_160# FILLER_0_6_37/a_36_472# 0.012692f
C15405 _162_ _062_ 0.033583f
C15406 net33 _107_ 0.001322f
C15407 _258_/a_36_160# _081_ 0.00776f
C15408 FILLER_0_7_72/a_2812_375# _028_ 0.003873f
C15409 net4 FILLER_0_12_220/a_124_375# 0.016485f
C15410 net73 fanout73/a_36_113# 0.02062f
C15411 net20 _277_/a_36_160# 0.015569f
C15412 FILLER_0_3_221/a_124_375# vdd 0.008869f
C15413 trim_mask\[1\] FILLER_0_6_90/a_484_472# 0.014443f
C15414 _058_ _227_/a_36_160# 0.008511f
C15415 mask\[4\] FILLER_0_18_177/a_1380_472# 0.016924f
C15416 net19 _001_ 0.018424f
C15417 _261_/a_36_160# FILLER_0_5_148/a_124_375# 0.005705f
C15418 _412_/a_2665_112# net5 0.042084f
C15419 FILLER_0_20_177/a_1380_472# vdd 0.009871f
C15420 FILLER_0_20_177/a_932_472# vss 0.001272f
C15421 FILLER_0_18_100/a_124_375# _438_/a_2248_156# 0.001068f
C15422 net28 net29 0.178557f
C15423 _440_/a_2248_156# net47 0.017063f
C15424 _119_ FILLER_0_8_156/a_124_375# 0.025304f
C15425 mask\[8\] FILLER_0_22_86/a_1468_375# 0.015339f
C15426 net35 FILLER_0_22_86/a_1020_375# 0.010202f
C15427 net69 _157_ 0.112249f
C15428 net52 _442_/a_1308_423# 0.017208f
C15429 _232_/a_67_603# vss 0.00988f
C15430 FILLER_0_14_263/a_36_472# vss 0.003195f
C15431 net57 _395_/a_36_488# 0.026081f
C15432 FILLER_0_16_89/a_36_472# _451_/a_2449_156# 0.001571f
C15433 _115_ trim_mask\[0\] 0.008966f
C15434 _057_ net21 0.143214f
C15435 _069_ _429_/a_1204_472# 0.025254f
C15436 fanout59/a_36_160# net64 0.006298f
C15437 _183_ _182_ 0.002134f
C15438 net74 _133_ 0.696379f
C15439 _077_ _426_/a_2665_112# 0.001392f
C15440 _429_/a_36_151# _043_ 0.002771f
C15441 net65 _425_/a_2665_112# 0.00628f
C15442 _321_/a_3662_472# _176_ 0.002006f
C15443 state\[0\] vdd 0.120171f
C15444 _186_ cal_count\[1\] 0.003341f
C15445 FILLER_0_18_177/a_1020_375# vdd 0.040478f
C15446 _095_ FILLER_0_14_107/a_932_472# 0.014431f
C15447 _128_ _426_/a_2248_156# 0.019019f
C15448 FILLER_0_13_290/a_36_472# result[3] 0.001069f
C15449 FILLER_0_9_223/a_124_375# _070_ 0.002989f
C15450 FILLER_0_2_101/a_124_375# _156_ 0.022015f
C15451 net44 FILLER_0_15_2/a_36_472# 0.007808f
C15452 net82 FILLER_0_3_212/a_124_375# 0.015932f
C15453 _150_ net14 0.001303f
C15454 ctln[5] _448_/a_1000_472# 0.007584f
C15455 output8/a_224_472# _413_/a_2665_112# 0.010726f
C15456 FILLER_0_10_78/a_484_472# net52 0.004421f
C15457 _192_/a_255_603# mask\[1\] 0.001059f
C15458 result[7] _419_/a_2665_112# 0.002471f
C15459 _131_ FILLER_0_17_56/a_572_375# 0.006224f
C15460 FILLER_0_2_127/a_36_472# vss 0.002567f
C15461 _091_ _098_ 1.501073f
C15462 FILLER_0_7_59/a_36_472# net67 0.021549f
C15463 FILLER_0_7_72/a_2812_375# trim_mask\[0\] 0.005302f
C15464 _128_ _113_ 0.002117f
C15465 FILLER_0_18_2/a_2276_472# net17 0.037088f
C15466 FILLER_0_14_91/a_572_375# vdd -0.011429f
C15467 _255_/a_224_552# _068_ 0.002412f
C15468 _057_ _070_ 0.033401f
C15469 FILLER_0_19_187/a_484_472# _434_/a_2665_112# 0.001868f
C15470 _105_ ctlp[1] 0.158795f
C15471 FILLER_0_5_117/a_36_472# _154_ 0.005034f
C15472 _138_ vss 0.006962f
C15473 vdd FILLER_0_10_94/a_484_472# 0.008627f
C15474 net15 FILLER_0_13_72/a_124_375# 0.006403f
C15475 _422_/a_2665_112# _009_ 0.061508f
C15476 mask\[8\] _437_/a_2665_112# 0.007907f
C15477 _453_/a_1000_472# vss 0.001738f
C15478 _095_ _451_/a_1353_112# 0.00475f
C15479 _348_/a_49_472# vss 0.002301f
C15480 _417_/a_1308_423# _006_ 0.022704f
C15481 _012_ FILLER_0_21_60/a_124_375# 0.016032f
C15482 output9/a_224_472# fanout76/a_36_160# 0.016067f
C15483 FILLER_0_13_212/a_1020_375# FILLER_0_12_220/a_124_375# 0.05841f
C15484 _429_/a_2248_156# FILLER_0_15_212/a_1468_375# 0.001068f
C15485 _091_ FILLER_0_13_212/a_1380_472# 0.003507f
C15486 input1/a_36_113# clk 0.001121f
C15487 result[8] FILLER_0_23_282/a_36_472# 0.001908f
C15488 FILLER_0_9_223/a_572_375# net20 0.03118f
C15489 _104_ net78 0.049954f
C15490 FILLER_0_11_101/a_572_375# cal_count\[3\] 0.002017f
C15491 FILLER_0_20_2/a_124_375# vdd 0.010886f
C15492 _114_ _117_ 0.008886f
C15493 ctln[4] net65 0.020799f
C15494 FILLER_0_5_212/a_124_375# vdd 0.024541f
C15495 _219_/a_36_160# _439_/a_2665_112# 0.002537f
C15496 FILLER_0_18_177/a_2276_472# net21 0.01016f
C15497 FILLER_0_3_2/a_124_375# output41/a_224_472# 0.030009f
C15498 _438_/a_2665_112# vdd 0.00587f
C15499 _438_/a_2248_156# vss 0.002607f
C15500 _274_/a_716_497# net64 0.007904f
C15501 _444_/a_448_472# net67 0.046278f
C15502 _129_ _125_ 0.069221f
C15503 net53 _427_/a_36_151# 0.13192f
C15504 FILLER_0_1_266/a_124_375# vdd -0.002281f
C15505 trim_mask\[1\] FILLER_0_5_88/a_124_375# 0.072632f
C15506 result[9] _420_/a_2665_112# 0.037019f
C15507 net82 _170_ 0.080348f
C15508 _430_/a_36_151# FILLER_0_18_177/a_2724_472# 0.001512f
C15509 FILLER_0_9_60/a_572_375# _439_/a_36_151# 0.001107f
C15510 _077_ _330_/a_224_472# 0.001921f
C15511 net52 _120_ 0.023363f
C15512 net57 calibrate 0.037299f
C15513 state\[2\] net74 0.024462f
C15514 output34/a_224_472# _094_ 0.002719f
C15515 FILLER_0_8_127/a_124_375# _124_ 0.022175f
C15516 FILLER_0_15_282/a_484_472# _006_ 0.00444f
C15517 _151_ _154_ 0.108571f
C15518 result[6] net78 0.027123f
C15519 _128_ _118_ 0.58787f
C15520 _127_ _124_ 0.035569f
C15521 trim[4] vss 0.033925f
C15522 _008_ _418_/a_1308_423# 0.027229f
C15523 fanout61/a_36_113# net78 0.009579f
C15524 _236_/a_36_160# _064_ 0.039922f
C15525 _130_ _131_ 0.005955f
C15526 _402_/a_1296_93# _401_/a_36_68# 0.001523f
C15527 _087_ FILLER_0_5_172/a_124_375# 0.003043f
C15528 net15 FILLER_0_9_72/a_124_375# 0.006492f
C15529 ctln[4] net59 0.10527f
C15530 _143_ _339_/a_36_160# 0.00507f
C15531 trimb[1] net55 0.017528f
C15532 net81 net37 0.18149f
C15533 _340_/a_36_160# vdd 0.006001f
C15534 trimb[1] _452_/a_3129_107# 0.007229f
C15535 mask\[4\] _346_/a_665_69# 0.001125f
C15536 net74 trim_mask\[4\] 0.548293f
C15537 FILLER_0_7_162/a_36_472# _074_ 0.003809f
C15538 FILLER_0_12_136/a_1020_375# vdd 0.017472f
C15539 FILLER_0_12_136/a_572_375# vss 0.006091f
C15540 ctln[1] net2 0.126801f
C15541 _144_ FILLER_0_18_107/a_1916_375# 0.003148f
C15542 _402_/a_56_567# vdd 0.014708f
C15543 _065_ output16/a_224_472# 0.049052f
C15544 FILLER_0_9_28/a_36_472# FILLER_0_10_28/a_36_472# 0.05841f
C15545 _114_ _225_/a_36_160# 0.003628f
C15546 result[5] result[6] 0.065361f
C15547 _114_ _308_/a_124_24# 0.052818f
C15548 _431_/a_448_472# net53 0.002087f
C15549 _444_/a_1308_423# FILLER_0_8_24/a_36_472# 0.009119f
C15550 net20 _418_/a_2665_112# 0.013517f
C15551 net53 _451_/a_2225_156# 0.011677f
C15552 _423_/a_1308_423# _012_ 0.01389f
C15553 net62 mask\[0\] 0.552008f
C15554 ctlp[4] mask\[7\] 0.080163f
C15555 result[5] fanout61/a_36_113# 0.001866f
C15556 cal_itt\[3\] _163_ 0.021146f
C15557 FILLER_0_1_98/a_124_375# _442_/a_2665_112# 0.003045f
C15558 net73 FILLER_0_19_111/a_572_375# 0.04458f
C15559 FILLER_0_17_104/a_484_472# net14 0.004272f
C15560 _307_/a_234_472# vdd 0.001209f
C15561 net79 _286_/a_224_472# 0.001276f
C15562 _031_ _369_/a_36_68# 0.050502f
C15563 _159_ vdd 0.025131f
C15564 _116_ _085_ 0.049304f
C15565 result[8] _048_ 0.006006f
C15566 _105_ _204_/a_67_603# 0.061486f
C15567 FILLER_0_3_172/a_2724_472# net22 0.012284f
C15568 net79 FILLER_0_12_220/a_124_375# 0.010895f
C15569 _427_/a_2665_112# _043_ 0.002612f
C15570 _081_ _163_ 0.427672f
C15571 net14 _156_ 0.184287f
C15572 _104_ ctlp[3] 0.025066f
C15573 mask\[5\] _141_ 0.241158f
C15574 _417_/a_2560_156# vdd 0.001658f
C15575 _417_/a_2665_112# vss 0.002571f
C15576 net62 _417_/a_1204_472# 0.001941f
C15577 ctln[1] cal 0.123834f
C15578 fanout51/a_36_113# FILLER_0_11_78/a_124_375# 0.005683f
C15579 output20/a_224_472# ctlp[2] 0.085373f
C15580 _424_/a_2248_156# _012_ 0.009377f
C15581 _412_/a_2248_156# cal_itt\[1\] 0.005868f
C15582 net48 _316_/a_124_24# 0.068708f
C15583 FILLER_0_18_2/a_124_375# vss 0.003207f
C15584 _130_ _428_/a_2665_112# 0.001241f
C15585 cal_count\[3\] _136_ 0.00703f
C15586 mask\[5\] _295_/a_36_472# 0.034027f
C15587 FILLER_0_18_53/a_572_375# vss 0.057185f
C15588 FILLER_0_18_53/a_36_472# vdd 0.089087f
C15589 _128_ _068_ 0.863174f
C15590 net35 FILLER_0_22_177/a_484_472# 0.00632f
C15591 FILLER_0_10_78/a_1468_375# vdd 0.001778f
C15592 FILLER_0_22_86/a_932_472# net71 0.005789f
C15593 FILLER_0_16_107/a_124_375# _451_/a_36_151# 0.001597f
C15594 output48/a_224_472# en 0.003074f
C15595 _415_/a_448_472# net27 0.05785f
C15596 _104_ net31 0.102776f
C15597 net20 FILLER_0_15_228/a_124_375# 0.047331f
C15598 FILLER_0_16_107/a_36_472# _040_ 0.015026f
C15599 _413_/a_36_151# _002_ 0.0076f
C15600 FILLER_0_3_172/a_2364_375# vdd -0.010717f
C15601 _052_ FILLER_0_21_28/a_2364_375# 0.002388f
C15602 FILLER_0_21_206/a_36_472# net21 0.132984f
C15603 net31 _421_/a_2665_112# 0.005428f
C15604 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3172_472# 0.013276f
C15605 FILLER_0_21_28/a_1020_375# net17 0.001134f
C15606 _438_/a_448_472# net14 0.020612f
C15607 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1380_472# 0.026657f
C15608 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_36_472# 0.002765f
C15609 _001_ cal_itt\[0\] 0.004843f
C15610 FILLER_0_13_212/a_1468_375# _043_ 0.01418f
C15611 _093_ FILLER_0_18_107/a_484_472# 0.008683f
C15612 net69 net13 0.005834f
C15613 en net5 0.892091f
C15614 _079_ FILLER_0_3_172/a_1828_472# 0.001638f
C15615 FILLER_0_11_142/a_36_472# _076_ 0.003047f
C15616 fanout69/a_36_113# net74 0.034782f
C15617 FILLER_0_12_2/a_36_472# vdd 0.104425f
C15618 FILLER_0_12_2/a_572_375# vss 0.017629f
C15619 net19 _044_ 0.138869f
C15620 _142_ _334_/a_36_160# 0.009001f
C15621 _412_/a_2248_156# vss 0.005692f
C15622 cal_count\[3\] _070_ 0.059233f
C15623 _098_ FILLER_0_15_212/a_484_472# 0.00912f
C15624 _444_/a_36_151# net47 0.016691f
C15625 _086_ _163_ 0.413768f
C15626 net31 result[6] 0.002094f
C15627 FILLER_0_8_138/a_124_375# vss 0.00629f
C15628 _093_ FILLER_0_16_89/a_932_472# 0.002018f
C15629 _079_ net37 0.408392f
C15630 _120_ _172_ 0.010275f
C15631 net56 FILLER_0_19_155/a_36_472# 0.00611f
C15632 _131_ _160_ 0.003984f
C15633 _005_ _416_/a_448_472# 0.04044f
C15634 net68 net49 0.607379f
C15635 _053_ FILLER_0_7_104/a_124_375# 0.012564f
C15636 _430_/a_448_472# vdd 0.002959f
C15637 vdd FILLER_0_4_91/a_124_375# 0.019812f
C15638 output27/a_224_472# FILLER_0_9_290/a_124_375# 0.02894f
C15639 _447_/a_2248_156# net69 0.001126f
C15640 _091_ _274_/a_3368_68# 0.001328f
C15641 _086_ _115_ 0.4112f
C15642 _415_/a_2665_112# net62 0.003644f
C15643 result[8] FILLER_0_24_290/a_124_375# 0.00562f
C15644 _277_/a_36_160# vss 0.030147f
C15645 _119_ _163_ 0.009297f
C15646 _267_/a_1568_472# _055_ 0.001681f
C15647 _166_ _034_ 0.001936f
C15648 _448_/a_448_472# net76 0.003937f
C15649 FILLER_0_4_49/a_124_375# _035_ 0.00215f
C15650 net65 net21 0.04444f
C15651 net52 FILLER_0_5_72/a_484_472# 0.050714f
C15652 net50 FILLER_0_5_72/a_1468_375# 0.001777f
C15653 _093_ _136_ 0.226819f
C15654 _445_/a_2665_112# trim_mask\[1\] 0.00183f
C15655 _119_ _115_ 0.06747f
C15656 _130_ _126_ 0.061836f
C15657 net22 _435_/a_448_472# 0.001929f
C15658 _093_ net21 0.032584f
C15659 mask\[0\] _429_/a_448_472# 0.061449f
C15660 FILLER_0_0_130/a_36_472# _442_/a_36_151# 0.001723f
C15661 _239_/a_36_160# net41 0.006002f
C15662 _011_ _009_ 0.035129f
C15663 mask\[4\] net31 0.499009f
C15664 _350_/a_49_472# vss 0.001319f
C15665 net31 net22 0.002533f
C15666 FILLER_0_7_195/a_124_375# cal_itt\[3\] 0.034632f
C15667 FILLER_0_15_116/a_36_472# _040_ 0.002896f
C15668 net51 _450_/a_2225_156# 0.009822f
C15669 FILLER_0_2_111/a_484_472# vss -0.001894f
C15670 FILLER_0_2_111/a_932_472# vdd 0.003808f
C15671 _043_ _278_/a_36_160# 0.004357f
C15672 _070_ _169_ 0.006335f
C15673 FILLER_0_20_177/a_572_375# _098_ 0.015373f
C15674 _428_/a_2248_156# _131_ 0.005621f
C15675 net73 vss 0.342554f
C15676 _092_ _291_/a_36_160# 0.03297f
C15677 _103_ _418_/a_36_151# 0.032388f
C15678 _398_/a_36_113# net44 0.011803f
C15679 FILLER_0_15_150/a_124_375# net53 0.041074f
C15680 FILLER_0_9_60/a_484_472# net51 0.061362f
C15681 fanout62/a_36_160# vdd 0.059299f
C15682 _414_/a_1308_423# vdd 0.004897f
C15683 _185_ _278_/a_36_160# 0.001237f
C15684 net78 _419_/a_2248_156# 0.001614f
C15685 _136_ FILLER_0_15_180/a_572_375# 0.001571f
C15686 FILLER_0_5_88/a_124_375# _164_ 0.006288f
C15687 mask\[8\] net71 0.424276f
C15688 FILLER_0_5_206/a_124_375# net22 0.019537f
C15689 net63 FILLER_0_20_177/a_484_472# 0.002172f
C15690 _093_ _356_/a_36_472# 0.009235f
C15691 FILLER_0_20_169/a_124_375# _434_/a_36_151# 0.026916f
C15692 net17 vss 0.940703f
C15693 _086_ _321_/a_3126_472# 0.001522f
C15694 net59 net21 0.157689f
C15695 net34 _435_/a_2248_156# 0.01519f
C15696 FILLER_0_3_2/a_36_472# _446_/a_36_151# 0.004032f
C15697 FILLER_0_7_72/a_572_375# net52 0.022624f
C15698 _415_/a_36_151# vdd 0.115639f
C15699 _012_ _098_ 0.002778f
C15700 _093_ FILLER_0_17_72/a_2364_375# 0.010888f
C15701 FILLER_0_18_2/a_2724_472# _452_/a_448_472# 0.008967f
C15702 net41 _445_/a_2665_112# 0.056125f
C15703 FILLER_0_10_78/a_36_472# vss 0.008832f
C15704 FILLER_0_22_86/a_1468_375# _211_/a_36_160# 0.010334f
C15705 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_484_472# 0.026657f
C15706 output35/a_224_472# net21 0.069263f
C15707 FILLER_0_7_162/a_124_375# net57 0.033245f
C15708 net81 _429_/a_796_472# 0.002847f
C15709 FILLER_0_8_107/a_36_472# vss 0.006371f
C15710 net63 FILLER_0_18_177/a_124_375# 0.001937f
C15711 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_124_375# 0.009654f
C15712 _430_/a_2248_156# _069_ 0.042876f
C15713 _053_ _372_/a_3662_472# 0.002006f
C15714 _413_/a_448_472# FILLER_0_1_192/a_36_472# 0.001462f
C15715 result[5] _418_/a_448_472# 0.007308f
C15716 fanout74/a_36_113# _371_/a_36_113# 0.01088f
C15717 FILLER_0_9_223/a_572_375# vss 0.00704f
C15718 _099_ _195_/a_255_603# 0.002146f
C15719 _105_ _201_/a_67_603# 0.003335f
C15720 _444_/a_2248_156# FILLER_0_6_37/a_124_375# 0.001101f
C15721 cal_count\[3\] FILLER_0_11_78/a_572_375# 0.010243f
C15722 _115_ FILLER_0_9_142/a_124_375# 0.010167f
C15723 _098_ FILLER_0_15_235/a_484_472# 0.004898f
C15724 _275_/a_224_472# _091_ 0.003461f
C15725 net45 output17/a_224_472# 0.01994f
C15726 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_36_472# 0.009654f
C15727 _256_/a_244_497# _128_ 0.002372f
C15728 _098_ _438_/a_448_472# 0.008962f
C15729 cal_count\[3\] FILLER_0_12_50/a_36_472# 0.063276f
C15730 net63 FILLER_0_19_171/a_1380_472# 0.003014f
C15731 _073_ _081_ 0.046537f
C15732 net58 net2 0.070564f
C15733 FILLER_0_15_150/a_36_472# net23 0.010444f
C15734 mask\[3\] _282_/a_36_160# 0.005823f
C15735 _452_/a_36_151# vss 0.02741f
C15736 _452_/a_448_472# vdd 0.019824f
C15737 _429_/a_1204_472# net22 0.001899f
C15738 net75 _415_/a_36_151# 0.024047f
C15739 _077_ net74 0.025882f
C15740 result[8] result[9] 0.242998f
C15741 net17 _452_/a_836_156# 0.002817f
C15742 FILLER_0_9_28/a_1020_375# net68 0.004803f
C15743 _450_/a_2225_156# net6 0.001143f
C15744 _143_ vss 0.02001f
C15745 FILLER_0_17_72/a_2724_472# vdd 0.007064f
C15746 FILLER_0_17_72/a_2276_472# vss -0.001288f
C15747 _028_ FILLER_0_7_104/a_124_375# 0.008248f
C15748 _425_/a_36_151# FILLER_0_8_247/a_484_472# 0.059367f
C15749 FILLER_0_16_37/a_36_472# vss 0.005874f
C15750 net58 _412_/a_448_472# 0.044616f
C15751 net32 net33 0.467071f
C15752 _274_/a_36_68# state\[0\] 0.001852f
C15753 _104_ net60 0.063407f
C15754 _053_ FILLER_0_5_54/a_1380_472# 0.00114f
C15755 FILLER_0_21_142/a_572_375# vdd 0.002442f
C15756 net60 _421_/a_2665_112# 0.044114f
C15757 _274_/a_1612_497# net4 0.00807f
C15758 FILLER_0_19_195/a_36_472# net21 0.009159f
C15759 _418_/a_2665_112# vss 0.003519f
C15760 _418_/a_2560_156# vdd 0.001506f
C15761 mask\[0\] _056_ 0.001878f
C15762 net15 _423_/a_1000_472# 0.001786f
C15763 _422_/a_2560_156# mask\[7\] 0.010664f
C15764 _390_/a_36_68# _171_ 0.001252f
C15765 net58 cal 0.001209f
C15766 _074_ _056_ 0.002397f
C15767 _426_/a_36_151# _425_/a_1308_423# 0.001518f
C15768 net57 _428_/a_1204_472# 0.015233f
C15769 _140_ _146_ 0.135012f
C15770 _091_ FILLER_0_15_212/a_932_472# 0.008749f
C15771 _450_/a_2449_156# net40 0.010265f
C15772 net61 _422_/a_1000_472# 0.001947f
C15773 net56 fanout54/a_36_160# 0.044466f
C15774 _000_ _080_ 0.002867f
C15775 result[7] net78 0.019651f
C15776 ctln[8] net14 0.001447f
C15777 output24/a_224_472# ctlp[7] 0.060657f
C15778 trimb[3] FILLER_0_20_2/a_484_472# 0.001829f
C15779 net31 _419_/a_2248_156# 0.001521f
C15780 _102_ net19 0.011979f
C15781 FILLER_0_4_213/a_484_472# net59 0.048997f
C15782 _253_/a_36_68# _082_ 0.013108f
C15783 _126_ _428_/a_2248_156# 0.001131f
C15784 en_co_clk _095_ 0.003753f
C15785 FILLER_0_17_72/a_1020_375# net36 0.001777f
C15786 result[6] net60 0.094624f
C15787 FILLER_0_12_28/a_36_472# vdd 0.095598f
C15788 FILLER_0_12_28/a_124_375# vss 0.013117f
C15789 net44 cal_count\[2\] 0.191151f
C15790 FILLER_0_16_89/a_124_375# _176_ 0.002781f
C15791 _028_ FILLER_0_5_72/a_932_472# 0.003042f
C15792 _428_/a_796_472# _043_ 0.007935f
C15793 _322_/a_124_24# _125_ 0.01165f
C15794 FILLER_0_18_177/a_3260_375# _047_ 0.030543f
C15795 _052_ _424_/a_1000_472# 0.007574f
C15796 _021_ _093_ 0.049589f
C15797 net34 FILLER_0_22_128/a_2276_472# 0.005532f
C15798 _441_/a_1308_423# vdd 0.002837f
C15799 _441_/a_448_472# vss 0.025073f
C15800 FILLER_0_21_150/a_36_472# _146_ 0.00236f
C15801 _098_ _434_/a_1204_472# 0.006257f
C15802 _235_/a_67_603# vss 0.002019f
C15803 FILLER_0_13_212/a_36_472# mask\[0\] 0.001366f
C15804 _449_/a_2665_112# en_co_clk 0.002966f
C15805 net72 _452_/a_448_472# 0.001296f
C15806 ctln[8] _447_/a_2665_112# 0.001271f
C15807 _442_/a_2665_112# trim_mask\[3\] 0.019514f
C15808 FILLER_0_4_152/a_124_375# trim_mask\[4\] 0.01182f
C15809 _394_/a_56_524# FILLER_0_15_59/a_484_472# 0.001033f
C15810 _394_/a_718_524# FILLER_0_15_59/a_572_375# 0.001447f
C15811 mask\[3\] FILLER_0_18_177/a_1916_375# 0.003052f
C15812 trim_mask\[2\] net17 0.084388f
C15813 _117_ _310_/a_49_472# 0.018229f
C15814 _193_/a_36_160# _044_ 0.025719f
C15815 mask\[5\] ctlp[2] 0.104304f
C15816 result[7] result[5] 0.016166f
C15817 FILLER_0_15_228/a_124_375# vss 0.006435f
C15818 FILLER_0_15_228/a_36_472# vdd 0.084606f
C15819 net79 _138_ 0.024731f
C15820 _412_/a_36_151# fanout81/a_36_160# 0.001725f
C15821 _238_/a_67_603# vss 0.008203f
C15822 _036_ _164_ 0.011115f
C15823 _176_ _390_/a_36_68# 0.005007f
C15824 net15 _029_ 0.111797f
C15825 FILLER_0_11_101/a_572_375# _120_ 0.006382f
C15826 _447_/a_1308_423# net17 0.002531f
C15827 _440_/a_1204_472# vss 0.007007f
C15828 _440_/a_2248_156# vdd -0.003421f
C15829 net55 FILLER_0_17_72/a_1380_472# 0.021108f
C15830 FILLER_0_19_142/a_124_375# vss 0.032026f
C15831 FILLER_0_19_142/a_36_472# vdd 0.107105f
C15832 FILLER_0_4_185/a_124_375# vss 0.024832f
C15833 _112_ _425_/a_448_472# 0.002335f
C15834 output29/a_224_472# net30 0.044542f
C15835 _439_/a_36_151# vss 0.032466f
C15836 _439_/a_448_472# vdd 0.006996f
C15837 fanout58/a_36_160# input4/a_36_68# 0.059453f
C15838 vdd FILLER_0_13_290/a_124_375# 0.031436f
C15839 mask\[7\] _350_/a_49_472# 0.035293f
C15840 _062_ _055_ 0.29425f
C15841 _092_ mask\[3\] 0.040554f
C15842 net54 _022_ 0.004106f
C15843 _443_/a_2665_112# _170_ 0.019855f
C15844 _061_ _060_ 0.066418f
C15845 _141_ _348_/a_49_472# 0.037821f
C15846 net76 FILLER_0_5_181/a_124_375# 0.031324f
C15847 cal_itt\[2\] _081_ 0.003204f
C15848 _327_/a_36_472# _016_ 0.04536f
C15849 FILLER_0_19_47/a_484_472# vdd 0.001133f
C15850 FILLER_0_19_47/a_36_472# vss 0.001559f
C15851 _131_ FILLER_0_17_104/a_484_472# 0.003483f
C15852 _176_ cal_count\[2\] 0.005783f
C15853 net36 mask\[2\] 0.871463f
C15854 net20 _078_ 0.105266f
C15855 _426_/a_36_151# FILLER_0_8_247/a_572_375# 0.059049f
C15856 net57 _069_ 0.026933f
C15857 _008_ net78 0.032202f
C15858 _414_/a_36_151# _057_ 0.003902f
C15859 net1 _081_ 0.111227f
C15860 FILLER_0_18_2/a_36_472# vdd 0.104532f
C15861 net56 FILLER_0_18_139/a_124_375# 0.00281f
C15862 FILLER_0_6_47/a_2276_472# vdd 0.002735f
C15863 FILLER_0_6_47/a_1828_472# vss 0.003457f
C15864 _316_/a_692_472# vdd 0.001634f
C15865 _175_ FILLER_0_15_72/a_572_375# 0.04785f
C15866 FILLER_0_4_144/a_36_472# net23 0.016933f
C15867 net39 vss 0.170972f
C15868 _428_/a_36_151# FILLER_0_14_107/a_124_375# 0.001597f
C15869 FILLER_0_21_206/a_124_375# _048_ 0.018458f
C15870 net50 FILLER_0_6_37/a_124_375# 0.003821f
C15871 _098_ _113_ 0.001472f
C15872 _201_/a_67_603# _047_ 0.013357f
C15873 net65 valid 0.074257f
C15874 vss _039_ 0.180364f
C15875 _010_ _108_ 0.002048f
C15876 FILLER_0_10_37/a_36_472# net68 0.005405f
C15877 _079_ _122_ 0.003853f
C15878 _161_ _163_ 0.024512f
C15879 output42/a_224_472# net38 0.066219f
C15880 FILLER_0_18_171/a_124_375# _091_ 0.034351f
C15881 _091_ _137_ 0.486022f
C15882 _412_/a_2665_112# en 0.015256f
C15883 mask\[0\] FILLER_0_12_196/a_124_375# 0.034009f
C15884 mask\[9\] FILLER_0_20_107/a_124_375# 0.004716f
C15885 _291_/a_36_160# vdd 0.010802f
C15886 FILLER_0_21_142/a_124_375# _433_/a_2560_156# 0.001178f
C15887 FILLER_0_15_205/a_36_472# net22 0.037011f
C15888 net53 FILLER_0_17_142/a_484_472# 0.001286f
C15889 _207_/a_67_603# vdd 0.034688f
C15890 result[5] _008_ 0.165753f
C15891 net54 FILLER_0_18_107/a_36_472# 0.002116f
C15892 net70 FILLER_0_14_123/a_36_472# 0.009456f
C15893 _367_/a_36_68# vdd 0.010246f
C15894 FILLER_0_22_86/a_484_472# net14 0.006746f
C15895 _091_ FILLER_0_19_171/a_36_472# 0.029168f
C15896 output14/a_224_472# vss 0.012129f
C15897 output46/a_224_472# FILLER_0_20_2/a_124_375# 0.030009f
C15898 _026_ net71 0.406369f
C15899 result[7] net31 0.231528f
C15900 net69 _160_ 0.077526f
C15901 FILLER_0_5_109/a_484_472# net47 0.002299f
C15902 _077_ FILLER_0_9_72/a_124_375# 0.008103f
C15903 _427_/a_1308_423# vss 0.030292f
C15904 net68 FILLER_0_8_37/a_36_472# 0.001088f
C15905 FILLER_0_9_223/a_572_375# net4 0.02077f
C15906 valid net59 0.577796f
C15907 _412_/a_796_472# cal_itt\[1\] 0.004226f
C15908 _406_/a_36_159# _185_ 0.001573f
C15909 _257_/a_36_472# vss 0.023401f
C15910 net65 net9 0.061456f
C15911 _053_ _414_/a_448_472# 0.065053f
C15912 _273_/a_36_68# _090_ 0.034955f
C15913 net75 _316_/a_692_472# 0.00138f
C15914 _448_/a_36_151# FILLER_0_2_177/a_124_375# 0.001597f
C15915 FILLER_0_9_28/a_1828_472# net68 0.048468f
C15916 _179_ cal_count\[1\] 0.088667f
C15917 vss FILLER_0_8_156/a_36_472# 0.00168f
C15918 vdd FILLER_0_8_156/a_484_472# 0.007249f
C15919 net76 vdd 1.272072f
C15920 mask\[4\] _433_/a_2665_112# 0.005353f
C15921 net20 _411_/a_448_472# 0.002167f
C15922 FILLER_0_16_107/a_484_472# _136_ 0.013449f
C15923 _449_/a_1308_423# _067_ 0.021042f
C15924 _033_ _444_/a_1000_472# 0.00692f
C15925 _165_ _444_/a_2665_112# 0.044447f
C15926 _110_ mask\[8\] 0.05045f
C15927 net49 net47 0.53353f
C15928 _068_ _311_/a_2700_473# 0.001846f
C15929 _211_/a_36_160# net71 0.035804f
C15930 net76 FILLER_0_6_177/a_572_375# 0.073022f
C15931 _058_ _062_ 1.676625f
C15932 _235_/a_67_603# trim_mask\[2\] 0.022726f
C15933 _370_/a_692_472# _081_ 0.00129f
C15934 _370_/a_848_380# _152_ 0.031499f
C15935 _108_ vdd 0.298249f
C15936 _177_ _176_ 0.226424f
C15937 _238_/a_67_603# FILLER_0_1_98/a_36_472# 0.02529f
C15938 net68 net47 0.063835f
C15939 _426_/a_36_151# _317_/a_36_113# 0.001082f
C15940 _070_ _120_ 0.838223f
C15941 cal_count\[3\] _373_/a_632_68# 0.004529f
C15942 _173_ vdd 0.080629f
C15943 net60 _418_/a_448_472# 0.055895f
C15944 net31 _008_ 0.292444f
C15945 _238_/a_67_603# trim_mask\[2\] 0.003021f
C15946 net60 _419_/a_2248_156# 0.047724f
C15947 net61 _419_/a_2560_156# 0.008214f
C15948 net58 FILLER_0_9_290/a_124_375# 0.001157f
C15949 _140_ _147_ 0.08953f
C15950 cal_count\[2\] _183_ 0.034303f
C15951 output29/a_224_472# FILLER_0_14_263/a_36_472# 0.0323f
C15952 FILLER_0_7_195/a_124_375# _161_ 0.005368f
C15953 trimb[3] vss 0.161605f
C15954 net27 _425_/a_2665_112# 0.001323f
C15955 FILLER_0_19_47/a_36_472# _424_/a_448_472# 0.004782f
C15956 FILLER_0_4_99/a_124_375# FILLER_0_4_91/a_572_375# 0.012001f
C15957 result[8] net61 0.001106f
C15958 en_co_clk net74 0.039096f
C15959 fanout73/a_36_113# net36 0.01199f
C15960 FILLER_0_7_59/a_124_375# vss 0.002006f
C15961 FILLER_0_7_59/a_572_375# vdd 0.005991f
C15962 FILLER_0_12_28/a_36_472# cal_count\[0\] 0.001662f
C15963 _430_/a_36_151# fanout80/a_36_113# 0.018169f
C15964 _086_ _121_ 0.049499f
C15965 net75 net76 0.106326f
C15966 _115_ _127_ 0.042389f
C15967 net35 FILLER_0_22_128/a_2364_375# 0.012732f
C15968 FILLER_0_9_28/a_1020_375# FILLER_0_10_37/a_36_472# 0.001597f
C15969 FILLER_0_1_204/a_124_375# vdd 0.047704f
C15970 _064_ output39/a_224_472# 0.107406f
C15971 net20 FILLER_0_6_231/a_36_472# 0.045553f
C15972 net68 FILLER_0_6_47/a_124_375# 0.002491f
C15973 _091_ _248_/a_36_68# 0.071763f
C15974 _092_ FILLER_0_17_218/a_124_375# 0.020704f
C15975 _002_ vss 0.08396f
C15976 _136_ FILLER_0_16_154/a_124_375# 0.00252f
C15977 trim_mask\[1\] FILLER_0_6_47/a_1020_375# 0.007169f
C15978 FILLER_0_9_142/a_36_472# _120_ 0.035902f
C15979 _119_ _121_ 0.007336f
C15980 _091_ net81 0.03653f
C15981 output15/a_224_472# _164_ 0.031363f
C15982 fanout51/a_36_113# net55 0.010147f
C15983 _114_ FILLER_0_12_136/a_1468_375# 0.006974f
C15984 net53 FILLER_0_14_99/a_124_375# 0.00494f
C15985 FILLER_0_5_109/a_36_472# _163_ 0.00319f
C15986 _086_ FILLER_0_7_104/a_124_375# 0.001629f
C15987 net38 net6 0.071232f
C15988 result[4] FILLER_0_15_290/a_36_472# 0.001422f
C15989 _070_ FILLER_0_9_105/a_572_375# 0.017191f
C15990 _165_ _160_ 0.008705f
C15991 FILLER_0_18_177/a_1380_472# _139_ 0.00195f
C15992 _444_/a_36_151# vdd 0.071209f
C15993 FILLER_0_22_86/a_484_472# _098_ 0.003294f
C15994 net20 net36 0.03843f
C15995 _095_ _181_ 0.008117f
C15996 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_36_472# 0.001723f
C15997 _091_ _060_ 0.085764f
C15998 _027_ _438_/a_36_151# 0.010763f
C15999 _150_ _438_/a_1308_423# 0.001472f
C16000 _421_/a_36_151# _419_/a_448_472# 0.002098f
C16001 _427_/a_36_151# net23 0.006844f
C16002 ctlp[0] vss 0.005302f
C16003 net55 _451_/a_2225_156# 0.031243f
C16004 _065_ _441_/a_2665_112# 0.003318f
C16005 FILLER_0_8_138/a_36_472# vdd 0.008749f
C16006 net69 _170_ 0.006468f
C16007 net15 FILLER_0_5_72/a_36_472# 0.006713f
C16008 _307_/a_672_472# _114_ 0.0018f
C16009 _065_ _447_/a_1000_472# 0.03162f
C16010 _446_/a_1000_472# _035_ 0.00349f
C16011 _273_/a_36_68# _076_ 0.001503f
C16012 FILLER_0_14_50/a_124_375# _179_ 0.021823f
C16013 net81 FILLER_0_9_270/a_36_472# 0.084422f
C16014 FILLER_0_21_125/a_124_375# mask\[7\] 0.00145f
C16015 FILLER_0_7_72/a_3260_375# _058_ 0.00258f
C16016 mask\[3\] vdd 0.340612f
C16017 _432_/a_2560_156# net80 0.01523f
C16018 fanout50/a_36_160# _168_ 0.033707f
C16019 net52 _384_/a_224_472# 0.001238f
C16020 FILLER_0_9_28/a_3260_375# vss 0.05542f
C16021 _015_ _426_/a_2560_156# 0.024461f
C16022 result[4] FILLER_0_17_282/a_36_472# 0.017375f
C16023 FILLER_0_12_50/a_124_375# _067_ 0.011869f
C16024 _067_ _450_/a_2225_156# 0.002584f
C16025 net42 vss 0.017902f
C16026 result[9] _103_ 0.034463f
C16027 FILLER_0_11_78/a_572_375# _120_ 0.01683f
C16028 FILLER_0_21_125/a_36_472# net54 0.016672f
C16029 _182_ _401_/a_36_68# 0.088487f
C16030 FILLER_0_9_72/a_36_472# vss 0.0392f
C16031 FILLER_0_9_72/a_484_472# vdd 0.005654f
C16032 net41 _450_/a_3129_107# 0.059083f
C16033 net27 _426_/a_796_472# 0.001678f
C16034 _070_ _227_/a_36_160# 0.00254f
C16035 _272_/a_36_472# _089_ 0.003862f
C16036 _171_ FILLER_0_10_94/a_484_472# 0.001446f
C16037 _131_ _118_ 0.001685f
C16038 net32 net18 0.028135f
C16039 _451_/a_836_156# net14 0.00174f
C16040 result[7] net60 0.778099f
C16041 net55 FILLER_0_13_72/a_36_472# 0.002172f
C16042 net55 net51 0.007067f
C16043 _057_ _228_/a_36_68# 0.002062f
C16044 _326_/a_36_160# FILLER_0_9_105/a_572_375# 0.005489f
C16045 FILLER_0_16_57/a_932_472# net55 0.00179f
C16046 FILLER_0_2_111/a_572_375# _160_ 0.001049f
C16047 _083_ vdd 0.157549f
C16048 _359_/a_36_488# vss 0.002427f
C16049 _078_ vss 0.367953f
C16050 fanout72/a_36_113# _067_ 0.005796f
C16051 output19/a_224_472# net19 0.030721f
C16052 net29 _196_/a_36_160# 0.073294f
C16053 FILLER_0_12_50/a_36_472# _120_ 0.005447f
C16054 FILLER_0_1_192/a_124_375# net59 0.014491f
C16055 output8/a_224_472# FILLER_0_3_221/a_36_472# 0.001699f
C16056 _390_/a_244_472# _136_ 0.001777f
C16057 FILLER_0_13_212/a_124_375# FILLER_0_13_206/a_124_375# 0.005439f
C16058 net44 FILLER_0_20_2/a_124_375# 0.001564f
C16059 FILLER_0_9_28/a_3172_472# FILLER_0_9_60/a_36_472# 0.013276f
C16060 net43 FILLER_0_20_15/a_572_375# 0.003924f
C16061 net57 FILLER_0_13_142/a_36_472# 0.011199f
C16062 _320_/a_1568_472# _043_ 0.00177f
C16063 net18 _417_/a_1204_472# 0.01349f
C16064 FILLER_0_4_152/a_124_375# _066_ 0.003354f
C16065 _432_/a_1000_472# _137_ 0.008914f
C16066 trimb[1] FILLER_0_18_2/a_1468_375# 0.002041f
C16067 fanout66/a_36_113# net49 0.001044f
C16068 FILLER_0_20_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001543f
C16069 FILLER_0_15_282/a_36_472# output30/a_224_472# 0.001711f
C16070 vss _416_/a_796_472# 0.001468f
C16071 net62 _416_/a_448_472# 0.009111f
C16072 _367_/a_244_472# _154_ 0.001775f
C16073 vss clkc 0.0311f
C16074 net68 fanout66/a_36_113# 0.01746f
C16075 _408_/a_728_93# _186_ 0.003815f
C16076 FILLER_0_20_169/a_36_472# _339_/a_36_160# 0.001448f
C16077 net65 _084_ 0.031674f
C16078 _105_ net33 0.202272f
C16079 mask\[2\] FILLER_0_16_154/a_1468_375# 0.014254f
C16080 FILLER_0_13_142/a_1020_375# _043_ 0.005672f
C16081 FILLER_0_19_125/a_124_375# _345_/a_36_160# 0.005398f
C16082 FILLER_0_14_91/a_572_375# _176_ 0.002444f
C16083 _035_ _034_ 1.26804f
C16084 _057_ calibrate 0.002047f
C16085 net48 _425_/a_448_472# 0.013011f
C16086 _094_ _045_ 0.102437f
C16087 _431_/a_1308_423# _427_/a_36_151# 0.001256f
C16088 _176_ FILLER_0_10_94/a_484_472# 0.009483f
C16089 _086_ FILLER_0_11_124/a_124_375# 0.016039f
C16090 _140_ FILLER_0_22_128/a_36_472# 0.050084f
C16091 net20 result[4] 0.001673f
C16092 mask\[0\] FILLER_0_15_212/a_1468_375# 0.001182f
C16093 net31 _006_ 0.307613f
C16094 FILLER_0_20_169/a_124_375# mask\[6\] 0.001178f
C16095 FILLER_0_18_76/a_124_375# net71 0.008427f
C16096 _428_/a_2665_112# _118_ 0.001007f
C16097 _141_ _143_ 0.192528f
C16098 FILLER_0_21_28/a_2724_472# vdd 0.001342f
C16099 FILLER_0_6_90/a_572_375# vdd 0.028324f
C16100 FILLER_0_22_128/a_3260_375# _146_ 0.004692f
C16101 ctlp[1] FILLER_0_24_274/a_1020_375# 0.004803f
C16102 _091_ _095_ 0.005006f
C16103 net69 _156_ 0.008057f
C16104 _286_/a_224_472# _005_ 0.001254f
C16105 net35 _436_/a_1204_472# 0.005186f
C16106 _008_ net60 0.314106f
C16107 net15 FILLER_0_5_54/a_484_472# 0.002186f
C16108 trim_mask\[4\] _370_/a_124_24# 0.015021f
C16109 net75 _083_ 0.055491f
C16110 _114_ _134_ 0.015298f
C16111 FILLER_0_18_2/a_1828_472# vdd 0.001953f
C16112 net52 FILLER_0_2_111/a_36_472# 0.0659f
C16113 _415_/a_2665_112# net18 0.004988f
C16114 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_36_472# 0.009654f
C16115 cal_itt\[2\] FILLER_0_3_221/a_484_472# 0.016997f
C16116 _372_/a_2034_472# _076_ 0.007461f
C16117 _372_/a_170_472# _068_ 0.037034f
C16118 _126_ _113_ 0.547055f
C16119 FILLER_0_21_28/a_572_375# FILLER_0_20_31/a_124_375# 0.026339f
C16120 _129_ _076_ 0.043637f
C16121 FILLER_0_11_282/a_36_472# vdd 0.106843f
C16122 FILLER_0_11_282/a_124_375# vss 0.005415f
C16123 FILLER_0_4_107/a_36_472# _157_ 0.005289f
C16124 _374_/a_36_68# FILLER_0_8_156/a_484_472# 0.002559f
C16125 _173_ cal_count\[0\] 0.517178f
C16126 _163_ FILLER_0_5_148/a_572_375# 0.001706f
C16127 fanout65/a_36_113# net5 0.027955f
C16128 _411_/a_448_472# vss 0.009447f
C16129 FILLER_0_17_72/a_36_472# _131_ 0.002672f
C16130 net57 net22 0.003595f
C16131 fanout82/a_36_113# net19 0.021188f
C16132 output19/a_224_472# _009_ 0.003174f
C16133 vss FILLER_0_14_235/a_572_375# 0.017196f
C16134 net82 net2 0.451147f
C16135 _425_/a_448_472# net19 0.034226f
C16136 FILLER_0_14_99/a_124_375# _451_/a_36_151# 0.001441f
C16137 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_484_472# 0.013276f
C16138 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_124_375# 0.009654f
C16139 net81 FILLER_0_15_212/a_484_472# 0.00169f
C16140 trim_mask\[1\] FILLER_0_6_79/a_36_472# 0.006265f
C16141 net38 FILLER_0_15_2/a_572_375# 0.007477f
C16142 _341_/a_665_69# net23 0.001508f
C16143 FILLER_0_14_181/a_36_472# _138_ 0.002748f
C16144 FILLER_0_21_28/a_572_375# FILLER_0_19_28/a_484_472# 0.001512f
C16145 FILLER_0_5_206/a_36_472# net37 0.009858f
C16146 _334_/a_36_160# vss 0.002713f
C16147 _053_ _377_/a_36_472# 0.023504f
C16148 FILLER_0_11_109/a_124_375# FILLER_0_9_105/a_484_472# 0.0027f
C16149 FILLER_0_16_89/a_36_472# _177_ 0.048163f
C16150 _412_/a_448_472# net82 0.030379f
C16151 FILLER_0_0_130/a_124_375# _031_ 0.001861f
C16152 _164_ FILLER_0_6_47/a_1020_375# 0.004285f
C16153 _431_/a_3041_156# vss 0.001312f
C16154 _037_ net22 0.079675f
C16155 FILLER_0_10_78/a_1468_375# _171_ 0.034647f
C16156 _147_ _435_/a_36_151# 0.003096f
C16157 _126_ _118_ 0.215385f
C16158 _253_/a_36_68# net19 0.019615f
C16159 ctlp[7] vss 0.036681f
C16160 _132_ FILLER_0_18_107/a_2364_375# 0.006403f
C16161 _079_ net8 0.001928f
C16162 _431_/a_2248_156# _136_ 0.030673f
C16163 _053_ FILLER_0_8_107/a_36_472# 0.013669f
C16164 FILLER_0_7_233/a_124_375# FILLER_0_6_231/a_484_472# 0.001684f
C16165 _320_/a_36_472# state\[1\] 0.013058f
C16166 FILLER_0_15_150/a_124_375# net23 0.03361f
C16167 _058_ FILLER_0_8_156/a_572_375# 0.007692f
C16168 FILLER_0_12_2/a_36_472# net44 0.011079f
C16169 FILLER_0_12_20/a_484_472# vss 0.001783f
C16170 net78 _007_ 0.054904f
C16171 FILLER_0_17_218/a_124_375# vdd 0.00593f
C16172 _432_/a_448_472# _093_ 0.048289f
C16173 _435_/a_2665_112# vdd 0.01769f
C16174 FILLER_0_8_263/a_124_375# vdd 0.032664f
C16175 vdd FILLER_0_6_231/a_484_472# 0.004642f
C16176 vss FILLER_0_6_231/a_36_472# 0.0048f
C16177 trim[4] _221_/a_36_160# 0.002685f
C16178 _396_/a_224_472# _095_ 0.001351f
C16179 FILLER_0_20_31/a_124_375# vdd 0.04619f
C16180 net67 FILLER_0_9_60/a_572_375# 0.011073f
C16181 cal_count\[3\] _228_/a_36_68# 0.01871f
C16182 _130_ net74 0.001655f
C16183 _423_/a_36_151# net40 0.004045f
C16184 _176_ FILLER_0_18_53/a_36_472# 0.001868f
C16185 _091_ net64 0.079488f
C16186 _181_ cal_count\[1\] 0.186904f
C16187 net70 FILLER_0_13_100/a_124_375# 0.017886f
C16188 FILLER_0_20_87/a_124_375# vss 0.00279f
C16189 FILLER_0_20_87/a_36_472# vdd 0.006784f
C16190 FILLER_0_16_107/a_572_375# net70 0.002193f
C16191 FILLER_0_10_78/a_1468_375# _176_ 0.013408f
C16192 _152_ _261_/a_36_160# 0.001102f
C16193 net16 _408_/a_1336_472# 0.022364f
C16194 net25 vss 0.528437f
C16195 _451_/a_3129_107# _040_ 0.004116f
C16196 _091_ mask\[1\] 0.064614f
C16197 _440_/a_448_472# _160_ 0.004748f
C16198 _414_/a_448_472# cal_itt\[3\] 0.109704f
C16199 FILLER_0_22_86/a_124_375# _437_/a_36_151# 0.001597f
C16200 result[5] _007_ 0.0249f
C16201 FILLER_0_20_193/a_484_472# FILLER_0_18_177/a_2364_375# 0.0027f
C16202 FILLER_0_0_198/a_124_375# net59 0.004565f
C16203 net36 vss 1.788802f
C16204 _136_ _043_ 0.040107f
C16205 net26 FILLER_0_23_44/a_932_472# 0.001889f
C16206 _098_ _146_ 0.004276f
C16207 _043_ net21 0.033824f
C16208 FILLER_0_19_28/a_484_472# vdd 0.010504f
C16209 output45/a_224_472# trimb[2] 0.045907f
C16210 _177_ FILLER_0_17_72/a_1468_375# 0.026469f
C16211 _414_/a_448_472# _081_ 0.024533f
C16212 _050_ FILLER_0_22_128/a_1468_375# 0.001661f
C16213 net23 _163_ 0.034799f
C16214 net57 _076_ 0.028356f
C16215 _276_/a_36_160# FILLER_0_18_209/a_484_472# 0.003913f
C16216 FILLER_0_15_2/a_484_472# vss 0.003267f
C16217 output38/a_224_472# net49 0.002434f
C16218 net38 net66 0.040578f
C16219 FILLER_0_4_123/a_36_472# _154_ 0.001043f
C16220 FILLER_0_21_28/a_2724_472# _424_/a_36_151# 0.001723f
C16221 FILLER_0_10_28/a_124_375# net17 0.00917f
C16222 _064_ net40 0.141744f
C16223 net4 _078_ 0.487587f
C16224 _126_ _068_ 0.01065f
C16225 _140_ _433_/a_2665_112# 0.001108f
C16226 _256_/a_2960_68# _056_ 0.001168f
C16227 _115_ net23 0.018953f
C16228 net64 FILLER_0_9_270/a_36_472# 0.014971f
C16229 _137_ _113_ 0.030279f
C16230 mask\[5\] _204_/a_67_603# 0.023791f
C16231 trim[0] _445_/a_36_151# 0.008302f
C16232 net38 _445_/a_1308_423# 0.006454f
C16233 net16 _034_ 0.096088f
C16234 net34 FILLER_0_22_177/a_124_375# 0.006974f
C16235 net81 FILLER_0_15_235/a_484_472# 0.0047f
C16236 net82 FILLER_0_3_172/a_2724_472# 0.007912f
C16237 net40 output41/a_224_472# 0.081551f
C16238 net75 FILLER_0_8_263/a_124_375# 0.001386f
C16239 _041_ vdd 0.19154f
C16240 net75 FILLER_0_6_231/a_484_472# 0.003485f
C16241 _009_ _299_/a_36_472# 0.006927f
C16242 net18 _418_/a_1204_472# 0.01349f
C16243 FILLER_0_4_185/a_36_472# vss 0.002627f
C16244 FILLER_0_5_54/a_1468_375# _440_/a_36_151# 0.059049f
C16245 _411_/a_36_151# net8 0.012319f
C16246 FILLER_0_15_116/a_124_375# _095_ 0.002659f
C16247 net52 _441_/a_36_151# 0.013755f
C16248 net72 FILLER_0_20_31/a_124_375# 0.011347f
C16249 net60 _006_ 0.006254f
C16250 FILLER_0_14_123/a_124_375# vss 0.004985f
C16251 FILLER_0_14_123/a_36_472# vdd 0.088525f
C16252 FILLER_0_9_28/a_2276_472# vss -0.001894f
C16253 net32 _109_ 0.038411f
C16254 fanout63/a_36_160# FILLER_0_15_228/a_124_375# 0.001177f
C16255 _308_/a_848_380# _058_ 0.031449f
C16256 _115_ _439_/a_2248_156# 0.003553f
C16257 _189_/a_67_603# FILLER_0_12_236/a_124_375# 0.00221f
C16258 FILLER_0_5_109/a_484_472# vdd 0.007355f
C16259 FILLER_0_16_107/a_572_375# _132_ 0.007439f
C16260 FILLER_0_19_55/a_124_375# vss 0.001882f
C16261 FILLER_0_19_55/a_36_472# vdd 0.085984f
C16262 FILLER_0_15_142/a_484_472# net56 0.003214f
C16263 net52 _440_/a_1000_472# 0.013793f
C16264 _287_/a_36_472# _094_ 0.029751f
C16265 calibrate _169_ 0.001883f
C16266 net62 _429_/a_2560_156# 0.002164f
C16267 net38 _067_ 0.062447f
C16268 net72 _394_/a_718_524# 0.001558f
C16269 net55 _394_/a_728_93# 0.0026f
C16270 _423_/a_2560_156# vss 0.002241f
C16271 _414_/a_448_472# _089_ 0.003905f
C16272 net54 FILLER_0_19_111/a_484_472# 0.00105f
C16273 FILLER_0_5_54/a_124_375# FILLER_0_6_47/a_932_472# 0.001597f
C16274 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_124_375# 0.009654f
C16275 mask\[4\] FILLER_0_19_171/a_484_472# 0.004669f
C16276 FILLER_0_2_101/a_36_472# net14 0.051153f
C16277 net65 calibrate 0.012434f
C16278 FILLER_0_19_155/a_36_472# _145_ 0.005521f
C16279 _104_ _420_/a_2560_156# 0.002734f
C16280 _077_ FILLER_0_9_105/a_124_375# 0.007189f
C16281 _116_ vss 0.235141f
C16282 _106_ FILLER_0_17_218/a_572_375# 0.022684f
C16283 net72 FILLER_0_19_28/a_484_472# 0.004312f
C16284 net55 FILLER_0_19_28/a_124_375# 0.002644f
C16285 _123_ net37 0.002942f
C16286 net74 _160_ 0.165289f
C16287 FILLER_0_20_169/a_36_472# vss 0.005112f
C16288 _132_ net70 0.534228f
C16289 net15 _453_/a_1308_423# 0.00293f
C16290 net20 _317_/a_36_113# 0.00189f
C16291 net69 FILLER_0_2_111/a_124_375# 0.010762f
C16292 FILLER_0_22_128/a_2724_472# vdd 0.005923f
C16293 FILLER_0_22_128/a_2276_472# vss 0.02979f
C16294 net20 FILLER_0_24_274/a_36_472# 0.009746f
C16295 output13/a_224_472# net22 0.022308f
C16296 _028_ FILLER_0_8_107/a_36_472# 0.002173f
C16297 net32 _421_/a_2248_156# 0.038586f
C16298 result[4] vss 0.306116f
C16299 ctln[1] input5/a_36_113# 0.01908f
C16300 net55 FILLER_0_13_80/a_36_472# 0.016536f
C16301 _178_ _402_/a_728_93# 0.050963f
C16302 _070_ FILLER_0_10_107/a_484_472# 0.007421f
C16303 _144_ _436_/a_36_151# 0.029716f
C16304 en_co_clk _389_/a_36_148# 0.001249f
C16305 _030_ vss 0.117034f
C16306 net49 vdd 0.872948f
C16307 _127_ _121_ 0.023125f
C16308 _086_ _267_/a_1792_472# 0.002715f
C16309 _442_/a_2248_156# vdd 0.038702f
C16310 net72 _041_ 0.467856f
C16311 FILLER_0_6_79/a_36_472# _164_ 0.008685f
C16312 _114_ _311_/a_66_473# 0.081048f
C16313 _183_ FILLER_0_18_53/a_36_472# 0.007412f
C16314 _452_/a_1040_527# _041_ 0.002066f
C16315 _053_ FILLER_0_6_47/a_1828_472# 0.006408f
C16316 _424_/a_36_151# FILLER_0_20_31/a_124_375# 0.012574f
C16317 net68 vdd 1.026897f
C16318 _273_/a_36_68# _128_ 0.005719f
C16319 FILLER_0_14_50/a_124_375# _181_ 0.00402f
C16320 fanout68/a_36_113# net50 0.020067f
C16321 FILLER_0_18_2/a_484_472# _452_/a_2225_156# 0.019521f
C16322 net29 FILLER_0_16_255/a_124_375# 0.085055f
C16323 _424_/a_2248_156# FILLER_0_21_60/a_572_375# 0.030666f
C16324 _424_/a_2665_112# FILLER_0_21_60/a_124_375# 0.010688f
C16325 output28/a_224_472# result[1] 0.054333f
C16326 FILLER_0_15_290/a_36_472# result[3] 0.014709f
C16327 _445_/a_2560_156# net17 0.010829f
C16328 FILLER_0_20_193/a_36_472# FILLER_0_19_187/a_572_375# 0.001543f
C16329 _428_/a_2248_156# net74 0.072805f
C16330 _421_/a_448_472# _010_ 0.039422f
C16331 _430_/a_2560_156# _092_ 0.001333f
C16332 output37/a_224_472# _425_/a_2665_112# 0.022027f
C16333 net69 fanout49/a_36_160# 0.005942f
C16334 FILLER_0_10_78/a_572_375# net52 0.003311f
C16335 _103_ _288_/a_224_472# 0.002992f
C16336 net55 FILLER_0_18_76/a_36_472# 0.003695f
C16337 FILLER_0_3_54/a_36_472# _164_ 0.012512f
C16338 _414_/a_1204_472# _074_ 0.003142f
C16339 FILLER_0_15_150/a_36_472# fanout53/a_36_160# 0.002059f
C16340 trim_val\[4\] _163_ 0.03439f
C16341 net55 _423_/a_2248_156# 0.001188f
C16342 _430_/a_36_151# _138_ 0.001123f
C16343 _253_/a_36_68# cal_itt\[0\] 0.001495f
C16344 _425_/a_796_472# vdd 0.002206f
C16345 net20 FILLER_0_12_220/a_1020_375# 0.047331f
C16346 FILLER_0_9_282/a_36_472# vss 0.002224f
C16347 FILLER_0_14_50/a_36_472# _174_ 0.015387f
C16348 output45/a_224_472# net40 0.001284f
C16349 mask\[7\] _435_/a_2248_156# 0.026974f
C16350 net70 FILLER_0_14_107/a_572_375# 0.018214f
C16351 _071_ _121_ 0.007734f
C16352 vss FILLER_0_22_107/a_484_472# 0.003617f
C16353 net34 net80 0.041846f
C16354 FILLER_0_15_212/a_484_472# mask\[1\] 0.007258f
C16355 net73 FILLER_0_17_133/a_36_472# 0.049294f
C16356 _070_ FILLER_0_10_94/a_572_375# 0.009837f
C16357 _050_ _436_/a_796_472# 0.007055f
C16358 FILLER_0_16_57/a_1468_375# _131_ 0.015859f
C16359 cal_count\[3\] FILLER_0_12_196/a_36_472# 0.079338f
C16360 output34/a_224_472# _102_ 0.008577f
C16361 net58 _412_/a_1204_472# 0.018724f
C16362 _426_/a_2248_156# _060_ 0.00106f
C16363 _257_/a_36_472# _053_ 0.00507f
C16364 _117_ vss 0.048946f
C16365 _174_ cal_count\[3\] 0.053844f
C16366 output31/a_224_472# _103_ 0.006731f
C16367 _333_/a_36_160# vdd 0.107883f
C16368 _189_/a_67_603# FILLER_0_13_228/a_124_375# 0.00744f
C16369 _320_/a_36_472# vdd 0.086964f
C16370 FILLER_0_4_107/a_484_472# _153_ 0.026082f
C16371 FILLER_0_4_107/a_1380_472# _154_ 0.005297f
C16372 _208_/a_36_160# vdd 0.014709f
C16373 _113_ _060_ 0.01991f
C16374 FILLER_0_5_206/a_36_472# _122_ 0.003017f
C16375 mask\[5\] _201_/a_67_603# 0.001222f
C16376 FILLER_0_20_15/a_932_472# vdd 0.002617f
C16377 _442_/a_36_151# _158_ 0.001257f
C16378 mask\[9\] _438_/a_36_151# 0.060632f
C16379 FILLER_0_15_142/a_36_472# _095_ 0.001526f
C16380 net16 FILLER_0_6_37/a_124_375# 0.010358f
C16381 FILLER_0_18_209/a_572_375# _201_/a_67_603# 0.008812f
C16382 FILLER_0_3_172/a_572_375# net22 0.013048f
C16383 FILLER_0_15_72/a_484_472# _451_/a_3129_107# 0.005866f
C16384 FILLER_0_13_65/a_36_472# fanout72/a_36_113# 0.193651f
C16385 _072_ state\[1\] 0.267762f
C16386 FILLER_0_18_2/a_36_472# net44 0.011079f
C16387 net75 _425_/a_796_472# 0.001146f
C16388 FILLER_0_4_177/a_484_472# _087_ 0.005486f
C16389 net79 _416_/a_796_472# 0.01137f
C16390 _322_/a_692_472# _070_ 0.002328f
C16391 _305_/a_36_159# net37 0.015682f
C16392 _128_ _129_ 0.029628f
C16393 FILLER_0_8_247/a_1020_375# vdd -0.002559f
C16394 FILLER_0_14_91/a_124_375# net53 0.065572f
C16395 net76 FILLER_0_2_177/a_572_375# 0.053951f
C16396 _016_ FILLER_0_12_124/a_36_472# 0.002661f
C16397 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_572_375# 0.086635f
C16398 _363_/a_36_68# _163_ 0.005627f
C16399 _057_ _069_ 0.053765f
C16400 _421_/a_36_151# vss 0.021759f
C16401 _421_/a_448_472# vdd 0.030898f
C16402 FILLER_0_6_239/a_36_472# fanout75/a_36_113# 0.00191f
C16403 FILLER_0_15_142/a_484_472# _095_ 0.001509f
C16404 _132_ FILLER_0_14_107/a_572_375# 0.007439f
C16405 net23 FILLER_0_22_128/a_1380_472# 0.0019f
C16406 _028_ _439_/a_36_151# 0.009268f
C16407 FILLER_0_13_212/a_1380_472# FILLER_0_13_228/a_36_472# 0.013277f
C16408 FILLER_0_14_107/a_484_472# _043_ 0.001641f
C16409 output43/a_224_472# trimb[2] 0.005445f
C16410 _225_/a_36_160# vss 0.003244f
C16411 FILLER_0_23_88/a_124_375# _437_/a_36_151# 0.002709f
C16412 _448_/a_2665_112# _037_ 0.042225f
C16413 net55 _067_ 0.053438f
C16414 output34/a_224_472# _198_/a_67_603# 0.00179f
C16415 _427_/a_2248_156# net36 0.004462f
C16416 FILLER_0_20_193/a_484_472# vss 0.002439f
C16417 ctln[2] net5 0.001249f
C16418 _118_ _060_ 0.002868f
C16419 FILLER_0_9_28/a_1020_375# vdd 0.033815f
C16420 fanout54/a_36_160# _145_ 0.009257f
C16421 _446_/a_448_472# net40 0.05302f
C16422 net75 _253_/a_672_68# 0.003771f
C16423 _274_/a_2960_68# _091_ 0.001338f
C16424 trim_mask\[2\] _030_ 1.467465f
C16425 _053_ FILLER_0_7_59/a_124_375# 0.015298f
C16426 net73 _022_ 0.003246f
C16427 _178_ net17 0.115251f
C16428 net2 clk 0.046099f
C16429 FILLER_0_5_198/a_484_472# net59 0.059394f
C16430 _210_/a_67_603# vdd 0.028101f
C16431 _345_/a_36_160# FILLER_0_19_125/a_36_472# 0.006647f
C16432 mask\[3\] _099_ 0.10534f
C16433 FILLER_0_17_104/a_1468_375# FILLER_0_16_115/a_124_375# 0.026339f
C16434 net60 _007_ 0.025806f
C16435 FILLER_0_18_139/a_1380_472# vss 0.009272f
C16436 mask\[5\] FILLER_0_19_187/a_36_472# 0.007596f
C16437 _447_/a_448_472# net68 0.012962f
C16438 net49 _440_/a_2560_156# 0.011378f
C16439 _064_ _445_/a_448_472# 0.080931f
C16440 _431_/a_36_151# fanout70/a_36_113# 0.016241f
C16441 net79 FILLER_0_11_282/a_124_375# 0.002239f
C16442 _152_ _062_ 0.097086f
C16443 _091_ _097_ 0.036863f
C16444 net64 FILLER_0_15_235/a_484_472# 0.005893f
C16445 FILLER_0_16_154/a_1468_375# vss 0.002071f
C16446 FILLER_0_16_154/a_36_472# vdd 0.00225f
C16447 _431_/a_36_151# FILLER_0_18_107/a_2724_472# 0.00271f
C16448 trim_mask\[4\] _031_ 0.001262f
C16449 FILLER_0_7_162/a_124_375# _169_ 0.00336f
C16450 FILLER_0_15_235/a_484_472# mask\[1\] 0.014415f
C16451 _116_ net4 0.00603f
C16452 mask\[7\] FILLER_0_22_128/a_2276_472# 0.004398f
C16453 output41/a_224_472# trim[3] 0.042209f
C16454 net75 FILLER_0_8_247/a_1020_375# 0.009573f
C16455 result[9] FILLER_0_24_274/a_124_375# 0.008195f
C16456 trimb[1] net43 0.004299f
C16457 trimb[1] output44/a_224_472# 0.046391f
C16458 cal clk 0.033015f
C16459 net80 mask\[2\] 0.048734f
C16460 _119_ FILLER_0_8_138/a_124_375# 0.006523f
C16461 _088_ net22 0.17798f
C16462 FILLER_0_7_104/a_1468_375# vdd 0.026224f
C16463 _095_ _113_ 0.004037f
C16464 net73 FILLER_0_18_107/a_36_472# 0.002425f
C16465 FILLER_0_7_72/a_1380_472# net50 0.077411f
C16466 output32/a_224_472# _419_/a_36_151# 0.129117f
C16467 net26 FILLER_0_21_28/a_1916_375# 0.008721f
C16468 FILLER_0_18_107/a_2364_375# vdd 0.017472f
C16469 _251_/a_244_472# net4 0.005273f
C16470 net39 _445_/a_2560_156# 0.003401f
C16471 _317_/a_36_113# FILLER_0_7_233/a_36_472# 0.003531f
C16472 net52 FILLER_0_9_72/a_1468_375# 0.003576f
C16473 trim_mask\[3\] vss 0.156544f
C16474 _217_/a_36_160# _052_ 0.016695f
C16475 net54 net23 0.084191f
C16476 net58 _412_/a_1000_472# 0.030238f
C16477 net54 FILLER_0_22_128/a_1916_375# 0.001933f
C16478 FILLER_0_18_139/a_124_375# _145_ 0.00346f
C16479 FILLER_0_18_37/a_1468_375# vss 0.054381f
C16480 FILLER_0_18_37/a_36_472# vdd 0.136723f
C16481 net67 vss 0.435869f
C16482 FILLER_0_16_89/a_1020_375# vdd 0.007416f
C16483 ctln[2] FILLER_0_1_266/a_572_375# 0.012126f
C16484 _320_/a_36_472# FILLER_0_13_206/a_36_472# 0.038251f
C16485 _131_ FILLER_0_17_64/a_36_472# 0.002638f
C16486 _010_ _419_/a_36_151# 0.002099f
C16487 FILLER_0_24_274/a_36_472# vss 0.001013f
C16488 FILLER_0_24_274/a_484_472# vdd 0.004641f
C16489 output39/a_224_472# _054_ 0.002121f
C16490 net39 _221_/a_36_160# 0.059979f
C16491 FILLER_0_9_28/a_484_472# net40 0.020293f
C16492 _178_ FILLER_0_16_37/a_36_472# 0.007425f
C16493 net57 _128_ 0.040656f
C16494 output12/a_224_472# ctln[5] 0.069673f
C16495 _087_ _079_ 0.251042f
C16496 _242_/a_36_160# _066_ 0.044262f
C16497 _065_ trim_val\[3\] 1.235816f
C16498 _122_ _123_ 0.242965f
C16499 _062_ net21 0.025648f
C16500 trim_mask\[1\] _154_ 0.004835f
C16501 _053_ _359_/a_36_488# 0.015831f
C16502 _053_ _078_ 0.137388f
C16503 _055_ _223_/a_36_160# 0.012271f
C16504 _011_ _422_/a_36_151# 0.015698f
C16505 mask\[3\] FILLER_0_17_218/a_36_472# 0.015535f
C16506 _000_ FILLER_0_3_221/a_1468_375# 0.054354f
C16507 _025_ FILLER_0_22_107/a_572_375# 0.090334f
C16508 result[9] FILLER_0_23_274/a_124_375# 0.003102f
C16509 _148_ FILLER_0_22_107/a_484_472# 0.004761f
C16510 _091_ FILLER_0_15_180/a_124_375# 0.001415f
C16511 net20 FILLER_0_3_221/a_572_375# 0.004331f
C16512 cal_count\[2\] _401_/a_36_68# 0.008136f
C16513 trim_mask\[4\] _371_/a_36_113# 0.007529f
C16514 _032_ _159_ 0.053405f
C16515 FILLER_0_10_37/a_36_472# vdd 0.141896f
C16516 FILLER_0_10_37/a_124_375# vss 0.006228f
C16517 _408_/a_1936_472# vdd 0.022538f
C16518 _413_/a_36_151# FILLER_0_3_172/a_2812_375# 0.059049f
C16519 output22/a_224_472# _435_/a_448_472# 0.010723f
C16520 output21/a_224_472# output19/a_224_472# 0.007877f
C16521 _070_ _062_ 0.06973f
C16522 FILLER_0_9_28/a_1468_375# net51 0.00111f
C16523 calibrate _120_ 0.001106f
C16524 _184_ vdd 0.202732f
C16525 output26/a_224_472# FILLER_0_23_44/a_36_472# 0.026108f
C16526 _379_/a_36_472# _166_ 0.038062f
C16527 _126_ FILLER_0_11_142/a_36_472# 0.001428f
C16528 output43/a_224_472# net40 0.014984f
C16529 FILLER_0_18_209/a_484_472# vss 0.005794f
C16530 _101_ vdd 0.02756f
C16531 net18 _416_/a_448_472# 0.05521f
C16532 _114_ _428_/a_36_151# 0.008132f
C16533 _069_ cal_count\[3\] 0.012382f
C16534 _242_/a_36_160# net37 0.02401f
C16535 net50 net40 0.005105f
C16536 net47 _385_/a_36_68# 0.011168f
C16537 net54 _025_ 0.00573f
C16538 _094_ net77 0.00405f
C16539 FILLER_0_3_78/a_36_472# _160_ 0.006564f
C16540 FILLER_0_12_220/a_1020_375# vss 0.004698f
C16541 FILLER_0_12_220/a_1468_375# vdd 0.002801f
C16542 output13/a_224_472# _448_/a_2665_112# 0.027303f
C16543 FILLER_0_7_72/a_2276_472# _053_ 0.016004f
C16544 FILLER_0_15_142/a_36_472# net74 0.003166f
C16545 net72 FILLER_0_18_37/a_36_472# 0.043427f
C16546 net55 FILLER_0_18_37/a_572_375# 0.007169f
C16547 FILLER_0_4_107/a_36_472# _160_ 0.009073f
C16548 _426_/a_2248_156# net64 0.01109f
C16549 result[7] _420_/a_2560_156# 0.001179f
C16550 FILLER_0_18_2/a_2724_472# net47 0.001551f
C16551 net20 _000_ 0.159624f
C16552 FILLER_0_17_72/a_124_375# vss 0.048053f
C16553 FILLER_0_17_72/a_572_375# vdd 0.002455f
C16554 FILLER_0_8_37/a_36_472# vdd 0.135405f
C16555 FILLER_0_8_37/a_572_375# vss 0.00282f
C16556 net47 FILLER_0_4_91/a_36_472# 0.005186f
C16557 _121_ net23 0.078786f
C16558 _072_ FILLER_0_7_233/a_124_375# 0.002279f
C16559 _053_ FILLER_0_6_90/a_124_375# 0.003061f
C16560 _105_ _109_ 0.107328f
C16561 net27 FILLER_0_10_256/a_36_472# 0.008331f
C16562 _061_ _311_/a_3740_473# 0.006728f
C16563 mask\[1\] _113_ 0.032744f
C16564 FILLER_0_9_28/a_1828_472# vdd 0.006263f
C16565 FILLER_0_13_100/a_124_375# vdd 0.039324f
C16566 FILLER_0_16_107/a_572_375# vdd 0.019922f
C16567 net38 _450_/a_448_472# 0.031891f
C16568 _419_/a_36_151# vdd -0.110366f
C16569 net57 _386_/a_1084_68# 0.005716f
C16570 _072_ vdd 0.715894f
C16571 _449_/a_2560_156# _038_ 0.010532f
C16572 net80 FILLER_0_22_177/a_1020_375# 0.00258f
C16573 trim[0] FILLER_0_3_2/a_36_472# 0.017429f
C16574 FILLER_0_15_59/a_572_375# vdd 0.03104f
C16575 FILLER_0_15_59/a_124_375# vss 0.003806f
C16576 fanout57/a_36_113# net57 0.004316f
C16577 _004_ _415_/a_1000_472# 0.005004f
C16578 _091_ _019_ 0.031681f
C16579 _326_/a_36_160# _062_ 0.007797f
C16580 _392_/a_36_68# _067_ 0.020085f
C16581 FILLER_0_17_72/a_1828_472# _136_ 0.004161f
C16582 net73 net53 0.094507f
C16583 net34 _106_ 0.013009f
C16584 FILLER_0_7_59/a_484_472# net68 0.002785f
C16585 fanout69/a_36_113# _371_/a_36_113# 0.259508f
C16586 _348_/a_257_69# mask\[6\] 0.00159f
C16587 net7 _065_ 0.0295f
C16588 result[7] _421_/a_1456_156# 0.001009f
C16589 FILLER_0_18_107/a_124_375# FILLER_0_20_107/a_36_472# 0.00108f
C16590 net70 vdd 0.858299f
C16591 _093_ _069_ 0.008325f
C16592 FILLER_0_17_200/a_124_375# FILLER_0_18_177/a_2724_472# 0.001597f
C16593 net74 FILLER_0_13_142/a_484_472# 0.001771f
C16594 _404_/a_36_472# _041_ 0.003068f
C16595 net73 _431_/a_2665_112# 0.001495f
C16596 FILLER_0_1_98/a_36_472# trim_mask\[3\] 0.106084f
C16597 FILLER_0_15_142/a_572_375# vdd -0.013698f
C16598 FILLER_0_9_28/a_2364_375# trim_val\[0\] 0.006639f
C16599 _116_ net79 0.081785f
C16600 net47 vdd 2.422992f
C16601 FILLER_0_1_266/a_124_375# net19 0.007016f
C16602 net62 _195_/a_67_603# 0.002422f
C16603 FILLER_0_7_195/a_36_472# _055_ 0.03271f
C16604 _437_/a_448_472# vss 0.001524f
C16605 _437_/a_1308_423# vdd 0.005139f
C16606 _441_/a_2248_156# _164_ 0.040396f
C16607 trim_val\[2\] _164_ 0.005847f
C16608 net47 _365_/a_244_472# 0.001431f
C16609 trim_mask\[4\] FILLER_0_2_111/a_1468_375# 0.001226f
C16610 _177_ fanout55/a_36_160# 0.002687f
C16611 FILLER_0_21_125/a_124_375# _022_ 0.007023f
C16612 _098_ FILLER_0_15_205/a_36_472# 0.010528f
C16613 ctln[1] rstn 0.62944f
C16614 _074_ FILLER_0_3_221/a_1380_472# 0.001341f
C16615 net26 net55 0.002901f
C16616 net15 _440_/a_796_472# 0.005848f
C16617 _415_/a_2248_156# net18 0.057604f
C16618 net54 _436_/a_1000_472# 0.002051f
C16619 output25/a_224_472# net35 0.016177f
C16620 net62 net30 0.339141f
C16621 vss result[3] 0.28152f
C16622 FILLER_0_16_73/a_484_472# _175_ 0.036868f
C16623 result[4] net79 0.048452f
C16624 _446_/a_36_151# net66 0.034846f
C16625 _242_/a_36_160# FILLER_0_5_148/a_484_472# 0.003699f
C16626 _064_ _446_/a_2248_156# 0.04774f
C16627 net80 _339_/a_36_160# 0.016897f
C16628 _112_ _316_/a_692_472# 0.001614f
C16629 net35 net22 0.001381f
C16630 FILLER_0_23_44/a_1468_375# vdd -0.013698f
C16631 _125_ _120_ 0.006198f
C16632 _077_ _453_/a_1308_423# 0.071515f
C16633 _236_/a_36_160# FILLER_0_8_2/a_36_472# 0.01395f
C16634 FILLER_0_16_107/a_484_472# _040_ 0.003828f
C16635 FILLER_0_4_197/a_1020_375# net76 0.006026f
C16636 FILLER_0_18_107/a_932_472# FILLER_0_16_115/a_124_375# 0.001512f
C16637 FILLER_0_5_72/a_572_375# _029_ 0.010208f
C16638 _091_ _429_/a_2248_156# 0.006148f
C16639 FILLER_0_6_47/a_124_375# vdd 0.008011f
C16640 net72 FILLER_0_15_59/a_572_375# 0.00799f
C16641 fanout63/a_36_160# net36 0.004435f
C16642 ctln[8] ctln[9] 0.003265f
C16643 mask\[5\] net23 0.002188f
C16644 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1468_375# 0.086635f
C16645 _321_/a_170_472# _126_ 0.018831f
C16646 net32 _048_ 0.008647f
C16647 net16 _052_ 0.022236f
C16648 _340_/a_36_160# mask\[6\] 0.010151f
C16649 net63 FILLER_0_20_193/a_36_472# 0.048818f
C16650 _372_/a_3662_472# net23 0.002864f
C16651 _132_ vdd 0.960634f
C16652 _144_ FILLER_0_22_128/a_3172_472# 0.001287f
C16653 _098_ _433_/a_2665_112# 0.01601f
C16654 FILLER_0_7_104/a_572_375# _154_ 0.020664f
C16655 _057_ _090_ 0.112325f
C16656 FILLER_0_4_152/a_124_375# _170_ 0.029927f
C16657 _257_/a_36_472# cal_itt\[3\] 0.136487f
C16658 net17 _450_/a_2225_156# 0.033342f
C16659 FILLER_0_9_60/a_124_375# vdd 0.005798f
C16660 net47 _452_/a_1040_527# 0.014695f
C16661 net41 _444_/a_1000_472# 0.002179f
C16662 net27 output28/a_224_472# 0.011692f
C16663 net26 _424_/a_796_472# 0.006496f
C16664 FILLER_0_15_290/a_124_375# vdd 0.028723f
C16665 FILLER_0_7_72/a_2276_472# _028_ 0.001777f
C16666 _174_ _120_ 0.002521f
C16667 _136_ FILLER_0_16_115/a_36_472# 0.013477f
C16668 _065_ net15 0.065255f
C16669 FILLER_0_4_144/a_36_472# trim_mask\[4\] 0.017557f
C16670 _226_/a_860_68# net21 0.00107f
C16671 FILLER_0_8_127/a_36_472# vdd 0.069117f
C16672 fanout69/a_36_113# FILLER_0_2_111/a_1468_375# 0.015816f
C16673 _322_/a_124_24# _128_ 0.02077f
C16674 _028_ FILLER_0_6_90/a_124_375# 0.012573f
C16675 _058_ FILLER_0_9_105/a_484_472# 0.00148f
C16676 _057_ net22 0.163773f
C16677 net74 _118_ 0.060991f
C16678 _112_ net76 0.011948f
C16679 _397_/a_36_472# net36 0.010045f
C16680 _282_/a_36_160# vdd 0.010099f
C16681 output47/a_224_472# net17 0.081437f
C16682 _408_/a_1936_472# cal_count\[0\] 0.001434f
C16683 FILLER_0_12_136/a_572_375# _127_ 0.00116f
C16684 _093_ FILLER_0_17_104/a_36_472# 0.014431f
C16685 net5 cal_itt\[1\] 0.057623f
C16686 _438_/a_2665_112# FILLER_0_19_111/a_36_472# 0.007491f
C16687 _106_ mask\[2\] 0.039965f
C16688 FILLER_0_17_282/a_124_375# vdd 0.004586f
C16689 _448_/a_448_472# vdd 0.02042f
C16690 valid output37/a_224_472# 0.039402f
C16691 _077_ _074_ 0.148596f
C16692 _114_ _085_ 0.056448f
C16693 _053_ FILLER_0_9_28/a_2276_472# 0.002243f
C16694 _315_/a_1229_68# _121_ 0.003401f
C16695 _398_/a_36_113# _278_/a_36_160# 0.001636f
C16696 _411_/a_448_472# ctln[3] 0.00336f
C16697 _430_/a_2665_112# net36 0.003477f
C16698 FILLER_0_14_107/a_124_375# vss 0.002674f
C16699 net55 FILLER_0_17_38/a_36_472# 0.010728f
C16700 cal_count\[2\] FILLER_0_15_10/a_124_375# 0.017594f
C16701 FILLER_0_14_107/a_572_375# vdd 0.021509f
C16702 _059_ vss 0.714648f
C16703 _063_ FILLER_0_6_37/a_124_375# 0.012149f
C16704 FILLER_0_22_177/a_124_375# vss 0.002674f
C16705 FILLER_0_22_177/a_572_375# vdd -0.003694f
C16706 output48/a_224_472# vss 0.006655f
C16707 net15 fanout51/a_36_113# 0.001562f
C16708 FILLER_0_21_133/a_124_375# vdd 0.010519f
C16709 net81 net2 1.204674f
C16710 sample net5 0.359975f
C16711 net4 FILLER_0_12_220/a_1020_375# 0.020782f
C16712 net66 FILLER_0_5_54/a_124_375# 0.002093f
C16713 FILLER_0_7_104/a_572_375# _058_ 0.006125f
C16714 mask\[5\] net33 0.251971f
C16715 net36 FILLER_0_15_212/a_572_375# 0.004606f
C16716 FILLER_0_3_221/a_572_375# vss 0.003292f
C16717 _000_ cal_itt\[1\] 0.012692f
C16718 _375_/a_36_68# vss 0.02182f
C16719 net5 vss 0.326032f
C16720 mask\[4\] FILLER_0_18_177/a_2276_472# 0.016876f
C16721 _261_/a_36_160# FILLER_0_5_148/a_36_472# 0.195478f
C16722 fanout66/a_36_113# vdd 0.049012f
C16723 FILLER_0_18_107/a_2364_375# _433_/a_36_151# 0.002106f
C16724 FILLER_0_5_54/a_1020_375# _029_ 0.024737f
C16725 _093_ _438_/a_36_151# 0.088469f
C16726 _440_/a_2560_156# net47 0.003888f
C16727 trim[4] net38 0.095379f
C16728 FILLER_0_16_107/a_36_472# net14 0.004691f
C16729 _119_ FILLER_0_8_156/a_36_472# 0.010504f
C16730 net35 FILLER_0_22_86/a_36_472# 0.00797f
C16731 mask\[8\] FILLER_0_22_86/a_484_472# 0.012439f
C16732 _031_ _157_ 0.104339f
C16733 _412_/a_448_472# net81 0.047334f
C16734 net52 _442_/a_1000_472# 0.016308f
C16735 _020_ _431_/a_1204_472# 0.002176f
C16736 net62 FILLER_0_14_263/a_36_472# 0.019591f
C16737 _054_ net40 0.072879f
C16738 net57 net14 0.05113f
C16739 FILLER_0_15_235/a_124_375# FILLER_0_14_235/a_124_375# 0.05841f
C16740 FILLER_0_15_150/a_124_375# fanout53/a_36_160# 0.004079f
C16741 net78 _420_/a_2665_112# 0.039469f
C16742 _276_/a_36_160# _106_ 0.009097f
C16743 net52 trim_mask\[1\] 0.04149f
C16744 _219_/a_36_160# net14 0.048037f
C16745 _449_/a_2248_156# net74 0.004565f
C16746 _000_ vss 0.205593f
C16747 _186_ _180_ 0.003034f
C16748 FILLER_0_18_177/a_1916_375# vdd 0.021f
C16749 _083_ _082_ 0.018442f
C16750 net27 calibrate 0.017426f
C16751 FILLER_0_9_223/a_124_375# _076_ 0.004399f
C16752 FILLER_0_4_107/a_36_472# _156_ 0.005297f
C16753 FILLER_0_12_28/a_36_472# _450_/a_3129_107# 0.009814f
C16754 ctln[5] _448_/a_2248_156# 0.004396f
C16755 _122_ _242_/a_36_160# 0.005377f
C16756 _192_/a_67_603# _044_ 0.002571f
C16757 _131_ _135_ 0.068855f
C16758 _131_ FILLER_0_17_56/a_484_472# 0.002672f
C16759 _136_ _451_/a_2449_156# 0.004653f
C16760 FILLER_0_14_91/a_36_472# vss 0.001729f
C16761 FILLER_0_14_91/a_484_472# vdd 0.00605f
C16762 _119_ _319_/a_234_472# 0.004559f
C16763 _057_ _076_ 0.041986f
C16764 state\[1\] vdd 0.544231f
C16765 FILLER_0_5_117/a_36_472# _153_ 0.028773f
C16766 _141_ FILLER_0_18_139/a_1380_472# 0.016119f
C16767 FILLER_0_18_2/a_932_472# vdd 0.002342f
C16768 net15 FILLER_0_13_72/a_36_472# 0.006713f
C16769 net15 net51 0.191328f
C16770 _415_/a_36_151# net19 0.05689f
C16771 _453_/a_2248_156# vss 0.031525f
C16772 _453_/a_2665_112# vdd 0.005481f
C16773 _092_ vdd 0.140213f
C16774 FILLER_0_16_57/a_932_472# net15 0.037807f
C16775 net57 net82 0.91473f
C16776 _417_/a_1000_472# _006_ 0.026299f
C16777 net69 FILLER_0_3_78/a_572_375# 0.002984f
C16778 _072_ _374_/a_36_68# 0.061028f
C16779 _012_ FILLER_0_21_60/a_36_472# 0.017483f
C16780 mask\[3\] FILLER_0_16_154/a_932_472# 0.002604f
C16781 FILLER_0_13_212/a_1468_375# FILLER_0_12_220/a_572_375# 0.05841f
C16782 net81 FILLER_0_12_236/a_572_375# 0.021025f
C16783 net69 FILLER_0_2_101/a_36_472# 0.00845f
C16784 output32/a_224_472# _010_ 0.001508f
C16785 _144_ _346_/a_257_69# 0.001089f
C16786 _408_/a_728_93# _181_ 0.018292f
C16787 FILLER_0_4_123/a_36_472# _152_ 0.003937f
C16788 _414_/a_1000_472# _003_ 0.002053f
C16789 _074_ net37 0.064705f
C16790 FILLER_0_11_101/a_484_472# cal_count\[3\] 0.00702f
C16791 FILLER_0_20_2/a_572_375# vss 0.001471f
C16792 FILLER_0_20_2/a_36_472# vdd 0.102471f
C16793 _176_ _394_/a_718_524# 0.00141f
C16794 cal_count\[3\] _090_ 0.243462f
C16795 FILLER_0_5_212/a_36_472# vss 0.00578f
C16796 FILLER_0_18_177/a_3172_472# net21 0.010321f
C16797 FILLER_0_4_197/a_1468_375# net76 0.007667f
C16798 FILLER_0_4_177/a_124_375# _163_ 0.004052f
C16799 _444_/a_796_472# net67 0.006859f
C16800 net53 _427_/a_1308_423# 0.007426f
C16801 FILLER_0_5_128/a_572_375# _133_ 0.00134f
C16802 FILLER_0_12_236/a_572_375# _060_ 0.001597f
C16803 trim_val\[1\] vss 0.029927f
C16804 FILLER_0_1_266/a_36_472# vdd 0.008551f
C16805 FILLER_0_1_266/a_572_375# vss 0.001919f
C16806 _414_/a_1000_472# net21 0.042244f
C16807 _407_/a_36_472# _184_ 0.004667f
C16808 _089_ _002_ 0.002349f
C16809 cal_itt\[3\] _078_ 0.024443f
C16810 net18 FILLER_0_9_282/a_124_375# 0.024657f
C16811 _231_/a_652_68# _062_ 0.001555f
C16812 _083_ _265_/a_244_68# 0.004022f
C16813 _151_ _153_ 0.027868f
C16814 net32 result[9] 0.001371f
C16815 _078_ _081_ 0.445443f
C16816 _413_/a_2248_156# FILLER_0_3_212/a_124_375# 0.030666f
C16817 _008_ _418_/a_1000_472# 0.01006f
C16818 cal_count\[2\] _278_/a_36_160# 0.023061f
C16819 _112_ _083_ 0.003571f
C16820 _104_ _093_ 0.109158f
C16821 _450_/a_2225_156# _039_ 0.034731f
C16822 net80 vss 0.347557f
C16823 mask\[9\] _140_ 0.00126f
C16824 net1 net18 0.047886f
C16825 net65 output27/a_224_472# 0.019729f
C16826 FILLER_0_12_2/a_572_375# net38 0.00609f
C16827 ctln[2] en 0.001355f
C16828 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1468_375# 0.086742f
C16829 _370_/a_124_24# _160_ 0.001126f
C16830 FILLER_0_21_206/a_36_472# net22 0.012952f
C16831 trimb[1] _452_/a_2449_156# 0.001681f
C16832 FILLER_0_10_78/a_572_375# FILLER_0_11_78/a_572_375# 0.05841f
C16833 output24/a_224_472# _436_/a_36_151# 0.053592f
C16834 FILLER_0_12_136/a_1468_375# vss 0.043987f
C16835 _402_/a_718_527# vdd 0.020893f
C16836 FILLER_0_17_142/a_124_375# _137_ 0.006974f
C16837 _412_/a_36_151# net18 0.011383f
C16838 _308_/a_848_380# _070_ 0.033275f
C16839 _069_ _120_ 0.030804f
C16840 net34 _144_ 0.029247f
C16841 _304_/a_224_472# vss 0.001746f
C16842 _423_/a_1000_472# _012_ 0.013415f
C16843 net73 FILLER_0_19_111/a_484_472# 0.007404f
C16844 _106_ net20 0.050151f
C16845 FILLER_0_21_286/a_124_375# _420_/a_36_151# 0.001597f
C16846 _413_/a_1204_472# net65 0.017514f
C16847 _274_/a_36_68# _072_ 0.001647f
C16848 output32/a_224_472# vdd 0.082664f
C16849 net57 _098_ 0.062604f
C16850 FILLER_0_19_111/a_124_375# vdd 0.005128f
C16851 net79 FILLER_0_12_220/a_1020_375# 0.010818f
C16852 _168_ vss 0.171346f
C16853 output26/a_224_472# vss 0.0137f
C16854 net65 net22 0.374917f
C16855 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1380_472# 0.013276f
C16856 net62 _417_/a_2665_112# 0.006083f
C16857 fanout67/a_36_160# trim_val\[0\] 0.003096f
C16858 _144_ _354_/a_49_472# 0.03742f
C16859 _431_/a_36_151# _093_ 0.004862f
C16860 fanout51/a_36_113# FILLER_0_11_78/a_36_472# 0.193759f
C16861 _119_ _359_/a_36_488# 0.003263f
C16862 mask\[7\] FILLER_0_22_177/a_124_375# 0.001315f
C16863 _424_/a_2560_156# _012_ 0.002513f
C16864 mask\[4\] _093_ 0.469687f
C16865 _093_ net22 0.041918f
C16866 _113_ FILLER_0_15_180/a_124_375# 0.001512f
C16867 _051_ vdd 0.036931f
C16868 FILLER_0_4_152/a_36_472# net47 0.007541f
C16869 cal_count\[3\] _038_ 0.682941f
C16870 _126_ _135_ 0.011447f
C16871 ctlp[4] net33 0.001734f
C16872 FILLER_0_18_53/a_484_472# vss 0.003579f
C16873 output38/a_224_472# vdd -0.006652f
C16874 FILLER_0_17_161/a_36_472# _137_ 0.013985f
C16875 FILLER_0_18_76/a_572_375# _438_/a_36_151# 0.059049f
C16876 net35 FILLER_0_22_177/a_1380_472# 0.01447f
C16877 _104_ FILLER_0_17_226/a_36_472# 0.013926f
C16878 _010_ vdd 0.121474f
C16879 _247_/a_36_160# vss 0.009308f
C16880 FILLER_0_5_181/a_124_375# vdd 0.009553f
C16881 FILLER_0_21_28/a_572_375# vdd 0.013051f
C16882 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1468_375# 0.086635f
C16883 net23 _348_/a_49_472# 0.0037f
C16884 net38 net17 1.634286f
C16885 FILLER_0_3_172/a_3260_375# vdd -0.013516f
C16886 _052_ FILLER_0_21_28/a_3260_375# 0.002388f
C16887 FILLER_0_16_241/a_124_375# net30 0.028559f
C16888 _239_/a_36_160# net68 0.043367f
C16889 FILLER_0_5_128/a_484_472# _152_ 0.002283f
C16890 net4 FILLER_0_3_221/a_572_375# 0.030599f
C16891 FILLER_0_5_117/a_124_375# _160_ 0.008534f
C16892 fanout75/a_36_113# net1 0.011428f
C16893 FILLER_0_11_64/a_124_375# _453_/a_2248_156# 0.001901f
C16894 FILLER_0_13_212/a_484_472# _043_ 0.011439f
C16895 _385_/a_36_68# vdd 0.01625f
C16896 _129_ _372_/a_170_472# 0.001985f
C16897 _093_ FILLER_0_18_107/a_1380_472# 0.001782f
C16898 net4 net5 0.104296f
C16899 _029_ _156_ 0.018258f
C16900 _131_ _129_ 0.017222f
C16901 _088_ FILLER_0_3_172/a_2276_472# 0.024532f
C16902 _035_ net40 0.068572f
C16903 FILLER_0_12_2/a_484_472# vss 0.001748f
C16904 net73 _431_/a_796_472# 0.002306f
C16905 net22 net59 0.195226f
C16906 _173_ _450_/a_3129_107# 0.00264f
C16907 mask\[9\] _149_ 0.040342f
C16908 _132_ _433_/a_36_151# 0.024768f
C16909 _098_ FILLER_0_15_212/a_1380_472# 0.009972f
C16910 _444_/a_1308_423# net47 0.040252f
C16911 state\[0\] _055_ 0.042917f
C16912 FILLER_0_18_2/a_2724_472# vdd 0.004348f
C16913 _442_/a_36_151# net69 0.048683f
C16914 net52 _164_ 0.313379f
C16915 _005_ _416_/a_796_472# 0.009162f
C16916 _036_ net49 0.005235f
C16917 _053_ FILLER_0_7_104/a_1020_375# 0.002671f
C16918 vss FILLER_0_4_91/a_572_375# 0.055113f
C16919 _447_/a_2560_156# net69 0.001774f
C16920 FILLER_0_4_99/a_36_472# net47 0.003903f
C16921 FILLER_0_7_59/a_124_375# FILLER_0_6_47/a_1468_375# 0.05841f
C16922 output35/a_224_472# net22 0.028095f
C16923 output36/a_224_472# vdd 0.145046f
C16924 _445_/a_2665_112# net49 0.03968f
C16925 net68 _036_ 0.168017f
C16926 _000_ net4 0.036895f
C16927 net35 _140_ 0.12583f
C16928 output34/a_224_472# output18/a_224_472# 0.002121f
C16929 FILLER_0_4_107/a_1380_472# _152_ 0.001297f
C16930 _432_/a_2665_112# FILLER_0_18_177/a_2276_472# 0.021761f
C16931 _101_ _099_ 0.198807f
C16932 _412_/a_2665_112# cal_itt\[1\] 0.015571f
C16933 net52 FILLER_0_5_72/a_1380_472# 0.001523f
C16934 net29 _094_ 0.313846f
C16935 net56 FILLER_0_17_142/a_124_375# 0.004803f
C16936 _183_ _041_ 0.001931f
C16937 net79 result[3] 0.138076f
C16938 _053_ net67 0.672744f
C16939 _255_/a_224_552# _057_ 0.024333f
C16940 net48 net76 0.069349f
C16941 mask\[0\] _429_/a_796_472# 0.007281f
C16942 net16 _042_ 0.012486f
C16943 net55 FILLER_0_18_53/a_572_375# 0.015895f
C16944 FILLER_0_7_233/a_124_375# vdd 0.03915f
C16945 ctln[1] net65 0.073241f
C16946 net38 _452_/a_36_151# 0.010095f
C16947 _175_ _040_ 0.00133f
C16948 FILLER_0_2_111/a_1380_472# vss 0.001679f
C16949 FILLER_0_12_136/a_572_375# net23 0.00281f
C16950 _105_ _048_ 0.02699f
C16951 _134_ vss 0.088213f
C16952 net72 FILLER_0_21_28/a_572_375# 0.005742f
C16953 _133_ _163_ 0.034905f
C16954 _428_/a_2560_156# _131_ 0.002853f
C16955 _043_ FILLER_0_12_196/a_36_472# 0.001526f
C16956 FILLER_0_20_177/a_1468_375# _098_ 0.012889f
C16957 net35 FILLER_0_21_150/a_36_472# 0.004456f
C16958 _132_ FILLER_0_19_134/a_124_375# 0.00141f
C16959 _103_ _418_/a_1308_423# 0.004778f
C16960 _379_/a_36_472# _035_ 0.002226f
C16961 FILLER_0_4_123/a_124_375# trim_mask\[4\] 0.004312f
C16962 _174_ _043_ 0.964645f
C16963 _136_ FILLER_0_15_180/a_484_472# 0.002128f
C16964 net81 net28 0.034606f
C16965 _412_/a_2665_112# vss 0.011887f
C16966 _207_/a_67_603# mask\[6\] 0.072291f
C16967 _376_/a_36_160# _163_ 0.006811f
C16968 net63 FILLER_0_20_177/a_1380_472# 0.011079f
C16969 FILLER_0_21_133/a_124_375# _433_/a_36_151# 0.059049f
C16970 net59 net11 0.016998f
C16971 net34 _435_/a_2560_156# 0.002967f
C16972 net50 FILLER_0_8_24/a_124_375# 0.001597f
C16973 FILLER_0_7_72/a_572_375# net50 0.012932f
C16974 _093_ FILLER_0_17_72/a_3260_375# 0.011936f
C16975 FILLER_0_18_2/a_2724_472# _452_/a_1040_527# 0.001138f
C16976 _325_/a_224_472# _086_ 0.003155f
C16977 _046_ net30 0.006105f
C16978 FILLER_0_23_60/a_36_472# vdd 0.090554f
C16979 FILLER_0_23_60/a_124_375# vss 0.004081f
C16980 FILLER_0_6_177/a_124_375# vss 0.002362f
C16981 FILLER_0_6_177/a_572_375# vdd 0.02743f
C16982 output20/a_224_472# _109_ 0.003452f
C16983 _428_/a_36_151# FILLER_0_13_100/a_36_472# 0.004032f
C16984 ctln[1] net59 0.053978f
C16985 net80 mask\[7\] 0.020051f
C16986 _052_ FILLER_0_21_60/a_124_375# 0.002308f
C16987 net81 _429_/a_1204_472# 0.005046f
C16988 net64 FILLER_0_12_236/a_572_375# 0.005704f
C16989 mask\[4\] FILLER_0_19_195/a_36_472# 0.004669f
C16990 net63 FILLER_0_18_177/a_1020_375# 0.007516f
C16991 net76 net19 0.02061f
C16992 _233_/a_36_160# net17 0.003831f
C16993 _441_/a_1204_472# _168_ 0.009437f
C16994 trim_mask\[2\] _168_ 0.00704f
C16995 net81 FILLER_0_10_247/a_124_375# 0.044906f
C16996 net16 FILLER_0_14_50/a_36_472# 0.001377f
C16997 net15 _394_/a_728_93# 0.085551f
C16998 result[5] _418_/a_796_472# 0.001983f
C16999 _343_/a_257_69# _141_ 0.001515f
C17000 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_124_375# 0.026339f
C17001 _076_ net59 0.005449f
C17002 net27 FILLER_0_9_270/a_572_375# 0.043797f
C17003 FILLER_0_16_107/a_36_472# _131_ 0.008817f
C17004 net27 _015_ 0.103416f
C17005 FILLER_0_19_47/a_124_375# _013_ 0.023766f
C17006 cal_count\[3\] FILLER_0_11_78/a_484_472# 0.011737f
C17007 _079_ FILLER_0_5_206/a_124_375# 0.009128f
C17008 _098_ FILLER_0_19_171/a_484_472# 0.010731f
C17009 FILLER_0_16_255/a_124_375# _006_ 0.02007f
C17010 net57 _131_ 0.030577f
C17011 FILLER_0_16_89/a_484_472# net36 0.003595f
C17012 _428_/a_448_472# net70 0.007116f
C17013 FILLER_0_5_109/a_572_375# net47 0.011047f
C17014 _085_ _310_/a_49_472# 0.001093f
C17015 net60 _420_/a_2665_112# 0.038894f
C17016 mask\[4\] _346_/a_49_472# 0.079347f
C17017 net16 cal_count\[3\] 0.082821f
C17018 _074_ _122_ 0.300373f
C17019 FILLER_0_9_60/a_484_472# FILLER_0_9_72/a_36_472# 0.002296f
C17020 _126_ _129_ 0.039006f
C17021 net15 FILLER_0_13_80/a_36_472# 0.001122f
C17022 _188_ FILLER_0_12_50/a_36_472# 0.006464f
C17023 _064_ _033_ 0.001986f
C17024 net75 vdd 1.265616f
C17025 ctln[0] net40 0.001334f
C17026 net54 FILLER_0_20_98/a_36_472# 0.059367f
C17027 net32 net61 0.056005f
C17028 net82 FILLER_0_3_172/a_572_375# 0.010972f
C17029 FILLER_0_7_72/a_1916_375# FILLER_0_6_90/a_36_472# 0.001684f
C17030 cal_itt\[3\] _116_ 0.001364f
C17031 _214_/a_36_160# _437_/a_36_151# 0.001542f
C17032 _430_/a_2248_156# FILLER_0_15_212/a_932_472# 0.035805f
C17033 FILLER_0_0_266/a_36_472# rstn 0.006108f
C17034 net72 vdd 1.425686f
C17035 _108_ mask\[6\] 0.032481f
C17036 _452_/a_1040_527# vdd 0.004153f
C17037 output20/a_224_472# _422_/a_448_472# 0.009204f
C17038 _058_ FILLER_0_10_94/a_484_472# 0.002096f
C17039 _406_/a_36_159# cal_count\[2\] 0.028829f
C17040 net55 net17 0.056153f
C17041 trim_mask\[4\] _163_ 0.003686f
C17042 FILLER_0_17_72/a_3172_472# vss 0.001338f
C17043 FILLER_0_7_146/a_36_472# _059_ 0.073041f
C17044 _028_ FILLER_0_7_104/a_1020_375# 0.004954f
C17045 _425_/a_448_472# FILLER_0_8_247/a_932_472# 0.012285f
C17046 _308_/a_124_24# trim_mask\[0\] 0.018998f
C17047 FILLER_0_9_223/a_124_375# _128_ 0.004252f
C17048 _077_ FILLER_0_8_156/a_124_375# 0.00407f
C17049 _430_/a_36_151# net36 0.003701f
C17050 net20 FILLER_0_1_204/a_36_472# 0.001278f
C17051 net38 net39 0.066083f
C17052 FILLER_0_10_37/a_124_375# FILLER_0_10_28/a_124_375# 0.003228f
C17053 net15 FILLER_0_18_76/a_36_472# 0.001341f
C17054 _057_ _128_ 0.036548f
C17055 FILLER_0_9_223/a_484_472# net20 0.002601f
C17056 net60 _421_/a_1288_156# 0.001147f
C17057 FILLER_0_18_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001597f
C17058 FILLER_0_4_49/a_572_375# _440_/a_36_151# 0.073306f
C17059 result[0] calibrate 0.00287f
C17060 net15 _423_/a_2248_156# 0.048449f
C17061 net38 _039_ 0.059899f
C17062 _390_/a_36_68# _172_ 0.033476f
C17063 net16 net40 0.039189f
C17064 _074_ _061_ 0.007152f
C17065 _350_/a_49_472# net23 0.002397f
C17066 net57 _428_/a_2665_112# 0.027291f
C17067 result[8] ctlp[3] 0.278543f
C17068 FILLER_0_21_133/a_36_472# net54 0.02286f
C17069 net61 _422_/a_2248_156# 0.027973f
C17070 net20 _080_ 0.093195f
C17071 _106_ vss 0.180823f
C17072 _132_ _428_/a_448_472# 0.034825f
C17073 FILLER_0_17_72/a_1916_375# net36 0.015395f
C17074 FILLER_0_6_37/a_36_472# _160_ 0.008686f
C17075 FILLER_0_16_73/a_124_375# vdd 0.008987f
C17076 FILLER_0_9_28/a_124_375# net47 0.006757f
C17077 FILLER_0_22_128/a_572_375# vdd 0.001473f
C17078 FILLER_0_6_239/a_36_472# net37 0.004187f
C17079 net25 FILLER_0_22_86/a_572_375# 0.002444f
C17080 net18 net30 0.09055f
C17081 _086_ _116_ 1.316798f
C17082 _048_ _047_ 0.007849f
C17083 _024_ vdd 0.091532f
C17084 _422_/a_36_151# _299_/a_36_472# 0.004432f
C17085 FILLER_0_21_142/a_124_375# net54 0.027551f
C17086 _424_/a_36_151# vdd 0.125156f
C17087 _432_/a_2665_112# _093_ 0.02266f
C17088 ctln[5] FILLER_0_0_198/a_36_472# 0.012298f
C17089 _131_ FILLER_0_10_107/a_572_375# 0.007252f
C17090 _052_ _424_/a_2248_156# 0.005116f
C17091 output15/a_224_472# net49 0.005626f
C17092 net15 net66 0.006618f
C17093 net34 FILLER_0_22_128/a_3172_472# 0.003953f
C17094 _287_/a_36_472# _102_ 0.028733f
C17095 _441_/a_796_472# vss 0.001231f
C17096 FILLER_0_5_88/a_124_375# net47 0.005083f
C17097 _098_ _434_/a_2665_112# 0.013854f
C17098 _099_ _282_/a_36_160# 0.005808f
C17099 FILLER_0_7_72/a_2364_375# net50 0.017301f
C17100 net55 _452_/a_36_151# 0.042427f
C17101 FILLER_0_13_206/a_36_472# vdd 0.011681f
C17102 FILLER_0_13_206/a_124_375# vss 0.051723f
C17103 _009_ _108_ 1.645945f
C17104 _193_/a_36_160# FILLER_0_13_290/a_124_375# 0.005732f
C17105 _447_/a_448_472# vdd 0.014537f
C17106 _447_/a_36_151# vss 0.001541f
C17107 _242_/a_36_160# _170_ 0.001933f
C17108 _117_ _310_/a_1133_69# 0.002654f
C17109 net58 _416_/a_36_151# 0.001558f
C17110 trimb[0] vss 0.097724f
C17111 _084_ _316_/a_124_24# 0.001501f
C17112 result[7] _093_ 0.001096f
C17113 net62 FILLER_0_15_228/a_124_375# 0.001408f
C17114 FILLER_0_11_101/a_484_472# _120_ 0.011393f
C17115 net63 _434_/a_3041_156# 0.001449f
C17116 _440_/a_2665_112# vss 0.008703f
C17117 result[2] output30/a_224_472# 0.045862f
C17118 _439_/a_1308_423# vss 0.009355f
C17119 net81 FILLER_0_15_205/a_36_472# 0.081574f
C17120 vss FILLER_0_13_290/a_36_472# 0.009561f
C17121 net45 net40 0.029947f
C17122 en cal_itt\[1\] 0.028447f
C17123 fanout56/a_36_113# vss 0.03072f
C17124 _088_ net82 0.160444f
C17125 net16 _379_/a_36_472# 0.01109f
C17126 trim_val\[0\] trim_mask\[1\] 0.003033f
C17127 net53 net36 3.423337f
C17128 _443_/a_2665_112# _037_ 0.004052f
C17129 calibrate _062_ 2.032477f
C17130 _077_ net51 0.76967f
C17131 output37/a_224_472# calibrate 0.013149f
C17132 net76 FILLER_0_3_172/a_484_472# 0.002542f
C17133 _131_ FILLER_0_17_104/a_1380_472# 0.004125f
C17134 _426_/a_36_151# FILLER_0_8_247/a_1468_375# 0.059049f
C17135 net57 _126_ 0.021705f
C17136 _431_/a_2665_112# net36 0.001523f
C17137 net56 _433_/a_2665_112# 0.003434f
C17138 net56 FILLER_0_18_139/a_1020_375# 0.018398f
C17139 FILLER_0_6_47/a_2724_472# vss 0.020876f
C17140 FILLER_0_6_47/a_3172_472# vdd 0.002089f
C17141 _175_ FILLER_0_15_72/a_484_472# 0.020589f
C17142 trim[1] vss 0.085436f
C17143 sample en 0.001572f
C17144 net67 _221_/a_36_160# 0.008581f
C17145 mask\[9\] net14 0.090939f
C17146 FILLER_0_12_124/a_36_472# FILLER_0_11_124/a_36_472# 0.05841f
C17147 net17 _381_/a_36_472# 0.002796f
C17148 net58 net65 1.468105f
C17149 net15 _067_ 0.042278f
C17150 vdd cal_count\[0\] 0.491891f
C17151 net35 _435_/a_36_151# 0.038368f
C17152 en vss 0.466499f
C17153 _425_/a_448_472# _014_ 0.013561f
C17154 FILLER_0_10_78/a_932_472# vss 0.002987f
C17155 _069_ _043_ 0.04044f
C17156 mask\[5\] FILLER_0_19_171/a_572_375# 0.007169f
C17157 _118_ _311_/a_3740_473# 0.001244f
C17158 _414_/a_2248_156# vdd 0.00901f
C17159 net72 _424_/a_36_151# 0.09381f
C17160 _418_/a_1000_472# _007_ 0.001051f
C17161 _431_/a_1308_423# net73 0.039024f
C17162 output39/a_224_472# _063_ 0.001019f
C17163 net39 _233_/a_36_160# 0.017979f
C17164 _311_/a_254_473# vdd 0.001207f
C17165 FILLER_0_24_130/a_36_472# _050_ 0.008605f
C17166 net63 _430_/a_448_472# 0.026599f
C17167 output42/a_224_472# FILLER_0_8_2/a_124_375# 0.030009f
C17168 _093_ _008_ 0.252609f
C17169 net53 FILLER_0_14_123/a_124_375# 0.003138f
C17170 input5/a_36_113# clk 0.01086f
C17171 FILLER_0_22_86/a_1380_472# net14 0.039176f
C17172 _091_ FILLER_0_19_171/a_932_472# 0.002509f
C17173 trimb[3] net38 0.002836f
C17174 _072_ _176_ 0.298077f
C17175 _301_/a_36_472# net25 0.003165f
C17176 _448_/a_2665_112# net59 0.005948f
C17177 _141_ net80 0.077957f
C17178 net20 _323_/a_36_113# 0.002161f
C17179 _176_ FILLER_0_15_59/a_572_375# 0.007169f
C17180 _072_ _306_/a_36_68# 0.042843f
C17181 _053_ _059_ 0.042128f
C17182 _086_ _117_ 0.010287f
C17183 _031_ _160_ 0.004547f
C17184 _258_/a_36_160# net37 0.006865f
C17185 _077_ FILLER_0_9_72/a_1020_375# 0.008103f
C17186 _374_/a_36_68# vdd 0.075685f
C17187 _427_/a_1000_472# vss 0.012657f
C17188 _321_/a_170_472# net74 0.020269f
C17189 _415_/a_1204_472# result[1] 0.004051f
C17190 net58 net59 0.066534f
C17191 output44/a_224_472# FILLER_0_19_28/a_124_375# 0.005166f
C17192 net28 mask\[1\] 0.572459f
C17193 FILLER_0_8_24/a_124_375# _054_ 0.008177f
C17194 _186_ _067_ 0.001907f
C17195 _273_/a_36_68# _060_ 0.010339f
C17196 output35/a_224_472# FILLER_0_22_177/a_1380_472# 0.002486f
C17197 _072_ _251_/a_1130_472# 0.004007f
C17198 _281_/a_672_472# vdd 0.001069f
C17199 _448_/a_36_151# FILLER_0_2_177/a_36_472# 0.04556f
C17200 _136_ FILLER_0_14_99/a_36_472# 0.01535f
C17201 _179_ _180_ 0.018662f
C17202 _331_/a_448_472# vdd 0.001343f
C17203 _038_ _120_ 0.00117f
C17204 _431_/a_36_151# FILLER_0_18_139/a_36_472# 0.002529f
C17205 net44 _450_/a_836_156# 0.006278f
C17206 FILLER_0_10_78/a_124_375# cal_count\[3\] 0.012197f
C17207 FILLER_0_7_72/a_1828_472# net52 0.00159f
C17208 FILLER_0_10_247/a_124_375# net64 0.001597f
C17209 _449_/a_1000_472# _067_ 0.021759f
C17210 _402_/a_1948_68# _182_ 0.016049f
C17211 FILLER_0_13_212/a_572_375# vdd 0.001551f
C17212 FILLER_0_13_212/a_124_375# vss 0.007116f
C17213 _033_ _444_/a_2248_156# 0.011578f
C17214 _081_ _265_/a_224_472# 0.008598f
C17215 _436_/a_448_472# vdd 0.038494f
C17216 _068_ _311_/a_3740_473# 0.001409f
C17217 net76 FILLER_0_6_177/a_484_472# 0.016333f
C17218 _125_ _062_ 0.061735f
C17219 _235_/a_255_603# trim_val\[2\] 0.002471f
C17220 output47/a_224_472# FILLER_0_15_2/a_484_472# 0.038484f
C17221 FILLER_0_11_142/a_572_375# cal_count\[3\] 0.014082f
C17222 _370_/a_1152_472# _152_ 0.001423f
C17223 _411_/a_2665_112# _073_ 0.009313f
C17224 _076_ _120_ 0.736844f
C17225 trim_mask\[2\] _447_/a_36_151# 0.022881f
C17226 FILLER_0_17_226/a_36_472# _008_ 0.001842f
C17227 _091_ mask\[0\] 0.04171f
C17228 vdd _433_/a_36_151# 0.086874f
C17229 _238_/a_67_603# _441_/a_2665_112# 0.015187f
C17230 cal_count\[3\] _373_/a_1254_68# 0.001391f
C17231 net60 _418_/a_796_472# 0.008602f
C17232 FILLER_0_18_2/a_2364_375# net40 0.002024f
C17233 net34 _210_/a_255_603# 0.002153f
C17234 _445_/a_2665_112# net47 0.041188f
C17235 net60 _419_/a_2560_156# 0.006989f
C17236 _337_/a_49_472# vdd 0.028131f
C17237 net38 net42 0.012245f
C17238 _132_ FILLER_0_17_104/a_124_375# 0.001918f
C17239 _407_/a_36_472# vdd 0.095308f
C17240 ctln[0] trim[3] 0.216084f
C17241 net35 net14 0.040959f
C17242 net57 _137_ 0.006142f
C17243 _440_/a_36_151# _029_ 0.00874f
C17244 mask\[7\] FILLER_0_22_128/a_124_375# 0.01319f
C17245 FILLER_0_20_193/a_36_472# net21 0.001099f
C17246 _077_ _115_ 0.131611f
C17247 FILLER_0_4_152/a_36_472# vdd 0.087397f
C17248 FILLER_0_7_59/a_36_472# vss 0.004006f
C17249 FILLER_0_7_59/a_484_472# vdd 0.00824f
C17250 net54 FILLER_0_22_86/a_1468_375# 0.001597f
C17251 _053_ FILLER_0_5_212/a_36_472# 0.007052f
C17252 net35 FILLER_0_22_128/a_3260_375# 0.012732f
C17253 mask\[9\] _098_ 0.256513f
C17254 FILLER_0_1_204/a_36_472# vss 0.002247f
C17255 net36 _451_/a_36_151# 0.02414f
C17256 _053_ trim_val\[1\] 0.00385f
C17257 FILLER_0_20_98/a_124_375# _437_/a_36_151# 0.059049f
C17258 FILLER_0_8_263/a_124_375# net19 0.039576f
C17259 _437_/a_2665_112# FILLER_0_22_107/a_572_375# 0.001597f
C17260 net68 FILLER_0_6_47/a_1020_375# 0.029857f
C17261 FILLER_0_9_223/a_484_472# vss 0.006102f
C17262 _092_ FILLER_0_17_218/a_36_472# 0.033277f
C17263 net75 _411_/a_1000_472# 0.03227f
C17264 _104_ FILLER_0_23_274/a_36_472# 0.001642f
C17265 _136_ FILLER_0_16_154/a_1020_375# 0.004387f
C17266 trim_mask\[1\] FILLER_0_6_47/a_1916_375# 0.007169f
C17267 FILLER_0_3_142/a_124_375# vdd 0.00167f
C17268 FILLER_0_7_72/a_2812_375# _077_ 0.002969f
C17269 FILLER_0_13_206/a_124_375# net4 0.031251f
C17270 _285_/a_36_472# net36 0.003032f
C17271 _086_ FILLER_0_7_104/a_1020_375# 0.00757f
C17272 _114_ FILLER_0_12_136/a_484_472# 0.003953f
C17273 vdd FILLER_0_19_134/a_124_375# 0.027957f
C17274 net38 clkc 0.088241f
C17275 FILLER_0_0_96/a_124_375# net14 0.077876f
C17276 _080_ vss 0.012982f
C17277 FILLER_0_7_195/a_36_472# net21 0.005469f
C17278 _070_ FILLER_0_9_105/a_484_472# 0.020248f
C17279 net58 result[1] 0.004614f
C17280 _033_ _166_ 0.004448f
C17281 _444_/a_1308_423# vdd 0.005677f
C17282 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1468_375# 0.086635f
C17283 trim_val\[0\] _164_ 0.133785f
C17284 _150_ _438_/a_1000_472# 0.003452f
C17285 _066_ _163_ 0.006401f
C17286 _444_/a_1204_472# net17 0.021952f
C17287 ctlp[1] _421_/a_36_151# 0.010453f
C17288 net54 _437_/a_2665_112# 0.061157f
C17289 _427_/a_1308_423# net23 0.004863f
C17290 fanout77/a_36_113# _419_/a_36_151# 0.002361f
C17291 FILLER_0_4_99/a_36_472# vdd 0.094733f
C17292 FILLER_0_4_99/a_124_375# vss 0.017518f
C17293 net1 fanout59/a_36_160# 0.002325f
C17294 net25 FILLER_0_23_88/a_36_472# 0.192699f
C17295 _446_/a_36_151# net17 0.006518f
C17296 FILLER_0_7_146/a_124_375# vdd 0.034288f
C17297 _065_ _447_/a_2248_156# 0.038629f
C17298 _316_/a_124_24# calibrate 0.016936f
C17299 _189_/a_67_603# net64 0.064691f
C17300 _073_ FILLER_0_3_221/a_1380_472# 0.045839f
C17301 FILLER_0_7_162/a_124_375# _062_ 0.010242f
C17302 result[5] _103_ 0.425479f
C17303 mask\[4\] FILLER_0_18_209/a_124_375# 0.020811f
C17304 net22 FILLER_0_18_209/a_124_375# 0.012909f
C17305 _322_/a_124_24# _126_ 0.019609f
C17306 output40/a_224_472# net40 0.0374f
C17307 FILLER_0_6_239/a_36_472# _122_ 0.01785f
C17308 net23 FILLER_0_8_156/a_36_472# 0.004939f
C17309 ctlp[4] ctlp[5] 0.001257f
C17310 FILLER_0_2_93/a_572_375# _030_ 0.001718f
C17311 FILLER_0_8_2/a_36_472# net40 0.002477f
C17312 _417_/a_36_151# net30 0.010021f
C17313 FILLER_0_16_89/a_124_375# _136_ 0.011795f
C17314 net27 output27/a_224_472# 0.046353f
C17315 net65 FILLER_0_3_172/a_2276_472# 0.001777f
C17316 _077_ FILLER_0_6_231/a_124_375# 0.009235f
C17317 _116_ _161_ 0.008003f
C17318 FILLER_0_18_2/a_932_472# net44 0.012286f
C17319 en net4 0.125535f
C17320 FILLER_0_11_78/a_484_472# _120_ 0.016839f
C17321 FILLER_0_9_72/a_1380_472# vdd 0.007659f
C17322 FILLER_0_9_72/a_932_472# vss 0.007033f
C17323 net34 output33/a_224_472# 0.077682f
C17324 _074_ net8 0.001023f
C17325 mask\[1\] FILLER_0_15_205/a_36_472# 0.006921f
C17326 fanout57/a_36_113# net65 0.035361f
C17327 _163_ net37 0.079552f
C17328 _076_ _227_/a_36_160# 0.004997f
C17329 fanout70/a_36_113# _131_ 0.003364f
C17330 _404_/a_36_472# vdd 0.034854f
C17331 _346_/a_49_472# _140_ 0.003436f
C17332 net16 _120_ 0.009918f
C17333 net48 _251_/a_468_472# 0.002731f
C17334 _326_/a_36_160# FILLER_0_9_105/a_484_472# 0.002647f
C17335 FILLER_0_2_111/a_1468_375# _160_ 0.001026f
C17336 _056_ _226_/a_1044_68# 0.002852f
C17337 _144_ vss 0.411237f
C17338 _094_ _418_/a_448_472# 0.042782f
C17339 net81 _412_/a_1204_472# 0.003435f
C17340 _105_ net61 0.020753f
C17341 FILLER_0_9_28/a_2724_472# trim_val\[0\] 0.001183f
C17342 net63 FILLER_0_15_228/a_36_472# 0.001669f
C17343 output8/a_224_472# FILLER_0_3_221/a_932_472# 0.001699f
C17344 net50 _033_ 0.003088f
C17345 _390_/a_244_472# _038_ 0.001278f
C17346 _390_/a_36_68# _136_ 0.032598f
C17347 output46/a_224_472# vdd 0.043652f
C17348 net44 FILLER_0_20_2/a_36_472# 0.037627f
C17349 _254_/a_448_472# net22 0.009088f
C17350 net58 _415_/a_2560_156# 0.002325f
C17351 net57 FILLER_0_13_142/a_932_472# 0.01158f
C17352 net57 net56 0.054294f
C17353 fanout52/a_36_160# vdd 0.026513f
C17354 _000_ ctln[3] 0.008418f
C17355 _406_/a_36_159# _402_/a_56_567# 0.001025f
C17356 FILLER_0_20_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001543f
C17357 vdd _416_/a_2248_156# 0.004325f
C17358 net24 vdd 0.223761f
C17359 _367_/a_36_68# _154_ 0.028801f
C17360 _431_/a_2665_112# FILLER_0_18_139/a_1380_472# 0.001008f
C17361 ctlp[6] FILLER_0_24_130/a_124_375# 0.021926f
C17362 _036_ fanout66/a_36_113# 0.014556f
C17363 _408_/a_1336_472# _095_ 0.011305f
C17364 mask\[2\] FILLER_0_16_154/a_484_472# 0.028444f
C17365 _122_ FILLER_0_8_156/a_124_375# 0.032617f
C17366 FILLER_0_13_142/a_36_472# _043_ 0.011974f
C17367 fanout57/a_36_113# net59 0.00178f
C17368 _053_ _385_/a_244_472# 0.00134f
C17369 FILLER_0_14_91/a_484_472# _176_ 0.003624f
C17370 net35 _098_ 0.017288f
C17371 _176_ state\[1\] 0.001641f
C17372 output28/a_224_472# fanout79/a_36_160# 0.022393f
C17373 _390_/a_36_68# _070_ 0.047478f
C17374 _142_ mask\[2\] 0.093231f
C17375 net31 _103_ 0.227588f
C17376 _306_/a_36_68# state\[1\] 0.028553f
C17377 _099_ vdd 0.326559f
C17378 _392_/a_36_68# _039_ 0.001522f
C17379 mask\[7\] _436_/a_36_151# 0.030028f
C17380 _430_/a_36_151# FILLER_0_18_209/a_484_472# 0.001043f
C17381 net58 output9/a_224_472# 0.050634f
C17382 _412_/a_2248_156# net18 0.05155f
C17383 FILLER_0_5_109/a_572_375# vdd 0.024724f
C17384 _328_/a_36_113# _135_ 0.005635f
C17385 FILLER_0_21_28/a_3172_472# vss 0.001574f
C17386 FILLER_0_6_90/a_36_472# vss 0.001409f
C17387 FILLER_0_6_90/a_484_472# vdd 0.003146f
C17388 _148_ _436_/a_36_151# 0.032004f
C17389 _360_/a_36_160# _152_ 0.040508f
C17390 _040_ FILLER_0_16_115/a_36_472# 0.001876f
C17391 net35 _436_/a_2665_112# 0.012468f
C17392 _428_/a_36_151# vss 0.00285f
C17393 _428_/a_448_472# vdd 0.034564f
C17394 net15 FILLER_0_5_54/a_1380_472# 0.047774f
C17395 net72 _404_/a_36_472# 0.019911f
C17396 net52 FILLER_0_2_111/a_932_472# 0.061249f
C17397 cal_itt\[2\] FILLER_0_3_221/a_1380_472# 0.015024f
C17398 _372_/a_358_69# _070_ 0.001293f
C17399 _077_ _073_ 0.009611f
C17400 net74 FILLER_0_5_136/a_36_472# 0.003704f
C17401 _258_/a_36_160# _122_ 0.00102f
C17402 _114_ vss 0.365613f
C17403 _043_ _090_ 0.001578f
C17404 _161_ _117_ 0.25528f
C17405 _163_ FILLER_0_5_148/a_484_472# 0.002734f
C17406 net37 FILLER_0_6_231/a_124_375# 0.001989f
C17407 fanout50/a_36_160# vss 0.009871f
C17408 FILLER_0_17_72/a_932_472# _131_ 0.002672f
C17409 net74 _135_ 0.002261f
C17410 _414_/a_796_472# vdd 0.001497f
C17411 vss FILLER_0_14_235/a_484_472# 0.003246f
C17412 net62 FILLER_0_14_235/a_572_375# 0.017549f
C17413 _443_/a_448_472# vdd 0.007773f
C17414 _443_/a_36_151# vss 0.019802f
C17415 net81 FILLER_0_15_212/a_1380_472# 0.003953f
C17416 _292_/a_36_160# net22 0.001864f
C17417 _165_ FILLER_0_6_37/a_124_375# 0.002884f
C17418 _341_/a_49_472# FILLER_0_17_161/a_36_472# 0.079018f
C17419 net38 FILLER_0_15_2/a_484_472# 0.003391f
C17420 FILLER_0_13_206/a_124_375# net79 0.009649f
C17421 _411_/a_1204_472# net8 0.001768f
C17422 _043_ net22 0.041447f
C17423 net49 FILLER_0_3_54/a_36_472# 0.00186f
C17424 FILLER_0_20_177/a_1468_375# _434_/a_2248_156# 0.001221f
C17425 FILLER_0_5_72/a_36_472# _440_/a_36_151# 0.001723f
C17426 _072_ FILLER_0_12_220/a_484_472# 0.028355f
C17427 _088_ FILLER_0_3_212/a_36_472# 0.005583f
C17428 _413_/a_2665_112# vdd 0.02286f
C17429 _069_ _062_ 0.029863f
C17430 net79 FILLER_0_13_290/a_36_472# 0.038324f
C17431 net68 FILLER_0_3_54/a_36_472# 0.049455f
C17432 _037_ net12 0.007817f
C17433 FILLER_0_9_223/a_484_472# net4 0.047334f
C17434 _414_/a_2665_112# _072_ 0.025361f
C17435 cal_count\[3\] net14 0.028995f
C17436 _155_ _151_ 0.10611f
C17437 output35/a_224_472# _435_/a_36_151# 0.001362f
C17438 _053_ FILLER_0_6_177/a_124_375# 0.009352f
C17439 FILLER_0_9_28/a_124_375# vdd -0.004893f
C17440 _093_ FILLER_0_19_155/a_484_472# 0.001236f
C17441 net16 FILLER_0_18_37/a_124_375# 0.017482f
C17442 _321_/a_1194_69# vss 0.0011f
C17443 FILLER_0_4_197/a_36_472# net21 0.011079f
C17444 _430_/a_2248_156# mask\[1\] 0.001498f
C17445 FILLER_0_2_177/a_572_375# vdd 0.022268f
C17446 FILLER_0_2_177/a_124_375# vss 0.00252f
C17447 net4 _080_ 0.076128f
C17448 _058_ FILLER_0_8_156/a_484_472# 0.013955f
C17449 net16 _446_/a_2248_156# 0.010032f
C17450 FILLER_0_17_218/a_572_375# vss 0.078608f
C17451 FILLER_0_17_218/a_36_472# vdd 0.084913f
C17452 _379_/a_36_472# _063_ 0.071695f
C17453 _139_ FILLER_0_15_180/a_572_375# 0.022254f
C17454 FILLER_0_5_88/a_124_375# vdd 0.020896f
C17455 _116_ _071_ 0.017991f
C17456 net71 FILLER_0_22_107/a_572_375# 0.006403f
C17457 _020_ FILLER_0_18_107/a_2364_375# 0.003755f
C17458 _412_/a_1000_472# net81 0.012828f
C17459 _435_/a_1288_156# vdd 0.001119f
C17460 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_572_375# 0.086635f
C17461 _130_ _427_/a_36_151# 0.001056f
C17462 FILLER_0_8_263/a_36_472# vss 0.001089f
C17463 FILLER_0_20_31/a_36_472# vss 0.004923f
C17464 net67 FILLER_0_9_60/a_484_472# 0.001345f
C17465 FILLER_0_13_65/a_36_472# net15 0.036527f
C17466 _360_/a_36_160# _070_ 0.012463f
C17467 net54 FILLER_0_21_150/a_124_375# 0.007123f
C17468 FILLER_0_17_200/a_484_472# _093_ 0.007492f
C17469 net20 _421_/a_1308_423# 0.012036f
C17470 FILLER_0_21_286/a_124_375# vss 0.005049f
C17471 FILLER_0_21_286/a_572_375# vdd 0.03062f
C17472 _181_ _180_ 0.216908f
C17473 net76 FILLER_0_5_198/a_572_375# 0.006974f
C17474 clk rstn 0.541051f
C17475 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_124_375# 0.005439f
C17476 _017_ FILLER_0_13_100/a_124_375# 0.001274f
C17477 FILLER_0_21_28/a_1828_472# _423_/a_36_151# 0.059367f
C17478 fanout70/a_36_113# FILLER_0_15_116/a_572_375# 0.003553f
C17479 _073_ net37 0.013152f
C17480 _421_/a_448_472# net19 0.058446f
C17481 net57 _095_ 0.07431f
C17482 FILLER_0_8_138/a_36_472# _313_/a_67_603# 0.005759f
C17483 _081_ _059_ 0.04053f
C17484 net54 net71 0.536043f
C17485 result[7] FILLER_0_24_274/a_572_375# 0.006125f
C17486 _451_/a_2449_156# _040_ 0.004434f
C17487 output48/a_224_472# _081_ 0.007705f
C17488 cal_itt\[3\] _375_/a_36_68# 0.005168f
C17489 FILLER_0_15_212/a_124_375# vdd -0.004549f
C17490 _077_ _067_ 0.090648f
C17491 net62 net36 0.034265f
C17492 output21/a_224_472# _108_ 0.005356f
C17493 _008_ _094_ 0.234346f
C17494 _144_ mask\[7\] 0.111088f
C17495 _093_ net14 0.11038f
C17496 trim[0] net66 0.376153f
C17497 FILLER_0_4_123/a_36_472# _153_ 0.001419f
C17498 mask\[4\] FILLER_0_20_177/a_484_472# 0.001215f
C17499 net70 _017_ 0.015488f
C17500 _144_ _148_ 0.038002f
C17501 _128_ _120_ 0.053476f
C17502 _106_ fanout63/a_36_160# 0.00715f
C17503 FILLER_0_10_78/a_124_375# _120_ 0.006134f
C17504 _093_ FILLER_0_17_161/a_124_375# 0.002431f
C17505 _072_ _250_/a_36_68# 0.007337f
C17506 net44 vdd 0.897202f
C17507 FILLER_0_7_72/a_2276_472# _439_/a_2248_156# 0.013656f
C17508 _171_ vdd 0.038202f
C17509 net34 FILLER_0_22_177/a_1020_375# 0.006974f
C17510 net20 FILLER_0_8_239/a_124_375# 0.004302f
C17511 trim[2] output41/a_224_472# 0.005452f
C17512 output40/a_224_472# trim[3] 0.122003f
C17513 net80 _434_/a_448_472# 0.113898f
C17514 _415_/a_1204_472# net27 0.006198f
C17515 mask\[4\] FILLER_0_18_177/a_124_375# 0.016093f
C17516 net65 net82 0.630327f
C17517 net60 _103_ 0.066266f
C17518 FILLER_0_11_142/a_572_375# _120_ 0.009014f
C17519 FILLER_0_17_72/a_1380_472# _150_ 0.014154f
C17520 FILLER_0_15_116/a_36_472# _095_ 0.001098f
C17521 _245_/a_234_472# net6 0.001301f
C17522 net50 _441_/a_36_151# 0.060777f
C17523 net52 _441_/a_1308_423# 0.059264f
C17524 FILLER_0_13_212/a_124_375# net79 0.007396f
C17525 FILLER_0_16_89/a_124_375# _451_/a_448_472# 0.001597f
C17526 _086_ _375_/a_36_68# 0.038443f
C17527 _096_ _320_/a_36_472# 0.052438f
C17528 comp vss 0.148428f
C17529 _429_/a_2248_156# FILLER_0_13_228/a_36_472# 0.035805f
C17530 _119_ _059_ 0.039711f
C17531 net63 mask\[3\] 0.37365f
C17532 result[7] FILLER_0_23_274/a_36_472# 0.014434f
C17533 net73 FILLER_0_17_104/a_1468_375# 0.002342f
C17534 net52 _440_/a_2248_156# 0.028463f
C17535 _033_ _054_ 0.003394f
C17536 _187_ vss 0.080956f
C17537 net52 _439_/a_448_472# 0.042072f
C17538 FILLER_0_8_138/a_36_472# _058_ 0.005325f
C17539 _129_ net74 0.476969f
C17540 _122_ _163_ 0.156898f
C17541 output20/a_224_472# result[9] 0.001884f
C17542 FILLER_0_17_104/a_124_375# vdd 0.030663f
C17543 FILLER_0_18_2/a_1468_375# net17 0.004803f
C17544 _323_/a_36_113# net4 0.005657f
C17545 FILLER_0_4_177/a_36_472# _074_ 0.002603f
C17546 mask\[4\] FILLER_0_19_171/a_1380_472# 0.002581f
C17547 FILLER_0_5_54/a_572_375# FILLER_0_6_47/a_1380_472# 0.001597f
C17548 net55 net36 0.273956f
C17549 _425_/a_36_151# net37 0.003145f
C17550 _119_ _375_/a_36_68# 0.007338f
C17551 _085_ vss 0.132721f
C17552 _176_ vdd 0.874707f
C17553 _077_ FILLER_0_9_105/a_36_472# 0.003177f
C17554 _106_ FILLER_0_17_218/a_484_472# 0.012952f
C17555 FILLER_0_5_164/a_572_375# vdd 0.0042f
C17556 net55 FILLER_0_19_28/a_36_472# 0.001572f
C17557 _239_/a_36_160# vdd 0.042369f
C17558 _010_ _420_/a_448_472# 0.027802f
C17559 net34 net20 0.003775f
C17560 _115_ _122_ 0.004082f
C17561 net82 net59 0.102279f
C17562 _321_/a_358_69# net23 0.001718f
C17563 _306_/a_36_68# vdd 0.044152f
C17564 _132_ _017_ 0.155924f
C17565 FILLER_0_5_212/a_36_472# _081_ 0.01062f
C17566 _335_/a_49_472# vdd 0.085394f
C17567 net69 FILLER_0_2_111/a_1020_375# 0.018655f
C17568 _031_ FILLER_0_2_111/a_124_375# 0.05482f
C17569 net52 FILLER_0_6_47/a_2276_472# 0.003298f
C17570 FILLER_0_22_128/a_3172_472# vss 0.006339f
C17571 output13/a_224_472# net12 0.002723f
C17572 net32 _421_/a_2560_156# 0.049213f
C17573 result[4] net62 0.050684f
C17574 net38 FILLER_0_20_15/a_484_472# 0.003376f
C17575 _018_ vss 0.022336f
C17576 _020_ net70 0.014391f
C17577 fanout71/a_36_113# net54 0.001194f
C17578 net1 net37 0.00519f
C17579 _251_/a_906_472# vss 0.0016f
C17580 _442_/a_2665_112# vss 0.001727f
C17581 _442_/a_2560_156# vdd 0.006195f
C17582 FILLER_0_15_142/a_484_472# FILLER_0_15_150/a_36_472# 0.013277f
C17583 _053_ FILLER_0_6_47/a_2724_472# 0.001777f
C17584 _036_ vdd 0.364747f
C17585 _131_ _451_/a_3129_107# 0.001608f
C17586 _144_ _433_/a_448_472# 0.075144f
C17587 mask\[0\] _113_ 0.01678f
C17588 _071_ _225_/a_36_160# 0.002808f
C17589 _428_/a_2248_156# _427_/a_36_151# 0.035837f
C17590 _445_/a_2665_112# vdd 0.055628f
C17591 FILLER_0_14_91/a_572_375# _136_ 0.049763f
C17592 _428_/a_2560_156# net74 0.002759f
C17593 mask\[5\] _048_ 0.062788f
C17594 net29 _044_ 0.01495f
C17595 net36 net23 0.028202f
C17596 _421_/a_796_472# _010_ 0.037434f
C17597 mask\[5\] FILLER_0_18_177/a_484_472# 0.001063f
C17598 _072_ net48 0.037795f
C17599 FILLER_0_19_55/a_124_375# net55 0.005311f
C17600 _104_ _422_/a_2665_112# 0.040586f
C17601 _322_/a_848_380# _118_ 0.047787f
C17602 net16 FILLER_0_17_38/a_572_375# 0.018281f
C17603 state\[0\] _070_ 0.009608f
C17604 _428_/a_36_151# _332_/a_36_472# 0.004432f
C17605 FILLER_0_14_181/a_124_375# vdd 0.040138f
C17606 FILLER_0_13_65/a_124_375# vdd 0.011301f
C17607 net55 _423_/a_2560_156# 0.002265f
C17608 _253_/a_36_68# _084_ 0.029805f
C17609 _425_/a_1204_472# vdd 0.015969f
C17610 output27/a_224_472# result[0] 0.031252f
C17611 state\[0\] FILLER_0_12_220/a_1380_472# 0.003733f
C17612 ctlp[7] _025_ 0.007483f
C17613 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_124_375# 0.012001f
C17614 _072_ _162_ 0.090175f
C17615 _100_ FILLER_0_12_236/a_572_375# 0.015109f
C17616 _093_ _098_ 0.556613f
C17617 FILLER_0_17_226/a_124_375# _093_ 0.001604f
C17618 net72 _176_ 0.059793f
C17619 _017_ FILLER_0_14_107/a_572_375# 0.003679f
C17620 mask\[7\] _435_/a_2560_156# 0.011544f
C17621 net70 FILLER_0_14_107/a_1468_375# 0.007955f
C17622 net16 _043_ 0.049385f
C17623 net58 net27 0.190417f
C17624 _114_ _332_/a_36_472# 0.021351f
C17625 FILLER_0_15_212/a_1380_472# mask\[1\] 0.041503f
C17626 net76 fanout76/a_36_160# 0.004503f
C17627 _122_ FILLER_0_6_231/a_124_375# 0.013183f
C17628 _070_ FILLER_0_10_94/a_484_472# 0.003573f
C17629 _050_ _436_/a_1204_472# 0.006724f
C17630 sample fanout65/a_36_113# 0.050978f
C17631 _159_ _152_ 0.035925f
C17632 FILLER_0_3_204/a_124_375# FILLER_0_4_197/a_932_472# 0.001597f
C17633 FILLER_0_16_57/a_484_472# _131_ 0.008223f
C17634 _094_ _006_ 0.090405f
C17635 FILLER_0_17_133/a_124_375# vdd 0.010519f
C17636 _020_ _132_ 0.037636f
C17637 _420_/a_448_472# vdd 0.010071f
C17638 _420_/a_36_151# vss 0.043027f
C17639 net16 _185_ 0.086347f
C17640 fanout65/a_36_113# vss 0.053899f
C17641 _162_ net47 0.004104f
C17642 _432_/a_36_151# mask\[3\] 0.002148f
C17643 _320_/a_672_472# vdd 0.008437f
C17644 _098_ FILLER_0_15_180/a_572_375# 0.01526f
C17645 net20 _419_/a_448_472# 0.025583f
C17646 _013_ FILLER_0_18_37/a_572_375# 0.003828f
C17647 net57 net74 2.360287f
C17648 net19 _419_/a_36_151# 0.009613f
C17649 _414_/a_36_151# FILLER_0_7_195/a_36_472# 0.001723f
C17650 FILLER_0_20_15/a_1380_472# vss 0.003678f
C17651 mask\[9\] _438_/a_1308_423# 0.044336f
C17652 _093_ FILLER_0_18_139/a_572_375# 0.008393f
C17653 FILLER_0_18_209/a_484_472# _201_/a_67_603# 0.001605f
C17654 FILLER_0_16_73/a_572_375# FILLER_0_17_72/a_572_375# 0.026339f
C17655 _087_ _074_ 0.004231f
C17656 _434_/a_36_151# vdd 0.104871f
C17657 FILLER_0_3_172/a_1468_375# net22 0.012895f
C17658 output35/a_224_472# _098_ 0.003653f
C17659 FILLER_0_13_142/a_124_375# vdd 0.02675f
C17660 _132_ FILLER_0_11_109/a_124_375# 0.008627f
C17661 FILLER_0_17_72/a_1828_472# _438_/a_36_151# 0.001221f
C17662 FILLER_0_16_73/a_124_375# _176_ 0.006386f
C17663 FILLER_0_21_133/a_124_375# FILLER_0_21_125/a_572_375# 0.012001f
C17664 output34/a_224_472# mask\[3\] 0.002385f
C17665 FILLER_0_17_200/a_572_375# vss 0.017327f
C17666 _430_/a_36_151# net80 0.082603f
C17667 _183_ vdd 0.109252f
C17668 net75 _425_/a_1204_472# 0.015778f
C17669 _144_ _141_ 0.095441f
C17670 _082_ vdd 0.191411f
C17671 net20 mask\[2\] 0.050364f
C17672 net79 _416_/a_1204_472# 0.006493f
C17673 output37/a_224_472# output27/a_224_472# 0.012653f
C17674 _322_/a_848_380# _068_ 0.009682f
C17675 FILLER_0_13_65/a_124_375# net72 0.002341f
C17676 _186_ _402_/a_728_93# 0.002381f
C17677 FILLER_0_8_247/a_1468_375# vss 0.054783f
C17678 FILLER_0_8_247/a_36_472# vdd 0.112197f
C17679 FILLER_0_14_91/a_36_472# net53 0.005849f
C17680 net76 FILLER_0_2_177/a_484_472# 0.012872f
C17681 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_484_472# 0.013277f
C17682 _057_ _126_ 0.022413f
C17683 _431_/a_1308_423# net36 0.002865f
C17684 fanout77/a_36_113# vdd 0.032109f
C17685 _132_ FILLER_0_14_107/a_1468_375# 0.019517f
C17686 net7 net17 0.050676f
C17687 comp input3/a_36_113# 0.022213f
C17688 net23 FILLER_0_22_128/a_2276_472# 0.011079f
C17689 FILLER_0_4_197/a_1020_375# vdd 0.002455f
C17690 FILLER_0_4_123/a_124_375# _160_ 0.038272f
C17691 net38 net67 1.762405f
C17692 cal_count\[2\] _402_/a_1948_68# 0.010022f
C17693 net63 FILLER_0_17_218/a_124_375# 0.040329f
C17694 FILLER_0_14_107/a_1380_472# _043_ 0.001641f
C17695 output25/a_224_472# ctlp[8] 0.018544f
C17696 _062_ _090_ 0.010805f
C17697 _426_/a_36_151# vss 0.003014f
C17698 _426_/a_448_472# vdd 0.042167f
C17699 en_co_clk _067_ 0.272082f
C17700 net63 _435_/a_2665_112# 0.039512f
C17701 cal_count\[3\] _405_/a_67_603# 0.011131f
C17702 _446_/a_796_472# net40 0.001504f
C17703 FILLER_0_1_98/a_36_472# _442_/a_2665_112# 0.002597f
C17704 _131_ cal_count\[3\] 0.035391f
C17705 trim_val\[2\] net49 0.00301f
C17706 _441_/a_2248_156# net49 0.048164f
C17707 _073_ _122_ 0.002157f
C17708 _053_ FILLER_0_7_59/a_36_472# 0.073877f
C17709 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001723f
C17710 _095_ FILLER_0_13_142/a_1380_472# 0.001782f
C17711 FILLER_0_21_142/a_484_472# _140_ 0.011035f
C17712 _074_ _068_ 0.011897f
C17713 _210_/a_255_603# vss 0.001246f
C17714 _250_/a_36_68# state\[1\] 0.103037f
C17715 FILLER_0_18_2/a_572_375# net44 0.072627f
C17716 trim_val\[3\] _441_/a_448_472# 0.00469f
C17717 _028_ FILLER_0_6_47/a_2724_472# 0.023218f
C17718 trim_val\[2\] net68 0.010894f
C17719 _013_ net26 0.174966f
C17720 _413_/a_36_151# FILLER_0_3_204/a_124_375# 0.035849f
C17721 FILLER_0_3_142/a_36_472# _443_/a_36_151# 0.001723f
C17722 _447_/a_796_472# net68 0.001593f
C17723 _447_/a_448_472# _036_ 0.015378f
C17724 _064_ _445_/a_796_472# 0.00673f
C17725 _293_/a_36_472# _105_ 0.004667f
C17726 _238_/a_67_603# trim_val\[3\] 0.024283f
C17727 FILLER_0_16_154/a_932_472# vdd 0.00549f
C17728 FILLER_0_16_154/a_484_472# vss 0.003464f
C17729 FILLER_0_3_172/a_2364_375# net21 0.004803f
C17730 _272_/a_36_472# net37 0.002669f
C17731 FILLER_0_8_239/a_124_375# vss 0.017196f
C17732 FILLER_0_8_239/a_36_472# vdd 0.079402f
C17733 _265_/a_244_68# vdd 0.022571f
C17734 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_124_375# 0.009654f
C17735 FILLER_0_7_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001723f
C17736 net41 _423_/a_36_151# 0.001134f
C17737 _142_ vss 0.121933f
C17738 net75 _082_ 0.417366f
C17739 FILLER_0_5_109/a_484_472# _154_ 0.039428f
C17740 net72 _183_ 0.093818f
C17741 FILLER_0_7_104/a_932_472# _134_ 0.004249f
C17742 FILLER_0_21_142/a_484_472# FILLER_0_21_150/a_36_472# 0.013277f
C17743 net75 FILLER_0_8_247/a_36_472# 0.002992f
C17744 result[9] FILLER_0_24_274/a_1020_375# 0.001657f
C17745 net38 FILLER_0_8_24/a_484_472# 0.001223f
C17746 _405_/a_67_603# net40 0.015326f
C17747 _112_ vdd 0.086153f
C17748 FILLER_0_7_104/a_36_472# vss 0.002797f
C17749 FILLER_0_7_104/a_484_472# vdd 0.021325f
C17750 net32 _419_/a_2665_112# 0.027035f
C17751 _118_ _124_ 0.652002f
C17752 fanout64/a_36_160# vdd 0.010802f
C17753 FILLER_0_12_136/a_572_375# state\[2\] 0.001955f
C17754 FILLER_0_12_136/a_1468_375# net53 0.002709f
C17755 net73 FILLER_0_18_107/a_932_472# 0.016711f
C17756 _430_/a_448_472# net21 0.03842f
C17757 _120_ net14 0.024442f
C17758 net75 _426_/a_448_472# 0.041705f
C17759 _081_ FILLER_0_6_177/a_124_375# 0.005524f
C17760 output32/a_224_472# _419_/a_1308_423# 0.005111f
C17761 _346_/a_49_472# _098_ 0.028579f
C17762 net26 FILLER_0_21_28/a_2812_375# 0.001905f
C17763 FILLER_0_18_107/a_2812_375# vss 0.002392f
C17764 FILLER_0_18_107/a_3260_375# vdd 0.004983f
C17765 FILLER_0_16_107/a_484_472# net14 0.001528f
C17766 output15/a_224_472# vdd 0.025731f
C17767 output20/a_224_472# net61 0.177946f
C17768 net41 _064_ 0.301777f
C17769 net52 FILLER_0_9_72/a_484_472# 0.049391f
C17770 _093_ _131_ 0.254316f
C17771 FILLER_0_14_107/a_124_375# _451_/a_36_151# 0.059049f
C17772 _116_ _056_ 0.30649f
C17773 net29 _102_ 0.056837f
C17774 output9/a_224_472# net82 0.003636f
C17775 _163_ _160_ 0.120564f
C17776 net27 FILLER_0_12_236/a_124_375# 0.044776f
C17777 output45/a_224_472# net46 0.005906f
C17778 _433_/a_2665_112# _145_ 0.018359f
C17779 _086_ _134_ 0.020487f
C17780 FILLER_0_18_37/a_932_472# vdd 0.01019f
C17781 fanout68/a_36_113# net69 0.046009f
C17782 net34 vss 0.481379f
C17783 net54 FILLER_0_20_107/a_36_472# 0.050184f
C17784 FILLER_0_16_241/a_124_375# net36 0.004069f
C17785 _375_/a_36_68# _161_ 0.028567f
C17786 FILLER_0_16_89/a_1468_375# vss 0.048986f
C17787 FILLER_0_16_89/a_36_472# vdd 0.040085f
C17788 _429_/a_2665_112# _098_ 0.003225f
C17789 ctln[2] FILLER_0_1_266/a_484_472# 0.019076f
C17790 net41 output41/a_224_472# 0.008587f
C17791 _196_/a_36_160# mask\[1\] 0.003254f
C17792 FILLER_0_24_274/a_932_472# vss 0.001001f
C17793 fanout82/a_36_113# calibrate 0.004982f
C17794 _104_ _011_ 0.021454f
C17795 _425_/a_36_151# _122_ 0.063131f
C17796 _425_/a_448_472# calibrate 0.105581f
C17797 ctln[7] _442_/a_2248_156# 0.006094f
C17798 net75 _265_/a_244_68# 0.046186f
C17799 _079_ _088_ 0.012529f
C17800 _289_/a_36_472# mask\[2\] 0.006392f
C17801 FILLER_0_4_49/a_484_472# _160_ 0.001336f
C17802 _053_ _359_/a_1492_488# 0.001437f
C17803 _233_/a_36_160# net67 0.001315f
C17804 _394_/a_56_524# _174_ 0.015122f
C17805 _011_ _422_/a_1308_423# 0.001997f
C17806 net50 fanout67/a_36_160# 0.007195f
C17807 ctlp[3] _107_ 0.132316f
C17808 fanout70/a_36_113# _095_ 0.003087f
C17809 _086_ FILLER_0_6_177/a_124_375# 0.043788f
C17810 _025_ FILLER_0_22_107/a_484_472# 0.00892f
C17811 _091_ FILLER_0_15_180/a_36_472# 0.00375f
C17812 net75 _112_ 0.041092f
C17813 FILLER_0_24_96/a_36_472# vdd 0.094828f
C17814 net20 FILLER_0_3_221/a_1468_375# 0.007234f
C17815 _414_/a_1308_423# net21 0.06986f
C17816 output33/a_224_472# vss 0.05089f
C17817 _320_/a_36_472# _055_ 0.001393f
C17818 net16 _402_/a_1296_93# 0.053493f
C17819 _072_ FILLER_0_10_214/a_124_375# 0.033245f
C17820 _245_/a_234_472# _067_ 0.005071f
C17821 _016_ FILLER_0_12_124/a_124_375# 0.007335f
C17822 output14/a_224_472# FILLER_0_0_130/a_124_375# 0.00515f
C17823 _076_ _062_ 0.978627f
C17824 _186_ net17 0.001172f
C17825 FILLER_0_22_177/a_572_375# mask\[6\] 0.002657f
C17826 net47 _386_/a_848_380# 0.003045f
C17827 _004_ net28 0.082388f
C17828 _413_/a_1000_472# vdd 0.002781f
C17829 output26/a_224_472# FILLER_0_23_44/a_932_472# 0.0323f
C17830 _379_/a_244_68# _160_ 0.001202f
C17831 net18 _416_/a_796_472# 0.007144f
C17832 FILLER_0_15_142/a_36_472# _427_/a_36_151# 0.001723f
C17833 _126_ cal_count\[3\] 0.418508f
C17834 net57 _097_ 0.100409f
C17835 _094_ _007_ 0.170362f
C17836 _449_/a_448_472# vdd 0.007757f
C17837 _449_/a_36_151# vss 0.014774f
C17838 FILLER_0_12_220/a_484_472# vdd 0.002383f
C17839 FILLER_0_12_220/a_36_472# vss 0.023702f
C17840 FILLER_0_10_247/a_124_375# _100_ 0.001804f
C17841 input1/a_36_113# net1 0.003795f
C17842 net55 FILLER_0_18_37/a_1468_375# 0.009059f
C17843 FILLER_0_18_139/a_1380_472# net23 0.013087f
C17844 FILLER_0_4_107/a_932_472# _160_ 0.014254f
C17845 _322_/a_124_24# net74 0.05722f
C17846 _426_/a_2560_156# net64 0.00801f
C17847 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_36_472# 0.001723f
C17848 net35 _434_/a_2248_156# 0.026885f
C17849 _414_/a_2665_112# vdd 0.006496f
C17850 FILLER_0_17_72/a_1020_375# vss 0.005441f
C17851 FILLER_0_17_72/a_1468_375# vdd 0.003316f
C17852 FILLER_0_8_37/a_484_472# vss 0.001267f
C17853 _308_/a_124_24# _439_/a_2248_156# 0.01963f
C17854 _004_ FILLER_0_10_247/a_124_375# 0.004573f
C17855 _412_/a_2248_156# fanout59/a_36_160# 0.007753f
C17856 _053_ FILLER_0_6_90/a_36_472# 0.002495f
C17857 result[2] _416_/a_36_151# 0.010509f
C17858 FILLER_0_8_247/a_124_375# calibrate 0.008393f
C17859 fanout54/a_36_160# net54 0.018583f
C17860 FILLER_0_15_142/a_484_472# _427_/a_36_151# 0.001723f
C17861 FILLER_0_8_107/a_36_472# _133_ 0.00589f
C17862 net35 _213_/a_67_603# 0.012955f
C17863 mask\[8\] _213_/a_255_603# 0.002776f
C17864 _231_/a_244_68# _059_ 0.004384f
C17865 _056_ _117_ 0.065147f
C17866 FILLER_0_22_86/a_124_375# vdd 0.024158f
C17867 output44/a_224_472# FILLER_0_18_2/a_124_375# 0.001168f
C17868 _116_ FILLER_0_12_196/a_124_375# 0.005332f
C17869 FILLER_0_13_100/a_36_472# vss 0.003094f
C17870 FILLER_0_4_197/a_1468_375# vdd 0.019672f
C17871 net38 _450_/a_1040_527# 0.027925f
C17872 _127_ _059_ 0.002878f
C17873 _419_/a_1308_423# vdd 0.007543f
C17874 result[9] net30 0.231442f
C17875 _430_/a_1308_423# net36 0.003317f
C17876 FILLER_0_5_117/a_36_472# FILLER_0_4_107/a_1020_375# 0.001684f
C17877 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_124_375# 0.001597f
C17878 clk net59 0.052607f
C17879 net80 FILLER_0_22_177/a_36_472# 0.018848f
C17880 net16 _033_ 0.042852f
C17881 FILLER_0_9_223/a_36_472# vss 0.019592f
C17882 FILLER_0_18_107/a_572_375# net14 0.00258f
C17883 FILLER_0_15_59/a_484_472# vdd 0.010447f
C17884 FILLER_0_15_59/a_36_472# vss 0.00459f
C17885 net18 FILLER_0_11_282/a_124_375# 0.042342f
C17886 fanout66/a_36_113# FILLER_0_3_54/a_36_472# 0.001645f
C17887 net82 _370_/a_848_380# 0.014538f
C17888 _453_/a_36_151# _042_ 0.035846f
C17889 FILLER_0_17_72/a_2724_472# _136_ 0.03065f
C17890 _431_/a_1204_472# _136_ 0.007382f
C17891 output24/a_224_472# vss 0.004078f
C17892 _210_/a_255_603# mask\[7\] 0.001329f
C17893 _443_/a_2665_112# net59 0.0434f
C17894 _017_ vdd 0.26981f
C17895 _413_/a_36_151# vss 0.003285f
C17896 cal_count\[2\] _452_/a_2225_156# 0.003086f
C17897 net15 _441_/a_448_472# 0.049213f
C17898 net59 FILLER_0_3_212/a_36_472# 0.058623f
C17899 output46/a_224_472# net44 0.003804f
C17900 mask\[2\] vss 0.536426f
C17901 FILLER_0_1_266/a_36_472# net19 0.07227f
C17902 _437_/a_1000_472# vdd 0.001777f
C17903 _441_/a_2560_156# _164_ 0.049213f
C17904 net47 _365_/a_36_68# 0.020511f
C17905 _449_/a_448_472# net72 0.01383f
C17906 _431_/a_36_151# FILLER_0_16_115/a_36_472# 0.004847f
C17907 _122_ _121_ 0.034975f
C17908 FILLER_0_7_195/a_36_472# calibrate 0.010951f
C17909 FILLER_0_4_213/a_124_375# vss 0.006145f
C17910 FILLER_0_4_213/a_572_375# vdd 0.026692f
C17911 FILLER_0_7_72/a_1916_375# vss 0.001259f
C17912 net15 _440_/a_1204_472# 0.01349f
C17913 _057_ net56 0.002158f
C17914 net54 _436_/a_2248_156# 0.043158f
C17915 net55 FILLER_0_17_72/a_124_375# 0.019544f
C17916 net62 result[3] 0.451989f
C17917 net15 _439_/a_36_151# 0.068183f
C17918 FILLER_0_22_177/a_124_375# _023_ 0.001195f
C17919 net79 _018_ 0.069992f
C17920 _446_/a_1308_423# net66 0.005976f
C17921 net47 FILLER_0_5_148/a_124_375# 0.008947f
C17922 FILLER_0_24_63/a_36_472# ctlp[9] 0.012298f
C17923 _064_ _446_/a_2560_156# 0.029586f
C17924 _250_/a_36_68# vdd 0.014409f
C17925 _032_ vdd 0.174834f
C17926 _341_/a_257_69# _137_ 0.004351f
C17927 FILLER_0_7_72/a_932_472# vss 0.002763f
C17928 FILLER_0_23_44/a_36_472# vss 0.002194f
C17929 FILLER_0_23_44/a_484_472# vdd 0.003276f
C17930 _077_ FILLER_0_10_94/a_36_472# 0.001114f
C17931 _141_ FILLER_0_22_128/a_3172_472# 0.01947f
C17932 net54 FILLER_0_18_139/a_124_375# 0.002807f
C17933 FILLER_0_4_152/a_124_375# net57 0.001947f
C17934 _077_ _453_/a_1000_472# 0.033726f
C17935 FILLER_0_21_125/a_572_375# vdd -0.013698f
C17936 FILLER_0_20_193/a_124_375# _098_ 0.009717f
C17937 FILLER_0_5_72/a_124_375# trim_mask\[1\] 0.010758f
C17938 FILLER_0_5_72/a_1468_375# _029_ 0.007876f
C17939 net15 FILLER_0_6_47/a_1828_472# 0.014911f
C17940 _091_ _429_/a_2560_156# 0.001502f
C17941 FILLER_0_6_47/a_1020_375# vdd 0.016637f
C17942 net72 FILLER_0_15_59/a_484_472# 0.008749f
C17943 _189_/a_67_603# _100_ 0.002818f
C17944 net58 result[0] 0.443436f
C17945 net26 _423_/a_448_472# 0.011612f
C17946 net34 mask\[7\] 0.901671f
C17947 _276_/a_36_160# vss 0.02914f
C17948 FILLER_0_18_171/a_36_472# mask\[3\] 0.00262f
C17949 vdd _450_/a_3129_107# 0.039939f
C17950 output7/a_224_472# vss 0.00746f
C17951 ctln[2] vss 0.256543f
C17952 FILLER_0_13_228/a_124_375# _043_ 0.133079f
C17953 FILLER_0_7_104/a_1468_375# _154_ 0.003683f
C17954 _057_ _060_ 0.033334f
C17955 net17 net43 0.144179f
C17956 cal_count\[3\] _453_/a_36_151# 0.023915f
C17957 _422_/a_36_151# _108_ 0.062205f
C17958 output44/a_224_472# net17 0.07836f
C17959 ctln[4] FILLER_0_1_204/a_124_375# 0.008283f
C17960 _370_/a_848_380# FILLER_0_5_136/a_124_375# 0.014613f
C17961 output32/a_224_472# net19 0.08441f
C17962 FILLER_0_9_60/a_36_472# vdd 0.08419f
C17963 FILLER_0_9_60/a_572_375# vss 0.022532f
C17964 net41 _444_/a_2248_156# 0.028267f
C17965 _020_ vdd 0.194776f
C17966 _096_ state\[1\] 0.083332f
C17967 net26 _424_/a_1204_472# 0.00194f
C17968 FILLER_0_15_290/a_36_472# vss 0.010015f
C17969 _065_ ctln[8] 0.193903f
C17970 net41 _446_/a_448_472# 0.040165f
C17971 _106_ ctlp[1] 0.002631f
C17972 output43/a_224_472# net46 0.0215f
C17973 _430_/a_2665_112# FILLER_0_17_218/a_572_375# 0.002362f
C17974 net66 _160_ 0.097885f
C17975 _086_ _311_/a_66_473# 0.007295f
C17976 output11/a_224_472# _000_ 0.006606f
C17977 ctln[8] FILLER_0_0_96/a_36_472# 0.012298f
C17978 _028_ FILLER_0_6_90/a_36_472# 0.013106f
C17979 FILLER_0_11_109/a_36_472# _134_ 0.007739f
C17980 FILLER_0_21_28/a_1380_472# _012_ 0.004453f
C17981 fanout70/a_36_113# net74 0.002663f
C17982 _010_ net19 0.408364f
C17983 _445_/a_36_151# _034_ 0.005488f
C17984 cal_itt\[1\] FILLER_0_3_221/a_1468_375# 0.020427f
C17985 trim_mask\[1\] _166_ 0.124855f
C17986 FILLER_0_11_109/a_124_375# vdd 0.079069f
C17987 _163_ _156_ 0.001616f
C17988 _411_/a_2248_156# ctln[3] 0.001208f
C17989 _076_ _226_/a_860_68# 0.001752f
C17990 _093_ FILLER_0_17_104/a_932_472# 0.014431f
C17991 FILLER_0_2_93/a_124_375# vdd 0.008901f
C17992 _255_/a_224_552# _062_ 0.009032f
C17993 _432_/a_36_151# _333_/a_36_160# 0.032942f
C17994 net48 FILLER_0_7_233/a_124_375# 0.013455f
C17995 _086_ _374_/a_244_472# 0.001496f
C17996 FILLER_0_11_135/a_124_375# vdd 0.042201f
C17997 _372_/a_3662_472# _122_ 0.002653f
C17998 FILLER_0_17_282/a_36_472# vss 0.007765f
C17999 _448_/a_796_472# vdd 0.002153f
C18000 _074_ FILLER_0_5_172/a_36_472# 0.016713f
C18001 net58 output37/a_224_472# 0.099539f
C18002 FILLER_0_14_81/a_36_472# _095_ 0.014706f
C18003 net38 FILLER_0_20_2/a_572_375# 0.004413f
C18004 _093_ _137_ 0.201779f
C18005 FILLER_0_14_107/a_1468_375# vdd 0.007687f
C18006 mask\[8\] mask\[9\] 0.078756f
C18007 FILLER_0_22_177/a_1468_375# vdd -0.007187f
C18008 net48 vdd 0.35704f
C18009 _167_ _160_ 0.157458f
C18010 net4 FILLER_0_12_220/a_36_472# 0.019348f
C18011 mask\[5\] _049_ 0.008296f
C18012 _423_/a_36_151# FILLER_0_23_44/a_572_375# 0.059049f
C18013 output23/a_224_472# FILLER_0_24_130/a_124_375# 0.006051f
C18014 FILLER_0_19_125/a_124_375# FILLER_0_18_107/a_2276_472# 0.001684f
C18015 output36/a_224_472# net19 0.106928f
C18016 _151_ net14 0.009212f
C18017 _086_ _331_/a_244_472# 0.001991f
C18018 net36 FILLER_0_15_212/a_1468_375# 0.005276f
C18019 FILLER_0_3_221/a_36_472# vdd 0.018263f
C18020 FILLER_0_3_221/a_1468_375# vss 0.004085f
C18021 _073_ net8 0.206839f
C18022 fanout73/a_36_113# vss 0.01873f
C18023 net16 FILLER_0_16_37/a_124_375# 0.033245f
C18024 _162_ vdd 0.073371f
C18025 net80 _023_ 0.261119f
C18026 _334_/a_36_160# FILLER_0_17_104/a_1468_375# 0.027706f
C18027 mask\[4\] FILLER_0_18_177/a_3172_472# 0.014657f
C18028 _072_ _055_ 0.083351f
C18029 FILLER_0_18_177/a_3172_472# net22 0.037136f
C18030 _131_ _120_ 0.191602f
C18031 _003_ net76 0.080782f
C18032 FILLER_0_19_55/a_36_472# _216_/a_67_603# 0.00254f
C18033 FILLER_0_5_54/a_572_375# trim_mask\[1\] 0.011664f
C18034 result[1] result[2] 0.072492f
C18035 _093_ _438_/a_1308_423# 0.001057f
C18036 net52 net49 0.092082f
C18037 _414_/a_1000_472# net22 0.001649f
C18038 FILLER_0_16_107/a_484_472# _131_ 0.008223f
C18039 FILLER_0_12_136/a_1468_375# _071_ 0.002023f
C18040 mask\[8\] FILLER_0_22_86/a_1380_472# 0.012151f
C18041 net35 FILLER_0_22_86/a_932_472# 0.007806f
C18042 _137_ FILLER_0_15_180/a_572_375# 0.028083f
C18043 net52 _442_/a_2248_156# 0.022954f
C18044 net20 FILLER_0_7_233/a_36_472# 0.035074f
C18045 net76 net21 0.041873f
C18046 FILLER_0_16_89/a_124_375# _040_ 0.006315f
C18047 _404_/a_36_472# _183_ 0.002637f
C18048 _430_/a_2560_156# net63 0.009628f
C18049 trim[4] FILLER_0_8_2/a_124_375# 0.028454f
C18050 _114_ trim_mask\[0\] 0.021887f
C18051 _027_ FILLER_0_18_76/a_124_375# 0.001285f
C18052 FILLER_0_15_235/a_572_375# FILLER_0_14_235/a_572_375# 0.05841f
C18053 FILLER_0_9_28/a_484_472# net41 0.042989f
C18054 _131_ _403_/a_224_472# 0.003274f
C18055 net50 trim_mask\[1\] 0.502622f
C18056 FILLER_0_9_223/a_36_472# net4 0.014911f
C18057 _205_/a_36_160# vdd 0.016131f
C18058 _057_ _095_ 0.001346f
C18059 FILLER_0_7_72/a_2364_375# net14 0.005919f
C18060 _053_ _251_/a_906_472# 0.001696f
C18061 FILLER_0_21_206/a_124_375# _434_/a_2665_112# 0.002259f
C18062 FILLER_0_18_177/a_2812_375# vdd 0.003766f
C18063 net15 FILLER_0_7_59/a_124_375# 0.004662f
C18064 net20 vss 1.402494f
C18065 result[4] net18 0.048179f
C18066 _081_ _080_ 0.003905f
C18067 result[8] net35 0.001362f
C18068 _339_/a_36_160# vss 0.027338f
C18069 _104_ _198_/a_67_603# 0.007168f
C18070 FILLER_0_18_2/a_2276_472# vss 0.001865f
C18071 _346_/a_257_69# _141_ 0.002092f
C18072 net32 net78 0.055231f
C18073 net19 vdd 2.167778f
C18074 _043_ net14 0.037706f
C18075 net20 _298_/a_224_472# 0.001861f
C18076 _076_ FILLER_0_8_156/a_572_375# 0.010751f
C18077 _010_ _009_ 0.030637f
C18078 FILLER_0_8_138/a_124_375# _077_ 0.007238f
C18079 _013_ FILLER_0_18_53/a_572_375# 0.015534f
C18080 _136_ _451_/a_1697_156# 0.001053f
C18081 net75 net48 0.10167f
C18082 FILLER_0_23_88/a_124_375# vdd 0.03583f
C18083 _453_/a_2560_156# vss 0.00337f
C18084 output16/a_224_472# _447_/a_36_151# 0.200384f
C18085 mask\[6\] vdd 0.573103f
C18086 _417_/a_2248_156# _006_ 0.039121f
C18087 net69 FILLER_0_3_78/a_484_472# 0.002068f
C18088 _439_/a_36_151# FILLER_0_6_47/a_2364_375# 0.002807f
C18089 FILLER_0_7_72/a_484_472# net52 0.049487f
C18090 FILLER_0_18_107/a_3260_375# FILLER_0_19_134/a_124_375# 0.026339f
C18091 net81 FILLER_0_12_236/a_484_472# 0.001419f
C18092 _131_ FILLER_0_9_105/a_572_375# 0.031928f
C18093 input2/a_36_113# vdd 0.096633f
C18094 _142_ _141_ 0.200324f
C18095 FILLER_0_6_79/a_36_472# vdd 0.087807f
C18096 FILLER_0_6_79/a_124_375# vss 0.007008f
C18097 net73 net71 0.033964f
C18098 FILLER_0_16_73/a_572_375# vdd 0.005054f
C18099 net47 _154_ 0.055128f
C18100 net41 net50 0.002438f
C18101 _176_ _394_/a_1936_472# 0.001255f
C18102 cal_count\[3\] _060_ 0.007037f
C18103 _079_ _260_/a_36_68# 0.043596f
C18104 _144_ _022_ 0.139742f
C18105 net53 _427_/a_1000_472# 0.008132f
C18106 FILLER_0_4_177/a_36_472# _163_ 0.002787f
C18107 FILLER_0_12_236/a_484_472# _060_ 0.002678f
C18108 FILLER_0_1_266/a_484_472# vss 0.001113f
C18109 _015_ FILLER_0_8_247/a_124_375# 0.00706f
C18110 FILLER_0_1_204/a_124_375# net21 0.008041f
C18111 net18 FILLER_0_9_282/a_36_472# 0.041571f
C18112 net3 _043_ 0.004313f
C18113 FILLER_0_3_204/a_124_375# vss 0.017795f
C18114 _360_/a_36_160# _153_ 0.006561f
C18115 _093_ net56 0.040124f
C18116 _128_ _062_ 0.025708f
C18117 mask\[8\] _352_/a_49_472# 0.002573f
C18118 FILLER_0_3_54/a_36_472# vdd 0.00827f
C18119 _114_ FILLER_0_13_142/a_572_375# 0.00191f
C18120 _359_/a_1044_488# _152_ 0.001339f
C18121 _095_ FILLER_0_13_72/a_572_375# 0.003559f
C18122 cal_itt\[2\] net8 0.057335f
C18123 net75 net19 1.345314f
C18124 mask\[8\] net35 2.631701f
C18125 net3 _185_ 0.004236f
C18126 _008_ _418_/a_2248_156# 0.047066f
C18127 _450_/a_1284_156# _039_ 0.001226f
C18128 _176_ _171_ 0.049997f
C18129 _450_/a_3129_107# cal_count\[0\] 0.020971f
C18130 net36 FILLER_0_15_235/a_572_375# 0.083299f
C18131 net65 FILLER_0_3_172/a_124_375# 0.021073f
C18132 FILLER_0_8_107/a_124_375# _134_ 0.007753f
C18133 FILLER_0_12_2/a_484_472# net38 0.002706f
C18134 net1 net8 0.00497f
C18135 net15 FILLER_0_9_72/a_36_472# 0.006905f
C18136 _059_ net23 0.265909f
C18137 _402_/a_728_93# _179_ 0.011717f
C18138 ctln[2] net4 0.039098f
C18139 net81 net65 0.083316f
C18140 result[9] _417_/a_2665_112# 0.060365f
C18141 _072_ _058_ 0.029688f
C18142 FILLER_0_14_91/a_124_375# en_co_clk 0.006788f
C18143 _174_ cal_count\[2\] 0.004821f
C18144 _274_/a_36_68# FILLER_0_12_220/a_484_472# 0.001048f
C18145 output24/a_224_472# _436_/a_1308_423# 0.005632f
C18146 net34 _295_/a_36_472# 0.032003f
C18147 _077_ FILLER_0_10_78/a_36_472# 0.002486f
C18148 net55 _453_/a_2248_156# 0.001546f
C18149 FILLER_0_12_136/a_484_472# vss 0.007054f
C18150 FILLER_0_12_136/a_932_472# vdd 0.005266f
C18151 FILLER_0_10_214/a_36_472# _247_/a_36_160# 0.004828f
C18152 FILLER_0_20_177/a_124_375# FILLER_0_20_169/a_124_375# 0.003732f
C18153 _431_/a_1456_156# net73 0.001304f
C18154 mask\[0\] FILLER_0_13_228/a_36_472# 0.002986f
C18155 _077_ FILLER_0_8_107/a_36_472# 0.007552f
C18156 _130_ FILLER_0_11_124/a_124_375# 0.001943f
C18157 _009_ vdd 0.693198f
C18158 FILLER_0_17_142/a_36_472# _137_ 0.003953f
C18159 output10/a_224_472# vdd 0.107357f
C18160 _126_ _120_ 0.055349f
C18161 _274_/a_2552_68# _070_ 0.001238f
C18162 _111_ vdd 0.3227f
C18163 _423_/a_2248_156# _012_ 0.011646f
C18164 FILLER_0_21_142/a_484_472# _098_ 0.001158f
C18165 _088_ _269_/a_36_472# 0.004438f
C18166 _114_ FILLER_0_11_101/a_124_375# 0.013348f
C18167 mask\[3\] net21 0.100738f
C18168 net54 _150_ 0.001162f
C18169 _164_ _166_ 0.002368f
C18170 FILLER_0_8_138/a_36_472# _070_ 0.001342f
C18171 _096_ vdd 0.557569f
C18172 FILLER_0_21_286/a_36_472# _420_/a_36_151# 0.059367f
C18173 _327_/a_36_472# FILLER_0_12_136/a_36_472# 0.096379f
C18174 FILLER_0_1_98/a_124_375# trim_val\[3\] 0.001628f
C18175 FILLER_0_3_172/a_124_375# net59 0.001045f
C18176 net31 net32 0.023293f
C18177 _421_/a_36_151# net18 0.00659f
C18178 FILLER_0_19_111/a_36_472# vdd 0.034386f
C18179 FILLER_0_19_111/a_572_375# vss 0.003337f
C18180 net81 net59 0.074175f
C18181 net79 FILLER_0_12_220/a_36_472# 0.005464f
C18182 FILLER_0_14_50/a_36_472# _095_ 0.013704f
C18183 _292_/a_36_160# _098_ 0.048643f
C18184 FILLER_0_19_187/a_572_375# vdd 0.023383f
C18185 fanout60/a_36_160# FILLER_0_17_282/a_124_375# 0.005489f
C18186 _446_/a_2665_112# _160_ 0.013745f
C18187 fanout78/a_36_113# vdd 0.061637f
C18188 _144_ _354_/a_665_69# 0.001518f
C18189 net14 FILLER_0_10_94/a_572_375# 0.047331f
C18190 _102_ _419_/a_2248_156# 0.001679f
C18191 FILLER_0_21_125/a_36_472# _436_/a_36_151# 0.001695f
C18192 ctlp[3] _422_/a_2248_156# 0.001888f
C18193 _098_ _043_ 0.032706f
C18194 FILLER_0_18_76/a_484_472# _438_/a_36_151# 0.001723f
C18195 net73 fanout71/a_36_113# 0.004833f
C18196 _177_ _040_ 0.061289f
C18197 net47 _278_/a_36_160# 0.001838f
C18198 FILLER_0_5_181/a_36_472# vss 0.001068f
C18199 cal_count\[3\] _095_ 0.06065f
C18200 FILLER_0_21_28/a_1468_375# vdd -0.008892f
C18201 FILLER_0_21_125/a_572_375# _433_/a_36_151# 0.059049f
C18202 FILLER_0_3_172/a_36_472# vss 0.001848f
C18203 FILLER_0_3_172/a_484_472# vdd 0.007258f
C18204 _386_/a_124_24# vss 0.009702f
C18205 _386_/a_848_380# vdd 0.054849f
C18206 output31/a_224_472# net30 0.149277f
C18207 _443_/a_36_151# _081_ 0.001923f
C18208 net4 FILLER_0_3_221/a_1468_375# 0.006974f
C18209 _115_ _118_ 1.045555f
C18210 FILLER_0_24_96/a_36_472# net24 0.028193f
C18211 FILLER_0_14_81/a_36_472# cal_count\[1\] 0.034486f
C18212 _264_/a_224_472# _084_ 0.007508f
C18213 FILLER_0_13_212/a_1380_472# _043_ 0.014431f
C18214 mask\[5\] _091_ 0.048311f
C18215 _093_ FILLER_0_18_107/a_2276_472# 0.001996f
C18216 fanout53/a_36_160# net36 0.028652f
C18217 _359_/a_36_488# _133_ 0.04287f
C18218 FILLER_0_18_100/a_124_375# vss 0.025563f
C18219 FILLER_0_18_100/a_36_472# vdd 0.012574f
C18220 _088_ FILLER_0_3_172/a_3172_472# 0.004381f
C18221 FILLER_0_22_177/a_124_375# net33 0.013581f
C18222 _091_ FILLER_0_18_209/a_572_375# 0.001343f
C18223 _087_ _163_ 0.004829f
C18224 _106_ _201_/a_67_603# 0.00327f
C18225 net12 net59 0.001028f
C18226 _449_/a_2665_112# cal_count\[3\] 0.001422f
C18227 mask\[9\] _026_ 0.002924f
C18228 _444_/a_1000_472# net47 0.036015f
C18229 _161_ _311_/a_66_473# 0.021817f
C18230 _091_ FILLER_0_12_220/a_124_375# 0.006907f
C18231 _120_ FILLER_0_10_107/a_124_375# 0.001834f
C18232 FILLER_0_10_214/a_124_375# vdd 0.018944f
C18233 _063_ _033_ 0.250192f
C18234 _442_/a_36_151# _031_ 0.013852f
C18235 net50 _164_ 0.080818f
C18236 _005_ _416_/a_1204_472# 0.014873f
C18237 FILLER_0_3_172/a_36_472# FILLER_0_2_171/a_124_375# 0.001723f
C18238 _053_ FILLER_0_7_104/a_36_472# 0.01752f
C18239 vss FILLER_0_4_91/a_484_472# 0.003328f
C18240 state\[0\] calibrate 0.001061f
C18241 FILLER_0_19_195/a_36_472# _434_/a_2248_156# 0.001731f
C18242 FILLER_0_14_81/a_124_375# _451_/a_3129_107# 0.009542f
C18243 FILLER_0_7_59/a_572_375# FILLER_0_6_47/a_1916_375# 0.05841f
C18244 _140_ _352_/a_665_69# 0.001363f
C18245 FILLER_0_3_142/a_124_375# _032_ 0.001153f
C18246 trimb[3] net43 0.221036f
C18247 _261_/a_36_160# FILLER_0_5_136/a_124_375# 0.003477f
C18248 _086_ _114_ 1.371271f
C18249 state\[1\] _055_ 0.067603f
C18250 fanout58/a_36_160# vdd 0.101571f
C18251 cal_itt\[1\] vss 0.327626f
C18252 cal_itt\[0\] vdd 0.438996f
C18253 _162_ _374_/a_36_68# 0.005729f
C18254 _095_ net40 0.674445f
C18255 net20 net4 0.650415f
C18256 FILLER_0_7_72/a_1020_375# FILLER_0_5_72/a_932_472# 0.001512f
C18257 FILLER_0_8_127/a_36_472# _058_ 0.003283f
C18258 net50 FILLER_0_5_72/a_1380_472# 0.002431f
C18259 trim_mask\[2\] FILLER_0_3_54/a_124_375# 0.015198f
C18260 _141_ mask\[2\] 0.084094f
C18261 net56 FILLER_0_17_142/a_36_472# 0.003603f
C18262 fanout55/a_36_160# vdd 0.016488f
C18263 valid net76 0.285892f
C18264 mask\[0\] _429_/a_1204_472# 0.005396f
C18265 _119_ _114_ 0.001581f
C18266 net55 FILLER_0_18_53/a_484_472# 0.012319f
C18267 _415_/a_36_151# FILLER_0_10_256/a_36_472# 0.004847f
C18268 _079_ net59 0.102335f
C18269 FILLER_0_7_233/a_36_472# vss 0.005354f
C18270 net38 _452_/a_1353_112# 0.005918f
C18271 _415_/a_2665_112# FILLER_0_9_290/a_124_375# 0.001597f
C18272 _321_/a_3126_472# _118_ 0.002754f
C18273 net63 FILLER_0_22_177/a_572_375# 0.001597f
C18274 FILLER_0_12_136/a_1468_375# net23 0.021046f
C18275 _193_/a_36_160# vdd 0.092266f
C18276 _401_/a_36_68# vdd 0.003745f
C18277 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3172_472# 0.013276f
C18278 sample vss 0.276162f
C18279 net72 FILLER_0_21_28/a_1468_375# 0.001823f
C18280 _068_ _163_ 0.04926f
C18281 FILLER_0_20_177/a_484_472# _098_ 0.009817f
C18282 _077_ _439_/a_36_151# 0.035432f
C18283 _104_ output19/a_224_472# 0.064818f
C18284 _103_ _418_/a_1000_472# 0.006239f
C18285 result[8] FILLER_0_21_206/a_36_472# 0.001292f
C18286 _115_ _068_ 0.889978f
C18287 _376_/a_36_160# FILLER_0_6_90/a_124_375# 0.005705f
C18288 _365_/a_36_68# vdd 0.004308f
C18289 _120_ _453_/a_36_151# 0.001848f
C18290 cal_count\[1\] _451_/a_3129_107# 0.028519f
C18291 ctlp[0] net43 0.003786f
C18292 result[7] _102_ 0.010818f
C18293 net50 FILLER_0_8_24/a_36_472# 0.015187f
C18294 _176_ _183_ 0.024038f
C18295 _427_/a_2665_112# state\[1\] 0.021573f
C18296 _093_ FILLER_0_17_72/a_484_472# 0.008637f
C18297 vdd FILLER_0_5_148/a_124_375# -0.011369f
C18298 FILLER_0_6_177/a_36_472# vss 0.001617f
C18299 FILLER_0_6_177/a_484_472# vdd 0.007991f
C18300 result[6] output19/a_224_472# 0.001526f
C18301 FILLER_0_17_72/a_124_375# FILLER_0_15_72/a_36_472# 0.001512f
C18302 result[4] _417_/a_36_151# 0.010571f
C18303 _327_/a_36_472# vdd 0.00142f
C18304 net15 net25 0.013745f
C18305 net81 _429_/a_2665_112# 0.012675f
C18306 net74 FILLER_0_13_72/a_572_375# 0.012891f
C18307 net64 FILLER_0_12_236/a_484_472# 0.010321f
C18308 _442_/a_36_151# _371_/a_36_113# 0.001089f
C18309 FILLER_0_2_171/a_124_375# vss 0.049142f
C18310 FILLER_0_2_171/a_36_472# vdd 0.029996f
C18311 net75 cal_itt\[0\] 0.032053f
C18312 net63 FILLER_0_18_177/a_1916_375# 0.040551f
C18313 _077_ _039_ 0.104126f
C18314 FILLER_0_15_290/a_36_472# net79 0.04083f
C18315 _411_/a_36_151# net65 0.001415f
C18316 _411_/a_1308_423# _000_ 0.004012f
C18317 net64 _416_/a_36_151# 0.013586f
C18318 net15 net36 0.265646f
C18319 _021_ mask\[3\] 0.036781f
C18320 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_36_472# 0.001723f
C18321 net41 _054_ 0.035503f
C18322 FILLER_0_7_72/a_124_375# vss 0.044754f
C18323 _144_ FILLER_0_21_125/a_36_472# 0.008287f
C18324 net20 FILLER_0_13_212/a_1020_375# 0.003962f
C18325 net27 FILLER_0_9_270/a_484_472# 0.023461f
C18326 FILLER_0_4_152/a_124_375# FILLER_0_4_144/a_572_375# 0.012001f
C18327 _217_/a_36_160# FILLER_0_19_28/a_572_375# 0.058908f
C18328 _095_ FILLER_0_12_20/a_124_375# 0.001588f
C18329 FILLER_0_19_47/a_36_472# _013_ 0.03573f
C18330 _435_/a_2665_112# net21 0.067461f
C18331 _053_ FILLER_0_8_37/a_484_472# 0.002095f
C18332 _408_/a_56_524# _190_/a_36_160# 0.004025f
C18333 _098_ FILLER_0_19_171/a_1380_472# 0.001764f
C18334 net16 _182_ 0.05291f
C18335 FILLER_0_16_89/a_1380_472# net36 0.001657f
C18336 _428_/a_448_472# _017_ 0.056f
C18337 _428_/a_36_151# net53 0.001124f
C18338 net63 _092_ 0.008819f
C18339 FILLER_0_21_28/a_1468_375# _424_/a_36_151# 0.059049f
C18340 FILLER_0_16_57/a_484_472# cal_count\[1\] 0.001664f
C18341 result[9] _418_/a_2665_112# 0.053489f
C18342 net72 _401_/a_36_68# 0.006818f
C18343 net80 net33 0.037227f
C18344 _413_/a_448_472# net65 0.044062f
C18345 ctln[0] trim[2] 0.011834f
C18346 net32 net60 0.509175f
C18347 output25/a_224_472# _423_/a_2665_112# 0.001396f
C18348 _114_ net53 0.001275f
C18349 _131_ _043_ 0.047425f
C18350 net82 FILLER_0_3_172/a_1468_375# 0.010439f
C18351 FILLER_0_2_165/a_36_472# vdd -0.003333f
C18352 FILLER_0_2_165/a_124_375# vss 0.008386f
C18353 _397_/a_36_472# FILLER_0_17_72/a_1020_375# 0.001781f
C18354 fanout75/a_36_113# _317_/a_36_113# 0.001442f
C18355 net65 net64 0.119915f
C18356 _185_ _405_/a_67_603# 0.060789f
C18357 _008_ _102_ 0.027578f
C18358 _257_/a_36_472# _077_ 0.019883f
C18359 _076_ FILLER_0_6_231/a_572_375# 0.001647f
C18360 _328_/a_36_113# cal_count\[3\] 0.006392f
C18361 _369_/a_692_472# vdd 0.003899f
C18362 fanout63/a_36_160# mask\[2\] 0.026642f
C18363 ctln[6] vdd 0.116327f
C18364 net52 net47 0.039912f
C18365 _267_/a_36_472# _121_ 0.041237f
C18366 _394_/a_1336_472# _095_ 0.031869f
C18367 _137_ FILLER_0_16_154/a_124_375# 0.007998f
C18368 _028_ FILLER_0_7_104/a_36_472# 0.006408f
C18369 _077_ FILLER_0_8_156/a_36_472# 0.00563f
C18370 _189_/a_67_603# mask\[0\] 0.043158f
C18371 trim_mask\[2\] FILLER_0_4_91/a_484_472# 0.0022f
C18372 FILLER_0_16_73/a_36_472# _394_/a_1336_472# 0.00108f
C18373 _415_/a_36_151# output28/a_224_472# 0.229574f
C18374 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_36_472# 0.001963f
C18375 net34 ctlp[2] 0.953441f
C18376 FILLER_0_2_171/a_124_375# FILLER_0_2_165/a_124_375# 0.003598f
C18377 _062_ net14 0.003317f
C18378 FILLER_0_4_49/a_484_472# _440_/a_36_151# 0.006095f
C18379 output27/a_224_472# FILLER_0_9_282/a_572_375# 0.029138f
C18380 FILLER_0_18_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001597f
C18381 net15 _423_/a_2560_156# 0.007083f
C18382 _175_ _131_ 0.050098f
C18383 _429_/a_36_151# vdd 0.076815f
C18384 _413_/a_448_472# net59 0.059041f
C18385 FILLER_0_10_78/a_1020_375# vdd 0.002901f
C18386 result[8] output35/a_224_472# 0.016867f
C18387 _350_/a_665_69# net23 0.001468f
C18388 net39 FILLER_0_8_2/a_124_375# 0.008405f
C18389 FILLER_0_14_50/a_36_472# cal_count\[1\] 0.030015f
C18390 net61 _422_/a_2560_156# 0.010748f
C18391 net74 cal_count\[3\] 0.040777f
C18392 _095_ FILLER_0_13_80/a_124_375# 0.001989f
C18393 net35 _211_/a_36_160# 0.009886f
C18394 FILLER_0_7_72/a_1916_375# _053_ 0.013335f
C18395 _443_/a_448_472# _032_ 0.036717f
C18396 net82 _001_ 0.044461f
C18397 _316_/a_848_380# net37 0.01216f
C18398 output9/a_224_472# net81 0.02825f
C18399 _132_ _428_/a_796_472# 0.001472f
C18400 _105_ net78 0.004705f
C18401 net64 net59 0.005832f
C18402 _441_/a_36_151# FILLER_0_3_78/a_124_375# 0.035849f
C18403 ctlp[1] FILLER_0_21_286/a_124_375# 0.025059f
C18404 _093_ mask\[8\] 0.004026f
C18405 mask\[1\] FILLER_0_15_180/a_572_375# 0.011186f
C18406 FILLER_0_16_89/a_36_472# _176_ 0.012173f
C18407 FILLER_0_7_72/a_932_472# _053_ 0.01339f
C18408 FILLER_0_22_128/a_1468_375# vdd 0.016807f
C18409 FILLER_0_22_128/a_1020_375# vss 0.003747f
C18410 _428_/a_2665_112# _043_ 0.021483f
C18411 net18 result[3] 0.237732f
C18412 net20 net79 0.046876f
C18413 FILLER_0_1_98/a_36_472# vss 0.002275f
C18414 _449_/a_2665_112# FILLER_0_13_80/a_124_375# 0.010688f
C18415 _086_ _085_ 0.374127f
C18416 _424_/a_448_472# vss 0.002076f
C18417 _424_/a_1308_423# vdd 0.002386f
C18418 output33/a_224_472# ctlp[2] 0.00175f
C18419 _052_ _424_/a_2560_156# 0.003401f
C18420 net15 _030_ 0.355335f
C18421 _441_/a_2248_156# vdd -0.003818f
C18422 _441_/a_1204_472# vss 0.011996f
C18423 trim_val\[2\] vdd 0.160419f
C18424 trim_mask\[2\] vss 0.182675f
C18425 FILLER_0_11_64/a_124_375# vss 0.021069f
C18426 FILLER_0_11_64/a_36_472# vdd 0.015144f
C18427 _106_ _199_/a_36_160# 0.003376f
C18428 mask\[5\] FILLER_0_20_177/a_572_375# 0.013294f
C18429 net55 _452_/a_1353_112# 0.030679f
C18430 _008_ _198_/a_67_603# 0.012332f
C18431 trim_val\[4\] _241_/a_224_472# 0.003005f
C18432 _053_ FILLER_0_6_47/a_572_375# 0.008213f
C18433 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_572_375# 0.026339f
C18434 mask\[3\] FILLER_0_18_177/a_36_472# 0.005668f
C18435 _447_/a_796_472# vdd 0.001959f
C18436 trim_val\[3\] trim_mask\[3\] 0.48462f
C18437 _141_ _339_/a_36_160# 0.011118f
C18438 FILLER_0_7_72/a_1916_375# FILLER_0_5_88/a_36_472# 0.0027f
C18439 net76 FILLER_0_1_192/a_124_375# 0.00275f
C18440 _075_ _072_ 0.024301f
C18441 _406_/a_36_159# net47 0.034933f
C18442 FILLER_0_13_142/a_1468_375# _225_/a_36_160# 0.027706f
C18443 _430_/a_2665_112# mask\[2\] 0.028551f
C18444 _112_ _425_/a_1204_472# 0.001132f
C18445 net68 trim_val\[0\] 0.052045f
C18446 _439_/a_1000_472# vss 0.032923f
C18447 net31 FILLER_0_16_255/a_36_472# 0.003056f
C18448 net62 FILLER_0_13_290/a_36_472# 0.003157f
C18449 input3/a_36_113# vss 0.043862f
C18450 net4 cal_itt\[1\] 0.048147f
C18451 _428_/a_36_151# FILLER_0_11_109/a_36_472# 0.001221f
C18452 _181_ _402_/a_728_93# 0.064373f
C18453 _142_ FILLER_0_17_133/a_36_472# 0.069383f
C18454 mask\[9\] FILLER_0_18_76/a_124_375# 0.004592f
C18455 _232_/a_67_603# _160_ 0.001684f
C18456 net76 FILLER_0_3_172/a_1380_472# 0.015215f
C18457 _414_/a_36_151# net76 0.037157f
C18458 _426_/a_36_151# FILLER_0_8_247/a_484_472# 0.001723f
C18459 output42/a_224_472# output6/a_224_472# 0.292612f
C18460 _055_ vdd 0.406945f
C18461 net4 FILLER_0_7_233/a_36_472# 0.036721f
C18462 _114_ FILLER_0_11_109/a_36_472# 0.023029f
C18463 mask\[7\] vss 0.85153f
C18464 net56 FILLER_0_18_139/a_36_472# 0.002172f
C18465 FILLER_0_10_28/a_36_472# net47 0.002783f
C18466 _091_ FILLER_0_18_177/a_572_375# 0.004285f
C18467 _428_/a_36_151# FILLER_0_14_107/a_36_472# 0.02628f
C18468 net26 _012_ 0.066032f
C18469 _155_ trim_mask\[1\] 0.006536f
C18470 fanout60/a_36_160# vdd 0.090968f
C18471 _148_ vss 0.025751f
C18472 _276_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C18473 _190_/a_36_160# _450_/a_36_151# 0.002486f
C18474 _350_/a_49_472# _049_ 0.025442f
C18475 output8/a_224_472# ctln[1] 0.020259f
C18476 _126_ _043_ 0.128227f
C18477 net4 vss 0.774455f
C18478 mask\[5\] FILLER_0_19_171/a_1468_375# 0.007169f
C18479 FILLER_0_18_107/a_2812_375# FILLER_0_17_133/a_36_472# 0.001543f
C18480 _430_/a_1000_472# net36 0.001836f
C18481 FILLER_0_15_10/a_124_375# vdd 0.021578f
C18482 _114_ FILLER_0_14_107/a_36_472# 0.00191f
C18483 net41 _217_/a_36_160# 0.004517f
C18484 FILLER_0_7_72/a_3260_375# net14 0.025344f
C18485 net19 _416_/a_2248_156# 0.024466f
C18486 _190_/a_36_160# _043_ 0.06415f
C18487 _269_/a_36_472# _260_/a_36_68# 0.002875f
C18488 _311_/a_1212_473# vdd 0.001387f
C18489 FILLER_0_15_142/a_124_375# vdd -0.003809f
C18490 _265_/a_244_68# _082_ 0.031951f
C18491 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_1020_375# 0.026339f
C18492 _428_/a_36_151# _451_/a_36_151# 0.003608f
C18493 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_36_472# 0.002296f
C18494 output31/a_224_472# _417_/a_2665_112# 0.011048f
C18495 net24 FILLER_0_23_88/a_124_375# 0.020193f
C18496 _154_ vdd 0.639978f
C18497 _313_/a_67_603# vdd -0.002183f
C18498 _343_/a_49_472# vdd 0.089707f
C18499 FILLER_0_9_28/a_3260_375# _077_ 0.01495f
C18500 _114_ _161_ 0.024297f
C18501 net41 _035_ 0.048883f
C18502 ctln[7] vdd 0.359832f
C18503 net51 output6/a_224_472# 0.006462f
C18504 _176_ FILLER_0_15_59/a_484_472# 0.007596f
C18505 net81 _094_ 0.004737f
C18506 _077_ FILLER_0_9_72/a_36_472# 0.006408f
C18507 net31 _105_ 0.054065f
C18508 _427_/a_2248_156# vss 0.018484f
C18509 _427_/a_2665_112# vdd 0.033395f
C18510 result[1] net64 0.048458f
C18511 result[4] _418_/a_36_151# 0.005556f
C18512 net70 FILLER_0_17_104/a_1020_375# 0.001894f
C18513 _050_ _140_ 0.001f
C18514 _102_ _006_ 0.006115f
C18515 output44/a_224_472# FILLER_0_19_28/a_36_472# 0.023414f
C18516 _077_ _078_ 0.069858f
C18517 FILLER_0_8_24/a_36_472# _054_ 0.007348f
C18518 _136_ _333_/a_36_160# 0.00842f
C18519 _322_/a_848_380# _129_ 0.048486f
C18520 _429_/a_36_151# FILLER_0_13_206/a_36_472# 0.059367f
C18521 _320_/a_36_472# net21 0.025762f
C18522 FILLER_0_7_72/a_1916_375# _028_ 0.003862f
C18523 _002_ FILLER_0_3_172/a_1828_472# 0.016749f
C18524 _429_/a_2665_112# net64 0.013014f
C18525 net20 fanout63/a_36_160# 0.084165f
C18526 FILLER_0_7_72/a_1828_472# net50 0.094122f
C18527 net5 net18 0.015361f
C18528 net38 _444_/a_448_472# 0.031117f
C18529 FILLER_0_14_50/a_124_375# cal_count\[3\] 0.002524f
C18530 FILLER_0_8_37/a_124_375# _054_ 0.014206f
C18531 net63 vdd 1.002883f
C18532 _076_ _223_/a_36_160# 0.001756f
C18533 _429_/a_2665_112# mask\[1\] 0.001022f
C18534 FILLER_0_7_72/a_932_472# _028_ 0.001777f
C18535 _449_/a_2248_156# _067_ 0.040648f
C18536 FILLER_0_13_212/a_1468_375# vdd -0.013698f
C18537 FILLER_0_21_142/a_36_472# _210_/a_67_603# 0.001547f
C18538 FILLER_0_13_212/a_1020_375# vss 0.041631f
C18539 net62 FILLER_0_13_212/a_124_375# 0.001597f
C18540 _378_/a_224_472# net67 0.00211f
C18541 _081_ _265_/a_916_472# 0.002264f
C18542 _012_ FILLER_0_23_44/a_124_375# 0.002474f
C18543 _106_ _294_/a_224_472# 0.001038f
C18544 _436_/a_796_472# vdd 0.005009f
C18545 net52 _453_/a_2665_112# 0.073881f
C18546 trimb[4] FILLER_0_15_2/a_124_375# 0.003305f
C18547 FILLER_0_11_142/a_484_472# cal_count\[3\] 0.014314f
C18548 _431_/a_2248_156# _137_ 0.01617f
C18549 FILLER_0_7_72/a_2276_472# _077_ 0.00475f
C18550 _447_/a_2665_112# _441_/a_36_151# 0.028591f
C18551 trim_val\[1\] FILLER_0_5_54/a_124_375# 0.001814f
C18552 _438_/a_36_151# _437_/a_36_151# 0.002668f
C18553 vss _433_/a_448_472# 0.005349f
C18554 _058_ vdd 0.511536f
C18555 _430_/a_36_151# FILLER_0_17_200/a_572_375# 0.059049f
C18556 _118_ _121_ 0.02882f
C18557 output32/a_224_472# output34/a_224_472# 0.001691f
C18558 net66 _440_/a_36_151# 0.041433f
C18559 FILLER_0_7_104/a_1468_375# _152_ 0.009263f
C18560 net20 FILLER_0_1_212/a_124_375# 0.084041f
C18561 _086_ _310_/a_49_472# 0.013039f
C18562 _394_/a_1336_472# cal_count\[1\] 0.018116f
C18563 FILLER_0_5_172/a_36_472# _163_ 0.006934f
C18564 FILLER_0_12_124/a_36_472# _132_ 0.00101f
C18565 net74 FILLER_0_13_80/a_124_375# 0.012889f
C18566 _132_ FILLER_0_17_104/a_1020_375# 0.009251f
C18567 _415_/a_2560_156# net64 0.066438f
C18568 output21/a_224_472# vdd 0.028725f
C18569 ctln[2] ctln[3] 0.012289f
C18570 net57 _267_/a_1120_472# 0.002885f
C18571 _127_ _428_/a_36_151# 0.030717f
C18572 ctlp[1] _420_/a_36_151# 0.067975f
C18573 mask\[7\] FILLER_0_22_128/a_1020_375# 0.035799f
C18574 FILLER_0_5_198/a_572_375# vdd 0.005402f
C18575 _053_ FILLER_0_6_79/a_124_375# 0.003818f
C18576 output6/a_224_472# net6 0.076605f
C18577 net35 FILLER_0_22_128/a_484_472# 0.004578f
C18578 net45 net46 0.038161f
C18579 FILLER_0_5_128/a_36_472# _133_ 0.001217f
C18580 _126_ FILLER_0_10_94/a_572_375# 0.027249f
C18581 _114_ _127_ 0.006414f
C18582 vdd _278_/a_36_160# 0.016488f
C18583 net36 _451_/a_1353_112# 0.01266f
C18584 FILLER_0_12_136/a_124_375# _428_/a_2665_112# 0.029834f
C18585 _106_ net33 0.001049f
C18586 _437_/a_2665_112# FILLER_0_22_107/a_484_472# 0.007376f
C18587 _137_ _043_ 0.007284f
C18588 net68 FILLER_0_6_47/a_1916_375# 0.00799f
C18589 FILLER_0_19_125/a_124_375# _145_ 0.006777f
C18590 _430_/a_2665_112# net20 0.005397f
C18591 _415_/a_448_472# vdd 0.005273f
C18592 _136_ FILLER_0_16_154/a_36_472# 0.00615f
C18593 output39/a_224_472# _445_/a_36_151# 0.11862f
C18594 _078_ net37 0.459092f
C18595 FILLER_0_1_266/a_572_375# net18 0.080358f
C18596 FILLER_0_3_142/a_36_472# vss 0.012379f
C18597 _053_ FILLER_0_7_72/a_2724_472# 0.016187f
C18598 _114_ FILLER_0_12_136/a_1380_472# 0.003953f
C18599 ctlp[6] net54 0.00409f
C18600 vss FILLER_0_19_134/a_36_472# 0.005204f
C18601 net16 trim_mask\[1\] 0.007065f
C18602 _432_/a_1204_472# _137_ 0.006554f
C18603 net15 net67 0.109181f
C18604 _444_/a_1000_472# vdd 0.004148f
C18605 _104_ output18/a_224_472# 0.08426f
C18606 _155_ FILLER_0_7_104/a_572_375# 0.002336f
C18607 _027_ _438_/a_1000_472# 0.010911f
C18608 ctlp[1] _421_/a_1308_423# 0.002417f
C18609 _427_/a_1000_472# net23 0.003046f
C18610 _035_ _164_ 0.056332f
C18611 _431_/a_448_472# FILLER_0_17_142/a_124_375# 0.006782f
C18612 net79 vss 0.770834f
C18613 _446_/a_1308_423# net17 0.033125f
C18614 FILLER_0_7_146/a_36_472# vss 0.029149f
C18615 _065_ _447_/a_2560_156# 0.012523f
C18616 FILLER_0_4_144/a_124_375# _370_/a_848_380# 0.005599f
C18617 _316_/a_848_380# _122_ 0.002234f
C18618 _316_/a_692_472# calibrate 0.006232f
C18619 _394_/a_1336_472# FILLER_0_13_72/a_124_375# 0.001597f
C18620 _068_ _121_ 0.008802f
C18621 _093_ _103_ 0.124026f
C18622 mask\[4\] FILLER_0_18_209/a_36_472# 0.018888f
C18623 _083_ _084_ 0.016693f
C18624 _148_ mask\[7\] 0.010238f
C18625 net22 FILLER_0_18_209/a_36_472# 0.018061f
C18626 fanout54/a_36_160# FILLER_0_19_142/a_124_375# 0.005489f
C18627 FILLER_0_18_177/a_2276_472# FILLER_0_19_195/a_124_375# 0.001684f
C18628 _114_ _071_ 0.040513f
C18629 FILLER_0_4_123/a_124_375# FILLER_0_4_107/a_1468_375# 0.012001f
C18630 _269_/a_36_472# net59 0.011985f
C18631 net31 _047_ 0.029502f
C18632 _432_/a_36_151# vdd 0.173104f
C18633 output40/a_224_472# trim[2] 0.025041f
C18634 _141_ vss 0.308762f
C18635 result[6] output18/a_224_472# 0.003068f
C18636 FILLER_0_6_239/a_124_375# _123_ 0.044771f
C18637 mask\[8\] FILLER_0_22_107/a_124_375# 0.015331f
C18638 FILLER_0_20_87/a_124_375# net71 0.003629f
C18639 FILLER_0_21_28/a_484_472# net40 0.022617f
C18640 net74 _442_/a_1308_423# 0.001618f
C18641 _272_/a_36_472# _087_ 0.048282f
C18642 _214_/a_36_160# _051_ 0.207388f
C18643 FILLER_0_2_93/a_36_472# net49 0.001451f
C18644 net41 net16 2.918931f
C18645 _417_/a_36_151# result[3] 0.006379f
C18646 _417_/a_1308_423# net30 0.007538f
C18647 FILLER_0_16_89/a_1020_375# _136_ 0.019549f
C18648 _431_/a_2248_156# net56 0.013627f
C18649 net65 FILLER_0_3_172/a_3172_472# 0.001777f
C18650 FILLER_0_7_104/a_1020_375# _133_ 0.008772f
C18651 _077_ FILLER_0_6_231/a_36_472# 0.075292f
C18652 _085_ _161_ 0.008926f
C18653 state\[2\] _225_/a_36_160# 0.037565f
C18654 net81 net27 1.118985f
C18655 vss _295_/a_36_472# 0.009751f
C18656 _372_/a_170_472# _062_ 0.014919f
C18657 _131_ _062_ 0.120189f
C18658 FILLER_0_12_136/a_124_375# _126_ 0.013041f
C18659 net36 net71 0.148833f
C18660 net63 _024_ 0.001348f
C18661 net57 _074_ 0.026184f
C18662 FILLER_0_10_107/a_124_375# FILLER_0_10_94/a_572_375# 0.003228f
C18663 FILLER_0_17_200/a_484_472# FILLER_0_18_177/a_3172_472# 0.026657f
C18664 _129_ _124_ 0.010499f
C18665 net58 output8/a_224_472# 0.018549f
C18666 net20 ctlp[2] 0.254928f
C18667 output34/a_224_472# vdd 0.094191f
C18668 FILLER_0_10_78/a_1380_472# _115_ 0.051132f
C18669 net27 _060_ 0.045136f
C18670 FILLER_0_18_107/a_124_375# mask\[9\] 0.006029f
C18671 _094_ _418_/a_796_472# 0.005889f
C18672 _105_ net60 0.042726f
C18673 mask\[4\] output18/a_224_472# 0.017718f
C18674 _390_/a_36_68# _038_ 0.019355f
C18675 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_124_375# 0.016748f
C18676 net43 FILLER_0_20_15/a_484_472# 0.001534f
C18677 FILLER_0_11_124/a_124_375# _118_ 0.030768f
C18678 output44/a_224_472# FILLER_0_20_15/a_484_472# 0.0323f
C18679 output31/a_224_472# _418_/a_2665_112# 0.008243f
C18680 net15 FILLER_0_17_72/a_124_375# 0.006492f
C18681 FILLER_0_20_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001543f
C18682 _257_/a_36_472# _122_ 0.007741f
C18683 FILLER_0_15_282/a_572_375# result[3] 0.038939f
C18684 vss _416_/a_2665_112# 0.002676f
C18685 vdd _416_/a_2560_156# 0.00165f
C18686 _420_/a_36_151# FILLER_0_23_282/a_124_375# 0.059049f
C18687 _430_/a_796_472# _091_ 0.005465f
C18688 _367_/a_36_68# _153_ 0.019803f
C18689 FILLER_0_9_28/a_2812_375# net68 0.012462f
C18690 _408_/a_56_524# _095_ 0.01643f
C18691 FILLER_0_20_169/a_124_375# _140_ 0.01799f
C18692 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_124_375# 0.005439f
C18693 _142_ net53 0.001961f
C18694 _122_ FILLER_0_8_156/a_36_472# 0.047846f
C18695 FILLER_0_13_142/a_932_472# _043_ 0.011974f
C18696 mask\[2\] FILLER_0_16_154/a_1380_472# 0.017868f
C18697 _056_ _311_/a_66_473# 0.026074f
C18698 FILLER_0_16_107/a_572_375# FILLER_0_18_107/a_484_472# 0.001512f
C18699 net10 vdd 0.227004f
C18700 net50 FILLER_0_4_91/a_124_375# 0.022557f
C18701 net58 _425_/a_448_472# 0.002474f
C18702 _432_/a_448_472# mask\[3\] 0.005831f
C18703 _152_ net47 0.242864f
C18704 net58 FILLER_0_9_282/a_572_375# 0.006142f
C18705 net15 FILLER_0_15_59/a_124_375# 0.007439f
C18706 FILLER_0_0_232/a_124_375# vdd 0.012494f
C18707 _028_ FILLER_0_6_79/a_124_375# 0.015932f
C18708 _392_/a_244_472# cal_count\[0\] 0.003287f
C18709 net34 ctlp[1] 0.127025f
C18710 _013_ net36 0.032392f
C18711 net74 _120_ 0.027885f
C18712 fanout81/a_36_160# ctln[2] 0.003798f
C18713 _308_/a_848_380# net14 0.021982f
C18714 FILLER_0_16_73/a_572_375# _176_ 0.006454f
C18715 FILLER_0_4_197/a_36_472# net22 0.003404f
C18716 _025_ _436_/a_36_151# 0.026707f
C18717 ctlp[1] FILLER_0_24_274/a_932_472# 0.003603f
C18718 _094_ mask\[1\] 0.49634f
C18719 _428_/a_796_472# vdd 0.003502f
C18720 net69 FILLER_0_2_127/a_124_375# 0.08337f
C18721 FILLER_0_9_28/a_2276_472# _077_ 0.003256f
C18722 _214_/a_36_160# vdd 0.010812f
C18723 FILLER_0_16_107/a_572_375# _136_ 0.006445f
C18724 _028_ FILLER_0_7_72/a_2724_472# 0.001777f
C18725 cal_count\[3\] _389_/a_36_148# 0.024777f
C18726 result[8] FILLER_0_24_274/a_572_375# 0.00726f
C18727 _430_/a_448_472# _069_ 0.047845f
C18728 fanout76/a_36_160# vdd 0.108854f
C18729 FILLER_0_15_72/a_572_375# vdd 0.003801f
C18730 FILLER_0_15_72/a_124_375# vss 0.048711f
C18731 net37 FILLER_0_6_231/a_36_472# 0.002982f
C18732 fanout63/a_36_160# vss 0.008974f
C18733 _064_ _444_/a_36_151# 0.001296f
C18734 _072_ net21 0.062333f
C18735 net52 vdd 1.32956f
C18736 output33/a_224_472# ctlp[1] 0.018552f
C18737 FILLER_0_17_72/a_1828_472# _131_ 0.004882f
C18738 _091_ _143_ 0.007204f
C18739 net62 FILLER_0_14_235/a_484_472# 0.017862f
C18740 _443_/a_1308_423# vss 0.031091f
C18741 _127_ _085_ 0.00179f
C18742 net75 net10 0.073869f
C18743 net70 _136_ 0.032219f
C18744 _053_ vss 0.85895f
C18745 _413_/a_36_151# FILLER_0_4_197/a_484_472# 0.001512f
C18746 net48 _082_ 0.003853f
C18747 FILLER_0_19_55/a_124_375# _013_ 0.009611f
C18748 net75 FILLER_0_0_232/a_124_375# 0.00217f
C18749 FILLER_0_7_72/a_1468_375# _164_ 0.003223f
C18750 _072_ _070_ 2.141346f
C18751 _374_/a_36_68# _058_ 0.010442f
C18752 _077_ _251_/a_244_472# 0.002492f
C18753 net19 _420_/a_448_472# 0.05745f
C18754 _036_ FILLER_0_3_54/a_36_472# 0.002156f
C18755 _414_/a_2560_156# vss 0.001078f
C18756 _412_/a_2665_112# net18 0.001321f
C18757 net2 _425_/a_36_151# 0.012359f
C18758 FILLER_0_1_212/a_36_472# vdd 0.10765f
C18759 FILLER_0_1_212/a_124_375# vss 0.011796f
C18760 net16 _164_ 0.015161f
C18761 _132_ _318_/a_224_472# 0.001097f
C18762 _216_/a_67_603# vdd 0.030831f
C18763 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_36_472# 0.086635f
C18764 _053_ FILLER_0_6_177/a_36_472# 0.00572f
C18765 _430_/a_36_151# mask\[2\] 0.016265f
C18766 net16 FILLER_0_18_37/a_1020_375# 0.005406f
C18767 _144_ net23 0.091811f
C18768 net55 FILLER_0_21_28/a_3172_472# 0.06297f
C18769 FILLER_0_7_72/a_1468_375# FILLER_0_5_72/a_1380_472# 0.00108f
C18770 _397_/a_36_472# vss 0.003673f
C18771 FILLER_0_7_72/a_2724_472# trim_mask\[0\] 0.006975f
C18772 FILLER_0_2_177/a_484_472# vdd 0.008489f
C18773 _320_/a_1568_472# state\[1\] 0.001531f
C18774 _101_ _045_ 0.001111f
C18775 FILLER_0_8_138/a_36_472# calibrate 0.047835f
C18776 _070_ net47 0.071795f
C18777 FILLER_0_17_218/a_484_472# vss 0.035317f
C18778 _139_ FILLER_0_15_180/a_484_472# 0.004763f
C18779 FILLER_0_5_88/a_36_472# vss 0.005793f
C18780 _053_ FILLER_0_7_72/a_124_375# 0.014569f
C18781 _085_ _071_ 0.127349f
C18782 _096_ _306_/a_36_68# 0.016266f
C18783 net71 FILLER_0_22_107/a_484_472# 0.00689f
C18784 output29/a_224_472# vss 0.013148f
C18785 FILLER_0_5_206/a_36_472# net59 0.060133f
C18786 net74 _370_/a_848_380# 0.004546f
C18787 FILLER_0_21_125/a_36_472# _354_/a_49_472# 0.063744f
C18788 ctlp[1] _419_/a_448_472# 0.020153f
C18789 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_484_472# 0.013276f
C18790 _096_ _335_/a_49_472# 0.00151f
C18791 result[8] FILLER_0_23_274/a_36_472# 0.001908f
C18792 output12/a_224_472# _448_/a_36_151# 0.069748f
C18793 _387_/a_36_113# vdd 0.041853f
C18794 _016_ _131_ 0.017461f
C18795 net1 net2 0.624657f
C18796 _161_ _310_/a_49_472# 0.022411f
C18797 output28/a_224_472# FILLER_0_11_282/a_36_472# 0.008834f
C18798 net63 _337_/a_49_472# 0.001801f
C18799 _093_ FILLER_0_17_142/a_572_375# 0.009547f
C18800 net79 net4 0.386068f
C18801 _065_ _383_/a_36_472# 0.02518f
C18802 _430_/a_2665_112# vss 0.031646f
C18803 _406_/a_36_159# vdd 0.020825f
C18804 net19 _082_ 0.029316f
C18805 _434_/a_36_151# mask\[6\] 0.048644f
C18806 FILLER_0_21_286/a_36_472# vss 0.004123f
C18807 FILLER_0_21_286/a_484_472# vdd 0.007903f
C18808 FILLER_0_24_63/a_36_472# output25/a_224_472# 0.002338f
C18809 net20 _421_/a_1000_472# 0.012469f
C18810 net76 FILLER_0_5_198/a_484_472# 0.00169f
C18811 net48 _265_/a_244_68# 0.00365f
C18812 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_36_472# 0.016748f
C18813 FILLER_0_21_28/a_2276_472# _423_/a_448_472# 0.008036f
C18814 FILLER_0_18_2/a_2812_375# net40 0.018463f
C18815 _421_/a_796_472# net19 0.009462f
C18816 fanout70/a_36_113# FILLER_0_15_116/a_484_472# 0.002001f
C18817 _132_ _136_ 0.034253f
C18818 _412_/a_36_151# net2 0.003823f
C18819 result[7] FILLER_0_24_274/a_1468_375# 0.006125f
C18820 FILLER_0_15_212/a_572_375# vss 0.005835f
C18821 FILLER_0_15_212/a_1020_375# vdd -0.00211f
C18822 _093_ FILLER_0_18_76/a_124_375# 0.061549f
C18823 _050_ net14 0.001835f
C18824 _412_/a_448_472# net1 0.035155f
C18825 FILLER_0_22_86/a_36_472# _437_/a_36_151# 0.059367f
C18826 net69 _384_/a_224_472# 0.002407f
C18827 FILLER_0_5_164/a_572_375# _386_/a_848_380# 0.001121f
C18828 _319_/a_672_472# _125_ 0.002725f
C18829 _128_ _223_/a_36_160# 0.012824f
C18830 net48 _112_ 0.284235f
C18831 trim_val\[3\] _168_ 0.271475f
C18832 _303_/a_36_472# _098_ 0.021192f
C18833 _131_ FILLER_0_16_115/a_36_472# 0.008241f
C18834 net16 cal_count\[2\] 0.041089f
C18835 state\[0\] _090_ 0.003121f
C18836 _078_ _122_ 0.185069f
C18837 _083_ calibrate 0.001446f
C18838 _075_ vdd 0.190898f
C18839 FILLER_0_10_28/a_124_375# vss 0.013087f
C18840 FILLER_0_10_28/a_36_472# vdd 0.092132f
C18841 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_36_472# 0.007947f
C18842 output20/a_224_472# net78 0.001495f
C18843 _095_ _043_ 2.807456f
C18844 cal net1 0.336092f
C18845 output33/a_224_472# _204_/a_67_603# 0.00401f
C18846 mask\[4\] FILLER_0_20_177/a_1380_472# 0.001215f
C18847 _449_/a_36_151# FILLER_0_12_50/a_124_375# 0.017882f
C18848 _096_ FILLER_0_14_181/a_124_375# 0.002455f
C18849 _124_ FILLER_0_10_107/a_572_375# 0.002135f
C18850 net53 mask\[2\] 0.005907f
C18851 _114_ net23 0.029535f
C18852 net38 _445_/a_2248_156# 0.029721f
C18853 net16 FILLER_0_8_37/a_124_375# 0.010358f
C18854 _095_ _185_ 0.034457f
C18855 FILLER_0_4_197/a_1380_472# _088_ 0.017451f
C18856 _172_ vdd 0.008764f
C18857 _016_ _428_/a_2665_112# 0.050481f
C18858 net34 FILLER_0_22_177/a_36_472# 0.003953f
C18859 _420_/a_448_472# _009_ 0.061681f
C18860 _445_/a_36_151# net40 0.007227f
C18861 net74 _390_/a_244_472# 0.001317f
C18862 net80 _434_/a_796_472# 0.039593f
C18863 mask\[4\] FILLER_0_18_177/a_1020_375# 0.015941f
C18864 ctln[5] _037_ 0.19244f
C18865 fanout72/a_36_113# _449_/a_36_151# 0.032681f
C18866 _144_ net33 0.042826f
C18867 net27 net64 1.364577f
C18868 _413_/a_1308_423# net65 0.022097f
C18869 net20 _081_ 0.024512f
C18870 FILLER_0_6_90/a_572_375# _439_/a_2665_112# 0.001646f
C18871 _443_/a_36_151# net23 0.012359f
C18872 FILLER_0_5_54/a_1380_472# _440_/a_36_151# 0.001723f
C18873 FILLER_0_11_142/a_484_472# _120_ 0.007893f
C18874 FILLER_0_17_72/a_1380_472# _027_ 0.00378f
C18875 FILLER_0_17_72/a_2276_472# _150_ 0.003968f
C18876 _030_ _157_ 0.011014f
C18877 _067_ output6/a_224_472# 0.001611f
C18878 net50 _441_/a_1308_423# 0.032656f
C18879 net52 _441_/a_1000_472# 0.011506f
C18880 _175_ _095_ 0.041931f
C18881 result[4] result[9] 0.101112f
C18882 FILLER_0_8_127/a_36_472# _070_ 0.005078f
C18883 FILLER_0_4_49/a_124_375# net66 0.017584f
C18884 FILLER_0_13_212/a_1020_375# net79 0.009597f
C18885 _176_ fanout55/a_36_160# 0.070942f
C18886 ctlp[2] vss 0.131085f
C18887 FILLER_0_12_136/a_932_472# FILLER_0_13_142/a_124_375# 0.001684f
C18888 FILLER_0_16_73/a_36_472# _175_ 0.006803f
C18889 _096_ _320_/a_672_472# 0.0082f
C18890 FILLER_0_18_61/a_124_375# vdd 0.022663f
C18891 _176_ _401_/a_36_68# 0.004263f
C18892 net52 _440_/a_2560_156# 0.004924f
C18893 _028_ vss 0.410396f
C18894 _077_ _308_/a_124_24# 0.018118f
C18895 FILLER_0_12_124/a_36_472# vdd 0.040515f
C18896 fanout74/a_36_113# _443_/a_36_151# 0.032681f
C18897 net50 _439_/a_448_472# 0.020872f
C18898 net52 _439_/a_796_472# 0.003099f
C18899 FILLER_0_17_104/a_1020_375# vdd 0.012531f
C18900 ctln[3] vss 0.133697f
C18901 FILLER_0_5_54/a_36_472# FILLER_0_6_47/a_932_472# 0.026657f
C18902 FILLER_0_5_54/a_1020_375# FILLER_0_6_47/a_1828_472# 0.001597f
C18903 _425_/a_1308_423# net37 0.002601f
C18904 FILLER_0_5_164/a_36_472# vss 0.001809f
C18905 FILLER_0_5_164/a_484_472# vdd 0.005235f
C18906 net41 output40/a_224_472# 0.018977f
C18907 _110_ net36 0.002287f
C18908 _413_/a_1308_423# net59 0.018948f
C18909 net47 _450_/a_2449_156# 0.004488f
C18910 ctln[1] FILLER_0_3_221/a_124_375# 0.001391f
C18911 net15 _453_/a_2248_156# 0.044493f
C18912 _133_ _059_ 0.039848f
C18913 net20 _274_/a_1164_497# 0.002879f
C18914 _432_/a_36_151# _337_/a_49_472# 0.002462f
C18915 net69 FILLER_0_2_111/a_36_472# 0.010759f
C18916 _031_ FILLER_0_2_111/a_1020_375# 0.016661f
C18917 net52 FILLER_0_6_47/a_3172_472# 0.047876f
C18918 FILLER_0_5_109/a_572_375# _154_ 0.014669f
C18919 FILLER_0_4_49/a_124_375# _167_ 0.009437f
C18920 _178_ _402_/a_2172_497# 0.003871f
C18921 _429_/a_36_151# FILLER_0_15_212/a_124_375# 0.059049f
C18922 output20/a_224_472# ctlp[3] 0.023589f
C18923 net18 FILLER_0_13_290/a_36_472# 0.079901f
C18924 _016_ _126_ 0.051451f
C18925 FILLER_0_19_171/a_124_375# vdd -0.009473f
C18926 FILLER_0_21_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001723f
C18927 _413_/a_2248_156# net65 0.036792f
C18928 FILLER_0_7_72/a_124_375# _028_ 0.017052f
C18929 _346_/a_49_472# _145_ 0.001141f
C18930 _114_ _311_/a_1660_473# 0.003304f
C18931 mask\[3\] FILLER_0_16_241/a_36_472# 0.00209f
C18932 FILLER_0_15_235/a_124_375# vdd -0.006807f
C18933 FILLER_0_18_177/a_1916_375# net21 0.004339f
C18934 _144_ _433_/a_796_472# 0.008448f
C18935 net64 _043_ 0.004021f
C18936 FILLER_0_18_171/a_36_472# vdd 0.010704f
C18937 FILLER_0_17_200/a_36_472# vss 0.001182f
C18938 FILLER_0_14_91/a_484_472# _136_ 0.038919f
C18939 _163_ FILLER_0_5_136/a_36_472# 0.007779f
C18940 trim_mask\[0\] vss 0.014228f
C18941 mask\[1\] _043_ 0.027561f
C18942 _053_ net4 0.013559f
C18943 _101_ _285_/a_244_68# 0.001153f
C18944 result[2] _044_ 0.393081f
C18945 state\[1\] net21 0.210202f
C18946 mask\[5\] FILLER_0_18_177/a_1380_472# 0.001063f
C18947 net73 FILLER_0_15_142/a_36_472# 0.001893f
C18948 _114_ _056_ 0.034246f
C18949 _322_/a_1152_472# _118_ 0.001235f
C18950 _322_/a_124_24# _124_ 0.041337f
C18951 en net18 0.32189f
C18952 _422_/a_36_151# _010_ 0.006787f
C18953 net16 FILLER_0_17_38/a_484_472# 0.032356f
C18954 FILLER_0_14_181/a_36_472# vss 0.002955f
C18955 _233_/a_36_160# _445_/a_2248_156# 0.00136f
C18956 _221_/a_36_160# vss 0.037067f
C18957 FILLER_0_19_125/a_36_472# _145_ 0.004858f
C18958 _253_/a_1732_68# cal_itt\[1\] 0.001829f
C18959 _063_ trim_mask\[1\] 0.127216f
C18960 _425_/a_2665_112# vdd 0.012933f
C18961 net20 FILLER_0_12_220/a_932_472# 0.007397f
C18962 _100_ FILLER_0_12_236/a_484_472# 0.00195f
C18963 _413_/a_2248_156# net59 0.05485f
C18964 _165_ _033_ 0.022734f
C18965 _077_ net67 0.073924f
C18966 net70 FILLER_0_14_107/a_484_472# 0.010987f
C18967 FILLER_0_20_98/a_124_375# vdd 0.0135f
C18968 _115_ _135_ 0.004345f
C18969 FILLER_0_14_91/a_484_472# _070_ 0.001773f
C18970 mask\[5\] _146_ 0.051687f
C18971 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1468_375# 0.086635f
C18972 FILLER_0_8_263/a_124_375# calibrate 0.006928f
C18973 _070_ state\[1\] 0.032046f
C18974 _122_ FILLER_0_6_231/a_36_472# 0.015997f
C18975 _050_ _436_/a_2665_112# 0.030939f
C18976 _103_ _094_ 0.280781f
C18977 FILLER_0_16_57/a_1380_472# _131_ 0.008223f
C18978 _098_ FILLER_0_14_235/a_124_375# 0.001228f
C18979 fanout73/a_36_113# net53 0.047141f
C18980 FILLER_0_17_133/a_36_472# vss 0.006791f
C18981 _420_/a_1308_423# vss 0.001461f
C18982 _321_/a_2034_472# _120_ 0.002489f
C18983 net15 _304_/a_224_472# 0.001451f
C18984 trim_val\[4\] _443_/a_36_151# 0.009986f
C18985 cal_itt\[0\] _082_ 0.018597f
C18986 net70 _451_/a_448_472# 0.043107f
C18987 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_124_375# 0.001597f
C18988 ctln[1] FILLER_0_1_266/a_124_375# 0.002958f
C18989 net20 ctlp[1] 0.024556f
C18990 _098_ FILLER_0_15_180/a_484_472# 0.014511f
C18991 FILLER_0_10_78/a_1020_375# _176_ 0.020379f
C18992 _013_ FILLER_0_18_37/a_1468_375# 0.017213f
C18993 net19 _419_/a_1308_423# 0.056469f
C18994 ctln[4] vdd 0.210384f
C18995 _432_/a_1308_423# net80 0.030835f
C18996 net41 _063_ 0.105528f
C18997 mask\[9\] _438_/a_1000_472# 0.056239f
C18998 _093_ FILLER_0_18_139/a_1468_375# 0.004939f
C18999 ctln[5] output13/a_224_472# 0.023159f
C19000 fanout81/a_36_160# cal_itt\[1\] 0.069457f
C19001 net81 _001_ 0.012492f
C19002 output36/a_224_472# FILLER_0_15_282/a_124_375# 0.002977f
C19003 fanout59/a_36_160# net5 0.05829f
C19004 _121_ _314_/a_224_472# 0.00323f
C19005 _434_/a_1308_423# vdd 0.033494f
C19006 net15 _168_ 0.04897f
C19007 FILLER_0_3_172/a_2364_375# net22 0.013028f
C19008 FILLER_0_13_142/a_1020_375# vdd 0.018221f
C19009 FILLER_0_13_142/a_572_375# vss 0.04084f
C19010 net57 FILLER_0_8_156/a_124_375# 0.001628f
C19011 FILLER_0_17_72/a_2724_472# _438_/a_36_151# 0.002529f
C19012 _285_/a_36_472# mask\[2\] 0.002447f
C19013 FILLER_0_10_256/a_124_375# _426_/a_36_151# 0.001597f
C19014 _429_/a_448_472# _018_ 0.035489f
C19015 net34 _023_ 0.00872f
C19016 _085_ net23 0.020463f
C19017 net74 _043_ 0.65119f
C19018 _424_/a_2665_112# _423_/a_2248_156# 0.001314f
C19019 FILLER_0_14_81/a_124_375# _175_ 0.005719f
C19020 net79 _416_/a_2665_112# 0.035115f
C19021 _075_ _414_/a_2248_156# 0.044302f
C19022 FILLER_0_8_247/a_484_472# vss -0.001894f
C19023 _322_/a_1152_472# _068_ 0.001502f
C19024 FILLER_0_8_247/a_932_472# vdd 0.008645f
C19025 net81 output37/a_224_472# 0.00641f
C19026 _421_/a_1204_472# vdd 0.002198f
C19027 FILLER_0_9_28/a_2364_375# _453_/a_36_151# 0.001597f
C19028 _132_ FILLER_0_14_107/a_484_472# 0.005391f
C19029 net23 FILLER_0_22_128/a_3172_472# 0.015058f
C19030 cal_count\[3\] _408_/a_728_93# 0.040643f
C19031 _430_/a_448_472# net22 0.036303f
C19032 _034_ 0 0.304805f
C19033 _160_ 0 1.542665f
C19034 _166_ 0 0.299751f
C19035 trim[3] 0 1.777626f
C19036 output41/a_224_472# 0 2.38465f
C19037 clkc 0 0.763769f
C19038 net6 0 1.112469f
C19039 output6/a_224_472# 0 2.38465f
C19040 FILLER_0_12_196/a_36_472# 0 0.417394f
C19041 FILLER_0_12_196/a_124_375# 0 0.246306f
C19042 result[3] 0 0.50376f
C19043 net30 0 1.81422f
C19044 output30/a_224_472# 0 2.38465f
C19045 _047_ 0 0.374694f
C19046 _201_/a_67_603# 0 0.345683f
C19047 _416_/a_2560_156# 0 0.016968f
C19048 _416_/a_2665_112# 0 0.62251f
C19049 _416_/a_2248_156# 0 0.371662f
C19050 _416_/a_1204_472# 0 0.012971f
C19051 _416_/a_1000_472# 0 0.291735f
C19052 _416_/a_796_472# 0 0.023206f
C19053 _416_/a_1308_423# 0 0.279043f
C19054 _416_/a_448_472# 0 0.684413f
C19055 _416_/a_36_151# 0 1.43589f
C19056 FILLER_0_13_290/a_36_472# 0 0.417394f
C19057 FILLER_0_13_290/a_124_375# 0 0.246306f
C19058 _278_/a_36_160# 0 0.696445f
C19059 _145_ 0 0.546455f
C19060 FILLER_0_13_72/a_484_472# 0 0.345058f
C19061 FILLER_0_13_72/a_36_472# 0 0.404746f
C19062 FILLER_0_13_72/a_572_375# 0 0.232991f
C19063 FILLER_0_13_72/a_124_375# 0 0.185089f
C19064 FILLER_0_14_235/a_484_472# 0 0.345058f
C19065 FILLER_0_14_235/a_36_472# 0 0.404746f
C19066 FILLER_0_14_235/a_572_375# 0 0.232991f
C19067 FILLER_0_14_235/a_124_375# 0 0.185089f
C19068 _156_ 0 0.593796f
C19069 _107_ 0 0.391583f
C19070 _295_/a_36_472# 0 0.031137f
C19071 _022_ 0 0.387773f
C19072 _433_/a_2560_156# 0 0.016968f
C19073 _433_/a_2665_112# 0 0.62251f
C19074 _433_/a_2248_156# 0 0.371662f
C19075 _433_/a_1204_472# 0 0.012971f
C19076 _433_/a_1000_472# 0 0.291735f
C19077 _433_/a_796_472# 0 0.023206f
C19078 _433_/a_1308_423# 0 0.279043f
C19079 _433_/a_448_472# 0 0.684413f
C19080 _433_/a_36_151# 0 1.43589f
C19081 FILLER_0_5_148/a_484_472# 0 0.345058f
C19082 FILLER_0_5_148/a_36_472# 0 0.404746f
C19083 FILLER_0_5_148/a_572_375# 0 0.232991f
C19084 FILLER_0_5_148/a_124_375# 0 0.185089f
C19085 _167_ 0 0.285904f
C19086 _381_/a_36_472# 0 0.031137f
C19087 trim[2] 0 0.79181f
C19088 net40 0 1.845219f
C19089 output40/a_224_472# 0 2.38465f
C19090 cal_count\[0\] 0 0.893784f
C19091 _039_ 0 0.412301f
C19092 _450_/a_2449_156# 0 0.049992f
C19093 _450_/a_2225_156# 0 0.434082f
C19094 _450_/a_3129_107# 0 0.58406f
C19095 _450_/a_836_156# 0 0.019766f
C19096 _450_/a_1040_527# 0 0.302082f
C19097 _450_/a_1353_112# 0 0.286513f
C19098 _450_/a_448_472# 0 1.21246f
C19099 _450_/a_36_151# 0 1.31409f
C19100 rstn 0 1.86494f
C19101 FILLER_0_8_156/a_484_472# 0 0.345058f
C19102 FILLER_0_8_156/a_36_472# 0 0.404746f
C19103 FILLER_0_8_156/a_572_375# 0 0.232991f
C19104 FILLER_0_8_156/a_124_375# 0 0.185089f
C19105 FILLER_0_6_37/a_36_472# 0 0.417394f
C19106 FILLER_0_6_37/a_124_375# 0 0.246306f
C19107 FILLER_0_21_60/a_484_472# 0 0.345058f
C19108 FILLER_0_21_60/a_36_472# 0 0.404746f
C19109 FILLER_0_21_60/a_572_375# 0 0.232991f
C19110 FILLER_0_21_60/a_124_375# 0 0.185089f
C19111 FILLER_0_22_107/a_484_472# 0 0.345058f
C19112 FILLER_0_22_107/a_36_472# 0 0.404746f
C19113 FILLER_0_22_107/a_572_375# 0 0.232991f
C19114 FILLER_0_22_107/a_124_375# 0 0.185089f
C19115 FILLER_0_16_115/a_36_472# 0 0.417394f
C19116 FILLER_0_16_115/a_124_375# 0 0.246306f
C19117 FILLER_0_19_134/a_36_472# 0 0.417394f
C19118 FILLER_0_19_134/a_124_375# 0 0.246306f
C19119 FILLER_0_3_212/a_36_472# 0 0.417394f
C19120 FILLER_0_3_212/a_124_375# 0 0.246306f
C19121 FILLER_0_10_94/a_484_472# 0 0.345058f
C19122 FILLER_0_10_94/a_36_472# 0 0.404746f
C19123 FILLER_0_10_94/a_572_375# 0 0.232991f
C19124 FILLER_0_10_94/a_124_375# 0 0.185089f
C19125 FILLER_0_4_91/a_484_472# 0 0.345058f
C19126 FILLER_0_4_91/a_36_472# 0 0.404746f
C19127 FILLER_0_4_91/a_572_375# 0 0.232991f
C19128 FILLER_0_4_91/a_124_375# 0 0.185089f
C19129 net14 0 1.508711f
C19130 _202_/a_36_160# 0 0.696445f
C19131 FILLER_0_6_231/a_484_472# 0 0.345058f
C19132 FILLER_0_6_231/a_36_472# 0 0.404746f
C19133 FILLER_0_6_231/a_572_375# 0 0.232991f
C19134 FILLER_0_6_231/a_124_375# 0 0.185089f
C19135 vss 0 65.60368f
C19136 vdd 0 1.086009p
C19137 _006_ 0 0.41456f
C19138 _417_/a_2560_156# 0 0.016968f
C19139 _417_/a_2665_112# 0 0.62251f
C19140 _417_/a_2248_156# 0 0.371662f
C19141 _417_/a_1204_472# 0 0.012971f
C19142 _417_/a_1000_472# 0 0.291735f
C19143 _417_/a_796_472# 0 0.023206f
C19144 _417_/a_1308_423# 0 0.279043f
C19145 _417_/a_448_472# 0 0.684413f
C19146 _417_/a_36_151# 0 1.43589f
C19147 _146_ 0 0.35443f
C19148 mask\[6\] 0 1.246962f
C19149 _348_/a_49_472# 0 0.054843f
C19150 _365_/a_36_68# 0 0.150048f
C19151 _023_ 0 0.345812f
C19152 _434_/a_2560_156# 0 0.016968f
C19153 _434_/a_2665_112# 0 0.62251f
C19154 _434_/a_2248_156# 0 0.371662f
C19155 _434_/a_1204_472# 0 0.012971f
C19156 _434_/a_1000_472# 0 0.291735f
C19157 _434_/a_796_472# 0 0.023206f
C19158 _434_/a_1308_423# 0 0.279043f
C19159 _434_/a_448_472# 0 0.684413f
C19160 _434_/a_36_151# 0 1.43589f
C19161 FILLER_0_5_136/a_36_472# 0 0.417394f
C19162 FILLER_0_5_136/a_124_375# 0 0.246306f
C19163 FILLER_0_18_209/a_484_472# 0 0.345058f
C19164 FILLER_0_18_209/a_36_472# 0 0.404746f
C19165 FILLER_0_18_209/a_572_375# 0 0.232991f
C19166 FILLER_0_18_209/a_124_375# 0 0.185089f
C19167 FILLER_0_12_28/a_36_472# 0 0.417394f
C19168 FILLER_0_12_28/a_124_375# 0 0.246306f
C19169 _040_ 0 0.355703f
C19170 _451_/a_2449_156# 0 0.049992f
C19171 _451_/a_2225_156# 0 0.434082f
C19172 _451_/a_3129_107# 0 0.58406f
C19173 _451_/a_836_156# 0 0.019766f
C19174 _451_/a_1040_527# 0 0.302082f
C19175 _451_/a_1353_112# 0 0.286513f
C19176 _451_/a_448_472# 0 1.21246f
C19177 _451_/a_36_151# 0 1.31409f
C19178 FILLER_0_6_47/a_3172_472# 0 0.345058f
C19179 FILLER_0_6_47/a_2724_472# 0 0.33241f
C19180 FILLER_0_6_47/a_2276_472# 0 0.33241f
C19181 FILLER_0_6_47/a_1828_472# 0 0.33241f
C19182 FILLER_0_6_47/a_1380_472# 0 0.33241f
C19183 FILLER_0_6_47/a_932_472# 0 0.33241f
C19184 FILLER_0_6_47/a_484_472# 0 0.33241f
C19185 FILLER_0_6_47/a_36_472# 0 0.404746f
C19186 FILLER_0_6_47/a_3260_375# 0 0.233093f
C19187 FILLER_0_6_47/a_2812_375# 0 0.17167f
C19188 FILLER_0_6_47/a_2364_375# 0 0.17167f
C19189 FILLER_0_6_47/a_1916_375# 0 0.17167f
C19190 FILLER_0_6_47/a_1468_375# 0 0.17167f
C19191 FILLER_0_6_47/a_1020_375# 0 0.17167f
C19192 FILLER_0_6_47/a_572_375# 0 0.17167f
C19193 FILLER_0_6_47/a_124_375# 0 0.185915f
C19194 FILLER_0_21_150/a_36_472# 0 0.417394f
C19195 FILLER_0_21_150/a_124_375# 0 0.246306f
C19196 FILLER_0_15_180/a_484_472# 0 0.345058f
C19197 FILLER_0_15_180/a_36_472# 0 0.404746f
C19198 FILLER_0_15_180/a_572_375# 0 0.232991f
C19199 FILLER_0_15_180/a_124_375# 0 0.185089f
C19200 FILLER_0_22_128/a_3172_472# 0 0.345058f
C19201 FILLER_0_22_128/a_2724_472# 0 0.33241f
C19202 FILLER_0_22_128/a_2276_472# 0 0.33241f
C19203 FILLER_0_22_128/a_1828_472# 0 0.33241f
C19204 FILLER_0_22_128/a_1380_472# 0 0.33241f
C19205 FILLER_0_22_128/a_932_472# 0 0.33241f
C19206 FILLER_0_22_128/a_484_472# 0 0.33241f
C19207 FILLER_0_22_128/a_36_472# 0 0.404746f
C19208 FILLER_0_22_128/a_3260_375# 0 0.233093f
C19209 FILLER_0_22_128/a_2812_375# 0 0.17167f
C19210 FILLER_0_22_128/a_2364_375# 0 0.17167f
C19211 FILLER_0_22_128/a_1916_375# 0 0.17167f
C19212 FILLER_0_22_128/a_1468_375# 0 0.17167f
C19213 FILLER_0_22_128/a_1020_375# 0 0.17167f
C19214 FILLER_0_22_128/a_572_375# 0 0.17167f
C19215 FILLER_0_22_128/a_124_375# 0 0.185915f
C19216 FILLER_0_19_111/a_484_472# 0 0.345058f
C19217 FILLER_0_19_111/a_36_472# 0 0.404746f
C19218 FILLER_0_19_111/a_572_375# 0 0.232991f
C19219 FILLER_0_19_111/a_124_375# 0 0.185089f
C19220 FILLER_0_19_155/a_484_472# 0 0.345058f
C19221 FILLER_0_19_155/a_36_472# 0 0.404746f
C19222 FILLER_0_19_155/a_572_375# 0 0.232991f
C19223 FILLER_0_19_155/a_124_375# 0 0.185089f
C19224 net11 0 1.328455f
C19225 net21 0 1.922829f
C19226 _007_ 0 0.309495f
C19227 net77 0 1.39077f
C19228 _418_/a_2560_156# 0 0.016968f
C19229 _418_/a_2665_112# 0 0.62251f
C19230 _418_/a_2248_156# 0 0.371662f
C19231 _418_/a_1204_472# 0 0.012971f
C19232 _418_/a_1000_472# 0 0.291735f
C19233 _418_/a_796_472# 0 0.023206f
C19234 _418_/a_1308_423# 0 0.279043f
C19235 _418_/a_448_472# 0 0.684413f
C19236 _418_/a_36_151# 0 1.43589f
C19237 _220_/a_67_603# 0 0.345683f
C19238 FILLER_0_9_282/a_484_472# 0 0.345058f
C19239 FILLER_0_9_282/a_36_472# 0 0.404746f
C19240 FILLER_0_9_282/a_572_375# 0 0.232991f
C19241 FILLER_0_9_282/a_124_375# 0 0.185089f
C19242 FILLER_0_18_37/a_1380_472# 0 0.345058f
C19243 FILLER_0_18_37/a_932_472# 0 0.33241f
C19244 FILLER_0_18_37/a_484_472# 0 0.33241f
C19245 FILLER_0_18_37/a_36_472# 0 0.404746f
C19246 FILLER_0_18_37/a_1468_375# 0 0.233029f
C19247 FILLER_0_18_37/a_1020_375# 0 0.171606f
C19248 FILLER_0_18_37/a_572_375# 0 0.171606f
C19249 FILLER_0_18_37/a_124_375# 0 0.185399f
C19250 FILLER_0_2_127/a_36_472# 0 0.417394f
C19251 FILLER_0_2_127/a_124_375# 0 0.246306f
C19252 _157_ 0 0.531763f
C19253 _435_/a_2560_156# 0 0.016968f
C19254 _435_/a_2665_112# 0 0.62251f
C19255 _435_/a_2248_156# 0 0.371662f
C19256 _435_/a_1204_472# 0 0.012971f
C19257 _435_/a_1000_472# 0 0.291735f
C19258 _435_/a_796_472# 0 0.023206f
C19259 _435_/a_1308_423# 0 0.279043f
C19260 _435_/a_448_472# 0 0.684413f
C19261 _435_/a_36_151# 0 1.43589f
C19262 _108_ 0 0.411979f
C19263 _297_/a_36_472# 0 0.031137f
C19264 trim_mask\[3\] 0 1.081535f
C19265 _164_ 0 1.3268f
C19266 _383_/a_36_472# 0 0.031137f
C19267 _041_ 0 0.299289f
C19268 _452_/a_2449_156# 0 0.049992f
C19269 _452_/a_2225_156# 0 0.434082f
C19270 _452_/a_3129_107# 0 0.58406f
C19271 _452_/a_836_156# 0 0.019766f
C19272 _452_/a_1040_527# 0 0.302082f
C19273 _452_/a_1353_112# 0 0.286513f
C19274 _452_/a_448_472# 0 1.21246f
C19275 _452_/a_36_151# 0 1.31409f
C19276 FILLER_0_6_79/a_36_472# 0 0.417394f
C19277 FILLER_0_6_79/a_124_375# 0 0.246306f
C19278 net59 0 5.044369f
C19279 FILLER_0_15_59/a_484_472# 0 0.345058f
C19280 FILLER_0_15_59/a_36_472# 0 0.404746f
C19281 FILLER_0_15_59/a_572_375# 0 0.232991f
C19282 FILLER_0_15_59/a_124_375# 0 0.185089f
C19283 FILLER_0_3_221/a_1380_472# 0 0.345058f
C19284 FILLER_0_3_221/a_932_472# 0 0.33241f
C19285 FILLER_0_3_221/a_484_472# 0 0.33241f
C19286 FILLER_0_3_221/a_36_472# 0 0.404746f
C19287 FILLER_0_3_221/a_1468_375# 0 0.233029f
C19288 FILLER_0_3_221/a_1020_375# 0 0.171606f
C19289 FILLER_0_3_221/a_572_375# 0 0.171606f
C19290 FILLER_0_3_221/a_124_375# 0 0.185399f
C19291 FILLER_0_19_187/a_484_472# 0 0.345058f
C19292 FILLER_0_19_187/a_36_472# 0 0.404746f
C19293 FILLER_0_19_187/a_572_375# 0 0.232991f
C19294 FILLER_0_19_187/a_124_375# 0 0.185089f
C19295 FILLER_0_20_15/a_1380_472# 0 0.345058f
C19296 FILLER_0_20_15/a_932_472# 0 0.33241f
C19297 FILLER_0_20_15/a_484_472# 0 0.33241f
C19298 FILLER_0_20_15/a_36_472# 0 0.404746f
C19299 FILLER_0_20_15/a_1468_375# 0 0.233029f
C19300 FILLER_0_20_15/a_1020_375# 0 0.171606f
C19301 FILLER_0_20_15/a_572_375# 0 0.171606f
C19302 FILLER_0_20_15/a_124_375# 0 0.185399f
C19303 _204_/a_67_603# 0 0.345683f
C19304 _419_/a_2560_156# 0 0.016968f
C19305 _419_/a_2665_112# 0 0.62251f
C19306 _419_/a_2248_156# 0 0.371662f
C19307 _419_/a_1204_472# 0 0.012971f
C19308 _419_/a_1000_472# 0 0.291735f
C19309 _419_/a_796_472# 0 0.023206f
C19310 _419_/a_1308_423# 0 0.279043f
C19311 _419_/a_448_472# 0 0.684413f
C19312 _419_/a_36_151# 0 1.43589f
C19313 _054_ 0 0.522819f
C19314 _221_/a_36_160# 0 0.386641f
C19315 FILLER_0_9_270/a_484_472# 0 0.345058f
C19316 FILLER_0_9_270/a_36_472# 0 0.404746f
C19317 FILLER_0_9_270/a_572_375# 0 0.232991f
C19318 FILLER_0_9_270/a_124_375# 0 0.185089f
C19319 FILLER_0_1_192/a_36_472# 0 0.417394f
C19320 FILLER_0_1_192/a_124_375# 0 0.246306f
C19321 FILLER_0_13_80/a_36_472# 0 0.417394f
C19322 FILLER_0_13_80/a_124_375# 0 0.246306f
C19323 _153_ 0 1.165862f
C19324 _154_ 0 1.167112f
C19325 _367_/a_36_68# 0 0.150048f
C19326 _436_/a_2560_156# 0 0.016968f
C19327 _436_/a_2665_112# 0 0.62251f
C19328 _436_/a_2248_156# 0 0.371662f
C19329 _436_/a_1204_472# 0 0.012971f
C19330 _436_/a_1000_472# 0 0.291735f
C19331 _436_/a_796_472# 0 0.023206f
C19332 _436_/a_1308_423# 0 0.279043f
C19333 _436_/a_448_472# 0 0.684413f
C19334 _436_/a_36_151# 0 1.43589f
C19335 FILLER_0_10_107/a_484_472# 0 0.345058f
C19336 FILLER_0_10_107/a_36_472# 0 0.404746f
C19337 FILLER_0_10_107/a_572_375# 0 0.232991f
C19338 FILLER_0_10_107/a_124_375# 0 0.185089f
C19339 _168_ 0 0.336537f
C19340 net51 0 2.105066f
C19341 _042_ 0 0.323587f
C19342 _453_/a_2560_156# 0 0.016968f
C19343 _453_/a_2665_112# 0 0.62251f
C19344 _453_/a_2248_156# 0 0.371662f
C19345 _453_/a_1204_472# 0 0.012971f
C19346 _453_/a_1000_472# 0 0.291735f
C19347 _453_/a_796_472# 0 0.023206f
C19348 _453_/a_1308_423# 0 0.279043f
C19349 _453_/a_448_472# 0 0.684413f
C19350 _453_/a_36_151# 0 1.43589f
C19351 FILLER_0_19_142/a_36_472# 0 0.417394f
C19352 FILLER_0_19_142/a_124_375# 0 0.246306f
C19353 _048_ 0 0.358805f
C19354 _205_/a_36_160# 0 0.696445f
C19355 net43 0 1.236377f
C19356 FILLER_0_3_78/a_484_472# 0 0.345058f
C19357 FILLER_0_3_78/a_36_472# 0 0.404746f
C19358 FILLER_0_3_78/a_572_375# 0 0.232991f
C19359 FILLER_0_3_78/a_124_375# 0 0.185089f
C19360 _437_/a_2560_156# 0 0.016968f
C19361 _437_/a_2665_112# 0 0.62251f
C19362 _437_/a_2248_156# 0 0.371662f
C19363 _437_/a_1204_472# 0 0.012971f
C19364 _437_/a_1000_472# 0 0.291735f
C19365 _437_/a_796_472# 0 0.023206f
C19366 _437_/a_1308_423# 0 0.279043f
C19367 _437_/a_448_472# 0 0.684413f
C19368 _437_/a_36_151# 0 1.43589f
C19369 _109_ 0 0.319326f
C19370 _299_/a_36_472# 0 0.031137f
C19371 net37 0 1.529713f
C19372 _385_/a_36_68# 0 0.112263f
C19373 FILLER_0_0_266/a_36_472# 0 0.417394f
C19374 FILLER_0_0_266/a_124_375# 0 0.246306f
C19375 net12 0 1.263595f
C19376 net22 0 2.108509f
C19377 FILLER_0_9_290/a_36_472# 0 0.417394f
C19378 FILLER_0_9_290/a_124_375# 0 0.246306f
C19379 _223_/a_36_160# 0 0.696445f
C19380 FILLER_0_14_263/a_36_472# 0 0.417394f
C19381 FILLER_0_14_263/a_124_375# 0 0.246306f
C19382 _158_ 0 0.309522f
C19383 _369_/a_36_68# 0 0.150048f
C19384 net71 0 1.420869f
C19385 _438_/a_2560_156# 0 0.016968f
C19386 _438_/a_2665_112# 0 0.62251f
C19387 _438_/a_2248_156# 0 0.371662f
C19388 _438_/a_1204_472# 0 0.012971f
C19389 _438_/a_1000_472# 0 0.291735f
C19390 _438_/a_796_472# 0 0.023206f
C19391 _438_/a_1308_423# 0 0.279043f
C19392 _438_/a_448_472# 0 0.684413f
C19393 _438_/a_36_151# 0 1.43589f
C19394 FILLER_0_23_274/a_36_472# 0 0.417394f
C19395 FILLER_0_23_274/a_124_375# 0 0.246306f
C19396 FILLER_0_17_282/a_36_472# 0 0.417394f
C19397 FILLER_0_17_282/a_124_375# 0 0.246306f
C19398 FILLER_0_5_198/a_484_472# 0 0.345058f
C19399 FILLER_0_5_198/a_36_472# 0 0.404746f
C19400 FILLER_0_5_198/a_572_375# 0 0.232991f
C19401 FILLER_0_5_198/a_124_375# 0 0.185089f
C19402 _163_ 0 1.03762f
C19403 _169_ 0 0.245383f
C19404 _386_/a_848_380# 0 0.40208f
C19405 _386_/a_124_24# 0 0.591898f
C19406 FILLER_0_20_2/a_484_472# 0 0.345058f
C19407 FILLER_0_20_2/a_36_472# 0 0.404746f
C19408 FILLER_0_20_2/a_572_375# 0 0.232991f
C19409 FILLER_0_20_2/a_124_375# 0 0.185089f
C19410 FILLER_0_16_154/a_1380_472# 0 0.345058f
C19411 FILLER_0_16_154/a_932_472# 0 0.33241f
C19412 FILLER_0_16_154/a_484_472# 0 0.33241f
C19413 FILLER_0_16_154/a_36_472# 0 0.404746f
C19414 FILLER_0_16_154/a_1468_375# 0 0.233029f
C19415 FILLER_0_16_154/a_1020_375# 0 0.171606f
C19416 FILLER_0_16_154/a_572_375# 0 0.171606f
C19417 FILLER_0_16_154/a_124_375# 0 0.185399f
C19418 FILLER_0_0_232/a_36_472# 0 0.417394f
C19419 FILLER_0_0_232/a_124_375# 0 0.246306f
C19420 FILLER_0_19_195/a_36_472# 0 0.417394f
C19421 FILLER_0_19_195/a_124_375# 0 0.246306f
C19422 _049_ 0 0.329957f
C19423 net33 0 1.934915f
C19424 _207_/a_67_603# 0 0.345683f
C19425 FILLER_0_3_54/a_36_472# 0 0.417394f
C19426 FILLER_0_3_54/a_124_375# 0 0.246306f
C19427 FILLER_0_2_101/a_36_472# 0 0.417394f
C19428 FILLER_0_2_101/a_124_375# 0 0.246306f
C19429 trim_mask\[0\] 0 0.605753f
C19430 _439_/a_2560_156# 0 0.016968f
C19431 _439_/a_2665_112# 0 0.62251f
C19432 _439_/a_2248_156# 0 0.371662f
C19433 _439_/a_1204_472# 0 0.012971f
C19434 _439_/a_1000_472# 0 0.291735f
C19435 _439_/a_796_472# 0 0.023206f
C19436 _439_/a_1308_423# 0 0.279043f
C19437 _439_/a_448_472# 0 0.684413f
C19438 _439_/a_36_151# 0 1.43589f
C19439 _066_ 0 0.333041f
C19440 FILLER_0_23_44/a_1380_472# 0 0.345058f
C19441 FILLER_0_23_44/a_932_472# 0 0.33241f
C19442 FILLER_0_23_44/a_484_472# 0 0.33241f
C19443 FILLER_0_23_44/a_36_472# 0 0.404746f
C19444 FILLER_0_23_44/a_1468_375# 0 0.233029f
C19445 FILLER_0_23_44/a_1020_375# 0 0.171606f
C19446 FILLER_0_23_44/a_572_375# 0 0.171606f
C19447 FILLER_0_23_44/a_124_375# 0 0.185399f
C19448 FILLER_0_23_88/a_36_472# 0 0.417394f
C19449 FILLER_0_23_88/a_124_375# 0 0.246306f
C19450 FILLER_0_5_164/a_484_472# 0 0.345058f
C19451 FILLER_0_5_164/a_36_472# 0 0.404746f
C19452 FILLER_0_5_164/a_572_375# 0 0.232991f
C19453 FILLER_0_5_164/a_124_375# 0 0.185089f
C19454 _060_ 0 2.485177f
C19455 _113_ 0 2.833205f
C19456 _090_ 0 2.629271f
C19457 _310_/a_49_472# 0 0.098072f
C19458 _037_ 0 0.467089f
C19459 _170_ 0 0.413995f
C19460 _387_/a_36_113# 0 0.418095f
C19461 _208_/a_36_160# 0 0.696445f
C19462 FILLER_0_18_76/a_484_472# 0 0.345058f
C19463 FILLER_0_18_76/a_36_472# 0 0.404746f
C19464 FILLER_0_18_76/a_572_375# 0 0.232991f
C19465 FILLER_0_18_76/a_124_375# 0 0.185089f
C19466 _225_/a_36_160# 0 0.386641f
C19467 FILLER_0_2_177/a_484_472# 0 0.345058f
C19468 FILLER_0_2_177/a_36_472# 0 0.404746f
C19469 FILLER_0_2_177/a_572_375# 0 0.232991f
C19470 FILLER_0_2_177/a_124_375# 0 0.185089f
C19471 FILLER_0_2_111/a_1380_472# 0 0.345058f
C19472 FILLER_0_2_111/a_932_472# 0 0.33241f
C19473 FILLER_0_2_111/a_484_472# 0 0.33241f
C19474 FILLER_0_2_111/a_36_472# 0 0.404746f
C19475 FILLER_0_2_111/a_1468_375# 0 0.233029f
C19476 FILLER_0_2_111/a_1020_375# 0 0.171606f
C19477 FILLER_0_2_111/a_572_375# 0 0.171606f
C19478 FILLER_0_2_111/a_124_375# 0 0.185399f
C19479 FILLER_0_15_228/a_36_472# 0 0.417394f
C19480 FILLER_0_15_228/a_124_375# 0 0.246306f
C19481 net47 0 2.314376f
C19482 _242_/a_36_160# 0 0.696445f
C19483 _117_ 0 1.266251f
C19484 _311_/a_66_473# 0 0.11665f
C19485 _043_ 0 0.487279f
C19486 _190_/a_36_160# 0 0.696445f
C19487 FILLER_0_9_105/a_484_472# 0 0.345058f
C19488 FILLER_0_9_105/a_36_472# 0 0.404746f
C19489 FILLER_0_9_105/a_572_375# 0 0.232991f
C19490 FILLER_0_9_105/a_124_375# 0 0.185089f
C19491 FILLER_0_13_100/a_36_472# 0 0.417394f
C19492 FILLER_0_13_100/a_124_375# 0 0.246306f
C19493 FILLER_0_22_177/a_1380_472# 0 0.345058f
C19494 FILLER_0_22_177/a_932_472# 0 0.33241f
C19495 FILLER_0_22_177/a_484_472# 0 0.33241f
C19496 FILLER_0_22_177/a_36_472# 0 0.404746f
C19497 FILLER_0_22_177/a_1468_375# 0 0.233029f
C19498 FILLER_0_22_177/a_1020_375# 0 0.171606f
C19499 FILLER_0_22_177/a_572_375# 0 0.171606f
C19500 FILLER_0_22_177/a_124_375# 0 0.185399f
C19501 FILLER_0_15_2/a_484_472# 0 0.345058f
C19502 FILLER_0_15_2/a_36_472# 0 0.404746f
C19503 FILLER_0_15_2/a_572_375# 0 0.232991f
C19504 FILLER_0_15_2/a_124_375# 0 0.185089f
C19505 FILLER_0_15_10/a_36_472# 0 0.417394f
C19506 FILLER_0_15_10/a_124_375# 0 0.246306f
C19507 FILLER_0_19_171/a_1380_472# 0 0.345058f
C19508 FILLER_0_19_171/a_932_472# 0 0.33241f
C19509 FILLER_0_19_171/a_484_472# 0 0.33241f
C19510 FILLER_0_19_171/a_36_472# 0 0.404746f
C19511 FILLER_0_19_171/a_1468_375# 0 0.233029f
C19512 FILLER_0_19_171/a_1020_375# 0 0.171606f
C19513 FILLER_0_19_171/a_572_375# 0 0.171606f
C19514 FILLER_0_19_171/a_124_375# 0 0.185399f
C19515 net13 0 1.176306f
C19516 net23 0 2.091399f
C19517 FILLER_0_20_87/a_36_472# 0 0.417394f
C19518 FILLER_0_20_87/a_124_375# 0 0.246306f
C19519 FILLER_0_20_98/a_36_472# 0 0.417394f
C19520 FILLER_0_20_98/a_124_375# 0 0.246306f
C19521 _055_ 0 1.782885f
C19522 FILLER_0_18_53/a_484_472# 0 0.345058f
C19523 FILLER_0_18_53/a_36_472# 0 0.404746f
C19524 FILLER_0_18_53/a_572_375# 0 0.232991f
C19525 FILLER_0_18_53/a_124_375# 0 0.185089f
C19526 FILLER_0_2_165/a_36_472# 0 0.417394f
C19527 FILLER_0_2_165/a_124_375# 0 0.246306f
C19528 FILLER_0_15_205/a_36_472# 0 0.417394f
C19529 FILLER_0_15_205/a_124_375# 0 0.246306f
C19530 FILLER_0_23_282/a_484_472# 0 0.345058f
C19531 FILLER_0_23_282/a_36_472# 0 0.404746f
C19532 FILLER_0_23_282/a_572_375# 0 0.232991f
C19533 FILLER_0_23_282/a_124_375# 0 0.185089f
C19534 net42 0 1.067446f
C19535 net17 0 2.210219f
C19536 _172_ 0 0.265782f
C19537 _171_ 0 0.300355f
C19538 _389_/a_36_148# 0 0.388358f
C19539 _080_ 0 0.328202f
C19540 _260_/a_36_68# 0 0.112263f
C19541 FILLER_0_0_96/a_36_472# 0 0.417394f
C19542 FILLER_0_0_96/a_124_375# 0 0.246306f
C19543 FILLER_0_9_72/a_1380_472# 0 0.345058f
C19544 FILLER_0_9_72/a_932_472# 0 0.33241f
C19545 FILLER_0_9_72/a_484_472# 0 0.33241f
C19546 FILLER_0_9_72/a_36_472# 0 0.404746f
C19547 FILLER_0_9_72/a_1468_375# 0 0.233029f
C19548 FILLER_0_9_72/a_1020_375# 0 0.171606f
C19549 FILLER_0_9_72/a_572_375# 0 0.171606f
C19550 FILLER_0_9_72/a_124_375# 0 0.185399f
C19551 FILLER_0_20_31/a_36_472# 0 0.417394f
C19552 FILLER_0_20_31/a_124_375# 0 0.246306f
C19553 _227_/a_36_160# 0 0.386641f
C19554 _120_ 0 1.533088f
C19555 _313_/a_67_603# 0 0.345683f
C19556 FILLER_0_5_172/a_36_472# 0 0.417394f
C19557 FILLER_0_5_172/a_124_375# 0 0.246306f
C19558 FILLER_0_12_20/a_484_472# 0 0.345058f
C19559 FILLER_0_12_20/a_36_472# 0 0.404746f
C19560 FILLER_0_12_20/a_572_375# 0 0.232991f
C19561 FILLER_0_12_20/a_124_375# 0 0.185089f
C19562 _134_ 0 0.365972f
C19563 _062_ 0 1.717773f
C19564 _059_ 0 1.686761f
C19565 _261_/a_36_160# 0 0.386641f
C19566 _044_ 0 0.388801f
C19567 mask\[1\] 0 1.295078f
C19568 _192_/a_67_603# 0 0.345683f
C19569 FILLER_0_13_142/a_1380_472# 0 0.345058f
C19570 FILLER_0_13_142/a_932_472# 0 0.33241f
C19571 FILLER_0_13_142/a_484_472# 0 0.33241f
C19572 FILLER_0_13_142/a_36_472# 0 0.404746f
C19573 FILLER_0_13_142/a_1468_375# 0 0.233029f
C19574 FILLER_0_13_142/a_1020_375# 0 0.171606f
C19575 FILLER_0_13_142/a_572_375# 0 0.171606f
C19576 FILLER_0_13_142/a_124_375# 0 0.185399f
C19577 FILLER_0_9_60/a_484_472# 0 0.345058f
C19578 FILLER_0_9_60/a_36_472# 0 0.404746f
C19579 FILLER_0_9_60/a_572_375# 0 0.232991f
C19580 FILLER_0_9_60/a_124_375# 0 0.185089f
C19581 FILLER_0_7_233/a_36_472# 0 0.417394f
C19582 FILLER_0_7_233/a_124_375# 0 0.246306f
C19583 _228_/a_36_68# 0 0.69549f
C19584 FILLER_0_21_206/a_36_472# 0 0.417394f
C19585 FILLER_0_21_206/a_124_375# 0 0.246306f
C19586 _067_ 0 0.851951f
C19587 _135_ 0 0.339478f
C19588 _193_/a_36_160# 0 0.696445f
C19589 _180_ 0 0.390598f
C19590 cal_count\[1\] 0 1.568289f
C19591 FILLER_0_4_213/a_484_472# 0 0.345058f
C19592 FILLER_0_4_213/a_36_472# 0 0.404746f
C19593 FILLER_0_4_213/a_572_375# 0 0.232991f
C19594 FILLER_0_4_213/a_124_375# 0 0.185089f
C19595 FILLER_0_11_282/a_36_472# 0 0.417394f
C19596 FILLER_0_11_282/a_124_375# 0 0.246306f
C19597 FILLER_0_18_61/a_36_472# 0 0.417394f
C19598 FILLER_0_18_61/a_124_375# 0 0.246306f
C19599 FILLER_0_15_235/a_484_472# 0 0.345058f
C19600 FILLER_0_15_235/a_36_472# 0 0.404746f
C19601 FILLER_0_15_235/a_572_375# 0 0.232991f
C19602 FILLER_0_15_235/a_124_375# 0 0.185089f
C19603 FILLER_0_23_290/a_36_472# 0 0.417394f
C19604 FILLER_0_23_290/a_124_375# 0 0.246306f
C19605 _121_ 0 0.532847f
C19606 _315_/a_36_68# 0 0.052951f
C19607 _246_/a_36_68# 0 0.69549f
C19608 FILLER_0_5_181/a_36_472# 0 0.417394f
C19609 FILLER_0_5_181/a_124_375# 0 0.246306f
C19610 _082_ 0 0.619901f
C19611 net8 0 1.163723f
C19612 net18 0 2.032159f
C19613 _332_/a_36_472# 0 0.031137f
C19614 _179_ 0 0.336984f
C19615 _401_/a_36_68# 0 0.112263f
C19616 FILLER_0_14_107/a_1380_472# 0 0.345058f
C19617 FILLER_0_14_107/a_932_472# 0 0.33241f
C19618 FILLER_0_14_107/a_484_472# 0 0.33241f
C19619 FILLER_0_14_107/a_36_472# 0 0.404746f
C19620 FILLER_0_14_107/a_1468_375# 0 0.233029f
C19621 FILLER_0_14_107/a_1020_375# 0 0.171606f
C19622 FILLER_0_14_107/a_572_375# 0 0.171606f
C19623 FILLER_0_14_107/a_124_375# 0 0.185399f
C19624 _097_ 0 0.592554f
C19625 FILLER_0_1_204/a_36_472# 0 0.417394f
C19626 FILLER_0_1_204/a_124_375# 0 0.246306f
C19627 FILLER_0_15_72/a_484_472# 0 0.345058f
C19628 FILLER_0_15_72/a_36_472# 0 0.404746f
C19629 FILLER_0_15_72/a_572_375# 0 0.232991f
C19630 FILLER_0_15_72/a_124_375# 0 0.185089f
C19631 FILLER_0_17_104/a_1380_472# 0 0.345058f
C19632 FILLER_0_17_104/a_932_472# 0 0.33241f
C19633 FILLER_0_17_104/a_484_472# 0 0.33241f
C19634 FILLER_0_17_104/a_36_472# 0 0.404746f
C19635 FILLER_0_17_104/a_1468_375# 0 0.233029f
C19636 FILLER_0_17_104/a_1020_375# 0 0.171606f
C19637 FILLER_0_17_104/a_572_375# 0 0.171606f
C19638 FILLER_0_17_104/a_124_375# 0 0.185399f
C19639 FILLER_0_8_37/a_484_472# 0 0.345058f
C19640 FILLER_0_8_37/a_36_472# 0 0.404746f
C19641 FILLER_0_8_37/a_572_375# 0 0.232991f
C19642 FILLER_0_8_37/a_124_375# 0 0.185089f
C19643 FILLER_0_15_212/a_1380_472# 0 0.345058f
C19644 FILLER_0_15_212/a_932_472# 0 0.33241f
C19645 FILLER_0_15_212/a_484_472# 0 0.33241f
C19646 FILLER_0_15_212/a_36_472# 0 0.404746f
C19647 FILLER_0_15_212/a_1468_375# 0 0.233029f
C19648 FILLER_0_15_212/a_1020_375# 0 0.171606f
C19649 FILLER_0_15_212/a_572_375# 0 0.171606f
C19650 FILLER_0_15_212/a_124_375# 0 0.185399f
C19651 FILLER_0_23_60/a_36_472# 0 0.417394f
C19652 FILLER_0_23_60/a_124_375# 0 0.246306f
C19653 _123_ 0 0.344874f
C19654 _122_ 0 0.600118f
C19655 calibrate 0 1.343796f
C19656 _316_/a_848_380# 0 0.40208f
C19657 _316_/a_124_24# 0 0.591898f
C19658 _247_/a_36_160# 0 0.696445f
C19659 FILLER_0_12_50/a_36_472# 0 0.417394f
C19660 FILLER_0_12_50/a_124_375# 0 0.246306f
C19661 _084_ 0 0.296163f
C19662 cal_itt\[0\] 0 1.831055f
C19663 cal_itt\[1\] 0 1.705665f
C19664 FILLER_0_11_109/a_36_472# 0 0.417394f
C19665 FILLER_0_11_109/a_124_375# 0 0.246306f
C19666 _182_ 0 0.34197f
C19667 _402_/a_1948_68# 0 0.022025f
C19668 _402_/a_718_527# 0 0.001795f
C19669 _402_/a_56_567# 0 0.424713f
C19670 _402_/a_728_93# 0 0.65929f
C19671 _402_/a_1296_93# 0 0.317801f
C19672 _045_ 0 0.349338f
C19673 mask\[2\] 0 1.335688f
C19674 _195_/a_67_603# 0 0.345683f
C19675 _333_/a_36_160# 0 0.386641f
C19676 _098_ 0 1.816151f
C19677 _147_ 0 0.322539f
C19678 _350_/a_49_472# 0 0.054843f
C19679 FILLER_0_12_236/a_484_472# 0 0.345058f
C19680 FILLER_0_12_236/a_36_472# 0 0.404746f
C19681 FILLER_0_12_236/a_572_375# 0 0.232991f
C19682 FILLER_0_12_236/a_124_375# 0 0.185089f
C19683 FILLER_0_2_171/a_36_472# 0 0.417394f
C19684 FILLER_0_2_171/a_124_375# 0 0.246306f
C19685 _014_ 0 0.363432f
C19686 _317_/a_36_113# 0 0.418095f
C19687 _248_/a_36_68# 0 0.69549f
C19688 FILLER_0_17_38/a_484_472# 0 0.345058f
C19689 FILLER_0_17_38/a_36_472# 0 0.404746f
C19690 FILLER_0_17_38/a_572_375# 0 0.232991f
C19691 FILLER_0_17_38/a_124_375# 0 0.185089f
C19692 _001_ 0 0.285216f
C19693 _265_/a_244_68# 0 0.138666f
C19694 _196_/a_36_160# 0 0.696445f
C19695 FILLER_0_6_90/a_484_472# 0 0.345058f
C19696 FILLER_0_6_90/a_36_472# 0 0.404746f
C19697 FILLER_0_6_90/a_572_375# 0 0.232991f
C19698 FILLER_0_6_90/a_124_375# 0 0.185089f
C19699 _183_ 0 0.356629f
C19700 _334_/a_36_160# 0 0.386641f
C19701 _282_/a_36_160# 0 0.386641f
C19702 _024_ 0 0.451815f
C19703 _009_ 0 0.397943f
C19704 _420_/a_2560_156# 0 0.016968f
C19705 _420_/a_2665_112# 0 0.62251f
C19706 _420_/a_2248_156# 0 0.371662f
C19707 _420_/a_1204_472# 0 0.012971f
C19708 _420_/a_1000_472# 0 0.291735f
C19709 _420_/a_796_472# 0 0.023206f
C19710 _420_/a_1308_423# 0 0.279043f
C19711 _420_/a_448_472# 0 0.684413f
C19712 _420_/a_36_151# 0 1.43589f
C19713 clk 0 1.162312f
C19714 FILLER_0_8_2/a_36_472# 0 0.417394f
C19715 FILLER_0_8_2/a_124_375# 0 0.246306f
C19716 FILLER_0_8_24/a_484_472# 0 0.345058f
C19717 FILLER_0_8_24/a_36_472# 0 0.404746f
C19718 FILLER_0_8_24/a_572_375# 0 0.232991f
C19719 FILLER_0_8_24/a_124_375# 0 0.185089f
C19720 _124_ 0 0.294081f
C19721 _118_ 0 1.378735f
C19722 _071_ 0 1.600488f
C19723 net9 0 1.13171f
C19724 net19 0 1.889339f
C19725 _138_ 0 0.33132f
C19726 _137_ 0 1.178616f
C19727 _335_/a_49_472# 0 0.054843f
C19728 _404_/a_36_472# 0 0.031137f
C19729 FILLER_0_20_107/a_36_472# 0 0.417394f
C19730 FILLER_0_20_107/a_124_375# 0 0.246306f
C19731 FILLER_0_9_142/a_36_472# 0 0.417394f
C19732 FILLER_0_9_142/a_124_375# 0 0.246306f
C19733 _099_ 0 1.152785f
C19734 _283_/a_36_472# 0 0.031137f
C19735 mask\[7\] 0 1.477838f
C19736 _352_/a_49_472# 0 0.054843f
C19737 _010_ 0 0.377779f
C19738 _421_/a_2560_156# 0 0.016968f
C19739 _421_/a_2665_112# 0 0.62251f
C19740 _421_/a_2248_156# 0 0.371662f
C19741 _421_/a_1204_472# 0 0.012971f
C19742 _421_/a_1000_472# 0 0.291735f
C19743 _421_/a_796_472# 0 0.023206f
C19744 _421_/a_1308_423# 0 0.279043f
C19745 _421_/a_448_472# 0 0.684413f
C19746 _421_/a_36_151# 0 1.43589f
C19747 FILLER_0_1_212/a_36_472# 0 0.417394f
C19748 FILLER_0_1_212/a_124_375# 0 0.246306f
C19749 FILLER_0_8_239/a_36_472# 0 0.417394f
C19750 FILLER_0_8_239/a_124_375# 0 0.246306f
C19751 _125_ 0 1.526603f
C19752 _058_ 0 1.483584f
C19753 FILLER_0_6_177/a_484_472# 0 0.345058f
C19754 FILLER_0_6_177/a_36_472# 0 0.404746f
C19755 FILLER_0_6_177/a_572_375# 0 0.232991f
C19756 FILLER_0_6_177/a_124_375# 0 0.185089f
C19757 state\[1\] 0 2.652405f
C19758 _267_/a_36_472# 0 0.137725f
C19759 _184_ 0 0.350066f
C19760 cal_count\[2\] 0 1.971854f
C19761 _405_/a_67_603# 0 0.345683f
C19762 _018_ 0 0.358633f
C19763 _046_ 0 0.361963f
C19764 _198_/a_67_603# 0 0.345683f
C19765 _094_ 0 1.263877f
C19766 _100_ 0 0.333135f
C19767 net36 0 2.262756f
C19768 FILLER_0_17_133/a_36_472# 0 0.417394f
C19769 FILLER_0_17_133/a_124_375# 0 0.246306f
C19770 _025_ 0 0.350324f
C19771 _148_ 0 0.325709f
C19772 _422_/a_2560_156# 0 0.016968f
C19773 _422_/a_2665_112# 0 0.62251f
C19774 _422_/a_2248_156# 0 0.371662f
C19775 _422_/a_1204_472# 0 0.012971f
C19776 _422_/a_1000_472# 0 0.291735f
C19777 _422_/a_796_472# 0 0.023206f
C19778 _422_/a_1308_423# 0 0.279043f
C19779 _422_/a_448_472# 0 0.684413f
C19780 _422_/a_36_151# 0 1.43589f
C19781 FILLER_0_1_266/a_484_472# 0 0.345058f
C19782 FILLER_0_1_266/a_36_472# 0 0.404746f
C19783 FILLER_0_1_266/a_572_375# 0 0.232991f
C19784 FILLER_0_1_266/a_124_375# 0 0.185089f
C19785 _152_ 0 0.918583f
C19786 _081_ 0 1.140656f
C19787 _370_/a_848_380# 0 0.40208f
C19788 _370_/a_124_24# 0 0.591898f
C19789 FILLER_0_24_274/a_1380_472# 0 0.345058f
C19790 FILLER_0_24_274/a_932_472# 0 0.33241f
C19791 FILLER_0_24_274/a_484_472# 0 0.33241f
C19792 FILLER_0_24_274/a_36_472# 0 0.404746f
C19793 FILLER_0_24_274/a_1468_375# 0 0.233029f
C19794 FILLER_0_24_274/a_1020_375# 0 0.171606f
C19795 FILLER_0_24_274/a_572_375# 0 0.171606f
C19796 FILLER_0_24_274/a_124_375# 0 0.185399f
C19797 _185_ 0 0.386917f
C19798 _406_/a_36_159# 0 0.374116f
C19799 _337_/a_49_472# 0 0.054843f
C19800 _199_/a_36_160# 0 0.696445f
C19801 _285_/a_36_472# 0 0.031137f
C19802 _354_/a_49_472# 0 0.054843f
C19803 _012_ 0 0.75195f
C19804 _423_/a_2560_156# 0 0.016968f
C19805 _423_/a_2665_112# 0 0.62251f
C19806 _423_/a_2248_156# 0 0.371662f
C19807 _423_/a_1204_472# 0 0.012971f
C19808 _423_/a_1000_472# 0 0.291735f
C19809 _423_/a_796_472# 0 0.023206f
C19810 _423_/a_1308_423# 0 0.279043f
C19811 _423_/a_448_472# 0 0.684413f
C19812 _423_/a_36_151# 0 1.43589f
C19813 FILLER_0_5_88/a_36_472# 0 0.417394f
C19814 FILLER_0_5_88/a_124_375# 0 0.246306f
C19815 trim_mask\[1\] 0 1.020743f
C19816 _029_ 0 0.308904f
C19817 _440_/a_2560_156# 0 0.016968f
C19818 _440_/a_2665_112# 0 0.62251f
C19819 _440_/a_2248_156# 0 0.371662f
C19820 _440_/a_1204_472# 0 0.012971f
C19821 _440_/a_1000_472# 0 0.291735f
C19822 _440_/a_796_472# 0 0.023206f
C19823 _440_/a_1308_423# 0 0.279043f
C19824 _440_/a_448_472# 0 0.684413f
C19825 _440_/a_36_151# 0 1.43589f
C19826 _159_ 0 0.351814f
C19827 _371_/a_36_113# 0 0.418095f
C19828 FILLER_0_17_56/a_484_472# 0 0.345058f
C19829 FILLER_0_17_56/a_36_472# 0 0.404746f
C19830 FILLER_0_17_56/a_572_375# 0 0.232991f
C19831 FILLER_0_17_56/a_124_375# 0 0.185089f
C19832 _083_ 0 0.527882f
C19833 _078_ 0 0.904554f
C19834 _269_/a_36_472# 0 0.031137f
C19835 _181_ 0 0.829168f
C19836 _407_/a_36_472# 0 0.031137f
C19837 _019_ 0 0.32907f
C19838 _139_ 0 0.346404f
C19839 FILLER_0_14_123/a_36_472# 0 0.417394f
C19840 FILLER_0_14_123/a_124_375# 0 0.246306f
C19841 _005_ 0 0.340993f
C19842 _101_ 0 0.280497f
C19843 _424_/a_2560_156# 0 0.016968f
C19844 _424_/a_2665_112# 0 0.62251f
C19845 _424_/a_2248_156# 0 0.371662f
C19846 _424_/a_1204_472# 0 0.012971f
C19847 _424_/a_1000_472# 0 0.291735f
C19848 _424_/a_796_472# 0 0.023206f
C19849 _424_/a_1308_423# 0 0.279043f
C19850 _424_/a_448_472# 0 0.684413f
C19851 _424_/a_36_151# 0 1.43589f
C19852 _026_ 0 0.320379f
C19853 _149_ 0 0.305496f
C19854 FILLER_0_5_54/a_1380_472# 0 0.345058f
C19855 FILLER_0_5_54/a_932_472# 0 0.33241f
C19856 FILLER_0_5_54/a_484_472# 0 0.33241f
C19857 FILLER_0_5_54/a_36_472# 0 0.404746f
C19858 FILLER_0_5_54/a_1468_375# 0 0.233029f
C19859 FILLER_0_5_54/a_1020_375# 0 0.171606f
C19860 FILLER_0_5_54/a_572_375# 0 0.171606f
C19861 FILLER_0_5_54/a_124_375# 0 0.185399f
C19862 FILLER_0_17_142/a_484_472# 0 0.345058f
C19863 FILLER_0_17_142/a_36_472# 0 0.404746f
C19864 FILLER_0_17_142/a_572_375# 0 0.232991f
C19865 FILLER_0_17_142/a_124_375# 0 0.185089f
C19866 _068_ 0 3.162692f
C19867 _076_ 0 3.812442f
C19868 _133_ 0 1.430901f
C19869 _070_ 0 3.115722f
C19870 _372_/a_170_472# 0 0.077257f
C19871 net49 0 5.140563f
C19872 _030_ 0 0.307083f
C19873 net66 0 1.472669f
C19874 _441_/a_2560_156# 0 0.016968f
C19875 _441_/a_2665_112# 0 0.62251f
C19876 _441_/a_2248_156# 0 0.371662f
C19877 _441_/a_1204_472# 0 0.012971f
C19878 _441_/a_1000_472# 0 0.291735f
C19879 _441_/a_796_472# 0 0.023206f
C19880 _441_/a_1308_423# 0 0.279043f
C19881 _441_/a_448_472# 0 0.684413f
C19882 _441_/a_36_151# 0 1.43589f
C19883 FILLER_0_5_206/a_36_472# 0 0.417394f
C19884 FILLER_0_5_206/a_124_375# 0 0.246306f
C19885 fanout49/a_36_160# 0 0.696445f
C19886 FILLER_0_8_247/a_1380_472# 0 0.345058f
C19887 FILLER_0_8_247/a_932_472# 0 0.33241f
C19888 FILLER_0_8_247/a_484_472# 0 0.33241f
C19889 FILLER_0_8_247/a_36_472# 0 0.404746f
C19890 FILLER_0_8_247/a_1468_375# 0 0.233029f
C19891 FILLER_0_8_247/a_1020_375# 0 0.171606f
C19892 FILLER_0_8_247/a_572_375# 0 0.171606f
C19893 FILLER_0_8_247/a_124_375# 0 0.185399f
C19894 FILLER_0_12_220/a_1380_472# 0 0.345058f
C19895 FILLER_0_12_220/a_932_472# 0 0.33241f
C19896 FILLER_0_12_220/a_484_472# 0 0.33241f
C19897 FILLER_0_12_220/a_36_472# 0 0.404746f
C19898 FILLER_0_12_220/a_1468_375# 0 0.233029f
C19899 FILLER_0_12_220/a_1020_375# 0 0.171606f
C19900 FILLER_0_12_220/a_572_375# 0 0.171606f
C19901 FILLER_0_12_220/a_124_375# 0 0.185399f
C19902 FILLER_0_21_286/a_484_472# 0 0.345058f
C19903 FILLER_0_21_286/a_36_472# 0 0.404746f
C19904 FILLER_0_21_286/a_572_375# 0 0.232991f
C19905 FILLER_0_21_286/a_124_375# 0 0.185089f
C19906 _140_ 0 1.276518f
C19907 _339_/a_36_160# 0 0.386641f
C19908 _095_ 0 2.689027f
C19909 _186_ 0 0.580923f
C19910 _408_/a_1936_472# 0 0.009918f
C19911 _408_/a_718_524# 0 0.005143f
C19912 _408_/a_56_524# 0 0.41096f
C19913 _408_/a_728_93# 0 0.654825f
C19914 _408_/a_1336_472# 0 0.316639f
C19915 FILLER_0_20_169/a_36_472# 0 0.417394f
C19916 FILLER_0_20_169/a_124_375# 0 0.246306f
C19917 _210_/a_67_603# 0 0.345683f
C19918 _425_/a_2560_156# 0 0.016968f
C19919 _425_/a_2665_112# 0 0.62251f
C19920 _425_/a_2248_156# 0 0.371662f
C19921 _425_/a_1204_472# 0 0.012971f
C19922 _425_/a_1000_472# 0 0.291735f
C19923 _425_/a_796_472# 0 0.023206f
C19924 _425_/a_1308_423# 0 0.279043f
C19925 _425_/a_448_472# 0 0.684413f
C19926 _425_/a_36_151# 0 1.43589f
C19927 net5 0 0.610761f
C19928 input5/a_36_113# 0 0.418095f
C19929 FILLER_0_11_78/a_484_472# 0 0.345058f
C19930 FILLER_0_11_78/a_36_472# 0 0.404746f
C19931 FILLER_0_11_78/a_572_375# 0 0.232991f
C19932 FILLER_0_11_78/a_124_375# 0 0.185089f
C19933 _102_ 0 0.335308f
C19934 _287_/a_36_472# 0 0.031137f
C19935 mask\[9\] 0 1.383606f
C19936 _356_/a_36_472# 0 0.031137f
C19937 _031_ 0 0.417351f
C19938 net69 0 1.020293f
C19939 _442_/a_2560_156# 0 0.016968f
C19940 _442_/a_2665_112# 0 0.62251f
C19941 _442_/a_2248_156# 0 0.371662f
C19942 _442_/a_1204_472# 0 0.012971f
C19943 _442_/a_1000_472# 0 0.291735f
C19944 _442_/a_796_472# 0 0.023206f
C19945 _442_/a_1308_423# 0 0.279043f
C19946 _442_/a_448_472# 0 0.684413f
C19947 _442_/a_36_151# 0 1.43589f
C19948 net64 0 2.598514f
C19949 fanout59/a_36_160# 0 0.696445f
C19950 FILLER_0_14_99/a_36_472# 0 0.417394f
C19951 FILLER_0_14_99/a_124_375# 0 0.246306f
C19952 _038_ 0 0.362839f
C19953 _136_ 0 1.345638f
C19954 _390_/a_36_68# 0 0.150048f
C19955 FILLER_0_15_282/a_484_472# 0 0.345058f
C19956 FILLER_0_15_282/a_36_472# 0 0.404746f
C19957 FILLER_0_15_282/a_572_375# 0 0.232991f
C19958 FILLER_0_15_282/a_124_375# 0 0.185089f
C19959 FILLER_0_11_124/a_36_472# 0 0.417394f
C19960 FILLER_0_11_124/a_124_375# 0 0.246306f
C19961 FILLER_0_11_135/a_36_472# 0 0.417394f
C19962 FILLER_0_11_135/a_124_375# 0 0.246306f
C19963 _188_ 0 0.349407f
C19964 cal_count\[3\] 0 1.862896f
C19965 _050_ 0 0.622354f
C19966 _211_/a_36_160# 0 0.386641f
C19967 net4 0 2.711508f
C19968 en 0 0.833743f
C19969 input4/a_36_68# 0 0.69549f
C19970 _426_/a_2560_156# 0 0.016968f
C19971 _426_/a_2665_112# 0 0.62251f
C19972 _426_/a_2248_156# 0 0.371662f
C19973 _426_/a_1204_472# 0 0.012971f
C19974 _426_/a_1000_472# 0 0.291735f
C19975 _426_/a_796_472# 0 0.023206f
C19976 _426_/a_1308_423# 0 0.279043f
C19977 _426_/a_448_472# 0 0.684413f
C19978 _426_/a_36_151# 0 1.43589f
C19979 _027_ 0 0.302949f
C19980 _150_ 0 0.320497f
C19981 FILLER_0_18_107/a_3172_472# 0 0.345058f
C19982 FILLER_0_18_107/a_2724_472# 0 0.33241f
C19983 FILLER_0_18_107/a_2276_472# 0 0.33241f
C19984 FILLER_0_18_107/a_1828_472# 0 0.33241f
C19985 FILLER_0_18_107/a_1380_472# 0 0.33241f
C19986 FILLER_0_18_107/a_932_472# 0 0.33241f
C19987 FILLER_0_18_107/a_484_472# 0 0.33241f
C19988 FILLER_0_18_107/a_36_472# 0 0.404746f
C19989 FILLER_0_18_107/a_3260_375# 0 0.233093f
C19990 FILLER_0_18_107/a_2812_375# 0 0.17167f
C19991 FILLER_0_18_107/a_2364_375# 0 0.17167f
C19992 FILLER_0_18_107/a_1916_375# 0 0.17167f
C19993 FILLER_0_18_107/a_1468_375# 0 0.17167f
C19994 FILLER_0_18_107/a_1020_375# 0 0.17167f
C19995 FILLER_0_18_107/a_572_375# 0 0.17167f
C19996 FILLER_0_18_107/a_124_375# 0 0.185915f
C19997 trim_mask\[4\] 0 0.987791f
C19998 _032_ 0 0.34876f
C19999 _443_/a_2560_156# 0 0.016968f
C20000 _443_/a_2665_112# 0 0.62251f
C20001 _443_/a_2248_156# 0 0.371662f
C20002 _443_/a_1204_472# 0 0.012971f
C20003 _443_/a_1000_472# 0 0.291735f
C20004 _443_/a_796_472# 0 0.023206f
C20005 _443_/a_1308_423# 0 0.279043f
C20006 _443_/a_448_472# 0 0.684413f
C20007 _443_/a_36_151# 0 1.43589f
C20008 _061_ 0 0.84986f
C20009 _056_ 0 2.393362f
C20010 _374_/a_36_68# 0 0.112263f
C20011 fanout58/a_36_160# 0 0.696445f
C20012 net74 0 1.237373f
C20013 fanout69/a_36_113# 0 0.418095f
C20014 _173_ 0 0.339446f
C20015 FILLER_0_3_142/a_36_472# 0 0.417394f
C20016 FILLER_0_3_142/a_124_375# 0 0.246306f
C20017 FILLER_0_17_64/a_36_472# 0 0.417394f
C20018 FILLER_0_17_64/a_124_375# 0 0.246306f
C20019 FILLER_0_11_101/a_484_472# 0 0.345058f
C20020 FILLER_0_11_101/a_36_472# 0 0.404746f
C20021 FILLER_0_11_101/a_572_375# 0 0.232991f
C20022 FILLER_0_11_101/a_124_375# 0 0.185089f
C20023 FILLER_0_22_86/a_1380_472# 0 0.345058f
C20024 FILLER_0_22_86/a_932_472# 0 0.33241f
C20025 FILLER_0_22_86/a_484_472# 0 0.33241f
C20026 FILLER_0_22_86/a_36_472# 0 0.404746f
C20027 FILLER_0_22_86/a_1468_375# 0 0.233029f
C20028 FILLER_0_22_86/a_1020_375# 0 0.171606f
C20029 FILLER_0_22_86/a_572_375# 0 0.171606f
C20030 FILLER_0_22_86/a_124_375# 0 0.185399f
C20031 net24 0 1.61895f
C20032 net3 0 0.740676f
C20033 input3/a_36_113# 0 0.418095f
C20034 _103_ 0 0.350464f
C20035 _289_/a_36_472# 0 0.031137f
C20036 _151_ 0 0.300777f
C20037 _427_/a_2560_156# 0 0.016968f
C20038 _427_/a_2665_112# 0 0.91969f
C20039 _427_/a_2248_156# 0 0.30886f
C20040 _427_/a_1204_472# 0 0.012971f
C20041 _427_/a_1000_472# 0 0.291735f
C20042 _427_/a_796_472# 0 0.023206f
C20043 _427_/a_1308_423# 0 0.279043f
C20044 _427_/a_448_472# 0 0.684413f
C20045 _427_/a_36_151# 0 1.43587f
C20046 FILLER_0_17_161/a_36_472# 0 0.417394f
C20047 FILLER_0_17_161/a_124_375# 0 0.246306f
C20048 FILLER_0_18_139/a_1380_472# 0 0.345058f
C20049 FILLER_0_18_139/a_932_472# 0 0.33241f
C20050 FILLER_0_18_139/a_484_472# 0 0.33241f
C20051 FILLER_0_18_139/a_36_472# 0 0.404746f
C20052 FILLER_0_18_139/a_1468_375# 0 0.233029f
C20053 FILLER_0_18_139/a_1020_375# 0 0.171606f
C20054 FILLER_0_18_139/a_572_375# 0 0.171606f
C20055 FILLER_0_18_139/a_124_375# 0 0.185399f
C20056 _161_ 0 0.592909f
C20057 _162_ 0 0.597238f
C20058 _375_/a_36_68# 0 0.048026f
C20059 trim_val\[0\] 0 0.742779f
C20060 net67 0 1.662327f
C20061 _444_/a_2560_156# 0 0.016968f
C20062 _444_/a_2665_112# 0 0.62251f
C20063 _444_/a_2248_156# 0 0.371662f
C20064 _444_/a_1204_472# 0 0.012971f
C20065 _444_/a_1000_472# 0 0.291735f
C20066 _444_/a_796_472# 0 0.023206f
C20067 _444_/a_1308_423# 0 0.279043f
C20068 _444_/a_448_472# 0 0.684413f
C20069 _444_/a_36_151# 0 1.43589f
C20070 net65 0 0.804072f
C20071 fanout57/a_36_113# 0 0.418095f
C20072 fanout68/a_36_113# 0 0.418095f
C20073 FILLER_0_12_2/a_484_472# 0 0.345058f
C20074 FILLER_0_12_2/a_36_472# 0 0.404746f
C20075 FILLER_0_12_2/a_572_375# 0 0.232991f
C20076 FILLER_0_12_2/a_124_375# 0 0.185089f
C20077 net79 0 1.584979f
C20078 fanout79/a_36_160# 0 0.386641f
C20079 _392_/a_36_68# 0 0.112263f
C20080 FILLER_0_13_228/a_36_472# 0 0.417394f
C20081 FILLER_0_13_228/a_124_375# 0 0.246306f
C20082 FILLER_0_13_206/a_36_472# 0 0.417394f
C20083 FILLER_0_13_206/a_124_375# 0 0.246306f
C20084 FILLER_0_20_177/a_1380_472# 0 0.345058f
C20085 FILLER_0_20_177/a_932_472# 0 0.33241f
C20086 FILLER_0_20_177/a_484_472# 0 0.33241f
C20087 FILLER_0_20_177/a_36_472# 0 0.404746f
C20088 FILLER_0_20_177/a_1468_375# 0 0.233029f
C20089 FILLER_0_20_177/a_1020_375# 0 0.171606f
C20090 FILLER_0_20_177/a_572_375# 0 0.171606f
C20091 FILLER_0_20_177/a_124_375# 0 0.185399f
C20092 _051_ 0 0.349381f
C20093 _213_/a_67_603# 0 0.345683f
C20094 net2 0 0.461658f
C20095 input2/a_36_113# 0 0.418095f
C20096 _129_ 0 0.926508f
C20097 _131_ 0 1.734297f
C20098 _359_/a_36_488# 0 0.101145f
C20099 FILLER_0_11_64/a_36_472# 0 0.417394f
C20100 FILLER_0_11_64/a_124_375# 0 0.246306f
C20101 state\[2\] 0 0.607433f
C20102 net53 0 4.483899f
C20103 _017_ 0 0.334329f
C20104 net70 0 1.238296f
C20105 _428_/a_2560_156# 0 0.016968f
C20106 _428_/a_2665_112# 0 0.62251f
C20107 _428_/a_2248_156# 0 0.371662f
C20108 _428_/a_1204_472# 0 0.012971f
C20109 _428_/a_1000_472# 0 0.291735f
C20110 _428_/a_796_472# 0 0.023206f
C20111 _428_/a_1308_423# 0 0.279043f
C20112 _428_/a_448_472# 0 0.684413f
C20113 _428_/a_36_151# 0 1.43589f
C20114 FILLER_0_5_72/a_1380_472# 0 0.345058f
C20115 FILLER_0_5_72/a_932_472# 0 0.33241f
C20116 FILLER_0_5_72/a_484_472# 0 0.33241f
C20117 FILLER_0_5_72/a_36_472# 0 0.404746f
C20118 FILLER_0_5_72/a_1468_375# 0 0.233029f
C20119 FILLER_0_5_72/a_1020_375# 0 0.171606f
C20120 FILLER_0_5_72/a_572_375# 0 0.171606f
C20121 FILLER_0_5_72/a_124_375# 0 0.185399f
C20122 _376_/a_36_160# 0 0.386641f
C20123 trim_val\[1\] 0 0.683578f
C20124 _445_/a_2560_156# 0 0.016968f
C20125 _445_/a_2665_112# 0 0.62251f
C20126 _445_/a_2248_156# 0 0.371662f
C20127 _445_/a_1204_472# 0 0.012971f
C20128 _445_/a_1000_472# 0 0.291735f
C20129 _445_/a_796_472# 0 0.023206f
C20130 _445_/a_1308_423# 0 0.279043f
C20131 _445_/a_448_472# 0 0.684413f
C20132 _445_/a_36_151# 0 1.43589f
C20133 fanout67/a_36_160# 0 0.386641f
C20134 fanout56/a_36_113# 0 0.418095f
C20135 net78 0 0.686263f
C20136 fanout78/a_36_113# 0 0.418095f
C20137 _174_ 0 0.979741f
C20138 FILLER_0_0_198/a_36_472# 0 0.417394f
C20139 FILLER_0_0_198/a_124_375# 0 0.246306f
C20140 FILLER_0_15_290/a_36_472# 0 0.417394f
C20141 FILLER_0_15_290/a_124_375# 0 0.246306f
C20142 FILLER_0_24_290/a_36_472# 0 0.417394f
C20143 FILLER_0_24_290/a_124_375# 0 0.246306f
C20144 FILLER_0_4_107/a_1380_472# 0 0.345058f
C20145 FILLER_0_4_107/a_932_472# 0 0.33241f
C20146 FILLER_0_4_107/a_484_472# 0 0.33241f
C20147 FILLER_0_4_107/a_36_472# 0 0.404746f
C20148 FILLER_0_4_107/a_1468_375# 0 0.233029f
C20149 FILLER_0_4_107/a_1020_375# 0 0.171606f
C20150 FILLER_0_4_107/a_572_375# 0 0.171606f
C20151 FILLER_0_4_107/a_124_375# 0 0.185399f
C20152 FILLER_0_7_104/a_1380_472# 0 0.345058f
C20153 FILLER_0_7_104/a_932_472# 0 0.33241f
C20154 FILLER_0_7_104/a_484_472# 0 0.33241f
C20155 FILLER_0_7_104/a_36_472# 0 0.404746f
C20156 FILLER_0_7_104/a_1468_375# 0 0.233029f
C20157 FILLER_0_7_104/a_1020_375# 0 0.171606f
C20158 FILLER_0_7_104/a_572_375# 0 0.171606f
C20159 FILLER_0_7_104/a_124_375# 0 0.185399f
C20160 _214_/a_36_160# 0 0.386641f
C20161 net1 0 0.364811f
C20162 input1/a_36_113# 0 0.418095f
C20163 _429_/a_2560_156# 0 0.016968f
C20164 _429_/a_2665_112# 0 0.62251f
C20165 _429_/a_2248_156# 0 0.371662f
C20166 _429_/a_1204_472# 0 0.012971f
C20167 _429_/a_1000_472# 0 0.291735f
C20168 _429_/a_796_472# 0 0.023206f
C20169 _429_/a_1308_423# 0 0.279043f
C20170 _429_/a_448_472# 0 0.684413f
C20171 _429_/a_36_151# 0 1.43589f
C20172 _011_ 0 0.278979f
C20173 _377_/a_36_472# 0 0.031137f
C20174 fanout66/a_36_113# 0 0.418095f
C20175 _035_ 0 0.327801f
C20176 _446_/a_2560_156# 0 0.016968f
C20177 _446_/a_2665_112# 0 0.62251f
C20178 _446_/a_2248_156# 0 0.371662f
C20179 _446_/a_1204_472# 0 0.012971f
C20180 _446_/a_1000_472# 0 0.291735f
C20181 _446_/a_796_472# 0 0.023206f
C20182 _446_/a_1308_423# 0 0.279043f
C20183 _446_/a_448_472# 0 0.684413f
C20184 _446_/a_36_151# 0 1.43589f
C20185 fanout77/a_36_113# 0 0.418095f
C20186 FILLER_0_5_212/a_36_472# 0 0.417394f
C20187 FILLER_0_5_212/a_124_375# 0 0.246306f
C20188 fanout55/a_36_160# 0 0.696445f
C20189 _175_ 0 0.344159f
C20190 _394_/a_1936_472# 0 0.009918f
C20191 _394_/a_718_524# 0 0.005143f
C20192 _394_/a_56_524# 0 0.41096f
C20193 _394_/a_728_93# 0 0.654825f
C20194 _394_/a_1336_472# 0 0.316639f
C20195 FILLER_0_3_172/a_3172_472# 0 0.345058f
C20196 FILLER_0_3_172/a_2724_472# 0 0.33241f
C20197 FILLER_0_3_172/a_2276_472# 0 0.33241f
C20198 FILLER_0_3_172/a_1828_472# 0 0.33241f
C20199 FILLER_0_3_172/a_1380_472# 0 0.33241f
C20200 FILLER_0_3_172/a_932_472# 0 0.33241f
C20201 FILLER_0_3_172/a_484_472# 0 0.33241f
C20202 FILLER_0_3_172/a_36_472# 0 0.404746f
C20203 FILLER_0_3_172/a_3260_375# 0 0.233093f
C20204 FILLER_0_3_172/a_2812_375# 0 0.17167f
C20205 FILLER_0_3_172/a_2364_375# 0 0.17167f
C20206 FILLER_0_3_172/a_1916_375# 0 0.17167f
C20207 FILLER_0_3_172/a_1468_375# 0 0.17167f
C20208 FILLER_0_3_172/a_1020_375# 0 0.17167f
C20209 FILLER_0_3_172/a_572_375# 0 0.17167f
C20210 FILLER_0_3_172/a_124_375# 0 0.185915f
C20211 FILLER_0_17_72/a_3172_472# 0 0.345058f
C20212 FILLER_0_17_72/a_2724_472# 0 0.33241f
C20213 FILLER_0_17_72/a_2276_472# 0 0.33241f
C20214 FILLER_0_17_72/a_1828_472# 0 0.33241f
C20215 FILLER_0_17_72/a_1380_472# 0 0.33241f
C20216 FILLER_0_17_72/a_932_472# 0 0.33241f
C20217 FILLER_0_17_72/a_484_472# 0 0.33241f
C20218 FILLER_0_17_72/a_36_472# 0 0.404746f
C20219 FILLER_0_17_72/a_3260_375# 0 0.233093f
C20220 FILLER_0_17_72/a_2812_375# 0 0.17167f
C20221 FILLER_0_17_72/a_2364_375# 0 0.17167f
C20222 FILLER_0_17_72/a_1916_375# 0 0.17167f
C20223 FILLER_0_17_72/a_1468_375# 0 0.17167f
C20224 FILLER_0_17_72/a_1020_375# 0 0.17167f
C20225 FILLER_0_17_72/a_572_375# 0 0.17167f
C20226 FILLER_0_17_72/a_124_375# 0 0.185915f
C20227 FILLER_0_2_93/a_484_472# 0 0.345058f
C20228 FILLER_0_2_93/a_36_472# 0 0.404746f
C20229 FILLER_0_2_93/a_572_375# 0 0.232991f
C20230 FILLER_0_2_93/a_124_375# 0 0.185089f
C20231 FILLER_0_11_142/a_484_472# 0 0.345058f
C20232 FILLER_0_11_142/a_36_472# 0 0.404746f
C20233 FILLER_0_11_142/a_572_375# 0 0.232991f
C20234 FILLER_0_11_142/a_124_375# 0 0.185089f
C20235 net25 0 1.803174f
C20236 _232_/a_67_603# 0 0.345683f
C20237 net35 0 1.844415f
C20238 mask\[8\] 0 1.276111f
C20239 _301_/a_36_472# 0 0.031137f
C20240 _033_ 0 0.323682f
C20241 _165_ 0 0.331995f
C20242 FILLER_0_3_2/a_36_472# 0 0.417394f
C20243 FILLER_0_3_2/a_124_375# 0 0.246306f
C20244 trim_val\[3\] 0 0.719615f
C20245 _036_ 0 0.369206f
C20246 net68 0 1.735004f
C20247 _447_/a_2560_156# 0 0.016968f
C20248 _447_/a_2665_112# 0 0.62251f
C20249 _447_/a_2248_156# 0 0.371662f
C20250 _447_/a_1204_472# 0 0.012971f
C20251 _447_/a_1000_472# 0 0.291735f
C20252 _447_/a_796_472# 0 0.023206f
C20253 _447_/a_1308_423# 0 0.279043f
C20254 _447_/a_448_472# 0 0.684413f
C20255 _447_/a_36_151# 0 1.43589f
C20256 FILLER_0_19_28/a_484_472# 0 0.345058f
C20257 FILLER_0_19_28/a_36_472# 0 0.404746f
C20258 FILLER_0_19_28/a_572_375# 0 0.232991f
C20259 FILLER_0_19_28/a_124_375# 0 0.185089f
C20260 fanout65/a_36_113# 0 0.418095f
C20261 fanout76/a_36_160# 0 0.386641f
C20262 net54 0 5.456963f
C20263 fanout54/a_36_160# 0 0.696445f
C20264 FILLER_0_4_49/a_484_472# 0 0.345058f
C20265 FILLER_0_4_49/a_36_472# 0 0.404746f
C20266 FILLER_0_4_49/a_572_375# 0 0.232991f
C20267 FILLER_0_4_49/a_124_375# 0 0.185089f
C20268 _176_ 0 0.804011f
C20269 _085_ 0 2.280803f
C20270 _116_ 0 1.959915f
C20271 _395_/a_36_488# 0 0.101145f
C20272 FILLER_0_14_50/a_36_472# 0 0.417394f
C20273 FILLER_0_14_50/a_124_375# 0 0.246306f
C20274 FILLER_0_8_263/a_36_472# 0 0.417394f
C20275 FILLER_0_8_263/a_124_375# 0 0.246306f
C20276 FILLER_0_0_130/a_36_472# 0 0.417394f
C20277 FILLER_0_0_130/a_124_375# 0 0.246306f
C20278 FILLER_0_16_255/a_36_472# 0 0.417394f
C20279 FILLER_0_16_255/a_124_375# 0 0.246306f
C20280 FILLER_0_7_59/a_484_472# 0 0.345058f
C20281 FILLER_0_7_59/a_36_472# 0 0.404746f
C20282 FILLER_0_7_59/a_572_375# 0 0.232991f
C20283 FILLER_0_7_59/a_124_375# 0 0.185089f
C20284 ctlp[2] 0 0.17528f
C20285 output19/a_224_472# 0 2.38465f
C20286 FILLER_0_7_146/a_36_472# 0 0.417394f
C20287 FILLER_0_7_146/a_124_375# 0 0.246306f
C20288 _216_/a_67_603# 0 0.345683f
C20289 FILLER_0_15_116/a_484_472# 0 0.345058f
C20290 FILLER_0_15_116/a_36_472# 0 0.404746f
C20291 FILLER_0_15_116/a_572_375# 0 0.232991f
C20292 FILLER_0_15_116/a_124_375# 0 0.185089f
C20293 _063_ 0 0.370155f
C20294 _233_/a_36_160# 0 0.386641f
C20295 FILLER_0_21_28/a_3172_472# 0 0.345058f
C20296 FILLER_0_21_28/a_2724_472# 0 0.33241f
C20297 FILLER_0_21_28/a_2276_472# 0 0.33241f
C20298 FILLER_0_21_28/a_1828_472# 0 0.33241f
C20299 FILLER_0_21_28/a_1380_472# 0 0.33241f
C20300 FILLER_0_21_28/a_932_472# 0 0.33241f
C20301 FILLER_0_21_28/a_484_472# 0 0.33241f
C20302 FILLER_0_21_28/a_36_472# 0 0.404746f
C20303 FILLER_0_21_28/a_3260_375# 0 0.233093f
C20304 FILLER_0_21_28/a_2812_375# 0 0.17167f
C20305 FILLER_0_21_28/a_2364_375# 0 0.17167f
C20306 FILLER_0_21_28/a_1916_375# 0 0.17167f
C20307 FILLER_0_21_28/a_1468_375# 0 0.17167f
C20308 FILLER_0_21_28/a_1020_375# 0 0.17167f
C20309 FILLER_0_21_28/a_572_375# 0 0.17167f
C20310 FILLER_0_21_28/a_124_375# 0 0.185915f
C20311 _110_ 0 0.323912f
C20312 _379_/a_36_472# 0 0.031137f
C20313 trim_val\[4\] 0 0.662409f
C20314 net76 0 1.454269f
C20315 _448_/a_2560_156# 0 0.016968f
C20316 _448_/a_2665_112# 0 0.62251f
C20317 _448_/a_2248_156# 0 0.371662f
C20318 _448_/a_1204_472# 0 0.012971f
C20319 _448_/a_1000_472# 0 0.291735f
C20320 _448_/a_796_472# 0 0.023206f
C20321 _448_/a_1308_423# 0 0.279043f
C20322 _448_/a_448_472# 0 0.684413f
C20323 _448_/a_36_151# 0 1.43589f
C20324 fanout64/a_36_160# 0 0.386641f
C20325 fanout75/a_36_113# 0 0.418095f
C20326 _250_/a_36_68# 0 0.69549f
C20327 net56 0 0.843396f
C20328 fanout53/a_36_160# 0 0.696445f
C20329 _177_ 0 0.358286f
C20330 result[2] 0 0.230851f
C20331 net29 0 1.802718f
C20332 output29/a_224_472# 0 2.38465f
C20333 ctlp[1] 0 0.17418f
C20334 output18/a_224_472# 0 2.38465f
C20335 FILLER_0_14_181/a_36_472# 0 0.417394f
C20336 FILLER_0_14_181/a_124_375# 0 0.246306f
C20337 _052_ 0 0.569133f
C20338 _217_/a_36_160# 0 0.386641f
C20339 net44 0 1.407054f
C20340 _303_/a_36_472# 0 0.031137f
C20341 en_co_clk 0 0.346872f
C20342 net55 0 5.119958f
C20343 net72 0 1.366255f
C20344 _449_/a_2560_156# 0 0.016968f
C20345 _449_/a_2665_112# 0 0.62251f
C20346 _449_/a_2248_156# 0 0.371662f
C20347 _449_/a_1204_472# 0 0.012971f
C20348 _449_/a_1000_472# 0 0.291735f
C20349 _449_/a_796_472# 0 0.023206f
C20350 _449_/a_1308_423# 0 0.279043f
C20351 _449_/a_448_472# 0 0.684413f
C20352 _449_/a_36_151# 0 1.43589f
C20353 fanout52/a_36_160# 0 0.696445f
C20354 net82 0 0.706042f
C20355 fanout74/a_36_113# 0 0.418095f
C20356 FILLER_0_10_28/a_36_472# 0 0.417394f
C20357 FILLER_0_10_28/a_124_375# 0 0.246306f
C20358 mask\[0\] 0 2.242948f
C20359 _320_/a_36_472# 0 0.137725f
C20360 fanout63/a_36_160# 0 0.696445f
C20361 FILLER_0_14_81/a_36_472# 0 0.417394f
C20362 FILLER_0_14_81/a_124_375# 0 0.246306f
C20363 _397_/a_36_472# 0 0.031137f
C20364 FILLER_0_13_212/a_1380_472# 0 0.345058f
C20365 FILLER_0_13_212/a_932_472# 0 0.33241f
C20366 FILLER_0_13_212/a_484_472# 0 0.33241f
C20367 FILLER_0_13_212/a_36_472# 0 0.404746f
C20368 FILLER_0_13_212/a_1468_375# 0 0.233029f
C20369 FILLER_0_13_212/a_1020_375# 0 0.171606f
C20370 FILLER_0_13_212/a_572_375# 0 0.171606f
C20371 FILLER_0_13_212/a_124_375# 0 0.185399f
C20372 trim[1] 0 0.793787f
C20373 net39 0 1.445128f
C20374 output39/a_224_472# 0 2.38465f
C20375 result[1] 0 0.229507f
C20376 net28 0 1.759728f
C20377 output28/a_224_472# 0 2.38465f
C20378 ctlp[0] 0 1.002286f
C20379 output17/a_224_472# 0 2.38465f
C20380 FILLER_0_16_37/a_36_472# 0 0.417394f
C20381 FILLER_0_16_37/a_124_375# 0 0.246306f
C20382 net26 0 1.671545f
C20383 _064_ 0 0.581481f
C20384 trim_val\[2\] 0 0.65354f
C20385 trim_mask\[2\] 0 0.92551f
C20386 _235_/a_67_603# 0 0.345683f
C20387 _013_ 0 0.48783f
C20388 _111_ 0 0.369652f
C20389 FILLER_0_18_177/a_3172_472# 0 0.345058f
C20390 FILLER_0_18_177/a_2724_472# 0 0.33241f
C20391 FILLER_0_18_177/a_2276_472# 0 0.33241f
C20392 FILLER_0_18_177/a_1828_472# 0 0.33241f
C20393 FILLER_0_18_177/a_1380_472# 0 0.33241f
C20394 FILLER_0_18_177/a_932_472# 0 0.33241f
C20395 FILLER_0_18_177/a_484_472# 0 0.33241f
C20396 FILLER_0_18_177/a_36_472# 0 0.404746f
C20397 FILLER_0_18_177/a_3260_375# 0 0.233093f
C20398 FILLER_0_18_177/a_2812_375# 0 0.17167f
C20399 FILLER_0_18_177/a_2364_375# 0 0.17167f
C20400 FILLER_0_18_177/a_1916_375# 0 0.17167f
C20401 FILLER_0_18_177/a_1468_375# 0 0.17167f
C20402 FILLER_0_18_177/a_1020_375# 0 0.17167f
C20403 FILLER_0_18_177/a_572_375# 0 0.17167f
C20404 FILLER_0_18_177/a_124_375# 0 0.185915f
C20405 FILLER_0_18_100/a_36_472# 0 0.417394f
C20406 FILLER_0_18_100/a_124_375# 0 0.246306f
C20407 _073_ 0 0.953711f
C20408 _126_ 0 2.036767f
C20409 _069_ 0 2.034557f
C20410 _321_/a_170_472# 0 0.077257f
C20411 fanout51/a_36_113# 0 0.418095f
C20412 net62 0 4.932099f
C20413 fanout62/a_36_160# 0 0.696445f
C20414 fanout73/a_36_113# 0 0.418095f
C20415 FILLER_0_19_47/a_484_472# 0 0.345058f
C20416 FILLER_0_19_47/a_36_472# 0 0.404746f
C20417 FILLER_0_19_47/a_572_375# 0 0.232991f
C20418 FILLER_0_19_47/a_124_375# 0 0.185089f
C20419 FILLER_0_14_91/a_484_472# 0 0.345058f
C20420 FILLER_0_14_91/a_36_472# 0 0.404746f
C20421 FILLER_0_14_91/a_572_375# 0 0.232991f
C20422 FILLER_0_14_91/a_124_375# 0 0.185089f
C20423 FILLER_0_10_214/a_36_472# 0 0.417394f
C20424 FILLER_0_10_214/a_124_375# 0 0.246306f
C20425 FILLER_0_10_247/a_36_472# 0 0.417394f
C20426 FILLER_0_10_247/a_124_375# 0 0.246306f
C20427 _178_ 0 1.252435f
C20428 _398_/a_36_113# 0 0.418095f
C20429 FILLER_0_16_241/a_36_472# 0 0.417394f
C20430 FILLER_0_16_241/a_124_375# 0 0.246306f
C20431 trim[0] 0 0.796081f
C20432 net38 0 1.529392f
C20433 output38/a_224_472# 0 2.38465f
C20434 ctln[9] 0 0.904836f
C20435 net16 0 1.295744f
C20436 output16/a_224_472# 0 2.38465f
C20437 result[0] 0 0.56622f
C20438 output27/a_224_472# 0 2.38465f
C20439 _219_/a_36_160# 0 0.386641f
C20440 FILLER_0_20_193/a_484_472# 0 0.345058f
C20441 FILLER_0_20_193/a_36_472# 0 0.404746f
C20442 FILLER_0_20_193/a_572_375# 0 0.232991f
C20443 FILLER_0_20_193/a_124_375# 0 0.185089f
C20444 _236_/a_36_160# 0 0.696445f
C20445 _112_ 0 0.308886f
C20446 _305_/a_36_159# 0 0.374116f
C20447 _074_ 0 1.813232f
C20448 _253_/a_36_68# 0 0.061249f
C20449 net50 0 4.486121f
C20450 net52 0 3.536016f
C20451 fanout50/a_36_160# 0 0.696445f
C20452 FILLER_0_10_37/a_36_472# 0 0.417394f
C20453 FILLER_0_10_37/a_124_375# 0 0.246306f
C20454 fanout72/a_36_113# 0 0.418095f
C20455 fanout61/a_36_113# 0 0.418095f
C20456 _128_ 0 0.447252f
C20457 _127_ 0 1.291729f
C20458 _322_/a_848_380# 0 0.40208f
C20459 _322_/a_124_24# 0 0.591898f
C20460 _088_ 0 0.457961f
C20461 _079_ 0 1.114894f
C20462 _087_ 0 0.601674f
C20463 _270_/a_36_472# 0 0.031137f
C20464 FILLER_0_4_123/a_36_472# 0 0.417394f
C20465 FILLER_0_4_123/a_124_375# 0 0.246306f
C20466 FILLER_0_17_218/a_484_472# 0 0.345058f
C20467 FILLER_0_17_218/a_36_472# 0 0.404746f
C20468 FILLER_0_17_218/a_572_375# 0 0.232991f
C20469 FILLER_0_17_218/a_124_375# 0 0.185089f
C20470 sample 0 0.508149f
C20471 output37/a_224_472# 0 2.38465f
C20472 valid 0 0.272072f
C20473 net48 0 1.219262f
C20474 output48/a_224_472# 0 2.38465f
C20475 ctln[8] 0 1.547984f
C20476 net15 0 1.440851f
C20477 output15/a_224_472# 0 2.38465f
C20478 ctlp[9] 0 0.73349f
C20479 output26/a_224_472# 0 2.38465f
C20480 FILLER_0_16_57/a_1380_472# 0 0.345058f
C20481 FILLER_0_16_57/a_932_472# 0 0.33241f
C20482 FILLER_0_16_57/a_484_472# 0 0.33241f
C20483 FILLER_0_16_57/a_36_472# 0 0.404746f
C20484 FILLER_0_16_57/a_1468_375# 0 0.233029f
C20485 FILLER_0_16_57/a_1020_375# 0 0.171606f
C20486 FILLER_0_16_57/a_572_375# 0 0.171606f
C20487 FILLER_0_16_57/a_124_375# 0 0.185399f
C20488 _306_/a_36_68# 0 0.69549f
C20489 _072_ 0 2.604301f
C20490 fanout82/a_36_113# 0 0.418095f
C20491 _015_ 0 0.406653f
C20492 _323_/a_36_113# 0 0.418095f
C20493 net60 0 5.024503f
C20494 net61 0 1.666523f
C20495 fanout60/a_36_160# 0 0.696445f
C20496 fanout71/a_36_113# 0 0.418095f
C20497 FILLER_0_6_239/a_36_472# 0 0.417394f
C20498 FILLER_0_6_239/a_124_375# 0 0.246306f
C20499 FILLER_0_4_99/a_36_472# 0 0.417394f
C20500 FILLER_0_4_99/a_124_375# 0 0.246306f
C20501 net57 0 1.383718f
C20502 FILLER_0_10_256/a_36_472# 0 0.417394f
C20503 FILLER_0_10_256/a_124_375# 0 0.246306f
C20504 cal_itt\[3\] 0 1.854962f
C20505 _340_/a_36_160# 0 0.386641f
C20506 FILLER_0_4_177/a_484_472# 0 0.345058f
C20507 FILLER_0_4_177/a_36_472# 0 0.404746f
C20508 FILLER_0_4_177/a_572_375# 0 0.232991f
C20509 FILLER_0_4_177/a_124_375# 0 0.185089f
C20510 FILLER_0_4_144/a_484_472# 0 0.345058f
C20511 FILLER_0_4_144/a_36_472# 0 0.404746f
C20512 FILLER_0_4_144/a_572_375# 0 0.232991f
C20513 FILLER_0_4_144/a_124_375# 0 0.185089f
C20514 ctln[7] 0 1.265946f
C20515 output14/a_224_472# 0 2.38465f
C20516 result[9] 0 0.8197f
C20517 output36/a_224_472# 0 2.38465f
C20518 trimb[4] 0 0.752332f
C20519 output47/a_224_472# 0 2.38465f
C20520 ctlp[8] 0 1.136333f
C20521 output25/a_224_472# 0 2.38465f
C20522 FILLER_0_12_136/a_1380_472# 0 0.345058f
C20523 FILLER_0_12_136/a_932_472# 0 0.33241f
C20524 FILLER_0_12_136/a_484_472# 0 0.33241f
C20525 FILLER_0_12_136/a_36_472# 0 0.404746f
C20526 FILLER_0_12_136/a_1468_375# 0 0.233029f
C20527 FILLER_0_12_136/a_1020_375# 0 0.171606f
C20528 FILLER_0_12_136/a_572_375# 0 0.171606f
C20529 FILLER_0_12_136/a_124_375# 0 0.185399f
C20530 FILLER_0_16_89/a_1380_472# 0 0.345058f
C20531 FILLER_0_16_89/a_932_472# 0 0.33241f
C20532 FILLER_0_16_89/a_484_472# 0 0.33241f
C20533 FILLER_0_16_89/a_36_472# 0 0.404746f
C20534 FILLER_0_16_89/a_1468_375# 0 0.233029f
C20535 FILLER_0_16_89/a_1020_375# 0 0.171606f
C20536 FILLER_0_16_89/a_572_375# 0 0.171606f
C20537 FILLER_0_16_89/a_124_375# 0 0.185399f
C20538 FILLER_0_21_125/a_484_472# 0 0.345058f
C20539 FILLER_0_21_125/a_36_472# 0 0.404746f
C20540 FILLER_0_21_125/a_572_375# 0 0.232991f
C20541 FILLER_0_21_125/a_124_375# 0 0.185089f
C20542 _238_/a_67_603# 0 0.345683f
C20543 _096_ 0 2.205532f
C20544 _093_ 0 1.893313f
C20545 FILLER_0_19_55/a_36_472# 0 0.417394f
C20546 FILLER_0_19_55/a_124_375# 0 0.246306f
C20547 net81 0 1.738987f
C20548 fanout81/a_36_160# 0 0.386641f
C20549 _057_ 0 1.600886f
C20550 _255_/a_224_552# 0 1.31114f
C20551 net73 0 1.058857f
C20552 fanout70/a_36_113# 0 0.418095f
C20553 _003_ 0 0.3064f
C20554 _089_ 0 0.36777f
C20555 _272_/a_36_472# 0 0.031137f
C20556 _187_ 0 0.311229f
C20557 _410_/a_36_68# 0 0.112263f
C20558 _141_ 0 1.249289f
C20559 mask\[3\] 0 1.26722f
C20560 _341_/a_49_472# 0 0.054843f
C20561 cal 0 0.793393f
C20562 FILLER_0_7_195/a_36_472# 0 0.417394f
C20563 FILLER_0_7_195/a_124_375# 0 0.246306f
C20564 FILLER_0_7_162/a_36_472# 0 0.417394f
C20565 FILLER_0_7_162/a_124_375# 0 0.246306f
C20566 ctln[6] 0 1.451644f
C20567 output13/a_224_472# 0 2.38465f
C20568 FILLER_0_18_2/a_3172_472# 0 0.345058f
C20569 FILLER_0_18_2/a_2724_472# 0 0.33241f
C20570 FILLER_0_18_2/a_2276_472# 0 0.33241f
C20571 FILLER_0_18_2/a_1828_472# 0 0.33241f
C20572 FILLER_0_18_2/a_1380_472# 0 0.33241f
C20573 FILLER_0_18_2/a_932_472# 0 0.33241f
C20574 FILLER_0_18_2/a_484_472# 0 0.33241f
C20575 FILLER_0_18_2/a_36_472# 0 0.404746f
C20576 FILLER_0_18_2/a_3260_375# 0 0.233093f
C20577 FILLER_0_18_2/a_2812_375# 0 0.17167f
C20578 FILLER_0_18_2/a_2364_375# 0 0.17167f
C20579 FILLER_0_18_2/a_1916_375# 0 0.17167f
C20580 FILLER_0_18_2/a_1468_375# 0 0.17167f
C20581 FILLER_0_18_2/a_1020_375# 0 0.17167f
C20582 FILLER_0_18_2/a_572_375# 0 0.17167f
C20583 FILLER_0_18_2/a_124_375# 0 0.185915f
C20584 trimb[3] 0 0.34698f
C20585 net46 0 1.13395f
C20586 output46/a_224_472# 0 2.38465f
C20587 result[8] 0 0.68837f
C20588 output35/a_224_472# 0 2.38465f
C20589 ctlp[7] 0 0.83567f
C20590 output24/a_224_472# 0 2.38465f
C20591 FILLER_0_8_107/a_36_472# 0 0.417394f
C20592 FILLER_0_8_107/a_124_375# 0 0.246306f
C20593 FILLER_0_12_124/a_36_472# 0 0.417394f
C20594 FILLER_0_12_124/a_124_375# 0 0.246306f
C20595 net41 0 1.746759f
C20596 _065_ 0 0.523724f
C20597 _239_/a_36_160# 0 0.696445f
C20598 FILLER_0_1_98/a_36_472# 0 0.417394f
C20599 FILLER_0_1_98/a_124_375# 0 0.246306f
C20600 _115_ 0 1.281516f
C20601 _114_ 0 2.293579f
C20602 _308_/a_848_380# 0 0.40208f
C20603 _308_/a_124_24# 0 0.591898f
C20604 _256_/a_36_68# 0 0.063181f
C20605 FILLER_0_10_78/a_1380_472# 0 0.345058f
C20606 FILLER_0_10_78/a_932_472# 0 0.33241f
C20607 FILLER_0_10_78/a_484_472# 0 0.33241f
C20608 FILLER_0_10_78/a_36_472# 0 0.404746f
C20609 FILLER_0_10_78/a_1468_375# 0 0.233029f
C20610 FILLER_0_10_78/a_1020_375# 0 0.171606f
C20611 FILLER_0_10_78/a_572_375# 0 0.171606f
C20612 FILLER_0_10_78/a_124_375# 0 0.185399f
C20613 _130_ 0 0.304085f
C20614 net80 0 1.375599f
C20615 fanout80/a_36_113# 0 0.418095f
C20616 net58 0 5.308423f
C20617 _000_ 0 0.382358f
C20618 net75 0 1.474299f
C20619 _411_/a_2560_156# 0 0.016968f
C20620 _411_/a_2665_112# 0 0.62251f
C20621 _411_/a_2248_156# 0 0.371662f
C20622 _411_/a_1204_472# 0 0.012971f
C20623 _411_/a_1000_472# 0 0.291735f
C20624 _411_/a_796_472# 0 0.023206f
C20625 _411_/a_1308_423# 0 0.279043f
C20626 _411_/a_448_472# 0 0.684413f
C20627 _411_/a_36_151# 0 1.43589f
C20628 state\[0\] 0 0.680109f
C20629 _273_/a_36_68# 0 0.69549f
C20630 _142_ 0 0.324372f
C20631 FILLER_0_9_223/a_484_472# 0 0.345058f
C20632 FILLER_0_9_223/a_36_472# 0 0.404746f
C20633 FILLER_0_9_223/a_572_375# 0 0.232991f
C20634 FILLER_0_9_223/a_124_375# 0 0.185089f
C20635 FILLER_0_4_197/a_1380_472# 0 0.345058f
C20636 FILLER_0_4_197/a_932_472# 0 0.33241f
C20637 FILLER_0_4_197/a_484_472# 0 0.33241f
C20638 FILLER_0_4_197/a_36_472# 0 0.404746f
C20639 FILLER_0_4_197/a_1468_375# 0 0.233029f
C20640 FILLER_0_4_197/a_1020_375# 0 0.171606f
C20641 FILLER_0_4_197/a_572_375# 0 0.171606f
C20642 FILLER_0_4_197/a_124_375# 0 0.185399f
C20643 FILLER_0_17_226/a_36_472# 0 0.417394f
C20644 FILLER_0_17_226/a_124_375# 0 0.246306f
C20645 FILLER_0_5_109/a_484_472# 0 0.345058f
C20646 FILLER_0_5_109/a_36_472# 0 0.404746f
C20647 FILLER_0_5_109/a_572_375# 0 0.232991f
C20648 FILLER_0_5_109/a_124_375# 0 0.185089f
C20649 ctln[5] 0 1.585113f
C20650 output12/a_224_472# 0 2.38465f
C20651 result[7] 0 0.24756f
C20652 net34 0 1.724665f
C20653 output34/a_224_472# 0 2.38465f
C20654 trimb[2] 0 0.839614f
C20655 net45 0 1.12041f
C20656 output45/a_224_472# 0 2.38465f
C20657 ctlp[6] 0 1.243017f
C20658 output23/a_224_472# 0 2.38465f
C20659 FILLER_0_15_142/a_484_472# 0 0.345058f
C20660 FILLER_0_15_142/a_36_472# 0 0.404746f
C20661 FILLER_0_15_142/a_572_375# 0 0.232991f
C20662 FILLER_0_15_142/a_124_375# 0 0.185089f
C20663 _077_ 0 1.645892f
C20664 _075_ 0 0.374516f
C20665 _257_/a_36_472# 0 0.031137f
C20666 _326_/a_36_160# 0 0.696445f
C20667 _412_/a_2560_156# 0 0.016968f
C20668 _412_/a_2665_112# 0 0.62251f
C20669 _412_/a_2248_156# 0 0.371662f
C20670 _412_/a_1204_472# 0 0.012971f
C20671 _412_/a_1000_472# 0 0.291735f
C20672 _412_/a_796_472# 0 0.023206f
C20673 _412_/a_1308_423# 0 0.279043f
C20674 _412_/a_448_472# 0 0.684413f
C20675 _412_/a_36_151# 0 1.43589f
C20676 _091_ 0 1.841339f
C20677 _274_/a_36_68# 0 0.063181f
C20678 _143_ 0 0.329289f
C20679 mask\[4\] 0 1.300438f
C20680 _343_/a_49_472# 0 0.054843f
C20681 FILLER_0_13_65/a_36_472# 0 0.417394f
C20682 FILLER_0_13_65/a_124_375# 0 0.246306f
C20683 _360_/a_36_160# 0 0.386641f
C20684 FILLER_0_4_185/a_36_472# 0 0.417394f
C20685 FILLER_0_4_185/a_124_375# 0 0.246306f
C20686 FILLER_0_4_152/a_36_472# 0 0.417394f
C20687 FILLER_0_4_152/a_124_375# 0 0.246306f
C20688 _291_/a_36_160# 0 0.386641f
C20689 ctln[2] 0 1.833091f
C20690 output9/a_224_472# 0 2.38465f
C20691 ctln[4] 0 1.461847f
C20692 output11/a_224_472# 0 2.38465f
C20693 trimb[1] 0 0.378532f
C20694 output44/a_224_472# 0 2.38465f
C20695 result[6] 0 0.19512f
C20696 output33/a_224_472# 0 2.38465f
C20697 ctlp[5] 0 1.282822f
C20698 output22/a_224_472# 0 2.38465f
C20699 FILLER_0_8_127/a_36_472# 0 0.417394f
C20700 FILLER_0_8_127/a_124_375# 0 0.246306f
C20701 FILLER_0_8_138/a_36_472# 0 0.417394f
C20702 FILLER_0_8_138/a_124_375# 0 0.246306f
C20703 FILLER_0_21_133/a_36_472# 0 0.417394f
C20704 FILLER_0_21_133/a_124_375# 0 0.246306f
C20705 FILLER_0_24_130/a_36_472# 0 0.417394f
C20706 FILLER_0_24_130/a_124_375# 0 0.246306f
C20707 FILLER_0_18_171/a_36_472# 0 0.417394f
C20708 FILLER_0_18_171/a_124_375# 0 0.246306f
C20709 _258_/a_36_160# 0 0.386641f
C20710 _016_ 0 0.314121f
C20711 _327_/a_36_472# 0 0.031137f
C20712 _189_/a_67_603# 0 0.345683f
C20713 FILLER_0_24_63/a_36_472# 0 0.417394f
C20714 FILLER_0_24_63/a_124_375# 0 0.246306f
C20715 FILLER_0_24_96/a_36_472# 0 0.417394f
C20716 FILLER_0_24_96/a_124_375# 0 0.246306f
C20717 cal_itt\[2\] 0 1.473514f
C20718 _002_ 0 0.289553f
C20719 _413_/a_2560_156# 0 0.016968f
C20720 _413_/a_2665_112# 0 0.62251f
C20721 _413_/a_2248_156# 0 0.371662f
C20722 _413_/a_1204_472# 0 0.012971f
C20723 _413_/a_1000_472# 0 0.291735f
C20724 _413_/a_796_472# 0 0.023206f
C20725 _413_/a_1308_423# 0 0.279043f
C20726 _413_/a_448_472# 0 0.684413f
C20727 _413_/a_36_151# 0 1.43589f
C20728 _092_ 0 0.680239f
C20729 FILLER_0_7_72/a_3172_472# 0 0.345058f
C20730 FILLER_0_7_72/a_2724_472# 0 0.33241f
C20731 FILLER_0_7_72/a_2276_472# 0 0.33241f
C20732 FILLER_0_7_72/a_1828_472# 0 0.33241f
C20733 FILLER_0_7_72/a_1380_472# 0 0.33241f
C20734 FILLER_0_7_72/a_932_472# 0 0.33241f
C20735 FILLER_0_7_72/a_484_472# 0 0.33241f
C20736 FILLER_0_7_72/a_36_472# 0 0.404746f
C20737 FILLER_0_7_72/a_3260_375# 0 0.233093f
C20738 FILLER_0_7_72/a_2812_375# 0 0.17167f
C20739 FILLER_0_7_72/a_2364_375# 0 0.17167f
C20740 FILLER_0_7_72/a_1916_375# 0 0.17167f
C20741 FILLER_0_7_72/a_1468_375# 0 0.17167f
C20742 FILLER_0_7_72/a_1020_375# 0 0.17167f
C20743 FILLER_0_7_72/a_572_375# 0 0.17167f
C20744 FILLER_0_7_72/a_124_375# 0 0.185915f
C20745 _086_ 0 2.45259f
C20746 _119_ 0 1.237181f
C20747 net63 0 5.362473f
C20748 _430_/a_2560_156# 0 0.016968f
C20749 _430_/a_2665_112# 0 0.62251f
C20750 _430_/a_2248_156# 0 0.371662f
C20751 _430_/a_1204_472# 0 0.012971f
C20752 _430_/a_1000_472# 0 0.291735f
C20753 _430_/a_796_472# 0 0.023206f
C20754 _430_/a_1308_423# 0 0.279043f
C20755 _430_/a_448_472# 0 0.684413f
C20756 _430_/a_36_151# 0 1.43589f
C20757 _292_/a_36_160# 0 0.386641f
C20758 comp 0 1.022965f
C20759 ctln[1] 0 1.11973f
C20760 output8/a_224_472# 0 2.38465f
C20761 ctln[3] 0 0.835391f
C20762 output10/a_224_472# 0 2.38465f
C20763 result[5] 0 0.206867f
C20764 net32 0 1.78884f
C20765 output32/a_224_472# 0 2.38465f
C20766 trimb[0] 0 0.847787f
C20767 output43/a_224_472# 0 2.38465f
C20768 ctlp[4] 0 0.37565f
C20769 output21/a_224_472# 0 2.38465f
C20770 _053_ 0 1.705161f
C20771 FILLER_0_16_107/a_484_472# 0 0.345058f
C20772 FILLER_0_16_107/a_36_472# 0 0.404746f
C20773 FILLER_0_16_107/a_572_375# 0 0.232991f
C20774 FILLER_0_16_107/a_124_375# 0 0.185089f
C20775 FILLER_0_3_204/a_36_472# 0 0.417394f
C20776 FILLER_0_3_204/a_124_375# 0 0.246306f
C20777 FILLER_0_9_28/a_3172_472# 0 0.345058f
C20778 FILLER_0_9_28/a_2724_472# 0 0.33241f
C20779 FILLER_0_9_28/a_2276_472# 0 0.33241f
C20780 FILLER_0_9_28/a_1828_472# 0 0.33241f
C20781 FILLER_0_9_28/a_1380_472# 0 0.33241f
C20782 FILLER_0_9_28/a_932_472# 0 0.33241f
C20783 FILLER_0_9_28/a_484_472# 0 0.33241f
C20784 FILLER_0_9_28/a_36_472# 0 0.404746f
C20785 FILLER_0_9_28/a_3260_375# 0 0.233093f
C20786 FILLER_0_9_28/a_2812_375# 0 0.17167f
C20787 FILLER_0_9_28/a_2364_375# 0 0.17167f
C20788 FILLER_0_9_28/a_1916_375# 0 0.17167f
C20789 FILLER_0_9_28/a_1468_375# 0 0.17167f
C20790 FILLER_0_9_28/a_1020_375# 0 0.17167f
C20791 FILLER_0_9_28/a_572_375# 0 0.17167f
C20792 FILLER_0_9_28/a_124_375# 0 0.185915f
C20793 _132_ 0 1.491425f
C20794 _328_/a_36_113# 0 0.418095f
C20795 _414_/a_2560_156# 0 0.016968f
C20796 _414_/a_2665_112# 0 0.62251f
C20797 _414_/a_2248_156# 0 0.371662f
C20798 _414_/a_1204_472# 0 0.012971f
C20799 _414_/a_1000_472# 0 0.291735f
C20800 _414_/a_796_472# 0 0.023206f
C20801 _414_/a_1308_423# 0 0.279043f
C20802 _414_/a_448_472# 0 0.684413f
C20803 _414_/a_36_151# 0 1.43589f
C20804 _276_/a_36_160# 0 0.386641f
C20805 _144_ 0 1.173846f
C20806 _345_/a_36_160# 0 0.386641f
C20807 _155_ 0 0.638535f
C20808 _020_ 0 0.316793f
C20809 _431_/a_2560_156# 0 0.016968f
C20810 _431_/a_2665_112# 0 0.62251f
C20811 _431_/a_2248_156# 0 0.371662f
C20812 _431_/a_1204_472# 0 0.012971f
C20813 _431_/a_1000_472# 0 0.291735f
C20814 _431_/a_796_472# 0 0.023206f
C20815 _431_/a_1308_423# 0 0.279043f
C20816 _431_/a_448_472# 0 0.684413f
C20817 _431_/a_36_151# 0 1.43589f
C20818 _105_ 0 1.21281f
C20819 _293_/a_36_472# 0 0.031137f
C20820 FILLER_0_5_128/a_484_472# 0 0.345058f
C20821 FILLER_0_5_128/a_36_472# 0 0.404746f
C20822 FILLER_0_5_128/a_572_375# 0 0.232991f
C20823 FILLER_0_5_128/a_124_375# 0 0.185089f
C20824 FILLER_0_5_117/a_36_472# 0 0.417394f
C20825 FILLER_0_5_117/a_124_375# 0 0.246306f
C20826 ctln[0] 0 1.423102f
C20827 net7 0 1.174913f
C20828 output7/a_224_472# 0 2.38465f
C20829 trim[4] 0 0.763069f
C20830 output42/a_224_472# 0 2.38465f
C20831 result[4] 0 0.038878f
C20832 net31 0 1.912935f
C20833 output31/a_224_472# 0 2.38465f
C20834 ctlp[3] 0 1.14968f
C20835 output20/a_224_472# 0 2.38465f
C20836 FILLER_0_16_73/a_484_472# 0 0.345058f
C20837 FILLER_0_16_73/a_36_472# 0 0.404746f
C20838 FILLER_0_16_73/a_572_375# 0 0.232991f
C20839 FILLER_0_16_73/a_124_375# 0 0.185089f
C20840 FILLER_0_21_142/a_484_472# 0 0.345058f
C20841 FILLER_0_21_142/a_36_472# 0 0.404746f
C20842 FILLER_0_21_142/a_572_375# 0 0.232991f
C20843 FILLER_0_21_142/a_124_375# 0 0.185089f
C20844 FILLER_0_15_150/a_36_472# 0 0.417394f
C20845 FILLER_0_15_150/a_124_375# 0 0.246306f
C20846 FILLER_0_19_125/a_36_472# 0 0.417394f
C20847 FILLER_0_19_125/a_124_375# 0 0.246306f
C20848 net10 0 1.480101f
C20849 net20 0 2.034189f
C20850 _277_/a_36_160# 0 0.386641f
C20851 net27 0 2.023744f
C20852 _004_ 0 0.390107f
C20853 _415_/a_2560_156# 0 0.016968f
C20854 _415_/a_2665_112# 0 0.62251f
C20855 _415_/a_2248_156# 0 0.371662f
C20856 _415_/a_1204_472# 0 0.012971f
C20857 _415_/a_1000_472# 0 0.291735f
C20858 _415_/a_796_472# 0 0.023206f
C20859 _415_/a_1308_423# 0 0.279043f
C20860 _415_/a_448_472# 0 0.684413f
C20861 _415_/a_36_151# 0 1.43589f
C20862 mask\[5\] 0 1.334568f
C20863 _346_/a_49_472# 0 0.054843f
C20864 _028_ 0 0.386029f
C20865 _363_/a_36_68# 0 0.150048f
C20866 _021_ 0 0.316776f
C20867 _432_/a_2560_156# 0 0.016968f
C20868 _432_/a_2665_112# 0 0.62251f
C20869 _432_/a_2248_156# 0 0.371662f
C20870 _432_/a_1204_472# 0 0.012971f
C20871 _432_/a_1000_472# 0 0.291735f
C20872 _432_/a_796_472# 0 0.023206f
C20873 _432_/a_1308_423# 0 0.279043f
C20874 _432_/a_448_472# 0 0.684413f
C20875 _432_/a_36_151# 0 1.43589f
C20876 _008_ 0 0.423631f
C20877 _104_ 0 1.435764f
C20878 _106_ 0 0.378703f
C20879 FILLER_0_17_200/a_484_472# 0 0.345058f
C20880 FILLER_0_17_200/a_36_472# 0 0.404746f
C20881 FILLER_0_17_200/a_572_375# 0 0.232991f
C20882 FILLER_0_17_200/a_124_375# 0 0.185089f
.ends

.subckt saradc trim3 trim2 trim0 trim1 trim4 trimb3 trimb2 trimb0 trimb1 trimb4 cmp_outn
+ cmp_outp cmp_vinn cmp_vinp vss ctlp2 ctlp1 ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9
+ ctlp0 vdd ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctln8 ctln9 ctln0 cmp_clkc sample
+ vinn rstn clk en cal valid vinp result0 result1 result2 result3 result4 result5
+ result6 result7 result8 result9
Xlatch_0 latch_0/Qn vdd cmp_outp cmp_outn latch_0/XM3$5_0/a_n211_n1582# latch_0/x3_0/out
+ latch_0/x4_0/out latch_0/XM4$5_0/a_540_n1607# vss latch
Xbuffer_0 buffer_0/in cmp_clkc buffer_0/inv$2_1/in vdd vss buffer
Xdacp_0 ctlp0 vinp vdd ctlp2 ctlp1 ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9 cmp_vinp
+ dacp_0/ndum dacp_0/n1 dacp_0/n2 dacp_0/n3 dacp_0/n4 dacp_0/n5 dacp_0/n6 dacp_0/n7
+ dacp_0/n8 dacp_0/n9 sample dacp_0/bootstrapped_sw_0/vbsl dacp_0/bootstrapped_sw_0/vbsh
+ dacp_0/n0 vdd vss dacp
Xdacn_0 vinn vdd ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctln8 ctln9 ctln0 cmp_vinn
+ dacn_0/ndum dacn_0/n1 dacn_0/n2 dacn_0/n3 dacn_0/n4 dacn_0/n5 dacn_0/n6 dacn_0/n7
+ dacn_0/n8 dacn_0/n9 dacn_0/n0 sample vdd dacn_0/bootstrapped_sw$1_0/vbsl dacn_0/bootstrapped_sw$1_0/vbsh
+ vss dacn
Xcomparator_0 vdd cmp_vinp cmp_vinn trimb0 comparator_0/diff comparator_0/ip comparator_0/trimb_0/n3
+ cmp_outn cmp_clkc trim4 cmp_outp trim3 trim2 comparator_0/trim_0/n3 trim1 trim0
+ comparator_0/in trimb4 comparator_0/trim_0/n4 trimb3 comparator_0/trimb_0/n2 comparator_0/trim_0/n2
+ trimb2 comparator_0/trimb_0/n4 vss trimb1 comparator
Xmim_cap_boss_0 vss vdd vss mim_cap_boss
Xmim_cap_boss_1 vss vdd vss mim_cap_boss
Xsarlogic_0 ctln0 ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln8 ctlp0 ctlp1 ctlp2 ctlp3
+ ctlp4 ctlp5 ctlp6 ctlp7 ctlp8 ctlp9 cal clk buffer_0/in vdd en result0 result1 result2
+ result3 result4 result5 result6 result7 result8 result9 rstn sample trim0 trim1
+ trim2 trim3 trim4 trimb0 trimb1 trimb2 trimb3 trimb4 valid sarlogic_0/output13/a_224_472#
+ sarlogic_0/output23/a_224_472# sarlogic_0/net27 sarlogic_0/output25/a_224_472# sarlogic_0/cal_itt\[1\]
+ ctln7 sarlogic_0/net15 sarlogic_0/net59 ctln9 sarlogic_0/output10/a_224_472# sarlogic_0/net24
+ sarlogic_0/output11/a_224_472# sarlogic_0/output21/a_224_472# sarlogic_0/net14 sarlogic_0/output12/a_224_472#
+ sarlogic_0/output22/a_224_472# vdd sarlogic_0/net62 sarlogic_0/net20 vss sarlogic
C0 cmp_outn buffer_0/inv$2_1/in 0.010101f
C1 cmp_vinn dacn_0/n7 0.210031p
C2 dacp_0/n6 dacp_0/n1 0.134562f
C3 trimb3 vdd 0.303807f
C4 ctln3 ctln2 4.188161f
C5 result0 vdd 7.663611f
C6 result8 vdd 8.332389f
C7 result8 result9 6.071793f
C8 ctln2 vdd 0.50039f
C9 dacn_0/n9 dacn_0/n7 29.516087f
C10 comparator_0/trim_0/n3 vdd 0.160823f
C11 sample result2 0.160984f
C12 dacn_0/n2 dacn_0/n8 0.770114f
C13 sample vdd 2.339275f
C14 sarlogic_0/output12/a_224_472# vdd 0.004511f
C15 sample result9 0.161326f
C16 dacn_0/n1 cmp_vinn 3.365905f
C17 dacp_0/n6 dacp_0/n3 0.336612f
C18 cmp_vinp dacp_0/n6 0.105055p
C19 dacp_0/n6 dacp_0/n8 11.2161f
C20 ctlp1 vdd 0.803166f
C21 comparator_0/ip comparator_0/trimb_0/n3 6.42492f
C22 dacn_0/n0 dacn_0/n6 0.025424f
C23 dacp_0/n6 dacp_0/n2 0.207877f
C24 trimb0 vdd 0.066096f
C25 cal sample 0.161292f
C26 dacp_0/n6 dacp_0/n0 0.025424f
C27 dacn_0/n1 dacn_0/n9 0.342393f
C28 ctlp8 vdd 0.232138f
C29 dacn_0/n4 dacn_0/n7 1.70387f
C30 dacp_0/n6 dacp_0/n5 28.589401f
C31 ctlp6 ctlp5 3.405441f
C32 comparator_0/trim_0/n0 comparator_0/trim_0/n1 0.032158f
C33 comparator_0/in comparator_0/trim_0/n1 1.60623f
C34 result7 vdd 7.905001f
C35 comparator_0/in vdd 0.276627f
C36 dacp_0/n7 dacp_0/n1 0.205173f
C37 dacn_0/n2 dacn_0/n5 0.207999f
C38 dacn_0/n2 dacn_0/ndum 0.041162f
C39 dacn_0/n1 dacn_0/n4 0.134826f
C40 ctlp3 ctlp4 3.92725f
C41 dacn_0/n6 cmp_vinn 0.105055p
C42 cmp_clkc cmp_outn 0.134865f
C43 dacp_0/n9 dacp_0/n1 0.342393f
C44 cmp_vinp dacp_0/n7 0.210031p
C45 dacp_0/n7 dacp_0/n3 0.891504f
C46 dacp_0/n8 dacp_0/n7 50.178104f
C47 dacn_0/n6 dacn_0/n9 14.716789f
C48 comparator_0/trimb_0/n1 comparator_0/trimb_0/n0 0.032158f
C49 dacp_0/n7 dacp_0/n2 0.485242f
C50 en vdd 7.929791f
C51 dacp_0/n7 dacp_0/n0 0.06073f
C52 dacn_0/n1 dacn_0/n7 0.205173f
C53 comparator_0/trimb_0/n2 vdd 0.035873f
C54 dacn_0/n0 dacn_0/n2 0.099202f
C55 dacp_0/n5 dacp_0/n7 3.36878f
C56 cmp_vinp dacp_0/n9 0.846155p
C57 cal en 6.091991f
C58 dacp_0/n9 dacp_0/n3 1.911224f
C59 dacp_0/n9 dacp_0/n8 87.10268f
C60 vdd rstn 9.38116f
C61 dacn_0/n8 dacn_0/n3 1.46111f
C62 ctlp1 ctlp2 4.44906f
C63 dacp_0/n9 dacp_0/n2 0.996568f
C64 result6 vdd 7.645501f
C65 dacp_0/n9 dacp_0/n0 0.184985f
C66 dacn_0/n4 dacn_0/n6 0.614078f
C67 trimb4 trimb1 2.933839f
C68 ctlp9 ctlp0 2.368197f
C69 ctln5 vdd 1.126741f
C70 dacp_0/n9 dacp_0/n5 7.399346f
C71 comparator_0/trim_0/n2 comparator_0/in 3.21246f
C72 comparator_0/trim_0/n4 comparator_0/trim_0/n1 0.032158f
C73 comparator_0/trim_0/n4 vdd 0.050918f
C74 dacp_0/n6 dacp_0/ndum 0.025424f
C75 ctlp3 vdd 0.357376f
C76 dacn_0/n6 dacn_0/n7 34.326103f
C77 comparator_0/ip comparator_0/trimb_0/n4 12.849839f
C78 trimb1 vdd 0.066886f
C79 result0 valid 2.38317f
C80 dacn_0/n2 cmp_vinn 6.640605f
C81 result4 vdd 7.126491f
C82 sarlogic_0/net20 vdd 0.003406f
C83 ctlp6 ctlp7 3.144531f
C84 ctln1 vdd 0.810505f
C85 sample clk 0.18099f
C86 ctlp4 vdd 0.688795f
C87 dacn_0/n5 dacn_0/n3 0.346757f
C88 dacn_0/ndum dacn_0/n3 0.025424f
C89 ctln0 trim3 0.097876f
C90 sample sarlogic_0/fanout65/a_36_113# 0.001365f
C91 sample valid 0.161748f
C92 dacn_0/n2 dacn_0/n9 0.996568f
C93 latch_0/XM4$5_0/a_540_n1607# vdd 0.002382f
C94 trim3 vdd 0.303807f
C95 dacn_0/n1 dacn_0/n6 0.134562f
C96 cmp_outp vdd 0.061575f
C97 trim0 vdd 0.066096f
C98 trimb3 ctlp0 0.087957f
C99 dacn_0/n2 dacn_0/n4 0.213096f
C100 dacn_0/n0 dacn_0/n3 0.051666f
C101 dacp_0/n7 dacp_0/ndum 0.06073f
C102 trimb4 vdd 0.098486f
C103 trimb3 trimb2 2.951539f
C104 comparator_0/trim_0/n2 comparator_0/trim_0/n4 0.128631f
C105 sample sarlogic_0/net27 0.004307f
C106 ctln0 vdd 0.206198f
C107 ctln7 vdd 0.374489f
C108 result2 vdd 6.553131f
C109 dacn_0/n2 dacn_0/n7 0.485242f
C110 dacp_0/n9 dacp_0/ndum 0.127951f
C111 ctln3 vdd 0.357376f
C112 sample sarlogic_0/net62 0.20203f
C113 ctlp3 ctlp2 4.188161f
C114 en clk 6.086483f
C115 result9 vdd 9.36568f
C116 ctln9 ctln0 2.368197f
C117 cal vdd 7.670291f
C118 trimb0 trimb2 3.097479f
C119 dacn_0/n3 cmp_vinn 13.201303f
C120 clk rstn 6.080953f
C121 ctln9 vdd 0.334729f
C122 cmp_outp latch_0/x4_0/out 0.005228f
C123 dacn_0/n2 dacn_0/n1 16.597801f
C124 dacn_0/n3 dacn_0/n9 1.911224f
C125 dacp_0/n4 dacp_0/n1 0.134826f
C126 cmp_outp latch_0/Qn 0.002019f
C127 dacp_0/n6 dacp_0/n7 34.326103f
C128 sample result3 0.160929f
C129 dacn_0/n8 dacn_0/n5 5.60732f
C130 dacn_0/n8 dacn_0/ndum 0.097254f
C131 dacp_0/n4 dacp_0/n3 25.8929f
C132 cmp_vinp dacp_0/n4 26.32268f
C133 cmp_clkc comparator_0/in 0.016561f
C134 dacp_0/n4 dacp_0/n8 2.84323f
C135 dacp_0/n6 dacp_0/n9 14.716789f
C136 dacn_0/n4 dacn_0/n3 25.8929f
C137 dacp_0/n4 dacp_0/n2 0.213096f
C138 latch_0/x4_0/out vdd 0.002021f
C139 dacp_0/n4 dacp_0/n0 0.040502f
C140 dacn_0/n2 dacn_0/n6 0.207877f
C141 comparator_0/trimb_0/n2 comparator_0/trimb_0/n4 0.128631f
C142 comparator_0/trim_0/n2 vdd 0.035873f
C143 comparator_0/trimb_0/n3 vdd 0.160824f
C144 comparator_0/trimb_0/n4 comparator_0/trimb_0/n0 0.032158f
C145 dacp_0/n4 dacp_0/n5 27.491999f
C146 ctlp2 vdd 0.54584f
C147 latch_0/Qn vdd 0.059458f
C148 dacn_0/n3 dacn_0/n7 0.891504f
C149 dacn_0/n0 dacn_0/n8 0.097254f
C150 cmp_vinp vdd 0.257757f
C151 ctlp8 ctlp9 2.62272f
C152 result5 sample 0.160929f
C153 sample sarlogic_0/cal_itt\[1\] 0.004307f
C154 dacn_0/ndum dacn_0/n5 0.025424f
C155 ctlp8 ctlp7 2.88363f
C156 ctln7 ctln8 2.88363f
C157 result0 result1 6.064423f
C158 buffer_0/in vdd 0.287466f
C159 ctln8 vdd 0.232138f
C160 ctlp4 ctlp5 3.66635f
C161 vinp vdd 12.3187f
C162 dacn_0/n1 dacn_0/n3 0.137399f
C163 sample result1 0.160984f
C164 dacp_0/n9 dacp_0/n7 29.516087f
C165 vdd sarlogic_0/net14 0.003601f
C166 ctln9 ctln8 2.62272f
C167 latch_0/x3_0/out vdd 0.084411f
C168 dacp_0/bootstrapped_sw_0/vbsl vinp 0.012179f
C169 clk vdd 8.18937f
C170 cmp_vinn vdd 0.257757f
C171 trim0 trim1 2.987179f
C172 dacn_0/n8 cmp_vinn 0.420151p
C173 ctln4 ctln5 3.66635f
C174 dacn_0/n0 dacn_0/n5 0.025424f
C175 sample result0 0.161748f
C176 sample result8 0.161003f
C177 cmp_outn cmp_outp 0.235348f
C178 valid vdd 8.159651f
C179 buffer_0/inv$2_1/in vdd 0.071983f
C180 trim2 trim3 2.959509f
C181 trim4 vdd 0.100841f
C182 dacn_0/n8 dacn_0/n9 87.10268f
C183 ctln6 ctln5 3.405441f
C184 cal valid 6.097543f
C185 dacp_0/n1 dacp_0/n3 0.137399f
C186 cmp_vinp dacp_0/n1 3.365905f
C187 dacp_0/n8 dacp_0/n1 0.278221f
C188 trim2 trim0 3.097479f
C189 dacn_0/n6 dacn_0/n3 0.336612f
C190 dacp_0/n2 dacp_0/n1 16.597801f
C191 comparator_0/ip comparator_0/trimb_0/n2 3.21246f
C192 sarlogic_0/output10/a_224_472# vdd 0.004573f
C193 dacp_0/n0 dacp_0/n1 8.469266f
C194 comparator_0/ip comparator_0/trimb_0/n0 1.60623f
C195 trim1 vdd 0.064237f
C196 dacp_0/n4 dacp_0/ndum 0.025424f
C197 result7 result8 6.077323f
C198 result4 result3 6.099443f
C199 ctlp5 vdd 1.126741f
C200 sarlogic_0/net24 vdd 0.003517f
C201 comparator_0/trimb_0/n1 comparator_0/trimb_0/n4 0.032158f
C202 dacn_0/n5 cmp_vinn 52.565514f
C203 dacn_0/n8 dacn_0/n4 2.84323f
C204 dacn_0/ndum cmp_vinn 1.640173f
C205 dacp_0/n5 dacp_0/n1 0.134705f
C206 cmp_vinp dacp_0/n3 13.201303f
C207 cmp_vinp dacp_0/n8 0.420151p
C208 ctlp0 vdd 0.206198f
C209 dacp_0/n8 dacp_0/n3 1.46111f
C210 comparator_0/in comparator_0/trim_0/n3 6.42492f
C211 result5 result6 6.088384f
C212 cmp_outn vdd 0.208f
C213 cmp_vinp dacp_0/n2 6.640605f
C214 dacp_0/n2 dacp_0/n3 22.8406f
C215 result7 sample 0.161003f
C216 dacp_0/n8 dacp_0/n2 0.770114f
C217 cmp_vinp dacp_0/n0 1.702731f
C218 dacp_0/n0 dacp_0/n3 0.051666f
C219 comparator_0/trimb_0/n4 vdd 0.050918f
C220 dacp_0/n8 dacp_0/n0 0.097254f
C221 dacn_0/n5 dacn_0/n9 7.399346f
C222 dacn_0/ndum dacn_0/n9 0.127951f
C223 dacp_0/n0 dacp_0/n2 0.099202f
C224 trim2 vdd 0.092754f
C225 dacn_0/n8 dacn_0/n7 50.178104f
C226 cmp_vinp dacp_0/n5 52.565514f
C227 dacp_0/n5 dacp_0/n3 0.346757f
C228 dacp_0/n5 dacp_0/n8 5.60732f
C229 trimb2 vdd 0.090104f
C230 dacp_0/n5 dacp_0/n2 0.207999f
C231 ctlp6 vdd 0.849567f
C232 dacp_0/n5 dacp_0/n0 0.025424f
C233 dacn_0/n0 cmp_vinn 1.702731f
C234 result5 result4 6.093913f
C235 comparator_0/in comparator_0/trim_0/n0 1.60623f
C236 dacn_0/n5 dacn_0/n4 27.491999f
C237 cmp_clkc vdd 0.060231f
C238 dacn_0/ndum dacn_0/n4 0.025424f
C239 ctln4 ctln3 3.92725f
C240 sample en 0.185896f
C241 dacn_0/n8 dacn_0/n1 0.278221f
C242 ctln4 vdd 0.687612f
C243 dacn_0/n2 dacn_0/n3 22.8406f
C244 dacn_0/n0 dacn_0/n9 0.184985f
C245 dacp_0/n4 dacp_0/n6 0.614078f
C246 ctln6 ctln7 3.144531f
C247 sample rstn 0.161326f
C248 result2 result3 6.064423f
C249 vinn dacn_0/bootstrapped_sw$1_0/vbsl 0.01281f
C250 buffer_0/in buffer_0/inv$2_1/in 0.003647f
C251 sample result6 0.161003f
C252 ctln6 vdd 0.849567f
C253 vdd result3 6.868131f
C254 dacn_0/n5 dacn_0/n7 3.36878f
C255 dacn_0/ndum dacn_0/n7 0.06073f
C256 sample sarlogic_0/net59 0.043318f
C257 comparator_0/trim_0/n3 comparator_0/trim_0/n4 0.241184f
C258 dacn_0/n0 dacn_0/n4 0.040502f
C259 comparator_0/ip comparator_0/trimb_0/n1 1.60623f
C260 comparator_0/trimb_0/n3 comparator_0/trimb_0/n4 0.241184f
C261 ctln2 ctln1 4.44906f
C262 dacp_0/ndum dacp_0/n1 8.161697f
C263 ctlp9 vdd 0.38096f
C264 ctlp7 vdd 0.368909f
C265 dacn_0/n5 dacn_0/n1 0.134705f
C266 dacn_0/ndum dacn_0/n1 8.161697f
C267 dacn_0/n8 dacn_0/n6 11.2161f
C268 dacn_0/n9 cmp_vinn 0.846155p
C269 result7 result6 6.082853f
C270 result4 sample 0.160929f
C271 comparator_0/ip vdd 0.276626f
C272 trimb0 trimb1 2.995159f
C273 dacn_0/n0 dacn_0/n7 0.06073f
C274 sarlogic_0/output22/a_224_472# vdd 0.004694f
C275 dacp_0/n4 dacp_0/n7 1.70387f
C276 cmp_vinp dacp_0/ndum 1.640173f
C277 result5 vdd 7.386001f
C278 dacp_0/ndum dacp_0/n3 0.025424f
C279 dacp_0/n8 dacp_0/ndum 0.097254f
C280 dacp_0/ndum dacp_0/n2 0.041162f
C281 comparator_0/trim_0/n4 comparator_0/trim_0/n0 0.032158f
C282 comparator_0/in comparator_0/trim_0/n4 12.849839f
C283 dacn_0/n4 cmp_vinn 26.32268f
C284 cmp_outn latch_0/x3_0/out 0.004541f
C285 result1 result2 6.299723f
C286 trim4 trim1 2.925859f
C287 dacp_0/n4 dacp_0/n9 3.740573f
C288 dacn_0/n0 dacn_0/n1 8.469266f
C289 dacp_0/n5 dacp_0/ndum 0.025424f
C290 result1 vdd 6.582241f
C291 vinn vdd 12.3187f
C292 dacn_0/n5 dacn_0/n6 28.589401f
C293 dacn_0/ndum dacn_0/n6 0.025424f
C294 dacn_0/n4 dacn_0/n9 3.740573f
C295 sarlogic_0/_034_ vss 0.304805f
C296 sarlogic_0/_160_ vss 1.542665f
C297 sarlogic_0/_166_ vss 0.299751f
C298 sarlogic_0/output41/a_224_472# vss 2.38465f
C299 sarlogic_0/net6 vss 1.112469f
C300 sarlogic_0/output6/a_224_472# vss 2.38465f
C301 sarlogic_0/FILLER_0_12_196/a_36_472# vss 0.417394f
C302 sarlogic_0/FILLER_0_12_196/a_124_375# vss 0.246306f
C303 result3 vss 16.620413f
C304 sarlogic_0/net30 vss 1.81422f
C305 sarlogic_0/output30/a_224_472# vss 2.38465f
C306 sarlogic_0/_047_ vss 0.374694f
C307 sarlogic_0/_201_/a_67_603# vss 0.345683f
C308 sarlogic_0/_416_/a_2560_156# vss 0.016968f
C309 sarlogic_0/_416_/a_2665_112# vss 0.62251f
C310 sarlogic_0/_416_/a_2248_156# vss 0.371662f
C311 sarlogic_0/_416_/a_1204_472# vss 0.012971f
C312 sarlogic_0/_416_/a_1000_472# vss 0.291735f
C313 sarlogic_0/_416_/a_796_472# vss 0.023206f
C314 sarlogic_0/_416_/a_1308_423# vss 0.279043f
C315 sarlogic_0/_416_/a_448_472# vss 0.684413f
C316 sarlogic_0/_416_/a_36_151# vss 1.43589f
C317 sarlogic_0/FILLER_0_13_290/a_36_472# vss 0.417394f
C318 sarlogic_0/FILLER_0_13_290/a_124_375# vss 0.246306f
C319 sarlogic_0/_278_/a_36_160# vss 0.696445f
C320 sarlogic_0/_145_ vss 0.546455f
C321 sarlogic_0/FILLER_0_13_72/a_484_472# vss 0.345058f
C322 sarlogic_0/FILLER_0_13_72/a_36_472# vss 0.404746f
C323 sarlogic_0/FILLER_0_13_72/a_572_375# vss 0.232991f
C324 sarlogic_0/FILLER_0_13_72/a_124_375# vss 0.185089f
C325 sarlogic_0/FILLER_0_14_235/a_484_472# vss 0.345058f
C326 sarlogic_0/FILLER_0_14_235/a_36_472# vss 0.404746f
C327 sarlogic_0/FILLER_0_14_235/a_572_375# vss 0.232991f
C328 sarlogic_0/FILLER_0_14_235/a_124_375# vss 0.185089f
C329 sarlogic_0/_156_ vss 0.593796f
C330 sarlogic_0/_107_ vss 0.391583f
C331 sarlogic_0/_295_/a_36_472# vss 0.031137f
C332 sarlogic_0/_022_ vss 0.387773f
C333 sarlogic_0/_433_/a_2560_156# vss 0.016968f
C334 sarlogic_0/_433_/a_2665_112# vss 0.62251f
C335 sarlogic_0/_433_/a_2248_156# vss 0.371662f
C336 sarlogic_0/_433_/a_1204_472# vss 0.012971f
C337 sarlogic_0/_433_/a_1000_472# vss 0.291735f
C338 sarlogic_0/_433_/a_796_472# vss 0.023206f
C339 sarlogic_0/_433_/a_1308_423# vss 0.279043f
C340 sarlogic_0/_433_/a_448_472# vss 0.684413f
C341 sarlogic_0/_433_/a_36_151# vss 1.43589f
C342 sarlogic_0/FILLER_0_5_148/a_484_472# vss 0.345058f
C343 sarlogic_0/FILLER_0_5_148/a_36_472# vss 0.404746f
C344 sarlogic_0/FILLER_0_5_148/a_572_375# vss 0.232991f
C345 sarlogic_0/FILLER_0_5_148/a_124_375# vss 0.185089f
C346 sarlogic_0/_167_ vss 0.285904f
C347 sarlogic_0/_381_/a_36_472# vss 0.031137f
C348 sarlogic_0/net40 vss 1.845219f
C349 sarlogic_0/output40/a_224_472# vss 2.38465f
C350 sarlogic_0/cal_count\[0\] vss 0.893784f
C351 sarlogic_0/_039_ vss 0.412301f
C352 sarlogic_0/_450_/a_2449_156# vss 0.049992f
C353 sarlogic_0/_450_/a_2225_156# vss 0.434082f
C354 sarlogic_0/_450_/a_3129_107# vss 0.58406f
C355 sarlogic_0/_450_/a_836_156# vss 0.019766f
C356 sarlogic_0/_450_/a_1040_527# vss 0.302082f
C357 sarlogic_0/_450_/a_1353_112# vss 0.286513f
C358 sarlogic_0/_450_/a_448_472# vss 1.21246f
C359 sarlogic_0/_450_/a_36_151# vss 1.31409f
C360 rstn vss 26.841475f
C361 sarlogic_0/FILLER_0_8_156/a_484_472# vss 0.345058f
C362 sarlogic_0/FILLER_0_8_156/a_36_472# vss 0.404746f
C363 sarlogic_0/FILLER_0_8_156/a_572_375# vss 0.232991f
C364 sarlogic_0/FILLER_0_8_156/a_124_375# vss 0.185089f
C365 sarlogic_0/FILLER_0_6_37/a_36_472# vss 0.417394f
C366 sarlogic_0/FILLER_0_6_37/a_124_375# vss 0.246306f
C367 sarlogic_0/FILLER_0_21_60/a_484_472# vss 0.345058f
C368 sarlogic_0/FILLER_0_21_60/a_36_472# vss 0.404746f
C369 sarlogic_0/FILLER_0_21_60/a_572_375# vss 0.232991f
C370 sarlogic_0/FILLER_0_21_60/a_124_375# vss 0.185089f
C371 sarlogic_0/FILLER_0_22_107/a_484_472# vss 0.345058f
C372 sarlogic_0/FILLER_0_22_107/a_36_472# vss 0.404746f
C373 sarlogic_0/FILLER_0_22_107/a_572_375# vss 0.232991f
C374 sarlogic_0/FILLER_0_22_107/a_124_375# vss 0.185089f
C375 sarlogic_0/FILLER_0_16_115/a_36_472# vss 0.417394f
C376 sarlogic_0/FILLER_0_16_115/a_124_375# vss 0.246306f
C377 sarlogic_0/FILLER_0_19_134/a_36_472# vss 0.417394f
C378 sarlogic_0/FILLER_0_19_134/a_124_375# vss 0.246306f
C379 sarlogic_0/FILLER_0_3_212/a_36_472# vss 0.417394f
C380 sarlogic_0/FILLER_0_3_212/a_124_375# vss 0.246306f
C381 sarlogic_0/FILLER_0_10_94/a_484_472# vss 0.345058f
C382 sarlogic_0/FILLER_0_10_94/a_36_472# vss 0.404746f
C383 sarlogic_0/FILLER_0_10_94/a_572_375# vss 0.232991f
C384 sarlogic_0/FILLER_0_10_94/a_124_375# vss 0.185089f
C385 sarlogic_0/FILLER_0_4_91/a_484_472# vss 0.345058f
C386 sarlogic_0/FILLER_0_4_91/a_36_472# vss 0.404746f
C387 sarlogic_0/FILLER_0_4_91/a_572_375# vss 0.232991f
C388 sarlogic_0/FILLER_0_4_91/a_124_375# vss 0.185089f
C389 sarlogic_0/net14 vss 1.508711f
C390 sarlogic_0/_202_/a_36_160# vss 0.696445f
C391 sarlogic_0/FILLER_0_6_231/a_484_472# vss 0.345058f
C392 sarlogic_0/FILLER_0_6_231/a_36_472# vss 0.404746f
C393 sarlogic_0/FILLER_0_6_231/a_572_375# vss 0.232991f
C394 sarlogic_0/FILLER_0_6_231/a_124_375# vss 0.185089f
C395 vdd vss 9.660555p
C396 sarlogic_0/_006_ vss 0.41456f
C397 sarlogic_0/_417_/a_2560_156# vss 0.016968f
C398 sarlogic_0/_417_/a_2665_112# vss 0.62251f
C399 sarlogic_0/_417_/a_2248_156# vss 0.371662f
C400 sarlogic_0/_417_/a_1204_472# vss 0.012971f
C401 sarlogic_0/_417_/a_1000_472# vss 0.291735f
C402 sarlogic_0/_417_/a_796_472# vss 0.023206f
C403 sarlogic_0/_417_/a_1308_423# vss 0.279043f
C404 sarlogic_0/_417_/a_448_472# vss 0.684413f
C405 sarlogic_0/_417_/a_36_151# vss 1.43589f
C406 sarlogic_0/_146_ vss 0.35443f
C407 sarlogic_0/mask\[6\] vss 1.246962f
C408 sarlogic_0/_348_/a_49_472# vss 0.054843f
C409 sarlogic_0/_365_/a_36_68# vss 0.150048f
C410 sarlogic_0/_023_ vss 0.345812f
C411 sarlogic_0/_434_/a_2560_156# vss 0.016968f
C412 sarlogic_0/_434_/a_2665_112# vss 0.62251f
C413 sarlogic_0/_434_/a_2248_156# vss 0.371662f
C414 sarlogic_0/_434_/a_1204_472# vss 0.012971f
C415 sarlogic_0/_434_/a_1000_472# vss 0.291735f
C416 sarlogic_0/_434_/a_796_472# vss 0.023206f
C417 sarlogic_0/_434_/a_1308_423# vss 0.279043f
C418 sarlogic_0/_434_/a_448_472# vss 0.684413f
C419 sarlogic_0/_434_/a_36_151# vss 1.43589f
C420 sarlogic_0/FILLER_0_5_136/a_36_472# vss 0.417394f
C421 sarlogic_0/FILLER_0_5_136/a_124_375# vss 0.246306f
C422 sarlogic_0/FILLER_0_18_209/a_484_472# vss 0.345058f
C423 sarlogic_0/FILLER_0_18_209/a_36_472# vss 0.404746f
C424 sarlogic_0/FILLER_0_18_209/a_572_375# vss 0.232991f
C425 sarlogic_0/FILLER_0_18_209/a_124_375# vss 0.185089f
C426 sarlogic_0/FILLER_0_12_28/a_36_472# vss 0.417394f
C427 sarlogic_0/FILLER_0_12_28/a_124_375# vss 0.246306f
C428 sarlogic_0/_040_ vss 0.355703f
C429 sarlogic_0/_451_/a_2449_156# vss 0.049992f
C430 sarlogic_0/_451_/a_2225_156# vss 0.434082f
C431 sarlogic_0/_451_/a_3129_107# vss 0.58406f
C432 sarlogic_0/_451_/a_836_156# vss 0.019766f
C433 sarlogic_0/_451_/a_1040_527# vss 0.302082f
C434 sarlogic_0/_451_/a_1353_112# vss 0.286513f
C435 sarlogic_0/_451_/a_448_472# vss 1.21246f
C436 sarlogic_0/_451_/a_36_151# vss 1.31409f
C437 sarlogic_0/FILLER_0_6_47/a_3172_472# vss 0.345058f
C438 sarlogic_0/FILLER_0_6_47/a_2724_472# vss 0.33241f
C439 sarlogic_0/FILLER_0_6_47/a_2276_472# vss 0.33241f
C440 sarlogic_0/FILLER_0_6_47/a_1828_472# vss 0.33241f
C441 sarlogic_0/FILLER_0_6_47/a_1380_472# vss 0.33241f
C442 sarlogic_0/FILLER_0_6_47/a_932_472# vss 0.33241f
C443 sarlogic_0/FILLER_0_6_47/a_484_472# vss 0.33241f
C444 sarlogic_0/FILLER_0_6_47/a_36_472# vss 0.404746f
C445 sarlogic_0/FILLER_0_6_47/a_3260_375# vss 0.233093f
C446 sarlogic_0/FILLER_0_6_47/a_2812_375# vss 0.17167f
C447 sarlogic_0/FILLER_0_6_47/a_2364_375# vss 0.17167f
C448 sarlogic_0/FILLER_0_6_47/a_1916_375# vss 0.17167f
C449 sarlogic_0/FILLER_0_6_47/a_1468_375# vss 0.17167f
C450 sarlogic_0/FILLER_0_6_47/a_1020_375# vss 0.17167f
C451 sarlogic_0/FILLER_0_6_47/a_572_375# vss 0.17167f
C452 sarlogic_0/FILLER_0_6_47/a_124_375# vss 0.185915f
C453 sarlogic_0/FILLER_0_21_150/a_36_472# vss 0.417394f
C454 sarlogic_0/FILLER_0_21_150/a_124_375# vss 0.246306f
C455 sarlogic_0/FILLER_0_15_180/a_484_472# vss 0.345058f
C456 sarlogic_0/FILLER_0_15_180/a_36_472# vss 0.404746f
C457 sarlogic_0/FILLER_0_15_180/a_572_375# vss 0.232991f
C458 sarlogic_0/FILLER_0_15_180/a_124_375# vss 0.185089f
C459 sarlogic_0/FILLER_0_22_128/a_3172_472# vss 0.345058f
C460 sarlogic_0/FILLER_0_22_128/a_2724_472# vss 0.33241f
C461 sarlogic_0/FILLER_0_22_128/a_2276_472# vss 0.33241f
C462 sarlogic_0/FILLER_0_22_128/a_1828_472# vss 0.33241f
C463 sarlogic_0/FILLER_0_22_128/a_1380_472# vss 0.33241f
C464 sarlogic_0/FILLER_0_22_128/a_932_472# vss 0.33241f
C465 sarlogic_0/FILLER_0_22_128/a_484_472# vss 0.33241f
C466 sarlogic_0/FILLER_0_22_128/a_36_472# vss 0.404746f
C467 sarlogic_0/FILLER_0_22_128/a_3260_375# vss 0.233093f
C468 sarlogic_0/FILLER_0_22_128/a_2812_375# vss 0.17167f
C469 sarlogic_0/FILLER_0_22_128/a_2364_375# vss 0.17167f
C470 sarlogic_0/FILLER_0_22_128/a_1916_375# vss 0.17167f
C471 sarlogic_0/FILLER_0_22_128/a_1468_375# vss 0.17167f
C472 sarlogic_0/FILLER_0_22_128/a_1020_375# vss 0.17167f
C473 sarlogic_0/FILLER_0_22_128/a_572_375# vss 0.17167f
C474 sarlogic_0/FILLER_0_22_128/a_124_375# vss 0.185915f
C475 sarlogic_0/FILLER_0_19_111/a_484_472# vss 0.345058f
C476 sarlogic_0/FILLER_0_19_111/a_36_472# vss 0.404746f
C477 sarlogic_0/FILLER_0_19_111/a_572_375# vss 0.232991f
C478 sarlogic_0/FILLER_0_19_111/a_124_375# vss 0.185089f
C479 sarlogic_0/FILLER_0_19_155/a_484_472# vss 0.345058f
C480 sarlogic_0/FILLER_0_19_155/a_36_472# vss 0.404746f
C481 sarlogic_0/FILLER_0_19_155/a_572_375# vss 0.232991f
C482 sarlogic_0/FILLER_0_19_155/a_124_375# vss 0.185089f
C483 sarlogic_0/net11 vss 1.328455f
C484 sarlogic_0/net21 vss 1.922829f
C485 sarlogic_0/_007_ vss 0.309495f
C486 sarlogic_0/net77 vss 1.39077f
C487 sarlogic_0/_418_/a_2560_156# vss 0.016968f
C488 sarlogic_0/_418_/a_2665_112# vss 0.62251f
C489 sarlogic_0/_418_/a_2248_156# vss 0.371662f
C490 sarlogic_0/_418_/a_1204_472# vss 0.012971f
C491 sarlogic_0/_418_/a_1000_472# vss 0.291735f
C492 sarlogic_0/_418_/a_796_472# vss 0.023206f
C493 sarlogic_0/_418_/a_1308_423# vss 0.279043f
C494 sarlogic_0/_418_/a_448_472# vss 0.684413f
C495 sarlogic_0/_418_/a_36_151# vss 1.43589f
C496 sarlogic_0/_220_/a_67_603# vss 0.345683f
C497 sarlogic_0/FILLER_0_9_282/a_484_472# vss 0.345058f
C498 sarlogic_0/FILLER_0_9_282/a_36_472# vss 0.404746f
C499 sarlogic_0/FILLER_0_9_282/a_572_375# vss 0.232991f
C500 sarlogic_0/FILLER_0_9_282/a_124_375# vss 0.185089f
C501 sarlogic_0/FILLER_0_18_37/a_1380_472# vss 0.345058f
C502 sarlogic_0/FILLER_0_18_37/a_932_472# vss 0.33241f
C503 sarlogic_0/FILLER_0_18_37/a_484_472# vss 0.33241f
C504 sarlogic_0/FILLER_0_18_37/a_36_472# vss 0.404746f
C505 sarlogic_0/FILLER_0_18_37/a_1468_375# vss 0.233029f
C506 sarlogic_0/FILLER_0_18_37/a_1020_375# vss 0.171606f
C507 sarlogic_0/FILLER_0_18_37/a_572_375# vss 0.171606f
C508 sarlogic_0/FILLER_0_18_37/a_124_375# vss 0.185399f
C509 sarlogic_0/FILLER_0_2_127/a_36_472# vss 0.417394f
C510 sarlogic_0/FILLER_0_2_127/a_124_375# vss 0.246306f
C511 sarlogic_0/_157_ vss 0.531763f
C512 sarlogic_0/_435_/a_2560_156# vss 0.016968f
C513 sarlogic_0/_435_/a_2665_112# vss 0.62251f
C514 sarlogic_0/_435_/a_2248_156# vss 0.371662f
C515 sarlogic_0/_435_/a_1204_472# vss 0.012971f
C516 sarlogic_0/_435_/a_1000_472# vss 0.291735f
C517 sarlogic_0/_435_/a_796_472# vss 0.023206f
C518 sarlogic_0/_435_/a_1308_423# vss 0.279043f
C519 sarlogic_0/_435_/a_448_472# vss 0.684413f
C520 sarlogic_0/_435_/a_36_151# vss 1.43589f
C521 sarlogic_0/_108_ vss 0.411979f
C522 sarlogic_0/_297_/a_36_472# vss 0.031137f
C523 sarlogic_0/trim_mask\[3\] vss 1.081535f
C524 sarlogic_0/_164_ vss 1.3268f
C525 sarlogic_0/_383_/a_36_472# vss 0.031137f
C526 sarlogic_0/_041_ vss 0.299289f
C527 sarlogic_0/_452_/a_2449_156# vss 0.049992f
C528 sarlogic_0/_452_/a_2225_156# vss 0.434082f
C529 sarlogic_0/_452_/a_3129_107# vss 0.58406f
C530 sarlogic_0/_452_/a_836_156# vss 0.019766f
C531 sarlogic_0/_452_/a_1040_527# vss 0.302082f
C532 sarlogic_0/_452_/a_1353_112# vss 0.286513f
C533 sarlogic_0/_452_/a_448_472# vss 1.21246f
C534 sarlogic_0/_452_/a_36_151# vss 1.31409f
C535 sarlogic_0/FILLER_0_6_79/a_36_472# vss 0.417394f
C536 sarlogic_0/FILLER_0_6_79/a_124_375# vss 0.246306f
C537 sarlogic_0/net59 vss 5.044369f
C538 sarlogic_0/FILLER_0_15_59/a_484_472# vss 0.345058f
C539 sarlogic_0/FILLER_0_15_59/a_36_472# vss 0.404746f
C540 sarlogic_0/FILLER_0_15_59/a_572_375# vss 0.232991f
C541 sarlogic_0/FILLER_0_15_59/a_124_375# vss 0.185089f
C542 sarlogic_0/FILLER_0_3_221/a_1380_472# vss 0.345058f
C543 sarlogic_0/FILLER_0_3_221/a_932_472# vss 0.33241f
C544 sarlogic_0/FILLER_0_3_221/a_484_472# vss 0.33241f
C545 sarlogic_0/FILLER_0_3_221/a_36_472# vss 0.404746f
C546 sarlogic_0/FILLER_0_3_221/a_1468_375# vss 0.233029f
C547 sarlogic_0/FILLER_0_3_221/a_1020_375# vss 0.171606f
C548 sarlogic_0/FILLER_0_3_221/a_572_375# vss 0.171606f
C549 sarlogic_0/FILLER_0_3_221/a_124_375# vss 0.185399f
C550 sarlogic_0/FILLER_0_19_187/a_484_472# vss 0.345058f
C551 sarlogic_0/FILLER_0_19_187/a_36_472# vss 0.404746f
C552 sarlogic_0/FILLER_0_19_187/a_572_375# vss 0.232991f
C553 sarlogic_0/FILLER_0_19_187/a_124_375# vss 0.185089f
C554 sarlogic_0/FILLER_0_20_15/a_1380_472# vss 0.345058f
C555 sarlogic_0/FILLER_0_20_15/a_932_472# vss 0.33241f
C556 sarlogic_0/FILLER_0_20_15/a_484_472# vss 0.33241f
C557 sarlogic_0/FILLER_0_20_15/a_36_472# vss 0.404746f
C558 sarlogic_0/FILLER_0_20_15/a_1468_375# vss 0.233029f
C559 sarlogic_0/FILLER_0_20_15/a_1020_375# vss 0.171606f
C560 sarlogic_0/FILLER_0_20_15/a_572_375# vss 0.171606f
C561 sarlogic_0/FILLER_0_20_15/a_124_375# vss 0.185399f
C562 sarlogic_0/_204_/a_67_603# vss 0.345683f
C563 sarlogic_0/_419_/a_2560_156# vss 0.016968f
C564 sarlogic_0/_419_/a_2665_112# vss 0.62251f
C565 sarlogic_0/_419_/a_2248_156# vss 0.371662f
C566 sarlogic_0/_419_/a_1204_472# vss 0.012971f
C567 sarlogic_0/_419_/a_1000_472# vss 0.291735f
C568 sarlogic_0/_419_/a_796_472# vss 0.023206f
C569 sarlogic_0/_419_/a_1308_423# vss 0.279043f
C570 sarlogic_0/_419_/a_448_472# vss 0.684413f
C571 sarlogic_0/_419_/a_36_151# vss 1.43589f
C572 sarlogic_0/_054_ vss 0.522819f
C573 sarlogic_0/_221_/a_36_160# vss 0.386641f
C574 sarlogic_0/FILLER_0_9_270/a_484_472# vss 0.345058f
C575 sarlogic_0/FILLER_0_9_270/a_36_472# vss 0.404746f
C576 sarlogic_0/FILLER_0_9_270/a_572_375# vss 0.232991f
C577 sarlogic_0/FILLER_0_9_270/a_124_375# vss 0.185089f
C578 sarlogic_0/FILLER_0_1_192/a_36_472# vss 0.417394f
C579 sarlogic_0/FILLER_0_1_192/a_124_375# vss 0.246306f
C580 sarlogic_0/FILLER_0_13_80/a_36_472# vss 0.417394f
C581 sarlogic_0/FILLER_0_13_80/a_124_375# vss 0.246306f
C582 sarlogic_0/_153_ vss 1.165862f
C583 sarlogic_0/_154_ vss 1.167112f
C584 sarlogic_0/_367_/a_36_68# vss 0.150048f
C585 sarlogic_0/_436_/a_2560_156# vss 0.016968f
C586 sarlogic_0/_436_/a_2665_112# vss 0.62251f
C587 sarlogic_0/_436_/a_2248_156# vss 0.371662f
C588 sarlogic_0/_436_/a_1204_472# vss 0.012971f
C589 sarlogic_0/_436_/a_1000_472# vss 0.291735f
C590 sarlogic_0/_436_/a_796_472# vss 0.023206f
C591 sarlogic_0/_436_/a_1308_423# vss 0.279043f
C592 sarlogic_0/_436_/a_448_472# vss 0.684413f
C593 sarlogic_0/_436_/a_36_151# vss 1.43589f
C594 sarlogic_0/FILLER_0_10_107/a_484_472# vss 0.345058f
C595 sarlogic_0/FILLER_0_10_107/a_36_472# vss 0.404746f
C596 sarlogic_0/FILLER_0_10_107/a_572_375# vss 0.232991f
C597 sarlogic_0/FILLER_0_10_107/a_124_375# vss 0.185089f
C598 sarlogic_0/_168_ vss 0.336537f
C599 sarlogic_0/net51 vss 2.105066f
C600 sarlogic_0/_042_ vss 0.323587f
C601 sarlogic_0/_453_/a_2560_156# vss 0.016968f
C602 sarlogic_0/_453_/a_2665_112# vss 0.62251f
C603 sarlogic_0/_453_/a_2248_156# vss 0.371662f
C604 sarlogic_0/_453_/a_1204_472# vss 0.012971f
C605 sarlogic_0/_453_/a_1000_472# vss 0.291735f
C606 sarlogic_0/_453_/a_796_472# vss 0.023206f
C607 sarlogic_0/_453_/a_1308_423# vss 0.279043f
C608 sarlogic_0/_453_/a_448_472# vss 0.684413f
C609 sarlogic_0/_453_/a_36_151# vss 1.43589f
C610 sarlogic_0/FILLER_0_19_142/a_36_472# vss 0.417394f
C611 sarlogic_0/FILLER_0_19_142/a_124_375# vss 0.246306f
C612 sarlogic_0/_048_ vss 0.358805f
C613 sarlogic_0/_205_/a_36_160# vss 0.696445f
C614 sarlogic_0/net43 vss 1.236377f
C615 sarlogic_0/FILLER_0_3_78/a_484_472# vss 0.345058f
C616 sarlogic_0/FILLER_0_3_78/a_36_472# vss 0.404746f
C617 sarlogic_0/FILLER_0_3_78/a_572_375# vss 0.232991f
C618 sarlogic_0/FILLER_0_3_78/a_124_375# vss 0.185089f
C619 sarlogic_0/_437_/a_2560_156# vss 0.016968f
C620 sarlogic_0/_437_/a_2665_112# vss 0.62251f
C621 sarlogic_0/_437_/a_2248_156# vss 0.371662f
C622 sarlogic_0/_437_/a_1204_472# vss 0.012971f
C623 sarlogic_0/_437_/a_1000_472# vss 0.291735f
C624 sarlogic_0/_437_/a_796_472# vss 0.023206f
C625 sarlogic_0/_437_/a_1308_423# vss 0.279043f
C626 sarlogic_0/_437_/a_448_472# vss 0.684413f
C627 sarlogic_0/_437_/a_36_151# vss 1.43589f
C628 sarlogic_0/_109_ vss 0.319326f
C629 sarlogic_0/_299_/a_36_472# vss 0.031137f
C630 sarlogic_0/net37 vss 1.529713f
C631 sarlogic_0/_385_/a_36_68# vss 0.112263f
C632 sarlogic_0/FILLER_0_0_266/a_36_472# vss 0.417394f
C633 sarlogic_0/FILLER_0_0_266/a_124_375# vss 0.246306f
C634 sarlogic_0/net12 vss 1.263595f
C635 sarlogic_0/net22 vss 2.108509f
C636 sarlogic_0/FILLER_0_9_290/a_36_472# vss 0.417394f
C637 sarlogic_0/FILLER_0_9_290/a_124_375# vss 0.246306f
C638 sarlogic_0/_223_/a_36_160# vss 0.696445f
C639 sarlogic_0/FILLER_0_14_263/a_36_472# vss 0.417394f
C640 sarlogic_0/FILLER_0_14_263/a_124_375# vss 0.246306f
C641 sarlogic_0/_158_ vss 0.309522f
C642 sarlogic_0/_369_/a_36_68# vss 0.150048f
C643 sarlogic_0/net71 vss 1.420869f
C644 sarlogic_0/_438_/a_2560_156# vss 0.016968f
C645 sarlogic_0/_438_/a_2665_112# vss 0.62251f
C646 sarlogic_0/_438_/a_2248_156# vss 0.371662f
C647 sarlogic_0/_438_/a_1204_472# vss 0.012971f
C648 sarlogic_0/_438_/a_1000_472# vss 0.291735f
C649 sarlogic_0/_438_/a_796_472# vss 0.023206f
C650 sarlogic_0/_438_/a_1308_423# vss 0.279043f
C651 sarlogic_0/_438_/a_448_472# vss 0.684413f
C652 sarlogic_0/_438_/a_36_151# vss 1.43589f
C653 sarlogic_0/FILLER_0_23_274/a_36_472# vss 0.417394f
C654 sarlogic_0/FILLER_0_23_274/a_124_375# vss 0.246306f
C655 sarlogic_0/FILLER_0_17_282/a_36_472# vss 0.417394f
C656 sarlogic_0/FILLER_0_17_282/a_124_375# vss 0.246306f
C657 sarlogic_0/FILLER_0_5_198/a_484_472# vss 0.345058f
C658 sarlogic_0/FILLER_0_5_198/a_36_472# vss 0.404746f
C659 sarlogic_0/FILLER_0_5_198/a_572_375# vss 0.232991f
C660 sarlogic_0/FILLER_0_5_198/a_124_375# vss 0.185089f
C661 sarlogic_0/_163_ vss 1.03762f
C662 sarlogic_0/_169_ vss 0.245383f
C663 sarlogic_0/_386_/a_848_380# vss 0.40208f
C664 sarlogic_0/_386_/a_124_24# vss 0.591898f
C665 sarlogic_0/FILLER_0_20_2/a_484_472# vss 0.345058f
C666 sarlogic_0/FILLER_0_20_2/a_36_472# vss 0.404746f
C667 sarlogic_0/FILLER_0_20_2/a_572_375# vss 0.232991f
C668 sarlogic_0/FILLER_0_20_2/a_124_375# vss 0.185089f
C669 sarlogic_0/FILLER_0_16_154/a_1380_472# vss 0.345058f
C670 sarlogic_0/FILLER_0_16_154/a_932_472# vss 0.33241f
C671 sarlogic_0/FILLER_0_16_154/a_484_472# vss 0.33241f
C672 sarlogic_0/FILLER_0_16_154/a_36_472# vss 0.404746f
C673 sarlogic_0/FILLER_0_16_154/a_1468_375# vss 0.233029f
C674 sarlogic_0/FILLER_0_16_154/a_1020_375# vss 0.171606f
C675 sarlogic_0/FILLER_0_16_154/a_572_375# vss 0.171606f
C676 sarlogic_0/FILLER_0_16_154/a_124_375# vss 0.185399f
C677 sarlogic_0/FILLER_0_0_232/a_36_472# vss 0.417394f
C678 sarlogic_0/FILLER_0_0_232/a_124_375# vss 0.246306f
C679 sarlogic_0/FILLER_0_19_195/a_36_472# vss 0.417394f
C680 sarlogic_0/FILLER_0_19_195/a_124_375# vss 0.246306f
C681 sarlogic_0/_049_ vss 0.329957f
C682 sarlogic_0/net33 vss 1.934915f
C683 sarlogic_0/_207_/a_67_603# vss 0.345683f
C684 sarlogic_0/FILLER_0_3_54/a_36_472# vss 0.417394f
C685 sarlogic_0/FILLER_0_3_54/a_124_375# vss 0.246306f
C686 sarlogic_0/FILLER_0_2_101/a_36_472# vss 0.417394f
C687 sarlogic_0/FILLER_0_2_101/a_124_375# vss 0.246306f
C688 sarlogic_0/trim_mask\[0\] vss 0.605753f
C689 sarlogic_0/_439_/a_2560_156# vss 0.016968f
C690 sarlogic_0/_439_/a_2665_112# vss 0.62251f
C691 sarlogic_0/_439_/a_2248_156# vss 0.371662f
C692 sarlogic_0/_439_/a_1204_472# vss 0.012971f
C693 sarlogic_0/_439_/a_1000_472# vss 0.291735f
C694 sarlogic_0/_439_/a_796_472# vss 0.023206f
C695 sarlogic_0/_439_/a_1308_423# vss 0.279043f
C696 sarlogic_0/_439_/a_448_472# vss 0.684413f
C697 sarlogic_0/_439_/a_36_151# vss 1.43589f
C698 sarlogic_0/_066_ vss 0.333041f
C699 sarlogic_0/FILLER_0_23_44/a_1380_472# vss 0.345058f
C700 sarlogic_0/FILLER_0_23_44/a_932_472# vss 0.33241f
C701 sarlogic_0/FILLER_0_23_44/a_484_472# vss 0.33241f
C702 sarlogic_0/FILLER_0_23_44/a_36_472# vss 0.404746f
C703 sarlogic_0/FILLER_0_23_44/a_1468_375# vss 0.233029f
C704 sarlogic_0/FILLER_0_23_44/a_1020_375# vss 0.171606f
C705 sarlogic_0/FILLER_0_23_44/a_572_375# vss 0.171606f
C706 sarlogic_0/FILLER_0_23_44/a_124_375# vss 0.185399f
C707 sarlogic_0/FILLER_0_23_88/a_36_472# vss 0.417394f
C708 sarlogic_0/FILLER_0_23_88/a_124_375# vss 0.246306f
C709 sarlogic_0/FILLER_0_5_164/a_484_472# vss 0.345058f
C710 sarlogic_0/FILLER_0_5_164/a_36_472# vss 0.404746f
C711 sarlogic_0/FILLER_0_5_164/a_572_375# vss 0.232991f
C712 sarlogic_0/FILLER_0_5_164/a_124_375# vss 0.185089f
C713 sarlogic_0/_060_ vss 2.485177f
C714 sarlogic_0/_113_ vss 2.833205f
C715 sarlogic_0/_090_ vss 2.629271f
C716 sarlogic_0/_310_/a_49_472# vss 0.098072f
C717 sarlogic_0/_037_ vss 0.467089f
C718 sarlogic_0/_170_ vss 0.413995f
C719 sarlogic_0/_387_/a_36_113# vss 0.418095f
C720 sarlogic_0/_208_/a_36_160# vss 0.696445f
C721 sarlogic_0/FILLER_0_18_76/a_484_472# vss 0.345058f
C722 sarlogic_0/FILLER_0_18_76/a_36_472# vss 0.404746f
C723 sarlogic_0/FILLER_0_18_76/a_572_375# vss 0.232991f
C724 sarlogic_0/FILLER_0_18_76/a_124_375# vss 0.185089f
C725 sarlogic_0/_225_/a_36_160# vss 0.386641f
C726 sarlogic_0/FILLER_0_2_177/a_484_472# vss 0.345058f
C727 sarlogic_0/FILLER_0_2_177/a_36_472# vss 0.404746f
C728 sarlogic_0/FILLER_0_2_177/a_572_375# vss 0.232991f
C729 sarlogic_0/FILLER_0_2_177/a_124_375# vss 0.185089f
C730 sarlogic_0/FILLER_0_2_111/a_1380_472# vss 0.345058f
C731 sarlogic_0/FILLER_0_2_111/a_932_472# vss 0.33241f
C732 sarlogic_0/FILLER_0_2_111/a_484_472# vss 0.33241f
C733 sarlogic_0/FILLER_0_2_111/a_36_472# vss 0.404746f
C734 sarlogic_0/FILLER_0_2_111/a_1468_375# vss 0.233029f
C735 sarlogic_0/FILLER_0_2_111/a_1020_375# vss 0.171606f
C736 sarlogic_0/FILLER_0_2_111/a_572_375# vss 0.171606f
C737 sarlogic_0/FILLER_0_2_111/a_124_375# vss 0.185399f
C738 sarlogic_0/FILLER_0_15_228/a_36_472# vss 0.417394f
C739 sarlogic_0/FILLER_0_15_228/a_124_375# vss 0.246306f
C740 sarlogic_0/net47 vss 2.314376f
C741 sarlogic_0/_242_/a_36_160# vss 0.696445f
C742 sarlogic_0/_117_ vss 1.266251f
C743 sarlogic_0/_311_/a_66_473# vss 0.11665f
C744 sarlogic_0/_043_ vss 0.487279f
C745 sarlogic_0/_190_/a_36_160# vss 0.696445f
C746 sarlogic_0/FILLER_0_9_105/a_484_472# vss 0.345058f
C747 sarlogic_0/FILLER_0_9_105/a_36_472# vss 0.404746f
C748 sarlogic_0/FILLER_0_9_105/a_572_375# vss 0.232991f
C749 sarlogic_0/FILLER_0_9_105/a_124_375# vss 0.185089f
C750 sarlogic_0/FILLER_0_13_100/a_36_472# vss 0.417394f
C751 sarlogic_0/FILLER_0_13_100/a_124_375# vss 0.246306f
C752 sarlogic_0/FILLER_0_22_177/a_1380_472# vss 0.345058f
C753 sarlogic_0/FILLER_0_22_177/a_932_472# vss 0.33241f
C754 sarlogic_0/FILLER_0_22_177/a_484_472# vss 0.33241f
C755 sarlogic_0/FILLER_0_22_177/a_36_472# vss 0.404746f
C756 sarlogic_0/FILLER_0_22_177/a_1468_375# vss 0.233029f
C757 sarlogic_0/FILLER_0_22_177/a_1020_375# vss 0.171606f
C758 sarlogic_0/FILLER_0_22_177/a_572_375# vss 0.171606f
C759 sarlogic_0/FILLER_0_22_177/a_124_375# vss 0.185399f
C760 sarlogic_0/FILLER_0_15_2/a_484_472# vss 0.345058f
C761 sarlogic_0/FILLER_0_15_2/a_36_472# vss 0.404746f
C762 sarlogic_0/FILLER_0_15_2/a_572_375# vss 0.232991f
C763 sarlogic_0/FILLER_0_15_2/a_124_375# vss 0.185089f
C764 sarlogic_0/FILLER_0_15_10/a_36_472# vss 0.417394f
C765 sarlogic_0/FILLER_0_15_10/a_124_375# vss 0.246306f
C766 sarlogic_0/FILLER_0_19_171/a_1380_472# vss 0.345058f
C767 sarlogic_0/FILLER_0_19_171/a_932_472# vss 0.33241f
C768 sarlogic_0/FILLER_0_19_171/a_484_472# vss 0.33241f
C769 sarlogic_0/FILLER_0_19_171/a_36_472# vss 0.404746f
C770 sarlogic_0/FILLER_0_19_171/a_1468_375# vss 0.233029f
C771 sarlogic_0/FILLER_0_19_171/a_1020_375# vss 0.171606f
C772 sarlogic_0/FILLER_0_19_171/a_572_375# vss 0.171606f
C773 sarlogic_0/FILLER_0_19_171/a_124_375# vss 0.185399f
C774 sarlogic_0/net13 vss 1.176306f
C775 sarlogic_0/net23 vss 2.091399f
C776 sarlogic_0/FILLER_0_20_87/a_36_472# vss 0.417394f
C777 sarlogic_0/FILLER_0_20_87/a_124_375# vss 0.246306f
C778 sarlogic_0/FILLER_0_20_98/a_36_472# vss 0.417394f
C779 sarlogic_0/FILLER_0_20_98/a_124_375# vss 0.246306f
C780 sarlogic_0/_055_ vss 1.782885f
C781 sarlogic_0/FILLER_0_18_53/a_484_472# vss 0.345058f
C782 sarlogic_0/FILLER_0_18_53/a_36_472# vss 0.404746f
C783 sarlogic_0/FILLER_0_18_53/a_572_375# vss 0.232991f
C784 sarlogic_0/FILLER_0_18_53/a_124_375# vss 0.185089f
C785 sarlogic_0/FILLER_0_2_165/a_36_472# vss 0.417394f
C786 sarlogic_0/FILLER_0_2_165/a_124_375# vss 0.246306f
C787 sarlogic_0/FILLER_0_15_205/a_36_472# vss 0.417394f
C788 sarlogic_0/FILLER_0_15_205/a_124_375# vss 0.246306f
C789 sarlogic_0/FILLER_0_23_282/a_484_472# vss 0.345058f
C790 sarlogic_0/FILLER_0_23_282/a_36_472# vss 0.404746f
C791 sarlogic_0/FILLER_0_23_282/a_572_375# vss 0.232991f
C792 sarlogic_0/FILLER_0_23_282/a_124_375# vss 0.185089f
C793 sarlogic_0/net42 vss 1.067446f
C794 sarlogic_0/net17 vss 2.210219f
C795 sarlogic_0/_172_ vss 0.265782f
C796 sarlogic_0/_171_ vss 0.300355f
C797 sarlogic_0/_389_/a_36_148# vss 0.388358f
C798 sarlogic_0/_080_ vss 0.328202f
C799 sarlogic_0/_260_/a_36_68# vss 0.112263f
C800 sarlogic_0/FILLER_0_0_96/a_36_472# vss 0.417394f
C801 sarlogic_0/FILLER_0_0_96/a_124_375# vss 0.246306f
C802 sarlogic_0/FILLER_0_9_72/a_1380_472# vss 0.345058f
C803 sarlogic_0/FILLER_0_9_72/a_932_472# vss 0.33241f
C804 sarlogic_0/FILLER_0_9_72/a_484_472# vss 0.33241f
C805 sarlogic_0/FILLER_0_9_72/a_36_472# vss 0.404746f
C806 sarlogic_0/FILLER_0_9_72/a_1468_375# vss 0.233029f
C807 sarlogic_0/FILLER_0_9_72/a_1020_375# vss 0.171606f
C808 sarlogic_0/FILLER_0_9_72/a_572_375# vss 0.171606f
C809 sarlogic_0/FILLER_0_9_72/a_124_375# vss 0.185399f
C810 sarlogic_0/FILLER_0_20_31/a_36_472# vss 0.417394f
C811 sarlogic_0/FILLER_0_20_31/a_124_375# vss 0.246306f
C812 sarlogic_0/_227_/a_36_160# vss 0.386641f
C813 sarlogic_0/_120_ vss 1.533088f
C814 sarlogic_0/_313_/a_67_603# vss 0.345683f
C815 sarlogic_0/FILLER_0_5_172/a_36_472# vss 0.417394f
C816 sarlogic_0/FILLER_0_5_172/a_124_375# vss 0.246306f
C817 sarlogic_0/FILLER_0_12_20/a_484_472# vss 0.345058f
C818 sarlogic_0/FILLER_0_12_20/a_36_472# vss 0.404746f
C819 sarlogic_0/FILLER_0_12_20/a_572_375# vss 0.232991f
C820 sarlogic_0/FILLER_0_12_20/a_124_375# vss 0.185089f
C821 sarlogic_0/_134_ vss 0.365972f
C822 sarlogic_0/_062_ vss 1.717773f
C823 sarlogic_0/_059_ vss 1.686761f
C824 sarlogic_0/_261_/a_36_160# vss 0.386641f
C825 sarlogic_0/_044_ vss 0.388801f
C826 sarlogic_0/mask\[1\] vss 1.295078f
C827 sarlogic_0/_192_/a_67_603# vss 0.345683f
C828 sarlogic_0/FILLER_0_13_142/a_1380_472# vss 0.345058f
C829 sarlogic_0/FILLER_0_13_142/a_932_472# vss 0.33241f
C830 sarlogic_0/FILLER_0_13_142/a_484_472# vss 0.33241f
C831 sarlogic_0/FILLER_0_13_142/a_36_472# vss 0.404746f
C832 sarlogic_0/FILLER_0_13_142/a_1468_375# vss 0.233029f
C833 sarlogic_0/FILLER_0_13_142/a_1020_375# vss 0.171606f
C834 sarlogic_0/FILLER_0_13_142/a_572_375# vss 0.171606f
C835 sarlogic_0/FILLER_0_13_142/a_124_375# vss 0.185399f
C836 sarlogic_0/FILLER_0_9_60/a_484_472# vss 0.345058f
C837 sarlogic_0/FILLER_0_9_60/a_36_472# vss 0.404746f
C838 sarlogic_0/FILLER_0_9_60/a_572_375# vss 0.232991f
C839 sarlogic_0/FILLER_0_9_60/a_124_375# vss 0.185089f
C840 sarlogic_0/FILLER_0_7_233/a_36_472# vss 0.417394f
C841 sarlogic_0/FILLER_0_7_233/a_124_375# vss 0.246306f
C842 sarlogic_0/_228_/a_36_68# vss 0.69549f
C843 sarlogic_0/FILLER_0_21_206/a_36_472# vss 0.417394f
C844 sarlogic_0/FILLER_0_21_206/a_124_375# vss 0.246306f
C845 sarlogic_0/_067_ vss 0.851951f
C846 sarlogic_0/_135_ vss 0.339478f
C847 sarlogic_0/_193_/a_36_160# vss 0.696445f
C848 sarlogic_0/_180_ vss 0.390598f
C849 sarlogic_0/cal_count\[1\] vss 1.568289f
C850 sarlogic_0/FILLER_0_4_213/a_484_472# vss 0.345058f
C851 sarlogic_0/FILLER_0_4_213/a_36_472# vss 0.404746f
C852 sarlogic_0/FILLER_0_4_213/a_572_375# vss 0.232991f
C853 sarlogic_0/FILLER_0_4_213/a_124_375# vss 0.185089f
C854 sarlogic_0/FILLER_0_11_282/a_36_472# vss 0.417394f
C855 sarlogic_0/FILLER_0_11_282/a_124_375# vss 0.246306f
C856 sarlogic_0/FILLER_0_18_61/a_36_472# vss 0.417394f
C857 sarlogic_0/FILLER_0_18_61/a_124_375# vss 0.246306f
C858 sarlogic_0/FILLER_0_15_235/a_484_472# vss 0.345058f
C859 sarlogic_0/FILLER_0_15_235/a_36_472# vss 0.404746f
C860 sarlogic_0/FILLER_0_15_235/a_572_375# vss 0.232991f
C861 sarlogic_0/FILLER_0_15_235/a_124_375# vss 0.185089f
C862 sarlogic_0/FILLER_0_23_290/a_36_472# vss 0.417394f
C863 sarlogic_0/FILLER_0_23_290/a_124_375# vss 0.246306f
C864 sarlogic_0/_121_ vss 0.532847f
C865 sarlogic_0/_315_/a_36_68# vss 0.052951f
C866 sarlogic_0/_246_/a_36_68# vss 0.69549f
C867 sarlogic_0/FILLER_0_5_181/a_36_472# vss 0.417394f
C868 sarlogic_0/FILLER_0_5_181/a_124_375# vss 0.246306f
C869 sarlogic_0/_082_ vss 0.619901f
C870 sarlogic_0/net8 vss 1.163723f
C871 sarlogic_0/net18 vss 2.032159f
C872 sarlogic_0/_332_/a_36_472# vss 0.031137f
C873 sarlogic_0/_179_ vss 0.336984f
C874 sarlogic_0/_401_/a_36_68# vss 0.112263f
C875 sarlogic_0/FILLER_0_14_107/a_1380_472# vss 0.345058f
C876 sarlogic_0/FILLER_0_14_107/a_932_472# vss 0.33241f
C877 sarlogic_0/FILLER_0_14_107/a_484_472# vss 0.33241f
C878 sarlogic_0/FILLER_0_14_107/a_36_472# vss 0.404746f
C879 sarlogic_0/FILLER_0_14_107/a_1468_375# vss 0.233029f
C880 sarlogic_0/FILLER_0_14_107/a_1020_375# vss 0.171606f
C881 sarlogic_0/FILLER_0_14_107/a_572_375# vss 0.171606f
C882 sarlogic_0/FILLER_0_14_107/a_124_375# vss 0.185399f
C883 sarlogic_0/_097_ vss 0.592554f
C884 sarlogic_0/FILLER_0_1_204/a_36_472# vss 0.417394f
C885 sarlogic_0/FILLER_0_1_204/a_124_375# vss 0.246306f
C886 sarlogic_0/FILLER_0_15_72/a_484_472# vss 0.345058f
C887 sarlogic_0/FILLER_0_15_72/a_36_472# vss 0.404746f
C888 sarlogic_0/FILLER_0_15_72/a_572_375# vss 0.232991f
C889 sarlogic_0/FILLER_0_15_72/a_124_375# vss 0.185089f
C890 sarlogic_0/FILLER_0_17_104/a_1380_472# vss 0.345058f
C891 sarlogic_0/FILLER_0_17_104/a_932_472# vss 0.33241f
C892 sarlogic_0/FILLER_0_17_104/a_484_472# vss 0.33241f
C893 sarlogic_0/FILLER_0_17_104/a_36_472# vss 0.404746f
C894 sarlogic_0/FILLER_0_17_104/a_1468_375# vss 0.233029f
C895 sarlogic_0/FILLER_0_17_104/a_1020_375# vss 0.171606f
C896 sarlogic_0/FILLER_0_17_104/a_572_375# vss 0.171606f
C897 sarlogic_0/FILLER_0_17_104/a_124_375# vss 0.185399f
C898 sarlogic_0/FILLER_0_8_37/a_484_472# vss 0.345058f
C899 sarlogic_0/FILLER_0_8_37/a_36_472# vss 0.404746f
C900 sarlogic_0/FILLER_0_8_37/a_572_375# vss 0.232991f
C901 sarlogic_0/FILLER_0_8_37/a_124_375# vss 0.185089f
C902 sarlogic_0/FILLER_0_15_212/a_1380_472# vss 0.345058f
C903 sarlogic_0/FILLER_0_15_212/a_932_472# vss 0.33241f
C904 sarlogic_0/FILLER_0_15_212/a_484_472# vss 0.33241f
C905 sarlogic_0/FILLER_0_15_212/a_36_472# vss 0.404746f
C906 sarlogic_0/FILLER_0_15_212/a_1468_375# vss 0.233029f
C907 sarlogic_0/FILLER_0_15_212/a_1020_375# vss 0.171606f
C908 sarlogic_0/FILLER_0_15_212/a_572_375# vss 0.171606f
C909 sarlogic_0/FILLER_0_15_212/a_124_375# vss 0.185399f
C910 sarlogic_0/FILLER_0_23_60/a_36_472# vss 0.417394f
C911 sarlogic_0/FILLER_0_23_60/a_124_375# vss 0.246306f
C912 sarlogic_0/_123_ vss 0.344874f
C913 sarlogic_0/_122_ vss 0.600118f
C914 sarlogic_0/calibrate vss 1.343796f
C915 sarlogic_0/_316_/a_848_380# vss 0.40208f
C916 sarlogic_0/_316_/a_124_24# vss 0.591898f
C917 sarlogic_0/_247_/a_36_160# vss 0.696445f
C918 sarlogic_0/FILLER_0_12_50/a_36_472# vss 0.417394f
C919 sarlogic_0/FILLER_0_12_50/a_124_375# vss 0.246306f
C920 sarlogic_0/_084_ vss 0.296163f
C921 sarlogic_0/cal_itt\[0\] vss 1.831055f
C922 sarlogic_0/cal_itt\[1\] vss 1.705665f
C923 sarlogic_0/FILLER_0_11_109/a_36_472# vss 0.417394f
C924 sarlogic_0/FILLER_0_11_109/a_124_375# vss 0.246306f
C925 sarlogic_0/_182_ vss 0.34197f
C926 sarlogic_0/_402_/a_1948_68# vss 0.022025f
C927 sarlogic_0/_402_/a_718_527# vss 0.001795f
C928 sarlogic_0/_402_/a_56_567# vss 0.424713f
C929 sarlogic_0/_402_/a_728_93# vss 0.65929f
C930 sarlogic_0/_402_/a_1296_93# vss 0.317801f
C931 sarlogic_0/_045_ vss 0.349338f
C932 sarlogic_0/mask\[2\] vss 1.335688f
C933 sarlogic_0/_195_/a_67_603# vss 0.345683f
C934 sarlogic_0/_333_/a_36_160# vss 0.386641f
C935 sarlogic_0/_098_ vss 1.816151f
C936 sarlogic_0/_147_ vss 0.322539f
C937 sarlogic_0/_350_/a_49_472# vss 0.054843f
C938 sarlogic_0/FILLER_0_12_236/a_484_472# vss 0.345058f
C939 sarlogic_0/FILLER_0_12_236/a_36_472# vss 0.404746f
C940 sarlogic_0/FILLER_0_12_236/a_572_375# vss 0.232991f
C941 sarlogic_0/FILLER_0_12_236/a_124_375# vss 0.185089f
C942 sarlogic_0/FILLER_0_2_171/a_36_472# vss 0.417394f
C943 sarlogic_0/FILLER_0_2_171/a_124_375# vss 0.246306f
C944 sarlogic_0/_014_ vss 0.363432f
C945 sarlogic_0/_317_/a_36_113# vss 0.418095f
C946 sarlogic_0/_248_/a_36_68# vss 0.69549f
C947 sarlogic_0/FILLER_0_17_38/a_484_472# vss 0.345058f
C948 sarlogic_0/FILLER_0_17_38/a_36_472# vss 0.404746f
C949 sarlogic_0/FILLER_0_17_38/a_572_375# vss 0.232991f
C950 sarlogic_0/FILLER_0_17_38/a_124_375# vss 0.185089f
C951 sarlogic_0/_001_ vss 0.285216f
C952 sarlogic_0/_265_/a_244_68# vss 0.138666f
C953 sarlogic_0/_196_/a_36_160# vss 0.696445f
C954 sarlogic_0/FILLER_0_6_90/a_484_472# vss 0.345058f
C955 sarlogic_0/FILLER_0_6_90/a_36_472# vss 0.404746f
C956 sarlogic_0/FILLER_0_6_90/a_572_375# vss 0.232991f
C957 sarlogic_0/FILLER_0_6_90/a_124_375# vss 0.185089f
C958 sarlogic_0/_183_ vss 0.356629f
C959 sarlogic_0/_334_/a_36_160# vss 0.386641f
C960 sarlogic_0/_282_/a_36_160# vss 0.386641f
C961 sarlogic_0/_024_ vss 0.451815f
C962 sarlogic_0/_009_ vss 0.397943f
C963 sarlogic_0/_420_/a_2560_156# vss 0.016968f
C964 sarlogic_0/_420_/a_2665_112# vss 0.62251f
C965 sarlogic_0/_420_/a_2248_156# vss 0.371662f
C966 sarlogic_0/_420_/a_1204_472# vss 0.012971f
C967 sarlogic_0/_420_/a_1000_472# vss 0.291735f
C968 sarlogic_0/_420_/a_796_472# vss 0.023206f
C969 sarlogic_0/_420_/a_1308_423# vss 0.279043f
C970 sarlogic_0/_420_/a_448_472# vss 0.684413f
C971 sarlogic_0/_420_/a_36_151# vss 1.43589f
C972 clk vss 18.686785f
C973 sarlogic_0/FILLER_0_8_2/a_36_472# vss 0.417394f
C974 sarlogic_0/FILLER_0_8_2/a_124_375# vss 0.246306f
C975 sarlogic_0/FILLER_0_8_24/a_484_472# vss 0.345058f
C976 sarlogic_0/FILLER_0_8_24/a_36_472# vss 0.404746f
C977 sarlogic_0/FILLER_0_8_24/a_572_375# vss 0.232991f
C978 sarlogic_0/FILLER_0_8_24/a_124_375# vss 0.185089f
C979 sarlogic_0/_124_ vss 0.294081f
C980 sarlogic_0/_118_ vss 1.378735f
C981 sarlogic_0/_071_ vss 1.600488f
C982 sarlogic_0/net9 vss 1.13171f
C983 sarlogic_0/net19 vss 1.889339f
C984 sarlogic_0/_138_ vss 0.33132f
C985 sarlogic_0/_137_ vss 1.178616f
C986 sarlogic_0/_335_/a_49_472# vss 0.054843f
C987 sarlogic_0/_404_/a_36_472# vss 0.031137f
C988 sarlogic_0/FILLER_0_20_107/a_36_472# vss 0.417394f
C989 sarlogic_0/FILLER_0_20_107/a_124_375# vss 0.246306f
C990 sarlogic_0/FILLER_0_9_142/a_36_472# vss 0.417394f
C991 sarlogic_0/FILLER_0_9_142/a_124_375# vss 0.246306f
C992 sarlogic_0/_099_ vss 1.152785f
C993 sarlogic_0/_283_/a_36_472# vss 0.031137f
C994 sarlogic_0/mask\[7\] vss 1.478045f
C995 sarlogic_0/_352_/a_49_472# vss 0.054843f
C996 sarlogic_0/_010_ vss 0.377779f
C997 sarlogic_0/_421_/a_2560_156# vss 0.016968f
C998 sarlogic_0/_421_/a_2665_112# vss 0.62251f
C999 sarlogic_0/_421_/a_2248_156# vss 0.371662f
C1000 sarlogic_0/_421_/a_1204_472# vss 0.012971f
C1001 sarlogic_0/_421_/a_1000_472# vss 0.291735f
C1002 sarlogic_0/_421_/a_796_472# vss 0.023206f
C1003 sarlogic_0/_421_/a_1308_423# vss 0.279043f
C1004 sarlogic_0/_421_/a_448_472# vss 0.684413f
C1005 sarlogic_0/_421_/a_36_151# vss 1.43589f
C1006 sarlogic_0/FILLER_0_1_212/a_36_472# vss 0.417394f
C1007 sarlogic_0/FILLER_0_1_212/a_124_375# vss 0.246306f
C1008 sarlogic_0/FILLER_0_8_239/a_36_472# vss 0.417394f
C1009 sarlogic_0/FILLER_0_8_239/a_124_375# vss 0.246306f
C1010 sarlogic_0/_125_ vss 1.526603f
C1011 sarlogic_0/_058_ vss 1.483584f
C1012 sarlogic_0/FILLER_0_6_177/a_484_472# vss 0.345058f
C1013 sarlogic_0/FILLER_0_6_177/a_36_472# vss 0.404746f
C1014 sarlogic_0/FILLER_0_6_177/a_572_375# vss 0.232991f
C1015 sarlogic_0/FILLER_0_6_177/a_124_375# vss 0.185089f
C1016 sarlogic_0/state\[1\] vss 2.652405f
C1017 sarlogic_0/_267_/a_36_472# vss 0.137725f
C1018 sarlogic_0/_184_ vss 0.350066f
C1019 sarlogic_0/cal_count\[2\] vss 1.971854f
C1020 sarlogic_0/_405_/a_67_603# vss 0.345683f
C1021 sarlogic_0/_018_ vss 0.358633f
C1022 sarlogic_0/_046_ vss 0.361963f
C1023 sarlogic_0/_198_/a_67_603# vss 0.345683f
C1024 sarlogic_0/_094_ vss 1.263877f
C1025 sarlogic_0/_100_ vss 0.333135f
C1026 sarlogic_0/net36 vss 2.262756f
C1027 sarlogic_0/FILLER_0_17_133/a_36_472# vss 0.417394f
C1028 sarlogic_0/FILLER_0_17_133/a_124_375# vss 0.246306f
C1029 sarlogic_0/_025_ vss 0.350324f
C1030 sarlogic_0/_148_ vss 0.325709f
C1031 sarlogic_0/_422_/a_2560_156# vss 0.016968f
C1032 sarlogic_0/_422_/a_2665_112# vss 0.62251f
C1033 sarlogic_0/_422_/a_2248_156# vss 0.371662f
C1034 sarlogic_0/_422_/a_1204_472# vss 0.012971f
C1035 sarlogic_0/_422_/a_1000_472# vss 0.291735f
C1036 sarlogic_0/_422_/a_796_472# vss 0.023206f
C1037 sarlogic_0/_422_/a_1308_423# vss 0.279043f
C1038 sarlogic_0/_422_/a_448_472# vss 0.684413f
C1039 sarlogic_0/_422_/a_36_151# vss 1.43589f
C1040 sarlogic_0/FILLER_0_1_266/a_484_472# vss 0.345058f
C1041 sarlogic_0/FILLER_0_1_266/a_36_472# vss 0.404746f
C1042 sarlogic_0/FILLER_0_1_266/a_572_375# vss 0.232991f
C1043 sarlogic_0/FILLER_0_1_266/a_124_375# vss 0.185089f
C1044 sarlogic_0/_152_ vss 0.918583f
C1045 sarlogic_0/_081_ vss 1.140656f
C1046 sarlogic_0/_370_/a_848_380# vss 0.40208f
C1047 sarlogic_0/_370_/a_124_24# vss 0.591898f
C1048 sarlogic_0/FILLER_0_24_274/a_1380_472# vss 0.345058f
C1049 sarlogic_0/FILLER_0_24_274/a_932_472# vss 0.33241f
C1050 sarlogic_0/FILLER_0_24_274/a_484_472# vss 0.33241f
C1051 sarlogic_0/FILLER_0_24_274/a_36_472# vss 0.404746f
C1052 sarlogic_0/FILLER_0_24_274/a_1468_375# vss 0.233029f
C1053 sarlogic_0/FILLER_0_24_274/a_1020_375# vss 0.171606f
C1054 sarlogic_0/FILLER_0_24_274/a_572_375# vss 0.171606f
C1055 sarlogic_0/FILLER_0_24_274/a_124_375# vss 0.185399f
C1056 sarlogic_0/_185_ vss 0.386917f
C1057 sarlogic_0/_406_/a_36_159# vss 0.374116f
C1058 sarlogic_0/_337_/a_49_472# vss 0.054843f
C1059 sarlogic_0/_199_/a_36_160# vss 0.696445f
C1060 sarlogic_0/_285_/a_36_472# vss 0.031137f
C1061 sarlogic_0/_354_/a_49_472# vss 0.054843f
C1062 sarlogic_0/_012_ vss 0.75195f
C1063 sarlogic_0/_423_/a_2560_156# vss 0.016968f
C1064 sarlogic_0/_423_/a_2665_112# vss 0.62251f
C1065 sarlogic_0/_423_/a_2248_156# vss 0.371662f
C1066 sarlogic_0/_423_/a_1204_472# vss 0.012971f
C1067 sarlogic_0/_423_/a_1000_472# vss 0.291735f
C1068 sarlogic_0/_423_/a_796_472# vss 0.023206f
C1069 sarlogic_0/_423_/a_1308_423# vss 0.279043f
C1070 sarlogic_0/_423_/a_448_472# vss 0.684413f
C1071 sarlogic_0/_423_/a_36_151# vss 1.43589f
C1072 sarlogic_0/FILLER_0_5_88/a_36_472# vss 0.417394f
C1073 sarlogic_0/FILLER_0_5_88/a_124_375# vss 0.246306f
C1074 sarlogic_0/trim_mask\[1\] vss 1.020743f
C1075 sarlogic_0/_029_ vss 0.308904f
C1076 sarlogic_0/_440_/a_2560_156# vss 0.016968f
C1077 sarlogic_0/_440_/a_2665_112# vss 0.62251f
C1078 sarlogic_0/_440_/a_2248_156# vss 0.371662f
C1079 sarlogic_0/_440_/a_1204_472# vss 0.012971f
C1080 sarlogic_0/_440_/a_1000_472# vss 0.291735f
C1081 sarlogic_0/_440_/a_796_472# vss 0.023206f
C1082 sarlogic_0/_440_/a_1308_423# vss 0.279043f
C1083 sarlogic_0/_440_/a_448_472# vss 0.684413f
C1084 sarlogic_0/_440_/a_36_151# vss 1.43589f
C1085 sarlogic_0/_159_ vss 0.351814f
C1086 sarlogic_0/_371_/a_36_113# vss 0.418095f
C1087 sarlogic_0/FILLER_0_17_56/a_484_472# vss 0.345058f
C1088 sarlogic_0/FILLER_0_17_56/a_36_472# vss 0.404746f
C1089 sarlogic_0/FILLER_0_17_56/a_572_375# vss 0.232991f
C1090 sarlogic_0/FILLER_0_17_56/a_124_375# vss 0.185089f
C1091 sarlogic_0/_083_ vss 0.527882f
C1092 sarlogic_0/_078_ vss 0.904554f
C1093 sarlogic_0/_269_/a_36_472# vss 0.031137f
C1094 sarlogic_0/_181_ vss 0.829168f
C1095 sarlogic_0/_407_/a_36_472# vss 0.031137f
C1096 sarlogic_0/_019_ vss 0.32907f
C1097 sarlogic_0/_139_ vss 0.346404f
C1098 sarlogic_0/FILLER_0_14_123/a_36_472# vss 0.417394f
C1099 sarlogic_0/FILLER_0_14_123/a_124_375# vss 0.246306f
C1100 sarlogic_0/_005_ vss 0.340993f
C1101 sarlogic_0/_101_ vss 0.280497f
C1102 sarlogic_0/_424_/a_2560_156# vss 0.016968f
C1103 sarlogic_0/_424_/a_2665_112# vss 0.62251f
C1104 sarlogic_0/_424_/a_2248_156# vss 0.371662f
C1105 sarlogic_0/_424_/a_1204_472# vss 0.012971f
C1106 sarlogic_0/_424_/a_1000_472# vss 0.291735f
C1107 sarlogic_0/_424_/a_796_472# vss 0.023206f
C1108 sarlogic_0/_424_/a_1308_423# vss 0.279043f
C1109 sarlogic_0/_424_/a_448_472# vss 0.684413f
C1110 sarlogic_0/_424_/a_36_151# vss 1.43589f
C1111 sarlogic_0/_026_ vss 0.320379f
C1112 sarlogic_0/_149_ vss 0.305496f
C1113 sarlogic_0/FILLER_0_5_54/a_1380_472# vss 0.345058f
C1114 sarlogic_0/FILLER_0_5_54/a_932_472# vss 0.33241f
C1115 sarlogic_0/FILLER_0_5_54/a_484_472# vss 0.33241f
C1116 sarlogic_0/FILLER_0_5_54/a_36_472# vss 0.404746f
C1117 sarlogic_0/FILLER_0_5_54/a_1468_375# vss 0.233029f
C1118 sarlogic_0/FILLER_0_5_54/a_1020_375# vss 0.171606f
C1119 sarlogic_0/FILLER_0_5_54/a_572_375# vss 0.171606f
C1120 sarlogic_0/FILLER_0_5_54/a_124_375# vss 0.185399f
C1121 sarlogic_0/FILLER_0_17_142/a_484_472# vss 0.345058f
C1122 sarlogic_0/FILLER_0_17_142/a_36_472# vss 0.404746f
C1123 sarlogic_0/FILLER_0_17_142/a_572_375# vss 0.232991f
C1124 sarlogic_0/FILLER_0_17_142/a_124_375# vss 0.185089f
C1125 sarlogic_0/_068_ vss 3.162692f
C1126 sarlogic_0/_076_ vss 3.812442f
C1127 sarlogic_0/_133_ vss 1.430901f
C1128 sarlogic_0/_070_ vss 3.115722f
C1129 sarlogic_0/_372_/a_170_472# vss 0.077257f
C1130 sarlogic_0/net49 vss 5.140563f
C1131 sarlogic_0/_030_ vss 0.307083f
C1132 sarlogic_0/net66 vss 1.472669f
C1133 sarlogic_0/_441_/a_2560_156# vss 0.016968f
C1134 sarlogic_0/_441_/a_2665_112# vss 0.62251f
C1135 sarlogic_0/_441_/a_2248_156# vss 0.371662f
C1136 sarlogic_0/_441_/a_1204_472# vss 0.012971f
C1137 sarlogic_0/_441_/a_1000_472# vss 0.291735f
C1138 sarlogic_0/_441_/a_796_472# vss 0.023206f
C1139 sarlogic_0/_441_/a_1308_423# vss 0.279043f
C1140 sarlogic_0/_441_/a_448_472# vss 0.684413f
C1141 sarlogic_0/_441_/a_36_151# vss 1.43589f
C1142 sarlogic_0/FILLER_0_5_206/a_36_472# vss 0.417394f
C1143 sarlogic_0/FILLER_0_5_206/a_124_375# vss 0.246306f
C1144 sarlogic_0/fanout49/a_36_160# vss 0.696445f
C1145 sarlogic_0/FILLER_0_8_247/a_1380_472# vss 0.345058f
C1146 sarlogic_0/FILLER_0_8_247/a_932_472# vss 0.33241f
C1147 sarlogic_0/FILLER_0_8_247/a_484_472# vss 0.33241f
C1148 sarlogic_0/FILLER_0_8_247/a_36_472# vss 0.404746f
C1149 sarlogic_0/FILLER_0_8_247/a_1468_375# vss 0.233029f
C1150 sarlogic_0/FILLER_0_8_247/a_1020_375# vss 0.171606f
C1151 sarlogic_0/FILLER_0_8_247/a_572_375# vss 0.171606f
C1152 sarlogic_0/FILLER_0_8_247/a_124_375# vss 0.185399f
C1153 sarlogic_0/FILLER_0_12_220/a_1380_472# vss 0.345058f
C1154 sarlogic_0/FILLER_0_12_220/a_932_472# vss 0.33241f
C1155 sarlogic_0/FILLER_0_12_220/a_484_472# vss 0.33241f
C1156 sarlogic_0/FILLER_0_12_220/a_36_472# vss 0.404746f
C1157 sarlogic_0/FILLER_0_12_220/a_1468_375# vss 0.233029f
C1158 sarlogic_0/FILLER_0_12_220/a_1020_375# vss 0.171606f
C1159 sarlogic_0/FILLER_0_12_220/a_572_375# vss 0.171606f
C1160 sarlogic_0/FILLER_0_12_220/a_124_375# vss 0.185399f
C1161 sarlogic_0/FILLER_0_21_286/a_484_472# vss 0.345058f
C1162 sarlogic_0/FILLER_0_21_286/a_36_472# vss 0.404746f
C1163 sarlogic_0/FILLER_0_21_286/a_572_375# vss 0.232991f
C1164 sarlogic_0/FILLER_0_21_286/a_124_375# vss 0.185089f
C1165 sarlogic_0/_140_ vss 1.276518f
C1166 sarlogic_0/_339_/a_36_160# vss 0.386641f
C1167 sarlogic_0/_095_ vss 2.689027f
C1168 sarlogic_0/_186_ vss 0.580923f
C1169 sarlogic_0/_408_/a_1936_472# vss 0.009918f
C1170 sarlogic_0/_408_/a_718_524# vss 0.005143f
C1171 sarlogic_0/_408_/a_56_524# vss 0.41096f
C1172 sarlogic_0/_408_/a_728_93# vss 0.654825f
C1173 sarlogic_0/_408_/a_1336_472# vss 0.316639f
C1174 sarlogic_0/FILLER_0_20_169/a_36_472# vss 0.417394f
C1175 sarlogic_0/FILLER_0_20_169/a_124_375# vss 0.246306f
C1176 sarlogic_0/_210_/a_67_603# vss 0.345683f
C1177 sarlogic_0/_425_/a_2560_156# vss 0.016968f
C1178 sarlogic_0/_425_/a_2665_112# vss 0.62251f
C1179 sarlogic_0/_425_/a_2248_156# vss 0.371662f
C1180 sarlogic_0/_425_/a_1204_472# vss 0.012971f
C1181 sarlogic_0/_425_/a_1000_472# vss 0.291735f
C1182 sarlogic_0/_425_/a_796_472# vss 0.023206f
C1183 sarlogic_0/_425_/a_1308_423# vss 0.279043f
C1184 sarlogic_0/_425_/a_448_472# vss 0.684413f
C1185 sarlogic_0/_425_/a_36_151# vss 1.43589f
C1186 sarlogic_0/net5 vss 0.610761f
C1187 sarlogic_0/input5/a_36_113# vss 0.418095f
C1188 sarlogic_0/FILLER_0_11_78/a_484_472# vss 0.345058f
C1189 sarlogic_0/FILLER_0_11_78/a_36_472# vss 0.404746f
C1190 sarlogic_0/FILLER_0_11_78/a_572_375# vss 0.232991f
C1191 sarlogic_0/FILLER_0_11_78/a_124_375# vss 0.185089f
C1192 sarlogic_0/_102_ vss 0.335308f
C1193 sarlogic_0/_287_/a_36_472# vss 0.031137f
C1194 sarlogic_0/mask\[9\] vss 1.383606f
C1195 sarlogic_0/_356_/a_36_472# vss 0.031137f
C1196 sarlogic_0/_031_ vss 0.417351f
C1197 sarlogic_0/net69 vss 1.020293f
C1198 sarlogic_0/_442_/a_2560_156# vss 0.016968f
C1199 sarlogic_0/_442_/a_2665_112# vss 0.62251f
C1200 sarlogic_0/_442_/a_2248_156# vss 0.371662f
C1201 sarlogic_0/_442_/a_1204_472# vss 0.012971f
C1202 sarlogic_0/_442_/a_1000_472# vss 0.291735f
C1203 sarlogic_0/_442_/a_796_472# vss 0.023206f
C1204 sarlogic_0/_442_/a_1308_423# vss 0.279043f
C1205 sarlogic_0/_442_/a_448_472# vss 0.684413f
C1206 sarlogic_0/_442_/a_36_151# vss 1.43589f
C1207 sarlogic_0/net64 vss 2.598514f
C1208 sarlogic_0/fanout59/a_36_160# vss 0.696445f
C1209 sarlogic_0/FILLER_0_14_99/a_36_472# vss 0.417394f
C1210 sarlogic_0/FILLER_0_14_99/a_124_375# vss 0.246306f
C1211 sarlogic_0/_038_ vss 0.362839f
C1212 sarlogic_0/_136_ vss 1.345638f
C1213 sarlogic_0/_390_/a_36_68# vss 0.150048f
C1214 sarlogic_0/FILLER_0_15_282/a_484_472# vss 0.345058f
C1215 sarlogic_0/FILLER_0_15_282/a_36_472# vss 0.404746f
C1216 sarlogic_0/FILLER_0_15_282/a_572_375# vss 0.232991f
C1217 sarlogic_0/FILLER_0_15_282/a_124_375# vss 0.185089f
C1218 sarlogic_0/FILLER_0_11_124/a_36_472# vss 0.417394f
C1219 sarlogic_0/FILLER_0_11_124/a_124_375# vss 0.246306f
C1220 sarlogic_0/FILLER_0_11_135/a_36_472# vss 0.417394f
C1221 sarlogic_0/FILLER_0_11_135/a_124_375# vss 0.246306f
C1222 sarlogic_0/_188_ vss 0.349407f
C1223 sarlogic_0/cal_count\[3\] vss 1.862896f
C1224 sarlogic_0/_050_ vss 0.622354f
C1225 sarlogic_0/_211_/a_36_160# vss 0.386641f
C1226 sarlogic_0/net4 vss 2.711508f
C1227 en vss 17.928204f
C1228 sarlogic_0/input4/a_36_68# vss 0.69549f
C1229 sarlogic_0/_426_/a_2560_156# vss 0.016968f
C1230 sarlogic_0/_426_/a_2665_112# vss 0.62251f
C1231 sarlogic_0/_426_/a_2248_156# vss 0.371662f
C1232 sarlogic_0/_426_/a_1204_472# vss 0.012971f
C1233 sarlogic_0/_426_/a_1000_472# vss 0.291735f
C1234 sarlogic_0/_426_/a_796_472# vss 0.023206f
C1235 sarlogic_0/_426_/a_1308_423# vss 0.279043f
C1236 sarlogic_0/_426_/a_448_472# vss 0.684413f
C1237 sarlogic_0/_426_/a_36_151# vss 1.43589f
C1238 sarlogic_0/_027_ vss 0.302949f
C1239 sarlogic_0/_150_ vss 0.320497f
C1240 sarlogic_0/FILLER_0_18_107/a_3172_472# vss 0.345058f
C1241 sarlogic_0/FILLER_0_18_107/a_2724_472# vss 0.33241f
C1242 sarlogic_0/FILLER_0_18_107/a_2276_472# vss 0.33241f
C1243 sarlogic_0/FILLER_0_18_107/a_1828_472# vss 0.33241f
C1244 sarlogic_0/FILLER_0_18_107/a_1380_472# vss 0.33241f
C1245 sarlogic_0/FILLER_0_18_107/a_932_472# vss 0.33241f
C1246 sarlogic_0/FILLER_0_18_107/a_484_472# vss 0.33241f
C1247 sarlogic_0/FILLER_0_18_107/a_36_472# vss 0.404746f
C1248 sarlogic_0/FILLER_0_18_107/a_3260_375# vss 0.233093f
C1249 sarlogic_0/FILLER_0_18_107/a_2812_375# vss 0.17167f
C1250 sarlogic_0/FILLER_0_18_107/a_2364_375# vss 0.17167f
C1251 sarlogic_0/FILLER_0_18_107/a_1916_375# vss 0.17167f
C1252 sarlogic_0/FILLER_0_18_107/a_1468_375# vss 0.17167f
C1253 sarlogic_0/FILLER_0_18_107/a_1020_375# vss 0.17167f
C1254 sarlogic_0/FILLER_0_18_107/a_572_375# vss 0.17167f
C1255 sarlogic_0/FILLER_0_18_107/a_124_375# vss 0.185915f
C1256 sarlogic_0/trim_mask\[4\] vss 0.987791f
C1257 sarlogic_0/_032_ vss 0.34876f
C1258 sarlogic_0/_443_/a_2560_156# vss 0.016968f
C1259 sarlogic_0/_443_/a_2665_112# vss 0.62251f
C1260 sarlogic_0/_443_/a_2248_156# vss 0.371662f
C1261 sarlogic_0/_443_/a_1204_472# vss 0.012971f
C1262 sarlogic_0/_443_/a_1000_472# vss 0.291735f
C1263 sarlogic_0/_443_/a_796_472# vss 0.023206f
C1264 sarlogic_0/_443_/a_1308_423# vss 0.279043f
C1265 sarlogic_0/_443_/a_448_472# vss 0.684413f
C1266 sarlogic_0/_443_/a_36_151# vss 1.43589f
C1267 sarlogic_0/_061_ vss 0.84986f
C1268 sarlogic_0/_056_ vss 2.393362f
C1269 sarlogic_0/_374_/a_36_68# vss 0.112263f
C1270 sarlogic_0/fanout58/a_36_160# vss 0.696445f
C1271 sarlogic_0/net74 vss 1.237373f
C1272 sarlogic_0/fanout69/a_36_113# vss 0.418095f
C1273 sarlogic_0/_173_ vss 0.339446f
C1274 sarlogic_0/FILLER_0_3_142/a_36_472# vss 0.417394f
C1275 sarlogic_0/FILLER_0_3_142/a_124_375# vss 0.246306f
C1276 sarlogic_0/FILLER_0_17_64/a_36_472# vss 0.417394f
C1277 sarlogic_0/FILLER_0_17_64/a_124_375# vss 0.246306f
C1278 sarlogic_0/FILLER_0_11_101/a_484_472# vss 0.345058f
C1279 sarlogic_0/FILLER_0_11_101/a_36_472# vss 0.404746f
C1280 sarlogic_0/FILLER_0_11_101/a_572_375# vss 0.232991f
C1281 sarlogic_0/FILLER_0_11_101/a_124_375# vss 0.185089f
C1282 sarlogic_0/FILLER_0_22_86/a_1380_472# vss 0.345058f
C1283 sarlogic_0/FILLER_0_22_86/a_932_472# vss 0.33241f
C1284 sarlogic_0/FILLER_0_22_86/a_484_472# vss 0.33241f
C1285 sarlogic_0/FILLER_0_22_86/a_36_472# vss 0.404746f
C1286 sarlogic_0/FILLER_0_22_86/a_1468_375# vss 0.233029f
C1287 sarlogic_0/FILLER_0_22_86/a_1020_375# vss 0.171606f
C1288 sarlogic_0/FILLER_0_22_86/a_572_375# vss 0.171606f
C1289 sarlogic_0/FILLER_0_22_86/a_124_375# vss 0.185399f
C1290 sarlogic_0/net24 vss 1.61895f
C1291 sarlogic_0/net3 vss 0.740676f
C1292 sarlogic_0/input3/a_36_113# vss 0.418095f
C1293 sarlogic_0/_103_ vss 0.350464f
C1294 sarlogic_0/_289_/a_36_472# vss 0.031137f
C1295 sarlogic_0/_151_ vss 0.300777f
C1296 sarlogic_0/_427_/a_2560_156# vss 0.016968f
C1297 sarlogic_0/_427_/a_2665_112# vss 0.91969f
C1298 sarlogic_0/_427_/a_2248_156# vss 0.30886f
C1299 sarlogic_0/_427_/a_1204_472# vss 0.012971f
C1300 sarlogic_0/_427_/a_1000_472# vss 0.291735f
C1301 sarlogic_0/_427_/a_796_472# vss 0.023206f
C1302 sarlogic_0/_427_/a_1308_423# vss 0.279043f
C1303 sarlogic_0/_427_/a_448_472# vss 0.684413f
C1304 sarlogic_0/_427_/a_36_151# vss 1.43587f
C1305 sarlogic_0/FILLER_0_17_161/a_36_472# vss 0.417394f
C1306 sarlogic_0/FILLER_0_17_161/a_124_375# vss 0.246306f
C1307 sarlogic_0/FILLER_0_18_139/a_1380_472# vss 0.345058f
C1308 sarlogic_0/FILLER_0_18_139/a_932_472# vss 0.33241f
C1309 sarlogic_0/FILLER_0_18_139/a_484_472# vss 0.33241f
C1310 sarlogic_0/FILLER_0_18_139/a_36_472# vss 0.404746f
C1311 sarlogic_0/FILLER_0_18_139/a_1468_375# vss 0.233029f
C1312 sarlogic_0/FILLER_0_18_139/a_1020_375# vss 0.171606f
C1313 sarlogic_0/FILLER_0_18_139/a_572_375# vss 0.171606f
C1314 sarlogic_0/FILLER_0_18_139/a_124_375# vss 0.185399f
C1315 sarlogic_0/_161_ vss 0.592909f
C1316 sarlogic_0/_162_ vss 0.597238f
C1317 sarlogic_0/_375_/a_36_68# vss 0.048026f
C1318 sarlogic_0/trim_val\[0\] vss 0.742779f
C1319 sarlogic_0/net67 vss 1.662327f
C1320 sarlogic_0/_444_/a_2560_156# vss 0.016968f
C1321 sarlogic_0/_444_/a_2665_112# vss 0.62251f
C1322 sarlogic_0/_444_/a_2248_156# vss 0.371662f
C1323 sarlogic_0/_444_/a_1204_472# vss 0.012971f
C1324 sarlogic_0/_444_/a_1000_472# vss 0.291735f
C1325 sarlogic_0/_444_/a_796_472# vss 0.023206f
C1326 sarlogic_0/_444_/a_1308_423# vss 0.279043f
C1327 sarlogic_0/_444_/a_448_472# vss 0.684413f
C1328 sarlogic_0/_444_/a_36_151# vss 1.43589f
C1329 sarlogic_0/net65 vss 0.804072f
C1330 sarlogic_0/fanout57/a_36_113# vss 0.418095f
C1331 sarlogic_0/fanout68/a_36_113# vss 0.418095f
C1332 sarlogic_0/FILLER_0_12_2/a_484_472# vss 0.345058f
C1333 sarlogic_0/FILLER_0_12_2/a_36_472# vss 0.404746f
C1334 sarlogic_0/FILLER_0_12_2/a_572_375# vss 0.232991f
C1335 sarlogic_0/FILLER_0_12_2/a_124_375# vss 0.185089f
C1336 sarlogic_0/net79 vss 1.584979f
C1337 sarlogic_0/fanout79/a_36_160# vss 0.386641f
C1338 sarlogic_0/_392_/a_36_68# vss 0.112263f
C1339 sarlogic_0/FILLER_0_13_228/a_36_472# vss 0.417394f
C1340 sarlogic_0/FILLER_0_13_228/a_124_375# vss 0.246306f
C1341 sarlogic_0/FILLER_0_13_206/a_36_472# vss 0.417394f
C1342 sarlogic_0/FILLER_0_13_206/a_124_375# vss 0.246306f
C1343 sarlogic_0/FILLER_0_20_177/a_1380_472# vss 0.345058f
C1344 sarlogic_0/FILLER_0_20_177/a_932_472# vss 0.33241f
C1345 sarlogic_0/FILLER_0_20_177/a_484_472# vss 0.33241f
C1346 sarlogic_0/FILLER_0_20_177/a_36_472# vss 0.404746f
C1347 sarlogic_0/FILLER_0_20_177/a_1468_375# vss 0.233029f
C1348 sarlogic_0/FILLER_0_20_177/a_1020_375# vss 0.171606f
C1349 sarlogic_0/FILLER_0_20_177/a_572_375# vss 0.171606f
C1350 sarlogic_0/FILLER_0_20_177/a_124_375# vss 0.185399f
C1351 sarlogic_0/_051_ vss 0.349381f
C1352 sarlogic_0/_213_/a_67_603# vss 0.345683f
C1353 sarlogic_0/net2 vss 0.461658f
C1354 sarlogic_0/input2/a_36_113# vss 0.418095f
C1355 sarlogic_0/_129_ vss 0.926508f
C1356 sarlogic_0/_131_ vss 1.734297f
C1357 sarlogic_0/_359_/a_36_488# vss 0.101145f
C1358 sarlogic_0/FILLER_0_11_64/a_36_472# vss 0.417394f
C1359 sarlogic_0/FILLER_0_11_64/a_124_375# vss 0.246306f
C1360 sarlogic_0/state\[2\] vss 0.607433f
C1361 sarlogic_0/net53 vss 4.483899f
C1362 sarlogic_0/_017_ vss 0.334329f
C1363 sarlogic_0/net70 vss 1.238296f
C1364 sarlogic_0/_428_/a_2560_156# vss 0.016968f
C1365 sarlogic_0/_428_/a_2665_112# vss 0.62251f
C1366 sarlogic_0/_428_/a_2248_156# vss 0.371662f
C1367 sarlogic_0/_428_/a_1204_472# vss 0.012971f
C1368 sarlogic_0/_428_/a_1000_472# vss 0.291735f
C1369 sarlogic_0/_428_/a_796_472# vss 0.023206f
C1370 sarlogic_0/_428_/a_1308_423# vss 0.279043f
C1371 sarlogic_0/_428_/a_448_472# vss 0.684413f
C1372 sarlogic_0/_428_/a_36_151# vss 1.43589f
C1373 sarlogic_0/FILLER_0_5_72/a_1380_472# vss 0.345058f
C1374 sarlogic_0/FILLER_0_5_72/a_932_472# vss 0.33241f
C1375 sarlogic_0/FILLER_0_5_72/a_484_472# vss 0.33241f
C1376 sarlogic_0/FILLER_0_5_72/a_36_472# vss 0.404746f
C1377 sarlogic_0/FILLER_0_5_72/a_1468_375# vss 0.233029f
C1378 sarlogic_0/FILLER_0_5_72/a_1020_375# vss 0.171606f
C1379 sarlogic_0/FILLER_0_5_72/a_572_375# vss 0.171606f
C1380 sarlogic_0/FILLER_0_5_72/a_124_375# vss 0.185399f
C1381 sarlogic_0/_376_/a_36_160# vss 0.386641f
C1382 sarlogic_0/trim_val\[1\] vss 0.683578f
C1383 sarlogic_0/_445_/a_2560_156# vss 0.016968f
C1384 sarlogic_0/_445_/a_2665_112# vss 0.62251f
C1385 sarlogic_0/_445_/a_2248_156# vss 0.371662f
C1386 sarlogic_0/_445_/a_1204_472# vss 0.012971f
C1387 sarlogic_0/_445_/a_1000_472# vss 0.291735f
C1388 sarlogic_0/_445_/a_796_472# vss 0.023206f
C1389 sarlogic_0/_445_/a_1308_423# vss 0.279043f
C1390 sarlogic_0/_445_/a_448_472# vss 0.684413f
C1391 sarlogic_0/_445_/a_36_151# vss 1.43589f
C1392 sarlogic_0/fanout67/a_36_160# vss 0.386641f
C1393 sarlogic_0/fanout56/a_36_113# vss 0.418095f
C1394 sarlogic_0/net78 vss 0.686263f
C1395 sarlogic_0/fanout78/a_36_113# vss 0.418095f
C1396 sarlogic_0/_174_ vss 0.979741f
C1397 sarlogic_0/FILLER_0_0_198/a_36_472# vss 0.417394f
C1398 sarlogic_0/FILLER_0_0_198/a_124_375# vss 0.246306f
C1399 sarlogic_0/FILLER_0_15_290/a_36_472# vss 0.417394f
C1400 sarlogic_0/FILLER_0_15_290/a_124_375# vss 0.246306f
C1401 sarlogic_0/FILLER_0_24_290/a_36_472# vss 0.417394f
C1402 sarlogic_0/FILLER_0_24_290/a_124_375# vss 0.246306f
C1403 sarlogic_0/FILLER_0_4_107/a_1380_472# vss 0.345058f
C1404 sarlogic_0/FILLER_0_4_107/a_932_472# vss 0.33241f
C1405 sarlogic_0/FILLER_0_4_107/a_484_472# vss 0.33241f
C1406 sarlogic_0/FILLER_0_4_107/a_36_472# vss 0.404746f
C1407 sarlogic_0/FILLER_0_4_107/a_1468_375# vss 0.233029f
C1408 sarlogic_0/FILLER_0_4_107/a_1020_375# vss 0.171606f
C1409 sarlogic_0/FILLER_0_4_107/a_572_375# vss 0.171606f
C1410 sarlogic_0/FILLER_0_4_107/a_124_375# vss 0.185399f
C1411 sarlogic_0/FILLER_0_7_104/a_1380_472# vss 0.345058f
C1412 sarlogic_0/FILLER_0_7_104/a_932_472# vss 0.33241f
C1413 sarlogic_0/FILLER_0_7_104/a_484_472# vss 0.33241f
C1414 sarlogic_0/FILLER_0_7_104/a_36_472# vss 0.404746f
C1415 sarlogic_0/FILLER_0_7_104/a_1468_375# vss 0.233029f
C1416 sarlogic_0/FILLER_0_7_104/a_1020_375# vss 0.171606f
C1417 sarlogic_0/FILLER_0_7_104/a_572_375# vss 0.171606f
C1418 sarlogic_0/FILLER_0_7_104/a_124_375# vss 0.185399f
C1419 sarlogic_0/_214_/a_36_160# vss 0.386641f
C1420 sarlogic_0/net1 vss 0.364811f
C1421 sarlogic_0/input1/a_36_113# vss 0.418095f
C1422 sarlogic_0/_429_/a_2560_156# vss 0.016968f
C1423 sarlogic_0/_429_/a_2665_112# vss 0.62251f
C1424 sarlogic_0/_429_/a_2248_156# vss 0.371662f
C1425 sarlogic_0/_429_/a_1204_472# vss 0.012971f
C1426 sarlogic_0/_429_/a_1000_472# vss 0.291735f
C1427 sarlogic_0/_429_/a_796_472# vss 0.023206f
C1428 sarlogic_0/_429_/a_1308_423# vss 0.279043f
C1429 sarlogic_0/_429_/a_448_472# vss 0.684413f
C1430 sarlogic_0/_429_/a_36_151# vss 1.43589f
C1431 sarlogic_0/_011_ vss 0.278979f
C1432 sarlogic_0/_377_/a_36_472# vss 0.031137f
C1433 sarlogic_0/fanout66/a_36_113# vss 0.418095f
C1434 sarlogic_0/_035_ vss 0.327801f
C1435 sarlogic_0/_446_/a_2560_156# vss 0.016968f
C1436 sarlogic_0/_446_/a_2665_112# vss 0.62251f
C1437 sarlogic_0/_446_/a_2248_156# vss 0.371662f
C1438 sarlogic_0/_446_/a_1204_472# vss 0.012971f
C1439 sarlogic_0/_446_/a_1000_472# vss 0.291735f
C1440 sarlogic_0/_446_/a_796_472# vss 0.023206f
C1441 sarlogic_0/_446_/a_1308_423# vss 0.279043f
C1442 sarlogic_0/_446_/a_448_472# vss 0.684413f
C1443 sarlogic_0/_446_/a_36_151# vss 1.43589f
C1444 sarlogic_0/fanout77/a_36_113# vss 0.418095f
C1445 sarlogic_0/FILLER_0_5_212/a_36_472# vss 0.417394f
C1446 sarlogic_0/FILLER_0_5_212/a_124_375# vss 0.246306f
C1447 sarlogic_0/fanout55/a_36_160# vss 0.696445f
C1448 sarlogic_0/_175_ vss 0.344159f
C1449 sarlogic_0/_394_/a_1936_472# vss 0.009918f
C1450 sarlogic_0/_394_/a_718_524# vss 0.005143f
C1451 sarlogic_0/_394_/a_56_524# vss 0.41096f
C1452 sarlogic_0/_394_/a_728_93# vss 0.654825f
C1453 sarlogic_0/_394_/a_1336_472# vss 0.316639f
C1454 sarlogic_0/FILLER_0_3_172/a_3172_472# vss 0.345058f
C1455 sarlogic_0/FILLER_0_3_172/a_2724_472# vss 0.33241f
C1456 sarlogic_0/FILLER_0_3_172/a_2276_472# vss 0.33241f
C1457 sarlogic_0/FILLER_0_3_172/a_1828_472# vss 0.33241f
C1458 sarlogic_0/FILLER_0_3_172/a_1380_472# vss 0.33241f
C1459 sarlogic_0/FILLER_0_3_172/a_932_472# vss 0.33241f
C1460 sarlogic_0/FILLER_0_3_172/a_484_472# vss 0.33241f
C1461 sarlogic_0/FILLER_0_3_172/a_36_472# vss 0.404746f
C1462 sarlogic_0/FILLER_0_3_172/a_3260_375# vss 0.233093f
C1463 sarlogic_0/FILLER_0_3_172/a_2812_375# vss 0.17167f
C1464 sarlogic_0/FILLER_0_3_172/a_2364_375# vss 0.17167f
C1465 sarlogic_0/FILLER_0_3_172/a_1916_375# vss 0.17167f
C1466 sarlogic_0/FILLER_0_3_172/a_1468_375# vss 0.17167f
C1467 sarlogic_0/FILLER_0_3_172/a_1020_375# vss 0.17167f
C1468 sarlogic_0/FILLER_0_3_172/a_572_375# vss 0.17167f
C1469 sarlogic_0/FILLER_0_3_172/a_124_375# vss 0.185915f
C1470 sarlogic_0/FILLER_0_17_72/a_3172_472# vss 0.345058f
C1471 sarlogic_0/FILLER_0_17_72/a_2724_472# vss 0.33241f
C1472 sarlogic_0/FILLER_0_17_72/a_2276_472# vss 0.33241f
C1473 sarlogic_0/FILLER_0_17_72/a_1828_472# vss 0.33241f
C1474 sarlogic_0/FILLER_0_17_72/a_1380_472# vss 0.33241f
C1475 sarlogic_0/FILLER_0_17_72/a_932_472# vss 0.33241f
C1476 sarlogic_0/FILLER_0_17_72/a_484_472# vss 0.33241f
C1477 sarlogic_0/FILLER_0_17_72/a_36_472# vss 0.404746f
C1478 sarlogic_0/FILLER_0_17_72/a_3260_375# vss 0.233093f
C1479 sarlogic_0/FILLER_0_17_72/a_2812_375# vss 0.17167f
C1480 sarlogic_0/FILLER_0_17_72/a_2364_375# vss 0.17167f
C1481 sarlogic_0/FILLER_0_17_72/a_1916_375# vss 0.17167f
C1482 sarlogic_0/FILLER_0_17_72/a_1468_375# vss 0.17167f
C1483 sarlogic_0/FILLER_0_17_72/a_1020_375# vss 0.17167f
C1484 sarlogic_0/FILLER_0_17_72/a_572_375# vss 0.17167f
C1485 sarlogic_0/FILLER_0_17_72/a_124_375# vss 0.185915f
C1486 sarlogic_0/FILLER_0_2_93/a_484_472# vss 0.345058f
C1487 sarlogic_0/FILLER_0_2_93/a_36_472# vss 0.404746f
C1488 sarlogic_0/FILLER_0_2_93/a_572_375# vss 0.232991f
C1489 sarlogic_0/FILLER_0_2_93/a_124_375# vss 0.185089f
C1490 sarlogic_0/FILLER_0_11_142/a_484_472# vss 0.345058f
C1491 sarlogic_0/FILLER_0_11_142/a_36_472# vss 0.404746f
C1492 sarlogic_0/FILLER_0_11_142/a_572_375# vss 0.232991f
C1493 sarlogic_0/FILLER_0_11_142/a_124_375# vss 0.185089f
C1494 sarlogic_0/net25 vss 1.803472f
C1495 sarlogic_0/_232_/a_67_603# vss 0.345683f
C1496 sarlogic_0/net35 vss 1.844415f
C1497 sarlogic_0/mask\[8\] vss 1.276233f
C1498 sarlogic_0/_301_/a_36_472# vss 0.031137f
C1499 sarlogic_0/_033_ vss 0.323682f
C1500 sarlogic_0/_165_ vss 0.331995f
C1501 sarlogic_0/FILLER_0_3_2/a_36_472# vss 0.417394f
C1502 sarlogic_0/FILLER_0_3_2/a_124_375# vss 0.246306f
C1503 sarlogic_0/trim_val\[3\] vss 0.719615f
C1504 sarlogic_0/_036_ vss 0.369206f
C1505 sarlogic_0/net68 vss 1.735004f
C1506 sarlogic_0/_447_/a_2560_156# vss 0.016968f
C1507 sarlogic_0/_447_/a_2665_112# vss 0.62251f
C1508 sarlogic_0/_447_/a_2248_156# vss 0.371662f
C1509 sarlogic_0/_447_/a_1204_472# vss 0.012971f
C1510 sarlogic_0/_447_/a_1000_472# vss 0.291735f
C1511 sarlogic_0/_447_/a_796_472# vss 0.023206f
C1512 sarlogic_0/_447_/a_1308_423# vss 0.279043f
C1513 sarlogic_0/_447_/a_448_472# vss 0.684413f
C1514 sarlogic_0/_447_/a_36_151# vss 1.43589f
C1515 sarlogic_0/FILLER_0_19_28/a_484_472# vss 0.345058f
C1516 sarlogic_0/FILLER_0_19_28/a_36_472# vss 0.404746f
C1517 sarlogic_0/FILLER_0_19_28/a_572_375# vss 0.232991f
C1518 sarlogic_0/FILLER_0_19_28/a_124_375# vss 0.185089f
C1519 sarlogic_0/fanout65/a_36_113# vss 0.418095f
C1520 sarlogic_0/fanout76/a_36_160# vss 0.386641f
C1521 sarlogic_0/net54 vss 5.456963f
C1522 sarlogic_0/fanout54/a_36_160# vss 0.696445f
C1523 sarlogic_0/FILLER_0_4_49/a_484_472# vss 0.345058f
C1524 sarlogic_0/FILLER_0_4_49/a_36_472# vss 0.404746f
C1525 sarlogic_0/FILLER_0_4_49/a_572_375# vss 0.232991f
C1526 sarlogic_0/FILLER_0_4_49/a_124_375# vss 0.185089f
C1527 sarlogic_0/_176_ vss 0.804011f
C1528 sarlogic_0/_085_ vss 2.280803f
C1529 sarlogic_0/_116_ vss 1.959915f
C1530 sarlogic_0/_395_/a_36_488# vss 0.101145f
C1531 sarlogic_0/FILLER_0_14_50/a_36_472# vss 0.417394f
C1532 sarlogic_0/FILLER_0_14_50/a_124_375# vss 0.246306f
C1533 sarlogic_0/FILLER_0_8_263/a_36_472# vss 0.417394f
C1534 sarlogic_0/FILLER_0_8_263/a_124_375# vss 0.246306f
C1535 sarlogic_0/FILLER_0_0_130/a_36_472# vss 0.417394f
C1536 sarlogic_0/FILLER_0_0_130/a_124_375# vss 0.246306f
C1537 sarlogic_0/FILLER_0_16_255/a_36_472# vss 0.417394f
C1538 sarlogic_0/FILLER_0_16_255/a_124_375# vss 0.246306f
C1539 sarlogic_0/FILLER_0_7_59/a_484_472# vss 0.345058f
C1540 sarlogic_0/FILLER_0_7_59/a_36_472# vss 0.404746f
C1541 sarlogic_0/FILLER_0_7_59/a_572_375# vss 0.232991f
C1542 sarlogic_0/FILLER_0_7_59/a_124_375# vss 0.185089f
C1543 sarlogic_0/output19/a_224_472# vss 2.38465f
C1544 sarlogic_0/FILLER_0_7_146/a_36_472# vss 0.417394f
C1545 sarlogic_0/FILLER_0_7_146/a_124_375# vss 0.246306f
C1546 sarlogic_0/_216_/a_67_603# vss 0.345683f
C1547 sarlogic_0/FILLER_0_15_116/a_484_472# vss 0.345058f
C1548 sarlogic_0/FILLER_0_15_116/a_36_472# vss 0.404746f
C1549 sarlogic_0/FILLER_0_15_116/a_572_375# vss 0.232991f
C1550 sarlogic_0/FILLER_0_15_116/a_124_375# vss 0.185089f
C1551 sarlogic_0/_063_ vss 0.370155f
C1552 sarlogic_0/_233_/a_36_160# vss 0.386641f
C1553 sarlogic_0/FILLER_0_21_28/a_3172_472# vss 0.345058f
C1554 sarlogic_0/FILLER_0_21_28/a_2724_472# vss 0.33241f
C1555 sarlogic_0/FILLER_0_21_28/a_2276_472# vss 0.33241f
C1556 sarlogic_0/FILLER_0_21_28/a_1828_472# vss 0.33241f
C1557 sarlogic_0/FILLER_0_21_28/a_1380_472# vss 0.33241f
C1558 sarlogic_0/FILLER_0_21_28/a_932_472# vss 0.33241f
C1559 sarlogic_0/FILLER_0_21_28/a_484_472# vss 0.33241f
C1560 sarlogic_0/FILLER_0_21_28/a_36_472# vss 0.404746f
C1561 sarlogic_0/FILLER_0_21_28/a_3260_375# vss 0.233093f
C1562 sarlogic_0/FILLER_0_21_28/a_2812_375# vss 0.17167f
C1563 sarlogic_0/FILLER_0_21_28/a_2364_375# vss 0.17167f
C1564 sarlogic_0/FILLER_0_21_28/a_1916_375# vss 0.17167f
C1565 sarlogic_0/FILLER_0_21_28/a_1468_375# vss 0.17167f
C1566 sarlogic_0/FILLER_0_21_28/a_1020_375# vss 0.17167f
C1567 sarlogic_0/FILLER_0_21_28/a_572_375# vss 0.17167f
C1568 sarlogic_0/FILLER_0_21_28/a_124_375# vss 0.185915f
C1569 sarlogic_0/_110_ vss 0.323912f
C1570 sarlogic_0/_379_/a_36_472# vss 0.031137f
C1571 sarlogic_0/trim_val\[4\] vss 0.662409f
C1572 sarlogic_0/net76 vss 1.454269f
C1573 sarlogic_0/_448_/a_2560_156# vss 0.016968f
C1574 sarlogic_0/_448_/a_2665_112# vss 0.62251f
C1575 sarlogic_0/_448_/a_2248_156# vss 0.371662f
C1576 sarlogic_0/_448_/a_1204_472# vss 0.012971f
C1577 sarlogic_0/_448_/a_1000_472# vss 0.291735f
C1578 sarlogic_0/_448_/a_796_472# vss 0.023206f
C1579 sarlogic_0/_448_/a_1308_423# vss 0.279043f
C1580 sarlogic_0/_448_/a_448_472# vss 0.684413f
C1581 sarlogic_0/_448_/a_36_151# vss 1.43589f
C1582 sarlogic_0/fanout64/a_36_160# vss 0.386641f
C1583 sarlogic_0/fanout75/a_36_113# vss 0.418095f
C1584 sarlogic_0/_250_/a_36_68# vss 0.69549f
C1585 sarlogic_0/net56 vss 0.843396f
C1586 sarlogic_0/fanout53/a_36_160# vss 0.696445f
C1587 sarlogic_0/_177_ vss 0.358286f
C1588 result2 vss 15.903303f
C1589 sarlogic_0/net29 vss 1.802718f
C1590 sarlogic_0/output29/a_224_472# vss 2.38465f
C1591 sarlogic_0/output18/a_224_472# vss 2.38465f
C1592 sarlogic_0/FILLER_0_14_181/a_36_472# vss 0.417394f
C1593 sarlogic_0/FILLER_0_14_181/a_124_375# vss 0.246306f
C1594 sarlogic_0/_052_ vss 0.569133f
C1595 sarlogic_0/_217_/a_36_160# vss 0.386641f
C1596 sarlogic_0/net44 vss 1.407054f
C1597 sarlogic_0/_303_/a_36_472# vss 0.031137f
C1598 sarlogic_0/en_co_clk vss 0.346872f
C1599 sarlogic_0/net55 vss 5.119958f
C1600 sarlogic_0/net72 vss 1.366255f
C1601 sarlogic_0/_449_/a_2560_156# vss 0.016968f
C1602 sarlogic_0/_449_/a_2665_112# vss 0.62251f
C1603 sarlogic_0/_449_/a_2248_156# vss 0.371662f
C1604 sarlogic_0/_449_/a_1204_472# vss 0.012971f
C1605 sarlogic_0/_449_/a_1000_472# vss 0.291735f
C1606 sarlogic_0/_449_/a_796_472# vss 0.023206f
C1607 sarlogic_0/_449_/a_1308_423# vss 0.279043f
C1608 sarlogic_0/_449_/a_448_472# vss 0.684413f
C1609 sarlogic_0/_449_/a_36_151# vss 1.43589f
C1610 sarlogic_0/fanout52/a_36_160# vss 0.696445f
C1611 sarlogic_0/net82 vss 0.706042f
C1612 sarlogic_0/fanout74/a_36_113# vss 0.418095f
C1613 sarlogic_0/FILLER_0_10_28/a_36_472# vss 0.417394f
C1614 sarlogic_0/FILLER_0_10_28/a_124_375# vss 0.246306f
C1615 sarlogic_0/mask\[0\] vss 2.242948f
C1616 sarlogic_0/_320_/a_36_472# vss 0.137725f
C1617 sarlogic_0/fanout63/a_36_160# vss 0.696445f
C1618 sarlogic_0/FILLER_0_14_81/a_36_472# vss 0.417394f
C1619 sarlogic_0/FILLER_0_14_81/a_124_375# vss 0.246306f
C1620 sarlogic_0/_397_/a_36_472# vss 0.031137f
C1621 sarlogic_0/FILLER_0_13_212/a_1380_472# vss 0.345058f
C1622 sarlogic_0/FILLER_0_13_212/a_932_472# vss 0.33241f
C1623 sarlogic_0/FILLER_0_13_212/a_484_472# vss 0.33241f
C1624 sarlogic_0/FILLER_0_13_212/a_36_472# vss 0.404746f
C1625 sarlogic_0/FILLER_0_13_212/a_1468_375# vss 0.233029f
C1626 sarlogic_0/FILLER_0_13_212/a_1020_375# vss 0.171606f
C1627 sarlogic_0/FILLER_0_13_212/a_572_375# vss 0.171606f
C1628 sarlogic_0/FILLER_0_13_212/a_124_375# vss 0.185399f
C1629 sarlogic_0/net39 vss 1.445128f
C1630 sarlogic_0/output39/a_224_472# vss 2.38465f
C1631 result1 vss 15.943958f
C1632 sarlogic_0/net28 vss 1.759728f
C1633 sarlogic_0/output28/a_224_472# vss 2.38465f
C1634 sarlogic_0/output17/a_224_472# vss 2.38465f
C1635 sarlogic_0/FILLER_0_16_37/a_36_472# vss 0.417394f
C1636 sarlogic_0/FILLER_0_16_37/a_124_375# vss 0.246306f
C1637 sarlogic_0/net26 vss 1.671545f
C1638 sarlogic_0/_064_ vss 0.581481f
C1639 sarlogic_0/trim_val\[2\] vss 0.65354f
C1640 sarlogic_0/trim_mask\[2\] vss 0.92551f
C1641 sarlogic_0/_235_/a_67_603# vss 0.345683f
C1642 sarlogic_0/_013_ vss 0.48783f
C1643 sarlogic_0/_111_ vss 0.369652f
C1644 sarlogic_0/FILLER_0_18_177/a_3172_472# vss 0.345058f
C1645 sarlogic_0/FILLER_0_18_177/a_2724_472# vss 0.33241f
C1646 sarlogic_0/FILLER_0_18_177/a_2276_472# vss 0.33241f
C1647 sarlogic_0/FILLER_0_18_177/a_1828_472# vss 0.33241f
C1648 sarlogic_0/FILLER_0_18_177/a_1380_472# vss 0.33241f
C1649 sarlogic_0/FILLER_0_18_177/a_932_472# vss 0.33241f
C1650 sarlogic_0/FILLER_0_18_177/a_484_472# vss 0.33241f
C1651 sarlogic_0/FILLER_0_18_177/a_36_472# vss 0.404746f
C1652 sarlogic_0/FILLER_0_18_177/a_3260_375# vss 0.233093f
C1653 sarlogic_0/FILLER_0_18_177/a_2812_375# vss 0.17167f
C1654 sarlogic_0/FILLER_0_18_177/a_2364_375# vss 0.17167f
C1655 sarlogic_0/FILLER_0_18_177/a_1916_375# vss 0.17167f
C1656 sarlogic_0/FILLER_0_18_177/a_1468_375# vss 0.17167f
C1657 sarlogic_0/FILLER_0_18_177/a_1020_375# vss 0.17167f
C1658 sarlogic_0/FILLER_0_18_177/a_572_375# vss 0.17167f
C1659 sarlogic_0/FILLER_0_18_177/a_124_375# vss 0.185915f
C1660 sarlogic_0/FILLER_0_18_100/a_36_472# vss 0.417394f
C1661 sarlogic_0/FILLER_0_18_100/a_124_375# vss 0.246306f
C1662 sarlogic_0/_073_ vss 0.953711f
C1663 sarlogic_0/_126_ vss 2.036767f
C1664 sarlogic_0/_069_ vss 2.034557f
C1665 sarlogic_0/_321_/a_170_472# vss 0.077257f
C1666 sarlogic_0/fanout51/a_36_113# vss 0.418095f
C1667 sarlogic_0/net62 vss 4.932099f
C1668 sarlogic_0/fanout62/a_36_160# vss 0.696445f
C1669 sarlogic_0/fanout73/a_36_113# vss 0.418095f
C1670 sarlogic_0/FILLER_0_19_47/a_484_472# vss 0.345058f
C1671 sarlogic_0/FILLER_0_19_47/a_36_472# vss 0.404746f
C1672 sarlogic_0/FILLER_0_19_47/a_572_375# vss 0.232991f
C1673 sarlogic_0/FILLER_0_19_47/a_124_375# vss 0.185089f
C1674 sarlogic_0/FILLER_0_14_91/a_484_472# vss 0.345058f
C1675 sarlogic_0/FILLER_0_14_91/a_36_472# vss 0.404746f
C1676 sarlogic_0/FILLER_0_14_91/a_572_375# vss 0.232991f
C1677 sarlogic_0/FILLER_0_14_91/a_124_375# vss 0.185089f
C1678 sarlogic_0/FILLER_0_10_214/a_36_472# vss 0.417394f
C1679 sarlogic_0/FILLER_0_10_214/a_124_375# vss 0.246306f
C1680 sarlogic_0/FILLER_0_10_247/a_36_472# vss 0.417394f
C1681 sarlogic_0/FILLER_0_10_247/a_124_375# vss 0.246306f
C1682 sarlogic_0/_178_ vss 1.252435f
C1683 sarlogic_0/_398_/a_36_113# vss 0.418095f
C1684 sarlogic_0/FILLER_0_16_241/a_36_472# vss 0.417394f
C1685 sarlogic_0/FILLER_0_16_241/a_124_375# vss 0.246306f
C1686 sarlogic_0/net38 vss 1.529392f
C1687 sarlogic_0/output38/a_224_472# vss 2.38465f
C1688 sarlogic_0/net16 vss 1.295744f
C1689 sarlogic_0/output16/a_224_472# vss 2.38465f
C1690 result0 vss 20.418947f
C1691 sarlogic_0/output27/a_224_472# vss 2.38465f
C1692 sarlogic_0/_219_/a_36_160# vss 0.386641f
C1693 sarlogic_0/FILLER_0_20_193/a_484_472# vss 0.345058f
C1694 sarlogic_0/FILLER_0_20_193/a_36_472# vss 0.404746f
C1695 sarlogic_0/FILLER_0_20_193/a_572_375# vss 0.232991f
C1696 sarlogic_0/FILLER_0_20_193/a_124_375# vss 0.185089f
C1697 sarlogic_0/_236_/a_36_160# vss 0.696445f
C1698 sarlogic_0/_112_ vss 0.308886f
C1699 sarlogic_0/_305_/a_36_159# vss 0.374116f
C1700 sarlogic_0/_074_ vss 1.813232f
C1701 sarlogic_0/_253_/a_36_68# vss 0.061249f
C1702 sarlogic_0/net50 vss 4.486121f
C1703 sarlogic_0/net52 vss 3.536016f
C1704 sarlogic_0/fanout50/a_36_160# vss 0.696445f
C1705 sarlogic_0/FILLER_0_10_37/a_36_472# vss 0.417394f
C1706 sarlogic_0/FILLER_0_10_37/a_124_375# vss 0.246306f
C1707 sarlogic_0/fanout72/a_36_113# vss 0.418095f
C1708 sarlogic_0/fanout61/a_36_113# vss 0.418095f
C1709 sarlogic_0/_128_ vss 0.447252f
C1710 sarlogic_0/_127_ vss 1.291729f
C1711 sarlogic_0/_322_/a_848_380# vss 0.40208f
C1712 sarlogic_0/_322_/a_124_24# vss 0.591898f
C1713 sarlogic_0/_088_ vss 0.457961f
C1714 sarlogic_0/_079_ vss 1.114894f
C1715 sarlogic_0/_087_ vss 0.601674f
C1716 sarlogic_0/_270_/a_36_472# vss 0.031137f
C1717 sarlogic_0/FILLER_0_4_123/a_36_472# vss 0.417394f
C1718 sarlogic_0/FILLER_0_4_123/a_124_375# vss 0.246306f
C1719 sarlogic_0/FILLER_0_17_218/a_484_472# vss 0.345058f
C1720 sarlogic_0/FILLER_0_17_218/a_36_472# vss 0.404746f
C1721 sarlogic_0/FILLER_0_17_218/a_572_375# vss 0.232991f
C1722 sarlogic_0/FILLER_0_17_218/a_124_375# vss 0.185089f
C1723 sarlogic_0/output37/a_224_472# vss 2.38465f
C1724 valid vss 20.613598f
C1725 sarlogic_0/net48 vss 1.219262f
C1726 sarlogic_0/output48/a_224_472# vss 2.38465f
C1727 sarlogic_0/net15 vss 1.447491f
C1728 sarlogic_0/output15/a_224_472# vss 2.38465f
C1729 sarlogic_0/output26/a_224_472# vss 2.38465f
C1730 sarlogic_0/FILLER_0_16_57/a_1380_472# vss 0.345058f
C1731 sarlogic_0/FILLER_0_16_57/a_932_472# vss 0.33241f
C1732 sarlogic_0/FILLER_0_16_57/a_484_472# vss 0.33241f
C1733 sarlogic_0/FILLER_0_16_57/a_36_472# vss 0.404746f
C1734 sarlogic_0/FILLER_0_16_57/a_1468_375# vss 0.233029f
C1735 sarlogic_0/FILLER_0_16_57/a_1020_375# vss 0.171606f
C1736 sarlogic_0/FILLER_0_16_57/a_572_375# vss 0.171606f
C1737 sarlogic_0/FILLER_0_16_57/a_124_375# vss 0.185399f
C1738 sarlogic_0/_306_/a_36_68# vss 0.69549f
C1739 sarlogic_0/_072_ vss 2.604301f
C1740 sarlogic_0/fanout82/a_36_113# vss 0.418095f
C1741 sarlogic_0/_015_ vss 0.406653f
C1742 sarlogic_0/_323_/a_36_113# vss 0.418095f
C1743 sarlogic_0/net60 vss 5.024503f
C1744 sarlogic_0/net61 vss 1.666523f
C1745 sarlogic_0/fanout60/a_36_160# vss 0.696445f
C1746 sarlogic_0/fanout71/a_36_113# vss 0.418095f
C1747 sarlogic_0/FILLER_0_6_239/a_36_472# vss 0.417394f
C1748 sarlogic_0/FILLER_0_6_239/a_124_375# vss 0.246306f
C1749 sarlogic_0/FILLER_0_4_99/a_36_472# vss 0.417394f
C1750 sarlogic_0/FILLER_0_4_99/a_124_375# vss 0.246306f
C1751 sarlogic_0/net57 vss 1.383718f
C1752 sarlogic_0/FILLER_0_10_256/a_36_472# vss 0.417394f
C1753 sarlogic_0/FILLER_0_10_256/a_124_375# vss 0.246306f
C1754 sarlogic_0/cal_itt\[3\] vss 1.854962f
C1755 sarlogic_0/_340_/a_36_160# vss 0.386641f
C1756 sarlogic_0/FILLER_0_4_177/a_484_472# vss 0.345058f
C1757 sarlogic_0/FILLER_0_4_177/a_36_472# vss 0.404746f
C1758 sarlogic_0/FILLER_0_4_177/a_572_375# vss 0.232991f
C1759 sarlogic_0/FILLER_0_4_177/a_124_375# vss 0.185089f
C1760 sarlogic_0/FILLER_0_4_144/a_484_472# vss 0.345058f
C1761 sarlogic_0/FILLER_0_4_144/a_36_472# vss 0.404746f
C1762 sarlogic_0/FILLER_0_4_144/a_572_375# vss 0.232991f
C1763 sarlogic_0/FILLER_0_4_144/a_124_375# vss 0.185089f
C1764 sarlogic_0/output14/a_224_472# vss 2.38465f
C1765 result9 vss 25.761324f
C1766 sarlogic_0/output36/a_224_472# vss 2.38465f
C1767 sarlogic_0/output47/a_224_472# vss 2.38465f
C1768 sarlogic_0/output25/a_224_472# vss 2.389677f
C1769 sarlogic_0/FILLER_0_12_136/a_1380_472# vss 0.345058f
C1770 sarlogic_0/FILLER_0_12_136/a_932_472# vss 0.33241f
C1771 sarlogic_0/FILLER_0_12_136/a_484_472# vss 0.33241f
C1772 sarlogic_0/FILLER_0_12_136/a_36_472# vss 0.404746f
C1773 sarlogic_0/FILLER_0_12_136/a_1468_375# vss 0.233029f
C1774 sarlogic_0/FILLER_0_12_136/a_1020_375# vss 0.171606f
C1775 sarlogic_0/FILLER_0_12_136/a_572_375# vss 0.171606f
C1776 sarlogic_0/FILLER_0_12_136/a_124_375# vss 0.185399f
C1777 sarlogic_0/FILLER_0_16_89/a_1380_472# vss 0.345058f
C1778 sarlogic_0/FILLER_0_16_89/a_932_472# vss 0.33241f
C1779 sarlogic_0/FILLER_0_16_89/a_484_472# vss 0.33241f
C1780 sarlogic_0/FILLER_0_16_89/a_36_472# vss 0.404746f
C1781 sarlogic_0/FILLER_0_16_89/a_1468_375# vss 0.233029f
C1782 sarlogic_0/FILLER_0_16_89/a_1020_375# vss 0.171606f
C1783 sarlogic_0/FILLER_0_16_89/a_572_375# vss 0.171606f
C1784 sarlogic_0/FILLER_0_16_89/a_124_375# vss 0.185399f
C1785 sarlogic_0/FILLER_0_21_125/a_484_472# vss 0.345058f
C1786 sarlogic_0/FILLER_0_21_125/a_36_472# vss 0.404746f
C1787 sarlogic_0/FILLER_0_21_125/a_572_375# vss 0.232991f
C1788 sarlogic_0/FILLER_0_21_125/a_124_375# vss 0.185089f
C1789 sarlogic_0/_238_/a_67_603# vss 0.345683f
C1790 sarlogic_0/_096_ vss 2.205532f
C1791 sarlogic_0/_093_ vss 1.893313f
C1792 sarlogic_0/FILLER_0_19_55/a_36_472# vss 0.417394f
C1793 sarlogic_0/FILLER_0_19_55/a_124_375# vss 0.246306f
C1794 sarlogic_0/net81 vss 1.738987f
C1795 sarlogic_0/fanout81/a_36_160# vss 0.386641f
C1796 sarlogic_0/_057_ vss 1.600886f
C1797 sarlogic_0/_255_/a_224_552# vss 1.31114f
C1798 sarlogic_0/net73 vss 1.058857f
C1799 sarlogic_0/fanout70/a_36_113# vss 0.418095f
C1800 sarlogic_0/_003_ vss 0.3064f
C1801 sarlogic_0/_089_ vss 0.36777f
C1802 sarlogic_0/_272_/a_36_472# vss 0.031137f
C1803 sarlogic_0/_187_ vss 0.311229f
C1804 sarlogic_0/_410_/a_36_68# vss 0.112263f
C1805 sarlogic_0/_141_ vss 1.249289f
C1806 sarlogic_0/mask\[3\] vss 1.26722f
C1807 sarlogic_0/_341_/a_49_472# vss 0.054843f
C1808 cal vss 17.663244f
C1809 sarlogic_0/FILLER_0_7_195/a_36_472# vss 0.417394f
C1810 sarlogic_0/FILLER_0_7_195/a_124_375# vss 0.246306f
C1811 sarlogic_0/FILLER_0_7_162/a_36_472# vss 0.417394f
C1812 sarlogic_0/FILLER_0_7_162/a_124_375# vss 0.246306f
C1813 sarlogic_0/output13/a_224_472# vss 2.391402f
C1814 sarlogic_0/FILLER_0_18_2/a_3172_472# vss 0.345058f
C1815 sarlogic_0/FILLER_0_18_2/a_2724_472# vss 0.33241f
C1816 sarlogic_0/FILLER_0_18_2/a_2276_472# vss 0.33241f
C1817 sarlogic_0/FILLER_0_18_2/a_1828_472# vss 0.33241f
C1818 sarlogic_0/FILLER_0_18_2/a_1380_472# vss 0.33241f
C1819 sarlogic_0/FILLER_0_18_2/a_932_472# vss 0.33241f
C1820 sarlogic_0/FILLER_0_18_2/a_484_472# vss 0.33241f
C1821 sarlogic_0/FILLER_0_18_2/a_36_472# vss 0.404746f
C1822 sarlogic_0/FILLER_0_18_2/a_3260_375# vss 0.233093f
C1823 sarlogic_0/FILLER_0_18_2/a_2812_375# vss 0.17167f
C1824 sarlogic_0/FILLER_0_18_2/a_2364_375# vss 0.17167f
C1825 sarlogic_0/FILLER_0_18_2/a_1916_375# vss 0.17167f
C1826 sarlogic_0/FILLER_0_18_2/a_1468_375# vss 0.17167f
C1827 sarlogic_0/FILLER_0_18_2/a_1020_375# vss 0.17167f
C1828 sarlogic_0/FILLER_0_18_2/a_572_375# vss 0.17167f
C1829 sarlogic_0/FILLER_0_18_2/a_124_375# vss 0.185915f
C1830 sarlogic_0/net46 vss 1.13395f
C1831 sarlogic_0/output46/a_224_472# vss 2.38465f
C1832 result8 vss 18.36624f
C1833 sarlogic_0/output35/a_224_472# vss 2.38465f
C1834 sarlogic_0/output24/a_224_472# vss 2.38465f
C1835 sarlogic_0/FILLER_0_8_107/a_36_472# vss 0.417394f
C1836 sarlogic_0/FILLER_0_8_107/a_124_375# vss 0.246306f
C1837 sarlogic_0/FILLER_0_12_124/a_36_472# vss 0.417394f
C1838 sarlogic_0/FILLER_0_12_124/a_124_375# vss 0.246306f
C1839 sarlogic_0/net41 vss 1.746759f
C1840 sarlogic_0/_065_ vss 0.523724f
C1841 sarlogic_0/_239_/a_36_160# vss 0.696445f
C1842 sarlogic_0/FILLER_0_1_98/a_36_472# vss 0.417394f
C1843 sarlogic_0/FILLER_0_1_98/a_124_375# vss 0.246306f
C1844 sarlogic_0/_115_ vss 1.281516f
C1845 sarlogic_0/_114_ vss 2.293579f
C1846 sarlogic_0/_308_/a_848_380# vss 0.40208f
C1847 sarlogic_0/_308_/a_124_24# vss 0.591898f
C1848 sarlogic_0/_256_/a_36_68# vss 0.063181f
C1849 sarlogic_0/FILLER_0_10_78/a_1380_472# vss 0.345058f
C1850 sarlogic_0/FILLER_0_10_78/a_932_472# vss 0.33241f
C1851 sarlogic_0/FILLER_0_10_78/a_484_472# vss 0.33241f
C1852 sarlogic_0/FILLER_0_10_78/a_36_472# vss 0.404746f
C1853 sarlogic_0/FILLER_0_10_78/a_1468_375# vss 0.233029f
C1854 sarlogic_0/FILLER_0_10_78/a_1020_375# vss 0.171606f
C1855 sarlogic_0/FILLER_0_10_78/a_572_375# vss 0.171606f
C1856 sarlogic_0/FILLER_0_10_78/a_124_375# vss 0.185399f
C1857 sarlogic_0/_130_ vss 0.304085f
C1858 sarlogic_0/net80 vss 1.375599f
C1859 sarlogic_0/fanout80/a_36_113# vss 0.418095f
C1860 sarlogic_0/net58 vss 5.308423f
C1861 sarlogic_0/_000_ vss 0.382358f
C1862 sarlogic_0/net75 vss 1.474299f
C1863 sarlogic_0/_411_/a_2560_156# vss 0.016968f
C1864 sarlogic_0/_411_/a_2665_112# vss 0.62251f
C1865 sarlogic_0/_411_/a_2248_156# vss 0.371662f
C1866 sarlogic_0/_411_/a_1204_472# vss 0.012971f
C1867 sarlogic_0/_411_/a_1000_472# vss 0.291735f
C1868 sarlogic_0/_411_/a_796_472# vss 0.023206f
C1869 sarlogic_0/_411_/a_1308_423# vss 0.279043f
C1870 sarlogic_0/_411_/a_448_472# vss 0.684413f
C1871 sarlogic_0/_411_/a_36_151# vss 1.43589f
C1872 sarlogic_0/state\[0\] vss 0.680109f
C1873 sarlogic_0/_273_/a_36_68# vss 0.69549f
C1874 sarlogic_0/_142_ vss 0.324372f
C1875 sarlogic_0/FILLER_0_9_223/a_484_472# vss 0.345058f
C1876 sarlogic_0/FILLER_0_9_223/a_36_472# vss 0.404746f
C1877 sarlogic_0/FILLER_0_9_223/a_572_375# vss 0.232991f
C1878 sarlogic_0/FILLER_0_9_223/a_124_375# vss 0.185089f
C1879 sarlogic_0/FILLER_0_4_197/a_1380_472# vss 0.345058f
C1880 sarlogic_0/FILLER_0_4_197/a_932_472# vss 0.33241f
C1881 sarlogic_0/FILLER_0_4_197/a_484_472# vss 0.33241f
C1882 sarlogic_0/FILLER_0_4_197/a_36_472# vss 0.404746f
C1883 sarlogic_0/FILLER_0_4_197/a_1468_375# vss 0.233029f
C1884 sarlogic_0/FILLER_0_4_197/a_1020_375# vss 0.171606f
C1885 sarlogic_0/FILLER_0_4_197/a_572_375# vss 0.171606f
C1886 sarlogic_0/FILLER_0_4_197/a_124_375# vss 0.185399f
C1887 sarlogic_0/FILLER_0_17_226/a_36_472# vss 0.417394f
C1888 sarlogic_0/FILLER_0_17_226/a_124_375# vss 0.246306f
C1889 sarlogic_0/FILLER_0_5_109/a_484_472# vss 0.345058f
C1890 sarlogic_0/FILLER_0_5_109/a_36_472# vss 0.404746f
C1891 sarlogic_0/FILLER_0_5_109/a_572_375# vss 0.232991f
C1892 sarlogic_0/FILLER_0_5_109/a_124_375# vss 0.185089f
C1893 sarlogic_0/output12/a_224_472# vss 2.38465f
C1894 result7 vss 17.357138f
C1895 sarlogic_0/net34 vss 1.724665f
C1896 sarlogic_0/output34/a_224_472# vss 2.38465f
C1897 sarlogic_0/net45 vss 1.12041f
C1898 sarlogic_0/output45/a_224_472# vss 2.38465f
C1899 sarlogic_0/output23/a_224_472# vss 2.390503f
C1900 sarlogic_0/FILLER_0_15_142/a_484_472# vss 0.345058f
C1901 sarlogic_0/FILLER_0_15_142/a_36_472# vss 0.404746f
C1902 sarlogic_0/FILLER_0_15_142/a_572_375# vss 0.232991f
C1903 sarlogic_0/FILLER_0_15_142/a_124_375# vss 0.185089f
C1904 sarlogic_0/_077_ vss 1.645892f
C1905 sarlogic_0/_075_ vss 0.374516f
C1906 sarlogic_0/_257_/a_36_472# vss 0.031137f
C1907 sarlogic_0/_326_/a_36_160# vss 0.696445f
C1908 sarlogic_0/_412_/a_2560_156# vss 0.016968f
C1909 sarlogic_0/_412_/a_2665_112# vss 0.62251f
C1910 sarlogic_0/_412_/a_2248_156# vss 0.371662f
C1911 sarlogic_0/_412_/a_1204_472# vss 0.012971f
C1912 sarlogic_0/_412_/a_1000_472# vss 0.291735f
C1913 sarlogic_0/_412_/a_796_472# vss 0.023206f
C1914 sarlogic_0/_412_/a_1308_423# vss 0.279043f
C1915 sarlogic_0/_412_/a_448_472# vss 0.684413f
C1916 sarlogic_0/_412_/a_36_151# vss 1.43589f
C1917 sarlogic_0/_091_ vss 1.841339f
C1918 sarlogic_0/_274_/a_36_68# vss 0.063181f
C1919 sarlogic_0/_143_ vss 0.329289f
C1920 sarlogic_0/mask\[4\] vss 1.300438f
C1921 sarlogic_0/_343_/a_49_472# vss 0.054843f
C1922 sarlogic_0/FILLER_0_13_65/a_36_472# vss 0.417394f
C1923 sarlogic_0/FILLER_0_13_65/a_124_375# vss 0.246306f
C1924 sarlogic_0/_360_/a_36_160# vss 0.386641f
C1925 sarlogic_0/FILLER_0_4_185/a_36_472# vss 0.417394f
C1926 sarlogic_0/FILLER_0_4_185/a_124_375# vss 0.246306f
C1927 sarlogic_0/FILLER_0_4_152/a_36_472# vss 0.417394f
C1928 sarlogic_0/FILLER_0_4_152/a_124_375# vss 0.246306f
C1929 sarlogic_0/_291_/a_36_160# vss 0.386641f
C1930 sarlogic_0/output9/a_224_472# vss 2.38465f
C1931 sarlogic_0/output11/a_224_472# vss 2.391497f
C1932 sarlogic_0/output44/a_224_472# vss 2.38465f
C1933 result6 vss 17.04347f
C1934 sarlogic_0/output33/a_224_472# vss 2.38465f
C1935 sarlogic_0/output22/a_224_472# vss 2.38465f
C1936 sarlogic_0/FILLER_0_8_127/a_36_472# vss 0.417394f
C1937 sarlogic_0/FILLER_0_8_127/a_124_375# vss 0.246306f
C1938 sarlogic_0/FILLER_0_8_138/a_36_472# vss 0.417394f
C1939 sarlogic_0/FILLER_0_8_138/a_124_375# vss 0.246306f
C1940 sarlogic_0/FILLER_0_21_133/a_36_472# vss 0.417394f
C1941 sarlogic_0/FILLER_0_21_133/a_124_375# vss 0.246306f
C1942 sarlogic_0/FILLER_0_24_130/a_36_472# vss 0.417394f
C1943 sarlogic_0/FILLER_0_24_130/a_124_375# vss 0.246306f
C1944 sarlogic_0/FILLER_0_18_171/a_36_472# vss 0.417394f
C1945 sarlogic_0/FILLER_0_18_171/a_124_375# vss 0.246306f
C1946 sarlogic_0/_258_/a_36_160# vss 0.386641f
C1947 sarlogic_0/_016_ vss 0.314121f
C1948 sarlogic_0/_327_/a_36_472# vss 0.031137f
C1949 sarlogic_0/_189_/a_67_603# vss 0.345683f
C1950 sarlogic_0/FILLER_0_24_63/a_36_472# vss 0.417394f
C1951 sarlogic_0/FILLER_0_24_63/a_124_375# vss 0.246306f
C1952 sarlogic_0/FILLER_0_24_96/a_36_472# vss 0.417394f
C1953 sarlogic_0/FILLER_0_24_96/a_124_375# vss 0.246306f
C1954 sarlogic_0/cal_itt\[2\] vss 1.473514f
C1955 sarlogic_0/_002_ vss 0.289553f
C1956 sarlogic_0/_413_/a_2560_156# vss 0.016968f
C1957 sarlogic_0/_413_/a_2665_112# vss 0.62251f
C1958 sarlogic_0/_413_/a_2248_156# vss 0.371662f
C1959 sarlogic_0/_413_/a_1204_472# vss 0.012971f
C1960 sarlogic_0/_413_/a_1000_472# vss 0.291735f
C1961 sarlogic_0/_413_/a_796_472# vss 0.023206f
C1962 sarlogic_0/_413_/a_1308_423# vss 0.279043f
C1963 sarlogic_0/_413_/a_448_472# vss 0.684413f
C1964 sarlogic_0/_413_/a_36_151# vss 1.43589f
C1965 sarlogic_0/_092_ vss 0.680239f
C1966 sarlogic_0/FILLER_0_7_72/a_3172_472# vss 0.345058f
C1967 sarlogic_0/FILLER_0_7_72/a_2724_472# vss 0.33241f
C1968 sarlogic_0/FILLER_0_7_72/a_2276_472# vss 0.33241f
C1969 sarlogic_0/FILLER_0_7_72/a_1828_472# vss 0.33241f
C1970 sarlogic_0/FILLER_0_7_72/a_1380_472# vss 0.33241f
C1971 sarlogic_0/FILLER_0_7_72/a_932_472# vss 0.33241f
C1972 sarlogic_0/FILLER_0_7_72/a_484_472# vss 0.33241f
C1973 sarlogic_0/FILLER_0_7_72/a_36_472# vss 0.404746f
C1974 sarlogic_0/FILLER_0_7_72/a_3260_375# vss 0.233093f
C1975 sarlogic_0/FILLER_0_7_72/a_2812_375# vss 0.17167f
C1976 sarlogic_0/FILLER_0_7_72/a_2364_375# vss 0.17167f
C1977 sarlogic_0/FILLER_0_7_72/a_1916_375# vss 0.17167f
C1978 sarlogic_0/FILLER_0_7_72/a_1468_375# vss 0.17167f
C1979 sarlogic_0/FILLER_0_7_72/a_1020_375# vss 0.17167f
C1980 sarlogic_0/FILLER_0_7_72/a_572_375# vss 0.17167f
C1981 sarlogic_0/FILLER_0_7_72/a_124_375# vss 0.185915f
C1982 sarlogic_0/_086_ vss 2.45259f
C1983 sarlogic_0/_119_ vss 1.237181f
C1984 sarlogic_0/net63 vss 5.362473f
C1985 sarlogic_0/_430_/a_2560_156# vss 0.016968f
C1986 sarlogic_0/_430_/a_2665_112# vss 0.62251f
C1987 sarlogic_0/_430_/a_2248_156# vss 0.371662f
C1988 sarlogic_0/_430_/a_1204_472# vss 0.012971f
C1989 sarlogic_0/_430_/a_1000_472# vss 0.291735f
C1990 sarlogic_0/_430_/a_796_472# vss 0.023206f
C1991 sarlogic_0/_430_/a_1308_423# vss 0.279043f
C1992 sarlogic_0/_430_/a_448_472# vss 0.684413f
C1993 sarlogic_0/_430_/a_36_151# vss 1.43589f
C1994 sarlogic_0/_292_/a_36_160# vss 0.386641f
C1995 sarlogic_0/output8/a_224_472# vss 2.38465f
C1996 sarlogic_0/output10/a_224_472# vss 2.38465f
C1997 result5 vss 16.794119f
C1998 sarlogic_0/net32 vss 1.789002f
C1999 sarlogic_0/output32/a_224_472# vss 2.38465f
C2000 sarlogic_0/output43/a_224_472# vss 2.38465f
C2001 sarlogic_0/output21/a_224_472# vss 2.39076f
C2002 sarlogic_0/_053_ vss 1.705161f
C2003 sarlogic_0/FILLER_0_16_107/a_484_472# vss 0.345058f
C2004 sarlogic_0/FILLER_0_16_107/a_36_472# vss 0.404746f
C2005 sarlogic_0/FILLER_0_16_107/a_572_375# vss 0.232991f
C2006 sarlogic_0/FILLER_0_16_107/a_124_375# vss 0.185089f
C2007 sarlogic_0/FILLER_0_3_204/a_36_472# vss 0.417394f
C2008 sarlogic_0/FILLER_0_3_204/a_124_375# vss 0.246306f
C2009 sarlogic_0/FILLER_0_9_28/a_3172_472# vss 0.345058f
C2010 sarlogic_0/FILLER_0_9_28/a_2724_472# vss 0.33241f
C2011 sarlogic_0/FILLER_0_9_28/a_2276_472# vss 0.33241f
C2012 sarlogic_0/FILLER_0_9_28/a_1828_472# vss 0.33241f
C2013 sarlogic_0/FILLER_0_9_28/a_1380_472# vss 0.33241f
C2014 sarlogic_0/FILLER_0_9_28/a_932_472# vss 0.33241f
C2015 sarlogic_0/FILLER_0_9_28/a_484_472# vss 0.33241f
C2016 sarlogic_0/FILLER_0_9_28/a_36_472# vss 0.404746f
C2017 sarlogic_0/FILLER_0_9_28/a_3260_375# vss 0.233093f
C2018 sarlogic_0/FILLER_0_9_28/a_2812_375# vss 0.17167f
C2019 sarlogic_0/FILLER_0_9_28/a_2364_375# vss 0.17167f
C2020 sarlogic_0/FILLER_0_9_28/a_1916_375# vss 0.17167f
C2021 sarlogic_0/FILLER_0_9_28/a_1468_375# vss 0.17167f
C2022 sarlogic_0/FILLER_0_9_28/a_1020_375# vss 0.17167f
C2023 sarlogic_0/FILLER_0_9_28/a_572_375# vss 0.17167f
C2024 sarlogic_0/FILLER_0_9_28/a_124_375# vss 0.185915f
C2025 sarlogic_0/_132_ vss 1.491425f
C2026 sarlogic_0/_328_/a_36_113# vss 0.418095f
C2027 sarlogic_0/_414_/a_2560_156# vss 0.016968f
C2028 sarlogic_0/_414_/a_2665_112# vss 0.62251f
C2029 sarlogic_0/_414_/a_2248_156# vss 0.371662f
C2030 sarlogic_0/_414_/a_1204_472# vss 0.012971f
C2031 sarlogic_0/_414_/a_1000_472# vss 0.291735f
C2032 sarlogic_0/_414_/a_796_472# vss 0.023206f
C2033 sarlogic_0/_414_/a_1308_423# vss 0.279043f
C2034 sarlogic_0/_414_/a_448_472# vss 0.684413f
C2035 sarlogic_0/_414_/a_36_151# vss 1.43589f
C2036 sarlogic_0/_276_/a_36_160# vss 0.386641f
C2037 sarlogic_0/_144_ vss 1.173846f
C2038 sarlogic_0/_345_/a_36_160# vss 0.386641f
C2039 sarlogic_0/_155_ vss 0.638535f
C2040 sarlogic_0/_020_ vss 0.316793f
C2041 sarlogic_0/_431_/a_2560_156# vss 0.016968f
C2042 sarlogic_0/_431_/a_2665_112# vss 0.62251f
C2043 sarlogic_0/_431_/a_2248_156# vss 0.371662f
C2044 sarlogic_0/_431_/a_1204_472# vss 0.012971f
C2045 sarlogic_0/_431_/a_1000_472# vss 0.291735f
C2046 sarlogic_0/_431_/a_796_472# vss 0.023206f
C2047 sarlogic_0/_431_/a_1308_423# vss 0.279043f
C2048 sarlogic_0/_431_/a_448_472# vss 0.684413f
C2049 sarlogic_0/_431_/a_36_151# vss 1.43589f
C2050 sarlogic_0/_105_ vss 1.21281f
C2051 sarlogic_0/_293_/a_36_472# vss 0.031137f
C2052 sarlogic_0/FILLER_0_5_128/a_484_472# vss 0.345058f
C2053 sarlogic_0/FILLER_0_5_128/a_36_472# vss 0.404746f
C2054 sarlogic_0/FILLER_0_5_128/a_572_375# vss 0.232991f
C2055 sarlogic_0/FILLER_0_5_128/a_124_375# vss 0.185089f
C2056 sarlogic_0/FILLER_0_5_117/a_36_472# vss 0.417394f
C2057 sarlogic_0/FILLER_0_5_117/a_124_375# vss 0.246306f
C2058 sarlogic_0/net7 vss 1.174913f
C2059 sarlogic_0/output7/a_224_472# vss 2.38465f
C2060 sarlogic_0/output42/a_224_472# vss 2.38465f
C2061 result4 vss 16.365028f
C2062 sarlogic_0/net31 vss 1.912935f
C2063 sarlogic_0/output31/a_224_472# vss 2.38465f
C2064 sarlogic_0/output20/a_224_472# vss 2.38465f
C2065 sarlogic_0/FILLER_0_16_73/a_484_472# vss 0.345058f
C2066 sarlogic_0/FILLER_0_16_73/a_36_472# vss 0.404746f
C2067 sarlogic_0/FILLER_0_16_73/a_572_375# vss 0.232991f
C2068 sarlogic_0/FILLER_0_16_73/a_124_375# vss 0.185089f
C2069 sarlogic_0/FILLER_0_21_142/a_484_472# vss 0.345058f
C2070 sarlogic_0/FILLER_0_21_142/a_36_472# vss 0.404746f
C2071 sarlogic_0/FILLER_0_21_142/a_572_375# vss 0.232991f
C2072 sarlogic_0/FILLER_0_21_142/a_124_375# vss 0.185089f
C2073 sarlogic_0/FILLER_0_15_150/a_36_472# vss 0.417394f
C2074 sarlogic_0/FILLER_0_15_150/a_124_375# vss 0.246306f
C2075 sarlogic_0/FILLER_0_19_125/a_36_472# vss 0.417394f
C2076 sarlogic_0/FILLER_0_19_125/a_124_375# vss 0.246306f
C2077 sarlogic_0/net10 vss 1.481359f
C2078 sarlogic_0/net20 vss 2.034189f
C2079 sarlogic_0/_277_/a_36_160# vss 0.386641f
C2080 sarlogic_0/net27 vss 2.023744f
C2081 sarlogic_0/_004_ vss 0.390107f
C2082 sarlogic_0/_415_/a_2560_156# vss 0.016968f
C2083 sarlogic_0/_415_/a_2665_112# vss 0.62251f
C2084 sarlogic_0/_415_/a_2248_156# vss 0.371662f
C2085 sarlogic_0/_415_/a_1204_472# vss 0.012971f
C2086 sarlogic_0/_415_/a_1000_472# vss 0.291735f
C2087 sarlogic_0/_415_/a_796_472# vss 0.023206f
C2088 sarlogic_0/_415_/a_1308_423# vss 0.279043f
C2089 sarlogic_0/_415_/a_448_472# vss 0.684413f
C2090 sarlogic_0/_415_/a_36_151# vss 1.43589f
C2091 sarlogic_0/mask\[5\] vss 1.334568f
C2092 sarlogic_0/_346_/a_49_472# vss 0.054843f
C2093 sarlogic_0/_028_ vss 0.386029f
C2094 sarlogic_0/_363_/a_36_68# vss 0.150048f
C2095 sarlogic_0/_021_ vss 0.316776f
C2096 sarlogic_0/_432_/a_2560_156# vss 0.016968f
C2097 sarlogic_0/_432_/a_2665_112# vss 0.62251f
C2098 sarlogic_0/_432_/a_2248_156# vss 0.371662f
C2099 sarlogic_0/_432_/a_1204_472# vss 0.012971f
C2100 sarlogic_0/_432_/a_1000_472# vss 0.291735f
C2101 sarlogic_0/_432_/a_796_472# vss 0.023206f
C2102 sarlogic_0/_432_/a_1308_423# vss 0.279043f
C2103 sarlogic_0/_432_/a_448_472# vss 0.684413f
C2104 sarlogic_0/_432_/a_36_151# vss 1.43589f
C2105 sarlogic_0/_008_ vss 0.423631f
C2106 sarlogic_0/_104_ vss 1.435764f
C2107 sarlogic_0/_106_ vss 0.378703f
C2108 sarlogic_0/FILLER_0_17_200/a_484_472# vss 0.345058f
C2109 sarlogic_0/FILLER_0_17_200/a_36_472# vss 0.404746f
C2110 sarlogic_0/FILLER_0_17_200/a_572_375# vss 0.232991f
C2111 sarlogic_0/FILLER_0_17_200/a_124_375# vss 0.185089f
C2112 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2113 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2114 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2115 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2116 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2117 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2118 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2119 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2120 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2121 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2122 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2123 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2124 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2125 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2126 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2127 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2128 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2129 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2130 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2131 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2132 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2133 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2134 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2135 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2136 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2137 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2138 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2139 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2140 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2141 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2142 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2143 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2144 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2145 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2146 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2147 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2148 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2149 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2150 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2151 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2152 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2153 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2154 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2155 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2156 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2157 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2158 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2159 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2160 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2161 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2162 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2163 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2164 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2165 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2166 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2167 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2168 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2169 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2170 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2171 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2172 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2173 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2174 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2175 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2176 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2177 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2178 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2179 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2180 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2181 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2182 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2183 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2184 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2185 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2186 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2187 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2188 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2189 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2190 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2191 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2192 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2193 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2194 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2195 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2196 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2197 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2198 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2199 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2200 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2201 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2202 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2203 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2204 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2205 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2206 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2207 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2208 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2209 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2210 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2211 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2212 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2213 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2214 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2215 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2216 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2217 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2218 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2219 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2220 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2221 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2222 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2223 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2224 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2225 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2226 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2227 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2228 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2229 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2230 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2231 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2232 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2233 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2234 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2235 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2236 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2237 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2238 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2239 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2240 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2241 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2242 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2243 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2244 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2245 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2246 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2247 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2248 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2249 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2250 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2251 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2252 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2253 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2254 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2255 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2256 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2257 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2258 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2259 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2260 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2261 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2262 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2263 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2264 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2265 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2266 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2267 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2268 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2269 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2270 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2271 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2272 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2273 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2274 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2275 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2276 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2277 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2278 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2279 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2280 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2281 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2282 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2283 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2284 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2285 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2286 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2287 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2288 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2289 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2290 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2291 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2292 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2293 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2294 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2295 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2296 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2297 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2298 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2299 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2300 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2301 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2302 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2303 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2304 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2305 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2306 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2307 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2308 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2309 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2310 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2311 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2312 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2313 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2314 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2315 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2316 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2317 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2318 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2319 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2320 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2321 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2322 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2323 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2324 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2325 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2326 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2327 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2328 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2329 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2330 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2331 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2332 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2333 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2334 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2335 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2336 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2337 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2338 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2339 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2340 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2341 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2342 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2343 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2344 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2345 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2346 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2347 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2348 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2349 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2350 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2351 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2352 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2353 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2354 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2355 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2356 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2357 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2358 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2359 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2360 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2361 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2362 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2363 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2364 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2365 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2366 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2367 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2368 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2369 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2370 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2371 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2372 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2373 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2374 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2375 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2376 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2377 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2378 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2379 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2380 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2381 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2382 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2383 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2384 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2385 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2386 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2387 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2388 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2389 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2390 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2391 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2392 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2393 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2394 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2395 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2396 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2397 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2398 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2399 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2400 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2401 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2402 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2403 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2404 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2405 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2406 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2407 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2408 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2409 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2410 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2411 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2412 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2413 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2414 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2415 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2416 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2417 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2418 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2419 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2420 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2421 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2422 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2423 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2424 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2425 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2426 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2427 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2428 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2429 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2430 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2431 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2432 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2433 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2434 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2435 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2436 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2437 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2438 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2439 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2440 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2441 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2442 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2443 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2444 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2445 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2446 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2447 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2448 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2449 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2450 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2451 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2452 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2453 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2454 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2455 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2456 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2457 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2458 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2459 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2460 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2461 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2462 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2463 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2464 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2465 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2466 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2467 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2468 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2469 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2470 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2471 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2472 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2473 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2474 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2475 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2476 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2477 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2478 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2479 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2480 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2481 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2482 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2483 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2484 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2485 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2486 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2487 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2488 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2489 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2490 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2491 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2492 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2493 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2494 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2495 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2496 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2497 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2498 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2499 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2500 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2501 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2502 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2503 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2504 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2505 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2506 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2507 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2508 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2509 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2510 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2511 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2512 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2513 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2514 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2515 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2516 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2517 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2518 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2519 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2520 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2521 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2522 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2523 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2524 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2525 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2526 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2527 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2528 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2529 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2530 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2531 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2532 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2533 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2534 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2535 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2536 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2537 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2538 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2539 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2540 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2541 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2542 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2543 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2544 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2545 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2546 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2547 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2548 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2549 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2550 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2551 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2552 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2553 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2554 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2555 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2556 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2557 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2558 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2559 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2560 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2561 mim_cap_boss_1/mim_cap1_0/mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2562 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2563 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2564 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2565 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2566 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2567 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2568 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2569 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2570 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2571 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2572 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2573 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2574 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_221/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2575 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_232/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2576 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2577 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2578 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2579 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2580 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2581 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2582 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2583 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2584 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2585 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2586 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2587 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2588 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_220/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2589 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2590 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_210/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2591 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2592 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2593 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2594 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2595 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2596 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2597 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2598 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2599 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2600 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2601 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_231/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2602 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2603 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2604 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2605 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2606 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2607 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2608 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2609 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2610 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_230/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2611 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2612 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2613 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2614 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2615 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2616 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2617 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2618 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2619 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2620 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2621 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2622 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2623 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2624 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2625 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2626 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2627 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2628 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2629 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2630 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2631 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2632 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2633 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2634 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2635 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2636 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2637 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2638 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2639 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_109/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2640 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2641 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2642 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2643 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2644 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2645 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2646 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_108/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2647 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_119/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2648 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2649 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2650 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2651 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2652 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2653 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2654 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2655 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_129/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2656 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_107/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2657 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_118/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2658 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2659 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2660 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2661 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2662 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2663 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2664 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2665 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2666 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_128/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2667 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_139/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2668 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_106/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2669 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_117/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2670 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2671 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2672 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2673 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2674 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2675 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2676 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2677 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2678 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2679 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_127/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2680 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_138/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2681 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_149/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2682 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_116/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2683 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_105/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2684 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2685 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2686 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2687 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2688 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_169/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2689 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2690 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2691 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2692 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2693 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2694 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_159/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2695 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_126/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2696 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_148/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2697 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_137/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2698 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_115/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2699 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_104/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2700 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2701 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2702 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2703 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2704 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2705 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2706 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2707 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2708 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2709 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2710 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2711 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2712 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_158/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2713 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_125/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2714 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_147/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2715 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_136/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2716 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_114/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2717 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_103/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2718 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2719 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2720 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2721 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2722 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2723 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2724 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2725 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2726 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2727 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_9/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2728 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2729 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2730 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2731 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2732 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2733 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2734 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2735 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_124/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2736 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_146/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2737 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_135/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2738 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_113/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2739 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_102/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2740 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_179/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2741 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2742 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2743 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_155/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2744 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2745 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2746 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2747 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2748 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2749 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2750 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2751 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2752 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_8/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2753 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_89/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2754 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_45/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2755 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_56/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2756 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_34/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2757 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_12/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2758 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_78/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2759 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_67/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2760 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_23/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2761 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_134/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2762 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_189/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2763 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_123/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2764 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_145/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2765 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_112/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2766 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_101/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2767 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_178/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2768 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_167/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2769 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2770 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2771 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2772 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2773 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2774 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2775 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2776 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_154/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2777 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2778 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2779 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_7/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2780 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_88/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2781 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_55/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2782 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_44/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2783 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_33/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2784 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_99/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2785 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_11/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2786 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_66/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2787 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_22/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2788 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_77/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2789 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_177/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2790 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_188/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2791 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_199/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2792 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_122/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2793 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_144/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2794 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_133/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2795 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_100/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2796 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_111/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2797 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_166/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2798 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2799 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2800 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2801 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2802 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2803 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2804 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2805 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2806 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2807 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_6/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2808 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_98/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2809 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_87/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2810 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_54/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2811 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_43/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2812 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_32/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2813 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_10/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2814 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_65/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2815 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_21/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2816 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_76/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2817 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_187/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2818 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_198/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2819 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_143/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2820 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_121/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2821 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_132/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2822 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_110/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2823 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_165/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2824 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_176/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2825 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2826 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2827 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2828 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2829 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2830 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2831 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2832 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_5/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2833 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_97/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2834 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_53/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2835 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_42/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2836 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_86/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2837 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_64/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2838 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_20/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2839 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_75/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2840 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_31/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2841 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_175/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2842 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_164/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2843 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_197/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2844 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_142/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2845 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_186/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2846 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_153/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2847 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_120/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2848 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_131/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2849 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2850 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2851 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2852 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2853 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2854 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2855 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2856 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_4/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2857 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_63/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2858 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_41/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2859 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_96/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2860 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_52/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2861 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_85/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2862 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_74/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2863 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_30/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2864 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_163/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2865 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_185/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2866 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_130/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2867 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_196/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2868 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_141/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2869 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_152/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2870 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_174/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2871 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2872 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2873 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_183/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2874 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2875 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2876 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2877 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_3/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2878 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_62/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2879 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_40/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2880 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_51/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2881 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_95/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2882 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_84/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2883 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_73/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2884 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_151/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2885 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_140/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2886 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_195/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2887 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_184/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2888 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_162/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2889 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_173/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2890 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2891 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2892 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2893 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2894 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2895 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_2/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2896 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_61/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2897 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_50/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2898 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_94/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2899 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_72/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2900 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_83/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2901 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_161/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2902 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_194/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2903 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_150/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2904 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_172/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2905 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2906 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2907 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2908 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_170/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2909 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_1/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2910 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_93/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2911 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_71/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2912 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_82/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2913 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_60/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2914 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_171/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2915 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_182/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2916 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_193/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2917 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_160/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2918 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2919 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2920 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2921 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_0/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2922 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_92/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2923 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_70/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2924 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_81/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2925 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_192/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2926 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_181/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2927 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2928 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_91/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2929 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_80/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2930 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_191/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2931 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_180/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2932 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_90/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2933 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2934 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_190/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2935 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2936 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2937 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_209/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2938 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2939 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2940 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2941 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_208/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2942 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_219/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2943 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_19/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2944 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2945 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2946 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2947 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2948 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_207/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2949 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_218/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2950 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_229/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2951 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_29/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2952 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_18/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2953 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2954 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2955 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2956 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_206/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2957 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_239/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2958 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_217/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2959 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_228/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2960 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_39/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2961 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_28/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2962 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_17/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2963 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2964 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2965 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_216/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2966 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_205/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2967 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_238/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2968 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_227/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2969 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_27/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2970 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_38/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2971 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_49/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2972 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_16/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2973 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2974 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2975 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_215/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2976 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_237/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2977 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_204/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2978 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_226/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2979 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_37/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2980 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_26/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2981 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_48/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2982 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_15/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2983 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_59/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2984 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2985 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2986 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_236/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2987 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_203/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2988 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_225/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2989 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_36/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2990 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_47/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2991 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_25/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2992 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_14/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2993 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_69/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2994 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_58/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2995 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_201/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2996 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_223/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2997 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_234/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2998 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_235/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C2999 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_202/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3000 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_224/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3001 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_35/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3002 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_46/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3003 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_24/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3004 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_13/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3005 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_79/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3006 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_57/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3007 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_68/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3008 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_211/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3009 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_200/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3010 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_222/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3011 mim_cap_boss_0/mim_cap1_0/mim_cap_30_30_flip_233/cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# vss 9.60519f
C3012 cmp_outn vss 4.515526f
C3013 comparator_0/trimb_0/n2 vss 1.980196f
C3014 comparator_0/trimb_0/n0 vss 0.677622f
C3015 comparator_0/trimb_0/n1 vss 0.716105f
C3016 comparator_0/trimb_0/n4 vss 4.186665f
C3017 comparator_0/ip vss -4.6307f
C3018 comparator_0/trimb_0/n3 vss 3.310455f
C3019 trimb0 vss 5.040359f
C3020 trimb3 vss 9.24535f
C3021 trimb1 vss 5.292398f
C3022 trimb2 vss 5.230265f
C3023 trimb4 vss 9.899878f
C3024 cmp_clkc vss 7.514944f
C3025 cmp_outp vss 5.193122f
C3026 comparator_0/trim_0/n4 vss 4.186665f
C3027 comparator_0/in vss -4.630677f
C3028 comparator_0/trim_0/n3 vss 3.310455f
C3029 comparator_0/trim_0/n2 vss 1.980196f
C3030 comparator_0/trim_0/n0 vss 0.677622f
C3031 comparator_0/trim_0/n1 vss 0.716105f
C3032 trim4 vss 9.866366f
C3033 trim1 vss 5.678721f
C3034 trim0 vss 4.946733f
C3035 trim2 vss 5.221713f
C3036 trim3 vss 10.704487f
C3037 comparator_0/diff vss 0.155718f
C3038 dacn_0/bootstrapped_sw$1_0/XM4$4_0/w_n2712_234# vss 1.968192f
C3039 vinn vss 34.380764f
C3040 dacn_0/bootstrapped_sw$1_0/vbsh vss 7.079245f
C3041 dacn_0/bootstrapped_sw$1_0/vbsl vss 8.446682f
C3042 dacn_0/bootstrapped_sw$1_0/enb vss 1.523612f
C3043 dacn_0/bootstrapped_sw$1_0/vs vss 0.065021f
C3044 sample vss 60.522945f
C3045 dacn_0/bootstrapped_sw$1_0/vg vss 1.1621f
C3046 ctln9 vss 7.919665f
C3047 dacn_0/inv_renketu$1_0/dummy$1_1/ZN vss 0.095951f
C3048 dacn_0/inv_renketu$1_0/dummy$1_1/I vss 0.604559f
C3049 ctln8 vss 8.606935f
C3050 dacn_0/inv_renketu$1_0/dummy$1_0/ZN vss 0.095951f
C3051 dacn_0/inv_renketu$1_0/dummy$1_0/I vss 0.604559f
C3052 ctln7 vss 8.370317f
C3053 ctln6 vss 8.535432f
C3054 ctln5 vss 8.783366f
C3055 ctln4 vss 11.40431f
C3056 ctln3 vss 15.672786f
C3057 ctln1 vss 22.054564f
C3058 dacn_0/inv_renketu$1_0/inv$1$1_9/VSS vss 2.848055f
C3059 dacn_0/inv_renketu$1_0/inv$1$1_9/VDD vss 2.113035f
C3060 ctln0 vss 11.169371f
C3061 dacn_0/inv_renketu$1_0/inv$1$1_9/VNW vss 14.066851f
C3062 ctln2 vss 17.726461f
C3063 dacn_0/ndum vss 13.878879f
C3064 dacn_0/n0 vss 16.631123f
C3065 dacn_0/n1 vss 17.119806f
C3066 dacn_0/n4 vss 39.311863f
C3067 dacn_0/n5 vss 47.33512f
C3068 dacn_0/n2 vss 30.111814f
C3069 dacn_0/n3 vss 33.594227f
C3070 dacn_0/n9 vss 14.292219f
C3071 cmp_vinn vss -0.682473p
C3072 dacn_0/n8 vss 39.909065f
C3073 dacn_0/n7 vss 56.191708f
C3074 dacn_0/n6 vss 52.976902f
C3075 dacp_0/inv_renketu_0/dummy_1/ZN vss 0.095951f
C3076 dacp_0/inv_renketu_0/dummy_1/I vss 0.604559f
C3077 dacp_0/inv_renketu_0/dummy_0/ZN vss 0.095951f
C3078 dacp_0/inv_renketu_0/dummy_0/I vss 0.604559f
C3079 ctlp8 vss 8.312423f
C3080 ctlp7 vss 7.94004f
C3081 ctlp6 vss 8.807449f
C3082 ctlp5 vss 8.561325f
C3083 ctlp4 vss 7.904063f
C3084 ctlp3 vss 15.988887f
C3085 ctlp1 vss 21.120407f
C3086 dacp_0/inv_renketu_0/inv$1_9/VSS vss 2.848055f
C3087 dacp_0/inv_renketu_0/inv$1_9/VDD vss 2.113035f
C3088 ctlp0 vss 10.240612f
C3089 dacp_0/inv_renketu_0/inv$1_9/VNW vss 14.066851f
C3090 ctlp2 vss 16.06865f
C3091 dacp_0/ndum vss 13.878879f
C3092 ctlp9 vss 7.20226f
C3093 dacp_0/n4 vss 39.311863f
C3094 dacp_0/n5 vss 47.33512f
C3095 dacp_0/n9 vss 14.292219f
C3096 cmp_vinp vss -0.682573p
C3097 dacp_0/n8 vss 39.909065f
C3098 dacp_0/n7 vss 56.191708f
C3099 dacp_0/n6 vss 52.976902f
C3100 dacp_0/n0 vss 16.631123f
C3101 dacp_0/n2 vss 30.111814f
C3102 dacp_0/n1 vss 17.119806f
C3103 dacp_0/n3 vss 33.594227f
C3104 dacp_0/bootstrapped_sw_0/vs vss 0.065021f
C3105 dacp_0/bootstrapped_sw_0/enb vss 1.523612f
C3106 dacp_0/bootstrapped_sw_0/XM4_0/w_n2712_234# vss 1.968192f
C3107 dacp_0/bootstrapped_sw_0/vbsh vss 7.079245f
C3108 dacp_0/bootstrapped_sw_0/vbsl vss 8.446682f
C3109 vinp vss 34.380108f
C3110 dacp_0/bootstrapped_sw_0/vg vss 1.1621f
C3111 buffer_0/inv$2_1/in vss 0.881074f
C3112 buffer_0/in vss 6.651137f
C3113 latch_0/x3_0/out vss 0.606965f
C3114 latch_0/XM3$5_0/a_n211_n1582# vss 0.069312f
C3115 latch_0/XM4$5_0/a_540_n1607# vss 0.069312f
C3116 latch_0/Qn vss 0.69036f
C3117 latch_0/x4_0/out vss 0.606901f
.ends

