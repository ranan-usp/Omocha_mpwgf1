* NGSPICE file created from latch.ext - technology: gf180mcuD

.subckt XM2_x4_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 G VSUBS 0.124686f
C2 w_n319_n356# VSUBS 1.48703f
.ends

.subckt XM1_x4_latch G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n302_n324# 0.365275f
.ends

.subckt x4_latch inv_out inv_in vdd vss
XXM2_x4_latch_0 inv_in inv_out vdd vdd vss XM2_x4_latch
XXM1_x4_latch_0 inv_in inv_out vss vss XM1_x4_latch
C0 vdd 0 1.6624f
C1 inv_out 0 0.399533f
C2 vss 0 0.289424f
C3 inv_in 0 0.606521f
.ends

.subckt XM2_x3_latch G D w_n319_n356# S VSUBS
X0 S G D w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 G VSUBS 0.124686f
C2 w_n319_n356# VSUBS 1.48703f
.ends

.subckt XM1_x3_latch G D a_n319_n324# S
X0 S G D a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n319_n324# 0.365275f
.ends

.subckt x3_latch inv_out vdd inv_in vss
XXM2_x3_latch_0 inv_in inv_out vdd vdd vss XM2_x3_latch
XXM1_x3_latch_0 inv_in inv_out vss vss XM1_x3_latch
C0 vdd 0 1.658401f
C1 vss 0 0.284019f
C2 inv_out 0 0.399533f
C3 inv_in 0 0.606521f
.ends

.subckt XM4_latch G D a_n319_n324# S a_n319_252#
X0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n319_n324# 0.365186f
.ends

.subckt XM2_x2_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186194f
C1 G VSUBS 0.124686f
C2 w_n319_n356# VSUBS 1.48655f
.ends

.subckt XM1_x2_latch G a_n320_n324# D a_n318_252# S
X0 D G S a_n320_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n320_n324# 0.365186f
.ends

.subckt x2_latch inv_out vdd inv_in XM1_x2_latch_0/a_n318_252# vss
XXM2_x2_latch_0 inv_in inv_out vdd vdd vss XM2_x2_latch
XXM1_x2_latch_0 inv_in vss inv_out XM1_x2_latch_0/a_n318_252# vss XM1_x2_latch
C0 vdd 0 1.678276f
C1 inv_out 0 0.40245f
C2 vss 0 0.292283f
C3 inv_in 0 0.607553f
.ends

.subckt XM3_latch G D a_n319_n324# S a_n319_252#
X0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n319_n324# 0.365186f
.ends

.subckt XM2_x1_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186194f
C1 G VSUBS 0.124686f
C2 w_n319_n356# VSUBS 1.48655f
.ends

.subckt XM1_x1_latch G D a_n318_n324# S
X0 D G S a_n318_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G a_n318_n324# 0.365186f
.ends

.subckt x1_latch inv_out inv_in vdd vss
XXM2_x1_latch_0 inv_in inv_out vdd vdd vss XM2_x1_latch
XXM1_x1_latch_0 inv_in inv_out vss vss XM1_x1_latch
C0 vdd 0 1.676557f
C1 inv_out 0 0.40245f
C2 vss 0 0.30318f
C3 inv_in 0 0.607553f
.ends

.subckt latch vss vdd Q Qn R S
Xx4_latch_0 XM3_latch_0/G S vdd vss x4_latch
Xx3_latch_0 XM4_latch_0/G vdd R vss x3_latch
XXM4_latch_0 XM4_latch_0/G Q vss vss vss XM4_latch
Xx2_latch_0 Qn vdd Q vss vss x2_latch
XXM3_latch_0 XM3_latch_0/G Qn vss vss vss XM3_latch
Xx1_latch_0 Q Qn vdd vss x1_latch
C0 vss XM4_latch_0/G 0.103577f
C1 XM3_latch_0/G vdd 0.186837f
C2 vss Qn 0.167238f
C3 vss Q 0.14016f
C4 Q Qn 0.886677f
C5 XM4_latch_0/G vdd 0.186732f
C6 vdd Qn 0.134494f
C7 vss XM3_latch_0/G 0.103577f
C8 Q vdd 0.457389f
C9 vdd 0 9.513767f
C10 Qn 0 0.887927f
C11 vss 0 1.296609f
C12 Q 0 0.846126f
C13 XM4_latch_0/G 0 0.717123f
C14 R 0 0.592286f
C15 XM3_latch_0/G 0 0.717027f
C16 S 0 0.592286f
.ends

