* NGSPICE file created from buffer.ext - technology: gf180mcuD

.subckt XM2_buffer_inv2 G D S
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM1_buffer_inv2 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt buffer_inv2 in vdd vss out
XXM2_buffer_inv2_0 in out vdd XM2_buffer_inv2
XXM1_buffer_inv2_0 in out vss XM1_buffer_inv2
.ends

.subckt XM1_buffer_inv1 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt buffer_inv1 in vdd vss out
XXM1_buffer_inv1_0 in out vss XM1_buffer_inv1
.ends

.subckt buffer middle out in vdd vss
Xbuffer_inv2_0 middle vdd vss out buffer_inv2
Xbuffer_inv1_0 in vdd vss middle buffer_inv1
.ends

