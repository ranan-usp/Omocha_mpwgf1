* NGSPICE file created from saradc.ext - technology: gf180mcuD

.subckt XM2_x4_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 D S 0.045397f
C2 G S 0.002389f
C3 D G 0.002389f
C4 w_n319_n356# S 0.019807f
C5 D w_n319_n356# 0.019528f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48703f
.ends

.subckt XM1_x4_latch G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 S D 0.038197f
C2 G D 0.002868f
C3 D a_n302_n324# 0.065984f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365275f
.ends

.subckt x4_latch inv_out inv_in vdd vss
XXM2_x4_latch_0 inv_in inv_out vdd vdd vss XM2_x4_latch
XXM1_x4_latch_0 inv_in inv_out vss vss XM1_x4_latch
C0 inv_out vdd 0.090362f
C1 vss inv_out 0.041091f
C2 vss vdd 0.042913f
C3 inv_in inv_out 0.075645f
C4 inv_in vdd 0.070585f
C5 inv_in vss 0.036044f
C6 vdd 0 1.6624f
C7 inv_out 0 0.399533f
C8 vss 0 0.289424f
C9 inv_in 0 0.606521f
.ends

.subckt XM2_x3_latch G D w_n319_n356# S VSUBS
X0 S G D w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 G S 0.002389f
C1 S w_n319_n356# 0.019807f
C2 D S 0.045397f
C3 G w_n319_n356# 0.186402f
C4 D G 0.002389f
C5 D w_n319_n356# 0.019528f
C6 S VSUBS 0.0454f
C7 D VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48703f
.ends

.subckt XM1_x3_latch G D a_n319_n324# S
X0 S G D a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D G 0.002868f
C1 S D 0.038197f
C2 S G 0.002868f
C3 S a_n319_n324# 0.066063f
C4 D a_n319_n324# 0.065984f
C5 G a_n319_n324# 0.365275f
.ends

.subckt x3_latch inv_out vdd inv_in vss
XXM2_x3_latch_0 inv_in inv_out vdd vdd vss XM2_x3_latch
XXM1_x3_latch_0 inv_in inv_out vss vss XM1_x3_latch
C0 vss vdd 0.041623f
C1 inv_out vdd 0.090362f
C2 inv_in vss 0.036044f
C3 inv_in inv_out 0.075645f
C4 vss inv_out 0.041091f
C5 inv_in vdd 0.070585f
C6 vdd 0 1.658401f
C7 vss 0 0.284019f
C8 inv_out 0 0.399533f
C9 inv_in 0 0.606521f
.ends

.subckt XM4_latch G D a_n319_n324# S a_n319_252#
X0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 S G 0.002868f
C2 S D 0.038197f
C3 D a_n319_n324# 0.065984f
C4 S a_n319_n324# 0.065984f
C5 G a_n319_n324# 0.365186f
.ends

.subckt XM2_x2_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 G D 0.002389f
C1 S G 0.002389f
C2 w_n319_n356# D 0.019528f
C3 w_n319_n356# S 0.019528f
C4 w_n319_n356# G 0.186194f
C5 S D 0.045397f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48655f
.ends

.subckt XM1_x2_latch G a_n320_n324# D a_n318_252# S
X0 D G S a_n320_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 S G 0.002868f
C2 S D 0.038197f
C3 D a_n320_n324# 0.065984f
C4 S a_n320_n324# 0.065984f
C5 G a_n320_n324# 0.365186f
.ends

.subckt x2_latch inv_out vdd inv_in XM1_x2_latch_0/a_n318_252# vss
XXM2_x2_latch_0 inv_in inv_out vdd vdd vss XM2_x2_latch
XXM1_x2_latch_0 inv_in vss inv_out XM1_x2_latch_0/a_n318_252# vss XM1_x2_latch
C0 vdd inv_in 0.070339f
C1 inv_out vdd 0.089967f
C2 vdd vss 0.040272f
C3 inv_out inv_in 0.075645f
C4 vss inv_in 0.034813f
C5 inv_out vss 0.038009f
C6 vdd 0 1.678276f
C7 inv_out 0 0.40245f
C8 vss 0 0.292283f
C9 inv_in 0 0.607553f
.ends

.subckt XM3_latch G D a_n319_n324# S a_n319_252#
X0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 S D 0.038197f
C2 G D 0.002868f
C3 D a_n319_n324# 0.065984f
C4 S a_n319_n324# 0.065984f
C5 G a_n319_n324# 0.365186f
.ends

.subckt XM2_x1_latch G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 G S 0.002389f
C1 S D 0.045397f
C2 G D 0.002389f
C3 w_n319_n356# S 0.019528f
C4 G w_n319_n356# 0.186194f
C5 w_n319_n356# D 0.019528f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48655f
.ends

.subckt XM1_x1_latch G D a_n318_n324# S
X0 D G S a_n318_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S D 0.038197f
C1 G D 0.002868f
C2 S G 0.002868f
C3 D a_n318_n324# 0.065984f
C4 S a_n318_n324# 0.065984f
C5 G a_n318_n324# 0.365186f
.ends

.subckt x1_latch inv_out inv_in vdd vss
XXM2_x1_latch_0 inv_in inv_out vdd vdd vss XM2_x1_latch
XXM1_x1_latch_0 inv_in inv_out vss vss XM1_x1_latch
C0 inv_out vdd 0.089967f
C1 inv_in inv_out 0.075645f
C2 vss vdd 0.042519f
C3 inv_in vss 0.034813f
C4 inv_in vdd 0.070339f
C5 inv_out vss 0.038009f
C6 vdd 0 1.676557f
C7 inv_out 0 0.40245f
C8 vss 0 0.30318f
C9 inv_in 0 0.607553f
.ends

.subckt latch Q Qn R S tutyuu1 tutyuu2 vdd vss
Xx4_latch_0 tutyuu1 S vdd vss x4_latch
Xx3_latch_0 tutyuu2 vdd R vss x3_latch
XXM4_latch_0 tutyuu2 Q vss vss vss XM4_latch
Xx2_latch_0 Qn vdd Q vss vss x2_latch
XXM3_latch_0 tutyuu1 Qn vss vss vss XM3_latch
Xx1_latch_0 Q Qn vdd vss x1_latch
C0 R tutyuu2 0.091043f
C1 Q tutyuu2 0.080738f
C2 vdd tutyuu1 0.186837f
C3 vdd Qn 0.134494f
C4 Qn tutyuu1 0.080688f
C5 vss vdd 0.035019f
C6 vss tutyuu1 0.103577f
C7 vdd S 0.069238f
C8 vss Qn 0.167238f
C9 R vdd 0.069238f
C10 tutyuu1 S 0.091043f
C11 Qn S 0.008621f
C12 vdd Q 0.457389f
C13 Q tutyuu1 0.04404f
C14 Q Qn 0.886677f
C15 vss S 0.034158f
C16 R vss 0.034158f
C17 vss Q 0.14016f
C18 vdd tutyuu2 0.186732f
C19 R Q 0.008667f
C20 Qn tutyuu2 0.043999f
C21 vss tutyuu2 0.103577f
C22 vdd 0 9.513767f
C23 Qn 0 0.887927f
C24 vss 0 1.296609f
C25 Q 0 0.846126f
C26 tutyuu2 0 0.717123f
C27 R 0 0.592286f
C28 tutyuu1 0 0.717027f
C29 S 0 0.592286f
.ends

.subckt XM1_inv2 VSUBS G D a_n319_n324# S
X0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n319_n324# 0.066063f
C4 S a_n319_n324# 0.065984f
C5 G a_n319_n324# 0.365275f
.ends

.subckt XM2_inv2 VSUBS G D S
X0 D G S VSUBS pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 S D 0.045397f
C1 G S 0.002389f
C2 G D 0.002389f
C3 D VSUBS 0.065207f
C4 S VSUBS 0.064928f
C5 G VSUBS 0.311088f
.ends

.subckt inv2 inv_out inv_in vss
XXM1_inv2_0 XM1_inv2_0/VSUBS inv_in inv_out vss vss XM1_inv2
XXM2_inv2_0 vss inv_in inv_out vss XM2_inv2
C0 inv_in vss 0.106611f
C1 inv_out inv_in 0.075645f
C2 inv_out vss 0.138038f
C3 inv_out 0 0.395231f
C4 vss 0 1.956022f
C5 inv_in 0 0.606537f
.ends

.subckt XM1_inv1 VSUBS G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S D 0.038197f
C1 G D 0.002868f
C2 S G 0.002868f
C3 D a_n302_n324# 0.065984f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365275f
.ends

.subckt XM2_inv1 VSUBS G D S
X0 D G S VSUBS pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 S G 0.002389f
C1 D S 0.045397f
C2 D G 0.002389f
C3 D VSUBS 0.064928f
C4 S VSUBS 0.065207f
C5 G VSUBS 0.311088f
.ends

.subckt inv1 inv_out inv_in vss
XXM1_inv1_0 XM1_inv1_0/VSUBS inv_in inv_out vss vss XM1_inv1
XXM2_inv1_0 vss inv_in inv_out vss XM2_inv1
C0 vss inv_out 0.131465f
C1 inv_in inv_out 0.075645f
C2 vss inv_in 0.106647f
C3 inv_out 0 0.399522f
C4 vss 0 1.951823f
C5 inv_in 0 0.606504f
.ends

.subckt buffer buf_in buf_out inv2_0/inv_in vss
Xinv2_0 buf_out inv2_0/inv_in vss inv2
Xinv1_0 inv2_0/inv_in buf_in vss inv1
C0 vss inv2_0/inv_in 0.215763f
C1 vss buf_out 0.067727f
C2 vss buf_in 0.095444f
C3 inv2_0/inv_in buf_out 0.153015f
C4 inv2_0/inv_in buf_in 0.110773f
C5 buf_in 0 0.674967f
C6 buf_out 0 0.447624f
C7 vss 0 3.711325f
C8 inv2_0/inv_in 0 0.832311f
.ends

.subckt inv_p VSS ZN I VDD VPW VNW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 I VDD 0.074838f
C1 VSS VDD 0.029045f
C2 VDD ZN 0.271625f
C3 I VSS 0.091531f
C4 I ZN 0.58604f
C5 VSS ZN 0.180794f
C6 VNW VDD 0.082022f
C7 I VNW 0.285482f
C8 VNW VSS 0.006277f
C9 VNW ZN 0.023676f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu_p inv_p_7/I inv_p_9/ZN inv_p_6/ZN inv_p_3/ZN inv_p_9/I inv_p_0/ZN
+ inv_p_0/I inv_p_2/I inv_p_10/I inv_p_4/I inv_p_8/ZN inv_p_2/ZN inv_p_5/ZN inv_p_6/I
+ inv_p_10/ZN inv_p_8/I inv_p_1/I inv_p_7/ZN inv_p_4/ZN inv_p_1/ZN inv_p_3/I vss inv_p_5/I
+ vdd
Xinv_p_0 vss inv_p_0/ZN inv_p_0/I vdd inv_p_0/VPW vdd vss inv_p
Xinv_p_1 vss inv_p_1/ZN inv_p_1/I vdd inv_p_1/VPW vdd vss inv_p
Xinv_p_2 vss inv_p_2/ZN inv_p_2/I vdd inv_p_2/VPW vdd vss inv_p
Xinv_p_3 vss inv_p_3/ZN inv_p_3/I vdd inv_p_3/VPW vdd vss inv_p
Xinv_p_4 vss inv_p_4/ZN inv_p_4/I vdd inv_p_4/VPW vdd vss inv_p
Xinv_p_5 vss inv_p_5/ZN inv_p_5/I vdd inv_p_5/VPW vdd vss inv_p
Xinv_p_6 vss inv_p_6/ZN inv_p_6/I vdd inv_p_6/VPW vdd vss inv_p
Xinv_p_7 vss inv_p_7/ZN inv_p_7/I vdd inv_p_7/VPW vdd vss inv_p
Xinv_p_8 vss inv_p_8/ZN inv_p_8/I vdd inv_p_8/VPW vdd vss inv_p
Xinv_p_9 vss inv_p_9/ZN inv_p_9/I vdd inv_p_9/VPW vdd vss inv_p
Xinv_p_10 vss inv_p_10/ZN inv_p_10/I vdd inv_p_10/VPW vdd vss inv_p
C0 inv_p_4/ZN inv_p_1/I 0.028928f
C1 vss inv_p_7/I 0.166388f
C2 vss inv_p_3/I 0.166388f
C3 vdd inv_p_2/I 0.035575f
C4 vss inv_p_0/I 0.170492f
C5 vdd inv_p_1/I 0.019437f
C6 inv_p_6/I inv_p_6/ZN 0.029333f
C7 vss inv_p_7/ZN 0.003326f
C8 inv_p_4/I inv_p_5/I 0.084161f
C9 vss inv_p_8/I 0.166388f
C10 vss inv_p_0/ZN 0.005399f
C11 vss inv_p_9/I 0.166388f
C12 vss inv_p_4/I 0.166388f
C13 inv_p_10/I inv_p_2/ZN 0.028928f
C14 inv_p_7/I vdd 0.019437f
C15 vdd inv_p_3/I 0.019437f
C16 vss inv_p_8/ZN 0.003326f
C17 vss inv_p_10/I 0.166388f
C18 vss inv_p_3/ZN 0.003326f
C19 inv_p_0/I vdd 0.026972f
C20 inv_p_4/ZN inv_p_4/I 0.029333f
C21 inv_p_1/I inv_p_3/I 0.084161f
C22 vss inv_p_9/ZN 0.003326f
C23 inv_p_4/I inv_p_5/ZN 0.028928f
C24 inv_p_10/ZN inv_p_2/ZN 0.080571f
C25 inv_p_7/ZN vdd 0.159176f
C26 vss inv_p_10/ZN 0.003326f
C27 vdd inv_p_8/I 0.019437f
C28 vdd inv_p_0/ZN 0.184001f
C29 inv_p_5/I inv_p_6/I 0.084161f
C30 vdd inv_p_9/I 0.019437f
C31 inv_p_4/I vdd 0.019437f
C32 inv_p_2/I inv_p_10/I 0.084161f
C33 vdd inv_p_8/ZN 0.159176f
C34 vdd inv_p_10/I 0.019437f
C35 inv_p_0/I inv_p_3/I 0.08416f
C36 vdd inv_p_3/ZN 0.159176f
C37 inv_p_4/I inv_p_1/I 0.084161f
C38 vss inv_p_6/I 0.166388f
C39 inv_p_5/I inv_p_6/ZN 0.028928f
C40 vdd inv_p_9/ZN 0.159176f
C41 inv_p_7/I inv_p_7/ZN 0.029333f
C42 inv_p_1/I inv_p_3/ZN 0.002086f
C43 vss inv_p_1/ZN 0.003326f
C44 inv_p_2/I inv_p_10/ZN 0.002086f
C45 inv_p_7/I inv_p_8/I 0.084161f
C46 inv_p_0/ZN inv_p_3/I 0.002086f
C47 vdd inv_p_10/ZN 0.159176f
C48 vss inv_p_6/ZN 0.003326f
C49 inv_p_0/I inv_p_0/ZN 0.029333f
C50 inv_p_6/I inv_p_5/ZN 0.002086f
C51 inv_p_4/ZN inv_p_1/ZN 0.080571f
C52 inv_p_7/ZN inv_p_8/I 0.002086f
C53 inv_p_7/I inv_p_8/ZN 0.028928f
C54 inv_p_3/ZN inv_p_3/I 0.029333f
C55 inv_p_6/ZN inv_p_5/ZN 0.080571f
C56 vdd inv_p_6/I 0.019437f
C57 inv_p_0/I inv_p_3/ZN 0.028928f
C58 inv_p_8/I inv_p_9/I 0.084161f
C59 inv_p_7/ZN inv_p_8/ZN 0.080571f
C60 vdd inv_p_1/ZN 0.159176f
C61 inv_p_8/I inv_p_8/ZN 0.029333f
C62 inv_p_0/ZN inv_p_3/ZN 0.080571f
C63 vdd inv_p_6/ZN 0.159176f
C64 inv_p_1/I inv_p_1/ZN 0.029333f
C65 inv_p_8/I inv_p_9/ZN 0.028928f
C66 inv_p_8/ZN inv_p_9/I 0.002086f
C67 inv_p_10/I inv_p_9/I 0.084161f
C68 inv_p_9/I inv_p_9/ZN 0.029333f
C69 vss inv_p_5/I 0.166388f
C70 inv_p_7/I inv_p_6/I 0.084161f
C71 inv_p_8/ZN inv_p_9/ZN 0.080571f
C72 inv_p_10/I inv_p_9/ZN 0.002086f
C73 inv_p_10/ZN inv_p_9/I 0.028928f
C74 inv_p_1/ZN inv_p_3/I 0.028928f
C75 vss inv_p_2/ZN 0.005014f
C76 inv_p_4/ZN inv_p_5/I 0.002086f
C77 inv_p_10/I inv_p_10/ZN 0.029333f
C78 inv_p_7/ZN inv_p_6/I 0.028928f
C79 inv_p_7/I inv_p_6/ZN 0.002086f
C80 inv_p_5/I inv_p_5/ZN 0.029333f
C81 inv_p_10/ZN inv_p_9/ZN 0.080571f
C82 vss inv_p_4/ZN 0.003326f
C83 inv_p_7/ZN inv_p_6/ZN 0.080571f
C84 vss inv_p_5/ZN 0.003326f
C85 vdd inv_p_5/I 0.019437f
C86 inv_p_4/I inv_p_1/ZN 0.002086f
C87 inv_p_2/I inv_p_2/ZN 0.029333f
C88 vdd inv_p_2/ZN 0.174722f
C89 inv_p_4/ZN inv_p_5/ZN 0.080571f
C90 vss inv_p_2/I 0.164788f
C91 inv_p_1/ZN inv_p_3/ZN 0.080571f
C92 vss vdd 0.009518f
C93 vss inv_p_1/I 0.166388f
C94 inv_p_4/ZN vdd 0.159176f
C95 vdd inv_p_5/ZN 0.159176f
C96 inv_p_10/ZN 0 0.131999f
C97 inv_p_10/I 0 0.64919f
C98 inv_p_9/ZN 0 0.131999f
C99 inv_p_9/I 0 0.64919f
C100 inv_p_8/ZN 0 0.131999f
C101 inv_p_8/I 0 0.64919f
C102 inv_p_7/ZN 0 0.131999f
C103 inv_p_7/I 0 0.64919f
C104 inv_p_6/ZN 0 0.131999f
C105 inv_p_6/I 0 0.64919f
C106 inv_p_5/ZN 0 0.131999f
C107 inv_p_5/I 0 0.64919f
C108 inv_p_4/ZN 0 0.131999f
C109 inv_p_4/I 0 0.64919f
C110 inv_p_3/ZN 0 0.131999f
C111 inv_p_3/I 0 0.64919f
C112 vss 0 3.02573f
C113 inv_p_2/ZN 0 0.206166f
C114 vdd 0 16.013325f
C115 inv_p_2/I 0 0.750024f
C116 inv_p_1/ZN 0 0.131999f
C117 inv_p_1/I 0 0.64919f
C118 inv_p_0/ZN 0 0.209411f
C119 inv_p_0/I 0 0.731246f
.ends

.subckt XM3_bs_p G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 G S 0.002389f
C1 D S 0.045397f
C2 D G 0.002389f
C3 w_n319_n356# S 0.021189f
C4 w_n319_n356# G 0.186402f
C5 D w_n319_n356# 0.019807f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMs2_bs_p G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D S 0.038197f
C2 D G 0.002868f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.068446f
C5 G a_n302_n324# 0.365186f
.ends

.subckt XM2_bs_inv_p G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 G S 0.002389f
C1 D S 0.045397f
C2 D G 0.002389f
C3 w_n319_n356# S 0.019807f
C4 w_n319_n356# G 0.186609f
C5 D w_n319_n356# 0.019807f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48751f
.ends

.subckt XM1_bs_inv_p G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S D 0.038197f
C1 G D 0.002868f
C2 G S 0.002868f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365365f
.ends

.subckt bs_inv_p inv_out vdd inv_in vss
XXM2_bs_inv_p_0 inv_in inv_out vdd vdd vss XM2_bs_inv_p
XXM1_bs_inv_p_0 inv_in inv_out vss vss XM1_bs_inv_p
C0 vss inv_in 0.037258f
C1 inv_out vdd 0.092565f
C2 inv_in vdd 0.07083f
C3 vss vdd 0.043239f
C4 inv_out inv_in 0.075645f
C5 inv_out vss 0.04895f
C6 vdd 0 1.650725f
C7 inv_out 0 0.392313f
C8 vss 0 0.277512f
C9 inv_in 0 0.605506f
.ends

.subckt XM4_bs_p G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 w_n319_n356# S 0.021189f
C2 w_n319_n356# D 0.019807f
C3 G S 0.002389f
C4 D G 0.002389f
C5 D S 0.045397f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt bs_cap_p I1_1_1_R0_BOT I1_1_1_R0_TOP VSUBS
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.339999u c_length=12.339999u
C0 I1_1_1_R0_BOT I1_1_1_R0_TOP 0.730455f
C1 I1_1_1_R0_TOP VSUBS 2.59113f
C2 I1_1_1_R0_BOT VSUBS 1.76085f
.ends

.subckt XMs_bs_p G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 G D 0.002868f
C2 S D 0.038197f
C3 D a_n302_n324# 0.061336f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361785f
.ends

.subckt XM1_bs_p G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM2_bs_p G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XMs1_bs_p G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 G D 0.002868f
C2 S D 0.038197f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365275f
.ends

.subckt bootstrapped_sw_p vdd en enb bs_in bs_out vg vs vbsh vbsl vss
XXM3_bs_p_0 enb vg vbsh vbsh vss XM3_bs_p
XXMs2_bs_p_0 enb vss vss vss vs XMs2_bs_p
Xbs_inv_p_0 enb vdd en vss bs_inv_p
XXM4_bs_p_0 vg vdd vbsh vbsh vss XM4_bs_p
Xbs_cap_p_0 vbsl vbsh vss bs_cap_p
Xbs_cap_p_1 vbsl vbsh vss bs_cap_p
Xbs_cap_p_2 vbsl vbsh vss bs_cap_p
Xbs_cap_p_3 vbsl vbsh vss bs_cap_p
Xbs_cap_p_4 vbsl vbsh vss bs_cap_p
XXMs_bs_p_0 vg bs_out vss bs_in XMs_bs_p
XXM1_bs_p_0 vg vbsl vss vss bs_in XM1_bs_p
XXM2_bs_p_0 enb vbsl vss vss vss XM2_bs_p
XXMs1_bs_p_0 vdd vs vss vg XMs1_bs_p
C0 vs enb 0.00173f
C1 enb bs_out 0.001285f
C2 vdd enb 0.426791f
C3 vg bs_in 0.079028f
C4 vdd bs_out 0.008497f
C5 vbsl enb 0.01529f
C6 en enb 0.018916f
C7 vbsl bs_out 0.057454f
C8 enb vbsh 0.0922f
C9 vbsl vdd 0.002507f
C10 vdd en 0.086628f
C11 vbsh bs_out 0.119559f
C12 vdd vbsh 0.205818f
C13 vs vg 0.007099f
C14 enb vg 0.583075f
C15 vbsl vbsh 0.870275f
C16 vg bs_out 0.066304f
C17 vdd vg 0.500479f
C18 vbsl vg 0.043332f
C19 en vg 0.002156f
C20 vbsl bs_in 0.256003f
C21 vg vbsh 0.283904f
C22 vbsh bs_in 0.013047f
C23 vs vss 0.042967f
C24 enb vss 1.703464f
C25 bs_out vss 0.895635f
C26 bs_in vss 0.389944f
C27 vg vss 1.576155f
C28 vbsh vss 14.292329f
C29 vbsl vss 8.158694f
C30 vdd vss 3.558326f
C31 en vss 0.896531f
.ends

.subckt dacp dac_in dum ctl7 ctl8 ctl9 ctl10 sample ctl2 ctl1 carray_p_0/n0 carray_p_0/ndum
+ ctl4 ctl6 bootstrapped_sw_p_0/enb dac_out ctl3 bootstrapped_sw_p_0/vg carray_p_0/n8
+ carray_p_0/n9 ctl5 carray_p_0/n7 vdd bootstrapped_sw_p_0/vbsh vss bootstrapped_sw_p_0/vbsl
Xinv_renketu_p_0 ctl6 carray_p_0/n8 carray_p_0/n5 carray_p_0/n1 ctl8 carray_p_0/ndum
+ dum ctl10 ctl9 ctl3 carray_p_0/n7 carray_p_0/n0 carray_p_0/n4 ctl5 carray_p_0/n9
+ ctl7 ctl2 carray_p_0/n6 carray_p_0/n3 carray_p_0/n2 ctl1 vss ctl4 vdd inv_renketu_p
Xbootstrapped_sw_p_0 vdd sample bootstrapped_sw_p_0/enb dac_in dac_out bootstrapped_sw_p_0/vg
+ bootstrapped_sw_p_0/vs bootstrapped_sw_p_0/vbsh bootstrapped_sw_p_0/vbsl vss bootstrapped_sw_p
C0 dac_out carray_p_0/n5 52.565514f
C1 carray_p_0/n0 carray_p_0/n5 0.025424f
C2 carray_p_0/n6 carray_p_0/n3 0.336612f
C3 ctl6 ctl5 0.104537f
C4 carray_p_0/n0 vdd 0.002151f
C5 carray_p_0/n8 carray_p_0/n7 50.51461f
C6 carray_p_0/n5 vdd 0.002151f
C7 carray_p_0/ndum carray_p_0/n2 0.041162f
C8 carray_p_0/n4 carray_p_0/n3 26.229403f
C9 carray_p_0/n9 carray_p_0/n3 1.911224f
C10 carray_p_0/n8 carray_p_0/n6 11.2161f
C11 dum ctl1 0.104537f
C12 carray_p_0/n1 carray_p_0/ndum 8.498201f
C13 carray_p_0/n7 carray_p_0/n2 0.485355f
C14 dac_out carray_p_0/n3 13.201303f
C15 ctl7 ctl6 0.104537f
C16 carray_p_0/n0 carray_p_0/n3 0.051666f
C17 ctl3 ctl4 0.104537f
C18 carray_p_0/n8 carray_p_0/n9 87.43918f
C19 carray_p_0/n8 carray_p_0/n4 2.84323f
C20 carray_p_0/n1 carray_p_0/n7 0.212822f
C21 ctl5 ctl4 0.104537f
C22 ctl9 ctl8 0.104537f
C23 carray_p_0/n5 carray_p_0/n3 0.346757f
C24 dac_out bootstrapped_sw_p_0/vbsh 0.280658f
C25 carray_p_0/n6 carray_p_0/n2 0.20799f
C26 vdd carray_p_0/n3 0.002151f
C27 carray_p_0/n8 dac_out 0.420151p
C28 sample carray_p_0/ndum 0.045492f
C29 carray_p_0/n8 carray_p_0/n0 0.097254f
C30 ctl10 ctl9 0.104537f
C31 carray_p_0/n6 carray_p_0/n1 0.142211f
C32 carray_p_0/n9 carray_p_0/n2 0.996681f
C33 carray_p_0/n4 carray_p_0/n2 0.213209f
C34 carray_p_0/n8 carray_p_0/n5 5.60732f
C35 carray_p_0/n7 carray_p_0/ndum 0.06073f
C36 carray_p_0/n8 vdd 0.002151f
C37 ctl2 ctl1 0.104537f
C38 carray_p_0/n1 carray_p_0/n4 0.142475f
C39 carray_p_0/n9 carray_p_0/n1 0.350042f
C40 dac_out carray_p_0/n2 6.640605f
C41 carray_p_0/n0 carray_p_0/n2 0.099314f
C42 carray_p_0/n6 carray_p_0/ndum 0.025424f
C43 dac_out carray_p_0/n1 3.367623f
C44 carray_p_0/n5 carray_p_0/n2 0.208112f
C45 carray_p_0/n0 carray_p_0/n1 8.476914f
C46 carray_p_0/n6 carray_p_0/n7 34.662605f
C47 vdd carray_p_0/n2 0.002151f
C48 carray_p_0/ndum carray_p_0/n4 0.025424f
C49 carray_p_0/n9 carray_p_0/ndum 0.127951f
C50 carray_p_0/n8 carray_p_0/n3 1.46111f
C51 carray_p_0/n1 carray_p_0/n5 0.142354f
C52 carray_p_0/n1 vdd 0.002151f
C53 carray_p_0/n7 carray_p_0/n4 1.70387f
C54 carray_p_0/n9 carray_p_0/n7 29.516087f
C55 dac_out carray_p_0/ndum 1.640173f
C56 dac_out bootstrapped_sw_p_0/vbsl 0.207261f
C57 carray_p_0/n5 carray_p_0/ndum 0.025424f
C58 carray_p_0/n3 carray_p_0/n2 23.177217f
C59 ctl2 ctl3 0.104537f
C60 dac_out carray_p_0/n7 0.210031p
C61 carray_p_0/n6 carray_p_0/n9 14.716789f
C62 carray_p_0/n6 carray_p_0/n4 0.614078f
C63 ctl7 ctl8 0.104537f
C64 carray_p_0/n0 carray_p_0/n7 0.06073f
C65 vdd carray_p_0/ndum 0.004405f
C66 sample vdd 0.00675f
C67 carray_p_0/n1 carray_p_0/n3 0.145048f
C68 carray_p_0/n5 carray_p_0/n7 3.36878f
C69 dac_out carray_p_0/n6 0.105055p
C70 carray_p_0/n9 carray_p_0/n4 3.740573f
C71 carray_p_0/n7 vdd 0.002151f
C72 carray_p_0/n0 carray_p_0/n6 0.025424f
C73 carray_p_0/n8 carray_p_0/n2 0.770227f
C74 carray_p_0/n6 carray_p_0/n5 28.925901f
C75 carray_p_0/n8 carray_p_0/n1 0.28587f
C76 dac_out carray_p_0/n9 0.846161p
C77 dac_out carray_p_0/n4 26.32268f
C78 carray_p_0/ndum carray_p_0/n3 0.025424f
C79 carray_p_0/n6 vdd 0.002151f
C80 carray_p_0/n0 carray_p_0/n4 0.040502f
C81 carray_p_0/n0 carray_p_0/n9 0.521489f
C82 carray_p_0/n5 carray_p_0/n4 27.828503f
C83 carray_p_0/n9 carray_p_0/n5 7.399346f
C84 carray_p_0/n7 carray_p_0/n3 0.891504f
C85 carray_p_0/n0 dac_out 1.750611f
C86 carray_p_0/n9 vdd 0.002151f
C87 vdd carray_p_0/n4 0.002151f
C88 carray_p_0/n8 carray_p_0/ndum 0.097254f
C89 carray_p_0/n1 carray_p_0/n2 16.941952f
C90 carray_p_0/n2 vss 30.783176f
C91 carray_p_0/n3 vss 34.265587f
C92 carray_p_0/n4 vss 39.983223f
C93 carray_p_0/n5 vss 48.00648f
C94 carray_p_0/n9 vss 14.963586f
C95 dac_out vss -0.684032p
C96 carray_p_0/n8 vss 40.580837f
C97 carray_p_0/n7 vss 56.915478f
C98 carray_p_0/n6 vss 53.64827f
C99 carray_p_0/n0 vss 17.632519f
C100 carray_p_0/n1 vss 17.795374f
C101 bootstrapped_sw_p_0/vs vss 0.053987f
C102 bootstrapped_sw_p_0/enb vss 1.502816f
C103 dac_in vss 0.376878f
C104 bootstrapped_sw_p_0/vg vss 1.498165f
C105 bootstrapped_sw_p_0/vbsh vss 14.27723f
C106 bootstrapped_sw_p_0/vbsl vss 7.956583f
C107 sample vss 20.84873f
C108 ctl9 vss 0.916847f
C109 ctl8 vss 0.916847f
C110 ctl7 vss 0.916847f
C111 ctl6 vss 0.916847f
C112 ctl5 vss 0.916847f
C113 ctl4 vss 0.916847f
C114 ctl3 vss 0.916847f
C115 ctl1 vss 0.916847f
C116 vdd vss 19.888897f
C117 ctl10 vss 1.146163f
C118 ctl2 vss 0.916847f
C119 carray_p_0/ndum vss 14.881693f
C120 dum vss 1.125528f
.ends

.subckt inv_n VSS ZN I VDD VPW VNW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VDD VNW 0.082022f
C1 ZN VSS 0.180794f
C2 I ZN 0.58604f
C3 VDD ZN 0.271625f
C4 I VSS 0.091531f
C5 VDD VSS 0.029045f
C6 VDD I 0.074838f
C7 ZN VNW 0.023676f
C8 VNW VSS 0.006277f
C9 I VNW 0.285482f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu_n inv_n_8/I inv_n_1/I inv_n_7/ZN inv_n_4/ZN inv_n_1/ZN inv_n_3/I
+ vdd inv_n_5/I inv_n_7/I inv_n_9/ZN inv_n_9/I inv_n_6/ZN inv_n_10/ZN inv_n_3/ZN inv_n_0/ZN
+ inv_n_0/I inv_n_10/I inv_n_2/I inv_n_4/I inv_n_8/ZN inv_n_5/ZN inv_n_6/I inv_n_2/ZN
+ vss
Xinv_n_0 vss inv_n_0/ZN inv_n_0/I vdd inv_n_0/VPW vdd vss inv_n
Xinv_n_1 vss inv_n_1/ZN inv_n_1/I vdd inv_n_1/VPW vdd vss inv_n
Xinv_n_2 vss inv_n_2/ZN inv_n_2/I vdd inv_n_2/VPW vdd vss inv_n
Xinv_n_3 vss inv_n_3/ZN inv_n_3/I vdd inv_n_3/VPW vdd vss inv_n
Xinv_n_4 vss inv_n_4/ZN inv_n_4/I vdd inv_n_4/VPW vdd vss inv_n
Xinv_n_5 vss inv_n_5/ZN inv_n_5/I vdd inv_n_5/VPW vdd vss inv_n
Xinv_n_6 vss inv_n_6/ZN inv_n_6/I vdd inv_n_6/VPW vdd vss inv_n
Xinv_n_7 vss inv_n_7/ZN inv_n_7/I vdd inv_n_7/VPW vdd vss inv_n
Xinv_n_8 vss inv_n_8/ZN inv_n_8/I vdd inv_n_8/VPW vdd vss inv_n
Xinv_n_9 vss inv_n_9/ZN inv_n_9/I vdd inv_n_9/VPW vdd vss inv_n
Xinv_n_10 vss inv_n_10/ZN inv_n_10/I vdd inv_n_10/VPW vdd vss inv_n
C0 vss inv_n_9/ZN 0.003326f
C1 inv_n_5/I inv_n_6/ZN 0.028928f
C2 vss inv_n_2/ZN 0.005014f
C3 vdd inv_n_5/I 0.019437f
C4 vss inv_n_2/I 0.164788f
C5 vss inv_n_5/ZN 0.003326f
C6 inv_n_4/I vss 0.166388f
C7 inv_n_7/I inv_n_6/ZN 0.002086f
C8 vdd inv_n_7/I 0.019437f
C9 inv_n_9/ZN inv_n_9/I 0.029333f
C10 vss inv_n_0/I 0.170492f
C11 vss inv_n_10/ZN 0.003326f
C12 inv_n_1/ZN vss 0.003326f
C13 inv_n_1/I inv_n_3/ZN 0.002086f
C14 vdd inv_n_1/I 0.019437f
C15 inv_n_8/I inv_n_8/ZN 0.029333f
C16 vdd inv_n_3/ZN 0.159176f
C17 vdd inv_n_6/ZN 0.159176f
C18 inv_n_5/ZN inv_n_4/ZN 0.080571f
C19 inv_n_6/I inv_n_5/ZN 0.002086f
C20 vss inv_n_8/ZN 0.003326f
C21 inv_n_4/I inv_n_4/ZN 0.029333f
C22 inv_n_3/I inv_n_0/I 0.08416f
C23 inv_n_7/ZN inv_n_8/ZN 0.080571f
C24 vdd inv_n_10/I 0.019437f
C25 vss inv_n_5/I 0.166388f
C26 inv_n_1/ZN inv_n_3/I 0.028928f
C27 inv_n_0/I inv_n_0/ZN 0.029333f
C28 inv_n_1/ZN inv_n_4/ZN 0.080571f
C29 inv_n_9/I inv_n_10/ZN 0.028928f
C30 inv_n_9/I inv_n_8/ZN 0.002086f
C31 inv_n_7/I inv_n_8/I 0.084161f
C32 vss inv_n_7/I 0.166388f
C33 inv_n_5/I inv_n_4/ZN 0.002086f
C34 inv_n_6/I inv_n_5/I 0.084161f
C35 inv_n_2/ZN inv_n_2/I 0.029333f
C36 inv_n_7/ZN inv_n_7/I 0.029333f
C37 vss inv_n_1/I 0.166388f
C38 vss inv_n_3/ZN 0.003326f
C39 vdd inv_n_8/I 0.019437f
C40 vss inv_n_6/ZN 0.003326f
C41 inv_n_9/ZN inv_n_10/ZN 0.080571f
C42 vss vdd 0.009518f
C43 inv_n_2/ZN inv_n_10/ZN 0.080571f
C44 inv_n_7/ZN inv_n_6/ZN 0.080571f
C45 inv_n_6/I inv_n_7/I 0.084161f
C46 vss inv_n_10/I 0.166388f
C47 inv_n_7/ZN vdd 0.159176f
C48 inv_n_4/I inv_n_5/ZN 0.028928f
C49 inv_n_9/ZN inv_n_8/ZN 0.080571f
C50 inv_n_3/I inv_n_1/I 0.084161f
C51 inv_n_10/ZN inv_n_2/I 0.002086f
C52 inv_n_3/I inv_n_3/ZN 0.029333f
C53 inv_n_1/I inv_n_4/ZN 0.028928f
C54 vdd inv_n_3/I 0.019437f
C55 inv_n_6/I inv_n_6/ZN 0.029333f
C56 inv_n_0/ZN inv_n_3/ZN 0.080571f
C57 inv_n_4/I inv_n_1/ZN 0.002086f
C58 vdd inv_n_4/ZN 0.159176f
C59 inv_n_6/I vdd 0.019437f
C60 vdd inv_n_0/ZN 0.184001f
C61 vdd inv_n_9/I 0.019437f
C62 inv_n_10/I inv_n_9/I 0.084161f
C63 inv_n_5/I inv_n_5/ZN 0.029333f
C64 inv_n_4/I inv_n_5/I 0.084161f
C65 vss inv_n_8/I 0.166388f
C66 inv_n_7/ZN inv_n_8/I 0.002086f
C67 vss inv_n_7/ZN 0.003326f
C68 vdd inv_n_9/ZN 0.159176f
C69 inv_n_2/ZN vdd 0.174722f
C70 vss inv_n_3/I 0.166388f
C71 inv_n_10/I inv_n_9/ZN 0.002086f
C72 vss inv_n_4/ZN 0.003326f
C73 inv_n_9/I inv_n_8/I 0.084161f
C74 inv_n_2/ZN inv_n_10/I 0.028928f
C75 vss inv_n_6/I 0.166388f
C76 vss inv_n_0/ZN 0.005399f
C77 vss inv_n_9/I 0.166388f
C78 inv_n_4/I inv_n_1/I 0.084161f
C79 vdd inv_n_2/I 0.035575f
C80 inv_n_6/ZN inv_n_5/ZN 0.080571f
C81 inv_n_7/ZN inv_n_6/I 0.028928f
C82 vdd inv_n_5/ZN 0.159176f
C83 inv_n_4/I vdd 0.019437f
C84 inv_n_10/I inv_n_2/I 0.084161f
C85 inv_n_0/I inv_n_3/ZN 0.028928f
C86 inv_n_7/I inv_n_8/ZN 0.028928f
C87 inv_n_1/ZN inv_n_1/I 0.029333f
C88 vdd inv_n_0/I 0.026972f
C89 inv_n_1/ZN inv_n_3/ZN 0.080571f
C90 vdd inv_n_10/ZN 0.159176f
C91 inv_n_1/ZN vdd 0.159176f
C92 inv_n_3/I inv_n_0/ZN 0.002086f
C93 inv_n_10/I inv_n_10/ZN 0.029333f
C94 vdd inv_n_8/ZN 0.159176f
C95 inv_n_9/ZN inv_n_8/I 0.028928f
C96 inv_n_10/ZN 0 0.131999f
C97 inv_n_10/I 0 0.64919f
C98 inv_n_9/ZN 0 0.131999f
C99 inv_n_9/I 0 0.64919f
C100 inv_n_8/ZN 0 0.131999f
C101 inv_n_8/I 0 0.64919f
C102 inv_n_7/ZN 0 0.131999f
C103 inv_n_7/I 0 0.64919f
C104 inv_n_6/ZN 0 0.131999f
C105 inv_n_6/I 0 0.64919f
C106 inv_n_5/ZN 0 0.131999f
C107 inv_n_5/I 0 0.64919f
C108 inv_n_4/ZN 0 0.131999f
C109 inv_n_4/I 0 0.64919f
C110 inv_n_3/ZN 0 0.131999f
C111 inv_n_3/I 0 0.64919f
C112 vss 0 3.02573f
C113 inv_n_2/ZN 0 0.206166f
C114 vdd 0 16.013325f
C115 inv_n_2/I 0 0.750024f
C116 inv_n_1/ZN 0 0.131999f
C117 inv_n_1/I 0 0.64919f
C118 inv_n_0/ZN 0 0.209411f
C119 inv_n_0/I 0 0.731246f
.ends

.subckt XM2_bs_n G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S G 0.002868f
C1 S D 0.038197f
C2 D G 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XMs1_bs_n G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 D G 0.002868f
C2 G S 0.002868f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365275f
.ends

.subckt XM3_bs_n G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 S G 0.002389f
C1 D w_n319_n356# 0.019807f
C2 S w_n319_n356# 0.021189f
C3 S D 0.045397f
C4 w_n319_n356# G 0.186402f
C5 D G 0.002389f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMs2_bs_n G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S G 0.002868f
C1 S D 0.038197f
C2 D G 0.002868f
C3 D a_n302_n324# 0.068446f
C4 S a_n302_n324# 0.068446f
C5 G a_n302_n324# 0.365186f
.ends

.subckt XM4_bs_n G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 S G 0.002389f
C1 D w_n319_n356# 0.019807f
C2 S w_n319_n356# 0.021189f
C3 S D 0.045397f
C4 w_n319_n356# G 0.186402f
C5 D G 0.002389f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XM1_bs_inv_n G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 D G 0.002868f
C2 G S 0.002868f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.066063f
C5 G a_n302_n324# 0.365365f
.ends

.subckt XM2_bs_inv_n G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 S G 0.002389f
C1 D w_n319_n356# 0.019807f
C2 S w_n319_n356# 0.019807f
C3 S D 0.045397f
C4 w_n319_n356# G 0.186609f
C5 D G 0.002389f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.48751f
.ends

.subckt bs_inv_n inv_out vdd inv_in vss
XXM1_bs_inv_n_0 inv_in inv_out vss vss XM1_bs_inv_n
XXM2_bs_inv_n_0 inv_in inv_out vdd vdd vss XM2_bs_inv_n
C0 inv_out vss 0.04895f
C1 vdd inv_in 0.07083f
C2 inv_out vdd 0.092565f
C3 inv_out inv_in 0.075645f
C4 vdd vss 0.043239f
C5 inv_in vss 0.037258f
C6 vdd 0 1.650725f
C7 inv_out 0 0.392313f
C8 vss 0 0.277512f
C9 inv_in 0 0.605506f
.ends

.subckt bs_cap_n I1_1_1_R0_BOT I1_1_1_R0_TOP VSUBS
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.339999u c_length=12.339999u
C0 I1_1_1_R0_BOT I1_1_1_R0_TOP 0.730455f
C1 I1_1_1_R0_TOP VSUBS 2.59113f
C2 I1_1_1_R0_BOT VSUBS 1.76085f
.ends

.subckt XMs_bs_n G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D G 0.002868f
C1 G S 0.002868f
C2 D S 0.038197f
C3 D a_n302_n324# 0.061336f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361785f
.ends

.subckt XM1_bs_n G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S D 0.038197f
C1 G D 0.002868f
C2 S G 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt bootstrapped_sw_n enb bs_in bs_out vg vs vdd en vbsl vss vbsh
XXM2_bs_n_0 enb vbsl vss vss vss XM2_bs_n
XXMs1_bs_n_0 vdd vs vss vg XMs1_bs_n
XXM3_bs_n_0 enb vg vbsh vbsh vss XM3_bs_n
XXMs2_bs_n_0 enb vss vss vss vs XMs2_bs_n
XXM4_bs_n_0 vg vdd vbsh vbsh vss XM4_bs_n
Xbs_inv_n_0 enb vdd en vss bs_inv_n
Xbs_cap_n_0 vbsl vbsh vss bs_cap_n
Xbs_cap_n_1 vbsl vbsh vss bs_cap_n
Xbs_cap_n_2 vbsl vbsh vss bs_cap_n
Xbs_cap_n_4 vbsl vbsh vss bs_cap_n
Xbs_cap_n_3 vbsl vbsh vss bs_cap_n
XXMs_bs_n_0 vg bs_out vss bs_in XMs_bs_n
XXM1_bs_n_0 vg vbsl vss vss bs_in XM1_bs_n
C0 vbsl vdd 0.002507f
C1 vbsh enb 0.0922f
C2 vg vdd 0.500479f
C3 vdd en 0.086628f
C4 enb vdd 0.426791f
C5 vbsh vdd 0.205818f
C6 vbsl bs_out 0.057454f
C7 vg bs_out 0.066304f
C8 vbsl bs_in 0.256003f
C9 vs vg 0.007099f
C10 bs_in vg 0.079028f
C11 bs_out enb 0.001285f
C12 vbsh bs_out 0.119559f
C13 vs enb 0.00173f
C14 vbsh bs_in 0.013047f
C15 bs_out vdd 0.008497f
C16 vbsl vg 0.043332f
C17 vg en 0.002156f
C18 vbsl enb 0.01529f
C19 vbsh vbsl 0.870275f
C20 vg enb 0.583075f
C21 vbsh vg 0.283904f
C22 enb en 0.018916f
C23 bs_out vss 0.895635f
C24 bs_in vss 0.389944f
C25 vg vss 1.576155f
C26 vbsh vss 14.292329f
C27 vbsl vss 8.158694f
C28 vdd vss 3.558326f
C29 en vss 0.896531f
C30 vs vss 0.042967f
C31 enb vss 1.703464f
.ends

.subckt dacn dac_in ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10 bootstrapped_sw_n_0/vg
+ bootstrapped_sw_n_0/enb carray_n_0/n9 sample carray_n_0/n7 carray_n_0/n0 vdd carray_n_0/n8
+ bootstrapped_sw_n_0/vbsh dac_out dum vss bootstrapped_sw_n_0/vbsl carray_n_0/ndum
Xinv_renketu_n_0 ctl7 ctl2 carray_n_0/n6 carray_n_0/n3 carray_n_0/n2 ctl1 vdd ctl4
+ ctl6 carray_n_0/n8 ctl8 carray_n_0/n5 carray_n_0/n9 carray_n_0/n1 carray_n_0/ndum
+ dum ctl9 ctl10 ctl3 carray_n_0/n7 carray_n_0/n4 ctl5 carray_n_0/n0 vss inv_renketu_n
Xbootstrapped_sw_n_0 bootstrapped_sw_n_0/enb dac_in dac_out bootstrapped_sw_n_0/vg
+ bootstrapped_sw_n_0/vs vdd sample bootstrapped_sw_n_0/vbsl vss bootstrapped_sw_n_0/vbsh
+ bootstrapped_sw_n
C0 sample carray_n_0/ndum 0.045492f
C1 carray_n_0/n2 carray_n_0/n0 0.099314f
C2 carray_n_0/n0 carray_n_0/n8 0.097254f
C3 carray_n_0/ndum carray_n_0/n9 0.127951f
C4 carray_n_0/n4 carray_n_0/n6 0.614078f
C5 carray_n_0/n7 dac_out 0.210031p
C6 carray_n_0/n3 carray_n_0/n2 23.177217f
C7 carray_n_0/n3 carray_n_0/n8 1.46111f
C8 carray_n_0/n5 dac_out 52.565514f
C9 carray_n_0/n2 carray_n_0/n8 0.770227f
C10 carray_n_0/ndum carray_n_0/n6 0.025424f
C11 carray_n_0/n1 carray_n_0/n7 0.212822f
C12 carray_n_0/n6 carray_n_0/n9 14.716789f
C13 carray_n_0/n5 carray_n_0/n1 0.142354f
C14 carray_n_0/n0 dac_out 1.750611f
C15 carray_n_0/n4 carray_n_0/n7 1.70387f
C16 vdd carray_n_0/n1 0.002151f
C17 bootstrapped_sw_n_0/vbsl dac_out 0.207261f
C18 carray_n_0/n5 carray_n_0/n4 27.828503f
C19 ctl5 ctl4 0.104537f
C20 ctl3 ctl4 0.104537f
C21 vdd carray_n_0/n4 0.002151f
C22 carray_n_0/n3 dac_out 13.201303f
C23 carray_n_0/n1 carray_n_0/n0 8.476914f
C24 carray_n_0/n2 dac_out 6.640605f
C25 carray_n_0/n8 dac_out 0.420151p
C26 ctl5 ctl6 0.104537f
C27 ctl9 ctl8 0.104537f
C28 carray_n_0/n4 carray_n_0/n0 0.040502f
C29 carray_n_0/ndum carray_n_0/n7 0.06073f
C30 carray_n_0/n3 carray_n_0/n1 0.145048f
C31 carray_n_0/n5 carray_n_0/ndum 0.025424f
C32 carray_n_0/n7 carray_n_0/n9 29.516087f
C33 vdd carray_n_0/ndum 0.004405f
C34 sample vdd 0.00675f
C35 carray_n_0/n5 carray_n_0/n9 7.399346f
C36 carray_n_0/n3 carray_n_0/n4 26.229403f
C37 carray_n_0/n2 carray_n_0/n1 16.941952f
C38 carray_n_0/n1 carray_n_0/n8 0.28587f
C39 bootstrapped_sw_n_0/vbsh dac_out 0.280658f
C40 vdd carray_n_0/n9 0.002151f
C41 ctl8 ctl7 0.104537f
C42 carray_n_0/n2 carray_n_0/n4 0.213209f
C43 ctl2 ctl1 0.104537f
C44 carray_n_0/n4 carray_n_0/n8 2.84323f
C45 carray_n_0/n0 carray_n_0/n9 0.521489f
C46 carray_n_0/n6 carray_n_0/n7 34.662605f
C47 carray_n_0/n3 carray_n_0/ndum 0.025424f
C48 carray_n_0/n5 carray_n_0/n6 28.925901f
C49 vdd carray_n_0/n6 0.002151f
C50 carray_n_0/n3 carray_n_0/n9 1.911224f
C51 carray_n_0/n2 carray_n_0/ndum 0.041162f
C52 carray_n_0/ndum carray_n_0/n8 0.097254f
C53 carray_n_0/n1 dac_out 3.367623f
C54 carray_n_0/n2 carray_n_0/n9 0.996681f
C55 carray_n_0/n8 carray_n_0/n9 87.43918f
C56 carray_n_0/n4 dac_out 26.32268f
C57 carray_n_0/n0 carray_n_0/n6 0.025424f
C58 carray_n_0/n3 carray_n_0/n6 0.336612f
C59 carray_n_0/n5 carray_n_0/n7 3.36878f
C60 carray_n_0/n4 carray_n_0/n1 0.142475f
C61 vdd carray_n_0/n7 0.002151f
C62 carray_n_0/n2 carray_n_0/n6 0.20799f
C63 carray_n_0/n6 carray_n_0/n8 11.2161f
C64 carray_n_0/n5 vdd 0.002151f
C65 carray_n_0/ndum dac_out 1.640173f
C66 ctl3 ctl2 0.104537f
C67 dac_out carray_n_0/n9 0.846161p
C68 carray_n_0/n0 carray_n_0/n7 0.06073f
C69 carray_n_0/n5 carray_n_0/n0 0.025424f
C70 carray_n_0/ndum carray_n_0/n1 8.498201f
C71 ctl10 ctl9 0.104537f
C72 vdd carray_n_0/n0 0.002151f
C73 carray_n_0/n3 carray_n_0/n7 0.891504f
C74 carray_n_0/n1 carray_n_0/n9 0.350042f
C75 ctl6 ctl7 0.104537f
C76 carray_n_0/n4 carray_n_0/ndum 0.025424f
C77 carray_n_0/n3 carray_n_0/n5 0.346757f
C78 carray_n_0/n2 carray_n_0/n7 0.485355f
C79 carray_n_0/n4 carray_n_0/n9 3.740573f
C80 carray_n_0/n3 vdd 0.002151f
C81 carray_n_0/n7 carray_n_0/n8 50.51461f
C82 carray_n_0/n6 dac_out 0.105055p
C83 carray_n_0/n5 carray_n_0/n2 0.208112f
C84 carray_n_0/n5 carray_n_0/n8 5.60732f
C85 vdd carray_n_0/n2 0.002151f
C86 vdd carray_n_0/n8 0.002151f
C87 carray_n_0/n3 carray_n_0/n0 0.051666f
C88 dum ctl1 0.104537f
C89 carray_n_0/n1 carray_n_0/n6 0.142211f
C90 carray_n_0/n9 vss 14.963586f
C91 dac_out vss -0.684032p
C92 carray_n_0/n8 vss 40.580837f
C93 carray_n_0/n7 vss 56.915478f
C94 carray_n_0/n6 vss 53.64827f
C95 carray_n_0/n0 vss 17.632519f
C96 carray_n_0/n1 vss 17.795374f
C97 carray_n_0/n2 vss 30.783176f
C98 carray_n_0/n3 vss 34.265587f
C99 carray_n_0/n4 vss 39.983223f
C100 carray_n_0/n5 vss 48.00648f
C101 dac_in vss 0.376878f
C102 bootstrapped_sw_n_0/vg vss 1.498165f
C103 bootstrapped_sw_n_0/vbsh vss 14.27723f
C104 bootstrapped_sw_n_0/vbsl vss 7.956583f
C105 sample vss 20.84873f
C106 bootstrapped_sw_n_0/vs vss 0.053987f
C107 bootstrapped_sw_n_0/enb vss 1.502816f
C108 ctl9 vss 0.916847f
C109 ctl8 vss 0.916847f
C110 ctl7 vss 0.916847f
C111 ctl6 vss 0.916847f
C112 ctl5 vss 0.916847f
C113 ctl4 vss 0.916847f
C114 ctl3 vss 0.916847f
C115 ctl1 vss 0.916847f
C116 vdd vss 19.888895f
C117 ctl10 vss 1.146163f
C118 ctl2 vss 0.916847f
C119 carray_n_0/ndum vss 14.881693f
C120 dum vss 1.125528f
.ends

.subckt XMdiff_cmp a_192_n100# a_n280_n100# a_n192_n183# a_n52_n100# a_n424_n324#
+ a_52_n183#
X0 a_192_n100# a_52_n183# a_n52_n100# a_n424_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n52_n100# a_n192_n183# a_n280_n100# a_n424_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
C0 a_52_n183# a_n52_n100# 0.002868f
C1 a_192_n100# a_n52_n100# 0.038197f
C2 a_52_n183# a_192_n100# 0.002868f
C3 a_n192_n183# a_n280_n100# 0.002868f
C4 a_n280_n100# a_n52_n100# 0.038197f
C5 a_n192_n183# a_n52_n100# 0.002868f
C6 a_n192_n183# a_52_n183# 0.039785f
C7 a_192_n100# a_n424_n324# 0.113177f
C8 a_n52_n100# a_n424_n324# 0.036353f
C9 a_n280_n100# a_n424_n324# 0.113177f
C10 a_52_n183# a_n424_n324# 0.342168f
C11 a_n192_n183# a_n424_n324# 0.342168f
.ends

.subckt XM3_trims_right a_n2052_n100# a_n2668_n324# a_n1808_n100# a_n1948_n183# a_n1564_n100#
+ a_n2524_n100# a_n1704_n183# a_n2296_n100# a_n2192_n183# a_n2436_n183#
X0 a_n2052_n100# a_n2192_n183# a_n2296_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n1564_n100# a_n1704_n183# a_n1808_n100# a_n2668_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X2 a_n1808_n100# a_n1948_n183# a_n2052_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_n2296_n100# a_n2436_n183# a_n2524_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
C0 a_n2296_n100# a_n2192_n183# 0.002868f
C1 a_n1948_n183# a_n1808_n100# 0.002868f
C2 a_n2052_n100# a_n1808_n100# 0.038197f
C3 a_n2296_n100# a_n2052_n100# 0.038197f
C4 a_n2296_n100# a_n2524_n100# 0.038197f
C5 a_n1564_n100# a_n1808_n100# 0.038197f
C6 a_n1704_n183# a_n1948_n183# 0.039785f
C7 a_n2436_n183# a_n2192_n183# 0.039785f
C8 a_n1704_n183# a_n1564_n100# 0.002868f
C9 a_n2436_n183# a_n2524_n100# 0.002868f
C10 a_n1704_n183# a_n1808_n100# 0.002868f
C11 a_n1948_n183# a_n2192_n183# 0.039785f
C12 a_n2052_n100# a_n2192_n183# 0.002868f
C13 a_n2296_n100# a_n2436_n183# 0.002868f
C14 a_n2052_n100# a_n1948_n183# 0.002868f
C15 a_n1564_n100# a_n2668_n324# 0.061257f
C16 a_n1808_n100# a_n2668_n324# 0.036353f
C17 a_n2052_n100# a_n2668_n324# 0.036353f
C18 a_n2296_n100# a_n2668_n324# 0.036353f
C19 a_n2524_n100# a_n2668_n324# 0.113177f
C20 a_n1704_n183# a_n2668_n324# 0.334286f
C21 a_n1948_n183# a_n2668_n324# 0.306841f
C22 a_n2192_n183# a_n2668_n324# 0.30709f
C23 a_n2436_n183# a_n2668_n324# 0.34169f
.ends

.subckt XM0_trims_right G D a_n5334_252# a_n5334_n324# S
X0 S G D a_n5334_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 S G 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 S a_n5334_n324# 0.061257f
C4 D a_n5334_n324# 0.061257f
C5 G a_n5334_n324# 0.361695f
.ends

.subckt XM2_trims_right a_n4456_n324# a_n3948_n183# a_n3808_n100# a_n4280_n100# a_n4052_n100#
+ a_n4192_n183# a_n4456_252#
X0 a_n4052_n100# a_n4192_n183# a_n4280_n100# a_n4456_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X1 a_n3808_n100# a_n3948_n183# a_n4052_n100# a_n4456_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_n4280_n100# a_n4192_n183# 0.002868f
C1 a_n3808_n100# a_n3948_n183# 0.002868f
C2 a_n4052_n100# a_n3948_n183# 0.002868f
C3 a_n4052_n100# a_n4192_n183# 0.002868f
C4 a_n4052_n100# a_n4280_n100# 0.038197f
C5 a_n4052_n100# a_n3808_n100# 0.038197f
C6 a_n3948_n183# a_n4192_n183# 0.039785f
C7 a_n3808_n100# a_n4456_n324# 0.061257f
C8 a_n4052_n100# a_n4456_n324# 0.036353f
C9 a_n4280_n100# a_n4456_n324# 0.061257f
C10 a_n3948_n183# a_n4456_n324# 0.334154f
C11 a_n4192_n183# a_n4456_n324# 0.334154f
.ends

.subckt XM4_trims_right a_436_n100# a_192_n100# a_n1188_n324# a_n296_n100# a_784_n183#
+ a_n192_n183# a_n436_n183# a_540_n183# a_n52_n100# a_924_n100# a_680_n100# a_n1012_n100#
+ a_n784_n100# a_n924_n183# a_n680_n183# a_n540_n100# a_296_n183# a_52_n183#
X0 a_436_n100# a_296_n183# a_192_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n784_n100# a_n924_n183# a_n1012_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X2 a_192_n100# a_52_n183# a_n52_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_680_n100# a_540_n183# a_436_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X4 a_924_n100# a_784_n183# a_680_n100# a_n1188_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X5 a_n52_n100# a_n192_n183# a_n296_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X6 a_n296_n100# a_n436_n183# a_n540_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X7 a_n540_n100# a_n680_n183# a_n784_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_n436_n183# a_n296_n100# 0.002868f
C1 a_52_n183# a_n52_n100# 0.002868f
C2 a_680_n100# a_540_n183# 0.002868f
C3 a_924_n100# a_784_n183# 0.002868f
C4 a_n192_n183# a_n296_n100# 0.002868f
C5 a_436_n100# a_680_n100# 0.038197f
C6 a_436_n100# a_540_n183# 0.002868f
C7 a_n784_n100# a_n680_n183# 0.002868f
C8 a_n436_n183# a_n540_n100# 0.002868f
C9 a_680_n100# a_784_n183# 0.002868f
C10 a_540_n183# a_784_n183# 0.039785f
C11 a_n540_n100# a_n680_n183# 0.002868f
C12 a_296_n183# a_540_n183# 0.039785f
C13 a_n784_n100# a_n1012_n100# 0.038197f
C14 a_436_n100# a_192_n100# 0.038197f
C15 a_436_n100# a_296_n183# 0.002868f
C16 a_52_n183# a_n192_n183# 0.039785f
C17 a_n540_n100# a_n296_n100# 0.038197f
C18 a_n924_n183# a_n680_n183# 0.039785f
C19 a_n784_n100# a_n540_n100# 0.038197f
C20 a_296_n183# a_192_n100# 0.002868f
C21 a_n192_n183# a_n52_n100# 0.002868f
C22 a_n924_n183# a_n1012_n100# 0.002868f
C23 a_n296_n100# a_n52_n100# 0.038197f
C24 a_n924_n183# a_n784_n100# 0.002868f
C25 a_52_n183# a_192_n100# 0.002868f
C26 a_52_n183# a_296_n183# 0.039785f
C27 a_n436_n183# a_n680_n183# 0.039785f
C28 a_n436_n183# a_n192_n183# 0.039785f
C29 a_924_n100# a_680_n100# 0.038197f
C30 a_192_n100# a_n52_n100# 0.038197f
C31 a_924_n100# a_n1188_n324# 0.113177f
C32 a_680_n100# a_n1188_n324# 0.036353f
C33 a_436_n100# a_n1188_n324# 0.036353f
C34 a_192_n100# a_n1188_n324# 0.036353f
C35 a_n52_n100# a_n1188_n324# 0.036353f
C36 a_n296_n100# a_n1188_n324# 0.036353f
C37 a_n540_n100# a_n1188_n324# 0.036353f
C38 a_n784_n100# a_n1188_n324# 0.036353f
C39 a_n1012_n100# a_n1188_n324# 0.061257f
C40 a_784_n183# a_n1188_n324# 0.34169f
C41 a_540_n183# a_n1188_n324# 0.30709f
C42 a_296_n183# a_n1188_n324# 0.306841f
C43 a_52_n183# a_n1188_n324# 0.306744f
C44 a_n192_n183# a_n1188_n324# 0.306698f
C45 a_n436_n183# a_n1188_n324# 0.306672f
C46 a_n680_n183# a_n1188_n324# 0.306613f
C47 a_n924_n183# a_n1188_n324# 0.334154f
.ends

.subckt XM1_trims_right G D a_n5302_n324# S a_n5302_252#
X0 D G S a_n5302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 G S 0.002868f
C2 S D 0.038197f
C3 D a_n5302_n324# 0.061257f
C4 S a_n5302_n324# 0.061257f
C5 G a_n5302_n324# 0.361695f
.ends

.subckt trim_switch_right d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 VSUBS
XXM3_trims_right_0 n3 VSUBS VSUBS d_3 n3 n3 d_3 VSUBS d_3 d_3 XM3_trims_right
XXM0_trims_right_0 d_0 n0 VSUBS VSUBS VSUBS XM0_trims_right
XXM2_trims_right_0 VSUBS d_2 n2 n2 VSUBS d_2 VSUBS XM2_trims_right
XXM4_trims_right_0 n4 VSUBS VSUBS VSUBS d_4 d_4 d_4 d_4 n4 n4 VSUBS n4 VSUBS d_4 d_4
+ n4 d_4 d_4 XM4_trims_right
XXM1_trims_right_0 d_1 n1 VSUBS VSUBS VSUBS XM1_trims_right
C0 d_2 n2 0.052339f
C1 n0 n2 0.068796f
C2 n3 n2 0.068796f
C3 d_1 d_0 0.106626f
C4 n0 n1 0.025226f
C5 d_2 d_0 0.047211f
C6 d_0 n0 0.05352f
C7 d_3 d_2 0.03061f
C8 d_3 n3 0.171874f
C9 d_1 n1 0.05352f
C10 n4 n1 0.068796f
C11 d_1 d_4 0.02706f
C12 d_4 n4 0.398929f
C13 n1 VSUBS 0.224565f
C14 d_1 VSUBS 0.520942f
C15 n4 VSUBS 2.074915f
C16 d_4 VSUBS 3.301902f
C17 n2 VSUBS 0.637701f
C18 d_2 VSUBS 0.94246f
C19 n0 VSUBS 0.224565f
C20 d_0 VSUBS 0.500402f
C21 n3 VSUBS 1.232816f
C22 d_3 VSUBS 1.769471f
.ends

.subckt trim_right d_0 d_4 d_1 d_2 d_3 drain n1 n4 n0 n2 n3 vss
Xtrim_switch_right_0 d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 vss trim_switch_right
C0 n3 n4 1.599582f
C1 drain n1 1.60623f
C2 d_0 n0 0.010314f
C3 drain n2 3.213024f
C4 drain n0 1.60623f
C5 d_4 n4 0.001311f
C6 n1 n2 0.092902f
C7 drain n3 6.427484f
C8 n1 n0 0.506269f
C9 n2 n0 0.116341f
C10 drain n4 12.877382f
C11 n1 n3 0.087807f
C12 n3 n2 0.584482f
C13 n1 d_1 0.009441f
C14 n1 n4 0.166777f
C15 n2 d_1 0.00105f
C16 n3 n0 0.087807f
C17 n2 n4 0.616308f
C18 n0 n4 0.166348f
C19 d_1 vss 0.446833f
C20 d_4 vss 2.753276f
C21 d_2 vss 0.774671f
C22 d_0 vss 0.431586f
C23 d_3 vss 1.473178f
C24 n0 vss 0.644951f
C25 n1 vss 0.660965f
C26 n4 vss 4.842311f
C27 drain vss -5.906306f
C28 n3 vss 3.481832f
C29 n2 vss 2.023079f
.ends

.subckt XMinp_cmp G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 G S 0.002868f
C2 G D 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM4_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.019807f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMl4_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.021497f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12132f
.ends

.subckt XMl3_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.021497f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XM3_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.021497f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XMinn_cmp G D a_n302_n324# a_n302_252# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 D S 0.038197f
C1 G S 0.002868f
C2 G D 0.002868f
C3 D a_n302_n324# 0.061257f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.361695f
.ends

.subckt XM2_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.19321f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.021497f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.043431f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.11767f
C9 w_n319_n356# VSUBS 2.12131f
.ends

.subckt XMl2_cmp G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 G D 0.002868f
C2 S D 0.038197f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.368221f
.ends

.subckt XM1_cmp G D w_n319_n356# S VSUBS
X0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
C0 w_n319_n356# G 0.186402f
C1 D S 0.045397f
C2 w_n319_n356# S 0.021189f
C3 w_n319_n356# D 0.019807f
C4 G S 0.002389f
C5 G D 0.002389f
C6 D VSUBS 0.0454f
C7 S VSUBS 0.0454f
C8 G VSUBS 0.124686f
C9 w_n319_n356# VSUBS 1.47408f
.ends

.subckt XMl1_cmp G D a_n302_n324# S
X0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 G D 0.002868f
C2 S D 0.038197f
C3 D a_n302_n324# 0.066063f
C4 S a_n302_n324# 0.061257f
C5 G a_n302_n324# 0.368221f
.ends

.subckt XM4_trims_left a_436_n100# a_192_n100# a_n1188_n324# a_n296_n100# a_784_n183#
+ a_n192_n183# a_n436_n183# a_540_n183# a_n52_n100# a_924_n100# a_680_n100# a_n1012_n100#
+ a_n784_n100# a_n924_n183# a_n680_n183# a_n540_n100# a_296_n183# a_52_n183#
X0 a_436_n100# a_296_n183# a_192_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n784_n100# a_n924_n183# a_n1012_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X2 a_192_n100# a_52_n183# a_n52_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_680_n100# a_540_n183# a_436_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X4 a_924_n100# a_784_n183# a_680_n100# a_n1188_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X5 a_n52_n100# a_n192_n183# a_n296_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X6 a_n296_n100# a_n436_n183# a_n540_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X7 a_n540_n100# a_n680_n183# a_n784_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_n52_n100# a_192_n100# 0.038197f
C1 a_n52_n100# a_n296_n100# 0.038197f
C2 a_784_n183# a_540_n183# 0.039785f
C3 a_680_n100# a_540_n183# 0.002868f
C4 a_52_n183# a_n192_n183# 0.039785f
C5 a_n924_n183# a_n680_n183# 0.039785f
C6 a_436_n100# a_540_n183# 0.002868f
C7 a_n784_n100# a_n540_n100# 0.038197f
C8 a_n784_n100# a_n1012_n100# 0.038197f
C9 a_n924_n183# a_n784_n100# 0.002868f
C10 a_52_n183# a_192_n100# 0.002868f
C11 a_n52_n100# a_52_n183# 0.002868f
C12 a_n192_n183# a_n436_n183# 0.039785f
C13 a_n540_n100# a_n436_n183# 0.002868f
C14 a_296_n183# a_436_n100# 0.002868f
C15 a_296_n183# a_192_n100# 0.002868f
C16 a_n784_n100# a_n680_n183# 0.002868f
C17 a_n296_n100# a_n436_n183# 0.002868f
C18 a_680_n100# a_784_n183# 0.002868f
C19 a_924_n100# a_784_n183# 0.002868f
C20 a_296_n183# a_540_n183# 0.039785f
C21 a_n52_n100# a_n192_n183# 0.002868f
C22 a_n296_n100# a_n192_n183# 0.002868f
C23 a_n296_n100# a_n540_n100# 0.038197f
C24 a_n924_n183# a_n1012_n100# 0.002868f
C25 a_924_n100# a_680_n100# 0.038197f
C26 a_436_n100# a_680_n100# 0.038197f
C27 a_n680_n183# a_n436_n183# 0.039785f
C28 a_296_n183# a_52_n183# 0.039785f
C29 a_436_n100# a_192_n100# 0.038197f
C30 a_n680_n183# a_n540_n100# 0.002868f
C31 a_924_n100# a_n1188_n324# 0.113177f
C32 a_680_n100# a_n1188_n324# 0.036353f
C33 a_436_n100# a_n1188_n324# 0.036353f
C34 a_192_n100# a_n1188_n324# 0.036353f
C35 a_n52_n100# a_n1188_n324# 0.036353f
C36 a_n296_n100# a_n1188_n324# 0.036353f
C37 a_n540_n100# a_n1188_n324# 0.036353f
C38 a_n784_n100# a_n1188_n324# 0.036353f
C39 a_n1012_n100# a_n1188_n324# 0.061257f
C40 a_784_n183# a_n1188_n324# 0.34169f
C41 a_540_n183# a_n1188_n324# 0.30709f
C42 a_296_n183# a_n1188_n324# 0.306841f
C43 a_52_n183# a_n1188_n324# 0.306744f
C44 a_n192_n183# a_n1188_n324# 0.306698f
C45 a_n436_n183# a_n1188_n324# 0.306672f
C46 a_n680_n183# a_n1188_n324# 0.306613f
C47 a_n924_n183# a_n1188_n324# 0.334154f
.ends

.subckt XM0_trims_left G D a_n5334_252# a_n5334_n324# S
X0 S G D a_n5334_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G D 0.002868f
C1 S G 0.002868f
C2 S D 0.038197f
C3 S a_n5334_n324# 0.061257f
C4 D a_n5334_n324# 0.061257f
C5 G a_n5334_n324# 0.361695f
.ends

.subckt XM1_trims_left G D a_n5302_n324# S a_n5302_252#
X0 D G S a_n5302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
C0 G S 0.002868f
C1 D G 0.002868f
C2 D S 0.038197f
C3 D a_n5302_n324# 0.061257f
C4 S a_n5302_n324# 0.061257f
C5 G a_n5302_n324# 0.361695f
.ends

.subckt XM2_trims_left a_n4456_n324# a_n3948_n183# a_n3808_n100# a_n4280_n100# a_n4052_n100#
+ a_n4192_n183# a_n4456_252#
X0 a_n4052_n100# a_n4192_n183# a_n4280_n100# a_n4456_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
X1 a_n3808_n100# a_n3948_n183# a_n4052_n100# a_n4456_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
C0 a_n3948_n183# a_n3808_n100# 0.002868f
C1 a_n4052_n100# a_n3808_n100# 0.038197f
C2 a_n4192_n183# a_n3948_n183# 0.039785f
C3 a_n4052_n100# a_n4192_n183# 0.002868f
C4 a_n4052_n100# a_n3948_n183# 0.002868f
C5 a_n4280_n100# a_n4192_n183# 0.002868f
C6 a_n4052_n100# a_n4280_n100# 0.038197f
C7 a_n3808_n100# a_n4456_n324# 0.061257f
C8 a_n4052_n100# a_n4456_n324# 0.036353f
C9 a_n4280_n100# a_n4456_n324# 0.061257f
C10 a_n3948_n183# a_n4456_n324# 0.334154f
C11 a_n4192_n183# a_n4456_n324# 0.334154f
.ends

.subckt XM3_trims_left a_n2052_n100# a_n2668_n324# a_n1808_n100# a_n1948_n183# a_n1564_n100#
+ a_n2524_n100# a_n1704_n183# a_n2296_n100# a_n2192_n183# a_n2436_n183#
X0 a_n2052_n100# a_n2192_n183# a_n2296_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X1 a_n1564_n100# a_n1704_n183# a_n1808_n100# a_n2668_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
X2 a_n1808_n100# a_n1948_n183# a_n2052_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
X3 a_n2296_n100# a_n2436_n183# a_n2524_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
C0 a_n1704_n183# a_n1564_n100# 0.002868f
C1 a_n2052_n100# a_n2296_n100# 0.038197f
C2 a_n1808_n100# a_n2052_n100# 0.038197f
C3 a_n2192_n183# a_n2052_n100# 0.002868f
C4 a_n2192_n183# a_n2296_n100# 0.002868f
C5 a_n2052_n100# a_n1948_n183# 0.002868f
C6 a_n1808_n100# a_n1948_n183# 0.002868f
C7 a_n2524_n100# a_n2296_n100# 0.038197f
C8 a_n2192_n183# a_n1948_n183# 0.039785f
C9 a_n1808_n100# a_n1564_n100# 0.038197f
C10 a_n2436_n183# a_n2296_n100# 0.002868f
C11 a_n2436_n183# a_n2192_n183# 0.039785f
C12 a_n2524_n100# a_n2436_n183# 0.002868f
C13 a_n1808_n100# a_n1704_n183# 0.002868f
C14 a_n1704_n183# a_n1948_n183# 0.039785f
C15 a_n1564_n100# a_n2668_n324# 0.061257f
C16 a_n1808_n100# a_n2668_n324# 0.036353f
C17 a_n2052_n100# a_n2668_n324# 0.036353f
C18 a_n2296_n100# a_n2668_n324# 0.036353f
C19 a_n2524_n100# a_n2668_n324# 0.113177f
C20 a_n1704_n183# a_n2668_n324# 0.334286f
C21 a_n1948_n183# a_n2668_n324# 0.306841f
C22 a_n2192_n183# a_n2668_n324# 0.30709f
C23 a_n2436_n183# a_n2668_n324# 0.34169f
.ends

.subckt trim_switch_left d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 VSUBS
XXM4_trims_left_0 n4 VSUBS VSUBS VSUBS d_4 d_4 d_4 d_4 n4 n4 VSUBS n4 VSUBS d_4 d_4
+ n4 d_4 d_4 XM4_trims_left
XXM0_trims_left_0 d_0 n0 VSUBS VSUBS VSUBS XM0_trims_left
XXM1_trims_left_0 d_1 n1 VSUBS VSUBS VSUBS XM1_trims_left
XXM2_trims_left_0 VSUBS d_2 n2 n2 VSUBS d_2 VSUBS XM2_trims_left
XXM3_trims_left_0 n3 VSUBS VSUBS d_3 n3 n3 d_3 VSUBS d_3 d_3 XM3_trims_left
C0 d_0 d_1 0.106626f
C1 d_1 d_4 0.02706f
C2 n3 n2 0.068796f
C3 d_0 n0 0.05352f
C4 n2 d_2 0.052339f
C5 d_1 n1 0.05352f
C6 n0 n1 0.025226f
C7 n2 n0 0.068796f
C8 d_4 n4 0.398929f
C9 n3 d_3 0.171874f
C10 d_0 d_2 0.047211f
C11 d_3 d_2 0.03061f
C12 n4 n1 0.068796f
C13 n3 VSUBS 1.232816f
C14 d_3 VSUBS 1.769471f
C15 n2 VSUBS 0.637701f
C16 d_2 VSUBS 0.94246f
C17 n1 VSUBS 0.224565f
C18 d_1 VSUBS 0.520942f
C19 n0 VSUBS 0.224565f
C20 d_0 VSUBS 0.500402f
C21 n4 VSUBS 2.074915f
C22 d_4 VSUBS 3.301902f
.ends

.subckt trim_left d_0 d_4 d_1 d_2 d_3 drain n1 n0 n2 n3 n4 vss
Xtrim_switch_left_0 d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 vss trim_switch_left
C0 n2 n1 0.092902f
C1 n3 n1 0.087807f
C2 n4 drain 12.877382f
C3 d_1 n2 0.00105f
C4 n0 drain 1.60623f
C5 n0 n4 0.166348f
C6 n3 n2 0.584482f
C7 drain n1 1.60623f
C8 n4 n1 0.166777f
C9 n0 n1 0.506269f
C10 d_4 n4 0.001311f
C11 drain n2 3.213024f
C12 n4 n2 0.616308f
C13 n0 d_0 0.010314f
C14 drain n3 6.427484f
C15 n4 n3 1.599582f
C16 n0 n2 0.116341f
C17 d_1 n1 0.009441f
C18 n0 n3 0.087807f
C19 n0 vss 0.644951f
C20 n1 vss 0.660965f
C21 n4 vss 4.842311f
C22 drain vss -5.906306f
C23 n3 vss 3.481832f
C24 n2 vss 2.023079f
C25 d_3 vss 1.473178f
C26 d_2 vss 0.774671f
C27 d_1 vss 0.446833f
C28 d_0 vss 0.431586f
C29 d_4 vss 2.753276f
.ends

.subckt comparator trim1 trim0 trim4 trimb4 trimb1 trimb0 trimb2 trimb3 vp vn in ip
+ diff trim_right_0/n3 trim_left_0/n4 trim_left_0/n2 trim_left_0/n3 clkc trim3 outp
+ trim2 vdd outn trim_right_0/n4 trim_right_0/n2 vss
XXMdiff_cmp_0 vss vss clkc diff vss clkc XMdiff_cmp
Xtrim_right_0 trimb0 trimb4 trimb1 trimb2 trimb3 ip trim_right_0/n1 trim_right_0/n4
+ trim_right_0/n0 trim_right_0/n2 trim_right_0/n3 vss trim_right
XXMinp_cmp_0 vp ip vss vss diff XMinp_cmp
XXM4_cmp_0 clkc ip vdd vdd vss XM4_cmp
XXMl4_cmp_0 outn outp vdd vdd vss XMl4_cmp
XXMl3_cmp_0 outp outn vdd vdd vss XMl3_cmp
XXM3_cmp_0 clkc outp vdd vdd vss XM3_cmp
XXMinn_cmp_0 vn in vss vss diff XMinn_cmp
XXM2_cmp_0 clkc outn vdd vdd vss XM2_cmp
XXMl2_cmp_0 outn outp vss ip XMl2_cmp
XXM1_cmp_0 clkc in vdd vdd vss XM1_cmp
XXMl1_cmp_0 outp outn vss in XMl1_cmp
Xtrim_left_0 trim0 trim4 trim1 trim2 trim3 in trim_left_0/n1 trim_left_0/n0 trim_left_0/n2
+ trim_left_0/n3 trim_left_0/n4 vss trim_left
C0 diff outn 0.002551f
C1 vp ip 0.448228f
C2 trim_right_0/n0 ip 1.606869f
C3 trim_left_0/n1 trim_left_0/n4 0.032158f
C4 in outp 0.018491f
C5 vdd outp 0.454873f
C6 trim_right_0/n1 trim_right_0/n0 0.032158f
C7 clkc ip 0.528032f
C8 vp outp 0.256864f
C9 trim_left_0/n2 in 3.218424f
C10 trim0 trim2 0.786004f
C11 trim0 trim1 0.713549f
C12 trim_left_0/n3 in 6.426837f
C13 trimb2 trimb4 0.001666f
C14 outn ip 0.018487f
C15 clkc outp 0.295692f
C16 trim_left_0/n4 trim1 0.001799f
C17 outp vn 0.19705f
C18 vdd in 0.108547f
C19 trim_left_0/n2 trim_left_0/n4 0.128631f
C20 trim4 trim2 0.001666f
C21 diff ip 0.098316f
C22 trim_right_0/n3 trim_right_0/n4 0.241184f
C23 trim4 trim1 0.397758f
C24 trimb0 trimb1 0.713549f
C25 trim_right_0/n4 trim_right_0/n2 0.128631f
C26 trim_left_0/n3 trim_left_0/n4 0.241184f
C27 ip trim_right_0/n3 6.426837f
C28 in trim_left_0/n4 12.853152f
C29 trimb1 trim_right_0/n4 0.001799f
C30 ip trim_right_0/n2 3.218424f
C31 vp vdd 0.069074f
C32 outn outp 1.39519f
C33 diff outp 0.005373f
C34 clkc in 0.528032f
C35 trim0 trim4 0.002527f
C36 trim_left_0/n0 trim_left_0/n1 0.032158f
C37 in vn 0.448228f
C38 trimb2 trimb3 0.902342f
C39 ip trim_right_0/n4 12.853152f
C40 vdd clkc 0.289807f
C41 vdd vn 0.069074f
C42 vp clkc 0.133362f
C43 trim_left_0/n4 trim4 0.002904f
C44 vp vn 0.125877f
C45 outn in 0.103141f
C46 trim_right_0/n1 trim_right_0/n4 0.032158f
C47 vdd outn 0.503383f
C48 diff in 0.098316f
C49 trimb2 trimb0 0.786004f
C50 trim_right_0/n1 ip 1.606869f
C51 vp outn 0.159375f
C52 ip outp 0.10316f
C53 clkc vn 0.133362f
C54 vp diff 0.009142f
C55 trim3 trim2 0.902342f
C56 outn clkc 0.29566f
C57 trim_left_0/n0 in 1.606869f
C58 outn vn 0.199287f
C59 trimb0 trimb4 0.002527f
C60 trimb1 trimb4 0.397758f
C61 diff clkc 0.076203f
C62 trim_left_0/n1 in 1.606869f
C63 diff vn 0.009142f
C64 trimb4 trim_right_0/n4 0.002904f
C65 vdd ip 0.108547f
C66 trim_right_0/n0 trim_right_0/n4 0.032158f
C67 trim_left_0/n0 trim_left_0/n4 0.032158f
C68 trim_left_0/n0 vss 0.627477f
C69 trim_left_0/n1 vss 0.643951f
C70 trim_left_0/n4 vss 4.718663f
C71 in vss -4.355123f
C72 trim_left_0/n3 vss 3.342805f
C73 trim_left_0/n2 vss 1.998525f
C74 trim3 vss 3.460291f
C75 trim2 vss 1.618011f
C76 trim1 vss 1.092722f
C77 trim0 vss 1.058742f
C78 trim4 vss 3.293701f
C79 outp vss 2.729559f
C80 outn vss 2.683582f
C81 vdd vss 9.2164f
C82 vn vss 1.234778f
C83 vp vss 1.219948f
C84 trimb1 vss 1.092722f
C85 trimb4 vss 3.293701f
C86 trimb2 vss 1.618011f
C87 trimb0 vss 1.058742f
C88 trimb3 vss 3.460291f
C89 trim_right_0/n0 vss 0.627477f
C90 trim_right_0/n1 vss 0.643951f
C91 trim_right_0/n4 vss 4.718663f
C92 ip vss -4.354997f
C93 trim_right_0/n3 vss 3.342805f
C94 trim_right_0/n2 vss 1.998525f
C95 diff vss 0.291624f
C96 clkc vss 5.191715f
.ends

.subckt cap_mim_2p0fF_RCWXT2$1 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3120_n3000# m4_n3240_n3120# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30_flip cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$1
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_RCWXT2 m4_n3120_n3000# m4_n3240_n3120# VSUBS
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3120_n3000# m4_n3240_n3120# 2.57661f
C1 m4_n3120_n3000# VSUBS 9.60519f
C2 m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap1 vss vdd VSUBS
Xmim_cap_30_30_flip_233 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_222 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_200 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_211 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_68 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_57 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_79 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_13 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_24 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_46 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_35 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_213 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_224 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_202 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_235 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_212 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_234 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_223 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_201 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_58 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_69 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_14 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_25 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_47 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_36 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_214 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_225 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_203 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_236 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_224 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_213 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_235 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_202 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_59 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_15 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_48 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_26 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_37 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_226 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_204 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_237 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_215 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_225 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_214 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_236 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_203 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_16 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_49 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_38 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_27 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_227 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_238 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_205 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_216 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_226 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_215 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_237 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_204 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_17 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_28 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_39 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_228 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_217 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_239 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_206 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_227 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_216 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_238 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_205 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_18 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_29 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_229 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_218 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_207 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_228 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_217 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_206 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_239 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_19 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_219 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_208 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_229 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_218 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_207 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_209 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_219 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_208 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_190 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_209 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_90 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_180 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_191 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_80 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_91 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_190 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_170 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_181 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_192 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_81 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_70 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_92 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_0 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_191 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_180 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_0 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_160 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_193 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_182 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_171 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_60 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_82 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_71 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_93 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_1 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_170 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_192 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_181 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_1 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_183 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_172 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_150 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_194 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_161 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_83 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_72 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_94 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_50 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_61 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_2 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_160 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_193 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_182 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_171 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_2 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_173 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_162 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_184 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_195 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_140 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_151 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_73 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_84 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_95 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_51 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_40 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_62 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_3 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_161 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_172 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_194 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_183 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_150 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_3 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_174 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_152 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_141 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_196 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_130 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_185 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_163 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_30 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_74 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_85 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_52 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_96 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_41 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_63 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_4 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_151 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_162 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_140 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_173 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_184 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_195 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_4 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_131 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_120 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_153 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_186 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_142 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_197 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_164 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_175 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_31 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_75 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_20 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_64 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_86 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_42 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_53 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_97 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_5 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_152 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_163 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_141 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_174 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_130 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_196 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_185 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_5 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_154 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_176 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_165 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_110 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_132 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_121 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_143 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_198 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_187 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_76 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_21 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_65 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_10 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_32 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_43 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_54 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_87 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_98 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_6 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_153 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_164 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_175 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_131 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_142 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_120 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_197 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_186 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_6 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_155 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_166 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_111 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_100 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_133 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_144 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_122 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_199 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_188 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_177 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_77 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_22 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_66 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_11 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_99 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_33 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_44 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_55 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_88 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_7 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_110 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_121 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_154 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_176 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_143 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_198 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_187 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_132 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_165 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_7 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_156 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_167 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_178 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_101 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_112 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_145 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_123 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_189 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_134 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_23 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_67 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_78 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_12 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_34 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_56 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_45 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_89 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_8 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_100 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_111 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_177 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_188 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_133 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_122 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_199 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_144 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_155 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_166 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_8 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_168 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_157 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_179 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_102 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_113 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_135 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_146 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_124 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_68 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_79 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_24 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_13 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_35 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_57 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_46 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_9 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_156 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_145 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_101 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_112 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_123 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_178 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_134 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_189 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_167 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_9 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_103 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_114 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_136 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_147 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_125 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_169 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_158 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_14 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_69 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_25 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_58 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_36 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_47 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_157 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_168 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_146 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_113 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_102 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_135 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_124 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_179 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_104 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_115 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_137 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_148 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_126 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_159 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_15 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_26 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_59 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_37 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_48 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_158 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_147 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_169 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_114 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_103 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_136 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_125 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_105 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_116 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_149 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_138 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_127 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_16 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_27 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_38 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_49 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_115 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_104 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_137 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_126 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_148 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_159 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_117 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_106 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_139 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_128 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_17 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_28 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_39 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_149 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_116 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_105 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_138 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_127 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_118 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_107 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_129 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_90 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_29 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_18 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_117 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_106 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_139 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_128 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_119 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_108 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_80 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_91 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_19 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_118 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_107 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_129 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_109 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_70 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_81 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_92 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_119 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_108 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_82 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_60 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_71 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_93 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_109 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_50 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_83 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_72 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_61 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_94 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_73 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_84 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_62 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_95 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_51 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_40 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_74 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_52 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_85 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_63 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_96 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_30 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_41 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_230 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_75 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_20 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_64 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_86 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_53 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_31 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_42 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_97 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_220 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_231 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_230 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_65 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_76 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_10 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_54 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_21 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_87 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_32 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_43 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_98 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_221 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_232 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_210 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_231 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_220 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_66 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_77 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_11 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_22 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_88 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_44 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_99 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_33 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_55 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_222 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_233 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_200 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_211 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_flip_232 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_221 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_flip_210 vss vdd VSUBS mim_cap_30_30_flip
Xmim_cap_30_30_67 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_12 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_23 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_56 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_78 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_89 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_45 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_34 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_212 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_234 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_223 vss vdd VSUBS mim_cap_30_30
Xmim_cap_30_30_201 vss vdd VSUBS mim_cap_30_30
C0 vss vdd 0.196596p
C1 vdd VSUBS 4.633771p
C2 vss VSUBS 2.2518p
.ends

.subckt cap_mim_2p0fF_DMYL6H m4_n114303_n17580# m4_n114183_n17460# VSUBS
X0 m4_n114183_n17460# m4_n114303_n17580# cap_mim_2f0fF c_width=100u c_length=100u
C0 m4_n114303_n17580# m4_n114183_n17460# 8.5013f
C1 m4_n114183_n17460# VSUBS 85.381996f
C2 m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ VSUBS cap_mim_2p0fF_DMYL6H
C0 cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# VSUBS 17.2586f
.ends

.subckt cap_mim_2p0fF_RCWXT2$2 m4_n3148_n3000# m4_n3268_n3120# VSUBS
X0 m4_n3148_n3000# m4_n3268_n3120# cap_mim_2f0fF c_width=30u c_length=30u
C0 m4_n3268_n3120# m4_n3148_n3000# 2.57661f
C1 m4_n3148_n3000# VSUBS 9.60519f
C2 m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt mim_cap_30_30$1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000#
+ VSUBS
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120#
+ VSUBS cap_mim_2p0fF_RCWXT2$2
C0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# VSUBS 9.60519f
C1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# VSUBS 5.38044f
.ends

.subckt cap_mim_2p0fF_DMYL6H$1 m4_93823_n2660# m4_93943_n2540# VSUBS
X0 m4_93943_n2540# m4_93823_n2660# cap_mim_2f0fF c_width=100u c_length=100u
C0 m4_93823_n2660# m4_93943_n2540# 8.5013f
C1 m4_93943_n2540# VSUBS 85.381996f
C2 m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap_100_100$1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ VSUBS cap_mim_2p0fF_DMYL6H$1
C0 cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540# VSUBS 85.381996f
C1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# VSUBS 17.2586f
.ends

.subckt mim_cap2 vss vdd VSUBS
Xmim_cap_100_100_0 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_1 vss vdd VSUBS mim_cap_100_100
Xmim_cap_100_100_2 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_20 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_0 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_3 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_21 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_22 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_1 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_10 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_11 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100_4 vss vdd VSUBS mim_cap_100_100
Xmim_cap_30_30$1_23 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_2 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_12 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_24 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_3 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_13 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_4 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_14 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_5 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_6 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_15 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_16 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_7 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_8 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_17 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_9 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_18 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_30_30$1_19 vss vdd VSUBS mim_cap_30_30$1
Xmim_cap_100_100$1_0 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_1 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_2 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_3 vss vdd VSUBS mim_cap_100_100$1
Xmim_cap_100_100$1_4 vss vdd VSUBS mim_cap_100_100$1
C0 vss vdd 0.263674p
C1 vdd VSUBS 1.472734p
C2 vss VSUBS 0.651945p
.ends

.subckt mim_cap_boss vss vdd VSUBS
Xmim_cap1_0 vss vdd VSUBS mim_cap1
Xmim_cap2_0 vss vdd VSUBS mim_cap2
C0 vdd vss 1.238065p
C1 vdd VSUBS 6.097546p
C2 vss VSUBS 3.284302p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VPW VNW a_36_472# a_572_375# a_124_375#
+ a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VDD VNW 0.11314f
C1 a_36_472# a_124_375# 0.285629f
C2 VSS a_484_472# 0.148682f
C3 a_572_375# a_124_375# 0.012222f
C4 VDD a_484_472# 0.179463f
C5 a_124_375# VNW 0.180172f
C6 VDD VSS 0.013184f
C7 a_36_472# VNW 0.025611f
C8 a_572_375# VNW 0.18122f
C9 a_124_375# a_484_472# 0.086742f
C10 a_36_472# a_484_472# 0.013276f
C11 a_572_375# a_484_472# 0.285629f
C12 a_124_375# VSS 0.136476f
C13 a_36_472# VSS 0.151218f
C14 VDD a_124_375# 0.12673f
C15 a_572_375# VSS 0.082563f
C16 a_484_472# VNW 0.024396f
C17 a_36_472# VDD 0.093681f
C18 a_572_375# VDD 0.129266f
C19 VSS VNW 0.008822f
C20 VSS VSUBS 0.360066f
C21 VDD VSUBS 0.286281f
C22 VNW VSUBS 1.65967f
C23 a_484_472# VSUBS 0.345058f
C24 a_36_472# VSUBS 0.404746f
C25 a_572_375# VSUBS 0.232991f
C26 a_124_375# VSUBS 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VPW VNW VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 VNW VDD 0.048519f
C1 VSS VDD 0.009725f
C2 VSS VNW 0.007461f
C3 I VDD 0.017439f
C4 VNW I 0.027206f
C5 VSS I 0.031625f
C6 VSS VSUBS 0.12617f
C7 VDD VSUBS 0.087026f
C8 I VSUBS 0.139667f
C9 VNW VSUBS 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VPW VNW a_224_472# VSUBS
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 a_224_472# A2 0.008979f
C1 ZN A2 0.378409f
C2 a_224_472# ZN 0.023693f
C3 A1 A2 0.037814f
C4 A1 ZN 0.579732f
C5 VSS VDD 0.023219f
C6 VNW VDD 0.093678f
C7 VSS A2 0.043352f
C8 VNW A2 0.128798f
C9 VSS ZN 0.08687f
C10 A1 VSS 0.168633f
C11 VNW ZN 0.019783f
C12 A1 VNW 0.136915f
C13 VDD A2 0.255318f
C14 a_224_472# VDD 0.013964f
C15 VDD ZN 0.117921f
C16 A1 VDD 0.028041f
C17 VSS VNW 0.010571f
C18 VSS VSUBS 0.331491f
C19 ZN VSUBS 0.058886f
C20 VDD VSUBS 0.218051f
C21 A1 VSUBS 0.331856f
C22 A2 VSUBS 0.334514f
C23 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VPW VNW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_1456_156#
+ a_1288_156# a_2248_156# a_2560_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 VSS a_1288_156# 0.001702f
C1 VDD a_2665_112# 0.102046f
C2 VNW Q 0.034443f
C3 a_1000_472# VSS 0.04356f
C4 a_1000_472# a_1308_423# 0.934191f
C5 D a_796_472# 0.082858f
C6 VNW a_448_472# 0.341284f
C7 VSS a_36_151# 0.291264f
C8 a_36_151# a_1308_423# 0.05539f
C9 a_1000_472# a_2248_156# 0.001232f
C10 VNW RN 0.329494f
C11 a_36_151# a_2248_156# 0.042802f
C12 a_2560_156# a_36_151# 0.003674f
C13 VNW a_1204_472# 0.016269f
C14 VNW a_796_472# 0.010232f
C15 a_1000_472# VDD 0.119211f
C16 VSS a_1308_423# 0.013866f
C17 a_36_151# VDD 0.417088f
C18 VSS a_2248_156# 0.030473f
C19 a_1308_423# a_2248_156# 0.056721f
C20 a_2560_156# VSS 0.128503f
C21 a_2560_156# a_2248_156# 0.119687f
C22 VSS VDD 0.01338f
C23 VDD a_1308_423# 0.094185f
C24 VDD a_2248_156# 1.11667f
C25 a_2560_156# VDD 0.00217f
C26 Q a_2665_112# 0.109436f
C27 a_36_151# CLK 0.669598f
C28 a_3041_156# a_2665_112# 0.001774f
C29 VSS a_1456_156# 0.001901f
C30 D VNW 0.128231f
C31 a_448_472# a_2665_112# 0.020455f
C32 a_2665_112# RN 0.336469f
C33 VSS CLK 0.021952f
C34 a_1288_156# a_448_472# 0.002067f
C35 a_1000_472# a_448_472# 0.361958f
C36 VDD CLK 0.02303f
C37 a_36_151# a_448_472# 0.536965f
C38 a_1000_472# RN 0.0832f
C39 a_36_151# RN 0.080102f
C40 VSS Q 0.113401f
C41 a_1000_472# a_1204_472# 0.66083f
C42 a_1000_472# a_796_472# 0.048436f
C43 VSS a_448_472# 1.20207f
C44 Q a_2248_156# 0.014355f
C45 a_36_151# a_1204_472# 0.006996f
C46 a_448_472# a_1308_423# 0.882105f
C47 a_36_151# a_796_472# 0.011851f
C48 VSS RN 0.441968f
C49 a_448_472# a_2248_156# 0.510371f
C50 a_1308_423# RN 0.079294f
C51 a_2560_156# a_448_472# 0.277491f
C52 a_2248_156# RN 0.094336f
C53 VDD Q 0.149344f
C54 VSS a_796_472# 0.05215f
C55 a_1204_472# a_1308_423# 0.026665f
C56 a_2560_156# RN 0.038779f
C57 VDD a_448_472# 0.456269f
C58 VDD RN 0.034984f
C59 VNW a_2665_112# 0.354715f
C60 VDD a_1204_472# 0.282626f
C61 a_448_472# a_1456_156# 0.00227f
C62 D a_36_151# 0.094113f
C63 a_448_472# CLK 0.002757f
C64 a_1000_472# VNW 0.241357f
C65 D VSS 0.064618f
C66 a_36_151# VNW 1.28833f
C67 VSS VNW 0.010602f
C68 VNW a_1308_423# 0.149014f
C69 D VDD 0.009367f
C70 VNW a_2248_156# 0.212431f
C71 a_2560_156# VNW 0.020165f
C72 a_3041_156# RN 0.01068f
C73 a_448_472# RN 0.078731f
C74 VDD VNW 0.503557f
C75 a_1204_472# a_448_472# 0.008996f
C76 a_448_472# a_796_472# 0.401636f
C77 a_1204_472# RN 0.021039f
C78 a_36_151# a_2665_112# 0.019043f
C79 VNW CLK 0.137037f
C80 VSS a_2665_112# 0.184997f
C81 a_2665_112# a_2248_156# 0.633318f
C82 a_1000_472# a_36_151# 0.08126f
C83 a_2560_156# a_2665_112# 0.116059f
C84 D a_448_472# 0.328788f
C85 Q VSUBS 0.114762f
C86 VSS VSUBS 1.26186f
C87 RN VSUBS 1.36673f
C88 D VSUBS 0.253406f
C89 VDD VSUBS 0.79945f
C90 CLK VSUBS 0.291241f
C91 VNW VSUBS 6.1377f
C92 a_2560_156# VSUBS 0.016968f
C93 a_2665_112# VSUBS 0.62251f
C94 a_2248_156# VSUBS 0.371662f
C95 a_1204_472# VSUBS 0.012971f
C96 a_1000_472# VSUBS 0.291735f
C97 a_796_472# VSUBS 0.023206f
C98 a_1308_423# VSUBS 0.279043f
C99 a_448_472# VSUBS 0.684413f
C100 a_36_151# VSUBS 1.43589f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VPW VNW a_36_68# a_244_472#
+ a_692_472# VSUBS
X0 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 B2 a_244_472# 0.002003f
C1 B1 a_244_472# 0.003598f
C2 ZN VDD 0.004634f
C3 A2 A1 0.038725f
C4 VNW A2 0.125671f
C5 A2 ZN 0.390894f
C6 VSS VDD 0.011512f
C7 a_36_68# A1 0.160084f
C8 a_692_472# VDD 0.004194f
C9 VNW a_36_68# 0.040298f
C10 B1 B2 0.036483f
C11 ZN a_36_68# 0.419486f
C12 A2 VSS 0.087422f
C13 VSS a_36_68# 0.392965f
C14 A2 VDD 0.019572f
C15 a_692_472# a_36_68# 0.015646f
C16 B1 A1 0.163724f
C17 VNW B2 0.133721f
C18 VNW B1 0.125926f
C19 a_36_68# VDD 0.787847f
C20 ZN B1 0.079f
C21 VDD a_244_472# 0.00636f
C22 A2 a_36_68# 0.340509f
C23 VSS B2 0.025295f
C24 B1 VSS 0.025138f
C25 VNW A1 0.115376f
C26 ZN A1 0.430191f
C27 VNW ZN 0.010694f
C28 B2 VDD 0.246452f
C29 a_36_68# a_244_472# 0.027448f
C30 B1 VDD 0.014643f
C31 VSS A1 0.084232f
C32 VNW VSS 0.010714f
C33 ZN VSS 0.085273f
C34 a_692_472# ZN 0.011665f
C35 VDD A1 0.014671f
C36 a_36_68# B2 0.369561f
C37 B1 a_36_68# 0.437534f
C38 VNW VDD 0.139306f
C39 VSS VSUBS 0.383233f
C40 ZN VSUBS 0.012598f
C41 VDD VSUBS 0.318857f
C42 A2 VSUBS 0.2826f
C43 A1 VSUBS 0.258579f
C44 B1 VSUBS 0.257485f
C45 B2 VSUBS 0.309037f
C46 VNW VSUBS 2.00777f
C47 a_36_68# VSUBS 0.150048f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VPW VNW a_49_472#
+ a_665_69# a_257_69# VSUBS
X0 ZN B1 a_257_69# VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
C0 A1 a_665_69# 0.002008f
C1 a_49_472# B1 0.069833f
C2 VNW VDD 0.112326f
C3 ZN B1 0.367665f
C4 A1 A2 0.392541f
C5 A1 a_49_472# 0.021757f
C6 A2 a_665_69# 0.006702f
C7 VSS VDD 0.00787f
C8 A1 ZN 0.447732f
C9 ZN a_665_69# 0.001059f
C10 VNW VSS 0.011011f
C11 A2 a_49_472# 0.075759f
C12 VDD B2 0.026097f
C13 A2 ZN 0.102518f
C14 VNW B2 0.129409f
C15 ZN a_49_472# 0.239204f
C16 VSS B2 0.06757f
C17 VDD B1 0.017923f
C18 VNW B1 0.109456f
C19 A1 VDD 0.013859f
C20 a_257_69# VSS 0.00576f
C21 VNW A1 0.10965f
C22 VSS B1 0.095385f
C23 a_257_69# B2 0.003563f
C24 A2 VDD 0.013575f
C25 VDD a_49_472# 0.887006f
C26 B1 B2 0.18297f
C27 A1 VSS 0.087393f
C28 a_665_69# VSS 0.003829f
C29 VNW A2 0.131727f
C30 VNW a_49_472# 0.026629f
C31 ZN VDD 0.004108f
C32 VNW ZN 0.017894f
C33 A2 VSS 0.150463f
C34 VSS a_49_472# 0.02154f
C35 a_257_69# B1 0.003901f
C36 ZN VSS 0.071892f
C37 a_49_472# B2 0.151151f
C38 ZN B2 0.001886f
C39 A1 B1 0.041046f
C40 VSS VSUBS 0.39457f
C41 ZN VSUBS 0.021794f
C42 VDD VSUBS 0.243433f
C43 A2 VSUBS 0.322629f
C44 A1 VSUBS 0.250967f
C45 B1 VSUBS 0.261124f
C46 B2 VSUBS 0.322244f
C47 VNW VSUBS 1.83372f
C48 a_49_472# VSUBS 0.054843f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VPW VNW a_36_160# VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VDD VNW 0.087464f
C1 a_36_160# Z 0.281838f
C2 I a_36_160# 0.545454f
C3 I Z 0.041707f
C4 VSS VNW 0.009324f
C5 VDD a_36_160# 0.2736f
C6 VDD Z 0.128274f
C7 VDD I 0.02612f
C8 VSS a_36_160# 0.074156f
C9 VSS Z 0.146199f
C10 VNW a_36_160# 0.170864f
C11 VNW Z 0.030347f
C12 VSS I 0.12329f
C13 VNW I 0.2276f
C14 VDD VSS 0.009574f
C15 VSS VSUBS 0.28275f
C16 Z VSUBS 0.10469f
C17 VDD VSUBS 0.178615f
C18 I VSUBS 0.323491f
C19 VNW VSUBS 1.31158f
C20 a_36_160# VSUBS 0.386641f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD ZN 0.098026f
C1 VDD VNW 0.076212f
C2 I VSS 0.058937f
C3 I ZN 0.47009f
C4 ZN VSS 0.077008f
C5 VNW I 0.135368f
C6 VNW VSS 0.011085f
C7 VDD I 0.157124f
C8 VDD VSS 0.025441f
C9 VNW ZN 0.031181f
C10 VSS VSUBS 0.242183f
C11 ZN VSUBS 0.095505f
C12 VDD VSUBS 0.182097f
C13 I VSUBS 0.355642f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VDD ZN 0.137375f
C1 VDD VNW 0.076257f
C2 I VSS 0.0533f
C3 I ZN 0.262199f
C4 ZN VSS 0.115297f
C5 VNW I 0.137757f
C6 VNW VSS 0.011339f
C7 VDD I 0.041847f
C8 VDD VSS 0.025626f
C9 VNW ZN 0.022202f
C10 VSS VSUBS 0.2316f
C11 ZN VSUBS 0.113404f
C12 VDD VSUBS 0.181139f
C13 I VSUBS 0.341982f
C14 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VPW VNW a_36_472# a_124_375# VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VNW VDD 0.061035f
C1 VNW a_124_375# 0.179924f
C2 a_36_472# VSS 0.150876f
C3 a_36_472# VDD 0.093681f
C4 VDD VSS 0.006592f
C5 a_124_375# a_36_472# 0.285629f
C6 a_124_375# VSS 0.082879f
C7 VNW a_36_472# 0.025989f
C8 VNW VSS 0.004411f
C9 a_124_375# VDD 0.126034f
C10 VSS VSUBS 0.218985f
C11 VDD VSUBS 0.182777f
C12 VNW VSUBS 0.96348f
C13 a_36_472# VSUBS 0.417394f
C14 a_124_375# VSUBS 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VPW VNW a_224_472# VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 I VDD 0.1311f
C1 VSS VDD 0.031131f
C2 I a_224_472# 0.796069f
C3 VNW Z 0.038011f
C4 VSS a_224_472# 0.659695f
C5 I VSS 0.158668f
C6 VNW VDD 0.305516f
C7 VDD Z 0.819024f
C8 a_224_472# VNW 1.14633f
C9 a_224_472# Z 2.29481f
C10 I VNW 0.55539f
C11 I Z 0.001907f
C12 VSS VNW 0.01282f
C13 VSS Z 0.70427f
C14 a_224_472# VDD 0.74621f
C15 VSS VSUBS 0.910368f
C16 Z VSUBS 0.18914f
C17 VDD VSUBS 0.724491f
C18 I VSUBS 1.16773f
C19 VNW VSUBS 4.79254f
C20 a_224_472# VSUBS 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VPW VNW a_36_472# a_244_68#
+ VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VSUBS nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
C0 A1 VSS 0.021732f
C1 A2 ZN 0.248411f
C2 ZN a_36_472# 0.088503f
C3 VNW VSS 0.009145f
C4 A2 a_36_472# 0.10395f
C5 VDD VSS 0.01275f
C6 ZN A1 0.245346f
C7 B VSS 0.080416f
C8 A2 A1 0.047589f
C9 VNW ZN 0.014655f
C10 A1 a_36_472# 0.104556f
C11 A2 VNW 0.128282f
C12 VDD ZN 0.003129f
C13 VNW a_36_472# 0.013943f
C14 VSS a_244_68# 0.00255f
C15 VDD A2 0.015143f
C16 B ZN 0.00761f
C17 VDD a_36_472# 0.581285f
C18 B a_36_472# 0.01027f
C19 VNW A1 0.122087f
C20 ZN a_244_68# 0.008784f
C21 VDD A1 0.0167f
C22 VDD VNW 0.11216f
C23 B A1 0.157699f
C24 ZN VSS 0.304078f
C25 A2 VSS 0.069479f
C26 B VNW 0.137038f
C27 a_36_472# VSS 0.004325f
C28 VDD B 0.071777f
C29 VSS VSUBS 0.361309f
C30 VDD VSUBS 0.259458f
C31 ZN VSUBS 0.040013f
C32 B VSUBS 0.378232f
C33 A1 VSUBS 0.264815f
C34 A2 VSUBS 0.3189f
C35 VNW VSUBS 1.65967f
C36 a_36_472# VSUBS 0.031137f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VPW VNW a_36_113# VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VDD a_36_113# 0.278283f
C1 Z I 0.031362f
C2 VSS VNW 0.009307f
C3 VSS a_36_113# 0.11114f
C4 VDD Z 0.085355f
C5 VSS Z 0.136942f
C6 VDD I 0.028968f
C7 VSS I 0.070302f
C8 VNW a_36_113# 0.160792f
C9 VSS VDD 0.009561f
C10 Z VNW 0.030118f
C11 Z a_36_113# 0.191876f
C12 I VNW 0.152645f
C13 I a_36_113# 0.476912f
C14 VDD VNW 0.088196f
C15 VSS VSUBS 0.283681f
C16 Z VSUBS 0.117185f
C17 VDD VSUBS 0.180237f
C18 I VSUBS 0.336876f
C19 VNW VSUBS 1.31158f
C20 a_36_113# VSUBS 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VPW VNW a_1916_375# a_1380_472#
+ a_3260_375# a_36_472# a_932_472# a_2812_375# a_2276_472# a_1828_472# a_3172_472#
+ a_572_375# a_2724_472# a_124_375# a_1468_375# a_1020_375# a_484_472# a_2364_375#
+ VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 VNW a_1468_375# 0.181468f
C1 VDD a_36_472# 0.093681f
C2 VDD a_1380_472# 0.179463f
C3 a_2364_375# VSS 0.131736f
C4 a_572_375# VSS 0.131736f
C5 VDD a_1020_375# 0.129962f
C6 VSS a_36_472# 0.142026f
C7 VDD a_2812_375# 0.129962f
C8 VSS a_1380_472# 0.142721f
C9 VNW a_484_472# 0.024018f
C10 VSS a_1020_375# 0.131736f
C11 VSS a_2812_375# 0.131736f
C12 a_3260_375# a_2812_375# 0.013103f
C13 a_1916_375# a_1468_375# 0.013103f
C14 a_1828_472# VDD 0.179463f
C15 a_1828_472# VSS 0.142721f
C16 a_2364_375# VNW 0.181468f
C17 a_572_375# VNW 0.181468f
C18 VNW a_36_472# 0.025611f
C19 VDD a_2724_472# 0.179463f
C20 VDD a_932_472# 0.179463f
C21 VNW a_1380_472# 0.024018f
C22 VNW a_1020_375# 0.181468f
C23 a_2724_472# VSS 0.142721f
C24 VNW a_2812_375# 0.181468f
C25 VSS a_932_472# 0.142721f
C26 a_3172_472# a_2812_375# 0.087174f
C27 VDD VSS 0.052737f
C28 a_2364_375# a_1916_375# 0.013103f
C29 VDD a_3260_375# 0.129266f
C30 a_1828_472# VNW 0.024018f
C31 a_3260_375# VSS 0.081304f
C32 a_124_375# a_484_472# 0.087174f
C33 a_2724_472# VNW 0.024018f
C34 VNW a_932_472# 0.024018f
C35 a_3172_472# a_2724_472# 0.013276f
C36 VDD VNW 0.425768f
C37 a_1828_472# a_1916_375# 0.285629f
C38 VSS VNW 0.035286f
C39 a_2364_375# a_2276_472# 0.285629f
C40 a_3172_472# VDD 0.179463f
C41 a_3260_375# VNW 0.18122f
C42 a_572_375# a_124_375# 0.013103f
C43 a_3172_472# VSS 0.139489f
C44 a_124_375# a_36_472# 0.285629f
C45 a_3172_472# a_3260_375# 0.285629f
C46 VDD a_1916_375# 0.129962f
C47 VSS a_1916_375# 0.131736f
C48 a_1828_472# a_2276_472# 0.013276f
C49 a_1380_472# a_1468_375# 0.285629f
C50 a_1020_375# a_1468_375# 0.013103f
C51 a_572_375# a_484_472# 0.285629f
C52 a_36_472# a_484_472# 0.013276f
C53 a_3172_472# VNW 0.024396f
C54 a_2724_472# a_2276_472# 0.013276f
C55 VDD a_2276_472# 0.179463f
C56 VNW a_1916_375# 0.181468f
C57 VSS a_2276_472# 0.142721f
C58 a_1828_472# a_1468_375# 0.087174f
C59 VDD a_124_375# 0.12673f
C60 VSS a_124_375# 0.131736f
C61 a_572_375# a_1020_375# 0.013103f
C62 a_2364_375# a_2812_375# 0.013103f
C63 a_1020_375# a_1380_472# 0.087174f
C64 a_932_472# a_484_472# 0.013276f
C65 VDD a_1468_375# 0.129962f
C66 VSS a_1468_375# 0.131736f
C67 VDD a_484_472# 0.179463f
C68 VNW a_2276_472# 0.024018f
C69 VSS a_484_472# 0.142721f
C70 a_124_375# VNW 0.180172f
C71 a_1828_472# a_1380_472# 0.013276f
C72 a_2364_375# a_2724_472# 0.087174f
C73 a_572_375# a_932_472# 0.087174f
C74 a_932_472# a_1380_472# 0.013276f
C75 a_932_472# a_1020_375# 0.285629f
C76 a_2724_472# a_2812_375# 0.285629f
C77 VDD a_2364_375# 0.129962f
C78 VDD a_572_375# 0.129962f
C79 a_1916_375# a_2276_472# 0.087174f
C80 VSS VSUBS 1.20585f
C81 VDD VSUBS 0.907304f
C82 VNW VSUBS 5.83682f
C83 a_3172_472# VSUBS 0.345058f
C84 a_2724_472# VSUBS 0.33241f
C85 a_2276_472# VSUBS 0.33241f
C86 a_1828_472# VSUBS 0.33241f
C87 a_1380_472# VSUBS 0.33241f
C88 a_932_472# VSUBS 0.33241f
C89 a_484_472# VSUBS 0.33241f
C90 a_36_472# VSUBS 0.404746f
C91 a_3260_375# VSUBS 0.233093f
C92 a_2812_375# VSUBS 0.17167f
C93 a_2364_375# VSUBS 0.17167f
C94 a_1916_375# VSUBS 0.17167f
C95 a_1468_375# VSUBS 0.17167f
C96 a_1020_375# VSUBS 0.17167f
C97 a_572_375# VSUBS 0.17167f
C98 a_124_375# VSUBS 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VPW VNW a_455_68# a_271_68#
+ VSUBS
X0 ZN A1 a_455_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 A2 a_271_68# 0.004027f
C1 VNW VDD 0.112537f
C2 VNW VSS 0.008577f
C3 ZN a_271_68# 0.001916f
C4 A2 A1 0.133044f
C5 VSS a_271_68# 0.006038f
C6 VNW A3 0.148237f
C7 ZN A1 0.384588f
C8 A1 VDD 0.022021f
C9 VSS A1 0.084906f
C10 ZN A2 0.078589f
C11 a_455_68# A1 0.004981f
C12 A2 VDD 0.023177f
C13 VNW A1 0.12917f
C14 A2 VSS 0.104901f
C15 ZN VDD 0.33173f
C16 ZN VSS 0.064021f
C17 VSS VDD 0.008734f
C18 A2 A3 0.117566f
C19 a_455_68# A2 0.005127f
C20 A2 VNW 0.121191f
C21 ZN A3 0.008403f
C22 ZN a_455_68# 0.002926f
C23 A3 VDD 0.079999f
C24 VSS A3 0.07804f
C25 ZN VNW 0.034322f
C26 a_455_68# VSS 0.006909f
C27 VSS VSUBS 0.307914f
C28 ZN VSUBS 0.133449f
C29 VDD VSUBS 0.241872f
C30 A1 VSUBS 0.287469f
C31 A2 VSUBS 0.25736f
C32 A3 VSUBS 0.326833f
C33 VNW VSUBS 1.48562f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VPW VNW a_245_68# VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
C0 VNW ZN 0.02653f
C1 VSS A1 0.131667f
C2 VDD ZN 0.240333f
C3 ZN A1 0.351362f
C4 a_245_68# A1 0.008831f
C5 ZN VSS 0.098328f
C6 A2 VNW 0.125396f
C7 a_245_68# VSS 0.002295f
C8 A2 VDD 0.039698f
C9 A2 A1 0.226398f
C10 VNW VDD 0.084263f
C11 A2 VSS 0.051087f
C12 VNW A1 0.119756f
C13 VNW VSS 0.006174f
C14 VDD A1 0.027485f
C15 A2 ZN 0.038658f
C16 VDD VSS 0.017706f
C17 VSS VSUBS 0.238729f
C18 ZN VSUBS 0.105772f
C19 VDD VSUBS 0.243067f
C20 A1 VSUBS 0.290957f
C21 A2 VSUBS 0.314823f
C22 VNW VSUBS 1.13753f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VPW VNW a_255_603# a_67_603#
+ VSUBS
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 A1 VNW 0.220003f
C1 VSS VNW 0.010039f
C2 VDD a_67_603# 0.307039f
C3 VDD A2 0.147628f
C4 VDD Z 0.196046f
C5 A1 VSS 0.050738f
C6 VDD a_255_603# 0.005359f
C7 a_67_603# VNW 0.157241f
C8 A2 VNW 0.216313f
C9 Z VNW 0.033884f
C10 A1 a_67_603# 0.540888f
C11 A1 A2 0.062395f
C12 VSS a_67_603# 0.250493f
C13 VSS A2 0.025748f
C14 VSS Z 0.158265f
C15 VDD VNW 0.11771f
C16 a_67_603# A2 0.505374f
C17 Z a_67_603# 0.181586f
C18 a_255_603# a_67_603# 0.007617f
C19 A1 VDD 0.01431f
C20 Z A2 0.027598f
C21 a_255_603# A2 0.001961f
C22 VDD VSS 0.008648f
C23 VSS VSUBS 0.359722f
C24 Z VSUBS 0.102754f
C25 VDD VSUBS 0.233025f
C26 A2 VSUBS 0.313441f
C27 A1 VSUBS 0.39469f
C28 VNW VSUBS 1.65967f
C29 a_67_603# VSUBS 0.345683f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VPW VNW a_36_68# a_1612_497#
+ a_2124_68# a_244_497# a_2960_68# a_3368_68# a_2552_68# a_1164_497# a_716_497# VSUBS
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
C0 a_1164_497# A2 0.009095f
C1 a_36_68# A2 0.108262f
C2 A1 VSS 0.060963f
C3 ZN VDD 2.06829f
C4 a_716_497# A2 0.00653f
C5 ZN a_1612_497# 0.024559f
C6 A1 ZN 1.37575f
C7 VSS VNW 0.004483f
C8 a_2960_68# a_36_68# 0.009506f
C9 a_36_68# VSS 3.64719f
C10 a_36_68# a_3368_68# 0.007478f
C11 a_36_68# a_2124_68# 0.012118f
C12 VSS C 0.092809f
C13 ZN VNW 0.056895f
C14 a_36_68# a_2552_68# 0.009506f
C15 ZN a_1164_497# 0.021094f
C16 VSS A2 0.060501f
C17 VDD B 0.100578f
C18 ZN a_36_68# 1.98502f
C19 a_244_497# A2 0.01347f
C20 ZN a_716_497# 0.027752f
C21 ZN C 0.514613f
C22 ZN A2 1.2828f
C23 a_2960_68# VSS 0.002422f
C24 a_1612_497# VDD 0.009792f
C25 VSS a_3368_68# 0.004815f
C26 a_2124_68# VSS 0.004133f
C27 A1 VDD 0.078657f
C28 VNW B 0.600992f
C29 VSS a_2552_68# 0.002422f
C30 a_36_68# B 1.37417f
C31 ZN VSS 0.006216f
C32 ZN a_244_497# 0.009475f
C33 C B 1.73339f
C34 VNW VDD 0.366897f
C35 A2 B 0.037299f
C36 VDD a_1164_497# 0.008664f
C37 a_36_68# VDD 0.021485f
C38 A1 VNW 0.51833f
C39 a_716_497# VDD 0.008599f
C40 C VDD 0.095093f
C41 A1 a_36_68# 0.065645f
C42 VDD A2 0.15752f
C43 a_2960_68# B 0.002626f
C44 a_1612_497# A2 0.010709f
C45 VSS B 0.072527f
C46 A1 A2 1.73987f
C47 a_36_68# VNW 0.004654f
C48 a_2552_68# B 0.002588f
C49 ZN B 0.426118f
C50 VSS VDD 0.005699f
C51 VNW C 0.636287f
C52 a_244_497# VDD 0.020528f
C53 VNW A2 0.590323f
C54 a_36_68# C 0.105844f
C55 VSS VSUBS 1.08055f
C56 ZN VSUBS 0.051826f
C57 VDD VSUBS 0.846798f
C58 C VSUBS 1.06351f
C59 B VSUBS 1.11555f
C60 A1 VSUBS 1.1956f
C61 A2 VSUBS 1.16629f
C62 VNW VSUBS 5.892971f
C63 a_36_68# VSUBS 0.063181f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VPW VNW a_36_160# VSUBS
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VSUBS nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VSUBS nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
C0 a_36_160# I 0.564508f
C1 VDD I 0.028233f
C2 VNW VSS 0.00834f
C3 VSS a_36_160# 0.114407f
C4 VNW a_36_160# 0.302514f
C5 VSS VDD 0.01316f
C6 VNW VDD 0.111398f
C7 Z I 0.016176f
C8 a_36_160# VDD 0.31851f
C9 VNW Z 0.021185f
C10 VSS Z 0.111496f
C11 a_36_160# Z 0.426617f
C12 VSS I 0.178818f
C13 VNW I 0.1633f
C14 VDD Z 0.161733f
C15 VSS VSUBS 0.397291f
C16 Z VSUBS 0.097163f
C17 VDD VSUBS 0.238155f
C18 I VSUBS 0.333888f
C19 VNW VSUBS 1.65967f
C20 a_36_160# VSUBS 0.696445f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VPW VNW a_1380_472# a_36_472#
+ a_932_472# a_572_375# a_124_375# a_1468_375# a_1020_375# a_484_472# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 VSS a_484_472# 0.148077f
C1 a_484_472# VNW 0.024018f
C2 VDD a_1020_375# 0.129962f
C3 a_572_375# VSS 0.134699f
C4 a_124_375# VSS 0.134699f
C5 VDD a_1380_472# 0.179463f
C6 VSS a_932_472# 0.148077f
C7 a_572_375# VNW 0.181468f
C8 a_124_375# VNW 0.180172f
C9 a_932_472# VNW 0.024018f
C10 a_1468_375# a_1020_375# 0.012552f
C11 a_1380_472# a_1468_375# 0.285629f
C12 a_572_375# a_1020_375# 0.012552f
C13 VDD a_36_472# 0.093681f
C14 a_1020_375# a_932_472# 0.285629f
C15 VDD a_1468_375# 0.129266f
C16 a_1380_472# a_932_472# 0.013276f
C17 VDD a_484_472# 0.179463f
C18 a_36_472# a_484_472# 0.013276f
C19 a_572_375# VDD 0.129962f
C20 VDD a_124_375# 0.12673f
C21 VDD a_932_472# 0.179463f
C22 a_124_375# a_36_472# 0.285629f
C23 VSS VNW 0.017643f
C24 a_572_375# a_484_472# 0.285629f
C25 a_124_375# a_484_472# 0.086905f
C26 a_932_472# a_484_472# 0.013276f
C27 a_572_375# a_124_375# 0.012552f
C28 a_572_375# a_932_472# 0.086905f
C29 VSS a_1020_375# 0.134699f
C30 a_1020_375# VNW 0.181468f
C31 a_1380_472# VSS 0.144845f
C32 a_1380_472# VNW 0.024396f
C33 VDD VSS 0.026369f
C34 VDD VNW 0.217349f
C35 a_36_472# VSS 0.147381f
C36 a_1380_472# a_1020_375# 0.086905f
C37 a_36_472# VNW 0.025611f
C38 VSS a_1468_375# 0.082091f
C39 a_1468_375# VNW 0.18122f
C40 VSS VSUBS 0.642184f
C41 VDD VSUBS 0.493288f
C42 VNW VSUBS 3.05206f
C43 a_1380_472# VSUBS 0.345058f
C44 a_932_472# VSUBS 0.33241f
C45 a_484_472# VSUBS 0.33241f
C46 a_36_472# VSUBS 0.404746f
C47 a_1468_375# VSUBS 0.233029f
C48 a_1020_375# VSUBS 0.171606f
C49 a_572_375# VSUBS 0.171606f
C50 a_124_375# VSUBS 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VPW VNW a_36_68# VSUBS
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VSUBS nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 VDD VSS 0.014283f
C1 Z I 0.018906f
C2 Z a_36_68# 0.432914f
C3 VDD I 0.029139f
C4 VDD a_36_68# 0.271105f
C5 I VSS 0.128735f
C6 VSS a_36_68# 0.156367f
C7 VNW Z 0.023138f
C8 I a_36_68# 0.731677f
C9 VNW VDD 0.114912f
C10 VNW VSS 0.009972f
C11 Z VDD 0.172592f
C12 VNW I 0.133333f
C13 VNW a_36_68# 0.296832f
C14 Z VSS 0.133443f
C15 VSS VSUBS 0.338876f
C16 Z VSUBS 0.103236f
C17 VDD VSUBS 0.234026f
C18 I VSUBS 0.298844f
C19 VNW VSUBS 1.65967f
C20 a_36_68# VSUBS 0.69549f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VPW VNW a_848_380# a_1084_68#
+ a_124_24# a_1152_472# a_692_472# VSUBS
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VSUBS nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VSUBS nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
C0 a_848_380# S 0.754833f
C1 VDD S 0.056165f
C2 a_124_24# a_1084_68# 0.002839f
C3 a_848_380# VNW 0.174516f
C4 a_848_380# VSS 0.130064f
C5 VDD VNW 0.182986f
C6 VDD VSS 0.028952f
C7 Z I1 0.027341f
C8 a_848_380# a_692_472# 0.003985f
C9 a_124_24# a_1152_472# 0.00128f
C10 VDD a_692_472# 0.009663f
C11 a_124_24# a_848_380# 0.302602f
C12 a_124_24# VDD 0.309232f
C13 I0 a_1084_68# 0.00492f
C14 S VNW 0.253706f
C15 S VSS 0.081531f
C16 VSS VNW 0.009598f
C17 a_848_380# I1 0.013444f
C18 a_692_472# S 0.002582f
C19 a_848_380# I0 0.082224f
C20 VDD I1 0.227359f
C21 I0 VDD 0.028914f
C22 a_124_24# S 0.245829f
C23 a_124_24# VNW 0.277682f
C24 a_124_24# VSS 0.501844f
C25 Z VDD 0.20273f
C26 a_124_24# a_692_472# 0.033243f
C27 I1 S 0.042269f
C28 I0 S 0.533789f
C29 a_692_68# VSS 0.001982f
C30 I1 VNW 0.127749f
C31 I1 VSS 0.026996f
C32 I0 VNW 0.103064f
C33 I0 VSS 0.124513f
C34 a_848_380# a_1152_472# 0.007362f
C35 a_1152_472# VDD 0.00645f
C36 a_692_472# I1 0.001219f
C37 Z VNW 0.020389f
C38 a_848_380# VDD 0.319708f
C39 Z VSS 0.129676f
C40 a_124_24# a_692_68# 0.006853f
C41 a_124_24# I1 0.564972f
C42 a_124_24# I0 0.004772f
C43 a_1084_68# S 0.001644f
C44 a_1084_68# VSS 0.009508f
C45 a_124_24# Z 0.219295f
C46 VSS VSUBS 0.565512f
C47 Z VSUBS 0.047467f
C48 VDD VSUBS 0.424967f
C49 I0 VSUBS 0.267152f
C50 S VSUBS 0.549493f
C51 I1 VSUBS 0.247562f
C52 VNW VSUBS 2.87801f
C53 a_848_380# VSUBS 0.40208f
C54 a_124_24# VSUBS 0.591898f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VPW VNW a_36_68# a_244_472#
+ VSUBS
X0 VSS B a_36_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 a_244_472# VDD 0.004051f
C1 B VDD 0.07579f
C2 a_36_68# ZN 0.56857f
C3 A1 VDD 0.014914f
C4 B VNW 0.163023f
C5 VNW A1 0.117811f
C6 a_36_68# A2 0.489122f
C7 A2 ZN 0.400775f
C8 a_36_68# VSS 0.117681f
C9 VSS ZN 0.088946f
C10 B A1 0.034707f
C11 A2 VSS 0.083821f
C12 a_36_68# VDD 0.753239f
C13 ZN VDD 0.006004f
C14 a_36_68# VNW 0.038286f
C15 VNW ZN 0.011308f
C16 A2 VDD 0.017122f
C17 A2 VNW 0.122386f
C18 VSS VDD 0.004855f
C19 a_36_68# a_244_472# 0.013419f
C20 VSS VNW 0.0064f
C21 ZN a_244_472# 0.014146f
C22 a_36_68# B 0.389329f
C23 a_36_68# A1 0.292244f
C24 ZN A1 0.496662f
C25 VNW VDD 0.117098f
C26 A2 A1 0.038725f
C27 B VSS 0.198567f
C28 VSS A1 0.090903f
C29 VSS VSUBS 0.342662f
C30 ZN VSUBS 0.011384f
C31 VDD VSUBS 0.256635f
C32 B VSUBS 0.339176f
C33 A1 VSUBS 0.256004f
C34 A2 VSUBS 0.28395f
C35 VNW VSUBS 1.65967f
C36 a_36_68# VSUBS 0.112263f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VPW VNW a_224_552# VSUBS
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
C0 a_224_552# VSS 0.331404f
C1 VNW VSS 0.009226f
C2 VDD a_224_552# 0.347549f
C3 Z VSS 0.275062f
C4 VDD VNW 0.176912f
C5 VDD Z 0.356369f
C6 I a_224_552# 0.421587f
C7 I VNW 0.376531f
C8 I Z 0.002319f
C9 a_224_552# VNW 0.5926f
C10 a_224_552# Z 1.17071f
C11 Z VNW 0.027266f
C12 VDD VSS 0.030201f
C13 I VSS 0.061715f
C14 VDD I 0.069894f
C15 VSS VSUBS 0.628617f
C16 Z VSUBS 0.102362f
C17 VDD VSUBS 0.415149f
C18 I VSUBS 0.471574f
C19 VNW VSUBS 2.70396f
C20 a_224_552# VSUBS 1.31114f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VPW VNW a_234_472# a_672_472#
+ VSUBS
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 a_234_472# VDD 0.0121f
C1 ZN VNW 0.03148f
C2 VSS A2 0.07211f
C3 A2 VDD 0.13595f
C4 VSS VDD 0.023993f
C5 A1 A2 0.636124f
C6 VSS A1 0.052992f
C7 A1 VDD 0.037494f
C8 ZN a_672_472# 0.023475f
C9 ZN a_234_472# 0.003154f
C10 ZN A2 0.509001f
C11 ZN VSS 0.460527f
C12 ZN VDD 0.517479f
C13 VNW A2 0.275679f
C14 VSS VNW 0.010681f
C15 VNW VDD 0.137685f
C16 ZN A1 0.274601f
C17 VNW A1 0.25895f
C18 A2 a_672_472# 0.0147f
C19 a_234_472# A2 0.018681f
C20 a_672_472# VDD 0.005379f
C21 VSS VSUBS 0.451405f
C22 ZN VSUBS 0.138491f
C23 VDD VSUBS 0.322159f
C24 A1 VSUBS 0.557317f
C25 A2 VSUBS 0.617688f
C26 VNW VSUBS 2.00777f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VPW VNW a_448_472# a_244_472#
+ VSUBS
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
C0 A3 A2 0.416588f
C1 ZN A3 0.035547f
C2 a_448_472# A2 0.012315f
C3 ZN a_448_472# 0.006209f
C4 A3 VDD 0.201466f
C5 a_448_472# VDD 0.013539f
C6 VNW A3 0.136756f
C7 A1 a_448_472# 0.012619f
C8 VSS A2 0.027728f
C9 ZN VSS 0.283414f
C10 VSS VDD 0.01583f
C11 VSS A1 0.025677f
C12 VNW VSS 0.008407f
C13 a_244_472# A2 0.003952f
C14 ZN a_244_472# 0.001803f
C15 a_244_472# VDD 0.006513f
C16 ZN A2 0.096665f
C17 A2 VDD 0.09496f
C18 A1 A2 0.145555f
C19 A3 VSS 0.058214f
C20 ZN VDD 0.116419f
C21 ZN A1 0.499849f
C22 VNW A2 0.116878f
C23 ZN VNW 0.040402f
C24 A1 VDD 0.095023f
C25 VNW VDD 0.11801f
C26 VNW A1 0.127941f
C27 a_244_472# A3 0.019089f
C28 VSS VSUBS 0.367618f
C29 ZN VSUBS 0.134331f
C30 VDD VSUBS 0.264623f
C31 A1 VSUBS 0.311038f
C32 A2 VSUBS 0.285534f
C33 A3 VSUBS 0.334053f
C34 VNW VSUBS 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VPW VNW a_36_68# a_1732_68#
+ a_244_68# a_1100_68# a_1528_68# a_672_68# VSUBS
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
C0 VSS a_1732_68# 0.002237f
C1 VDD A3 0.107959f
C2 A3 a_1100_68# 0.003385f
C3 A1 a_36_68# 0.118844f
C4 A2 A3 1.65768f
C5 a_1732_68# a_36_68# 0.011094f
C6 VNW A3 0.599629f
C7 VDD ZN 1.57207f
C8 ZN A2 1.77619f
C9 VNW ZN 0.095885f
C10 VDD A2 0.124271f
C11 VSS a_672_68# 0.003125f
C12 VNW VDD 0.292073f
C13 VSS a_244_68# 0.006268f
C14 VNW A2 0.630933f
C15 a_672_68# a_36_68# 0.012389f
C16 VSS A3 0.09506f
C17 a_36_68# a_244_68# 0.009768f
C18 VSS ZN 0.00864f
C19 A3 a_36_68# 1.03106f
C20 VDD VSS 0.004708f
C21 A1 A3 0.001696f
C22 ZN a_36_68# 0.885472f
C23 VSS a_1100_68# 0.003125f
C24 VSS A2 0.070822f
C25 VNW VSS 0.003704f
C26 A1 ZN 1.266f
C27 VDD a_36_68# 0.029088f
C28 a_36_68# a_1100_68# 0.012396f
C29 ZN a_1732_68# 0.002613f
C30 A2 a_36_68# 0.223434f
C31 VNW a_36_68# 0.007741f
C32 A1 VDD 0.115489f
C33 A1 A2 0.077487f
C34 VNW A1 0.700258f
C35 A3 a_672_68# 0.003442f
C36 VSS a_1528_68# 0.003775f
C37 a_1528_68# a_36_68# 0.012072f
C38 VSS a_36_68# 2.77545f
C39 ZN A3 0.150755f
C40 A1 VSS 0.065524f
C41 VSS VSUBS 0.861061f
C42 ZN VSUBS 0.103891f
C43 VDD VSUBS 0.701563f
C44 A1 VSUBS 1.27704f
C45 A3 VSUBS 1.11693f
C46 A2 VSUBS 1.08692f
C47 VNW VSUBS 4.73584f
C48 a_36_68# VSUBS 0.061249f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VPW VNW a_36_159# VSUBS
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VSUBS nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VSUBS nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
C0 VNW a_36_159# 0.162496f
C1 VNW A1 0.206765f
C2 a_244_159# VSS 0.001449f
C3 VDD Z 0.158212f
C4 A2 Z 0.020174f
C5 VDD a_36_159# 0.130189f
C6 Z VSS 0.102819f
C7 A2 a_36_159# 0.472781f
C8 VDD A1 0.04397f
C9 A2 A1 0.061431f
C10 VDD VNW 0.125609f
C11 VNW A2 0.20463f
C12 a_36_159# VSS 0.244357f
C13 a_244_159# a_36_159# 0.003343f
C14 A1 VSS 0.010276f
C15 VNW VSS 0.007925f
C16 Z a_36_159# 0.215269f
C17 VDD A2 0.184025f
C18 VNW Z 0.032842f
C19 VDD VSS 0.014131f
C20 A1 a_36_159# 0.377122f
C21 A2 VSS 0.011099f
C22 VSS VSUBS 0.35312f
C23 Z VSUBS 0.096476f
C24 VDD VSUBS 0.251252f
C25 A2 VSUBS 0.262264f
C26 A1 VSUBS 0.321274f
C27 VNW VSUBS 1.65967f
C28 a_36_159# VSUBS 0.374116f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VPW VNW a_2590_472#
+ a_170_472# a_1602_69# a_786_69# a_3126_472# a_1194_69# a_3662_472# a_2034_472# a_358_69#
+ VSUBS
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VSUBS nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VSUBS nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VSUBS nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VSUBS nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
C0 A2 B 0.05388f
C1 B a_3126_472# 0.007345f
C2 B C 1.34577f
C3 a_2590_472# a_170_472# 0.013379f
C4 VDD a_2590_472# 0.007681f
C5 VNW B 0.617219f
C6 a_170_472# a_2034_472# 0.020753f
C7 VDD a_2034_472# 0.008673f
C8 A2 VNW 0.513788f
C9 a_170_472# A1 0.0698f
C10 VDD A1 0.051939f
C11 a_170_472# VSS 0.00801f
C12 VDD VSS 0.016824f
C13 a_170_472# ZN 0.818521f
C14 VDD ZN 0.008843f
C15 a_358_69# A1 0.001641f
C16 a_1602_69# VSS 0.005669f
C17 a_358_69# VSS 0.005318f
C18 a_1602_69# ZN 0.008113f
C19 a_358_69# ZN 0.011344f
C20 VNW C 0.61926f
C21 VSS a_1194_69# 0.005069f
C22 a_1194_69# ZN 0.00847f
C23 a_3662_472# a_170_472# 0.013628f
C24 VDD a_3662_472# 0.007223f
C25 B a_2590_472# 0.007345f
C26 B a_2034_472# 0.008709f
C27 a_786_69# A1 0.001203f
C28 a_786_69# VSS 0.003966f
C29 a_786_69# ZN 0.008749f
C30 B A1 0.001644f
C31 B VSS 0.119454f
C32 B ZN 0.231932f
C33 A2 A1 1.72617f
C34 A2 VSS 0.104058f
C35 A2 ZN 1.83822f
C36 B a_3662_472# 0.007338f
C37 A1 C 0.001754f
C38 VNW A1 0.480244f
C39 VSS C 0.088883f
C40 VNW VSS 0.012025f
C41 C ZN 1.79111f
C42 VNW ZN 0.045695f
C43 VDD a_170_472# 2.96356f
C44 B a_170_472# 2.12702f
C45 B VDD 0.110239f
C46 VSS A1 0.087217f
C47 A1 ZN 1.40746f
C48 VSS ZN 1.77446f
C49 A2 a_170_472# 0.109943f
C50 A2 VDD 0.052548f
C51 a_3126_472# a_170_472# 0.01307f
C52 a_3126_472# VDD 0.00779f
C53 a_170_472# C 0.075372f
C54 VNW a_170_472# 0.018375f
C55 VDD C 0.089678f
C56 VNW VDD 0.393677f
C57 VSS VSUBS 1.33264f
C58 VDD VSUBS 0.809429f
C59 ZN VSUBS 0.171181f
C60 C VSUBS 1.26656f
C61 B VSUBS 1.19887f
C62 A1 VSUBS 1.12703f
C63 A2 VSUBS 1.09165f
C64 VNW VSUBS 6.53302f
C65 a_170_472# VSUBS 0.077257f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VPW VNW a_1792_472# a_224_472#
+ a_1568_472# a_36_472# a_1120_472# a_672_472# VSUBS
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
C0 a_1120_472# VDD 0.011157f
C1 a_224_472# VDD 0.010911f
C2 VNW a_36_472# 0.031928f
C3 A2 VNW 0.539636f
C4 a_36_472# ZN 0.362263f
C5 A2 ZN 0.250963f
C6 a_1568_472# VDD 0.005385f
C7 a_1792_472# ZN 0.004144f
C8 a_1120_472# a_36_472# 0.01951f
C9 a_224_472# a_36_472# 0.01823f
C10 A2 a_1120_472# 0.002647f
C11 A2 a_224_472# 0.002647f
C12 VNW ZN 0.046016f
C13 A1 a_1568_472# 0.002055f
C14 A3 VSS 0.10353f
C15 A3 VDD 0.09322f
C16 VSS VDD 0.012739f
C17 a_1568_472# a_36_472# 0.025433f
C18 A2 a_1568_472# 0.004974f
C19 A3 A1 0.008795f
C20 A1 VSS 0.115774f
C21 A1 VDD 0.054887f
C22 a_672_472# VDD 0.01105f
C23 A3 a_36_472# 0.100976f
C24 A2 A3 1.6562f
C25 a_36_472# VSS 0.020716f
C26 A2 VSS 0.128956f
C27 a_36_472# VDD 1.90933f
C28 A2 VDD 0.082489f
C29 A3 VNW 0.478769f
C30 a_1792_472# VDD 0.002998f
C31 A1 a_36_472# 0.174868f
C32 A2 A1 0.085569f
C33 VNW VSS 0.009996f
C34 VNW VDD 0.286001f
C35 a_672_472# a_36_472# 0.01823f
C36 A2 a_672_472# 0.002647f
C37 A3 ZN 1.42151f
C38 a_1792_472# A1 0.006624f
C39 VSS ZN 2.18568f
C40 A1 VNW 0.520086f
C41 ZN VDD 0.005367f
C42 A2 a_36_472# 0.993181f
C43 A1 ZN 1.56829f
C44 a_1792_472# a_36_472# 0.022081f
C45 VSS VSUBS 0.918064f
C46 ZN VSUBS 0.159858f
C47 VDD VSUBS 0.61695f
C48 A1 VSUBS 1.35739f
C49 A3 VSUBS 1.33073f
C50 A2 VSUBS 1.29013f
C51 VNW VSUBS 4.79254f
C52 a_36_472# VSUBS 0.137725f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VPW VNW a_468_472# a_244_472#
+ a_1130_472# a_906_472# VSUBS
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 a_244_472# ZN 0.019831f
C1 a_468_472# VDD 0.00502f
C2 VSS ZN 1.3936f
C3 VNW ZN 0.031771f
C4 ZN a_906_472# 0.002855f
C5 A2 VDD 0.038421f
C6 A1 VDD 0.038139f
C7 a_468_472# ZN 0.015602f
C8 A3 a_1130_472# 0.016495f
C9 A3 VDD 0.178286f
C10 A2 ZN 0.694728f
C11 A1 ZN 0.084783f
C12 VSS VNW 0.007164f
C13 VDD a_1130_472# 0.011629f
C14 A3 ZN 1.03634f
C15 VSS A2 0.043139f
C16 a_1130_472# ZN 0.001342f
C17 VSS A1 0.044587f
C18 VDD ZN 0.579119f
C19 A2 VNW 0.241313f
C20 A1 VNW 0.254404f
C21 a_244_472# A3 0.010666f
C22 A3 VSS 0.0525f
C23 A3 VNW 0.28584f
C24 A3 a_906_472# 0.017829f
C25 A2 A1 0.570018f
C26 A3 a_468_472# 0.010018f
C27 a_244_472# VDD 0.00632f
C28 VSS VDD 0.009106f
C29 VDD VNW 0.178574f
C30 VDD a_906_472# 0.011614f
C31 A3 A2 0.624599f
C32 A3 A1 0.292395f
C33 VSS VSUBS 0.509614f
C34 ZN VSUBS 0.172636f
C35 VDD VSUBS 0.441158f
C36 A1 VSUBS 0.622214f
C37 A2 VSUBS 0.627317f
C38 A3 VSUBS 0.692739f
C39 VNW VSUBS 2.70396f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VPW VNW a_1492_488#
+ a_244_68# a_1044_488# a_636_68# a_36_488# VSUBS
X0 VSS B ZN VSUBS nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VSUBS nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
C0 B a_36_488# 0.80489f
C1 VDD a_36_488# 1.67897f
C2 B A2 0.036672f
C3 a_636_68# ZN 0.00593f
C4 VNW VSS 0.008434f
C5 B C 0.560408f
C6 VDD A2 0.02614f
C7 VDD A1 0.026261f
C8 C VDD 0.040747f
C9 VSS ZN 0.708286f
C10 B a_1044_488# 0.012375f
C11 A1 a_244_68# 0.003444f
C12 a_636_68# VSS 0.002222f
C13 VDD a_1044_488# 0.004195f
C14 VNW B 0.298561f
C15 VNW VDD 0.191798f
C16 B ZN 0.413891f
C17 VDD ZN 0.004894f
C18 A2 a_36_488# 0.076279f
C19 A1 a_36_488# 0.031215f
C20 a_1492_488# B 0.007233f
C21 ZN a_244_68# 0.001328f
C22 C a_36_488# 0.041645f
C23 B VSS 0.089442f
C24 A2 A1 0.652956f
C25 a_1492_488# VDD 0.00909f
C26 VSS VDD 0.009527f
C27 a_36_488# a_1044_488# 0.018358f
C28 VSS a_244_68# 0.004878f
C29 VNW a_36_488# 0.010653f
C30 VNW A2 0.280457f
C31 VNW A1 0.25321f
C32 ZN a_36_488# 0.459425f
C33 B VDD 0.04259f
C34 VNW C 0.268332f
C35 ZN A2 0.752866f
C36 ZN A1 0.372797f
C37 C ZN 0.191881f
C38 a_1492_488# a_36_488# 0.017313f
C39 VSS a_36_488# 0.005331f
C40 VSS A2 0.077665f
C41 VSS A1 0.090485f
C42 C VSS 0.05406f
C43 VNW ZN 0.028815f
C44 VSS VSUBS 0.653933f
C45 VDD VSUBS 0.406726f
C46 ZN VSUBS 0.089692f
C47 C VSUBS 0.626227f
C48 B VSUBS 0.654892f
C49 A1 VSUBS 0.552174f
C50 A2 VSUBS 0.559992f
C51 VNW VSUBS 3.2261f
C52 a_36_488# VSUBS 0.101145f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VPW VNW a_244_524# a_2215_68#
+ a_56_524# a_718_524# a_728_93# a_1936_472# a_1336_472# VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
C0 a_1936_472# VDD 0.595117f
C1 a_56_524# A1 0.569057f
C2 a_728_93# VDD 0.575073f
C3 a_1936_472# a_1336_472# 0.004622f
C4 VSS VDD 0.013872f
C5 a_728_93# A2 0.416172f
C6 a_1336_472# a_728_93# 0.62718f
C7 a_1936_472# A3 0.018144f
C8 a_1524_472# a_1336_472# 0.001046f
C9 A2 VSS 0.047538f
C10 a_1936_472# Z 0.337902f
C11 a_1336_472# VSS 0.326133f
C12 a_718_524# a_56_524# 0.009198f
C13 a_728_93# A3 0.720358f
C14 a_1936_472# VNW 0.004015f
C15 a_718_524# A1 0.026418f
C16 a_728_93# Z 0.402606f
C17 VSS A3 0.056027f
C18 a_728_93# VNW 0.346549f
C19 Z VSS 0.277351f
C20 VSS VNW 0.007756f
C21 a_56_524# VDD 0.049641f
C22 a_2215_68# VSS 0.004309f
C23 A1 VDD 0.018915f
C24 A2 a_56_524# 0.908796f
C25 A2 A1 0.321942f
C26 a_718_524# VDD 0.554575f
C27 a_56_524# VNW 0.188846f
C28 VNW A1 0.293766f
C29 a_718_524# A2 0.107911f
C30 a_1936_472# a_728_93# 0.105997f
C31 a_1524_472# a_728_93# 0.007139f
C32 A2 VDD 0.208821f
C33 a_718_524# VNW 0.020055f
C34 a_1336_472# VDD 0.033982f
C35 a_728_93# VSS 0.709567f
C36 a_244_524# VDD 0.004322f
C37 VDD A3 0.028848f
C38 a_1336_472# A2 0.001757f
C39 Z VDD 0.01058f
C40 a_728_93# a_952_93# 0.00421f
C41 a_244_524# A2 0.004824f
C42 VNW VDD 0.360391f
C43 a_1336_472# A3 0.490376f
C44 a_1336_472# Z 0.021039f
C45 A2 VNW 0.369075f
C46 a_1336_472# VNW 0.144065f
C47 a_728_93# a_56_524# 0.016741f
C48 Z A3 0.259021f
C49 a_728_93# A1 0.12992f
C50 VNW A3 0.268193f
C51 a_56_524# VSS 0.214447f
C52 VSS A1 0.139902f
C53 Z VNW 0.028011f
C54 a_2215_68# Z 0.008507f
C55 a_728_93# a_718_524# 0.329834f
C56 VSS VSUBS 0.861752f
C57 Z VSUBS 0.085787f
C58 A1 VSUBS 0.602985f
C59 A2 VSUBS 0.640744f
C60 VDD VSUBS 0.543474f
C61 A3 VSUBS 0.593976f
C62 VNW VSUBS 4.270391f
C63 a_1936_472# VSUBS 0.009918f
C64 a_718_524# VSUBS 0.005143f
C65 a_56_524# VSUBS 0.41096f
C66 a_728_93# VSUBS 0.654825f
C67 a_1336_472# VSUBS 0.316639f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VPW VNW a_652_68# a_244_68#
+ VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
C0 ZN A2 0.891023f
C1 ZN a_652_68# 0.008436f
C2 VSS VDD 0.020712f
C3 A1 A2 0.708017f
C4 VDD VNW 0.123338f
C5 VSS A2 0.057292f
C6 VSS a_652_68# 0.003855f
C7 A2 VNW 0.277885f
C8 ZN A1 0.363066f
C9 ZN a_244_68# 0.001926f
C10 A2 VDD 0.070487f
C11 ZN VSS 0.2597f
C12 a_244_68# A1 0.004867f
C13 ZN VNW 0.033841f
C14 VSS A1 0.115936f
C15 A1 VNW 0.232646f
C16 a_244_68# VSS 0.006834f
C17 VSS VNW 0.008805f
C18 ZN VDD 0.409997f
C19 A1 VDD 0.050088f
C20 VSS VSUBS 0.385688f
C21 ZN VSUBS 0.120217f
C22 VDD VSUBS 0.305683f
C23 A1 VSUBS 0.522064f
C24 A2 VSUBS 0.568932f
C25 VNW VSUBS 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VPW VNW a_36_68# a_1612_497#
+ a_692_497# a_1388_497# a_960_497# VSUBS
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
C0 a_692_497# A2 0.001398f
C1 A2 a_960_497# 0.003506f
C2 A3 a_36_68# 0.036843f
C3 A1 ZN 0.619225f
C4 VNW VDD 0.248379f
C5 VSS VNW 0.008187f
C6 A2 VNW 0.281901f
C7 ZN A3 1.02771f
C8 B VNW 0.309147f
C9 A1 A3 0.206693f
C10 A1 a_1612_497# 0.003158f
C11 a_1612_497# A3 0.030605f
C12 a_1388_497# ZN 0.001168f
C13 a_1388_497# A3 0.02079f
C14 a_36_68# VDD 0.001802f
C15 VSS a_36_68# 2.0408f
C16 A2 a_36_68# 0.032025f
C17 B a_36_68# 0.184521f
C18 ZN VDD 1.08837f
C19 A1 VDD 0.091309f
C20 VSS ZN 0.006088f
C21 ZN A2 0.152712f
C22 A1 VSS 0.032188f
C23 B ZN 0.244028f
C24 A1 A2 0.703324f
C25 A3 VDD 0.555327f
C26 a_1612_497# VDD 0.009412f
C27 VSS A3 0.03178f
C28 A2 A3 1.11591f
C29 B A3 0.036798f
C30 a_1612_497# A2 0.006056f
C31 ZN a_692_497# 0.018589f
C32 a_36_68# VNW 0.001442f
C33 a_1388_497# VDD 0.005409f
C34 ZN a_960_497# 0.012124f
C35 a_1388_497# A2 0.008156f
C36 a_692_497# A3 0.019827f
C37 A3 a_960_497# 0.014254f
C38 ZN VNW 0.025446f
C39 A1 VNW 0.279057f
C40 A3 VNW 0.297068f
C41 VSS VDD 0.010407f
C42 A2 VDD 0.030601f
C43 B VDD 0.119783f
C44 VSS A2 0.030287f
C45 B VSS 0.047409f
C46 a_692_497# VDD 0.00542f
C47 ZN a_36_68# 1.49222f
C48 A1 a_36_68# 0.158235f
C49 a_960_497# VDD 0.003264f
C50 VSS VSUBS 0.663038f
C51 ZN VSUBS 0.080495f
C52 VDD VSUBS 0.512998f
C53 A1 VSUBS 0.643779f
C54 A2 VSUBS 0.561227f
C55 A3 VSUBS 0.573818f
C56 B VSUBS 0.585725f
C57 VNW VSUBS 3.48825f
C58 a_36_68# VSUBS 0.048026f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VPW VNW a_2665_112# a_448_472#
+ a_796_472# a_36_151# a_1204_472# a_3041_156# a_1000_472# a_1308_423# a_2248_156#
+ a_2560_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 VNW a_2665_112# 0.486803f
C1 a_448_472# RN 0.078731f
C2 a_2248_156# RN 0.080362f
C3 a_448_472# a_796_472# 0.401636f
C4 a_448_472# a_2248_156# 0.510371f
C5 CLK VSS 0.021952f
C6 VNW VDD 0.546785f
C7 VNW a_2560_156# 0.019282f
C8 a_2665_112# VSS 0.21484f
C9 VNW a_1308_423# 0.149014f
C10 a_2248_156# Q 0.013765f
C11 VNW a_1000_472# 0.241357f
C12 VNW a_36_151# 1.28833f
C13 a_2665_112# a_3041_156# 0.001841f
C14 VDD VSS 0.02167f
C15 VSS a_1308_423# 0.013866f
C16 a_2560_156# VSS 0.128503f
C17 a_2665_112# RN 0.322698f
C18 VDD a_1204_472# 0.282626f
C19 a_448_472# CLK 0.002757f
C20 a_1204_472# a_1308_423# 0.026665f
C21 VDD D 0.009367f
C22 a_1000_472# VSS 0.04356f
C23 a_448_472# a_2665_112# 0.020455f
C24 a_36_151# VSS 0.291264f
C25 a_2665_112# a_2248_156# 0.63615f
C26 a_1000_472# a_1204_472# 0.66083f
C27 a_1456_156# VSS 0.001901f
C28 a_36_151# a_1204_472# 0.006996f
C29 a_36_151# D 0.094113f
C30 VDD RN 0.035003f
C31 RN a_2560_156# 0.038779f
C32 RN a_1308_423# 0.079294f
C33 a_1288_156# VSS 0.001702f
C34 a_2665_112# Q 0.263315f
C35 a_448_472# VDD 0.456269f
C36 VDD a_2248_156# 1.12036f
C37 a_448_472# a_1308_423# 0.882105f
C38 a_448_472# a_2560_156# 0.277491f
C39 a_1000_472# RN 0.0832f
C40 a_2248_156# a_2560_156# 0.119687f
C41 a_2248_156# a_1308_423# 0.056721f
C42 a_36_151# RN 0.080119f
C43 a_1000_472# a_796_472# 0.048436f
C44 a_796_472# a_36_151# 0.011851f
C45 a_448_472# a_1000_472# 0.361958f
C46 a_448_472# a_36_151# 0.536965f
C47 a_1000_472# a_2248_156# 0.001232f
C48 a_36_151# a_2248_156# 0.042802f
C49 VDD Q 0.260055f
C50 a_448_472# a_1456_156# 0.00227f
C51 a_448_472# a_1288_156# 0.002067f
C52 VNW VSS 0.012596f
C53 VDD CLK 0.02303f
C54 VNW a_1204_472# 0.016269f
C55 a_2665_112# VDD 0.152571f
C56 VNW D 0.128231f
C57 a_2665_112# a_2560_156# 0.116229f
C58 a_36_151# CLK 0.669598f
C59 a_2665_112# a_36_151# 0.019033f
C60 VNW RN 0.304626f
C61 VDD a_1308_423# 0.094185f
C62 VNW a_796_472# 0.010232f
C63 VDD a_2560_156# 0.00302f
C64 D VSS 0.064618f
C65 VNW a_448_472# 0.341284f
C66 VNW a_2248_156# 0.181292f
C67 a_3041_156# VSS 0.004935f
C68 VDD a_1000_472# 0.119211f
C69 VDD a_36_151# 0.417101f
C70 a_1000_472# a_1308_423# 0.934191f
C71 a_36_151# a_2560_156# 0.003674f
C72 a_36_151# a_1308_423# 0.05539f
C73 RN VSS 0.436942f
C74 VNW Q 0.026596f
C75 a_796_472# VSS 0.05215f
C76 a_1000_472# a_36_151# 0.08126f
C77 RN a_1204_472# 0.021039f
C78 a_448_472# VSS 1.20207f
C79 a_2248_156# VSS 0.030372f
C80 a_448_472# a_1204_472# 0.008996f
C81 a_796_472# D 0.082858f
C82 a_3041_156# RN 0.014924f
C83 a_448_472# D 0.328788f
C84 VNW CLK 0.137037f
C85 VSS Q 0.170514f
C86 Q VSUBS 0.061347f
C87 VSS VSUBS 1.33519f
C88 RN VSUBS 1.37098f
C89 D VSUBS 0.253406f
C90 VDD VSUBS 0.859994f
C91 CLK VSUBS 0.291241f
C92 VNW VSUBS 6.48579f
C93 a_2560_156# VSUBS 0.016968f
C94 a_2665_112# VSUBS 0.91969f
C95 a_2248_156# VSUBS 0.30886f
C96 a_1204_472# VSUBS 0.012971f
C97 a_1000_472# VSUBS 0.291735f
C98 a_796_472# VSUBS 0.023206f
C99 a_1308_423# VSUBS 0.279043f
C100 a_448_472# VSUBS 0.684413f
C101 a_36_151# VSUBS 1.43587f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VPW VNW a_438_68#
+ a_244_68# a_1254_68# a_1060_68# a_632_68# a_1458_68# VSUBS
X0 a_1458_68# A3 a_1254_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
C0 a_1060_68# VSS 0.001868f
C1 A4 VNW 0.388525f
C2 VDD VSS 0.004026f
C3 a_1254_68# ZN 0.008913f
C4 A1 ZN 0.071728f
C5 A4 VSS 0.056757f
C6 A1 VDD 0.044019f
C7 A3 ZN 0.881941f
C8 a_438_68# VSS 0.00542f
C9 A3 a_1060_68# 0.004303f
C10 A4 A1 0.451294f
C11 A3 VDD 0.040467f
C12 a_1458_68# VSS 0.002548f
C13 a_244_68# VSS 0.007139f
C14 A4 A3 0.297972f
C15 a_1060_68# ZN 0.007219f
C16 VDD ZN 1.39778f
C17 A3 a_438_68# 0.007312f
C18 A2 VNW 0.317841f
C19 A4 ZN 1.94271f
C20 a_632_68# VSS 0.005832f
C21 A2 VSS 0.036637f
C22 A3 a_244_68# 0.007f
C23 A4 VDD 0.047422f
C24 VNW VSS 0.006403f
C25 a_1458_68# ZN 0.01082f
C26 A1 A2 0.516286f
C27 A3 a_632_68# 0.0083f
C28 A1 VNW 0.345207f
C29 A3 A2 0.40854f
C30 a_1254_68# VSS 0.002331f
C31 A1 VSS 0.037456f
C32 A3 VNW 0.300046f
C33 a_632_68# ZN 0.001673f
C34 A2 ZN 0.068627f
C35 A3 VSS 0.248503f
C36 VNW ZN 0.062752f
C37 A2 VDD 0.041932f
C38 A3 a_1254_68# 0.004873f
C39 A3 A1 0.831807f
C40 VDD VNW 0.1769f
C41 ZN VSS 0.89636f
C42 A4 A2 0.762551f
C43 VSS VSUBS 0.597574f
C44 VDD VSUBS 0.397078f
C45 ZN VSUBS 0.12583f
C46 A1 VSUBS 0.558392f
C47 A2 VSUBS 0.513744f
C48 A3 VSUBS 0.547819f
C49 A4 VSUBS 0.580825f
C50 VNW VSUBS 3.05206f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
C0 I VSS 0.071429f
C1 I VNW 0.283715f
C2 ZN VDD 0.24022f
C3 ZN VSS 0.15979f
C4 VDD VSS 0.022662f
C5 VNW ZN 0.025997f
C6 VNW VDD 0.103267f
C7 I ZN 0.614595f
C8 VNW VSS 0.01054f
C9 I VDD 0.164681f
C10 VSS VSUBS 0.345063f
C11 ZN VSUBS 0.094435f
C12 VDD VSUBS 0.235951f
C13 I VSUBS 0.642286f
C14 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VPW VNW a_468_472#
+ a_224_472# a_244_68# a_916_472# VSUBS
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
C0 A3 A2 0.129823f
C1 VDD VSS 0.027141f
C2 A3 VNW 0.13805f
C3 B2 a_244_68# 0.29062f
C4 a_468_472# A2 0.002382f
C5 ZN B1 0.457921f
C6 A1 VSS 0.029231f
C7 B1 VNW 0.116377f
C8 VDD A1 0.015114f
C9 a_244_68# VSS 0.329999f
C10 A3 a_224_472# 0.012212f
C11 B2 ZN 0.371232f
C12 VDD a_244_68# 0.520053f
C13 B2 VNW 0.125762f
C14 a_244_68# A1 0.480797f
C15 VDD a_916_472# 0.004169f
C16 VSS A2 0.030842f
C17 ZN VSS 0.069913f
C18 VSS VNW 0.013582f
C19 VDD A2 0.071137f
C20 ZN VDD 0.006472f
C21 VDD VNW 0.158216f
C22 a_244_68# a_916_472# 0.018012f
C23 A1 A2 0.038953f
C24 ZN A1 0.164807f
C25 A1 VNW 0.125824f
C26 a_224_472# VSS 0.00124f
C27 a_244_68# A2 0.356992f
C28 ZN a_244_68# 0.2576f
C29 B2 B1 0.038725f
C30 a_244_68# VNW 0.043485f
C31 a_224_472# VDD 0.016257f
C32 ZN a_916_472# 0.008827f
C33 A3 VSS 0.046517f
C34 B1 VSS 0.072063f
C35 A3 VDD 0.236688f
C36 a_224_472# a_244_68# 0.004752f
C37 A2 VNW 0.121626f
C38 ZN VNW 0.012941f
C39 a_468_472# VDD 0.005594f
C40 B1 VDD 0.015317f
C41 a_468_472# A1 0.001494f
C42 B1 A1 0.13457f
C43 B2 VSS 0.072128f
C44 A3 a_244_68# 0.010697f
C45 a_468_472# a_244_68# 0.022611f
C46 B1 a_244_68# 0.212448f
C47 a_224_472# A2 0.014544f
C48 B2 VDD 0.018546f
C49 VSS VSUBS 0.474343f
C50 ZN VSUBS 0.00986f
C51 VDD VSUBS 0.363224f
C52 B2 VSUBS 0.282623f
C53 B1 VSUBS 0.257203f
C54 A1 VSUBS 0.255736f
C55 A2 VSUBS 0.254473f
C56 A3 VSUBS 0.308666f
C57 VNW VSUBS 2.35586f
C58 a_244_68# VSUBS 0.138666f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VPW VNW a_244_567# a_718_527#
+ a_2172_497# a_56_567# a_1948_68# a_728_93# a_1296_93# VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
C0 a_56_567# a_718_527# 0.00772f
C1 ZN VDD 0.47211f
C2 VDD a_244_567# 0.006111f
C3 ZN a_1296_93# 0.029802f
C4 ZN a_728_93# 0.663929f
C5 ZN VNW 0.032895f
C6 ZN A3 0.033406f
C7 VDD A2 0.210416f
C8 a_1296_93# A2 0.002759f
C9 ZN a_1948_68# 0.381585f
C10 ZN VSS 0.004739f
C11 a_952_93# a_728_93# 0.003723f
C12 a_952_93# VSS 0.003841f
C13 VDD a_1296_93# 0.030892f
C14 a_244_567# a_56_567# 0.00105f
C15 a_728_93# A2 0.516752f
C16 VNW A2 0.388997f
C17 ZN a_2172_497# 0.03345f
C18 A1 A2 0.757944f
C19 VSS A2 0.051212f
C20 A2 a_718_527# 0.141128f
C21 a_728_93# VDD 0.78216f
C22 a_728_93# a_1296_93# 0.624643f
C23 VNW VDD 0.370487f
C24 VNW a_1296_93# 0.155715f
C25 VDD A3 0.022483f
C26 A3 a_1296_93# 0.356198f
C27 VDD A1 0.022573f
C28 a_1948_68# VDD 0.001604f
C29 a_56_567# A2 0.174541f
C30 VSS VDD 0.011823f
C31 a_1948_68# a_1296_93# 0.005923f
C32 VSS a_1296_93# 0.379749f
C33 VDD a_718_527# 0.618394f
C34 a_1296_93# a_1504_93# 0.003723f
C35 a_728_93# VNW 0.385878f
C36 a_728_93# A3 0.721889f
C37 VDD a_56_567# 0.056918f
C38 VNW A3 0.298581f
C39 a_728_93# A1 0.281966f
C40 a_728_93# a_1948_68# 0.02618f
C41 a_728_93# VSS 0.328386f
C42 VNW A1 0.342048f
C43 VNW a_1948_68# 0.002346f
C44 VNW VSS 0.009921f
C45 a_1948_68# A3 0.069927f
C46 VSS A3 0.047056f
C47 VDD a_2172_497# 0.010751f
C48 a_728_93# a_718_527# 0.21558f
C49 VSS A1 0.0538f
C50 VSS a_1948_68# 0.719859f
C51 VNW a_718_527# 0.020227f
C52 A1 a_718_527# 0.023145f
C53 a_728_93# a_56_567# 0.070648f
C54 a_244_567# A2 0.004089f
C55 VNW a_56_567# 0.187311f
C56 VSS a_1504_93# 0.003902f
C57 a_56_567# A1 0.368741f
C58 VSS a_56_567# 0.400197f
C59 a_728_93# a_2172_497# 0.010602f
C60 VSS VSUBS 0.875791f
C61 ZN VSUBS 0.08517f
C62 A1 VSUBS 0.604039f
C63 A2 VSUBS 0.633287f
C64 VDD VSUBS 0.584594f
C65 A3 VSUBS 0.573218f
C66 VNW VSUBS 4.42794f
C67 a_1948_68# VSUBS 0.022025f
C68 a_718_527# VSUBS 0.001795f
C69 a_56_567# VSUBS 0.424713f
C70 a_728_93# VSUBS 0.65929f
C71 a_1296_93# VSUBS 0.317801f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VPW VNW a_36_68# a_244_497#
+ a_1657_68# a_1229_68# a_716_497# VSUBS
X0 a_1229_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
C0 ZN C 0.501479f
C1 ZN VDD 0.761655f
C2 A2 a_36_68# 0.091399f
C3 B ZN 0.3603f
C4 C a_36_68# 0.055076f
C5 ZN A1 0.622246f
C6 ZN a_716_497# 0.025301f
C7 VDD a_36_68# 0.019083f
C8 A2 VNW 0.30827f
C9 ZN VSS 0.004788f
C10 B a_36_68# 0.587375f
C11 a_1229_68# a_36_68# 0.011792f
C12 VNW C 0.309331f
C13 A1 a_36_68# 0.039393f
C14 a_1657_68# a_36_68# 0.009002f
C15 VNW VDD 0.219901f
C16 VSS a_36_68# 2.1107f
C17 ZN a_244_497# 0.006285f
C18 B VNW 0.311256f
C19 VNW A1 0.269127f
C20 A2 VDD 0.147417f
C21 VNW VSS 0.005994f
C22 B A2 0.037237f
C23 C VDD 0.056662f
C24 A2 A1 0.722847f
C25 A2 a_716_497# 0.010693f
C26 A2 VSS 0.030494f
C27 B C 0.698524f
C28 B VDD 0.089771f
C29 VDD A1 0.033883f
C30 C VSS 0.04168f
C31 B a_1229_68# 0.003462f
C32 VDD a_716_497# 0.008883f
C33 VDD VSS 0.007619f
C34 B a_1657_68# 0.002626f
C35 A2 a_244_497# 0.020646f
C36 B VSS 0.032629f
C37 VSS a_1229_68# 0.002856f
C38 A1 VSS 0.031008f
C39 VSS a_1657_68# 0.002208f
C40 VDD a_244_497# 0.016799f
C41 ZN a_36_68# 0.528658f
C42 ZN VNW 0.042076f
C43 ZN A2 1.02528f
C44 VNW a_36_68# 0.00468f
C45 VSS VSUBS 0.620026f
C46 ZN VSUBS 0.062404f
C47 VDD VSUBS 0.531064f
C48 C VSUBS 0.529789f
C49 B VSUBS 0.589191f
C50 A1 VSUBS 0.58772f
C51 A2 VSUBS 0.613706f
C52 VNW VSUBS 3.34705f
C53 a_36_68# VSUBS 0.052951f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VPW VNW a_428_148# a_36_148#
+ VSUBS
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VSUBS nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VSUBS nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VSUBS nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VSUBS nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
C0 VDD VSS 0.012823f
C1 VDD Z 0.164783f
C2 a_36_148# VNW 0.194548f
C3 A2 VSS 0.004456f
C4 VNW A1 0.214361f
C5 VNW VDD 0.134134f
C6 VSS A3 0.005273f
C7 VNW A2 0.189332f
C8 A3 Z 0.001054f
C9 VNW A3 0.213241f
C10 VSS Z 0.093779f
C11 a_36_148# a_244_148# 0.004781f
C12 a_36_148# a_428_148# 0.007047f
C13 a_244_148# A1 0.002081f
C14 VNW VSS 0.007319f
C15 VNW Z 0.033257f
C16 a_36_148# A1 0.205722f
C17 a_36_148# VDD 0.556761f
C18 VDD A1 0.021719f
C19 a_36_148# A2 0.141951f
C20 A2 A1 0.307806f
C21 a_428_148# A3 0.001335f
C22 A2 VDD 0.022493f
C23 a_36_148# A3 0.477475f
C24 VDD A3 0.022574f
C25 a_36_148# VSS 0.798993f
C26 a_36_148# Z 0.156534f
C27 A2 A3 0.340591f
C28 VSS A1 0.00434f
C29 VSS VSUBS 0.415001f
C30 Z VSUBS 0.095371f
C31 VDD VSUBS 0.277732f
C32 A3 VSUBS 0.275015f
C33 A2 VSUBS 0.257076f
C34 A1 VSUBS 0.330738f
C35 VNW VSUBS 2.00777f
C36 a_36_148# VSUBS 0.388358f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VPW VNW a_1044_68# a_452_68#
+ a_276_68# a_860_68# VSUBS
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VSUBS nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 ZN VDD 0.550625f
C1 ZN VNW 0.034063f
C2 A3 ZN 1.24554f
C3 A1 ZN 0.430404f
C4 VSS a_452_68# 0.003244f
C5 VSS A2 0.130985f
C6 VSS a_276_68# 0.003438f
C7 VDD VNW 0.172362f
C8 VSS a_1044_68# 0.00861f
C9 VSS a_860_68# 0.005864f
C10 A3 VDD 0.099291f
C11 A3 VNW 0.347673f
C12 A1 VDD 0.041745f
C13 A2 a_1044_68# 0.006328f
C14 A1 VNW 0.280755f
C15 a_860_68# A2 0.003842f
C16 VSS ZN 0.476547f
C17 A3 A1 0.037905f
C18 ZN a_452_68# 0.007752f
C19 ZN A2 0.082264f
C20 ZN a_276_68# 0.007178f
C21 ZN a_1044_68# 0.001223f
C22 a_860_68# ZN 0.001808f
C23 VSS VDD 0.009236f
C24 VSS VNW 0.007349f
C25 A2 VDD 0.041181f
C26 A2 VNW 0.279783f
C27 A3 VSS 0.074424f
C28 A1 VSS 0.050488f
C29 A3 A2 1.13496f
C30 A1 a_452_68# 0.001247f
C31 A1 A2 0.708241f
C32 VSS VSUBS 0.511432f
C33 ZN VSUBS 0.112753f
C34 VDD VSUBS 0.407724f
C35 A1 VSUBS 0.540441f
C36 A2 VSUBS 0.524145f
C37 A3 VSUBS 0.582222f
C38 VNW VSUBS 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VPW VNW a_692_473#
+ a_254_473# a_66_473# a_2700_473# a_1660_473# a_3220_473# a_1212_473# a_2180_473#
+ a_3740_473# a_1920_473# VSUBS
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
C0 A1 VSS 0.093176f
C1 ZN a_2180_473# 0.018904f
C2 VDD a_1920_473# 0.004058f
C3 a_66_473# A2 0.182327f
C4 a_1660_473# ZN 0.00216f
C5 VNW ZN 0.038639f
C6 A3 VSS 0.078892f
C7 A1 a_66_473# 0.077909f
C8 a_254_473# a_66_473# 0.016207f
C9 VDD A4 0.110338f
C10 A3 a_66_473# 1.66251f
C11 ZN a_3220_473# 0.019778f
C12 a_2700_473# ZN 0.019492f
C13 a_1920_473# a_66_473# 0.023791f
C14 VSS A4 0.099821f
C15 VSS VDD 0.009708f
C16 a_66_473# A4 0.100571f
C17 VDD a_66_473# 3.19476f
C18 ZN A2 2.14591f
C19 A1 ZN 1.60655f
C20 VSS a_66_473# 0.01197f
C21 VDD a_1212_473# 0.014305f
C22 A3 ZN 0.417545f
C23 a_3740_473# A2 0.010293f
C24 a_1920_473# ZN 0.017667f
C25 VNW A2 0.584134f
C26 A1 VNW 0.553741f
C27 a_1660_473# A3 0.0054f
C28 A3 VNW 0.567739f
C29 ZN A4 1.44735f
C30 a_66_473# a_1212_473# 0.018664f
C31 VDD ZN 0.007051f
C32 VDD a_3740_473# 0.003118f
C33 VDD a_2180_473# 0.00368f
C34 VNW A4 0.513548f
C35 VSS ZN 4.39577f
C36 a_1660_473# VDD 0.008572f
C37 VDD VNW 0.394018f
C38 ZN a_66_473# 0.956309f
C39 a_692_473# VDD 0.017923f
C40 a_3740_473# a_66_473# 0.028219f
C41 VDD a_3220_473# 0.003326f
C42 A1 A2 2.13585f
C43 a_2700_473# VDD 0.003457f
C44 VSS VNW 0.006947f
C45 a_66_473# a_2180_473# 0.020817f
C46 A3 A2 0.0303f
C47 a_1660_473# a_66_473# 0.035002f
C48 VNW a_66_473# 0.040351f
C49 a_692_473# a_66_473# 0.022803f
C50 a_66_473# a_3220_473# 0.021354f
C51 a_2700_473# a_66_473# 0.021497f
C52 VDD A2 0.054912f
C53 A1 VDD 0.055928f
C54 A3 A4 1.96796f
C55 VDD a_254_473# 0.012952f
C56 A3 VDD 0.086829f
C57 a_3740_473# ZN 0.004594f
C58 VSS A2 0.076134f
C59 VSS VSUBS 1.3434f
C60 ZN VSUBS 0.240026f
C61 VDD VSUBS 0.844436f
C62 A1 VSUBS 1.40024f
C63 A2 VSUBS 1.30271f
C64 A4 VSUBS 1.33565f
C65 A3 VSUBS 1.29175f
C66 VNW VSUBS 6.70706f
C67 a_66_473# VSUBS 0.11665f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VPW VNW a_49_472# a_1133_69#
+ a_741_69# VSUBS
X0 VSS A2 a_1133_69# VSUBS nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VSUBS nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VSUBS nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
C0 VDD A2 0.029358f
C1 a_1133_69# A1 0.003427f
C2 a_49_472# VSS 0.01207f
C3 A1 a_49_472# 0.03417f
C4 ZN VSS 0.784804f
C5 A2 a_49_472# 0.086717f
C6 A1 ZN 0.182845f
C7 A1 VSS 0.129775f
C8 ZN A2 0.800412f
C9 A2 VSS 0.047574f
C10 VDD B 0.045174f
C11 VDD VNW 0.151549f
C12 A1 A2 0.809974f
C13 a_49_472# B 0.234399f
C14 VNW a_49_472# 0.012852f
C15 ZN B 0.20884f
C16 ZN VNW 0.025755f
C17 B VSS 0.061328f
C18 VNW VSS 0.0086f
C19 A1 VNW 0.241301f
C20 A2 B 0.029994f
C21 A2 VNW 0.272677f
C22 ZN a_741_69# 0.006341f
C23 a_741_69# VSS 0.002035f
C24 VDD a_49_472# 1.09818f
C25 a_741_69# A2 0.001142f
C26 VDD ZN 0.008463f
C27 VDD VSS 0.009099f
C28 a_1133_69# ZN 0.001193f
C29 VDD A1 0.028601f
C30 a_1133_69# VSS 0.00441f
C31 VNW B 0.260678f
C32 ZN a_49_472# 0.475008f
C33 VSS VSUBS 0.510011f
C34 ZN VSUBS 0.070911f
C35 VDD VSUBS 0.327438f
C36 A1 VSUBS 0.556927f
C37 A2 VSUBS 0.56333f
C38 B VSUBS 0.662515f
C39 VNW VSUBS 2.52991f
C40 a_49_472# VSUBS 0.098072f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VPW VNW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 VSS VNW 0.010163f
C1 VNW I 0.285482f
C2 VSS I 0.091531f
C3 VNW ZN 0.027829f
C4 VSS ZN 0.179304f
C5 ZN I 0.58604f
C6 VNW VDD 0.097124f
C7 VSS VDD 0.023187f
C8 I VDD 0.074838f
C9 ZN VDD 0.266247f
C10 VSS VSUBS 0.308828f
C11 ZN VSUBS 0.100523f
C12 VDD VSUBS 0.240805f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VPW VNW a_448_472#
+ a_36_151# a_1293_527# a_3081_151# a_1284_156# a_1040_527# a_1353_112# a_836_156#
+ a_1697_156# a_2449_156# a_3129_107# a_2225_156# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VSUBS nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VSUBS nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VSUBS nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VSUBS nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VSUBS nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VSUBS nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
C0 D VNW 0.1615f
C1 a_36_151# VSS 0.286331f
C2 VSS a_1284_156# 0.003637f
C3 a_836_156# VSS 0.050008f
C4 D VDD 0.004944f
C5 Q a_3129_107# 0.179468f
C6 VSS a_448_472# 1.07431f
C7 VNW CLK 0.136589f
C8 a_836_156# a_36_151# 0.015697f
C9 VDD CLK 0.022091f
C10 a_36_151# a_448_472# 0.473132f
C11 a_1284_156# a_448_472# 0.002691f
C12 a_836_156# a_448_472# 0.427756f
C13 a_1040_527# VSS 0.060221f
C14 SETN VSS 0.008083f
C15 a_2449_156# a_3129_107# 0.00955f
C16 VNW VSS 0.009462f
C17 a_36_151# a_1040_527# 0.206392f
C18 a_836_156# a_1040_527# 0.068207f
C19 VSS VDD 0.013814f
C20 a_36_151# SETN 0.077775f
C21 a_36_151# VNW 0.909435f
C22 a_1040_527# a_448_472# 0.869605f
C23 a_836_156# VNW 0.01368f
C24 SETN a_448_472# 0.083903f
C25 a_36_151# VDD 1.41468f
C26 VNW a_448_472# 0.400964f
C27 VDD a_448_472# 0.624585f
C28 VSS a_2225_156# 1.18908f
C29 a_1040_527# SETN 0.063241f
C30 a_1040_527# VNW 0.223863f
C31 VNW SETN 0.811046f
C32 a_36_151# a_2225_156# 0.153684f
C33 a_1040_527# VDD 0.039677f
C34 SETN VDD 0.127822f
C35 a_2225_156# a_448_472# 0.153996f
C36 VNW VDD 0.539099f
C37 a_2449_156# a_3081_151# 0.001203f
C38 a_1697_156# a_448_472# 0.007618f
C39 SETN a_2225_156# 0.070597f
C40 VSS a_3129_107# 0.136769f
C41 a_36_151# a_1293_527# 0.008379f
C42 VNW a_2225_156# 0.209033f
C43 a_2225_156# VDD 0.073415f
C44 a_1040_527# a_1293_527# 0.00215f
C45 Q VSS 0.131272f
C46 SETN a_3129_107# 0.089288f
C47 VSS a_1353_112# 0.027348f
C48 VNW a_3129_107# 0.323464f
C49 a_3129_107# VDD 0.351307f
C50 a_36_151# a_1353_112# 0.840879f
C51 a_448_472# a_1353_112# 0.317251f
C52 a_36_151# a_2449_156# 0.005967f
C53 a_2225_156# a_3129_107# 0.514036f
C54 Q VNW 0.031621f
C55 a_1040_527# a_1353_112# 0.387423f
C56 a_2449_156# a_448_472# 0.056679f
C57 SETN a_1353_112# 0.072983f
C58 Q VDD 0.282179f
C59 VNW a_1353_112# 0.219511f
C60 D VSS 0.067877f
C61 VDD a_1353_112# 0.016257f
C62 a_2449_156# SETN 0.302222f
C63 a_2449_156# VNW 0.043816f
C64 a_36_151# D 0.092705f
C65 a_836_156# D 0.108102f
C66 VSS CLK 0.021941f
C67 a_2449_156# VDD 0.208631f
C68 D a_448_472# 0.400104f
C69 a_2225_156# a_1353_112# 0.152869f
C70 a_36_151# CLK 0.700974f
C71 a_3081_151# a_2225_156# 0.004129f
C72 a_1697_156# a_1353_112# 0.002752f
C73 CLK a_448_472# 0.001313f
C74 a_2449_156# a_2225_156# 0.569174f
C75 Q VSUBS 0.105566f
C76 VSS VSUBS 1.35707f
C77 SETN VSUBS 0.710246f
C78 D VSUBS 0.247102f
C79 VDD VSUBS 0.833181f
C80 CLK VSUBS 0.290467f
C81 VNW VSUBS 6.44257f
C82 a_2449_156# VSUBS 0.049992f
C83 a_2225_156# VSUBS 0.434082f
C84 a_3129_107# VSUBS 0.58406f
C85 a_836_156# VSUBS 0.019766f
C86 a_1040_527# VSUBS 0.302082f
C87 a_1353_112# VSUBS 0.286513f
C88 a_448_472# VSUBS 1.21246f
C89 a_36_151# VSUBS 1.31409f
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[3] ctln[4] ctln[5] ctln[6] ctln[8] ctlp[0] ctlp[1]
+ ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8] ctlp[9] clk clkc comp en
+ result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7]
+ result[8] result[9] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0]
+ trimb[1] trimb[2] trimb[3] trimb[4] valid net10 output13/a_224_472# output23/a_224_472#
+ net59 net16 net27 output25/a_224_472# cal_itt\[1\] fanout65/a_36_113# ctln[2] ctln[7]
+ net15 ctln[9] output10/a_224_472# net26 net24 output11/a_224_472# output21/a_224_472#
+ net14 output12/a_224_472# output22/a_224_472# cal net62 net20 vss vdd
XFILLER_0_17_200 vdd vss FILLER_0_17_200/VPW vdd FILLER_0_17_200/a_36_472# FILLER_0_17_200/a_572_375#
+ FILLER_0_17_200/a_124_375# FILLER_0_17_200/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd ANTENNA_fanout56_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_294_ vdd vss _008_ _104_ _106_ _294_/VPW vdd _294_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_432_ _021_ mask\[3\] net63 vss net80 vdd _432_/VPW vdd _432_/a_2665_112# _432_/a_448_472#
+ _432_/a_796_472# _432_/a_36_151# _432_/a_1204_472# _432_/a_3041_156# _432_/a_1000_472#
+ _432_/a_1308_423# _432_/a_1456_156# _432_/a_1288_156# _432_/a_2248_156# _432_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ _363_/VPW vdd _363_/a_36_68# _363_/a_244_472#
+ _363_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ _346_/VPW vdd _346_/a_49_472#
+ _346_/a_665_69# _346_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd _415_/VPW vdd _415_/a_2665_112# _415_/a_448_472#
+ _415_/a_796_472# _415_/a_36_151# _415_/a_1204_472# _415_/a_3041_156# _415_/a_1000_472#
+ _415_/a_1308_423# _415_/a_1456_156# _415_/a_1288_156# _415_/a_2248_156# _415_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd _277_/VPW vdd _277_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 _200_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd _329_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss FILLER_0_19_125/VPW vdd FILLER_0_19_125/a_36_472# FILLER_0_19_125/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd ANTENNA__392__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss FILLER_0_15_150/VPW vdd FILLER_0_15_150/a_36_472# FILLER_0_15_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss FILLER_0_21_142/VPW vdd FILLER_0_21_142/a_36_472# FILLER_0_21_142/a_572_375#
+ FILLER_0_21_142/a_124_375# FILLER_0_21_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss FILLER_0_16_73/VPW vdd FILLER_0_16_73/a_36_472# FILLER_0_16_73/a_572_375#
+ FILLER_0_16_73/a_124_375# FILLER_0_16_73/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss output20/VPW vdd output20/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss output31/VPW vdd output31/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss output42/VPW vdd output42/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 ctln[0] net7 vdd vss output7/VPW vdd output7/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss FILLER_0_5_117/VPW vdd FILLER_0_5_117/a_36_472# FILLER_0_5_117/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss FILLER_0_5_128/VPW vdd FILLER_0_5_128/a_36_472# FILLER_0_5_128/a_572_375#
+ FILLER_0_5_128/a_124_375# FILLER_0_5_128/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_293_ net31 vdd vss _106_ mask\[4\] _105_ _293_/VPW vdd _293_/a_36_472# _293_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_431_ _020_ mask\[2\] net53 vss net70 vdd _431_/VPW vdd _431_/a_2665_112# _431_/a_448_472#
+ _431_/a_796_472# _431_/a_36_151# _431_/a_1204_472# _431_/a_3041_156# _431_/a_1000_472#
+ _431_/a_1308_423# _431_/a_1456_156# _431_/a_1288_156# _431_/a_2248_156# _431_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_362_ vdd vss trim_mask\[1\] _155_ _362_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_345_ vss _144_ _132_ vdd _345_/VPW vdd _345_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ vss _093_ _092_ vdd _276_/VPW vdd _276_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd _414_/VPW vdd _414_/a_2665_112# _414_/a_448_472#
+ _414_/a_796_472# _414_/a_36_151# _414_/a_1204_472# _414_/a_3041_156# _414_/a_1000_472#
+ _414_/a_1308_423# _414_/a_1456_156# _414_/a_1288_156# _414_/a_2248_156# _414_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd _328_/VPW vdd _328_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss FILLER_0_9_28/VPW vdd FILLER_0_9_28/a_1916_375# FILLER_0_9_28/a_1380_472#
+ FILLER_0_9_28/a_3260_375# FILLER_0_9_28/a_36_472# FILLER_0_9_28/a_932_472# FILLER_0_9_28/a_2812_375#
+ FILLER_0_9_28/a_2276_472# FILLER_0_9_28/a_1828_472# FILLER_0_9_28/a_3172_472# FILLER_0_9_28/a_572_375#
+ FILLER_0_9_28/a_2724_472# FILLER_0_9_28/a_124_375# FILLER_0_9_28/a_1468_375# FILLER_0_9_28/a_1020_375#
+ FILLER_0_9_28/a_484_472# FILLER_0_9_28/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_204 vdd vss FILLER_0_3_204/VPW vdd FILLER_0_3_204/a_36_472# FILLER_0_3_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _078_ vdd vss _080_ _073_ _076_ _259_/VPW vdd _259_/a_455_68# _259_/a_271_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd vss FILLER_0_16_107/VPW vdd FILLER_0_16_107/a_36_472# FILLER_0_16_107/a_572_375#
+ FILLER_0_16_107/a_124_375# FILLER_0_16_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd ANTENNA_fanout79_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd ANTENNA__358__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss output21/VPW vdd output21/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss output43/VPW vdd output43/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss output32/VPW vdd output32/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss output10/VPW vdd output10/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss output8/VPW vdd output8/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd ANTENNA_input3_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ vss _105_ _098_ vdd _292_/VPW vdd _292_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_430_ _019_ mask\[1\] net63 vss net80 vdd _430_/VPW vdd _430_/a_2665_112# _430_/a_448_472#
+ _430_/a_796_472# _430_/a_36_151# _430_/a_1204_472# _430_/a_3041_156# _430_/a_1000_472#
+ _430_/a_1308_423# _430_/a_1456_156# _430_/a_1288_156# _430_/a_2248_156# _430_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_361_ vdd vss _154_ _086_ _119_ _361_/VPW vdd _361_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss FILLER_0_7_72/VPW vdd FILLER_0_7_72/a_1916_375# FILLER_0_7_72/a_1380_472#
+ FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472# FILLER_0_7_72/a_932_472# FILLER_0_7_72/a_2812_375#
+ FILLER_0_7_72/a_2276_472# FILLER_0_7_72/a_1828_472# FILLER_0_7_72/a_3172_472# FILLER_0_7_72/a_572_375#
+ FILLER_0_7_72/a_2724_472# FILLER_0_7_72/a_124_375# FILLER_0_7_72/a_1468_375# FILLER_0_7_72/a_1020_375#
+ FILLER_0_7_72/a_484_472# FILLER_0_7_72/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ _344_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ _275_/VPW vdd _275_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__191__I vss net17 vdd ANTENNA__191__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd _413_/VPW vdd _413_/a_2665_112# _413_/a_448_472#
+ _413_/a_796_472# _413_/a_36_151# _413_/a_1204_472# _413_/a_3041_156# _413_/a_1000_472#
+ _413_/a_1308_423# _413_/a_1456_156# _413_/a_1288_156# _413_/a_2248_156# _413_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_96 vdd vss FILLER_0_24_96/VPW vdd FILLER_0_24_96/a_36_472# FILLER_0_24_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss FILLER_0_24_63/VPW vdd FILLER_0_24_63/a_36_472# FILLER_0_24_63/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ vdd vss _043_ net27 mask\[0\] _189_/VPW vdd _189_/a_255_603# _189_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_327_ _131_ vdd vss _016_ _127_ _130_ _327_/VPW vdd _327_/a_36_472# _327_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ vss _079_ _078_ vdd _258_/VPW vdd _258_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss FILLER_0_18_171/VPW vdd FILLER_0_18_171/a_36_472# FILLER_0_18_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss FILLER_0_24_130/VPW vdd FILLER_0_24_130/a_36_472# FILLER_0_24_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd ANTENNA__377__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss FILLER_0_21_133/VPW vdd FILLER_0_21_133/a_36_472# FILLER_0_21_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss FILLER_0_8_138/VPW vdd FILLER_0_8_138/a_36_472# FILLER_0_8_138/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss FILLER_0_8_127/VPW vdd FILLER_0_8_127/a_36_472# FILLER_0_8_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 ctlp[5] net22 vdd vss output22/VPW vdd output22/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 result[6] net33 vdd vss output33/VPW vdd output33/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss output44/VPW vdd output44/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss output11/VPW vdd output11/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss output9/VPW vdd output9/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd ANTENNA__194__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd _291_/VPW vdd _291_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss FILLER_0_4_152/VPW vdd FILLER_0_4_152/a_36_472# FILLER_0_4_152/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss FILLER_0_4_185/VPW vdd FILLER_0_4_185/a_36_472# FILLER_0_4_185/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd _360_/VPW vdd _360_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss FILLER_0_13_65/VPW vdd FILLER_0_13_65/a_36_472# FILLER_0_13_65/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ _343_/VPW vdd _343_/a_49_472#
+ _343_/a_665_69# _343_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ _274_/VPW vdd _274_/a_36_68# _274_/a_1612_497#
+ _274_/a_2124_68# _274_/a_244_497# _274_/a_2960_68# _274_/a_3368_68# _274_/a_2552_68#
+ _274_/a_1164_497# _274_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd _412_/VPW vdd _412_/a_2665_112# _412_/a_448_472#
+ _412_/a_796_472# _412_/a_36_151# _412_/a_1204_472# _412_/a_3041_156# _412_/a_1000_472#
+ _412_/a_1308_423# _412_/a_1456_156# _412_/a_1288_156# _412_/a_2248_156# _412_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__292__I vss _098_ vdd ANTENNA__292__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ _326_/VPW vdd _326_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ _257_/VPW vdd _257_/a_36_472# _257_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd _309_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd ANTENNA__197__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__301__A2 vss _098_ vdd ANTENNA__301__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss FILLER_0_15_142/VPW vdd FILLER_0_15_142/a_36_472# FILLER_0_15_142/a_572_375#
+ FILLER_0_15_142/a_124_375# FILLER_0_15_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 ctlp[6] net23 vdd vss output23/VPW vdd output23/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss output45/VPW vdd output45/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss output34/VPW vdd output34/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss output12/VPW vdd output12/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss FILLER_0_5_109/VPW vdd FILLER_0_5_109/a_36_472# FILLER_0_5_109/a_572_375#
+ FILLER_0_5_109/a_124_375# FILLER_0_5_109/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss FILLER_0_17_226/VPW vdd FILLER_0_17_226/a_36_472# FILLER_0_17_226/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss FILLER_0_4_197/VPW vdd FILLER_0_4_197/a_1380_472# FILLER_0_4_197/a_36_472#
+ FILLER_0_4_197/a_932_472# FILLER_0_4_197/a_572_375# FILLER_0_4_197/a_124_375# FILLER_0_4_197/a_1468_375#
+ FILLER_0_4_197/a_1020_375# FILLER_0_4_197/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ _290_/VPW vdd _290_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss FILLER_0_9_223/VPW vdd FILLER_0_9_223/a_36_472# FILLER_0_9_223/a_572_375#
+ FILLER_0_9_223/a_124_375# FILLER_0_9_223/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ _342_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_273_ vss _090_ state\[0\] vdd _273_/VPW vdd _273_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd _411_/VPW vdd _411_/a_2665_112# _411_/a_448_472#
+ _411_/a_796_472# _411_/a_36_151# _411_/a_1204_472# _411_/a_3041_156# _411_/a_1000_472#
+ _411_/a_1308_423# _411_/a_1456_156# _411_/a_1288_156# _411_/a_2248_156# _411_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout80 vss net80 net81 vdd fanout80/VPW vdd fanout80/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_325_ vdd vss _130_ _118_ _129_ _325_/VPW vdd _325_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd vss FILLER_0_10_78/VPW vdd FILLER_0_10_78/a_1380_472# FILLER_0_10_78/a_36_472#
+ FILLER_0_10_78/a_932_472# FILLER_0_10_78/a_572_375# FILLER_0_10_78/a_124_375# FILLER_0_10_78/a_1468_375#
+ FILLER_0_10_78/a_1020_375# FILLER_0_10_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ _256_/VPW vdd _256_/a_36_68# _256_/a_1612_497#
+ _256_/a_2124_68# _256_/a_244_497# _256_/a_2960_68# _256_/a_3368_68# _256_/a_2552_68#
+ _256_/a_1164_497# _256_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ _308_/VPW vdd _308_/a_848_380# _308_/a_1084_68#
+ _308_/a_124_24# _308_/a_1152_472# _308_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss FILLER_0_1_98/VPW vdd FILLER_0_1_98/a_36_472# FILLER_0_1_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ _239_/VPW vdd _239_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss FILLER_0_12_124/VPW vdd FILLER_0_12_124/a_36_472# FILLER_0_12_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss FILLER_0_8_107/VPW vdd FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 ctlp[7] net24 vdd vss output24/VPW vdd output24/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss output35/VPW vdd output35/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss output46/VPW vdd output46/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss FILLER_0_18_2/VPW vdd FILLER_0_18_2/a_1916_375# FILLER_0_18_2/a_1380_472#
+ FILLER_0_18_2/a_3260_375# FILLER_0_18_2/a_36_472# FILLER_0_18_2/a_932_472# FILLER_0_18_2/a_2812_375#
+ FILLER_0_18_2/a_2276_472# FILLER_0_18_2/a_1828_472# FILLER_0_18_2/a_3172_472# FILLER_0_18_2/a_572_375#
+ FILLER_0_18_2/a_2724_472# FILLER_0_18_2/a_124_375# FILLER_0_18_2/a_1468_375# FILLER_0_18_2/a_1020_375#
+ FILLER_0_18_2/a_484_472# FILLER_0_18_2/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 ctln[6] net13 vdd vss output13/VPW vdd output13/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss FILLER_0_7_162/VPW vdd FILLER_0_7_162/a_36_472# FILLER_0_7_162/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss FILLER_0_7_195/VPW vdd FILLER_0_7_195/a_36_472# FILLER_0_7_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd ANTENNA_input1_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd ANTENNA__414__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ _341_/VPW vdd _341_/a_49_472#
+ _341_/a_665_69# _341_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss _410_/VPW vdd _410_/a_36_68# _410_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ _272_/VPW vdd _272_/a_36_472# _272_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd fanout70/VPW vdd fanout70/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ _076_ vss vdd _057_ _255_/VPW vdd _255_/a_224_552# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_324_ vdd vss _129_ calibrate _062_ _324_/VPW vdd _324_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output40_I vss net40 vdd ANTENNA_output40_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 vss net81 net82 vdd fanout81/VPW vdd fanout81/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_55 vdd vss FILLER_0_19_55/VPW vdd FILLER_0_19_55/a_36_472# FILLER_0_19_55/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A1 vss _093_ vdd ANTENNA__304__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_307_ vdd vss _114_ _113_ _096_ _307_/VPW vdd _307_/a_234_472# _307_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] _238_/VPW vdd _238_/a_255_603# _238_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss FILLER_0_21_125/VPW vdd FILLER_0_21_125/a_36_472# FILLER_0_21_125/a_572_375#
+ FILLER_0_21_125/a_124_375# FILLER_0_21_125/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss FILLER_0_16_89/VPW vdd FILLER_0_16_89/a_1380_472# FILLER_0_16_89/a_36_472#
+ FILLER_0_16_89/a_932_472# FILLER_0_16_89/a_572_375# FILLER_0_16_89/a_124_375# FILLER_0_16_89/a_1468_375#
+ FILLER_0_16_89/a_1020_375# FILLER_0_16_89/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss FILLER_0_12_136/VPW vdd FILLER_0_12_136/a_1380_472# FILLER_0_12_136/a_36_472#
+ FILLER_0_12_136/a_932_472# FILLER_0_12_136/a_572_375# FILLER_0_12_136/a_124_375#
+ FILLER_0_12_136/a_1468_375# FILLER_0_12_136/a_1020_375# FILLER_0_12_136/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 ctlp[8] net25 vdd vss output25/VPW vdd output25/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss output47/VPW vdd output47/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 result[9] net36 vdd vss output36/VPW vdd output36/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss output14/VPW vdd output14/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss FILLER_0_4_144/VPW vdd FILLER_0_4_144/a_36_472# FILLER_0_4_144/a_572_375#
+ FILLER_0_4_144/a_124_375# FILLER_0_4_144/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss FILLER_0_4_177/VPW vdd FILLER_0_4_177/a_36_472# FILLER_0_4_177/a_572_375#
+ FILLER_0_4_177/a_124_375# FILLER_0_4_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd _340_/VPW vdd _340_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ _271_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd ANTENNA__356__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss FILLER_0_10_256/VPW vdd FILLER_0_10_256/a_36_472# FILLER_0_10_256/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__200__I vss net20 vdd ANTENNA__200__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd ANTENNA_fanout52_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_99 vdd vss FILLER_0_4_99/VPW vdd FILLER_0_4_99/a_36_472# FILLER_0_4_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss FILLER_0_6_239/VPW vdd FILLER_0_6_239/a_36_472# FILLER_0_6_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout71 vss net71 net73 vdd fanout71/VPW vdd fanout71/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 net60 vss vdd net61 fanout60/VPW vdd fanout60/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_323_ vss _015_ _128_ vdd _323_/VPW vdd _323_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd fanout82/VPW vdd fanout82/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ _254_/VPW vdd _254_/a_448_472# _254_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_237_ vdd vss net40 net45 _237_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_306_ vss _113_ _057_ vdd _306_/VPW vdd _306_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_57 vdd vss FILLER_0_16_57/VPW vdd FILLER_0_16_57/a_1380_472# FILLER_0_16_57/a_36_472#
+ FILLER_0_16_57/a_932_472# FILLER_0_16_57/a_572_375# FILLER_0_16_57/a_124_375# FILLER_0_16_57/a_1468_375#
+ FILLER_0_16_57/a_1020_375# FILLER_0_16_57/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss output26/VPW vdd output26/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss output15/VPW vdd output15/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss output48/VPW vdd output48/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss output37/VPW vdd output37/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss FILLER_0_17_218/VPW vdd FILLER_0_17_218/a_36_472# FILLER_0_17_218/a_572_375#
+ FILLER_0_17_218/a_124_375# FILLER_0_17_218/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss FILLER_0_4_123/VPW vdd FILLER_0_4_123/a_36_472# FILLER_0_4_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd ANTENNA__203__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ _270_/VPW vdd _270_/a_36_472# _270_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ _399_/VPW vdd _399_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ _322_/VPW vdd _322_/a_848_380# _322_/a_1084_68#
+ _322_/a_124_24# _322_/a_1152_472# _322_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd fanout61/VPW vdd fanout61/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd fanout72/VPW vdd fanout72/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd vss FILLER_0_10_37/VPW vdd FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net50 vss vdd net52 fanout50/VPW vdd fanout50/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] _253_/VPW vdd _253_/a_36_68#
+ _253_/a_1732_68# _253_/a_244_68# _253_/a_1100_68# _253_/a_1528_68# _253_/a_672_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_305_ vdd vss _112_ net1 _081_ _305_/VPW vdd _305_/a_36_159# vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ net40 vss vdd _064_ _236_/VPW vdd _236_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vss net22 vdd ANTENNA__206__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss FILLER_0_20_193/VPW vdd FILLER_0_20_193/a_36_472# FILLER_0_20_193/a_572_375#
+ FILLER_0_20_193/a_124_375# FILLER_0_20_193/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd _219_/VPW vdd _219_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss output27/VPW vdd output27/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss output16/VPW vdd output16/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss output38/VPW vdd output38/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss FILLER_0_16_241/VPW vdd FILLER_0_16_241/a_36_472# FILLER_0_16_241/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd _398_/VPW vdd _398_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vss FILLER_0_10_247/VPW vdd FILLER_0_10_247/a_36_472# FILLER_0_10_247/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_214 vdd vss FILLER_0_10_214/VPW vdd FILLER_0_10_214/a_36_472# FILLER_0_10_214/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_91 vdd vss FILLER_0_14_91/VPW vdd FILLER_0_14_91/a_36_472# FILLER_0_14_91/a_572_375#
+ FILLER_0_14_91/a_124_375# FILLER_0_14_91/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__209__I vss net23 vdd ANTENNA__209__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I vss net19 vdd ANTENNA_output19_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss FILLER_0_19_47/VPW vdd FILLER_0_19_47/a_36_472# FILLER_0_19_47/a_572_375#
+ FILLER_0_19_47/a_124_375# FILLER_0_19_47/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd fanout73/VPW vdd fanout73/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 net62 vss vdd net64 fanout62/VPW vdd fanout62/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vss net51 net52 vdd fanout51/VPW vdd fanout51/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ _321_/VPW vdd _321_/a_2590_472# _321_/a_170_472#
+ _321_/a_1602_69# _321_/a_786_69# _321_/a_3126_472# _321_/a_1194_69# _321_/a_3662_472#
+ _321_/a_2034_472# _321_/a_358_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_252_ vdd vss cal_itt\[0\] _073_ _252_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_100 vdd vss FILLER_0_18_100/VPW vdd FILLER_0_18_100/a_36_472# FILLER_0_18_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss FILLER_0_18_177/VPW vdd FILLER_0_18_177/a_1916_375# FILLER_0_18_177/a_1380_472#
+ FILLER_0_18_177/a_3260_375# FILLER_0_18_177/a_36_472# FILLER_0_18_177/a_932_472#
+ FILLER_0_18_177/a_2812_375# FILLER_0_18_177/a_2276_472# FILLER_0_18_177/a_1828_472#
+ FILLER_0_18_177/a_3172_472# FILLER_0_18_177/a_572_375# FILLER_0_18_177/a_2724_472#
+ FILLER_0_18_177/a_124_375# FILLER_0_18_177/a_1468_375# FILLER_0_18_177/a_1020_375#
+ FILLER_0_18_177/a_484_472# FILLER_0_18_177/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ _304_/VPW vdd _304_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] _235_/VPW vdd _235_/a_255_603# _235_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd _218_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss FILLER_0_16_37/VPW vdd FILLER_0_16_37/a_36_472# FILLER_0_16_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss output17/VPW vdd output17/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss output28/VPW vdd output28/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss output39/VPW vdd output39/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss FILLER_0_13_212/VPW vdd FILLER_0_13_212/a_1380_472# FILLER_0_13_212/a_36_472#
+ FILLER_0_13_212/a_932_472# FILLER_0_13_212/a_572_375# FILLER_0_13_212/a_124_375#
+ FILLER_0_13_212/a_1468_375# FILLER_0_13_212/a_1020_375# FILLER_0_13_212/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ _397_/VPW vdd _397_/a_36_472# _397_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss FILLER_0_14_81/VPW vdd FILLER_0_14_81/a_36_472# FILLER_0_14_81/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout63 net63 vss vdd net64 fanout63/VPW vdd fanout63/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ _320_/VPW vdd _320_/a_1792_472# _320_/a_224_472#
+ _320_/a_1568_472# _320_/a_36_472# _320_/a_1120_472# _320_/a_672_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_28 vdd vss FILLER_0_10_28/VPW vdd FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 vss net74 net82 vdd fanout74/VPW vdd fanout74/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net52 vss vdd net57 fanout52/VPW vdd fanout52/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ _251_/VPW vdd _251_/a_468_472# _251_/a_244_472#
+ _251_/a_1130_472# _251_/a_906_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_449_ _038_ en_co_clk net55 vss net72 vdd _449_/VPW vdd _449_/a_2665_112# _449_/a_448_472#
+ _449_/a_796_472# _449_/a_36_151# _449_/a_1204_472# _449_/a_3041_156# _449_/a_1000_472#
+ _449_/a_1308_423# _449_/a_1456_156# _449_/a_1288_156# _449_/a_2248_156# _449_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ _303_/VPW vdd _303_/a_36_472# _303_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd _234_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_217_ vss net26 _052_ vdd _217_/VPW vdd _217_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_181 vdd vss FILLER_0_14_181/VPW vdd FILLER_0_14_181/a_36_472# FILLER_0_14_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 ctlp[1] net18 vdd vss output18/VPW vdd output18/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss output29/VPW vdd output29/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd ANTENNA_fanout80_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ _396_/VPW vdd _396_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout53 net53 vss vdd net56 fanout53/VPW vdd fanout53/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_250_ vss _072_ _071_ vdd _250_/VPW vdd _250_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 vss net75 net76 vdd fanout75/VPW vdd fanout75/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd fanout64/VPW vdd fanout64/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd _448_/VPW vdd _448_/a_2665_112# _448_/a_448_472#
+ _448_/a_796_472# _448_/a_36_151# _448_/a_1204_472# _448_/a_3041_156# _448_/a_1000_472#
+ _448_/a_1308_423# _448_/a_1456_156# _448_/a_1288_156# _448_/a_2248_156# _448_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ _379_/VPW vdd _379_/a_36_472#
+ _379_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_302_ vdd vss _012_ _093_ _110_ _302_/VPW vdd _302_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss FILLER_0_21_28/VPW vdd FILLER_0_21_28/a_1916_375# FILLER_0_21_28/a_1380_472#
+ FILLER_0_21_28/a_3260_375# FILLER_0_21_28/a_36_472# FILLER_0_21_28/a_932_472# FILLER_0_21_28/a_2812_375#
+ FILLER_0_21_28/a_2276_472# FILLER_0_21_28/a_1828_472# FILLER_0_21_28/a_3172_472#
+ FILLER_0_21_28/a_572_375# FILLER_0_21_28/a_2724_472# FILLER_0_21_28/a_124_375# FILLER_0_21_28/a_1468_375#
+ FILLER_0_21_28/a_1020_375# FILLER_0_21_28/a_484_472# FILLER_0_21_28/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__216__A2 vss net36 vdd ANTENNA__216__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ vss net39 _063_ vdd _233_/VPW vdd _233_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss FILLER_0_15_116/VPW vdd FILLER_0_15_116/a_36_472# FILLER_0_15_116/a_572_375#
+ FILLER_0_15_116/a_124_375# FILLER_0_15_116/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd ANTENNA__373__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_216_ vdd vss _052_ mask\[9\] net36 _216_/VPW vdd _216_/a_255_603# _216_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_146 vdd vss FILLER_0_7_146/VPW vdd FILLER_0_7_146/a_36_472# FILLER_0_7_146/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 ctlp[2] net19 vdd vss output19/VPW vdd output19/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss FILLER_0_7_59/VPW vdd FILLER_0_7_59/a_36_472# FILLER_0_7_59/a_572_375#
+ FILLER_0_7_59/a_124_375# FILLER_0_7_59/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss FILLER_0_16_255/VPW vdd FILLER_0_16_255/a_36_472# FILLER_0_16_255/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss FILLER_0_0_130/VPW vdd FILLER_0_0_130/a_36_472# FILLER_0_0_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss FILLER_0_8_263/VPW vdd FILLER_0_8_263/a_36_472# FILLER_0_8_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss FILLER_0_14_50/VPW vdd FILLER_0_14_50/a_36_472# FILLER_0_14_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ _395_/VPW vdd _395_/a_1492_488# _395_/a_244_68#
+ _395_/a_1044_488# _395_/a_636_68# _395_/a_36_488# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss FILLER_0_4_49/VPW vdd FILLER_0_4_49/a_36_472# FILLER_0_4_49/a_572_375#
+ FILLER_0_4_49/a_124_375# FILLER_0_4_49/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 fanout54/VPW vdd fanout54/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd fanout76/VPW vdd fanout76/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd fanout65/VPW vdd fanout65/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss FILLER_0_19_28/VPW vdd FILLER_0_19_28/a_36_472# FILLER_0_19_28/a_572_375#
+ FILLER_0_19_28/a_124_375# FILLER_0_19_28/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd _447_/VPW vdd _447_/a_2665_112# _447_/a_448_472#
+ _447_/a_796_472# _447_/a_36_151# _447_/a_1204_472# _447_/a_3041_156# _447_/a_1000_472#
+ _447_/a_1308_423# _447_/a_1456_156# _447_/a_1288_156# _447_/a_2248_156# _447_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_2 vdd vss FILLER_0_3_2/VPW vdd FILLER_0_3_2/a_36_472# FILLER_0_3_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ vdd vss _033_ _160_ _165_ _378_/VPW vdd _378_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ _301_/VPW vdd _301_/a_36_472# _301_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd ANTENNA_output17_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] _232_/VPW vdd _232_/a_255_603# _232_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd _215_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss FILLER_0_11_142/VPW vdd FILLER_0_11_142/a_36_472# FILLER_0_11_142/a_572_375#
+ FILLER_0_11_142/a_124_375# FILLER_0_11_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss FILLER_0_2_93/VPW vdd FILLER_0_2_93/a_36_472# FILLER_0_2_93/a_572_375#
+ FILLER_0_2_93/a_124_375# FILLER_0_2_93/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss FILLER_0_17_72/VPW vdd FILLER_0_17_72/a_1916_375# FILLER_0_17_72/a_1380_472#
+ FILLER_0_17_72/a_3260_375# FILLER_0_17_72/a_36_472# FILLER_0_17_72/a_932_472# FILLER_0_17_72/a_2812_375#
+ FILLER_0_17_72/a_2276_472# FILLER_0_17_72/a_1828_472# FILLER_0_17_72/a_3172_472#
+ FILLER_0_17_72/a_572_375# FILLER_0_17_72/a_2724_472# FILLER_0_17_72/a_124_375# FILLER_0_17_72/a_1468_375#
+ FILLER_0_17_72/a_1020_375# FILLER_0_17_72/a_484_472# FILLER_0_17_72/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss FILLER_0_3_172/VPW vdd FILLER_0_3_172/a_1916_375# FILLER_0_3_172/a_1380_472#
+ FILLER_0_3_172/a_3260_375# FILLER_0_3_172/a_36_472# FILLER_0_3_172/a_932_472# FILLER_0_3_172/a_2812_375#
+ FILLER_0_3_172/a_2276_472# FILLER_0_3_172/a_1828_472# FILLER_0_3_172/a_3172_472#
+ FILLER_0_3_172/a_572_375# FILLER_0_3_172/a_2724_472# FILLER_0_3_172/a_124_375# FILLER_0_3_172/a_1468_375#
+ FILLER_0_3_172/a_1020_375# FILLER_0_3_172/a_484_472# FILLER_0_3_172/a_2364_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd ANTENNA_output47_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] _394_/VPW vdd _394_/a_244_524# _394_/a_2215_68#
+ _394_/a_56_524# _394_/a_718_524# _394_/a_728_93# _394_/a_1936_472# _394_/a_1336_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 fanout55/VPW vdd fanout55/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss FILLER_0_5_212/VPW vdd FILLER_0_5_212/a_36_472# FILLER_0_5_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd fanout77/VPW vdd fanout77/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd _446_/VPW vdd _446_/a_2665_112# _446_/a_448_472#
+ _446_/a_796_472# _446_/a_36_151# _446_/a_1204_472# _446_/a_3041_156# _446_/a_1000_472#
+ _446_/a_1308_423# _446_/a_1456_156# _446_/a_1288_156# _446_/a_2248_156# _446_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout66 vss net66 net68 vdd fanout66/VPW vdd fanout66/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ _377_/VPW vdd _377_/a_36_472# _377_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd vss _011_ _104_ _109_ _300_/VPW vdd _300_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ _231_/VPW vdd _231_/a_652_68# _231_/a_244_68# vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd _429_/VPW vdd _429_/a_2665_112# _429_/a_448_472#
+ _429_/a_796_472# _429_/a_36_151# _429_/a_1204_472# _429_/a_3041_156# _429_/a_1000_472#
+ _429_/a_1308_423# _429_/a_1456_156# _429_/a_1288_156# _429_/a_2248_156# _429_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd input1/VPW vdd input1/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd _214_/VPW vdd _214_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss FILLER_0_7_104/VPW vdd FILLER_0_7_104/a_1380_472# FILLER_0_7_104/a_36_472#
+ FILLER_0_7_104/a_932_472# FILLER_0_7_104/a_572_375# FILLER_0_7_104/a_124_375# FILLER_0_7_104/a_1468_375#
+ FILLER_0_7_104/a_1020_375# FILLER_0_7_104/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss FILLER_0_4_107/VPW vdd FILLER_0_4_107/a_1380_472# FILLER_0_4_107/a_36_472#
+ FILLER_0_4_107/a_932_472# FILLER_0_4_107/a_572_375# FILLER_0_4_107/a_124_375# FILLER_0_4_107/a_1468_375#
+ FILLER_0_4_107/a_1020_375# FILLER_0_4_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss FILLER_0_24_290/VPW vdd FILLER_0_24_290/a_36_472# FILLER_0_24_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss FILLER_0_15_290/VPW vdd FILLER_0_15_290/a_36_472# FILLER_0_15_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss FILLER_0_0_198/VPW vdd FILLER_0_0_198/a_36_472# FILLER_0_0_198/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ _393_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd fanout78/VPW vdd fanout78/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd fanout56/VPW vdd fanout56/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd fanout67/VPW vdd fanout67/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd _445_/VPW vdd _445_/a_2665_112# _445_/a_448_472#
+ _445_/a_796_472# _445_/a_36_151# _445_/a_1204_472# _445_/a_3041_156# _445_/a_1000_472#
+ _445_/a_1308_423# _445_/a_1456_156# _445_/a_1288_156# _445_/a_2248_156# _445_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vss _164_ _163_ vdd _376_/VPW vdd _376_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd vss _062_ _060_ _061_ _230_/VPW vdd _230_/a_652_68# _230_/a_244_68# vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vss FILLER_0_5_72/VPW vdd FILLER_0_5_72/a_1380_472# FILLER_0_5_72/a_36_472#
+ FILLER_0_5_72/a_932_472# FILLER_0_5_72/a_572_375# FILLER_0_5_72/a_124_375# FILLER_0_5_72/a_1468_375#
+ FILLER_0_5_72/a_1020_375# FILLER_0_5_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ _017_ state\[2\] net53 vss net70 vdd _428_/VPW vdd _428_/a_2665_112# _428_/a_448_472#
+ _428_/a_796_472# _428_/a_36_151# _428_/a_1204_472# _428_/a_3041_156# _428_/a_1000_472#
+ _428_/a_1308_423# _428_/a_1456_156# _428_/a_1288_156# _428_/a_2248_156# _428_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd vss FILLER_0_11_64/VPW vdd FILLER_0_11_64/a_36_472# FILLER_0_11_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ _359_/VPW vdd _359_/a_1492_488# _359_/a_244_68#
+ _359_/a_1044_488# _359_/a_636_68# _359_/a_36_488# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vss net2 clk vdd input2/VPW vdd input2/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output22_I vss net22 vdd ANTENNA_output22_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 _213_/VPW vdd _213_/a_255_603# _213_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_177 vdd vss FILLER_0_20_177/VPW vdd FILLER_0_20_177/a_1380_472# FILLER_0_20_177/a_36_472#
+ FILLER_0_20_177/a_932_472# FILLER_0_20_177/a_572_375# FILLER_0_20_177/a_124_375#
+ FILLER_0_20_177/a_1468_375# FILLER_0_20_177/a_1020_375# FILLER_0_20_177/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_206 vdd vss FILLER_0_13_206/VPW vdd FILLER_0_13_206/a_36_472# FILLER_0_13_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss FILLER_0_13_228/VPW vdd FILLER_0_13_228/a_36_472# FILLER_0_13_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss _392_/VPW vdd _392_/a_36_68# _392_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__282__I vss _098_ vdd ANTENNA__282__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 vss net79 net81 vdd fanout79/VPW vdd fanout79/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_2 vdd vss FILLER_0_12_2/VPW vdd FILLER_0_12_2/a_36_472# FILLER_0_12_2/a_572_375#
+ FILLER_0_12_2/a_124_375# FILLER_0_12_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout68 vss net68 net69 vdd fanout68/VPW vdd fanout68/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 vss net57 net65 vdd fanout57/VPW vdd fanout57/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd _444_/VPW vdd _444_/a_2665_112# _444_/a_448_472#
+ _444_/a_796_472# _444_/a_36_151# _444_/a_1204_472# _444_/a_3041_156# _444_/a_1000_472#
+ _444_/a_1308_423# _444_/a_1456_156# _444_/a_1288_156# _444_/a_2248_156# _444_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] _375_/VPW vdd _375_/a_36_68# _375_/a_1612_497#
+ _375_/a_692_497# _375_/a_1388_497# _375_/a_960_497# vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__277__I vss _093_ vdd ANTENNA__277__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd vss FILLER_0_18_139/VPW vdd FILLER_0_18_139/a_1380_472# FILLER_0_18_139/a_36_472#
+ FILLER_0_18_139/a_932_472# FILLER_0_18_139/a_572_375# FILLER_0_18_139/a_124_375#
+ FILLER_0_18_139/a_1468_375# FILLER_0_18_139/a_1020_375# FILLER_0_18_139/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_161 vdd vss FILLER_0_17_161/VPW vdd FILLER_0_17_161/a_36_472# FILLER_0_17_161/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ _016_ state\[1\] net53 vdd vss net70 _427_/VPW vdd _427_/a_2665_112# _427_/a_448_472#
+ _427_/a_796_472# _427_/a_36_151# _427_/a_1204_472# _427_/a_3041_156# _427_/a_1000_472#
+ _427_/a_1308_423# _427_/a_2248_156# _427_/a_2560_156# vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_358_ vdd vss _053_ _151_ _358_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd ANTENNA__385__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ _289_/VPW vdd _289_/a_36_472# _289_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd input3/VPW vdd input3/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd _212_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd ANTENNA_output15_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss FILLER_0_22_86/VPW vdd FILLER_0_22_86/a_1380_472# FILLER_0_22_86/a_36_472#
+ FILLER_0_22_86/a_932_472# FILLER_0_22_86/a_572_375# FILLER_0_22_86/a_124_375# FILLER_0_22_86/a_1468_375#
+ FILLER_0_22_86/a_1020_375# FILLER_0_22_86/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss FILLER_0_11_101/VPW vdd FILLER_0_11_101/a_36_472# FILLER_0_11_101/a_572_375#
+ FILLER_0_11_101/a_124_375# FILLER_0_11_101/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss FILLER_0_17_64/VPW vdd FILLER_0_17_64/a_36_472# FILLER_0_17_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss FILLER_0_3_142/VPW vdd FILLER_0_3_142/a_36_472# FILLER_0_3_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ _391_/VPW vdd _391_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 vss net69 net74 vdd fanout69/VPW vdd fanout69/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net58 vss vdd net59 fanout58/VPW vdd fanout58/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_374_ vdd _061_ _056_ _162_ calibrate vss _374_/VPW vdd _374_/a_36_68# _374_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd _443_/VPW vdd _443_/a_2665_112# _443_/a_448_472#
+ _443_/a_796_472# _443_/a_36_151# _443_/a_1204_472# _443_/a_3041_156# _443_/a_1000_472#
+ _443_/a_1308_423# _443_/a_1456_156# _443_/a_1288_156# _443_/a_2248_156# _443_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_107 vdd vss FILLER_0_18_107/VPW vdd FILLER_0_18_107/a_1916_375# FILLER_0_18_107/a_1380_472#
+ FILLER_0_18_107/a_3260_375# FILLER_0_18_107/a_36_472# FILLER_0_18_107/a_932_472#
+ FILLER_0_18_107/a_2812_375# FILLER_0_18_107/a_2276_472# FILLER_0_18_107/a_1828_472#
+ FILLER_0_18_107/a_3172_472# FILLER_0_18_107/a_572_375# FILLER_0_18_107/a_2724_472#
+ FILLER_0_18_107/a_124_375# FILLER_0_18_107/a_1468_375# FILLER_0_18_107/a_1020_375#
+ FILLER_0_18_107/a_484_472# FILLER_0_18_107/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd ANTENNA__394__A3/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ _288_/VPW vdd _288_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ _357_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ _015_ state\[0\] net64 vss net81 vdd _426_/VPW vdd _426_/a_2665_112# _426_/a_448_472#
+ _426_/a_796_472# _426_/a_36_151# _426_/a_1204_472# _426_/a_3041_156# _426_/a_1000_472#
+ _426_/a_1308_423# _426_/a_1456_156# _426_/a_1288_156# _426_/a_2248_156# _426_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 vss net4 en vdd input4/VPW vdd input4/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_211_ vss net24 _050_ vdd _211_/VPW vdd _211_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ _409_/VPW vdd _409_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd vss FILLER_0_11_135/VPW vdd FILLER_0_11_135/a_36_472# FILLER_0_11_135/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vss FILLER_0_11_124/VPW vdd FILLER_0_11_124/a_36_472# FILLER_0_11_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss FILLER_0_15_282/VPW vdd FILLER_0_15_282/a_36_472# FILLER_0_15_282/a_572_375#
+ FILLER_0_15_282/a_124_375# FILLER_0_15_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd ANTENNA__413__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ _390_/VPW vdd _390_/a_36_68# _390_/a_244_472#
+ _390_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss FILLER_0_14_99/VPW vdd FILLER_0_14_99/a_36_472# FILLER_0_14_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 fanout59/VPW vdd fanout59/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ _373_/VPW vdd _373_/a_438_68#
+ _373_/a_244_68# _373_/a_1254_68# _373_/a_1060_68# _373_/a_632_68# _373_/a_1458_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd _442_/VPW vdd _442_/a_2665_112# _442_/a_448_472#
+ _442_/a_796_472# _442_/a_36_151# _442_/a_1204_472# _442_/a_3041_156# _442_/a_1000_472#
+ _442_/a_1308_423# _442_/a_1456_156# _442_/a_1288_156# _442_/a_2248_156# _442_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ _356_/VPW vdd _356_/a_36_472# _356_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ _287_/VPW vdd _287_/a_36_472# _287_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss FILLER_0_11_78/VPW vdd FILLER_0_11_78/a_36_472# FILLER_0_11_78/a_572_375#
+ FILLER_0_11_78/a_124_375# FILLER_0_11_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd input5/VPW vdd input5/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd _425_/VPW vdd _425_/a_2665_112# _425_/a_448_472#
+ _425_/a_796_472# _425_/a_36_151# _425_/a_1204_472# _425_/a_3041_156# _425_/a_1000_472#
+ _425_/a_1308_423# _425_/a_1456_156# _425_/a_1288_156# _425_/a_2248_156# _425_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 _210_/VPW vdd _210_/a_255_603# _210_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss FILLER_0_20_169/VPW vdd FILLER_0_20_169/a_36_472# FILLER_0_20_169/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] _408_/VPW vdd _408_/a_244_524# _408_/a_2215_68#
+ _408_/a_56_524# _408_/a_718_524# _408_/a_728_93# _408_/a_1936_472# _408_/a_1336_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd _339_/VPW vdd _339_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd ANTENNA_output20_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss FILLER_0_21_286/VPW vdd FILLER_0_21_286/a_36_472# FILLER_0_21_286/a_572_375#
+ FILLER_0_21_286/a_124_375# FILLER_0_21_286/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss FILLER_0_12_220/VPW vdd FILLER_0_12_220/a_1380_472# FILLER_0_12_220/a_36_472#
+ FILLER_0_12_220/a_932_472# FILLER_0_12_220/a_572_375# FILLER_0_12_220/a_124_375#
+ FILLER_0_12_220/a_1468_375# FILLER_0_12_220/a_1020_375# FILLER_0_12_220/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss FILLER_0_8_247/VPW vdd FILLER_0_8_247/a_1380_472# FILLER_0_8_247/a_36_472#
+ FILLER_0_8_247/a_932_472# FILLER_0_8_247/a_572_375# FILLER_0_8_247/a_124_375# FILLER_0_8_247/a_1468_375#
+ FILLER_0_8_247/a_1020_375# FILLER_0_8_247/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 net49 vss vdd net50 fanout49/VPW vdd fanout49/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_206 vdd vss FILLER_0_5_206/VPW vdd FILLER_0_5_206/a_36_472# FILLER_0_5_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd _441_/VPW vdd _441_/a_2665_112# _441_/a_448_472#
+ _441_/a_796_472# _441_/a_36_151# _441_/a_1204_472# _441_/a_3041_156# _441_/a_1000_472#
+ _441_/a_1308_423# _441_/a_1456_156# _441_/a_1288_156# _441_/a_2248_156# _441_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ _372_/VPW vdd _372_/a_2590_472# _372_/a_170_472#
+ _372_/a_1602_69# _372_/a_786_69# _372_/a_3126_472# _372_/a_1194_69# _372_/a_3662_472#
+ _372_/a_2034_472# _372_/a_358_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__303__A2 vss _098_ vdd ANTENNA__303__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vss FILLER_0_17_142/VPW vdd FILLER_0_17_142/a_36_472# FILLER_0_17_142/a_572_375#
+ FILLER_0_17_142/a_124_375# FILLER_0_17_142/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_54 vdd vss FILLER_0_5_54/VPW vdd FILLER_0_5_54/a_1380_472# FILLER_0_5_54/a_36_472#
+ FILLER_0_5_54/a_932_472# FILLER_0_5_54/a_572_375# FILLER_0_5_54/a_124_375# FILLER_0_5_54/a_1468_375#
+ FILLER_0_5_54/a_1020_375# FILLER_0_5_54/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_355_ vdd vss _149_ _026_ _355_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd _424_/VPW vdd _424_/a_2665_112# _424_/a_448_472#
+ _424_/a_796_472# _424_/a_36_151# _424_/a_1204_472# _424_/a_3041_156# _424_/a_1000_472#
+ _424_/a_1308_423# _424_/a_1456_156# _424_/a_1288_156# _424_/a_2248_156# _424_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ vdd vss _005_ _094_ _101_ _286_/VPW vdd _286_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_123 vdd vss FILLER_0_14_123/VPW vdd FILLER_0_14_123/a_36_472# FILLER_0_14_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ _338_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ _407_/VPW vdd _407_/a_36_472# _407_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ _269_/VPW vdd _269_/a_36_472# _269_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss FILLER_0_17_56/VPW vdd FILLER_0_17_56/a_36_472# FILLER_0_17_56/a_572_375#
+ FILLER_0_17_56/a_124_375# FILLER_0_17_56/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd ANTENNA_input4_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vss _032_ _159_ vdd _371_/VPW vdd _371_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd _440_/VPW vdd _440_/a_2665_112# _440_/a_448_472#
+ _440_/a_796_472# _440_/a_36_151# _440_/a_1204_472# _440_/a_3041_156# _440_/a_1000_472#
+ _440_/a_1308_423# _440_/a_1456_156# _440_/a_1288_156# _440_/a_2248_156# _440_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd vss FILLER_0_5_88/VPW vdd FILLER_0_5_88/a_36_472# FILLER_0_5_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ _012_ net35 net55 vss net72 vdd _423_/VPW vdd _423_/a_2665_112# _423_/a_448_472#
+ _423_/a_796_472# _423_/a_36_151# _423_/a_1204_472# _423_/a_3041_156# _423_/a_1000_472#
+ _423_/a_1308_423# _423_/a_1456_156# _423_/a_1288_156# _423_/a_2248_156# _423_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ _354_/VPW vdd _354_/a_49_472#
+ _354_/a_665_69# _354_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_285_ net28 vdd vss _101_ mask\[1\] _099_ _285_/VPW vdd _285_/a_36_472# _285_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_199_ net20 vss vdd _046_ _199_/VPW vdd _199_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ _337_/VPW vdd _337_/a_49_472#
+ _337_/a_665_69# _337_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] _406_/VPW vdd _406_/a_36_159# vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ _268_/VPW vdd _268_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss FILLER_0_24_274/VPW vdd FILLER_0_24_274/a_1380_472# FILLER_0_24_274/a_36_472#
+ FILLER_0_24_274/a_932_472# FILLER_0_24_274/a_572_375# FILLER_0_24_274/a_124_375#
+ FILLER_0_24_274/a_1468_375# FILLER_0_24_274/a_1020_375# FILLER_0_24_274/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ _370_/VPW vdd _370_/a_848_380# _370_/a_1084_68#
+ _370_/a_124_24# _370_/a_1152_472# _370_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd ANTENNA_fanout55_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss FILLER_0_1_266/VPW vdd FILLER_0_1_266/a_36_472# FILLER_0_1_266/a_572_375#
+ FILLER_0_1_266/a_124_375# FILLER_0_1_266/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_422_ _011_ net34 net61 vss net78 vdd _422_/VPW vdd _422_/a_2665_112# _422_/a_448_472#
+ _422_/a_796_472# _422_/a_36_151# _422_/a_1204_472# _422_/a_3041_156# _422_/a_1000_472#
+ _422_/a_1308_423# _422_/a_1456_156# _422_/a_1288_156# _422_/a_2248_156# _422_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_353_ vdd vss _148_ _025_ _353_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss FILLER_0_17_133/VPW vdd FILLER_0_17_133/a_36_472# FILLER_0_17_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output36_I vss net36 vdd ANTENNA_output36_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_284_ vdd vss _004_ _094_ _100_ _284_/VPW vdd _284_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_198_ vdd vss _046_ mask\[3\] net30 _198_/VPW vdd _198_/a_255_603# _198_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_336_ vdd vss _138_ _018_ _336_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] _405_/VPW vdd _405_/a_255_603# _405_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] _267_/VPW vdd _267_/a_1792_472# _267_/a_224_472#
+ _267_/a_1568_472# _267_/a_36_472# _267_/a_1120_472# _267_/a_672_472# vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss FILLER_0_6_177/VPW vdd FILLER_0_6_177/a_36_472# FILLER_0_6_177/a_572_375#
+ FILLER_0_6_177/a_124_375# FILLER_0_6_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ _319_/VPW vdd _319_/a_234_472# _319_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss FILLER_0_8_239/VPW vdd FILLER_0_8_239/a_36_472# FILLER_0_8_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss FILLER_0_1_212/VPW vdd FILLER_0_1_212/a_36_472# FILLER_0_1_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd _421_/VPW vdd _421_/a_2665_112# _421_/a_448_472#
+ _421_/a_796_472# _421_/a_36_151# _421_/a_1204_472# _421_/a_3041_156# _421_/a_1000_472#
+ _421_/a_1308_423# _421_/a_1456_156# _421_/a_1288_156# _421_/a_2248_156# _421_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ _352_/VPW vdd _352_/a_49_472#
+ _352_/a_665_69# _352_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ _283_/VPW vdd _283_/a_36_472# _283_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vdd vss FILLER_0_9_142/VPW vdd FILLER_0_9_142/a_36_472# FILLER_0_9_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vss FILLER_0_20_107/VPW vdd FILLER_0_20_107/a_36_472# FILLER_0_20_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ _404_/VPW vdd _404_/a_36_472# _404_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ _335_/VPW vdd _335_/a_49_472#
+ _335_/a_665_69# _335_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_266_ vdd vss _055_ _085_ _266_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_197_ vdd vss net19 net9 _197_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd _249_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vss cal_count\[3\] vdd ANTENNA__409__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd vss _124_ _115_ _118_ _318_/VPW vdd _318_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd vss FILLER_0_8_24/VPW vdd FILLER_0_8_24/a_36_472# FILLER_0_8_24/a_572_375#
+ FILLER_0_8_24/a_124_375# FILLER_0_8_24/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd ANTENNA__251__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss FILLER_0_8_2/VPW vdd FILLER_0_8_2/a_36_472# FILLER_0_8_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd ANTENNA_input2_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd _420_/VPW vdd _420_/a_2665_112# _420_/a_448_472#
+ _420_/a_796_472# _420_/a_36_151# _420_/a_1204_472# _420_/a_3041_156# _420_/a_1000_472#
+ _420_/a_1308_423# _420_/a_1456_156# _420_/a_1288_156# _420_/a_2248_156# _420_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ _351_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd _282_/VPW vdd _282_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd ANTENNA__390__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_334_ vss _137_ _132_ vdd _334_/VPW vdd _334_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_403_ vdd vss _183_ cal_count\[2\] _176_ _403_/VPW vdd _403_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vss net41 vdd ANTENNA_output41_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vss FILLER_0_6_90/VPW vdd FILLER_0_6_90/a_36_472# FILLER_0_6_90/a_572_375#
+ FILLER_0_6_90/a_124_375# FILLER_0_6_90/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net19 vss vdd _045_ _196_/VPW vdd _196_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ _265_/VPW vdd _265_/a_468_472#
+ _265_/a_224_472# _265_/a_244_68# _265_/a_916_472# vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd ANTENNA__395__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd vss FILLER_0_17_38/VPW vdd FILLER_0_17_38/a_36_472# FILLER_0_17_38/a_572_375#
+ FILLER_0_17_38/a_124_375# FILLER_0_17_38/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_248_ vss _070_ _069_ vdd _248_/VPW vdd _248_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__409__A2 vss _077_ vdd ANTENNA__409__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd _317_/VPW vdd _317_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss FILLER_0_2_171/VPW vdd FILLER_0_2_171/a_36_472# FILLER_0_2_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss FILLER_0_12_236/VPW vdd FILLER_0_12_236/a_36_472# FILLER_0_12_236/a_572_375#
+ FILLER_0_12_236/a_124_375# FILLER_0_12_236/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ _350_/VPW vdd _350_/a_49_472#
+ _350_/a_665_69# _350_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ _281_/VPW vdd _281_/a_234_472# _281_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd ANTENNA__237__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd _333_/VPW vdd _333_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 _195_/VPW vdd _195_/a_255_603# _195_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] _402_/VPW vdd _402_/a_244_567# _402_/a_718_527#
+ _402_/a_2172_497# _402_/a_56_567# _402_/a_1948_68# _402_/a_728_93# _402_/a_1296_93#
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss FILLER_0_11_109/VPW vdd FILLER_0_11_109/a_36_472# FILLER_0_11_109/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] _264_/VPW vdd _264_/a_224_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd ANTENNA__372__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss FILLER_0_12_50/VPW vdd FILLER_0_12_50/a_36_472# FILLER_0_12_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ _247_/VPW vdd _247_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate _316_/VPW vdd _316_/a_848_380# _316_/a_1084_68#
+ _316_/a_124_24# _316_/a_1152_472# _316_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_60 vdd vss FILLER_0_23_60/VPW vdd FILLER_0_23_60/a_36_472# FILLER_0_23_60/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vss FILLER_0_15_212/VPW vdd FILLER_0_15_212/a_1380_472# FILLER_0_15_212/a_36_472#
+ FILLER_0_15_212/a_932_472# FILLER_0_15_212/a_572_375# FILLER_0_15_212/a_124_375#
+ FILLER_0_15_212/a_1468_375# FILLER_0_15_212/a_1020_375# FILLER_0_15_212/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vss FILLER_0_8_37/VPW vdd FILLER_0_8_37/a_36_472# FILLER_0_8_37/a_572_375#
+ FILLER_0_8_37/a_124_375# FILLER_0_8_37/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss FILLER_0_17_104/VPW vdd FILLER_0_17_104/a_1380_472# FILLER_0_17_104/a_36_472#
+ FILLER_0_17_104/a_932_472# FILLER_0_17_104/a_572_375# FILLER_0_17_104/a_124_375#
+ FILLER_0_17_104/a_1468_375# FILLER_0_17_104/a_1020_375# FILLER_0_17_104/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_72 vdd vss FILLER_0_15_72/VPW vdd FILLER_0_15_72/a_36_472# FILLER_0_15_72/a_572_375#
+ FILLER_0_15_72/a_124_375# FILLER_0_15_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd vss FILLER_0_1_204/VPW vdd FILLER_0_1_204/a_36_472# FILLER_0_1_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ _280_/VPW vdd _280_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss FILLER_0_14_107/VPW vdd FILLER_0_14_107/a_1380_472# FILLER_0_14_107/a_36_472#
+ FILLER_0_14_107/a_932_472# FILLER_0_14_107/a_572_375# FILLER_0_14_107/a_124_375#
+ FILLER_0_14_107/a_1468_375# FILLER_0_14_107/a_1020_375# FILLER_0_14_107/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ vdd _180_ _179_ _181_ _174_ vss _401_/VPW vdd _401_/a_36_68# _401_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_332_ _126_ vdd vss _017_ _127_ _135_ _332_/VPW vdd _332_/a_36_472# _332_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_194_ vss net8 net18 vdd _194_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ _263_/VPW vdd _263_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss FILLER_0_5_181/VPW vdd FILLER_0_5_181/a_36_472# FILLER_0_5_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_246_ vss _068_ _055_ vdd _246_/VPW vdd _246_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss _315_/VPW vdd _315_/a_36_68# _315_/a_244_497#
+ _315_/a_1657_68# _315_/a_1229_68# _315_/a_716_497# vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_290 vdd vss FILLER_0_23_290/VPW vdd FILLER_0_23_290/a_36_472# FILLER_0_23_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss FILLER_0_15_235/VPW vdd FILLER_0_15_235/a_36_472# FILLER_0_15_235/a_572_375#
+ FILLER_0_15_235/a_124_375# FILLER_0_15_235/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ _229_/VPW vdd _229_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss FILLER_0_18_61/VPW vdd FILLER_0_18_61/a_36_472# FILLER_0_18_61/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss FILLER_0_11_282/VPW vdd FILLER_0_11_282/a_36_472# FILLER_0_11_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd ANTENNA_fanout76_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss FILLER_0_4_213/VPW vdd FILLER_0_4_213/a_36_472# FILLER_0_4_213/a_572_375#
+ FILLER_0_4_213/a_124_375# FILLER_0_4_213/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ vdd vss _180_ cal_count\[1\] _178_ _400_/VPW vdd _400_/a_245_68# vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_193_ net18 vss vdd _044_ _193_/VPW vdd _193_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_331_ _134_ vdd vss _135_ _086_ _132_ _331_/VPW vdd _331_/a_448_472# _331_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ _262_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd ANTENNA__303__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ vdd vss _121_ _085_ _069_ _314_/VPW vdd _314_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_245_ vdd vss net6 _067_ net67 _245_/VPW vdd _245_/a_234_472# _245_/a_672_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_206 vdd vss FILLER_0_21_206/VPW vdd FILLER_0_21_206/a_36_472# FILLER_0_21_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd _228_/VPW vdd _228_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss FILLER_0_7_233/VPW vdd FILLER_0_7_233/a_36_472# FILLER_0_7_233/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss FILLER_0_9_60/VPW vdd FILLER_0_9_60/a_36_472# FILLER_0_9_60/a_572_375#
+ FILLER_0_9_60/a_124_375# FILLER_0_9_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vss FILLER_0_13_142/VPW vdd FILLER_0_13_142/a_1380_472# FILLER_0_13_142/a_36_472#
+ FILLER_0_13_142/a_932_472# FILLER_0_13_142/a_572_375# FILLER_0_13_142/a_124_375#
+ FILLER_0_13_142/a_1468_375# FILLER_0_13_142/a_1020_375# FILLER_0_13_142/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ vdd vss _044_ mask\[1\] net28 _192_/VPW vdd _192_/a_255_603# _192_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_261_ vss _081_ _059_ vdd _261_/VPW vdd _261_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_330_ vdd vss _134_ _133_ _062_ _330_/VPW vdd _330_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss FILLER_0_12_20/VPW vdd FILLER_0_12_20/a_36_472# FILLER_0_12_20/a_572_375#
+ FILLER_0_12_20/a_124_375# FILLER_0_12_20/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss FILLER_0_5_172/VPW vdd FILLER_0_5_172/a_36_472# FILLER_0_5_172/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ vdd vss en_co_clk _067_ _244_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__190__I vss _043_ vdd ANTENNA__190__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_313_ vdd vss _120_ _059_ _119_ _313_/VPW vdd _313_/a_255_603# _313_/a_67_603# vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__257__A1 vss _053_ vdd ANTENNA__257__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd _227_/VPW vdd _227_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd ANTENNA__402__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss FILLER_0_20_31/VPW vdd FILLER_0_20_31/a_36_472# FILLER_0_20_31/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss FILLER_0_9_72/VPW vdd FILLER_0_9_72/a_1380_472# FILLER_0_9_72/a_36_472#
+ FILLER_0_9_72/a_932_472# FILLER_0_9_72/a_572_375# FILLER_0_9_72/a_124_375# FILLER_0_9_72/a_1468_375#
+ FILLER_0_9_72/a_1020_375# FILLER_0_9_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss FILLER_0_0_96/VPW vdd FILLER_0_0_96/a_36_472# FILLER_0_0_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss _260_/VPW vdd _260_/a_36_68# _260_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ _389_/VPW vdd _389_/a_428_148# _389_/a_36_148#
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 _191_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ _312_/VPW vdd _312_/a_234_472# _312_/a_672_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd vss net47 net42 _243_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd vss FILLER_0_23_282/VPW vdd FILLER_0_23_282/a_36_472# FILLER_0_23_282/a_572_375#
+ FILLER_0_23_282/a_124_375# FILLER_0_23_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss FILLER_0_15_205/VPW vdd FILLER_0_15_205/a_36_472# FILLER_0_15_205/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss FILLER_0_2_165/VPW vdd FILLER_0_2_165/a_36_472# FILLER_0_2_165/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss FILLER_0_18_53/VPW vdd FILLER_0_18_53/a_36_472# FILLER_0_18_53/a_572_375#
+ FILLER_0_18_53/a_124_375# FILLER_0_18_53/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ _226_/VPW vdd _226_/a_1044_68# _226_/a_452_68#
+ _226_/a_276_68# _226_/a_860_68# vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd ANTENNA__426__CLK/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_98 vdd vss FILLER_0_20_98/VPW vdd FILLER_0_20_98/a_36_472# FILLER_0_20_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_87 vdd vss FILLER_0_20_87/VPW vdd FILLER_0_20_87/a_36_472# FILLER_0_20_87/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 _209_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss FILLER_0_19_171/VPW vdd FILLER_0_19_171/a_1380_472# FILLER_0_19_171/a_36_472#
+ FILLER_0_19_171/a_932_472# FILLER_0_19_171/a_572_375# FILLER_0_19_171/a_124_375#
+ FILLER_0_19_171/a_1468_375# FILLER_0_19_171/a_1020_375# FILLER_0_19_171/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd ANTENNA__302__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss FILLER_0_15_10/VPW vdd FILLER_0_15_10/a_36_472# FILLER_0_15_10/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss FILLER_0_15_2/VPW vdd FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_572_375#
+ FILLER_0_15_2/a_124_375# FILLER_0_15_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss FILLER_0_22_177/VPW vdd FILLER_0_22_177/a_1380_472# FILLER_0_22_177/a_36_472#
+ FILLER_0_22_177/a_932_472# FILLER_0_22_177/a_572_375# FILLER_0_22_177/a_124_375#
+ FILLER_0_22_177/a_1468_375# FILLER_0_22_177/a_1020_375# FILLER_0_22_177/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss FILLER_0_13_100/VPW vdd FILLER_0_13_100/a_36_472# FILLER_0_13_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss FILLER_0_9_105/VPW vdd FILLER_0_9_105/a_36_472# FILLER_0_9_105/a_572_375#
+ FILLER_0_9_105/a_124_375# FILLER_0_9_105/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ _190_/VPW vdd _190_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ _388_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd ANTENNA_output18_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ _311_/VPW vdd _311_/a_692_473# _311_/a_254_473#
+ _311_/a_66_473# _311_/a_2700_473# _311_/a_1660_473# _311_/a_3220_473# _311_/a_1212_473#
+ _311_/a_2180_473# _311_/a_3740_473# _311_/a_1920_473# vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_242_ net47 vss vdd _066_ _242_/VPW vdd _242_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_228 vdd vss FILLER_0_15_228/VPW vdd FILLER_0_15_228/a_36_472# FILLER_0_15_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss FILLER_0_2_111/VPW vdd FILLER_0_2_111/a_1380_472# FILLER_0_2_111/a_36_472#
+ FILLER_0_2_111/a_932_472# FILLER_0_2_111/a_572_375# FILLER_0_2_111/a_124_375# FILLER_0_2_111/a_1468_375#
+ FILLER_0_2_111/a_1020_375# FILLER_0_2_111/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss FILLER_0_2_177/VPW vdd FILLER_0_2_177/a_36_472# FILLER_0_2_177/a_572_375#
+ FILLER_0_2_177/a_124_375# FILLER_0_2_177/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd _225_/VPW vdd _225_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss FILLER_0_18_76/VPW vdd FILLER_0_18_76/a_36_472# FILLER_0_18_76/a_572_375#
+ FILLER_0_18_76/a_124_375# FILLER_0_18_76/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ _208_/VPW vdd _208_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd _387_/VPW vdd _387_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_310_ _090_ vdd vss _117_ _060_ _113_ _310_/VPW vdd _310_/a_49_472# _310_/a_1133_69#
+ _310_/a_741_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_164 vdd vss FILLER_0_5_164/VPW vdd FILLER_0_5_164/a_36_472# FILLER_0_5_164/a_572_375#
+ FILLER_0_5_164/a_124_375# FILLER_0_5_164/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd vss FILLER_0_23_88/VPW vdd FILLER_0_23_88/a_36_472# FILLER_0_23_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss FILLER_0_23_44/VPW vdd FILLER_0_23_44/a_1380_472# FILLER_0_23_44/a_36_472#
+ FILLER_0_23_44/a_932_472# FILLER_0_23_44/a_572_375# FILLER_0_23_44/a_124_375# FILLER_0_23_44/a_1468_375#
+ FILLER_0_23_44/a_1020_375# FILLER_0_23_44/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] _241_/VPW vdd _241_/a_224_472# vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd _439_/VPW vdd _439_/a_2665_112# _439_/a_448_472#
+ _439_/a_796_472# _439_/a_36_151# _439_/a_1204_472# _439_/a_3041_156# _439_/a_1000_472#
+ _439_/a_1308_423# _439_/a_1456_156# _439_/a_1288_156# _439_/a_2248_156# _439_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd vss FILLER_0_2_101/VPW vdd FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss FILLER_0_3_54/VPW vdd FILLER_0_3_54/a_36_472# FILLER_0_3_54/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd _224_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd vss _049_ mask\[6\] net33 _207_/VPW vdd _207_/a_255_603# _207_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss FILLER_0_19_195/VPW vdd FILLER_0_19_195/a_36_472# FILLER_0_19_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss FILLER_0_0_232/VPW vdd FILLER_0_0_232/a_36_472# FILLER_0_0_232/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss FILLER_0_16_154/VPW vdd FILLER_0_16_154/a_1380_472# FILLER_0_16_154/a_36_472#
+ FILLER_0_16_154/a_932_472# FILLER_0_16_154/a_572_375# FILLER_0_16_154/a_124_375#
+ FILLER_0_16_154/a_1468_375# FILLER_0_16_154/a_1020_375# FILLER_0_16_154/a_484_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd ANTENNA__257__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd ANTENNA__220__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss FILLER_0_20_2/VPW vdd FILLER_0_20_2/a_36_472# FILLER_0_20_2/a_572_375#
+ FILLER_0_20_2/a_124_375# FILLER_0_20_2/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ _386_/VPW vdd _386_/a_848_380# _386_/a_1084_68#
+ _386_/a_124_24# _386_/a_1152_472# _386_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss FILLER_0_5_198/VPW vdd FILLER_0_5_198/a_36_472# FILLER_0_5_198/a_572_375#
+ FILLER_0_5_198/a_124_375# FILLER_0_5_198/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_240_ vdd vss net41 net46 _240_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_282 vdd vss FILLER_0_17_282/VPW vdd FILLER_0_17_282/a_36_472# FILLER_0_17_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_274 vdd vss FILLER_0_23_274/VPW vdd FILLER_0_23_274/a_36_472# FILLER_0_23_274/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd _438_/VPW vdd _438_/a_2665_112# _438_/a_448_472#
+ _438_/a_796_472# _438_/a_36_151# _438_/a_1204_472# _438_/a_3041_156# _438_/a_1000_472#
+ _438_/a_1308_423# _438_/a_1456_156# _438_/a_1288_156# _438_/a_2248_156# _438_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ _369_/VPW vdd _369_/a_36_68# _369_/a_244_472#
+ _369_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd ANTENNA_output23_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss FILLER_0_14_263/VPW vdd FILLER_0_14_263/a_36_472# FILLER_0_14_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] _223_/VPW vdd _223_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss FILLER_0_9_290/VPW vdd FILLER_0_9_290/a_36_472# FILLER_0_9_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 _206_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss FILLER_0_0_266/VPW vdd FILLER_0_0_266/a_36_472# FILLER_0_0_266/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss _385_/VPW vdd _385_/a_36_68# _385_/a_244_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ _299_/VPW vdd _299_/a_36_472# _299_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd _437_/VPW vdd _437_/a_2665_112# _437_/a_448_472#
+ _437_/a_796_472# _437_/a_36_151# _437_/a_1204_472# _437_/a_3041_156# _437_/a_1000_472#
+ _437_/a_1308_423# _437_/a_1456_156# _437_/a_1288_156# _437_/a_2248_156# _437_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_78 vdd vss FILLER_0_3_78/VPW vdd FILLER_0_3_78/a_36_472# FILLER_0_3_78/a_572_375#
+ FILLER_0_3_78/a_124_375# FILLER_0_3_78/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_368_ vdd vss trim_mask\[4\] _158_ _368_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_222_ vdd vss net38 net43 _222_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ _205_/VPW vdd _205_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss FILLER_0_19_142/VPW vdd FILLER_0_19_142/a_36_472# FILLER_0_19_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd _453_/VPW vdd _453_/a_2665_112# _453_/a_448_472#
+ _453_/a_796_472# _453_/a_36_151# _453_/a_1204_472# _453_/a_3041_156# _453_/a_1000_472#
+ _453_/a_1308_423# _453_/a_1456_156# _453_/a_1288_156# _453_/a_2248_156# _453_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ _384_/VPW vdd _384_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss FILLER_0_10_107/VPW vdd FILLER_0_10_107/a_36_472# FILLER_0_10_107/a_572_375#
+ FILLER_0_10_107/a_124_375# FILLER_0_10_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ _298_/VPW vdd _298_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd _436_/VPW vdd _436_/a_2665_112# _436_/a_448_472#
+ _436_/a_796_472# _436_/a_36_151# _436_/a_1204_472# _436_/a_3041_156# _436_/a_1000_472#
+ _436_/a_1308_423# _436_/a_1456_156# _436_/a_1288_156# _436_/a_2248_156# _436_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd ANTENNA__408__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ _367_/VPW vdd _367_/a_36_68# _367_/a_244_472#
+ _367_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss FILLER_0_13_80/VPW vdd FILLER_0_13_80/a_36_472# FILLER_0_13_80/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss FILLER_0_1_192/VPW vdd FILLER_0_1_192/a_36_472# FILLER_0_1_192/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd vss FILLER_0_9_270/VPW vdd FILLER_0_9_270/a_36_472# FILLER_0_9_270/a_572_375#
+ FILLER_0_9_270/a_124_375# FILLER_0_9_270/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vss net38 _054_ vdd _221_/VPW vdd _221_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ _008_ net31 net60 vss net77 vdd _419_/VPW vdd _419_/a_2665_112# _419_/a_448_472#
+ _419_/a_796_472# _419_/a_36_151# _419_/a_1204_472# _419_/a_3041_156# _419_/a_1000_472#
+ _419_/a_1308_423# _419_/a_1456_156# _419_/a_1288_156# _419_/a_2248_156# _419_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 _204_/VPW vdd _204_/a_255_603# _204_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss FILLER_0_20_15/VPW vdd FILLER_0_20_15/a_1380_472# FILLER_0_20_15/a_36_472#
+ FILLER_0_20_15/a_932_472# FILLER_0_20_15/a_572_375# FILLER_0_20_15/a_124_375# FILLER_0_20_15/a_1468_375#
+ FILLER_0_20_15/a_1020_375# FILLER_0_20_15/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss FILLER_0_19_187/VPW vdd FILLER_0_19_187/a_36_472# FILLER_0_19_187/a_572_375#
+ FILLER_0_19_187/a_124_375# FILLER_0_19_187/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss FILLER_0_3_221/VPW vdd FILLER_0_3_221/a_1380_472# FILLER_0_3_221/a_36_472#
+ FILLER_0_3_221/a_932_472# FILLER_0_3_221/a_572_375# FILLER_0_3_221/a_124_375# FILLER_0_3_221/a_1468_375#
+ FILLER_0_3_221/a_1020_375# FILLER_0_3_221/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss FILLER_0_15_59/VPW vdd FILLER_0_15_59/a_36_472# FILLER_0_15_59/a_572_375#
+ FILLER_0_15_59/a_124_375# FILLER_0_15_59/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vss net59 vdd ANTENNA_fanout58_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd vss FILLER_0_6_79/VPW vdd FILLER_0_6_79/a_36_472# FILLER_0_6_79/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 _452_/VPW vdd _452_/a_448_472# _452_/a_36_151#
+ _452_/a_1293_527# _452_/a_3081_151# _452_/a_1284_156# _452_/a_1040_527# _452_/a_1353_112#
+ _452_/a_836_156# _452_/a_1697_156# _452_/a_2449_156# _452_/a_3129_107# _452_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ _383_/VPW vdd _383_/a_36_472#
+ _383_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ _297_/VPW vdd _297_/a_36_472# _297_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd _435_/VPW vdd _435_/a_2665_112# _435_/a_448_472#
+ _435_/a_796_472# _435_/a_36_151# _435_/a_1204_472# _435_/a_3041_156# _435_/a_1000_472#
+ _435_/a_1308_423# _435_/a_1456_156# _435_/a_1288_156# _435_/a_2248_156# _435_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A2 vss cal_count\[3\] vdd ANTENNA__408__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ vdd vss trim_mask\[3\] _157_ _366_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_127 vdd vss FILLER_0_2_127/VPW vdd FILLER_0_2_127/a_36_472# FILLER_0_2_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vss FILLER_0_18_37/VPW vdd FILLER_0_18_37/a_1380_472# FILLER_0_18_37/a_36_472#
+ FILLER_0_18_37/a_932_472# FILLER_0_18_37/a_572_375# FILLER_0_18_37/a_124_375# FILLER_0_18_37/a_1468_375#
+ FILLER_0_18_37/a_1020_375# FILLER_0_18_37/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vss FILLER_0_9_282/VPW vdd FILLER_0_9_282/a_36_472# FILLER_0_9_282/a_572_375#
+ FILLER_0_9_282/a_124_375# FILLER_0_9_282/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd vss _054_ trim_val\[0\] _053_ _220_/VPW vdd _220_/a_255_603# _220_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_349_ vdd vss _146_ _023_ _349_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _007_ net30 net60 vss net77 vdd _418_/VPW vdd _418_/a_2665_112# _418_/a_448_472#
+ _418_/a_796_472# _418_/a_36_151# _418_/a_1204_472# _418_/a_3041_156# _418_/a_1000_472#
+ _418_/a_1308_423# _418_/a_1456_156# _418_/a_1288_156# _418_/a_2248_156# _418_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output21_I vss net21 vdd ANTENNA_output21_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 _203_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss FILLER_0_19_155/VPW vdd FILLER_0_19_155/a_36_472# FILLER_0_19_155/a_572_375#
+ FILLER_0_19_155/a_124_375# FILLER_0_19_155/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss FILLER_0_19_111/VPW vdd FILLER_0_19_111/a_36_472# FILLER_0_19_111/a_572_375#
+ FILLER_0_19_111/a_124_375# FILLER_0_19_111/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss FILLER_0_22_128/VPW vdd FILLER_0_22_128/a_1916_375# FILLER_0_22_128/a_1380_472#
+ FILLER_0_22_128/a_3260_375# FILLER_0_22_128/a_36_472# FILLER_0_22_128/a_932_472#
+ FILLER_0_22_128/a_2812_375# FILLER_0_22_128/a_2276_472# FILLER_0_22_128/a_1828_472#
+ FILLER_0_22_128/a_3172_472# FILLER_0_22_128/a_572_375# FILLER_0_22_128/a_2724_472#
+ FILLER_0_22_128/a_124_375# FILLER_0_22_128/a_1468_375# FILLER_0_22_128/a_1020_375#
+ FILLER_0_22_128/a_484_472# FILLER_0_22_128/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss FILLER_0_15_180/VPW vdd FILLER_0_15_180/a_36_472# FILLER_0_15_180/a_572_375#
+ FILLER_0_15_180/a_124_375# FILLER_0_15_180/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss FILLER_0_21_150/VPW vdd FILLER_0_21_150/a_36_472# FILLER_0_21_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss FILLER_0_6_47/VPW vdd FILLER_0_6_47/a_1916_375# FILLER_0_6_47/a_1380_472#
+ FILLER_0_6_47/a_3260_375# FILLER_0_6_47/a_36_472# FILLER_0_6_47/a_932_472# FILLER_0_6_47/a_2812_375#
+ FILLER_0_6_47/a_2276_472# FILLER_0_6_47/a_1828_472# FILLER_0_6_47/a_3172_472# FILLER_0_6_47/a_572_375#
+ FILLER_0_6_47/a_2724_472# FILLER_0_6_47/a_124_375# FILLER_0_6_47/a_1468_375# FILLER_0_6_47/a_1020_375#
+ FILLER_0_6_47/a_484_472# FILLER_0_6_47/a_2364_375# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 _451_/VPW vdd _451_/a_448_472# _451_/a_36_151#
+ _451_/a_1293_527# _451_/a_3081_151# _451_/a_1284_156# _451_/a_1040_527# _451_/a_1353_112#
+ _451_/a_836_156# _451_/a_1697_156# _451_/a_2449_156# _451_/a_3129_107# _451_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_28 vdd vss FILLER_0_12_28/VPW vdd FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd vss _035_ _160_ _167_ _382_/VPW vdd _382_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss FILLER_0_18_209/VPW vdd FILLER_0_18_209/a_36_472# FILLER_0_18_209/a_572_375#
+ FILLER_0_18_209/a_124_375# FILLER_0_18_209/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss FILLER_0_5_136/VPW vdd FILLER_0_5_136/a_36_472# FILLER_0_5_136/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ _296_/VPW vdd _296_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd _434_/VPW vdd _434_/a_2665_112# _434_/a_448_472#
+ _434_/a_796_472# _434_/a_36_151# _434_/a_1204_472# _434_/a_3041_156# _434_/a_1000_472#
+ _434_/a_1308_423# _434_/a_1456_156# _434_/a_1288_156# _434_/a_2248_156# _434_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ _365_/VPW vdd _365_/a_36_68# _365_/a_244_472#
+ _365_/a_692_472# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd ANTENNA__280__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd ANTENNA__240__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ _348_/VPW vdd _348_/a_49_472#
+ _348_/a_665_69# _348_/a_257_69# vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd _417_/VPW vdd _417_/a_2665_112# _417_/a_448_472#
+ _417_/a_796_472# _417_/a_36_151# _417_/a_1204_472# _417_/a_3041_156# _417_/a_1000_472#
+ _417_/a_1308_423# _417_/a_1456_156# _417_/a_1288_156# _417_/a_2248_156# _417_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_279_ vdd vss _096_ _090_ state\[1\] _279_/VPW vdd _279_/a_652_68# _279_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_231 vdd vss FILLER_0_6_231/VPW vdd FILLER_0_6_231/a_36_472# FILLER_0_6_231/a_572_375#
+ FILLER_0_6_231/a_124_375# FILLER_0_6_231/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ _202_/VPW vdd _202_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output14_I vss net14 vdd ANTENNA_output14_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd vss FILLER_0_4_91/VPW vdd FILLER_0_4_91/a_36_472# FILLER_0_4_91/a_572_375#
+ FILLER_0_4_91/a_124_375# FILLER_0_4_91/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_94 vdd vss FILLER_0_10_94/VPW vdd FILLER_0_10_94/a_36_472# FILLER_0_10_94/a_572_375#
+ FILLER_0_10_94/a_124_375# FILLER_0_10_94/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss FILLER_0_3_212/VPW vdd FILLER_0_3_212/a_36_472# FILLER_0_3_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss FILLER_0_19_134/VPW vdd FILLER_0_19_134/a_36_472# FILLER_0_19_134/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss FILLER_0_16_115/VPW vdd FILLER_0_16_115/a_36_472# FILLER_0_16_115/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss FILLER_0_22_107/VPW vdd FILLER_0_22_107/a_36_472# FILLER_0_22_107/a_572_375#
+ FILLER_0_22_107/a_124_375# FILLER_0_22_107/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss FILLER_0_21_60/VPW vdd FILLER_0_21_60/a_36_472# FILLER_0_21_60/a_572_375#
+ FILLER_0_21_60/a_124_375# FILLER_0_21_60/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss FILLER_0_6_37/VPW vdd FILLER_0_6_37/a_36_472# FILLER_0_6_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd vss FILLER_0_8_156/VPW vdd FILLER_0_8_156/a_36_472# FILLER_0_8_156/a_572_375#
+ FILLER_0_8_156/a_124_375# FILLER_0_8_156/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I vss rstn vdd ANTENNA_input5_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__243__I vss net47 vdd ANTENNA__243__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 _450_/VPW vdd _450_/a_448_472# _450_/a_36_151#
+ _450_/a_1293_527# _450_/a_3081_151# _450_/a_1284_156# _450_/a_1040_527# _450_/a_1353_112#
+ _450_/a_836_156# _450_/a_1697_156# _450_/a_2449_156# _450_/a_3129_107# _450_/a_2225_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xoutput40 trim[2] net40 vdd vss output40/VPW vdd output40/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ _381_/VPW vdd _381_/a_36_472#
+ _381_/a_244_68# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_148 vdd vss FILLER_0_5_148/VPW vdd FILLER_0_5_148/a_36_472# FILLER_0_5_148/a_572_375#
+ FILLER_0_5_148/a_124_375# FILLER_0_5_148/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd _433_/VPW vdd _433_/a_2665_112# _433_/a_448_472#
+ _433_/a_796_472# _433_/a_36_151# _433_/a_1204_472# _433_/a_3041_156# _433_/a_1000_472#
+ _433_/a_1308_423# _433_/a_1456_156# _433_/a_1288_156# _433_/a_2248_156# _433_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ _295_/VPW vdd _295_/a_36_472# _295_/a_244_68#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ _364_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss FILLER_0_14_235/VPW vdd FILLER_0_14_235/a_36_472# FILLER_0_14_235/a_572_375#
+ FILLER_0_14_235/a_124_375# FILLER_0_14_235/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss FILLER_0_13_72/VPW vdd FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_572_375#
+ FILLER_0_13_72/a_124_375# FILLER_0_13_72/a_484_472# vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_347_ vdd vss _145_ _022_ _347_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 _278_/VPW vdd _278_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_290 vdd vss FILLER_0_13_290/VPW vdd FILLER_0_13_290/a_36_472# FILLER_0_13_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ _005_ net28 net62 vss net79 vdd _416_/VPW vdd _416_/a_2665_112# _416_/a_448_472#
+ _416_/a_796_472# _416_/a_36_151# _416_/a_1204_472# _416_/a_3041_156# _416_/a_1000_472#
+ _416_/a_1308_423# _416_/a_1456_156# _416_/a_1288_156# _416_/a_2248_156# _416_/a_2560_156#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_201_ vdd vss _047_ mask\[4\] net31 _201_/VPW vdd _201_/a_255_603# _201_/a_67_603#
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd ANTENNA__448__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 result[3] net30 vdd vss output30/VPW vdd output30/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_196 vdd vss FILLER_0_12_196/VPW vdd FILLER_0_12_196/a_36_472# FILLER_0_12_196/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 clkc net6 vdd vss output6/VPW vdd output6/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss output41/VPW vdd output41/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ _380_/VPW vdd _380_/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
C0 net52 _386_/a_124_24# 0.001051f
C1 mask\[8\] _437_/a_2665_112# 0.007907f
C2 _012_ FILLER_0_23_60/a_36_472# 0.001572f
C3 FILLER_0_21_28/a_1468_375# vdd -0.008892f
C4 _129_ _160_ 0.001631f
C5 _320_/a_36_472# _043_ 0.019162f
C6 net15 vss 1.330044f
C7 _132_ FILLER_0_16_115/a_124_375# 0.033245f
C8 FILLER_0_11_78/a_484_472# vdd 0.001756f
C9 FILLER_0_11_78/a_36_472# vss 0.00471f
C10 ctlp[2] _420_/a_2665_112# 0.01544f
C11 net55 FILLER_0_21_28/a_3172_472# 0.06297f
C12 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_572_375# 0.086635f
C13 _265_/a_244_68# cal_itt\[0\] 0.003127f
C14 net82 FILLER_0_4_213/a_36_472# 0.003042f
C15 FILLER_0_17_200/a_484_472# mask\[3\] 0.014805f
C16 FILLER_0_7_162/a_124_375# _169_ 0.00336f
C17 net17 trim[3] 0.001664f
C18 net66 _167_ 0.016569f
C19 net63 _435_/a_1308_423# 0.003621f
C20 FILLER_0_22_86/a_932_472# _026_ 0.001587f
C21 net28 _094_ 0.007842f
C22 _055_ _113_ 0.153988f
C23 _125_ _062_ 0.061735f
C24 FILLER_0_8_127/a_36_472# _070_ 0.005078f
C25 _093_ FILLER_0_17_104/a_1468_375# 0.010965f
C26 FILLER_0_23_44/a_1380_472# vss 0.003905f
C27 net39 _054_ 0.049797f
C28 FILLER_0_4_107/a_1020_375# net47 0.011446f
C29 _414_/a_1308_423# cal_itt\[3\] 0.044184f
C30 FILLER_0_12_136/a_124_375# state\[2\] 0.001029f
C31 FILLER_0_12_136/a_1020_375# net53 0.002709f
C32 _051_ net71 0.001617f
C33 FILLER_0_5_164/a_572_375# net37 0.014025f
C34 FILLER_0_18_209/a_124_375# _047_ 0.006317f
C35 FILLER_0_6_90/a_36_472# vdd 0.00366f
C36 FILLER_0_6_90/a_572_375# vss 0.006421f
C37 FILLER_0_2_171/a_124_375# net22 0.009924f
C38 _091_ net57 0.006076f
C39 _328_/a_36_113# FILLER_0_11_109/a_36_472# 0.0161f
C40 _159_ FILLER_0_2_127/a_124_375# 0.020951f
C41 net29 _005_ 0.020239f
C42 mask\[5\] FILLER_0_20_177/a_572_375# 0.013294f
C43 _418_/a_2248_156# vdd 0.00423f
C44 _273_/a_36_68# net4 0.06843f
C45 fanout74/a_36_113# FILLER_0_3_142/a_124_375# 0.002073f
C46 output14/a_224_472# _442_/a_36_151# 0.172111f
C47 _305_/a_36_159# _425_/a_36_151# 0.001404f
C48 _132_ FILLER_0_19_111/a_572_375# 0.01675f
C49 FILLER_0_18_2/a_1916_375# net38 0.006403f
C50 mask\[8\] net14 0.040566f
C51 net52 FILLER_0_9_72/a_36_472# 0.014911f
C52 _116_ _071_ 0.017991f
C53 _122_ FILLER_0_5_181/a_36_472# 0.003016f
C54 ctlp[6] net23 0.006951f
C55 net81 FILLER_0_15_235/a_36_472# 0.001855f
C56 FILLER_0_13_142/a_1468_375# net23 0.011746f
C57 _445_/a_2665_112# net17 0.006445f
C58 _036_ _446_/a_2248_156# 0.001763f
C59 ctlp[1] FILLER_0_24_290/a_124_375# 0.050488f
C60 net39 vss 0.170972f
C61 net20 _418_/a_2248_156# 0.003507f
C62 FILLER_0_1_266/a_484_472# vss 0.001113f
C63 _445_/a_2665_112# trim_val\[1\] 0.015206f
C64 net51 vss 0.21065f
C65 _126_ _113_ 0.547055f
C66 _425_/a_448_472# net37 0.002755f
C67 _077_ FILLER_0_8_156/a_124_375# 0.00407f
C68 FILLER_0_24_274/a_36_472# FILLER_0_23_274/a_36_472# 0.05841f
C69 FILLER_0_16_89/a_36_472# _176_ 0.012173f
C70 FILLER_0_7_72/a_2364_375# net50 0.017301f
C71 cal_count\[3\] _134_ 0.011364f
C72 net32 mask\[7\] 0.01969f
C73 ctlp[5] _140_ 0.002123f
C74 net81 vss 0.766885f
C75 ctln[2] net65 0.113266f
C76 FILLER_0_18_2/a_932_472# net44 0.012286f
C77 net52 _453_/a_2248_156# 0.011419f
C78 FILLER_0_18_2/a_1828_472# vdd 0.001953f
C79 FILLER_0_18_2/a_1380_472# vss -0.001894f
C80 _144_ net35 0.036236f
C81 FILLER_0_4_177/a_124_375# _386_/a_848_380# 0.001277f
C82 FILLER_0_11_109/a_36_472# _120_ 0.014554f
C83 _432_/a_36_151# net80 0.035794f
C84 _402_/a_1948_68# cal_count\[1\] 0.037053f
C85 _137_ FILLER_0_19_155/a_572_375# 0.030256f
C86 _360_/a_36_160# _163_ 0.008593f
C87 cal_itt\[3\] FILLER_0_6_177/a_572_375# 0.00225f
C88 _413_/a_796_472# vdd 0.001569f
C89 FILLER_0_1_98/a_36_472# vdd 0.009937f
C90 net82 net37 0.037195f
C91 result[5] net61 0.092275f
C92 FILLER_0_19_125/a_124_375# net73 0.005414f
C93 _442_/a_36_151# FILLER_0_2_127/a_36_472# 0.012873f
C94 net48 calibrate 0.482314f
C95 net64 mask\[2\] 0.046428f
C96 net82 FILLER_0_3_221/a_1468_375# 0.009095f
C97 _119_ _118_ 0.001596f
C98 _140_ _433_/a_36_151# 0.020943f
C99 _350_/a_49_472# vss 0.001319f
C100 FILLER_0_8_247/a_1020_375# calibrate 0.008393f
C101 vdd _022_ 0.082842f
C102 trim_val\[4\] net59 0.062701f
C103 result[7] FILLER_0_23_274/a_36_472# 0.014434f
C104 FILLER_0_9_223/a_124_375# net4 0.061757f
C105 ctlp[1] FILLER_0_24_274/a_1380_472# 0.008573f
C106 _065_ _447_/a_448_472# 0.049072f
C107 FILLER_0_1_204/a_124_375# vdd 0.047704f
C108 _079_ _263_/a_224_472# 0.002505f
C109 output26/a_224_472# _423_/a_36_151# 0.011936f
C110 FILLER_0_5_212/a_36_472# vss 0.00578f
C111 FILLER_0_3_172/a_2724_472# net22 0.012284f
C112 FILLER_0_8_37/a_484_472# _220_/a_67_603# 0.005759f
C113 ctln[1] net65 0.073241f
C114 _094_ net77 0.00405f
C115 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_36_472# 0.086635f
C116 FILLER_0_12_136/a_1380_472# _127_ 0.001432f
C117 _106_ vss 0.180823f
C118 _422_/a_2560_156# mask\[7\] 0.010664f
C119 FILLER_0_12_20/a_572_375# net40 0.007477f
C120 FILLER_0_19_55/a_36_472# _012_ 0.001667f
C121 net35 net25 0.129685f
C122 _181_ _185_ 0.061846f
C123 net35 net23 0.04007f
C124 FILLER_0_19_125/a_36_472# _132_ 0.008568f
C125 _412_/a_2560_156# en 0.049213f
C126 net30 result[3] 0.002746f
C127 net38 vdd 0.906502f
C128 FILLER_0_15_290/a_124_375# net79 0.051113f
C129 _427_/a_796_472# _095_ 0.007281f
C130 net62 FILLER_0_15_290/a_36_472# 0.009046f
C131 net75 FILLER_0_8_247/a_1380_472# 0.020589f
C132 _232_/a_67_603# _160_ 0.001684f
C133 net16 _186_ 0.225785f
C134 _228_/a_36_68# vss 0.031389f
C135 FILLER_0_4_123/a_36_472# _160_ 0.050308f
C136 net38 FILLER_0_20_15/a_484_472# 0.003376f
C137 FILLER_0_13_65/a_36_472# FILLER_0_13_72/a_36_472# 0.002765f
C138 net74 FILLER_0_13_142/a_36_472# 0.003568f
C139 mask\[4\] _069_ 0.001182f
C140 FILLER_0_2_171/a_124_375# vdd 0.042659f
C141 FILLER_0_5_54/a_932_472# FILLER_0_6_47/a_1828_472# 0.026657f
C142 _428_/a_796_472# _017_ 0.025239f
C143 _158_ vdd 0.131365f
C144 trimb[2] net17 0.007637f
C145 _211_/a_36_160# _436_/a_36_151# 0.068534f
C146 _013_ FILLER_0_21_28/a_1828_472# 0.003978f
C147 _444_/a_36_151# net47 0.016691f
C148 net81 fanout76/a_36_160# 0.041089f
C149 output33/a_224_472# _421_/a_2665_112# 0.010726f
C150 _127_ FILLER_0_11_124/a_36_472# 0.001641f
C151 _141_ mask\[6\] 0.009844f
C152 _322_/a_1084_68# _129_ 0.00419f
C153 _390_/a_36_68# _070_ 0.047478f
C154 FILLER_0_18_107/a_484_472# vdd 0.035309f
C155 FILLER_0_18_107/a_36_472# vss 0.003245f
C156 _103_ mask\[2\] 0.002168f
C157 net57 _306_/a_36_68# 0.042596f
C158 _434_/a_1000_472# mask\[6\] 0.021582f
C159 net24 FILLER_0_22_86/a_1380_472# 0.003096f
C160 _302_/a_224_472# vss 0.005149f
C161 _414_/a_448_472# _003_ 0.023209f
C162 FILLER_0_10_78/a_932_472# net52 0.00207f
C163 output29/a_224_472# net19 0.09445f
C164 FILLER_0_7_104/a_36_472# vss 0.002797f
C165 FILLER_0_7_104/a_484_472# vdd 0.021325f
C166 ctlp[3] net61 0.007397f
C167 _424_/a_36_151# vdd 0.125156f
C168 FILLER_0_18_139/a_1380_472# _145_ 0.002077f
C169 net66 vdd 0.646189f
C170 _426_/a_36_151# net19 0.04851f
C171 _277_/a_36_160# vss 0.030147f
C172 _074_ _162_ 0.112872f
C173 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_124_375# 0.003732f
C174 net81 _195_/a_67_603# 0.002322f
C175 net55 FILLER_0_21_60/a_484_472# 0.098472f
C176 _067_ vdd 0.853589f
C177 net78 net77 0.252376f
C178 mask\[3\] output34/a_224_472# 0.002385f
C179 net50 _441_/a_36_151# 0.060777f
C180 net52 _441_/a_1308_423# 0.059264f
C181 FILLER_0_4_107/a_124_375# _153_ 0.073219f
C182 FILLER_0_4_107/a_1020_375# _154_ 0.013746f
C183 FILLER_0_12_28/a_124_375# net40 0.047331f
C184 FILLER_0_19_47/a_36_472# FILLER_0_18_37/a_1020_375# 0.001684f
C185 _088_ FILLER_0_3_212/a_36_472# 0.005583f
C186 FILLER_0_12_236/a_36_472# _060_ 0.014046f
C187 _068_ _160_ 0.003424f
C188 _053_ trim_mask\[0\] 0.007667f
C189 fanout60/a_36_160# vdd 0.090968f
C190 _162_ _076_ 0.008623f
C191 _407_/a_36_472# _181_ 0.035594f
C192 net2 vss 0.213737f
C193 _030_ _168_ 0.015729f
C194 _181_ cal_count\[0\] 0.001114f
C195 net18 _417_/a_448_472# 0.03772f
C196 _417_/a_36_151# result[3] 0.006379f
C197 _417_/a_1308_423# net30 0.007538f
C198 output10/a_224_472# _411_/a_36_151# 0.001362f
C199 _091_ FILLER_0_13_212/a_932_472# 0.008749f
C200 _086_ _151_ 0.002442f
C201 _072_ _375_/a_1612_497# 0.002646f
C202 ctlp[1] _010_ 0.002794f
C203 _441_/a_796_472# _030_ 0.024278f
C204 _256_/a_1164_497# net4 0.004729f
C205 net31 mask\[4\] 0.499009f
C206 cal net58 0.001209f
C207 _437_/a_2248_156# vdd 0.054674f
C208 result[7] FILLER_0_24_274/a_1468_375# 0.006125f
C209 fanout75/a_36_113# _081_ 0.015843f
C210 _115_ _439_/a_2248_156# 0.003553f
C211 en_co_clk _390_/a_244_472# 0.001238f
C212 net61 _422_/a_448_472# 0.006042f
C213 FILLER_0_3_172/a_2724_472# vdd 0.006405f
C214 _129_ _133_ 0.080636f
C215 _105_ net32 2.08459f
C216 _308_/a_848_380# net14 0.021982f
C217 _415_/a_2248_156# result[1] 0.010922f
C218 _035_ net40 0.068572f
C219 mask\[3\] FILLER_0_18_171/a_124_375# 0.001156f
C220 _127_ _428_/a_2665_112# 0.001162f
C221 FILLER_0_19_171/a_932_472# _434_/a_36_151# 0.00271f
C222 FILLER_0_23_282/a_124_375# FILLER_0_23_274/a_124_375# 0.003732f
C223 fanout61/a_36_113# net62 0.031315f
C224 output9/a_224_472# en 0.011047f
C225 _258_/a_36_160# _080_ 0.261387f
C226 state\[1\] _113_ 0.107642f
C227 mask\[8\] _148_ 0.356546f
C228 _077_ _439_/a_2665_112# 0.035688f
C229 _012_ FILLER_0_23_44/a_572_375# 0.002827f
C230 net80 fanout80/a_36_113# 0.004615f
C231 result[7] _093_ 0.001096f
C232 FILLER_0_4_213/a_572_375# net59 0.061684f
C233 cal_count\[3\] FILLER_0_12_196/a_124_375# 0.007717f
C234 net41 FILLER_0_23_44/a_124_375# 0.001526f
C235 FILLER_0_3_54/a_124_375# vdd 0.029897f
C236 FILLER_0_10_78/a_572_375# vss 0.004588f
C237 _144_ _433_/a_2665_112# 0.030413f
C238 vdd rstn 0.160093f
C239 _044_ _416_/a_2665_112# 0.01372f
C240 _430_/a_1308_423# mask\[2\] 0.020226f
C241 _114_ _061_ 0.123371f
C242 net57 _395_/a_36_488# 0.026081f
C243 vss clkc 0.0311f
C244 FILLER_0_7_72/a_124_375# _053_ 0.014569f
C245 _077_ FILLER_0_8_138/a_124_375# 0.007238f
C246 _114_ _311_/a_66_473# 0.081048f
C247 _093_ _198_/a_67_603# 0.004447f
C248 FILLER_0_7_72/a_2724_472# _077_ 0.004635f
C249 FILLER_0_22_177/a_36_472# _146_ 0.002f
C250 _098_ _023_ 0.004191f
C251 _045_ vss 0.032891f
C252 FILLER_0_7_72/a_124_375# FILLER_0_6_47/a_2812_375# 0.026339f
C253 FILLER_0_22_177/a_124_375# _435_/a_36_151# 0.059049f
C254 ctlp[1] FILLER_0_23_282/a_36_472# 0.003169f
C255 FILLER_0_14_181/a_36_472# vss 0.002955f
C256 _098_ FILLER_0_20_98/a_124_375# 0.012779f
C257 net57 FILLER_0_13_142/a_1468_375# 0.011369f
C258 net61 _108_ 0.030767f
C259 net69 _160_ 0.077526f
C260 FILLER_0_2_171/a_124_375# FILLER_0_2_165/a_124_375# 0.003598f
C261 FILLER_0_15_205/a_36_472# net21 0.007503f
C262 _115_ _315_/a_244_497# 0.00153f
C263 net75 _253_/a_1100_68# 0.001047f
C264 valid vss 0.308766f
C265 _140_ FILLER_0_22_128/a_3172_472# 0.005458f
C266 net61 net19 0.132027f
C267 _322_/a_848_380# FILLER_0_9_142/a_36_472# 0.011591f
C268 net23 _433_/a_2665_112# 0.015555f
C269 FILLER_0_18_107/a_124_375# net14 0.005202f
C270 net15 _095_ 0.056214f
C271 fanout76/a_36_160# net2 0.023033f
C272 net64 FILLER_0_12_220/a_1468_375# 0.01836f
C273 net71 _436_/a_36_151# 0.03535f
C274 _002_ net59 0.016205f
C275 FILLER_0_8_247/a_36_472# vss 0.003706f
C276 FILLER_0_8_247/a_484_472# vdd 0.005485f
C277 _114_ FILLER_0_11_101/a_484_472# 0.025975f
C278 _144_ vdd 0.40911f
C279 FILLER_0_4_49/a_572_375# _440_/a_36_151# 0.073306f
C280 _075_ _414_/a_2248_156# 0.044302f
C281 _256_/a_1612_497# _068_ 0.002759f
C282 _050_ _140_ 0.001f
C283 FILLER_0_16_73/a_124_375# vss 0.026383f
C284 _269_/a_36_472# _260_/a_36_68# 0.002875f
C285 _426_/a_2248_156# _060_ 0.00106f
C286 net55 FILLER_0_18_37/a_1468_375# 0.009059f
C287 _066_ vdd 0.14893f
C288 _114_ _072_ 0.078148f
C289 FILLER_0_12_136/a_1468_375# cal_count\[3\] 0.004337f
C290 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_36_472# 0.086635f
C291 net15 _036_ 0.036489f
C292 _322_/a_848_380# _128_ 0.012288f
C293 net78 _421_/a_448_472# 0.025808f
C294 _168_ trim_mask\[3\] 0.007154f
C295 net47 _054_ 0.171966f
C296 FILLER_0_8_138/a_124_375# _120_ 0.12254f
C297 FILLER_0_16_255/a_36_472# _094_ 0.005892f
C298 _152_ _160_ 0.286108f
C299 net75 _015_ 0.025217f
C300 _374_/a_36_68# _056_ 0.011052f
C301 FILLER_0_9_28/a_484_472# vdd 0.010868f
C302 mask\[5\] FILLER_0_21_206/a_36_472# 0.019416f
C303 _430_/a_36_151# _093_ 0.00184f
C304 _075_ net37 0.001054f
C305 net38 _450_/a_1353_112# 0.02208f
C306 _011_ _422_/a_1308_423# 0.001997f
C307 _086_ _162_ 0.107276f
C308 net47 _278_/a_36_160# 0.001838f
C309 cal clk 0.033015f
C310 net4 _269_/a_36_472# 0.033296f
C311 _430_/a_2560_156# _092_ 0.001333f
C312 net25 vdd 0.195306f
C313 net23 vdd 1.576398f
C314 net45 ctlp[0] 0.001134f
C315 output26/a_224_472# FILLER_0_23_44/a_1380_472# 0.0323f
C316 trim_mask\[4\] vss 0.641217f
C317 FILLER_0_4_49/a_36_472# _160_ 0.00202f
C318 net58 sample 0.006906f
C319 comp net3 0.05248f
C320 FILLER_0_14_50/a_124_375# _181_ 0.00402f
C321 net58 net37 0.15273f
C322 FILLER_0_13_80/a_124_375# FILLER_0_13_72/a_572_375# 0.012001f
C323 _444_/a_2560_156# net67 0.012781f
C324 net47 vss 0.919407f
C325 _091_ net36 0.067629f
C326 _178_ net47 0.09023f
C327 net52 _443_/a_2560_156# 0.020855f
C328 _430_/a_448_472# mask\[2\] 0.045973f
C329 output6/a_224_472# net6 0.076605f
C330 _086_ _131_ 0.886615f
C331 FILLER_0_16_57/a_1468_375# vss 0.062643f
C332 FILLER_0_16_57/a_36_472# vdd 0.088011f
C333 _315_/a_716_497# _120_ 0.001321f
C334 output13/a_224_472# vss 0.108144f
C335 _387_/a_36_113# _037_ 0.003577f
C336 net35 _436_/a_2248_156# 0.014499f
C337 _091_ _429_/a_1204_472# 0.024554f
C338 FILLER_0_7_72/a_124_375# FILLER_0_5_72/a_36_472# 0.001512f
C339 _112_ _316_/a_124_24# 0.032665f
C340 _414_/a_2248_156# net21 0.00415f
C341 _322_/a_1084_68# _068_ 0.001022f
C342 _127_ _070_ 0.031272f
C343 net15 _449_/a_448_472# 0.040076f
C344 _012_ vss 0.454371f
C345 sample calibrate 0.001861f
C346 net41 vdd 1.983262f
C347 fanout54/a_36_160# FILLER_0_19_155/a_124_375# 0.005705f
C348 FILLER_0_15_212/a_36_472# vss 0.002853f
C349 FILLER_0_15_212/a_1020_375# mask\[1\] 0.017527f
C350 FILLER_0_10_214/a_124_375# _090_ 0.072741f
C351 net72 _452_/a_36_151# 0.040035f
C352 _093_ _303_/a_36_472# 0.096502f
C353 calibrate net37 0.101109f
C354 FILLER_0_11_109/a_124_375# vdd 0.079069f
C355 net16 _063_ 0.038576f
C356 fanout71/a_36_113# FILLER_0_20_107/a_36_472# 0.001645f
C357 _195_/a_67_603# _045_ 0.004028f
C358 _363_/a_36_68# _153_ 0.008003f
C359 net32 _419_/a_2248_156# 0.034827f
C360 FILLER_0_4_197/a_36_472# _079_ 0.002448f
C361 FILLER_0_5_172/a_36_472# vdd 0.092294f
C362 FILLER_0_5_172/a_124_375# vss 0.028247f
C363 _110_ _423_/a_2665_112# 0.001668f
C364 FILLER_0_20_169/a_36_472# _098_ 0.007354f
C365 net79 FILLER_0_15_282/a_572_375# 0.01043f
C366 trim_mask\[1\] FILLER_0_6_47/a_2364_375# 0.007169f
C367 net62 FILLER_0_15_282/a_36_472# 0.013655f
C368 _083_ _001_ 0.002625f
C369 _067_ _450_/a_1353_112# 0.007106f
C370 _025_ _352_/a_49_472# 0.003933f
C371 _258_/a_36_160# vss 0.005039f
C372 _287_/a_36_472# _099_ 0.030964f
C373 net37 net21 0.03272f
C374 ctln[1] FILLER_0_0_232/a_124_375# 0.012033f
C375 _171_ _172_ 0.104216f
C376 _052_ FILLER_0_18_53/a_572_375# 0.001631f
C377 _065_ _441_/a_2665_112# 0.003318f
C378 _074_ _076_ 0.03553f
C379 FILLER_0_15_59/a_484_472# vss 0.007866f
C380 output45/a_224_472# net43 0.024629f
C381 _254_/a_448_472# _074_ 0.002163f
C382 net32 result[8] 0.024881f
C383 ctln[5] net76 0.001707f
C384 result[6] fanout61/a_36_113# 0.003917f
C385 output48/a_224_472# net48 0.001786f
C386 FILLER_0_11_101/a_36_472# _070_ 0.033113f
C387 net65 net18 0.879399f
C388 _105_ _420_/a_2665_112# 0.001159f
C389 _133_ _068_ 0.002552f
C390 net35 FILLER_0_22_128/a_1020_375# 0.010202f
C391 net74 vss 0.589483f
C392 trim_val\[4\] FILLER_0_3_172/a_932_472# 0.001407f
C393 _415_/a_796_472# vdd 0.001842f
C394 net73 _427_/a_448_472# 0.00132f
C395 _414_/a_2560_156# cal_itt\[3\] 0.007141f
C396 _207_/a_67_603# mask\[6\] 0.072291f
C397 _376_/a_36_160# FILLER_0_6_79/a_36_472# 0.003913f
C398 _411_/a_448_472# net65 0.006279f
C399 _079_ _080_ 0.022852f
C400 net50 net16 0.015448f
C401 net58 _264_/a_224_472# 0.001803f
C402 _064_ _445_/a_1000_472# 0.015908f
C403 net57 net22 0.003595f
C404 mask\[4\] _140_ 0.001697f
C405 _397_/a_36_472# net55 0.039732f
C406 _174_ FILLER_0_15_59/a_124_375# 0.00622f
C407 net73 _145_ 0.009144f
C408 _253_/a_36_68# vss 0.002481f
C409 net61 _419_/a_448_472# 0.024246f
C410 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_572_375# 0.086635f
C411 FILLER_0_17_104/a_124_375# vdd 0.030663f
C412 _415_/a_36_151# net79 0.001156f
C413 FILLER_0_5_88/a_124_375# net47 0.005083f
C414 mask\[1\] FILLER_0_15_205/a_36_472# 0.006921f
C415 FILLER_0_15_116/a_484_472# _131_ 0.042796f
C416 ctln[2] FILLER_0_1_266/a_572_375# 0.012126f
C417 _430_/a_36_151# _136_ 0.02044f
C418 _450_/a_1040_527# clkc 0.001412f
C419 output28/a_224_472# output29/a_224_472# 0.00289f
C420 _440_/a_36_151# _029_ 0.00874f
C421 mask\[9\] _140_ 0.00126f
C422 _091_ _128_ 0.003717f
C423 trim_mask\[4\] FILLER_0_2_165/a_36_472# 0.265591f
C424 FILLER_0_12_220/a_932_472# vss 0.003677f
C425 FILLER_0_12_220/a_1380_472# vdd 0.002025f
C426 _058_ FILLER_0_8_156/a_36_472# 0.011885f
C427 _139_ net21 0.004991f
C428 FILLER_0_11_109/a_124_375# _135_ 0.009057f
C429 net58 FILLER_0_9_282/a_572_375# 0.006142f
C430 _173_ vss 0.063821f
C431 _088_ net22 0.17798f
C432 _202_/a_36_160# _047_ 0.02265f
C433 output25/a_224_472# _051_ 0.019651f
C434 _074_ FILLER_0_5_164/a_484_472# 0.003556f
C435 net39 _445_/a_796_472# 0.002296f
C436 FILLER_0_7_72/a_1916_375# FILLER_0_5_88/a_36_472# 0.0027f
C437 FILLER_0_5_72/a_932_472# _029_ 0.007801f
C438 FILLER_0_5_72/a_1468_375# trim_mask\[1\] 0.017105f
C439 FILLER_0_22_177/a_1380_472# vss 0.001502f
C440 net81 output37/a_224_472# 0.00641f
C441 net20 FILLER_0_12_220/a_1380_472# 0.029747f
C442 ctln[1] FILLER_0_1_266/a_572_375# 0.004319f
C443 _159_ vss 0.102545f
C444 mask\[9\] _424_/a_2665_112# 0.015491f
C445 FILLER_0_15_150/a_124_375# vdd 0.026143f
C446 net75 _084_ 0.045583f
C447 mask\[2\] FILLER_0_16_154/a_484_472# 0.028444f
C448 ctln[4] FILLER_0_1_204/a_36_472# 0.006408f
C449 FILLER_0_4_107/a_1380_472# _160_ 0.020979f
C450 _452_/a_1353_112# net40 0.003745f
C451 net79 _136_ 0.00111f
C452 net52 FILLER_0_0_130/a_36_472# 0.002743f
C453 FILLER_0_4_49/a_124_375# _232_/a_67_603# 0.002082f
C454 trimb[1] _452_/a_2225_156# 0.004072f
C455 FILLER_0_6_37/a_124_375# _160_ 0.04948f
C456 _016_ state\[2\] 0.002937f
C457 FILLER_0_9_223/a_484_472# _060_ 0.001529f
C458 _418_/a_1000_472# _007_ 0.001051f
C459 FILLER_0_22_86/a_36_472# _098_ 0.182093f
C460 FILLER_0_17_72/a_2812_375# _131_ 0.006589f
C461 net62 net79 1.615103f
C462 _150_ net14 0.001303f
C463 _414_/a_448_472# net76 0.002346f
C464 net55 FILLER_0_13_72/a_36_472# 0.002172f
C465 vdd FILLER_0_19_134/a_124_375# 0.027957f
C466 _154_ vss 0.200253f
C467 FILLER_0_17_72/a_3172_472# net14 0.046864f
C468 fanout73/a_36_113# vdd 0.048166f
C469 _449_/a_2665_112# vss 0.007395f
C470 _074_ _081_ 0.070546f
C471 FILLER_0_20_87/a_36_472# net71 0.003995f
C472 FILLER_0_16_107/a_572_375# _132_ 0.007439f
C473 net64 FILLER_0_9_282/a_124_375# 0.046477f
C474 mask\[0\] FILLER_0_15_212/a_1020_375# 0.001158f
C475 _151_ _163_ 0.501188f
C476 FILLER_0_3_142/a_36_472# vdd 0.10948f
C477 FILLER_0_3_142/a_124_375# vss 0.008128f
C478 _028_ FILLER_0_6_90/a_484_472# 0.01566f
C479 FILLER_0_4_144/a_124_375# _059_ 0.031451f
C480 FILLER_0_5_54/a_124_375# vdd 0.007387f
C481 _086_ _074_ 0.186795f
C482 _076_ _081_ 0.010091f
C483 _133_ _152_ 0.124374f
C484 _141_ FILLER_0_17_161/a_36_472# 0.011708f
C485 _451_/a_3129_107# _040_ 0.004116f
C486 _053_ net15 0.041871f
C487 _442_/a_1308_423# vdd 0.00782f
C488 _442_/a_448_472# vss 0.001428f
C489 FILLER_0_18_177/a_124_375# FILLER_0_20_177/a_36_472# 0.0027f
C490 _183_ _179_ 0.017086f
C491 _043_ net14 0.037706f
C492 net34 _435_/a_796_472# 0.002288f
C493 _321_/a_170_472# _129_ 0.024601f
C494 output34/a_224_472# _421_/a_2665_112# 0.00151f
C495 _070_ trim_mask\[0\] 0.006144f
C496 net15 FILLER_0_6_47/a_2812_375# 0.002944f
C497 fanout55/a_36_160# _043_ 0.019538f
C498 _098_ FILLER_0_14_235/a_124_375# 0.001228f
C499 _176_ FILLER_0_15_72/a_484_472# 0.00753f
C500 _074_ net65 0.002666f
C501 trim[0] _445_/a_36_151# 0.008302f
C502 net38 _445_/a_1308_423# 0.006454f
C503 _126_ FILLER_0_14_181/a_124_375# 0.004632f
C504 _086_ _076_ 0.79237f
C505 _413_/a_2665_112# vdd 0.02286f
C506 FILLER_0_4_152/a_36_472# net23 0.047194f
C507 _449_/a_36_151# _067_ 0.031377f
C508 ctlp[1] vss 0.32843f
C509 net68 FILLER_0_3_54/a_36_472# 0.049455f
C510 net57 vdd 1.260693f
C511 result[7] result[6] 0.119475f
C512 FILLER_0_19_47/a_36_472# _013_ 0.03573f
C513 _411_/a_2560_156# vdd 0.001315f
C514 _115_ FILLER_0_10_107/a_572_375# 0.040198f
C515 FILLER_0_14_181/a_36_472# _095_ 0.071989f
C516 _132_ _428_/a_1456_156# 0.001009f
C517 FILLER_0_19_155/a_36_472# vss 0.004125f
C518 FILLER_0_19_155/a_484_472# vdd 0.003341f
C519 _425_/a_36_151# _014_ 0.12681f
C520 _328_/a_36_113# _017_ 0.006485f
C521 fanout82/a_36_113# _122_ 0.007118f
C522 FILLER_0_7_72/a_2724_472# _308_/a_848_380# 0.001797f
C523 FILLER_0_13_65/a_36_472# net15 0.036527f
C524 _053_ FILLER_0_6_90/a_572_375# 0.073688f
C525 _413_/a_2665_112# net20 0.015855f
C526 _415_/a_36_151# net75 0.024047f
C527 _436_/a_2248_156# vdd 0.011151f
C528 FILLER_0_3_221/a_932_472# vdd 0.005654f
C529 FILLER_0_3_221/a_484_472# vss 0.005602f
C530 FILLER_0_11_124/a_36_472# _118_ 0.002798f
C531 _115_ FILLER_0_9_142/a_36_472# 0.00336f
C532 _439_/a_1204_472# vss 0.006567f
C533 _026_ net14 0.010792f
C534 net62 _429_/a_2560_156# 0.002164f
C535 _088_ vdd 0.140259f
C536 _079_ vss 0.124667f
C537 FILLER_0_22_128/a_484_472# _433_/a_36_151# 0.001653f
C538 _427_/a_3041_156# net23 0.001305f
C539 _428_/a_36_151# _043_ 0.027757f
C540 ctln[5] ctln[4] 0.031901f
C541 net20 FILLER_0_3_221/a_932_472# 0.054476f
C542 net68 _164_ 0.189377f
C543 trimb[4] vdd 0.081023f
C544 net19 FILLER_0_23_274/a_36_472# 0.075097f
C545 net56 _145_ 0.009307f
C546 _068_ _121_ 0.008802f
C547 net62 FILLER_0_13_290/a_124_375# 0.032026f
C548 net20 _088_ 0.001704f
C549 _115_ _128_ 0.263909f
C550 net14 _156_ 0.184287f
C551 _081_ FILLER_0_5_164/a_484_472# 0.001105f
C552 _004_ _415_/a_36_151# 0.013592f
C553 _093_ FILLER_0_17_133/a_124_375# 0.009649f
C554 _069_ net23 0.418375f
C555 _350_/a_49_472# _147_ 0.016114f
C556 _341_/a_49_472# mask\[3\] 0.00631f
C557 net44 FILLER_0_12_2/a_36_472# 0.011079f
C558 _443_/a_448_472# _170_ 0.056211f
C559 _077_ FILLER_0_9_72/a_1468_375# 0.008273f
C560 FILLER_0_12_2/a_484_472# vss 0.001748f
C561 _177_ vss 0.074896f
C562 net53 FILLER_0_13_142/a_572_375# 0.001597f
C563 mask\[5\] _339_/a_36_160# 0.007734f
C564 output14/a_224_472# _031_ 0.001077f
C565 net16 _039_ 0.031852f
C566 _119_ net74 0.02813f
C567 FILLER_0_10_37/a_36_472# vss 0.003659f
C568 result[4] result[3] 0.089939f
C569 FILLER_0_24_274/a_124_375# vss 0.002674f
C570 _448_/a_1308_423# _037_ 0.034533f
C571 net63 FILLER_0_18_177/a_572_375# 0.004407f
C572 _095_ net47 0.508892f
C573 trimb[1] net44 0.089379f
C574 net15 FILLER_0_5_72/a_36_472# 0.006713f
C575 _077_ _453_/a_1204_472# 0.011124f
C576 _348_/a_257_69# mask\[6\] 0.00159f
C577 FILLER_0_22_128/a_1020_375# vdd 0.002503f
C578 FILLER_0_22_128/a_572_375# vss 0.00243f
C579 _052_ FILLER_0_19_28/a_572_375# 0.011078f
C580 _217_/a_36_160# FILLER_0_19_28/a_484_472# 0.006053f
C581 _428_/a_2665_112# _118_ 0.001007f
C582 _053_ FILLER_0_5_212/a_36_472# 0.007052f
C583 _301_/a_36_472# net35 0.051887f
C584 _019_ vss 0.10954f
C585 _139_ mask\[1\] 0.017315f
C586 FILLER_0_20_15/a_1020_375# net40 0.005742f
C587 _162_ _163_ 0.011497f
C588 _257_/a_36_472# cal_itt\[3\] 0.136487f
C589 _441_/a_36_151# FILLER_0_3_78/a_124_375# 0.035849f
C590 cal_itt\[1\] vss 0.327626f
C591 cal_itt\[0\] vdd 0.438996f
C592 _359_/a_636_68# _062_ 0.001578f
C593 trim[4] net38 0.095379f
C594 _088_ FILLER_0_3_172/a_2812_375# 0.002239f
C595 FILLER_0_8_138/a_124_375# _125_ 0.001589f
C596 _031_ FILLER_0_2_127/a_36_472# 0.016207f
C597 net58 net8 0.175026f
C598 net79 net4 0.386068f
C599 _187_ vdd 0.194575f
C600 _086_ _081_ 0.033115f
C601 _028_ FILLER_0_7_104/a_932_472# 0.003084f
C602 FILLER_0_5_181/a_124_375# net37 0.005396f
C603 FILLER_0_21_206/a_36_472# _434_/a_2665_112# 0.00243f
C604 _070_ _060_ 0.822179f
C605 _140_ _022_ 0.001997f
C606 _412_/a_36_151# net75 0.060039f
C607 net67 _164_ 0.030648f
C608 _421_/a_2248_156# mask\[7\] 0.016229f
C609 _004_ net62 0.001201f
C610 _064_ _160_ 0.006705f
C611 net57 FILLER_0_2_165/a_124_375# 0.007153f
C612 _414_/a_1308_423# net22 0.011978f
C613 result[5] net62 0.041722f
C614 net29 _102_ 0.056837f
C615 ctln[6] FILLER_0_0_130/a_36_472# 0.023355f
C616 valid output37/a_224_472# 0.039402f
C617 _420_/a_36_151# FILLER_0_23_274/a_36_472# 0.001723f
C618 FILLER_0_9_282/a_484_472# vss 0.00561f
C619 FILLER_0_6_47/a_2276_472# vdd 0.002735f
C620 FILLER_0_6_47/a_1828_472# vss 0.003457f
C621 FILLER_0_7_72/a_2276_472# FILLER_0_6_90/a_124_375# 0.001684f
C622 output48/a_224_472# net37 0.095886f
C623 FILLER_0_20_31/a_124_375# net40 0.011967f
C624 FILLER_0_19_125/a_124_375# _145_ 0.006777f
C625 _141_ FILLER_0_18_139/a_1468_375# 0.005239f
C626 _053_ FILLER_0_7_104/a_36_472# 0.01752f
C627 _321_/a_170_472# FILLER_0_11_135/a_124_375# 0.001153f
C628 net74 _095_ 0.04188f
C629 cal_count\[2\] _402_/a_1948_68# 0.010022f
C630 _119_ _154_ 0.01697f
C631 FILLER_0_7_104/a_1020_375# _151_ 0.002336f
C632 net32 _421_/a_1000_472# 0.002275f
C633 mask\[0\] FILLER_0_13_206/a_124_375# 0.005989f
C634 net75 _316_/a_848_380# 0.044673f
C635 FILLER_0_13_212/a_484_472# vss 0.002397f
C636 _443_/a_36_151# net69 0.069715f
C637 net80 _339_/a_36_160# 0.016897f
C638 net55 _423_/a_36_151# 0.001124f
C639 net26 FILLER_0_21_28/a_1916_375# 0.008721f
C640 ctlp[1] _420_/a_796_472# 0.001468f
C641 _056_ net59 0.001756f
C642 _116_ _070_ 0.166494f
C643 _238_/a_67_603# output15/a_224_472# 0.019027f
C644 FILLER_0_5_109/a_484_472# vss 0.00212f
C645 FILLER_0_16_37/a_124_375# _181_ 0.001198f
C646 _446_/a_2248_156# net17 0.008375f
C647 net9 cal_itt\[0\] 0.110446f
C648 _072_ _395_/a_1492_488# 0.003088f
C649 net63 _093_ 0.109689f
C650 _136_ FILLER_0_17_133/a_124_375# 0.001315f
C651 net20 FILLER_0_13_212/a_932_472# 0.003007f
C652 vdd FILLER_0_5_148/a_572_375# -0.009701f
C653 vss FILLER_0_5_148/a_124_375# 0.018465f
C654 FILLER_0_19_187/a_484_472# vss 0.004504f
C655 output27/a_224_472# FILLER_0_9_270/a_124_375# 0.001274f
C656 net36 net22 0.034258f
C657 net73 FILLER_0_18_107/a_2812_375# 0.018753f
C658 _141_ _343_/a_257_69# 0.001515f
C659 net55 FILLER_0_17_72/a_36_472# 0.020422f
C660 _381_/a_244_68# _167_ 0.001153f
C661 FILLER_0_12_20/a_124_375# _450_/a_448_472# 0.001597f
C662 FILLER_0_2_111/a_484_472# vdd 0.005951f
C663 _429_/a_1204_472# net22 0.001899f
C664 net54 _098_ 0.116416f
C665 FILLER_0_4_91/a_484_472# _160_ 0.009925f
C666 _028_ net14 0.066292f
C667 net50 _030_ 0.073046f
C668 _242_/a_36_160# net37 0.02401f
C669 net47 _385_/a_36_68# 0.011168f
C670 trimb[3] trimb[2] 0.369908f
C671 _443_/a_36_151# _152_ 0.002345f
C672 FILLER_0_4_152/a_36_472# net57 0.015332f
C673 _440_/a_1000_472# vss 0.031704f
C674 FILLER_0_14_99/a_124_375# FILLER_0_13_100/a_36_472# 0.001597f
C675 net18 _418_/a_796_472# 0.003044f
C676 _070_ _118_ 0.302298f
C677 _340_/a_36_160# vdd 0.006001f
C678 _423_/a_36_151# net17 0.002865f
C679 _006_ result[3] 0.016909f
C680 _049_ FILLER_0_22_128/a_3172_472# 0.01125f
C681 _068_ net59 0.001388f
C682 _392_/a_36_68# cal_count\[3\] 0.003072f
C683 net16 net72 0.367221f
C684 _028_ _164_ 0.019799f
C685 output21/a_224_472# ctlp[4] 0.052556f
C686 net82 _443_/a_796_472# 0.00219f
C687 _127_ calibrate 0.004656f
C688 FILLER_0_21_28/a_1380_472# _012_ 0.004453f
C689 net72 _176_ 0.059793f
C690 net75 net4 0.031823f
C691 FILLER_0_21_286/a_484_472# net18 0.001956f
C692 _431_/a_36_151# FILLER_0_17_133/a_124_375# 0.059049f
C693 _017_ FILLER_0_14_107/a_1020_375# 0.001363f
C694 net70 FILLER_0_14_107/a_36_472# 0.054561f
C695 net44 FILLER_0_20_2/a_36_472# 0.037627f
C696 fanout79/a_36_160# vss 0.002268f
C697 net41 FILLER_0_21_28/a_932_472# 0.014034f
C698 output32/a_224_472# output34/a_224_472# 0.001691f
C699 FILLER_0_5_54/a_1380_472# trim_mask\[1\] 0.01205f
C700 net60 _102_ 0.008212f
C701 _414_/a_1308_423# vdd 0.004897f
C702 FILLER_0_1_266/a_572_375# net18 0.080358f
C703 _438_/a_448_472# vss 0.00615f
C704 _432_/a_2560_156# net80 0.01523f
C705 FILLER_0_0_96/a_124_375# vdd 0.034959f
C706 ctlp[1] _419_/a_1000_472# 0.005263f
C707 net15 _098_ 0.003965f
C708 net52 FILLER_0_5_72/a_124_375# 0.029702f
C709 _086_ _090_ 0.065807f
C710 FILLER_0_16_73/a_36_472# net15 0.005297f
C711 _093_ FILLER_0_17_161/a_124_375# 0.002431f
C712 FILLER_0_12_2/a_572_375# net3 0.001872f
C713 _451_/a_2225_156# vss 0.003848f
C714 _369_/a_36_68# _160_ 0.015312f
C715 _414_/a_36_151# _074_ 0.070632f
C716 FILLER_0_5_72/a_124_375# net49 0.001158f
C717 _415_/a_36_151# net19 0.05689f
C718 FILLER_0_4_152/a_124_375# _066_ 0.003354f
C719 FILLER_0_9_28/a_1020_375# FILLER_0_10_37/a_36_472# 0.001597f
C720 net38 net43 0.016358f
C721 FILLER_0_15_2/a_124_375# vdd 0.010829f
C722 ctln[2] cal 0.009784f
C723 trim_val\[1\] FILLER_0_6_37/a_36_472# 0.011347f
C724 _077_ cal_count\[3\] 0.176576f
C725 FILLER_0_17_56/a_124_375# FILLER_0_18_53/a_484_472# 0.001597f
C726 _074_ FILLER_0_7_233/a_36_472# 0.001341f
C727 net57 _069_ 0.026933f
C728 cal_itt\[2\] _253_/a_244_68# 0.001073f
C729 _088_ FILLER_0_5_198/a_572_375# 0.001374f
C730 _079_ FILLER_0_5_198/a_36_472# 0.012251f
C731 FILLER_0_19_28/a_572_375# net40 0.00139f
C732 FILLER_0_18_2/a_2364_375# output44/a_224_472# 0.032639f
C733 net68 FILLER_0_5_54/a_572_375# 0.040374f
C734 FILLER_0_5_109/a_572_375# vdd 0.024724f
C735 _077_ _059_ 0.020736f
C736 net15 FILLER_0_7_59/a_124_375# 0.004662f
C737 _096_ _055_ 0.047639f
C738 mask\[4\] FILLER_0_18_177/a_2812_375# 0.013557f
C739 _068_ _122_ 0.096251f
C740 net51 cal_count\[0\] 0.030963f
C741 _126_ FILLER_0_13_206/a_36_472# 0.026561f
C742 _328_/a_36_113# cal_count\[3\] 0.006392f
C743 trim[0] FILLER_0_3_2/a_36_472# 0.017429f
C744 FILLER_0_20_177/a_572_375# mask\[6\] 0.001158f
C745 FILLER_0_6_177/a_124_375# vss 0.002362f
C746 _073_ _070_ 0.001892f
C747 FILLER_0_6_177/a_572_375# vdd 0.02743f
C748 _074_ _163_ 0.446493f
C749 net36 FILLER_0_15_235/a_572_375# 0.083299f
C750 FILLER_0_4_152/a_124_375# net23 0.039975f
C751 _153_ _156_ 0.539362f
C752 _070_ _330_/a_224_472# 0.001096f
C753 _408_/a_718_524# net17 0.012884f
C754 _068_ _227_/a_36_160# 0.053563f
C755 _348_/a_49_472# vdd 0.038046f
C756 _417_/a_1308_423# _006_ 0.022704f
C757 FILLER_0_7_104/a_1020_375# _131_ 0.016404f
C758 _301_/a_36_472# vdd 0.013061f
C759 _438_/a_36_151# _437_/a_36_151# 0.002668f
C760 FILLER_0_18_2/a_1468_375# _452_/a_448_472# 0.001597f
C761 result[5] result[6] 0.065361f
C762 cal ctln[1] 0.123834f
C763 mask\[5\] _434_/a_2248_156# 0.003462f
C764 _052_ FILLER_0_21_28/a_3260_375# 0.002388f
C765 FILLER_0_9_28/a_2364_375# trim_val\[0\] 0.006639f
C766 _144_ _140_ 0.415736f
C767 net36 vdd 0.939735f
C768 _128_ net22 0.03249f
C769 net32 net18 0.028135f
C770 _076_ _163_ 0.030003f
C771 FILLER_0_18_37/a_932_472# vdd 0.01019f
C772 _086_ _321_/a_2034_472# 0.001815f
C773 net81 _098_ 0.029506f
C774 _429_/a_1000_472# vss 0.006901f
C775 output32/a_224_472# _418_/a_36_151# 0.07368f
C776 _093_ FILLER_0_16_89/a_36_472# 0.001338f
C777 net50 trim_mask\[3\] 0.001654f
C778 net39 FILLER_0_8_2/a_36_472# 0.010296f
C779 net74 _332_/a_36_472# 0.003752f
C780 net62 net19 0.352148f
C781 _092_ vss 0.346097f
C782 FILLER_0_16_107/a_484_472# vdd 0.02929f
C783 _096_ _126_ 0.258912f
C784 _053_ net47 0.011652f
C785 FILLER_0_9_72/a_36_472# _453_/a_2665_112# 0.001167f
C786 cal_count\[3\] _120_ 4.687877f
C787 cal_count\[3\] _038_ 0.682941f
C788 net20 net36 0.03843f
C789 net79 _416_/a_1308_423# 0.030119f
C790 _044_ net30 0.005104f
C791 mask\[4\] _137_ 0.086066f
C792 _059_ _120_ 0.0127f
C793 _415_/a_1308_423# FILLER_0_9_270/a_124_375# 0.001064f
C794 _193_/a_36_160# vdd 0.092266f
C795 _093_ FILLER_0_17_72/a_2724_472# 0.02416f
C796 _061_ _311_/a_3740_473# 0.006728f
C797 net70 vss 0.175272f
C798 net26 _424_/a_448_472# 0.063966f
C799 _142_ _137_ 1.401722f
C800 _431_/a_1204_472# _136_ 0.007382f
C801 FILLER_0_3_204/a_36_472# FILLER_0_3_212/a_36_472# 0.002296f
C802 _390_/a_36_68# _171_ 0.001252f
C803 _430_/a_2248_156# net36 0.001198f
C804 _140_ net23 0.06742f
C805 _086_ _318_/a_224_472# 0.007024f
C806 FILLER_0_10_247/a_124_375# vss 0.006235f
C807 FILLER_0_10_247/a_36_472# vdd 0.111658f
C808 _177_ _095_ 0.004392f
C809 input4/a_36_68# net5 0.004765f
C810 result[7] _419_/a_36_151# 0.001036f
C811 output44/a_224_472# vss 0.014054f
C812 mask\[5\] _202_/a_36_160# 0.00164f
C813 FILLER_0_9_105/a_484_472# FILLER_0_10_107/a_124_375# 0.001543f
C814 _412_/a_36_151# net19 0.03393f
C815 FILLER_0_21_206/a_124_375# net33 0.001579f
C816 _086_ _314_/a_224_472# 0.003715f
C817 vss FILLER_0_22_107/a_484_472# 0.003617f
C818 FILLER_0_22_86/a_572_375# net71 0.002239f
C819 output44/a_224_472# FILLER_0_20_15/a_932_472# 0.0323f
C820 FILLER_0_5_72/a_1020_375# _164_ 0.018398f
C821 FILLER_0_10_107/a_124_375# vss 0.003015f
C822 FILLER_0_10_107/a_572_375# vdd 0.043678f
C823 _327_/a_36_472# _127_ 0.002934f
C824 FILLER_0_15_228/a_124_375# vss 0.006435f
C825 FILLER_0_15_228/a_36_472# vdd 0.084606f
C826 FILLER_0_12_50/a_36_472# _067_ 0.011087f
C827 _452_/a_36_151# vdd 0.109842f
C828 net15 net55 1.200864f
C829 net55 FILLER_0_11_78/a_36_472# 0.059367f
C830 net67 FILLER_0_12_20/a_124_375# 0.007044f
C831 FILLER_0_6_239/a_36_472# _316_/a_124_24# 0.002228f
C832 _413_/a_2665_112# cal_itt\[2\] 0.003007f
C833 FILLER_0_4_197/a_932_472# net76 0.003693f
C834 net16 FILLER_0_17_38/a_484_472# 0.032356f
C835 net72 _041_ 0.467856f
C836 FILLER_0_5_164/a_484_472# _163_ 0.029894f
C837 _016_ _043_ 0.030341f
C838 net32 _048_ 0.008647f
C839 en vdd 0.282941f
C840 net61 _009_ 0.042703f
C841 FILLER_0_2_93/a_484_472# net69 0.0127f
C842 _414_/a_36_151# _081_ 0.016708f
C843 net20 FILLER_0_15_228/a_36_472# 0.020589f
C844 FILLER_0_12_124/a_124_375# vdd -0.00168f
C845 _425_/a_1204_472# calibrate 0.009749f
C846 output34/a_224_472# _094_ 0.002719f
C847 FILLER_0_9_142/a_36_472# vdd 0.107619f
C848 FILLER_0_9_142/a_124_375# vss 0.006851f
C849 FILLER_0_5_128/a_484_472# _081_ 0.00169f
C850 _072_ _311_/a_3740_473# 0.005483f
C851 FILLER_0_4_197/a_1468_375# vss 0.057762f
C852 _053_ net74 0.09773f
C853 _424_/a_2560_156# _012_ 0.002513f
C854 net38 FILLER_0_15_10/a_36_472# 0.020589f
C855 _378_/a_224_472# net67 0.00211f
C856 cal_itt\[2\] FILLER_0_3_221/a_932_472# 0.016327f
C857 FILLER_0_12_136/a_932_472# net23 0.004375f
C858 _086_ _414_/a_36_151# 0.002687f
C859 FILLER_0_9_28/a_124_375# net47 0.006757f
C860 _417_/a_2248_156# vdd 0.004032f
C861 net57 _385_/a_244_472# 0.001506f
C862 net19 _316_/a_848_380# 0.00558f
C863 _024_ _435_/a_796_472# 0.006511f
C864 FILLER_0_9_72/a_1020_375# vdd -0.014642f
C865 FILLER_0_9_72/a_572_375# vss 0.007993f
C866 mask\[5\] FILLER_0_20_193/a_124_375# 0.015793f
C867 net73 FILLER_0_19_111/a_36_472# 0.001412f
C868 _093_ FILLER_0_18_139/a_1020_375# 0.003529f
C869 _115_ _176_ 1.300336f
C870 cal_itt\[2\] _088_ 0.010847f
C871 _128_ vdd 0.217501f
C872 input1/a_36_113# vdd 0.099655f
C873 _073_ _082_ 0.009987f
C874 _421_/a_2248_156# _419_/a_2248_156# 0.001364f
C875 _081_ _163_ 0.427672f
C876 _085_ _310_/a_49_472# 0.001093f
C877 _002_ _270_/a_244_68# 0.001153f
C878 _073_ net82 0.028504f
C879 _119_ _313_/a_255_603# 0.001151f
C880 net35 FILLER_0_22_86/a_1380_472# 0.00813f
C881 FILLER_0_5_72/a_36_472# net47 0.003953f
C882 FILLER_0_7_72/a_2364_375# vdd 0.018287f
C883 FILLER_0_21_28/a_1020_375# net17 0.001134f
C884 cal fanout58/a_36_160# 0.047586f
C885 FILLER_0_13_65/a_36_472# net74 0.014937f
C886 FILLER_0_13_212/a_1380_472# _043_ 0.014431f
C887 _127_ FILLER_0_11_142/a_124_375# 0.00205f
C888 cal_count\[2\] FILLER_0_15_2/a_572_375# 0.015401f
C889 _015_ _426_/a_796_472# 0.007696f
C890 _053_ _372_/a_2034_472# 0.00181f
C891 mask\[4\] FILLER_0_17_200/a_484_472# 0.001701f
C892 _086_ _163_ 0.413768f
C893 state\[2\] cal_count\[3\] 0.005312f
C894 net52 FILLER_0_2_101/a_124_375# 0.007787f
C895 net55 net51 0.007067f
C896 net20 _128_ 0.041f
C897 FILLER_0_16_89/a_36_472# _136_ 0.00722f
C898 ctln[1] FILLER_0_3_221/a_1468_375# 0.001235f
C899 _028_ _153_ 0.008011f
C900 net46 output44/a_224_472# 0.003211f
C901 FILLER_0_18_177/a_2724_472# net22 0.004297f
C902 _000_ FILLER_0_3_221/a_1380_472# 0.025567f
C903 net47 _166_ 0.034342f
C904 _337_/a_257_69# _137_ 0.001822f
C905 FILLER_0_18_2/a_1380_472# net55 0.007469f
C906 _430_/a_796_472# net63 0.002914f
C907 net65 _163_ 0.013462f
C908 _098_ _437_/a_1204_472# 0.005729f
C909 net58 FILLER_0_8_263/a_124_375# 0.001876f
C910 mask\[8\] _213_/a_67_603# 0.039626f
C911 net54 FILLER_0_22_128/a_932_472# 0.014735f
C912 _115_ _124_ 0.045023f
C913 mask\[5\] FILLER_0_18_177/a_1020_375# 0.001604f
C914 FILLER_0_14_91/a_484_472# FILLER_0_14_99/a_36_472# 0.013276f
C915 FILLER_0_17_72/a_2724_472# _136_ 0.03065f
C916 FILLER_0_4_185/a_124_375# net76 0.053929f
C917 _131_ FILLER_0_16_115/a_36_472# 0.008241f
C918 vss _433_/a_448_472# 0.005349f
C919 mask\[0\] _429_/a_1308_423# 0.019225f
C920 _093_ FILLER_0_18_76/a_484_472# 0.024853f
C921 _132_ net71 0.099427f
C922 _027_ _438_/a_448_472# 0.053901f
C923 net4 net19 0.050898f
C924 FILLER_0_3_172/a_572_375# net22 0.013048f
C925 FILLER_0_20_98/a_36_472# _437_/a_36_151# 0.001723f
C926 _094_ _418_/a_36_151# 0.041823f
C927 _394_/a_1336_472# FILLER_0_15_72/a_124_375# 0.016876f
C928 _052_ _424_/a_1000_472# 0.007574f
C929 _185_ net47 0.185634f
C930 FILLER_0_16_57/a_572_375# _131_ 0.015859f
C931 cal_itt\[2\] cal_itt\[0\] 0.011453f
C932 net39 net17 0.099429f
C933 FILLER_0_8_263/a_124_375# calibrate 0.006928f
C934 FILLER_0_11_142/a_36_472# _076_ 0.003047f
C935 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_124_375# 0.012001f
C936 _395_/a_1044_488# _085_ 0.00391f
C937 _395_/a_36_488# _176_ 0.010116f
C938 _053_ _154_ 0.41707f
C939 net17 net51 0.026974f
C940 net72 FILLER_0_17_64/a_124_375# 0.002236f
C941 FILLER_0_7_162/a_36_472# _074_ 0.003809f
C942 _096_ state\[1\] 0.083332f
C943 _131_ _183_ 0.227229f
C944 net23 FILLER_0_21_150/a_36_472# 0.016375f
C945 result[6] net19 0.834308f
C946 FILLER_0_19_195/a_36_472# vss 0.005146f
C947 FILLER_0_7_104/a_1468_375# _133_ 0.003206f
C948 trim[1] _033_ 0.015549f
C949 FILLER_0_18_2/a_1380_472# net17 0.003603f
C950 net15 _216_/a_67_603# 0.060076f
C951 output27/a_224_472# vdd 0.070751f
C952 _411_/a_1204_472# net8 0.001768f
C953 FILLER_0_20_177/a_124_375# vdd 0.001964f
C954 fanout52/a_36_160# _443_/a_2665_112# 0.007884f
C955 FILLER_0_4_152/a_124_375# net57 0.001947f
C956 fanout72/a_36_113# _043_ 0.017862f
C957 net81 _425_/a_448_472# 0.056225f
C958 FILLER_0_14_181/a_36_472# _098_ 0.004669f
C959 FILLER_0_5_206/a_36_472# _081_ 0.014328f
C960 _104_ result[7] 0.475003f
C961 ctlp[3] _422_/a_36_151# 0.002627f
C962 _093_ FILLER_0_18_209/a_36_472# 0.007068f
C963 _414_/a_2560_156# net22 0.00603f
C964 output16/a_224_472# _447_/a_448_472# 0.003175f
C965 trim_val\[0\] FILLER_0_6_47/a_484_472# 0.001215f
C966 _086_ _117_ 0.010287f
C967 net15 _111_ 0.049514f
C968 _365_/a_36_68# vss 0.029516f
C969 FILLER_0_16_89/a_932_472# net36 0.001709f
C970 FILLER_0_24_63/a_36_472# output25/a_224_472# 0.002338f
C971 FILLER_0_21_142/a_124_375# FILLER_0_22_128/a_1828_472# 0.001543f
C972 net81 _082_ 0.001633f
C973 _413_/a_36_151# FILLER_0_3_172/a_3172_472# 0.001723f
C974 _035_ _445_/a_36_151# 0.002276f
C975 _429_/a_36_151# FILLER_0_15_212/a_1020_375# 0.035849f
C976 net81 net82 0.063498f
C977 FILLER_0_20_15/a_124_375# vdd 0.006513f
C978 _057_ _161_ 1.09228f
C979 net65 FILLER_0_1_266/a_572_375# 0.002969f
C980 mask\[7\] _297_/a_36_472# 0.003196f
C981 _104_ _198_/a_67_603# 0.007168f
C982 _095_ _451_/a_2225_156# 0.001102f
C983 _181_ _179_ 0.011848f
C984 _114_ net23 0.029535f
C985 _141_ FILLER_0_21_150/a_124_375# 0.02192f
C986 cal_count\[2\] _452_/a_448_472# 0.003314f
C987 _062_ _310_/a_49_472# 0.020509f
C988 ctlp[2] _109_ 0.059999f
C989 FILLER_0_17_38/a_484_472# _041_ 0.009607f
C990 _028_ FILLER_0_7_72/a_2724_472# 0.001777f
C991 net74 FILLER_0_11_124/a_36_472# 0.020589f
C992 _441_/a_36_151# vdd 0.098562f
C993 _415_/a_36_151# output28/a_224_472# 0.229574f
C994 _092_ _275_/a_224_472# 0.002138f
C995 net69 _369_/a_244_472# 0.002456f
C996 _060_ net21 0.074356f
C997 net78 _418_/a_36_151# 0.003648f
C998 FILLER_0_16_89/a_36_472# net53 0.004701f
C999 _058_ FILLER_0_9_105/a_124_375# 0.014234f
C1000 mask\[3\] net30 0.451388f
C1001 net27 net37 0.003648f
C1002 FILLER_0_18_177/a_2724_472# vdd 0.002749f
C1003 net52 _442_/a_2248_156# 0.022954f
C1004 _005_ _416_/a_1000_472# 0.027013f
C1005 FILLER_0_24_130/a_124_375# net54 0.001269f
C1006 _053_ _079_ 0.007118f
C1007 FILLER_0_2_101/a_36_472# trim_mask\[3\] 0.013363f
C1008 result[9] _419_/a_1204_472# 0.019627f
C1009 net56 FILLER_0_16_154/a_932_472# 0.001401f
C1010 _441_/a_1308_423# _168_ 0.044302f
C1011 valid fanout64/a_36_160# 0.001811f
C1012 FILLER_0_9_60/a_484_472# vdd 0.005181f
C1013 FILLER_0_9_60/a_36_472# vss 0.001327f
C1014 _140_ FILLER_0_19_155/a_484_472# 0.004155f
C1015 net18 _419_/a_2560_156# 0.008155f
C1016 fanout75/a_36_113# net37 0.010418f
C1017 ctlp[1] _421_/a_1308_423# 0.002417f
C1018 FILLER_0_21_206/a_36_472# mask\[6\] 0.015735f
C1019 vdd _295_/a_36_472# 0.0083f
C1020 _114_ FILLER_0_11_109/a_124_375# 0.009676f
C1021 FILLER_0_17_104/a_932_472# net14 0.002113f
C1022 _429_/a_2248_156# _043_ 0.001001f
C1023 _069_ net36 0.032818f
C1024 FILLER_0_3_172/a_572_375# vdd 0.007121f
C1025 _100_ mask\[1\] 0.002229f
C1026 FILLER_0_17_218/a_484_472# vdd 0.004777f
C1027 FILLER_0_17_218/a_36_472# vss 0.006061f
C1028 net48 _074_ 1.192591f
C1029 _425_/a_2560_156# vdd 0.001827f
C1030 _425_/a_2665_112# vss 0.002983f
C1031 mask\[7\] FILLER_0_22_128/a_2724_472# 0.001055f
C1032 net63 FILLER_0_20_177/a_1020_375# 0.005919f
C1033 _069_ _429_/a_1204_472# 0.025254f
C1034 _443_/a_2248_156# net22 0.001984f
C1035 result[6] _420_/a_36_151# 0.011901f
C1036 _432_/a_36_151# FILLER_0_17_161/a_36_472# 0.004847f
C1037 mask\[2\] FILLER_0_15_180/a_484_472# 0.00848f
C1038 FILLER_0_20_31/a_124_375# FILLER_0_20_15/a_1468_375# 0.012001f
C1039 _116_ calibrate 0.018482f
C1040 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1468_375# 0.086742f
C1041 FILLER_0_14_181/a_36_472# FILLER_0_15_180/a_124_375# 0.001723f
C1042 state\[2\] _427_/a_2665_112# 0.007007f
C1043 _012_ _098_ 0.002778f
C1044 _013_ FILLER_0_18_61/a_36_472# 0.01628f
C1045 net48 _076_ 0.077031f
C1046 _423_/a_36_151# FILLER_0_23_44/a_1468_375# 0.059049f
C1047 fanout62/a_36_160# result[1] 0.036633f
C1048 net62 output28/a_224_472# 0.206137f
C1049 FILLER_0_5_72/a_124_375# FILLER_0_5_54/a_1468_375# 0.005439f
C1050 _017_ _043_ 0.02569f
C1051 cal net18 0.123815f
C1052 net26 _217_/a_36_160# 0.021067f
C1053 _098_ FILLER_0_15_212/a_36_472# 0.011079f
C1054 _428_/a_2665_112# net74 0.048822f
C1055 _429_/a_36_151# FILLER_0_15_205/a_36_472# 0.001723f
C1056 net50 _439_/a_2560_156# 0.006321f
C1057 _323_/a_36_113# _223_/a_36_160# 0.238626f
C1058 vdd _416_/a_36_151# 0.142481f
C1059 FILLER_0_4_144/a_484_472# net23 0.01239f
C1060 mask\[4\] output34/a_224_472# 0.001777f
C1061 _029_ _163_ 0.007545f
C1062 _256_/a_2960_68# _076_ 0.001292f
C1063 _422_/a_36_151# _108_ 0.062205f
C1064 _116_ net21 0.036746f
C1065 _086_ FILLER_0_11_142/a_36_472# 0.006774f
C1066 _415_/a_2248_156# net64 0.051575f
C1067 result[2] FILLER_0_15_282/a_124_375# 0.001114f
C1068 trim[0] trim[2] 0.002289f
C1069 net16 _167_ 0.001124f
C1070 FILLER_0_3_204/a_36_472# net22 0.036788f
C1071 _422_/a_36_151# net19 0.033614f
C1072 FILLER_0_7_162/a_36_472# _081_ 0.002493f
C1073 output46/a_224_472# FILLER_0_20_15/a_572_375# 0.00135f
C1074 _261_/a_36_160# vss 0.05095f
C1075 net70 _095_ 0.222423f
C1076 _028_ FILLER_0_6_47/a_2724_472# 0.023218f
C1077 _086_ FILLER_0_7_104/a_1020_375# 0.00757f
C1078 _098_ _434_/a_1308_423# 0.007057f
C1079 _210_/a_67_603# mask\[7\] 0.039004f
C1080 _117_ _090_ 0.041465f
C1081 FILLER_0_22_86/a_1380_472# vdd 0.008224f
C1082 FILLER_0_22_86/a_932_472# vss -0.001553f
C1083 net16 _235_/a_67_603# 0.038585f
C1084 _199_/a_36_160# vss 0.004608f
C1085 mask\[4\] FILLER_0_19_171/a_484_472# 0.004669f
C1086 output13/a_224_472# _387_/a_36_113# 0.020974f
C1087 en_co_clk _172_ 0.025699f
C1088 net31 net36 0.00943f
C1089 _415_/a_1308_423# vdd 0.004258f
C1090 mask\[4\] FILLER_0_18_171/a_124_375# 0.008445f
C1091 result[5] _419_/a_36_151# 0.006539f
C1092 net2 _082_ 0.034094f
C1093 FILLER_0_9_223/a_36_472# vdd 0.030289f
C1094 _118_ net21 0.007371f
C1095 net82 net2 0.451147f
C1096 _061_ _055_ 0.853642f
C1097 _036_ _381_/a_36_472# 0.023012f
C1098 FILLER_0_7_146/a_124_375# net23 0.00129f
C1099 FILLER_0_13_65/a_124_375# fanout72/a_36_113# 0.005467f
C1100 _030_ FILLER_0_3_78/a_124_375# 0.010439f
C1101 _055_ _311_/a_66_473# 0.040326f
C1102 _070_ net47 0.071795f
C1103 _069_ FILLER_0_9_142/a_36_472# 0.035528f
C1104 _320_/a_224_472# vdd 0.001757f
C1105 _053_ FILLER_0_6_47/a_1828_472# 0.006408f
C1106 FILLER_0_0_198/a_36_472# net11 0.056269f
C1107 FILLER_0_16_73/a_124_375# net55 0.007695f
C1108 net52 FILLER_0_6_79/a_36_472# 0.012286f
C1109 net28 net36 0.002537f
C1110 net82 FILLER_0_3_172/a_2276_472# 0.007729f
C1111 FILLER_0_21_206/a_124_375# net22 0.05301f
C1112 _105_ _297_/a_36_472# 0.03208f
C1113 _411_/a_36_151# ctln[4] 0.0022f
C1114 net58 _073_ 0.057725f
C1115 net34 FILLER_0_22_128/a_2364_375# 0.009656f
C1116 _093_ FILLER_0_18_107/a_2724_472# 0.00308f
C1117 _405_/a_67_603# vdd 0.034681f
C1118 vdd FILLER_0_14_235/a_484_472# 0.010228f
C1119 vss FILLER_0_14_235/a_36_472# 0.001602f
C1120 FILLER_0_4_197/a_124_375# _079_ 0.004772f
C1121 net27 FILLER_0_9_282/a_572_375# 0.002809f
C1122 _442_/a_2665_112# trim_mask\[3\] 0.019514f
C1123 _173_ cal_count\[0\] 0.517178f
C1124 _292_/a_36_160# net22 0.001864f
C1125 _128_ _069_ 0.018491f
C1126 _057_ _056_ 0.167928f
C1127 FILLER_0_4_152/a_124_375# FILLER_0_5_148/a_572_375# 0.05841f
C1128 calibrate _123_ 0.016296f
C1129 net61 net33 0.043271f
C1130 _443_/a_1204_472# vss 0.005425f
C1131 _443_/a_2248_156# vdd 0.010579f
C1132 FILLER_0_22_86/a_484_472# _437_/a_36_151# 0.013806f
C1133 fanout54/a_36_160# net54 0.018583f
C1134 FILLER_0_14_99/a_124_375# _451_/a_1040_527# 0.010005f
C1135 _255_/a_224_552# _311_/a_66_473# 0.002588f
C1136 _009_ FILLER_0_23_274/a_36_472# 0.005531f
C1137 FILLER_0_5_164/a_124_375# _066_ 0.006762f
C1138 FILLER_0_5_128/a_124_375# _160_ 0.001157f
C1139 ctln[2] net8 0.057281f
C1140 _072_ _055_ 0.083351f
C1141 _446_/a_448_472# net66 0.017696f
C1142 FILLER_0_24_130/a_36_472# output24/a_224_472# 0.023414f
C1143 net48 _081_ 0.137029f
C1144 _429_/a_36_151# FILLER_0_13_206/a_124_375# 0.001597f
C1145 _414_/a_36_151# _163_ 0.001186f
C1146 result[7] net60 0.778099f
C1147 net55 net47 0.049398f
C1148 _000_ _411_/a_36_151# 0.023297f
C1149 _449_/a_2248_156# FILLER_0_13_80/a_124_375# 0.001068f
C1150 FILLER_0_24_130/a_36_472# vss 0.001687f
C1151 FILLER_0_5_128/a_484_472# _163_ 0.009861f
C1152 _033_ _164_ 0.007117f
C1153 FILLER_0_16_57/a_1468_375# net55 0.006307f
C1154 FILLER_0_16_57/a_932_472# net72 0.004262f
C1155 _425_/a_36_151# FILLER_0_8_247/a_484_472# 0.059367f
C1156 _423_/a_1308_423# vss 0.001726f
C1157 _423_/a_796_472# vdd 0.001494f
C1158 sample net18 0.103617f
C1159 FILLER_0_16_89/a_572_375# vdd 0.005006f
C1160 _032_ net69 0.347645f
C1161 FILLER_0_3_204/a_36_472# vdd 0.092654f
C1162 valid net82 0.060784f
C1163 cal_count\[3\] _389_/a_428_148# 0.001072f
C1164 net57 _428_/a_2248_156# 0.022587f
C1165 mask\[0\] _100_ 0.005921f
C1166 net55 _012_ 0.060122f
C1167 net74 _070_ 0.394108f
C1168 _016_ FILLER_0_12_136/a_484_472# 0.001516f
C1169 _057_ _068_ 0.393271f
C1170 _126_ FILLER_0_11_101/a_484_472# 0.001488f
C1171 ctln[1] net8 0.678616f
C1172 net56 FILLER_0_19_155/a_124_375# 0.006762f
C1173 _077_ net52 0.047585f
C1174 FILLER_0_15_72/a_572_375# cal_count\[1\] 0.135344f
C1175 _142_ _334_/a_36_160# 0.009001f
C1176 _114_ net57 0.22998f
C1177 FILLER_0_9_28/a_2364_375# _453_/a_36_151# 0.001597f
C1178 FILLER_0_17_72/a_1380_472# vdd 0.001762f
C1179 FILLER_0_17_72/a_932_472# vss 0.002754f
C1180 _072_ _126_ 0.012566f
C1181 _214_/a_36_160# _437_/a_36_151# 0.001542f
C1182 FILLER_0_5_136/a_124_375# vss 0.053395f
C1183 FILLER_0_5_136/a_36_472# vdd 0.092379f
C1184 _430_/a_36_151# net80 0.082603f
C1185 FILLER_0_16_107/a_124_375# FILLER_0_18_107/a_36_472# 0.001512f
C1186 FILLER_0_4_107/a_484_472# _369_/a_36_68# 0.001049f
C1187 FILLER_0_12_20/a_572_375# _039_ 0.005679f
C1188 FILLER_0_7_195/a_36_472# _062_ 0.0045f
C1189 _119_ _319_/a_672_472# 0.00488f
C1190 net17 net47 2.009509f
C1191 ctln[5] _448_/a_36_151# 0.009209f
C1192 FILLER_0_3_78/a_572_375# _164_ 0.055492f
C1193 _427_/a_2248_156# vdd -0.002315f
C1194 _427_/a_1204_472# vss 0.0041f
C1195 _032_ _152_ 0.001206f
C1196 trim_mask\[4\] _370_/a_1084_68# 0.005157f
C1197 trim_val\[1\] net47 0.34878f
C1198 _415_/a_2560_156# vss 0.001286f
C1199 FILLER_0_5_172/a_124_375# FILLER_0_5_164/a_572_375# 0.012001f
C1200 _028_ _376_/a_36_160# 0.026437f
C1201 _372_/a_170_472# _133_ 0.031518f
C1202 cal_count\[3\] cal_count\[2\] 0.005307f
C1203 _340_/a_36_160# _140_ 0.062613f
C1204 net16 vdd 2.255325f
C1205 net58 net81 0.375649f
C1206 net76 FILLER_0_3_172/a_1020_375# 0.007439f
C1207 _085_ vss 0.132721f
C1208 FILLER_0_12_220/a_932_472# _070_ 0.001282f
C1209 _176_ vdd 0.874707f
C1210 ctlp[1] _098_ 0.0012f
C1211 _091_ FILLER_0_15_212/a_1380_472# 0.002787f
C1212 net50 _440_/a_2665_112# 0.009767f
C1213 FILLER_0_5_212/a_124_375# net59 0.045135f
C1214 FILLER_0_21_206/a_124_375# vdd 0.038521f
C1215 mask\[4\] FILLER_0_20_177/a_1380_472# 0.001215f
C1216 mask\[3\] FILLER_0_18_177/a_36_472# 0.005668f
C1217 net82 trim_mask\[4\] 0.21475f
C1218 FILLER_0_8_24/a_36_472# net42 0.010665f
C1219 net55 net74 0.048927f
C1220 _137_ net23 0.031218f
C1221 _144_ _049_ 0.100508f
C1222 net15 trim_mask\[2\] 0.026132f
C1223 _077_ FILLER_0_8_239/a_124_375# 0.001772f
C1224 _100_ _099_ 0.03589f
C1225 net52 _120_ 0.023363f
C1226 net52 _038_ 0.001152f
C1227 fanout57/a_36_113# trim_mask\[4\] 0.002404f
C1228 _292_/a_36_160# vdd 0.01694f
C1229 trim[1] _444_/a_36_151# 0.001391f
C1230 mask\[7\] _109_ 0.028117f
C1231 FILLER_0_18_107/a_2812_375# _145_ 0.030158f
C1232 net15 FILLER_0_23_44/a_1468_375# 0.001307f
C1233 trim_val\[0\] _453_/a_36_151# 0.001629f
C1234 net81 calibrate 0.047274f
C1235 FILLER_0_18_171/a_36_472# _141_ 0.002037f
C1236 _077_ FILLER_0_9_223/a_124_375# 0.008762f
C1237 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_36_472# 0.007947f
C1238 _447_/a_2560_156# vss 0.00126f
C1239 _053_ FILLER_0_6_177/a_124_375# 0.009352f
C1240 net81 FILLER_0_10_256/a_124_375# 0.026113f
C1241 FILLER_0_4_144/a_484_472# net57 0.003724f
C1242 mask\[5\] FILLER_0_19_171/a_572_375# 0.007169f
C1243 FILLER_0_16_57/a_1380_472# cal_count\[1\] 0.001568f
C1244 _124_ vdd 0.040228f
C1245 FILLER_0_11_64/a_124_375# _453_/a_2248_156# 0.001901f
C1246 net54 mask\[7\] 0.262465f
C1247 net81 net21 0.185411f
C1248 mask\[0\] FILLER_0_14_235/a_124_375# 0.009674f
C1249 _414_/a_2248_156# _074_ 0.013023f
C1250 net23 _049_ 0.215528f
C1251 _086_ _325_/a_224_472# 0.003155f
C1252 FILLER_0_9_72/a_124_375# _439_/a_36_151# 0.059049f
C1253 FILLER_0_5_72/a_1020_375# _440_/a_2248_156# 0.001068f
C1254 FILLER_0_7_72/a_3172_472# _219_/a_36_160# 0.035111f
C1255 net19 _419_/a_36_151# 0.009613f
C1256 net60 net79 0.113281f
C1257 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_484_472# 0.013277f
C1258 FILLER_0_5_212/a_124_375# _122_ 0.001352f
C1259 FILLER_0_12_28/a_124_375# _039_ 0.004669f
C1260 _405_/a_255_603# cal_count\[2\] 0.001576f
C1261 FILLER_0_18_100/a_36_472# net14 0.046864f
C1262 _432_/a_448_472# mask\[3\] 0.005831f
C1263 mask\[5\] _346_/a_49_472# 0.037629f
C1264 fanout71/a_36_113# vdd 0.028178f
C1265 _257_/a_36_472# vdd -0.001779f
C1266 _431_/a_36_151# FILLER_0_18_107/a_2724_472# 0.00271f
C1267 FILLER_0_5_117/a_36_472# _160_ 0.005314f
C1268 FILLER_0_2_111/a_1468_375# _160_ 0.001026f
C1269 net74 _370_/a_1084_68# 0.001301f
C1270 _214_/a_36_160# _051_ 0.207388f
C1271 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_572_375# 0.001597f
C1272 _216_/a_67_603# _012_ 0.001014f
C1273 _444_/a_2560_156# _054_ 0.003269f
C1274 _140_ _348_/a_49_472# 0.023816f
C1275 net75 _426_/a_1308_423# 0.002552f
C1276 net15 FILLER_0_18_61/a_124_375# 0.001179f
C1277 _061_ state\[1\] 0.02716f
C1278 net71 _437_/a_1308_423# 0.023981f
C1279 _074_ net37 0.064705f
C1280 FILLER_0_16_57/a_1468_375# _111_ 0.001371f
C1281 net36 _282_/a_36_160# 0.002754f
C1282 _435_/a_1308_423# vdd 0.012856f
C1283 net38 _444_/a_448_472# 0.031117f
C1284 mask\[0\] _060_ 0.002039f
C1285 net82 net74 0.007059f
C1286 FILLER_0_10_78/a_36_472# FILLER_0_9_72/a_572_375# 0.001543f
C1287 _019_ _098_ 0.010193f
C1288 trim_mask\[1\] FILLER_0_5_88/a_36_472# 0.038642f
C1289 net38 FILLER_0_8_24/a_124_375# 0.001013f
C1290 cal_count\[3\] _043_ 0.721078f
C1291 _103_ _418_/a_1000_472# 0.006239f
C1292 FILLER_0_3_204/a_124_375# _413_/a_36_151# 0.035849f
C1293 _449_/a_2665_112# net55 0.057694f
C1294 _076_ net37 0.072179f
C1295 FILLER_0_18_76/a_124_375# vdd 0.019258f
C1296 FILLER_0_16_73/a_572_375# vss 0.030752f
C1297 _414_/a_2665_112# _072_ 0.025361f
C1298 _134_ FILLER_0_9_105/a_124_375# 0.005919f
C1299 _253_/a_36_68# _082_ 0.013108f
C1300 _424_/a_2665_112# net36 0.028938f
C1301 net52 fanout52/a_36_160# 0.036543f
C1302 _253_/a_36_68# net82 0.016638f
C1303 _228_/a_36_68# net21 0.055313f
C1304 ctlp[3] _104_ 0.025066f
C1305 cal net65 0.023638f
C1306 net7 ctln[9] 0.005103f
C1307 net41 _446_/a_448_472# 0.040165f
C1308 _062_ vss 0.58133f
C1309 net69 _367_/a_36_68# 0.008893f
C1310 _088_ _083_ 0.007169f
C1311 net58 net2 0.070564f
C1312 _440_/a_3041_156# _164_ 0.001221f
C1313 net38 _452_/a_2225_156# 0.034415f
C1314 mask\[3\] _046_ 0.018595f
C1315 _438_/a_2560_156# net14 0.049389f
C1316 _072_ state\[1\] 0.267762f
C1317 fanout81/a_36_160# net81 0.025745f
C1318 _096_ FILLER_0_15_180/a_572_375# 0.001972f
C1319 output8/a_224_472# net4 0.015359f
C1320 ctln[8] vss 0.351742f
C1321 FILLER_0_21_28/a_2364_375# vdd -0.011393f
C1322 net82 _159_ 0.001393f
C1323 net2 calibrate 0.003482f
C1324 _041_ vdd 0.19154f
C1325 _104_ _422_/a_448_472# 0.001955f
C1326 FILLER_0_15_290/a_36_472# FILLER_0_15_282/a_484_472# 0.013277f
C1327 _430_/a_2665_112# net63 0.075661f
C1328 _265_/a_244_68# _084_ 0.016463f
C1329 net57 FILLER_0_5_164/a_124_375# 0.040872f
C1330 _148_ FILLER_0_22_128/a_36_472# 0.010386f
C1331 net63 _435_/a_1000_472# 0.002536f
C1332 _105_ _109_ 0.107328f
C1333 FILLER_0_24_96/a_36_472# net14 0.002882f
C1334 net36 _451_/a_36_151# 0.02414f
C1335 net54 _437_/a_448_472# 0.004418f
C1336 _093_ FILLER_0_17_104/a_484_472# 0.014431f
C1337 FILLER_0_5_212/a_124_375# FILLER_0_5_206/a_124_375# 0.005439f
C1338 FILLER_0_4_107/a_36_472# net47 0.002982f
C1339 _267_/a_36_472# vdd 0.005477f
C1340 FILLER_0_12_136/a_1020_375# state\[2\] 0.001952f
C1341 FILLER_0_5_164/a_484_472# net37 0.013857f
C1342 FILLER_0_16_255/a_36_472# net36 0.034335f
C1343 FILLER_0_18_209/a_36_472# _047_ 0.002672f
C1344 FILLER_0_6_90/a_484_472# vss 0.00243f
C1345 _091_ FILLER_0_18_177/a_572_375# 0.004285f
C1346 mask\[7\] _350_/a_49_472# 0.035293f
C1347 _414_/a_2248_156# _081_ 0.002027f
C1348 FILLER_0_16_107/a_484_472# _451_/a_36_151# 0.027244f
C1349 result[2] _005_ 0.060821f
C1350 mask\[5\] FILLER_0_20_177/a_1468_375# 0.013222f
C1351 _418_/a_2560_156# vdd 0.001506f
C1352 _418_/a_2665_112# vss 0.003519f
C1353 net82 FILLER_0_3_142/a_124_375# 0.018696f
C1354 FILLER_0_3_172/a_2276_472# net21 0.003603f
C1355 net14 FILLER_0_10_94/a_124_375# 0.007086f
C1356 _433_/a_1288_156# _022_ 0.001147f
C1357 _190_/a_36_160# _450_/a_36_151# 0.002486f
C1358 _132_ FILLER_0_19_111/a_484_472# 0.004619f
C1359 net52 FILLER_0_9_72/a_932_472# 0.008749f
C1360 _085_ _071_ 0.127349f
C1361 _131_ FILLER_0_18_37/a_1468_375# 0.001151f
C1362 FILLER_0_16_107/a_36_472# _131_ 0.008817f
C1363 net55 _177_ 0.327874f
C1364 net70 _451_/a_448_472# 0.043107f
C1365 FILLER_0_13_142/a_484_472# net23 0.006746f
C1366 _256_/a_3368_68# net22 0.001285f
C1367 trim[1] vss 0.085436f
C1368 net58 valid 0.149817f
C1369 output37/a_224_472# _425_/a_2665_112# 0.022027f
C1370 _057_ _113_ 0.339862f
C1371 _274_/a_36_68# net4 0.037848f
C1372 _104_ _108_ 0.02837f
C1373 result[7] FILLER_0_23_290/a_124_375# 0.018455f
C1374 _077_ FILLER_0_8_156/a_36_472# 0.00563f
C1375 FILLER_0_9_60/a_572_375# _439_/a_36_151# 0.001107f
C1376 _081_ net37 1.274337f
C1377 _415_/a_2665_112# _416_/a_36_151# 0.001602f
C1378 _104_ net19 0.159483f
C1379 _104_ net63 0.005363f
C1380 net81 mask\[1\] 2.509493f
C1381 net57 _137_ 0.006142f
C1382 _077_ _229_/a_224_472# 0.001293f
C1383 FILLER_0_18_2/a_2724_472# vdd 0.004348f
C1384 FILLER_0_18_2/a_2276_472# vss 0.001865f
C1385 FILLER_0_4_177/a_36_472# _386_/a_848_380# 0.007646f
C1386 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_36_472# 0.001963f
C1387 _086_ net37 0.039329f
C1388 FILLER_0_11_64/a_36_472# cal_count\[3\] 0.0081f
C1389 output27/a_224_472# FILLER_0_9_290/a_36_472# 0.001711f
C1390 valid calibrate 0.002363f
C1391 result[5] net60 0.16275f
C1392 fanout60/a_36_160# _418_/a_36_151# 0.029017f
C1393 output29/a_224_472# vdd 0.103437f
C1394 _011_ _299_/a_36_472# 0.004407f
C1395 sample net65 0.148853f
C1396 net82 FILLER_0_3_221/a_484_472# 0.013492f
C1397 net48 FILLER_0_7_233/a_36_472# 0.01015f
C1398 _426_/a_36_151# vdd 0.086652f
C1399 _098_ _438_/a_448_472# 0.008962f
C1400 net65 net37 0.008382f
C1401 ctlp[8] net35 0.001859f
C1402 net2 clk 0.046099f
C1403 FILLER_0_8_247/a_36_472# calibrate 0.008647f
C1404 FILLER_0_12_220/a_36_472# _090_ 0.023446f
C1405 FILLER_0_1_204/a_36_472# vss 0.002247f
C1406 _065_ _447_/a_796_472# 0.007495f
C1407 _079_ _082_ 0.709481f
C1408 net65 FILLER_0_3_221/a_1468_375# 0.001695f
C1409 _427_/a_2665_112# _043_ 0.002612f
C1410 _094_ _007_ 0.170362f
C1411 output36/a_224_472# result[9] 0.059164f
C1412 FILLER_0_12_20/a_484_472# FILLER_0_12_28/a_36_472# 0.013277f
C1413 _106_ mask\[1\] 0.005728f
C1414 FILLER_0_2_93/a_124_375# net14 0.007439f
C1415 net72 FILLER_0_17_38/a_124_375# 0.041464f
C1416 _175_ FILLER_0_15_72/a_572_375# 0.04785f
C1417 fanout66/a_36_113# _160_ 0.015681f
C1418 FILLER_0_12_20/a_484_472# net40 0.003391f
C1419 _341_/a_49_472# _142_ 0.011026f
C1420 output7/a_224_472# vss 0.00746f
C1421 mask\[3\] _143_ 0.023322f
C1422 _377_/a_36_472# trim_val\[0\] 0.135527f
C1423 FILLER_0_17_64/a_124_375# vdd 0.027957f
C1424 result[9] net30 0.231442f
C1425 net18 net8 0.072251f
C1426 net64 FILLER_0_8_247/a_1468_375# 0.002559f
C1427 FILLER_0_17_142/a_124_375# vss 0.008753f
C1428 FILLER_0_17_142/a_572_375# vdd 0.012885f
C1429 _053_ _365_/a_36_68# 0.001572f
C1430 _120_ FILLER_0_8_156/a_36_472# 0.005842f
C1431 fanout81/a_36_160# net2 0.044793f
C1432 FILLER_0_6_47/a_124_375# vdd 0.008011f
C1433 net38 net44 0.523774f
C1434 trim[0] vdd 0.125774f
C1435 mask\[5\] _108_ 0.036539f
C1436 _427_/a_1204_472# _095_ 0.006692f
C1437 _069_ _176_ 0.766885f
C1438 _288_/a_224_472# _102_ 0.002528f
C1439 FILLER_0_4_177/a_124_375# net22 0.006125f
C1440 output35/a_224_472# FILLER_0_21_206/a_36_472# 0.0323f
C1441 _193_/a_36_160# output30/a_224_472# 0.018f
C1442 _411_/a_448_472# net8 0.04545f
C1443 _446_/a_1000_472# trim[3] 0.001257f
C1444 mask\[5\] net63 0.112147f
C1445 FILLER_0_16_255/a_124_375# _417_/a_2665_112# 0.003856f
C1446 FILLER_0_4_197/a_484_472# net22 0.007955f
C1447 _091_ _093_ 0.035503f
C1448 _428_/a_1204_472# _017_ 0.005148f
C1449 FILLER_0_2_171/a_36_472# vss 0.002909f
C1450 FILLER_0_5_54/a_1380_472# FILLER_0_6_47/a_2276_472# 0.026657f
C1451 _412_/a_1308_423# net81 0.006961f
C1452 _161_ _056_ 0.065732f
C1453 _443_/a_36_151# _442_/a_36_151# 0.06169f
C1454 _050_ _436_/a_36_151# 0.037103f
C1455 FILLER_0_12_236/a_572_375# FILLER_0_14_235/a_484_472# 0.001026f
C1456 FILLER_0_16_37/a_124_375# net47 0.002638f
C1457 _444_/a_1308_423# net47 0.040252f
C1458 FILLER_0_15_10/a_124_375# FILLER_0_15_2/a_572_375# 0.012001f
C1459 fanout50/a_36_160# vss 0.009871f
C1460 _133_ _313_/a_67_603# 0.002974f
C1461 net51 output6/a_224_472# 0.006462f
C1462 FILLER_0_8_24/a_572_375# net47 0.0353f
C1463 _127_ _131_ 0.470047f
C1464 FILLER_0_18_107/a_1380_472# vdd 0.009462f
C1465 cal_itt\[1\] _082_ 0.921465f
C1466 _434_/a_2248_156# mask\[6\] 0.022666f
C1467 _119_ _062_ 0.080398f
C1468 _110_ vss 0.131865f
C1469 net29 net19 0.305661f
C1470 FILLER_0_7_72/a_2812_375# trim_mask\[0\] 0.005302f
C1471 net82 cal_itt\[1\] 0.396149f
C1472 FILLER_0_7_104/a_1380_472# vdd 0.011752f
C1473 _424_/a_448_472# vss 0.002076f
C1474 _424_/a_1308_423# vdd 0.002386f
C1475 _030_ vdd 0.244909f
C1476 net41 _444_/a_448_472# 0.031876f
C1477 result[2] _416_/a_448_472# 0.003015f
C1478 net65 _264_/a_224_472# 0.001866f
C1479 net44 _067_ 0.001203f
C1480 _150_ FILLER_0_18_76/a_572_375# 0.008337f
C1481 net78 _007_ 0.054904f
C1482 FILLER_0_16_57/a_1380_472# _175_ 0.002834f
C1483 _397_/a_36_472# _131_ 0.012338f
C1484 net50 _441_/a_1308_423# 0.032656f
C1485 net52 _441_/a_1000_472# 0.011506f
C1486 _412_/a_36_151# _265_/a_244_68# 0.072351f
C1487 _129_ FILLER_0_11_135/a_124_375# 0.009882f
C1488 FILLER_0_19_47/a_484_472# FILLER_0_18_37/a_1468_375# 0.001684f
C1489 _106_ _105_ 0.038327f
C1490 net27 _100_ 0.006783f
C1491 net61 vdd 0.46584f
C1492 _161_ _068_ 0.026092f
C1493 net81 output48/a_224_472# 0.040059f
C1494 net18 _417_/a_796_472# 0.006722f
C1495 _417_/a_1000_472# net30 0.004556f
C1496 ctln[5] vss 0.132862f
C1497 net5 rstn 0.101356f
C1498 _028_ FILLER_0_7_72/a_3260_375# 0.003505f
C1499 FILLER_0_12_136/a_124_375# vss 0.004063f
C1500 FILLER_0_12_136/a_572_375# vdd 0.016972f
C1501 mask\[3\] net64 0.002654f
C1502 FILLER_0_4_197/a_1020_375# net59 0.008989f
C1503 FILLER_0_21_28/a_2276_472# _423_/a_36_151# 0.013806f
C1504 _437_/a_2665_112# vss 0.002056f
C1505 _437_/a_2560_156# vdd 0.0026f
C1506 net31 _292_/a_36_160# 0.010041f
C1507 _114_ FILLER_0_12_124/a_124_375# 0.006974f
C1508 _428_/a_36_151# FILLER_0_14_107/a_36_472# 0.02628f
C1509 result[7] FILLER_0_24_274/a_484_472# 0.006641f
C1510 FILLER_0_3_172/a_36_472# FILLER_0_2_171/a_124_375# 0.001723f
C1511 net20 net61 0.014444f
C1512 net69 FILLER_0_2_111/a_572_375# 0.015789f
C1513 en_co_clk _390_/a_36_68# 0.086301f
C1514 FILLER_0_3_172/a_3172_472# vss 0.003689f
C1515 _129_ _068_ 0.104827f
C1516 output32/a_224_472# net30 0.001139f
C1517 ctlp[1] ctlp[2] 0.002331f
C1518 result[6] _009_ 0.095754f
C1519 _141_ FILLER_0_19_171/a_36_472# 0.001292f
C1520 net65 FILLER_0_9_282/a_572_375# 0.001388f
C1521 net81 mask\[0\] 0.320022f
C1522 _239_/a_36_160# _064_ 0.001292f
C1523 _065_ trim_val\[2\] 0.002278f
C1524 FILLER_0_9_28/a_1380_472# net16 0.005297f
C1525 _098_ FILLER_0_15_228/a_124_375# 0.080662f
C1526 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_124_375# 0.009654f
C1527 output9/a_224_472# net4 0.042449f
C1528 _367_/a_244_472# _157_ 0.002529f
C1529 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_124_375# 0.012221f
C1530 mask\[8\] _025_ 0.036686f
C1531 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_124_375# 0.009654f
C1532 _307_/a_672_472# _113_ 0.006607f
C1533 _012_ FILLER_0_23_44/a_1468_375# 0.002827f
C1534 net63 net80 0.337396f
C1535 FILLER_0_4_213/a_484_472# net59 0.048997f
C1536 FILLER_0_9_28/a_1468_375# vdd 0.009854f
C1537 net55 _451_/a_2225_156# 0.031243f
C1538 FILLER_0_3_54/a_36_472# vss 0.002818f
C1539 FILLER_0_4_177/a_124_375# vdd 0.021637f
C1540 _114_ _128_ 0.047516f
C1541 _074_ net8 0.001023f
C1542 input2/a_36_113# net2 0.015844f
C1543 FILLER_0_4_197/a_484_472# vdd 0.002749f
C1544 _432_/a_2665_112# _139_ 0.004089f
C1545 FILLER_0_7_72/a_3172_472# _058_ 0.001085f
C1546 net34 _108_ 0.297364f
C1547 output31/a_224_472# _418_/a_2665_112# 0.008243f
C1548 _053_ _414_/a_1204_472# 0.003935f
C1549 FILLER_0_14_91/a_572_375# _176_ 0.002444f
C1550 _359_/a_36_488# vdd 0.083138f
C1551 _045_ mask\[1\] 0.024178f
C1552 FILLER_0_22_177/a_1020_375# _435_/a_36_151# 0.059049f
C1553 FILLER_0_19_155/a_124_375# _145_ 0.006057f
C1554 _372_/a_170_472# _122_ 0.018399f
C1555 net63 net34 0.050865f
C1556 net34 net19 0.039959f
C1557 _091_ _136_ 0.075998f
C1558 FILLER_0_6_239/a_124_375# FILLER_0_8_239/a_36_472# 0.001512f
C1559 net57 FILLER_0_13_142/a_484_472# 0.011685f
C1560 vss net14 1.003274f
C1561 _406_/a_36_159# vdd 0.020825f
C1562 FILLER_0_14_181/a_36_472# mask\[1\] 0.006352f
C1563 net75 _265_/a_916_472# 0.001686f
C1564 FILLER_0_8_127/a_124_375# _124_ 0.022175f
C1565 _031_ _160_ 0.004547f
C1566 FILLER_0_15_72/a_124_375# vdd 0.020511f
C1567 FILLER_0_2_171/a_36_472# FILLER_0_2_165/a_36_472# 0.003468f
C1568 fanout55/a_36_160# vss 0.005203f
C1569 _091_ net62 0.019946f
C1570 _115_ _315_/a_36_68# 0.001683f
C1571 net75 _253_/a_1732_68# 0.001047f
C1572 net60 net19 0.102311f
C1573 FILLER_0_21_125/a_36_472# _149_ 0.008849f
C1574 net43 FILLER_0_20_15/a_124_375# 0.005925f
C1575 trim_mask\[3\] vdd 0.233305f
C1576 _164_ vss 0.597051f
C1577 mask\[3\] _103_ 0.055796f
C1578 net81 FILLER_0_15_212/a_124_375# 0.005049f
C1579 net27 FILLER_0_8_263/a_124_375# 0.016669f
C1580 net81 _099_ 0.140011f
C1581 FILLER_0_8_247/a_1380_472# vdd 0.036604f
C1582 FILLER_0_4_49/a_484_472# _440_/a_36_151# 0.006095f
C1583 net47 FILLER_0_4_91/a_124_375# 0.009482f
C1584 _093_ FILLER_0_18_100/a_124_375# 0.011632f
C1585 net27 FILLER_0_14_235/a_124_375# 0.002299f
C1586 _305_/a_36_159# net59 0.007898f
C1587 _323_/a_36_113# net64 0.06154f
C1588 net55 FILLER_0_18_37/a_484_472# 0.006153f
C1589 _069_ _267_/a_36_472# 0.003607f
C1590 FILLER_0_12_136/a_484_472# cal_count\[3\] 0.007275f
C1591 net80 FILLER_0_17_161/a_124_375# 0.021914f
C1592 _011_ vss 0.003987f
C1593 net72 FILLER_0_17_56/a_572_375# 0.004473f
C1594 net32 _420_/a_2665_112# 0.002753f
C1595 _070_ FILLER_0_10_107/a_124_375# 0.009848f
C1596 ctlp[8] vdd 0.115254f
C1597 _441_/a_2248_156# _164_ 0.040396f
C1598 _374_/a_36_68# _061_ 0.026111f
C1599 FILLER_0_3_221/a_36_472# net59 0.075858f
C1600 _093_ FILLER_0_17_72/a_572_375# 0.005609f
C1601 _428_/a_448_472# vdd 0.034564f
C1602 _098_ _433_/a_448_472# 0.027678f
C1603 _428_/a_36_151# vss 0.00285f
C1604 net38 _450_/a_836_156# 0.0039f
C1605 _011_ _422_/a_1000_472# 0.005583f
C1606 FILLER_0_14_181/a_124_375# _097_ 0.001668f
C1607 output48/a_224_472# net2 0.06309f
C1608 net13 vdd 0.264116f
C1609 _129_ _152_ 0.041257f
C1610 net27 _060_ 0.045136f
C1611 net1 _265_/a_468_472# 0.002612f
C1612 cal FILLER_0_1_266/a_572_375# 0.001707f
C1613 output44/a_224_472# net55 0.011586f
C1614 _422_/a_36_151# _009_ 0.015085f
C1615 output6/a_224_472# clkc 0.017846f
C1616 FILLER_0_16_57/a_484_472# vss 0.004107f
C1617 FILLER_0_16_57/a_932_472# vdd 0.005518f
C1618 _170_ _037_ 0.05171f
C1619 _274_/a_3368_68# vss 0.001714f
C1620 net35 _436_/a_2560_156# 0.003198f
C1621 _091_ _429_/a_2665_112# 0.002597f
C1622 _112_ _316_/a_692_472# 0.001614f
C1623 _127_ _076_ 0.137964f
C1624 net15 _449_/a_796_472# 0.006722f
C1625 cal_itt\[3\] _058_ 0.002207f
C1626 _008_ vss 0.355468f
C1627 _056_ _068_ 0.127175f
C1628 fanout54/a_36_160# FILLER_0_19_155/a_36_472# 0.193804f
C1629 FILLER_0_15_212/a_1380_472# vdd 0.003213f
C1630 FILLER_0_15_212/a_932_472# vss 0.019114f
C1631 _246_/a_36_68# vdd 0.047419f
C1632 FILLER_0_15_212/a_36_472# mask\[1\] 0.006865f
C1633 _327_/a_36_472# net74 0.009344f
C1634 FILLER_0_11_109/a_36_472# vss 0.003131f
C1635 _093_ _438_/a_2665_112# 0.003293f
C1636 _072_ _374_/a_36_68# 0.061028f
C1637 output36/a_224_472# _094_ 0.001477f
C1638 result[7] FILLER_0_23_282/a_124_375# 0.016009f
C1639 net32 _419_/a_2560_156# 0.029586f
C1640 _094_ net30 0.188507f
C1641 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_124_375# 0.026339f
C1642 _141_ vss 0.308762f
C1643 net54 _436_/a_448_472# 0.006129f
C1644 net57 _386_/a_1084_68# 0.005716f
C1645 net79 FILLER_0_15_282/a_484_472# 0.006575f
C1646 net36 _137_ 0.048198f
C1647 trim_mask\[1\] FILLER_0_6_47/a_3260_375# 0.003764f
C1648 _434_/a_1204_472# vdd 0.005382f
C1649 net20 FILLER_0_15_212/a_1380_472# 0.001449f
C1650 net75 _112_ 0.041092f
C1651 ctln[1] _073_ 0.001457f
C1652 FILLER_0_5_88/a_124_375# _164_ 0.006288f
C1653 FILLER_0_9_28/a_2364_375# _042_ 0.001216f
C1654 _087_ _122_ 0.007241f
C1655 output44/a_224_472# net17 0.07836f
C1656 _163_ net37 0.079552f
C1657 _277_/a_36_160# _099_ 0.001628f
C1658 net17 _381_/a_36_472# 0.002796f
C1659 _091_ FILLER_0_19_171/a_124_375# 0.028992f
C1660 FILLER_0_1_212/a_124_375# FILLER_0_1_204/a_124_375# 0.003732f
C1661 net57 fanout56/a_36_113# 0.079542f
C1662 _416_/a_36_151# output30/a_224_472# 0.012025f
C1663 FILLER_0_2_171/a_36_472# FILLER_0_2_177/a_36_472# 0.003468f
C1664 output48/a_224_472# valid 0.046397f
C1665 _115_ _219_/a_36_160# 0.001218f
C1666 _091_ _430_/a_796_472# 0.005465f
C1667 FILLER_0_15_290/a_124_375# vdd 0.028723f
C1668 net65 net8 0.203388f
C1669 _446_/a_2665_112# _160_ 0.013745f
C1670 _079_ net21 0.065561f
C1671 vss FILLER_0_8_156/a_124_375# 0.001766f
C1672 vdd FILLER_0_8_156/a_572_375# 0.014611f
C1673 cal_count\[3\] FILLER_0_12_50/a_124_375# 0.060164f
C1674 net35 FILLER_0_22_128/a_1916_375# 0.014552f
C1675 _028_ FILLER_0_7_72/a_1828_472# 0.001777f
C1676 output23/a_224_472# vss 0.075684f
C1677 mask\[0\] FILLER_0_14_181/a_36_472# 0.001234f
C1678 FILLER_0_18_100/a_124_375# _136_ 0.002528f
C1679 net58 cal_itt\[1\] 0.79493f
C1680 _064_ _445_/a_2248_156# 0.013127f
C1681 net68 FILLER_0_6_47/a_572_375# 0.007672f
C1682 _254_/a_244_472# _072_ 0.001552f
C1683 _091_ net4 0.125608f
C1684 FILLER_0_4_123/a_36_472# net69 0.001015f
C1685 net15 _439_/a_448_472# 0.038829f
C1686 output20/a_224_472# net61 0.177946f
C1687 _093_ net35 0.00127f
C1688 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_124_375# 0.001597f
C1689 net61 _419_/a_796_472# 0.00438f
C1690 net60 _419_/a_448_472# 0.05959f
C1691 FILLER_0_21_133/a_36_472# FILLER_0_21_125/a_484_472# 0.013276f
C1692 FILLER_0_4_177/a_572_375# net76 0.009573f
C1693 _360_/a_36_160# net47 0.011731f
C1694 FILLER_0_17_104/a_1020_375# vdd 0.012531f
C1695 net47 output6/a_224_472# 0.070584f
C1696 _013_ FILLER_0_18_37/a_1020_375# 0.023067f
C1697 _161_ _113_ 0.201931f
C1698 FILLER_0_16_89/a_124_375# _451_/a_448_472# 0.001597f
C1699 ctln[2] FILLER_0_1_266/a_484_472# 0.019076f
C1700 _148_ vss 0.025751f
C1701 net54 _354_/a_49_472# 0.002169f
C1702 ctlp[1] FILLER_0_21_286/a_572_375# 0.026009f
C1703 _147_ _435_/a_448_472# 0.001008f
C1704 _450_/a_2225_156# net6 0.001143f
C1705 FILLER_0_9_28/a_1916_375# vdd 0.01295f
C1706 FILLER_0_10_78/a_1468_375# vss 0.054053f
C1707 _432_/a_1308_423# _093_ 0.016365f
C1708 net28 output29/a_224_472# 0.028512f
C1709 ctln[2] net81 0.003762f
C1710 net28 _426_/a_36_151# 0.004878f
C1711 _019_ net21 0.065941f
C1712 FILLER_0_4_123/a_36_472# _152_ 0.003937f
C1713 net16 FILLER_0_8_37/a_124_375# 0.010358f
C1714 net58 FILLER_0_9_282/a_484_472# 0.091905f
C1715 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_124_375# 0.003228f
C1716 net63 _434_/a_2665_112# 0.120476f
C1717 _317_/a_36_113# _014_ 0.037134f
C1718 _015_ vdd 0.27747f
C1719 FILLER_0_15_116/a_124_375# net36 0.003055f
C1720 net39 _445_/a_1204_472# 0.002681f
C1721 FILLER_0_5_72/a_484_472# trim_mask\[1\] 0.012321f
C1722 FILLER_0_5_206/a_36_472# net37 0.009858f
C1723 ctln[1] FILLER_0_1_266/a_484_472# 0.002068f
C1724 net68 net49 0.607379f
C1725 FILLER_0_16_89/a_1380_472# net14 0.049391f
C1726 _426_/a_3041_156# net64 0.001046f
C1727 mask\[2\] FILLER_0_16_154/a_1380_472# 0.017868f
C1728 trim_mask\[4\] _241_/a_224_472# 0.009431f
C1729 _233_/a_36_160# net67 0.001315f
C1730 _452_/a_836_156# net40 0.023204f
C1731 _086_ _127_ 0.042698f
C1732 net25 _051_ 0.090798f
C1733 fanout64/a_36_160# _425_/a_2665_112# 0.005704f
C1734 mask\[3\] mask\[2\] 0.077703f
C1735 FILLER_0_18_171/a_36_472# _432_/a_36_151# 0.059367f
C1736 net20 _015_ 0.005917f
C1737 output42/a_224_472# _221_/a_36_160# 0.017421f
C1738 FILLER_0_22_86/a_932_472# _098_ 0.001442f
C1739 _176_ _451_/a_36_151# 0.003176f
C1740 trim_mask\[1\] _160_ 0.051511f
C1741 FILLER_0_17_72/a_36_472# _131_ 0.002672f
C1742 _035_ _167_ 0.01574f
C1743 _053_ _062_ 0.185944f
C1744 _106_ output18/a_224_472# 0.005393f
C1745 vss FILLER_0_19_134/a_36_472# 0.005204f
C1746 _369_/a_36_68# _367_/a_36_68# 0.038188f
C1747 _153_ vss 0.256017f
C1748 FILLER_0_15_116/a_572_375# net70 0.050592f
C1749 _116_ _162_ 0.00156f
C1750 FILLER_0_23_274/a_124_375# vss 0.017196f
C1751 FILLER_0_23_274/a_36_472# vdd 0.010289f
C1752 output10/a_224_472# net19 0.037774f
C1753 _230_/a_244_68# _070_ 0.001641f
C1754 net26 _423_/a_1000_472# 0.001338f
C1755 net64 FILLER_0_9_282/a_36_472# 0.031302f
C1756 _360_/a_36_160# net74 0.001912f
C1757 _086_ FILLER_0_11_135/a_36_472# 0.004074f
C1758 FILLER_0_5_54/a_572_375# vss 0.002617f
C1759 FILLER_0_5_54/a_1020_375# vdd -0.014642f
C1760 FILLER_0_17_72/a_1468_375# net36 0.047507f
C1761 _412_/a_448_472# net59 0.001462f
C1762 _068_ _152_ 0.006744f
C1763 _451_/a_2449_156# _040_ 0.004434f
C1764 _157_ _160_ 0.010231f
C1765 _442_/a_1000_472# vdd 0.003088f
C1766 FILLER_0_18_177/a_572_375# FILLER_0_20_177/a_484_472# 0.0027f
C1767 _356_/a_36_472# _438_/a_36_151# 0.004432f
C1768 result[6] net33 0.363421f
C1769 net34 _435_/a_1204_472# 0.004285f
C1770 mask\[9\] FILLER_0_20_87/a_36_472# 0.00596f
C1771 _093_ net22 0.041918f
C1772 _321_/a_2590_472# _129_ 0.005391f
C1773 net31 net61 0.053131f
C1774 _242_/a_36_160# net47 0.028264f
C1775 _178_ _402_/a_1948_68# 0.00815f
C1776 FILLER_0_18_177/a_572_375# vdd 0.031241f
C1777 FILLER_0_18_177/a_124_375# vss 0.00364f
C1778 _449_/a_1308_423# _067_ 0.021042f
C1779 net79 FILLER_0_11_282/a_124_375# 0.002239f
C1780 _036_ FILLER_0_3_54/a_36_472# 0.002156f
C1781 net62 FILLER_0_11_282/a_36_472# 0.00149f
C1782 FILLER_0_12_20/a_572_375# vdd 0.013384f
C1783 state\[0\] vss 0.126943f
C1784 _162_ _118_ 0.005444f
C1785 _115_ FILLER_0_10_107/a_484_472# 0.017642f
C1786 _095_ net14 0.043065f
C1787 FILLER_0_18_2/a_36_472# trimb[1] 0.010728f
C1788 _431_/a_1308_423# vdd 0.002397f
C1789 fanout55/a_36_160# _095_ 0.00409f
C1790 FILLER_0_5_128/a_572_375# vss 0.057605f
C1791 _341_/a_49_472# net23 0.031763f
C1792 _053_ FILLER_0_6_90/a_484_472# 0.011443f
C1793 fanout81/a_36_160# cal_itt\[1\] 0.069457f
C1794 _436_/a_2665_112# vss 0.007905f
C1795 FILLER_0_3_221/a_1380_472# vss 0.002804f
C1796 FILLER_0_4_99/a_36_472# net47 0.003903f
C1797 _131_ _118_ 0.001685f
C1798 mask\[7\] FILLER_0_22_128/a_572_375# 0.01909f
C1799 net72 FILLER_0_20_31/a_124_375# 0.011347f
C1800 FILLER_0_3_204/a_124_375# vss 0.017795f
C1801 net74 FILLER_0_13_100/a_36_472# 0.003924f
C1802 net20 _274_/a_716_497# 0.001321f
C1803 output31/a_224_472# _008_ 0.051074f
C1804 FILLER_0_9_28/a_1828_472# net51 0.001502f
C1805 _239_/a_36_160# _065_ 0.032139f
C1806 net63 FILLER_0_20_193/a_572_375# 0.015818f
C1807 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1468_375# 0.086635f
C1808 _439_/a_2665_112# vss 0.003954f
C1809 FILLER_0_22_128/a_1380_472# _433_/a_36_151# 0.001973f
C1810 FILLER_0_19_171/a_1380_472# FILLER_0_19_187/a_36_472# 0.013277f
C1811 _444_/a_2248_156# FILLER_0_8_37/a_484_472# 0.013656f
C1812 ctln[2] net2 0.004284f
C1813 _379_/a_36_472# _063_ 0.071695f
C1814 net36 _040_ 0.429029f
C1815 _428_/a_1308_423# _043_ 0.024052f
C1816 _036_ _164_ 0.011115f
C1817 FILLER_0_21_28/a_1828_472# _424_/a_36_151# 0.001723f
C1818 trimb[4] net44 0.127019f
C1819 ctln[3] FILLER_0_0_232/a_36_472# 0.015594f
C1820 _445_/a_448_472# net49 0.00122f
C1821 net15 FILLER_0_21_60/a_572_375# 0.03167f
C1822 _335_/a_49_472# vdd 0.085394f
C1823 _221_/a_36_160# net40 0.002952f
C1824 FILLER_0_7_162/a_36_472# net37 0.090785f
C1825 net79 FILLER_0_13_290/a_36_472# 0.038324f
C1826 _313_/a_67_603# _227_/a_36_160# 0.032438f
C1827 FILLER_0_16_57/a_124_375# FILLER_0_15_59/a_36_472# 0.001543f
C1828 FILLER_0_8_138/a_124_375# vss 0.00629f
C1829 FILLER_0_16_107/a_484_472# _040_ 0.003828f
C1830 net69 _152_ 0.002532f
C1831 _008_ _419_/a_1000_472# 0.003267f
C1832 _141_ FILLER_0_16_154/a_1020_375# 0.003441f
C1833 mask\[3\] FILLER_0_16_154/a_484_472# 0.002067f
C1834 _126_ net23 0.030487f
C1835 _072_ _121_ 0.041039f
C1836 _114_ _176_ 0.147182f
C1837 _428_/a_36_151# _095_ 0.006658f
C1838 _411_/a_2248_156# cal_itt\[0\] 0.006897f
C1839 _002_ FILLER_0_3_172/a_1828_472# 0.016749f
C1840 net15 _440_/a_36_151# 0.016061f
C1841 _077_ FILLER_0_9_72/a_484_472# 0.004472f
C1842 _119_ FILLER_0_8_156/a_124_375# 0.025304f
C1843 FILLER_0_10_28/a_36_472# net40 0.020589f
C1844 fanout62/a_36_160# net64 0.052109f
C1845 state\[2\] FILLER_0_13_142/a_572_375# 0.007511f
C1846 _056_ _113_ 0.052362f
C1847 net53 FILLER_0_13_142/a_1468_375# 0.002334f
C1848 net57 FILLER_0_3_172/a_36_472# 0.001007f
C1849 _144_ _346_/a_257_69# 0.001089f
C1850 result[4] result[9] 0.101112f
C1851 net81 fanout58/a_36_160# 0.005575f
C1852 _190_/a_36_160# _039_ 0.003926f
C1853 net27 net81 1.118985f
C1854 ctln[1] net2 0.126801f
C1855 FILLER_0_24_274/a_1020_375# vss 0.003553f
C1856 _448_/a_2248_156# _170_ 0.00254f
C1857 _448_/a_1000_472# _037_ 0.03564f
C1858 net63 FILLER_0_18_177/a_1468_375# 0.020059f
C1859 FILLER_0_12_28/a_124_375# vdd 0.040988f
C1860 vss output40/a_224_472# 0.002459f
C1861 _375_/a_36_68# _062_ 0.012855f
C1862 _437_/a_2248_156# _436_/a_36_151# 0.001837f
C1863 _105_ ctlp[1] 0.158795f
C1864 _077_ _453_/a_2665_112# 0.002824f
C1865 FILLER_0_22_128/a_1468_375# vss 0.006619f
C1866 _052_ FILLER_0_19_28/a_484_472# 0.003325f
C1867 net71 FILLER_0_22_107/a_124_375# 0.018295f
C1868 FILLER_0_15_142/a_572_375# net23 0.006327f
C1869 _408_/a_1936_472# cal_count\[0\] 0.001434f
C1870 _207_/a_67_603# vss 0.00837f
C1871 _019_ mask\[1\] 0.007797f
C1872 FILLER_0_3_204/a_124_375# FILLER_0_3_172/a_3260_375# 0.012001f
C1873 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1380_472# 0.013276f
C1874 _084_ vdd 0.134578f
C1875 _441_/a_36_151# FILLER_0_3_78/a_36_472# 0.001723f
C1876 _028_ net52 0.150861f
C1877 _131_ _330_/a_224_472# 0.001186f
C1878 _093_ vdd 1.439861f
C1879 _087_ FILLER_0_3_172/a_932_472# 0.001947f
C1880 _420_/a_36_151# FILLER_0_23_290/a_124_375# 0.026277f
C1881 net61 net77 0.986569f
C1882 _096_ _097_ 0.038778f
C1883 net82 FILLER_0_3_172/a_124_375# 0.011418f
C1884 _077_ FILLER_0_9_28/a_3260_375# 0.01495f
C1885 _035_ vdd 0.215473f
C1886 _093_ FILLER_0_18_107/a_572_375# 0.008393f
C1887 FILLER_0_15_282/a_124_375# vss 0.004893f
C1888 FILLER_0_15_282/a_572_375# vdd 0.002928f
C1889 _120_ FILLER_0_9_72/a_484_472# 0.001645f
C1890 net20 _093_ 0.398457f
C1891 FILLER_0_17_38/a_124_375# vdd 0.01443f
C1892 _065_ trim_val\[3\] 1.235816f
C1893 _064_ _034_ 1.397143f
C1894 FILLER_0_3_172/a_124_375# fanout57/a_36_113# 0.006548f
C1895 _016_ vss 0.069165f
C1896 FILLER_0_7_59/a_572_375# trim_mask\[1\] 0.001548f
C1897 _127_ _321_/a_2034_472# 0.003159f
C1898 net15 _131_ 0.037758f
C1899 _087_ FILLER_0_5_181/a_36_472# 0.154469f
C1900 _132_ _433_/a_36_151# 0.024768f
C1901 input4/a_36_68# net59 0.003625f
C1902 _120_ _453_/a_2665_112# 0.002925f
C1903 net63 _024_ 0.001348f
C1904 FILLER_0_14_123/a_36_472# vdd 0.088525f
C1905 FILLER_0_14_123/a_124_375# vss 0.004985f
C1906 FILLER_0_6_47/a_2724_472# vss 0.020876f
C1907 FILLER_0_6_47/a_3172_472# vdd 0.002089f
C1908 net48 net37 0.081653f
C1909 net56 net54 0.018493f
C1910 _250_/a_36_68# cal_count\[3\] 0.004136f
C1911 _070_ FILLER_0_5_136/a_124_375# 0.001083f
C1912 _053_ FILLER_0_7_104/a_932_472# 0.002529f
C1913 net57 FILLER_0_13_100/a_124_375# 0.012636f
C1914 net72 FILLER_0_19_28/a_572_375# 0.010026f
C1915 FILLER_0_0_266/a_124_375# rstn 0.073089f
C1916 _411_/a_448_472# _073_ 0.004279f
C1917 _119_ _153_ 0.001741f
C1918 _077_ FILLER_0_9_105/a_124_375# 0.007189f
C1919 net32 _421_/a_2248_156# 0.038586f
C1920 _402_/a_1948_68# _401_/a_36_68# 0.012664f
C1921 _115_ FILLER_0_10_78/a_932_472# 0.013773f
C1922 _144_ _436_/a_36_151# 0.029716f
C1923 FILLER_0_12_2/a_572_375# net6 0.058881f
C1924 FILLER_0_15_142/a_124_375# net74 0.005931f
C1925 output48/a_224_472# _079_ 0.003556f
C1926 FILLER_0_22_177/a_36_472# _434_/a_448_472# 0.012285f
C1927 fanout78/a_36_113# _094_ 0.01312f
C1928 fanout56/a_36_113# net36 0.021321f
C1929 FILLER_0_13_212/a_1380_472# vss 0.010223f
C1930 output12/a_224_472# FILLER_0_1_192/a_124_375# 0.032639f
C1931 _443_/a_36_151# _031_ 0.014344f
C1932 _443_/a_1308_423# net69 0.004128f
C1933 _032_ _442_/a_36_151# 0.005632f
C1934 FILLER_0_10_256/a_124_375# FILLER_0_10_247/a_124_375# 0.002036f
C1935 net26 FILLER_0_21_28/a_2812_375# 0.001905f
C1936 _116_ _076_ 0.008283f
C1937 _085_ _070_ 0.058787f
C1938 output46/a_224_472# net40 0.002542f
C1939 FILLER_0_17_200/a_124_375# net21 0.048656f
C1940 _412_/a_1308_423# cal_itt\[1\] 0.009991f
C1941 _415_/a_36_151# vdd 0.115639f
C1942 _446_/a_2560_156# net17 0.00101f
C1943 _000_ _411_/a_796_472# 0.044697f
C1944 _104_ _009_ 0.284256f
C1945 _402_/a_56_567# net47 0.026503f
C1946 vss FILLER_0_5_148/a_36_472# 0.029152f
C1947 _189_/a_67_603# net79 0.008944f
C1948 net2 fanout58/a_36_160# 0.010424f
C1949 net73 FILLER_0_18_107/a_36_472# 0.002425f
C1950 net55 FILLER_0_17_72/a_932_472# 0.024922f
C1951 _001_ net59 0.001439f
C1952 FILLER_0_12_20/a_36_472# _450_/a_448_472# 0.058631f
C1953 FILLER_0_2_111/a_932_472# vss -0.001894f
C1954 FILLER_0_2_111/a_1380_472# vdd 0.002688f
C1955 fanout69/a_36_113# _371_/a_36_113# 0.259508f
C1956 FILLER_0_9_142/a_124_375# calibrate 0.001505f
C1957 _115_ _058_ 0.038308f
C1958 net41 _402_/a_728_93# 0.032823f
C1959 _440_/a_2248_156# vss 0.010006f
C1960 _440_/a_2665_112# vdd -0.002297f
C1961 result[9] _006_ 0.05748f
C1962 en fanout59/a_36_160# 0.242369f
C1963 net15 FILLER_0_13_80/a_36_472# 0.001122f
C1964 net18 _418_/a_1204_472# 0.01349f
C1965 _430_/a_1000_472# vss 0.001626f
C1966 _029_ _365_/a_244_472# 0.001956f
C1967 _076_ _118_ 0.06281f
C1968 _448_/a_448_472# FILLER_0_3_172/a_572_375# 0.00123f
C1969 _448_/a_36_151# FILLER_0_3_172/a_1020_375# 0.001512f
C1970 net62 FILLER_0_15_235/a_572_375# 0.001315f
C1971 trim_mask\[2\] _381_/a_36_472# 0.034251f
C1972 _428_/a_36_151# _332_/a_36_472# 0.004432f
C1973 net57 FILLER_0_16_154/a_1468_375# 0.217874f
C1974 FILLER_0_22_86/a_1468_375# _211_/a_36_160# 0.010334f
C1975 FILLER_0_19_55/a_36_472# FILLER_0_18_53/a_124_375# 0.001684f
C1976 _219_/a_36_160# vdd 0.013125f
C1977 _136_ vdd 1.020301f
C1978 _020_ vss 0.008954f
C1979 state\[1\] net23 0.075055f
C1980 result[9] _103_ 0.034463f
C1981 net82 _443_/a_1204_472# 0.004056f
C1982 FILLER_0_21_28/a_2276_472# _012_ 0.023696f
C1983 net57 _055_ 0.008619f
C1984 output38/a_224_472# _034_ 0.039873f
C1985 net38 _160_ 0.00247f
C1986 net53 FILLER_0_14_107/a_1468_375# 0.001642f
C1987 net70 FILLER_0_14_107/a_932_472# 0.008396f
C1988 FILLER_0_4_107/a_484_472# _031_ 0.002521f
C1989 _114_ _267_/a_36_472# 0.011923f
C1990 net81 _429_/a_36_151# 0.018551f
C1991 net62 vdd 1.53102f
C1992 FILLER_0_1_266/a_572_375# net8 0.016292f
C1993 FILLER_0_1_266/a_484_472# net18 0.010423f
C1994 FILLER_0_15_142/a_572_375# FILLER_0_15_150/a_124_375# 0.012001f
C1995 FILLER_0_13_142/a_124_375# vdd 0.02675f
C1996 fanout72/a_36_113# vss 0.053396f
C1997 ctlp[1] _419_/a_2248_156# 0.028734f
C1998 _438_/a_796_472# vss 0.001171f
C1999 FILLER_0_0_96/a_36_472# vss 0.00344f
C2000 net35 _352_/a_49_472# 0.02594f
C2001 mask\[8\] _352_/a_257_69# 0.003259f
C2002 net52 FILLER_0_5_72/a_1020_375# 0.00799f
C2003 mask\[5\] _009_ 0.001095f
C2004 fanout78/a_36_113# net78 0.004202f
C2005 cal_count\[2\] net40 0.313209f
C2006 net81 net18 0.102876f
C2007 _053_ net14 0.713784f
C2008 _077_ _251_/a_468_472# 0.002497f
C2009 FILLER_0_24_274/a_484_472# _420_/a_36_151# 0.002841f
C2010 _119_ FILLER_0_8_138/a_124_375# 0.006523f
C2011 cal_count\[3\] _310_/a_49_472# 0.00277f
C2012 net16 _182_ 0.05291f
C2013 _158_ _160_ 0.018681f
C2014 _089_ _003_ 0.014763f
C2015 net20 net62 0.058892f
C2016 _176_ _182_ 0.008217f
C2017 FILLER_0_5_72/a_1020_375# net49 0.002208f
C2018 net75 net1 0.098901f
C2019 _311_/a_254_473# net21 0.003733f
C2020 FILLER_0_4_185/a_124_375# vss 0.024832f
C2021 _074_ _123_ 0.157299f
C2022 output29/a_224_472# output30/a_224_472# 0.005147f
C2023 net44 FILLER_0_15_2/a_124_375# 0.017852f
C2024 result[8] ctlp[1] 0.049662f
C2025 _053_ _164_ 0.058788f
C2026 output19/a_224_472# _108_ 0.005075f
C2027 FILLER_0_15_2/a_36_472# vdd 0.104741f
C2028 FILLER_0_15_2/a_572_375# vss 0.055203f
C2029 _077_ _188_ 0.1656f
C2030 _115_ _389_/a_36_148# 0.029505f
C2031 FILLER_0_17_56/a_36_472# FILLER_0_18_53/a_484_472# 0.026657f
C2032 net57 _126_ 0.021705f
C2033 _431_/a_36_151# vdd 0.145005f
C2034 FILLER_0_4_107/a_1380_472# _152_ 0.001297f
C2035 _074_ _073_ 0.040339f
C2036 _412_/a_36_151# vdd 0.080326f
C2037 net4 net22 0.036966f
C2038 output19/a_224_472# net19 0.030721f
C2039 FILLER_0_19_28/a_484_472# net40 0.020293f
C2040 mask\[4\] FILLER_0_18_177/a_36_472# 0.018019f
C2041 _450_/a_448_472# net40 0.00222f
C2042 _414_/a_448_472# _053_ 0.065053f
C2043 _095_ FILLER_0_12_20/a_124_375# 0.001588f
C2044 net66 _160_ 0.097885f
C2045 result[7] _420_/a_448_472# 0.003274f
C2046 FILLER_0_20_177/a_1468_375# mask\[6\] 0.001162f
C2047 FILLER_0_6_177/a_36_472# vss 0.001617f
C2048 _073_ _076_ 0.011358f
C2049 FILLER_0_6_177/a_484_472# vdd 0.007991f
C2050 net36 FILLER_0_15_235/a_484_472# 0.019725f
C2051 _411_/a_36_151# vss 0.035447f
C2052 _376_/a_36_160# vss 0.03081f
C2053 _070_ _062_ 0.06973f
C2054 _072_ FILLER_0_7_233/a_124_375# 0.002279f
C2055 _417_/a_1000_472# _006_ 0.026299f
C2056 FILLER_0_7_104/a_1468_375# _129_ 0.001165f
C2057 FILLER_0_7_104/a_36_472# _131_ 0.002019f
C2058 FILLER_0_7_146/a_36_472# _062_ 0.011622f
C2059 FILLER_0_18_2/a_2812_375# _452_/a_36_151# 0.001597f
C2060 _086_ _116_ 1.316798f
C2061 FILLER_0_18_37/a_1380_472# vss 0.002042f
C2062 FILLER_0_4_49/a_124_375# trim_mask\[1\] 0.006676f
C2063 _335_/a_257_69# _043_ 0.001043f
C2064 _250_/a_36_68# _427_/a_2665_112# 0.002152f
C2065 _014_ _122_ 0.001529f
C2066 _086_ _321_/a_3126_472# 0.001522f
C2067 _429_/a_2248_156# vss 0.040729f
C2068 _429_/a_2665_112# vdd 0.010552f
C2069 _093_ FILLER_0_16_89/a_932_472# 0.002018f
C2070 output32/a_224_472# _006_ 0.001009f
C2071 FILLER_0_17_56/a_124_375# vss 0.00143f
C2072 FILLER_0_17_56/a_572_375# vdd 0.003489f
C2073 _057_ _096_ 0.001547f
C2074 FILLER_0_13_212/a_484_472# mask\[0\] 0.001794f
C2075 _014_ FILLER_0_7_233/a_124_375# 0.00143f
C2076 net19 FILLER_0_23_282/a_124_375# 0.001668f
C2077 _188_ _120_ 0.046757f
C2078 _316_/a_124_24# vss 0.00516f
C2079 _316_/a_848_380# vdd 0.048727f
C2080 FILLER_0_19_195/a_36_472# net21 0.009159f
C2081 net79 _416_/a_1000_472# 0.024811f
C2082 net68 _165_ 0.002748f
C2083 trimb[3] FILLER_0_20_2/a_484_472# 0.001829f
C2084 FILLER_0_15_142/a_484_472# vdd 0.001097f
C2085 _044_ result[3] 0.00251f
C2086 output32/a_224_472# _103_ 0.090957f
C2087 FILLER_0_16_73/a_572_375# net55 0.015207f
C2088 net20 _429_/a_2665_112# 0.062922f
C2089 net53 vdd 0.78288f
C2090 _017_ vss 0.022624f
C2091 FILLER_0_7_72/a_484_472# net52 0.049487f
C2092 net26 _424_/a_796_472# 0.006496f
C2093 _186_ cal_count\[1\] 0.003341f
C2094 _453_/a_36_151# _042_ 0.035846f
C2095 _043_ net40 0.031043f
C2096 _390_/a_36_68# _172_ 0.033476f
C2097 result[8] FILLER_0_24_274/a_124_375# 0.00726f
C2098 FILLER_0_3_54/a_124_375# _160_ 0.004602f
C2099 FILLER_0_20_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001543f
C2100 _086_ _118_ 0.166544f
C2101 _294_/a_224_472# mask\[2\] 0.001715f
C2102 _091_ _430_/a_2665_112# 0.016404f
C2103 en net5 0.892091f
C2104 _386_/a_124_24# vdd 0.014293f
C2105 result[7] _419_/a_1308_423# 0.015718f
C2106 _260_/a_36_68# vdd 0.011119f
C2107 output42/a_224_472# net67 0.05585f
C2108 _090_ _060_ 0.396493f
C2109 FILLER_0_19_171/a_124_375# vdd -0.009473f
C2110 _412_/a_36_151# net9 0.005212f
C2111 FILLER_0_22_86/a_1468_375# net71 0.010224f
C2112 net15 FILLER_0_13_72/a_124_375# 0.006403f
C2113 net58 _425_/a_2665_112# 0.069807f
C2114 _432_/a_2248_156# net21 0.002329f
C2115 _451_/a_448_472# net14 0.04399f
C2116 net36 _437_/a_36_151# 0.002694f
C2117 FILLER_0_10_107/a_36_472# vss 0.003894f
C2118 FILLER_0_10_107/a_484_472# vdd 0.034172f
C2119 _069_ _315_/a_36_68# 0.002242f
C2120 mask\[1\] FILLER_0_15_228/a_124_375# 0.013558f
C2121 FILLER_0_11_282/a_36_472# _416_/a_1308_423# 0.001295f
C2122 _093_ _069_ 0.008325f
C2123 net34 _009_ 0.325819f
C2124 net2 net18 0.030437f
C2125 _108_ mask\[6\] 0.032481f
C2126 _452_/a_1353_112# vdd 0.008539f
C2127 net20 _260_/a_36_68# 0.033776f
C2128 net67 FILLER_0_12_20/a_36_472# 0.054453f
C2129 net63 mask\[6\] 0.146994f
C2130 FILLER_0_7_72/a_572_375# net52 0.022624f
C2131 net68 net40 0.036106f
C2132 _320_/a_1792_472# net79 0.002091f
C2133 net4 vdd 1.218939f
C2134 _211_/a_36_160# net71 0.035804f
C2135 FILLER_0_18_177/a_2276_472# net21 0.01016f
C2136 net60 _009_ 0.006086f
C2137 output18/a_224_472# ctlp[1] 0.039734f
C2138 fanout63/a_36_160# vss 0.008974f
C2139 _164_ _166_ 0.002368f
C2140 FILLER_0_12_124/a_36_472# vss 0.001443f
C2141 _155_ trim_mask\[1\] 0.006536f
C2142 _425_/a_2665_112# calibrate 0.029064f
C2143 FILLER_0_12_136/a_124_375# _428_/a_2665_112# 0.029834f
C2144 _081_ _123_ 0.007811f
C2145 _248_/a_36_68# vss 0.027935f
C2146 _230_/a_244_68# net21 0.00165f
C2147 _067_ FILLER_0_13_80/a_124_375# 0.001857f
C2148 _165_ net67 0.045827f
C2149 _012_ FILLER_0_21_60/a_572_375# 0.011991f
C2150 FILLER_0_16_89/a_124_375# FILLER_0_17_72/a_1916_375# 0.026339f
C2151 _440_/a_36_151# net47 0.013626f
C2152 _073_ _081_ 0.046537f
C2153 _105_ _092_ 0.006701f
C2154 _016_ _095_ 0.034744f
C2155 FILLER_0_14_107/a_124_375# vdd 0.013327f
C2156 _417_/a_2665_112# vss 0.002571f
C2157 _417_/a_2560_156# vdd 0.001658f
C2158 net20 net4 0.650415f
C2159 FILLER_0_9_72/a_36_472# vdd 0.109576f
C2160 FILLER_0_9_72/a_1468_375# vss 0.013085f
C2161 net75 FILLER_0_6_239/a_36_472# 0.009325f
C2162 _114_ FILLER_0_12_136/a_572_375# 0.006974f
C2163 result[6] vdd 0.513079f
C2164 _110_ _098_ 0.09704f
C2165 _420_/a_36_151# FILLER_0_23_282/a_124_375# 0.059049f
C2166 mask\[5\] FILLER_0_20_193/a_36_472# 0.013533f
C2167 _182_ _041_ 0.08834f
C2168 _093_ FILLER_0_18_139/a_36_472# 0.008761f
C2169 _077_ _308_/a_692_472# 0.002268f
C2170 _421_/a_2665_112# _419_/a_2665_112# 0.002588f
C2171 _116_ _090_ 0.122467f
C2172 _091_ FILLER_0_18_209/a_572_375# 0.001343f
C2173 _002_ _087_ 0.00636f
C2174 FILLER_0_5_72/a_932_472# net47 0.003953f
C2175 _095_ FILLER_0_14_123/a_124_375# 0.014486f
C2176 FILLER_0_16_73/a_124_375# _131_ 0.015859f
C2177 _453_/a_2248_156# vdd 0.010767f
C2178 _127_ FILLER_0_11_142/a_36_472# 0.004538f
C2179 net20 result[6] 0.026511f
C2180 _311_/a_1660_473# vdd 0.001435f
C2181 FILLER_0_22_128/a_3172_472# _146_ 0.008065f
C2182 cal_count\[2\] FILLER_0_15_2/a_484_472# 0.015036f
C2183 _015_ _426_/a_1204_472# 0.008883f
C2184 _073_ net65 0.775972f
C2185 net22 _047_ 0.132529f
C2186 _053_ _372_/a_3126_472# 0.001056f
C2187 net23 _160_ 0.030085f
C2188 net31 _093_ 0.274432f
C2189 _432_/a_36_151# vss 0.003647f
C2190 FILLER_0_16_89/a_932_472# _136_ 0.045229f
C2191 net57 state\[1\] 0.154183f
C2192 FILLER_0_18_2/a_124_375# vss 0.003207f
C2193 net63 FILLER_0_19_171/a_1020_375# 0.004794f
C2194 net73 net74 0.016949f
C2195 net54 FILLER_0_22_86/a_1020_375# 0.001597f
C2196 FILLER_0_18_2/a_2276_472# net55 0.006033f
C2197 _136_ FILLER_0_16_154/a_572_375# 0.003842f
C2198 _196_/a_36_160# _045_ 0.036714f
C2199 _162_ net47 0.004104f
C2200 _088_ FILLER_0_3_221/a_124_375# 0.002378f
C2201 _098_ _437_/a_2665_112# 0.003567f
C2202 net62 _283_/a_36_472# 0.002309f
C2203 valid net18 0.03851f
C2204 fanout60/a_36_160# _417_/a_36_151# 0.062739f
C2205 _352_/a_49_472# vdd 0.077542f
C2206 output40/a_224_472# output41/a_224_472# 0.292611f
C2207 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_36_472# 0.002765f
C2208 _308_/a_848_380# FILLER_0_9_105/a_124_375# 0.005599f
C2209 net67 net40 0.886781f
C2210 net54 FILLER_0_22_128/a_1828_472# 0.009504f
C2211 _301_/a_36_472# _051_ 0.001277f
C2212 net35 _213_/a_255_603# 0.001597f
C2213 mask\[5\] FILLER_0_18_177/a_1916_375# 0.002014f
C2214 output27/a_224_472# net5 0.008663f
C2215 FILLER_0_16_89/a_572_375# _040_ 0.004252f
C2216 _118_ _090_ 0.005469f
C2217 mask\[0\] _429_/a_1000_472# 0.020553f
C2218 _448_/a_2665_112# net59 0.005948f
C2219 _270_/a_36_472# _079_ 0.036715f
C2220 _005_ vss 0.01812f
C2221 _005_ _192_/a_255_603# 0.001058f
C2222 net41 _160_ 0.006523f
C2223 _027_ _438_/a_796_472# 0.031292f
C2224 _150_ _438_/a_1204_472# 0.003696f
C2225 FILLER_0_3_172/a_1468_375# net22 0.012895f
C2226 net4 net9 0.008183f
C2227 FILLER_0_18_53/a_572_375# vdd 0.018416f
C2228 _091_ mask\[5\] 0.048311f
C2229 _094_ _418_/a_1308_423# 0.029276f
C2230 _394_/a_728_93# FILLER_0_15_72/a_572_375# 0.02852f
C2231 _094_ _006_ 0.090405f
C2232 _052_ _424_/a_2248_156# 0.005116f
C2233 FILLER_0_16_57/a_1468_375# _131_ 0.015859f
C2234 _285_/a_36_472# mask\[2\] 0.002447f
C2235 _142_ _132_ 0.006253f
C2236 FILLER_0_7_72/a_1020_375# net52 0.00799f
C2237 FILLER_0_18_107/a_2364_375# _433_/a_36_151# 0.002106f
C2238 cal_itt\[2\] _084_ 0.061303f
C2239 _053_ _153_ 0.015583f
C2240 _414_/a_1204_472# net21 0.007637f
C2241 _103_ _094_ 0.280781f
C2242 FILLER_0_4_107/a_484_472# _157_ 0.027364f
C2243 _151_ _154_ 0.108571f
C2244 net74 _390_/a_244_472# 0.001317f
C2245 _132_ mask\[9\] 0.203851f
C2246 _445_/a_448_472# net40 0.044285f
C2247 _307_/a_672_472# _096_ 0.001367f
C2248 _104_ net33 0.037008f
C2249 FILLER_0_24_63/a_124_375# ctlp[8] 0.005758f
C2250 result[9] _420_/a_2248_156# 0.046636f
C2251 FILLER_0_21_28/a_484_472# net40 0.022617f
C2252 net70 FILLER_0_13_100/a_36_472# 0.00585f
C2253 net79 _043_ 0.393702f
C2254 _320_/a_36_472# net21 0.025762f
C2255 FILLER_0_18_2/a_2276_472# net17 0.037088f
C2256 FILLER_0_8_263/a_36_472# net64 0.00399f
C2257 net1 net19 0.024768f
C2258 FILLER_0_13_142/a_572_375# _043_ 0.009328f
C2259 FILLER_0_20_177/a_1020_375# vdd 0.005483f
C2260 net64 FILLER_0_14_235/a_572_375# 0.008689f
C2261 _098_ net14 0.061285f
C2262 _343_/a_49_472# vdd 0.089707f
C2263 state\[0\] _426_/a_2248_156# 0.001198f
C2264 mask\[8\] _423_/a_2248_156# 0.001648f
C2265 net62 _069_ 0.010033f
C2266 _176_ _040_ 0.272465f
C2267 net16 _447_/a_448_472# 0.063057f
C2268 _398_/a_36_113# vdd 0.030449f
C2269 _431_/a_796_472# _137_ 0.002195f
C2270 net41 FILLER_0_18_37/a_124_375# 0.004639f
C2271 fanout72/a_36_113# _095_ 0.001842f
C2272 FILLER_0_10_78/a_932_472# vdd 0.005517f
C2273 _429_/a_36_151# FILLER_0_15_212/a_36_472# 0.001723f
C2274 FILLER_0_20_15/a_1020_375# vdd 0.005198f
C2275 output11/a_224_472# net59 0.002364f
C2276 _426_/a_36_151# _425_/a_36_151# 0.006252f
C2277 net65 FILLER_0_1_266/a_484_472# 0.004635f
C2278 mask\[4\] _143_ 0.352305f
C2279 _422_/a_36_151# vdd 0.177717f
C2280 _432_/a_2248_156# mask\[1\] 0.002293f
C2281 output7/a_224_472# net17 0.001164f
C2282 _115_ _134_ 0.051655f
C2283 _384_/a_224_472# vss 0.004801f
C2284 _432_/a_2665_112# _337_/a_49_472# 0.001051f
C2285 output11/a_224_472# FILLER_0_0_198/a_124_375# 0.00363f
C2286 net81 net65 0.083316f
C2287 cal_count\[2\] _452_/a_1040_527# 0.002003f
C2288 FILLER_0_5_212/a_36_472# _081_ 0.01062f
C2289 _441_/a_1308_423# vdd 0.002837f
C2290 _441_/a_448_472# vss 0.025073f
C2291 _415_/a_36_151# net28 0.001195f
C2292 _131_ net74 0.227843f
C2293 _233_/a_36_160# _033_ 0.017573f
C2294 vdd _047_ 0.175913f
C2295 _031_ _369_/a_244_472# 0.002741f
C2296 net69 _369_/a_36_68# 0.008024f
C2297 net55 _424_/a_448_472# 0.005273f
C2298 trim_val\[2\] _446_/a_2665_112# 0.012621f
C2299 mask\[5\] net33 0.251971f
C2300 _288_/a_224_472# net19 0.002252f
C2301 FILLER_0_16_89/a_932_472# net53 0.012534f
C2302 FILLER_0_16_57/a_1380_472# _394_/a_728_93# 0.001627f
C2303 net75 net76 0.106326f
C2304 _058_ FILLER_0_9_105/a_36_472# 0.011426f
C2305 _415_/a_2560_156# net58 0.002325f
C2306 FILLER_0_2_111/a_124_375# _154_ 0.004032f
C2307 FILLER_0_8_138/a_36_472# _058_ 0.005325f
C2308 net20 _422_/a_36_151# 0.083307f
C2309 output33/a_224_472# net61 0.04987f
C2310 FILLER_0_18_177/a_3172_472# vss 0.002639f
C2311 net52 _442_/a_2560_156# 0.008682f
C2312 _255_/a_224_552# FILLER_0_6_177/a_572_375# 0.001776f
C2313 _053_ _439_/a_2665_112# 0.006037f
C2314 _005_ _416_/a_2248_156# 0.036714f
C2315 FILLER_0_4_152/a_36_472# _386_/a_124_24# 0.004755f
C2316 _176_ FILLER_0_10_94/a_572_375# 0.011743f
C2317 _441_/a_1000_472# _168_ 0.036305f
C2318 _058_ vdd 0.511536f
C2319 _077_ FILLER_0_11_64/a_124_375# 0.013507f
C2320 _356_/a_36_472# mask\[9\] 0.047632f
C2321 net32 _297_/a_36_472# 0.001843f
C2322 ctlp[1] _421_/a_1000_472# 0.007039f
C2323 _091_ net80 0.23053f
C2324 FILLER_0_17_142/a_572_375# _137_ 0.006974f
C2325 FILLER_0_20_31/a_124_375# vdd 0.04619f
C2326 fanout77/a_36_113# vdd 0.032109f
C2327 _028_ FILLER_0_6_79/a_124_375# 0.015932f
C2328 FILLER_0_3_172/a_1468_375# vdd 0.045181f
C2329 _129_ _372_/a_170_472# 0.001985f
C2330 _089_ net76 0.017609f
C2331 FILLER_0_7_72/a_2724_472# _053_ 0.016187f
C2332 FILLER_0_15_290/a_124_375# output30/a_224_472# 0.02894f
C2333 result[6] _420_/a_1308_423# 0.008756f
C2334 _431_/a_36_151# FILLER_0_18_139/a_36_472# 0.002529f
C2335 _070_ net14 0.536953f
C2336 _079_ fanout75/a_36_113# 0.059598f
C2337 net16 _444_/a_448_472# 0.038803f
C2338 fanout80/a_36_113# vss 0.003526f
C2339 FILLER_0_4_123/a_124_375# trim_mask\[4\] 0.004312f
C2340 cal_count\[3\] _278_/a_36_160# 0.008398f
C2341 _147_ _207_/a_67_603# 0.001123f
C2342 net54 _145_ 0.087336f
C2343 _423_/a_36_151# FILLER_0_23_44/a_484_472# 0.001723f
C2344 net62 net28 0.05491f
C2345 net82 FILLER_0_2_171/a_36_472# 0.001777f
C2346 cal net8 0.271166f
C2347 net26 _052_ 0.100927f
C2348 _098_ FILLER_0_15_212/a_932_472# 0.011837f
C2349 FILLER_0_4_123/a_124_375# net47 0.011322f
C2350 _430_/a_36_151# FILLER_0_18_209/a_484_472# 0.001043f
C2351 FILLER_0_15_142/a_572_375# net36 0.006382f
C2352 vdd _416_/a_1308_423# 0.002623f
C2353 vss _416_/a_448_472# 0.004806f
C2354 FILLER_0_7_104/a_1468_375# _152_ 0.009263f
C2355 _422_/a_1308_423# _108_ 0.019345f
C2356 cal_count\[3\] vss 1.35143f
C2357 _033_ net49 0.003904f
C2358 _178_ cal_count\[3\] 0.002061f
C2359 net52 fanout74/a_36_113# 0.001514f
C2360 _141_ _098_ 0.0697f
C2361 FILLER_0_11_64/a_124_375# _120_ 0.004514f
C2362 net46 FILLER_0_20_15/a_572_375# 0.029486f
C2363 output31/a_224_472# _417_/a_2665_112# 0.011048f
C2364 _059_ vss 0.714648f
C2365 FILLER_0_19_47/a_484_472# _012_ 0.001667f
C2366 _017_ _095_ 0.002789f
C2367 _098_ _434_/a_1000_472# 0.00725f
C2368 _089_ FILLER_0_5_198/a_124_375# 0.001517f
C2369 net15 _029_ 0.111797f
C2370 trim_mask\[4\] _170_ 0.09738f
C2371 _415_/a_2665_112# net62 0.003644f
C2372 net74 FILLER_0_13_80/a_36_472# 0.00679f
C2373 _295_/a_244_68# _107_ 0.00123f
C2374 FILLER_0_14_91/a_572_375# _136_ 0.049763f
C2375 _131_ _154_ 0.019221f
C2376 net47 _170_ 0.010131f
C2377 _389_/a_36_148# vdd 0.039639f
C2378 _117_ _060_ 0.149558f
C2379 net79 FILLER_0_12_236/a_124_375# 0.010367f
C2380 _434_/a_36_151# _023_ 0.035162f
C2381 FILLER_0_4_49/a_124_375# net66 0.017584f
C2382 fanout58/a_36_160# cal_itt\[1\] 0.010654f
C2383 mask\[4\] FILLER_0_19_171/a_1380_472# 0.002581f
C2384 output13/a_224_472# _170_ 0.024999f
C2385 output28/a_224_472# FILLER_0_11_282/a_124_375# 0.002977f
C2386 _074_ net47 0.012724f
C2387 net55 fanout55/a_36_160# 0.028425f
C2388 FILLER_0_7_72/a_3260_375# vss 0.053035f
C2389 _128_ _055_ 1.887595f
C2390 _413_/a_1000_472# net82 0.002029f
C2391 trim_mask\[4\] _076_ 0.001824f
C2392 net80 net33 0.037227f
C2393 trim[0] _446_/a_448_472# 0.007307f
C2394 _030_ FILLER_0_3_78/a_36_472# 0.007376f
C2395 net49 FILLER_0_3_78/a_572_375# 0.066078f
C2396 _069_ net4 0.07542f
C2397 _055_ _311_/a_692_473# 0.003127f
C2398 _076_ net47 0.00115f
C2399 FILLER_0_12_124/a_124_375# _126_ 0.02249f
C2400 net2 net65 0.035908f
C2401 _009_ FILLER_0_23_290/a_124_375# 0.002666f
C2402 _291_/a_36_160# vdd 0.010802f
C2403 _320_/a_1120_472# vdd 0.001676f
C2404 _053_ FILLER_0_6_47/a_2724_472# 0.001777f
C2405 net50 FILLER_0_6_79/a_36_472# 0.001614f
C2406 _213_/a_67_603# vss 0.019344f
C2407 net82 FILLER_0_3_172/a_3172_472# 0.007677f
C2408 net34 FILLER_0_22_128/a_3260_375# 0.006974f
C2409 output29/a_224_472# FILLER_0_14_263/a_36_472# 0.0323f
C2410 FILLER_0_4_123/a_124_375# net74 0.002449f
C2411 _074_ FILLER_0_5_172/a_124_375# 0.068565f
C2412 net27 FILLER_0_9_282/a_484_472# 0.006955f
C2413 FILLER_0_22_86/a_484_472# FILLER_0_23_88/a_124_375# 0.001684f
C2414 net34 net33 0.509436f
C2415 FILLER_0_3_172/a_2276_472# net65 0.001777f
C2416 FILLER_0_7_72/a_2276_472# _439_/a_2248_156# 0.013656f
C2417 net20 _291_/a_36_160# 0.002375f
C2418 _111_ _110_ 0.00195f
C2419 _093_ _424_/a_2665_112# 0.001854f
C2420 net55 _404_/a_36_472# 0.001746f
C2421 _070_ FILLER_0_11_109/a_36_472# 0.001091f
C2422 net62 net77 0.122747f
C2423 _128_ _126_ 0.008298f
C2424 _057_ _061_ 0.030546f
C2425 _094_ mask\[2\] 0.089828f
C2426 _132_ _022_ 0.001404f
C2427 net60 net33 0.008865f
C2428 _443_/a_2665_112# vss 0.007913f
C2429 _057_ _311_/a_66_473# 0.042545f
C2430 FILLER_0_5_164/a_36_472# _066_ 0.00611f
C2431 _096_ _161_ 0.00104f
C2432 _123_ FILLER_0_7_233/a_36_472# 0.002812f
C2433 _228_/a_36_68# _090_ 0.018462f
C2434 FILLER_0_9_223/a_484_472# state\[0\] 0.007034f
C2435 FILLER_0_12_220/a_124_375# _248_/a_36_68# 0.005308f
C2436 net17 _164_ 0.007595f
C2437 calibrate _062_ 2.032477f
C2438 FILLER_0_19_28/a_572_375# vdd 0.034691f
C2439 _426_/a_36_151# FILLER_0_9_270/a_36_472# 0.008172f
C2440 _092_ output18/a_224_472# 0.002205f
C2441 trimb[1] FILLER_0_20_2/a_124_375# 0.003431f
C2442 _446_/a_796_472# net66 0.002296f
C2443 trim_val\[1\] _164_ 0.100504f
C2444 cal_count\[3\] _373_/a_438_68# 0.003743f
C2445 ctlp[1] net18 0.088706f
C2446 _413_/a_2248_156# vdd -0.006767f
C2447 _155_ FILLER_0_7_104/a_484_472# 0.003068f
C2448 FILLER_0_16_57/a_484_472# net55 0.001797f
C2449 _425_/a_448_472# FILLER_0_8_247/a_932_472# 0.012285f
C2450 FILLER_0_14_181/a_124_375# _138_ 0.001663f
C2451 FILLER_0_16_89/a_1468_375# vdd 0.038266f
C2452 _062_ net21 0.025648f
C2453 output14/a_224_472# trim_mask\[3\] 0.001155f
C2454 _032_ _031_ 0.013851f
C2455 _070_ FILLER_0_8_156/a_124_375# 0.004329f
C2456 net57 _428_/a_2560_156# 0.010877f
C2457 result[2] net79 0.077934f
C2458 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_124_375# 0.012222f
C2459 output45/a_224_472# ctlp[0] 0.007867f
C2460 _177_ _131_ 0.058938f
C2461 net75 ctln[4] 0.00718f
C2462 net20 _413_/a_2248_156# 0.002515f
C2463 _118_ _117_ 0.032074f
C2464 output45/a_224_472# net45 0.019483f
C2465 net60 FILLER_0_17_282/a_124_375# 0.039003f
C2466 cal_itt\[2\] _260_/a_36_68# 0.004081f
C2467 _214_/a_36_160# FILLER_0_23_88/a_124_375# 0.005398f
C2468 _253_/a_36_68# _074_ 0.026327f
C2469 net56 FILLER_0_19_155/a_36_472# 0.00611f
C2470 _077_ net50 0.312283f
C2471 FILLER_0_4_123/a_124_375# _159_ 0.023643f
C2472 valid net65 0.074257f
C2473 FILLER_0_14_91/a_572_375# net53 0.063988f
C2474 FILLER_0_15_72/a_484_472# cal_count\[1\] 0.013337f
C2475 net36 state\[1\] 0.004105f
C2476 _440_/a_36_151# FILLER_0_6_47/a_1828_472# 0.001512f
C2477 _057_ _072_ 0.048392f
C2478 net31 result[6] 0.002094f
C2479 _083_ _265_/a_224_472# 0.003404f
C2480 FILLER_0_17_72/a_1828_472# vss 0.001443f
C2481 FILLER_0_17_72/a_2276_472# vdd 0.001409f
C2482 _181_ _402_/a_718_527# 0.00461f
C2483 FILLER_0_22_86/a_124_375# net14 0.003962f
C2484 FILLER_0_9_28/a_3260_375# net68 0.009969f
C2485 FILLER_0_21_142/a_36_472# net23 0.001629f
C2486 _419_/a_36_151# vdd -0.110366f
C2487 _065_ net69 0.051511f
C2488 FILLER_0_12_20/a_484_472# _039_ 0.006288f
C2489 FILLER_0_21_142/a_124_375# net54 0.027551f
C2490 mask\[5\] net35 0.003646f
C2491 FILLER_0_19_125/a_36_472# _433_/a_36_151# 0.059367f
C2492 _413_/a_796_472# net59 0.006163f
C2493 _396_/a_224_472# net36 0.00114f
C2494 ctln[5] _448_/a_1308_423# 0.004061f
C2495 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2724_472# 0.026657f
C2496 FILLER_0_3_78/a_484_472# _164_ 0.05311f
C2497 output20/a_224_472# _422_/a_36_151# 0.053592f
C2498 FILLER_0_6_239/a_124_375# net76 0.001286f
C2499 _427_/a_2665_112# vss 0.01229f
C2500 trim_mask\[4\] _081_ 0.111668f
C2501 cal_itt\[2\] net4 0.333682f
C2502 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_36_472# 0.026657f
C2503 net19 _420_/a_448_472# 0.05745f
C2504 FILLER_0_17_142/a_36_472# FILLER_0_19_142/a_124_375# 0.001512f
C2505 ctln[9] vdd 0.221231f
C2506 _372_/a_2034_472# _076_ 0.007461f
C2507 _372_/a_170_472# _068_ 0.037034f
C2508 net74 FILLER_0_13_72/a_124_375# 0.014594f
C2509 _269_/a_36_472# _078_ 0.033601f
C2510 _190_/a_36_160# vdd 0.031799f
C2511 net20 _419_/a_36_151# 0.001225f
C2512 net10 output10/a_224_472# 0.012455f
C2513 _081_ net47 1.302193f
C2514 _000_ net75 0.096899f
C2515 output15/a_224_472# net15 0.028578f
C2516 net76 FILLER_0_3_172/a_1916_375# 0.019901f
C2517 FILLER_0_1_204/a_124_375# net59 0.00999f
C2518 _017_ _332_/a_36_472# 0.033837f
C2519 _077_ FILLER_0_7_72/a_3172_472# 0.001923f
C2520 FILLER_0_21_206/a_36_472# vss 0.004971f
C2521 mask\[3\] FILLER_0_18_177/a_932_472# 0.005654f
C2522 _321_/a_1194_69# vss 0.0011f
C2523 en_co_clk net74 0.039096f
C2524 net26 net40 0.001136f
C2525 net76 net19 0.02061f
C2526 FILLER_0_13_65/a_36_472# fanout72/a_36_113# 0.193651f
C2527 FILLER_0_6_90/a_572_375# _163_ 0.007844f
C2528 net39 _444_/a_1000_472# 0.001323f
C2529 FILLER_0_4_49/a_572_375# net47 0.00654f
C2530 mask\[7\] _435_/a_448_472# 0.064472f
C2531 _394_/a_1336_472# cal_count\[1\] 0.018116f
C2532 net55 _217_/a_36_160# 0.001311f
C2533 cal_count\[3\] _071_ 0.214649f
C2534 net57 _374_/a_36_68# 0.001052f
C2535 net22 FILLER_0_18_209/a_572_375# 0.005202f
C2536 _053_ FILLER_0_6_177/a_36_472# 0.00572f
C2537 net25 FILLER_0_22_86/a_572_375# 0.002444f
C2538 cal_itt\[1\] net18 0.026586f
C2539 FILLER_0_8_107/a_124_375# FILLER_0_7_104/a_484_472# 0.001597f
C2540 _320_/a_36_472# mask\[0\] 0.001026f
C2541 _053_ _376_/a_36_160# 0.005109f
C2542 _069_ _047_ 0.001975f
C2543 _119_ _059_ 0.039711f
C2544 mask\[5\] FILLER_0_19_171/a_1468_375# 0.007169f
C2545 _443_/a_2665_112# FILLER_0_2_165/a_36_472# 0.007491f
C2546 _258_/a_36_160# _081_ 0.00776f
C2547 _149_ vdd 0.379674f
C2548 FILLER_0_2_171/a_124_375# net59 0.006603f
C2549 _086_ FILLER_0_5_172/a_124_375# 0.007355f
C2550 net23 FILLER_0_22_128/a_1380_472# 0.0019f
C2551 result[2] FILLER_0_13_290/a_124_375# 0.015011f
C2552 FILLER_0_18_139/a_572_375# vdd 0.004039f
C2553 FILLER_0_18_139/a_124_375# vss 0.006869f
C2554 mask\[0\] FILLER_0_14_235/a_36_472# 0.287093f
C2555 _408_/a_728_93# _067_ 0.006262f
C2556 FILLER_0_12_124/a_36_472# _332_/a_36_472# 0.004546f
C2557 FILLER_0_9_72/a_1020_375# _439_/a_36_151# 0.059049f
C2558 net78 _420_/a_2248_156# 0.001534f
C2559 _036_ _384_/a_224_472# 0.001921f
C2560 FILLER_0_5_72/a_1468_375# _440_/a_2665_112# 0.001077f
C2561 _121_ net23 0.078786f
C2562 FILLER_0_15_282/a_572_375# output30/a_224_472# 0.029138f
C2563 net19 _419_/a_1308_423# 0.056469f
C2564 FILLER_0_0_130/a_36_472# vdd 0.050082f
C2565 FILLER_0_0_130/a_124_375# vss 0.018073f
C2566 net32 _109_ 0.038411f
C2567 _233_/a_36_160# _444_/a_36_151# 0.032942f
C2568 net74 _081_ 0.093806f
C2569 _430_/a_2665_112# vdd 0.021353f
C2570 FILLER_0_4_152/a_124_375# _386_/a_124_24# 0.010472f
C2571 _016_ _428_/a_2665_112# 0.050481f
C2572 FILLER_0_1_98/a_36_472# FILLER_0_2_93/a_484_472# 0.026657f
C2573 FILLER_0_12_136/a_932_472# FILLER_0_13_142/a_124_375# 0.001684f
C2574 FILLER_0_1_204/a_36_472# net21 0.076466f
C2575 net75 _426_/a_1000_472# 0.002727f
C2576 FILLER_0_16_107/a_124_375# net14 0.004684f
C2577 net71 _437_/a_1000_472# 0.014459f
C2578 result[6] net77 0.111093f
C2579 _435_/a_1000_472# vdd 0.032539f
C2580 mask\[5\] net22 0.04021f
C2581 _086_ net74 0.058077f
C2582 _096_ _056_ 0.001946f
C2583 net63 output35/a_224_472# 0.148302f
C2584 _136_ _451_/a_36_151# 0.043941f
C2585 net38 _444_/a_796_472# 0.002641f
C2586 state\[0\] _070_ 0.009608f
C2587 net80 net35 0.028982f
C2588 result[4] fanout60/a_36_160# 0.027276f
C2589 state\[2\] _225_/a_36_160# 0.037565f
C2590 _430_/a_2665_112# net20 0.005397f
C2591 FILLER_0_20_87/a_36_472# _438_/a_1308_423# 0.010224f
C2592 net38 FILLER_0_8_24/a_36_472# 0.015829f
C2593 _103_ _418_/a_2248_156# 0.012186f
C2594 _443_/a_36_151# net23 0.012359f
C2595 _449_/a_2665_112# en_co_clk 0.002966f
C2596 _003_ _414_/a_796_472# 0.006511f
C2597 FILLER_0_18_76/a_572_375# vss 0.007413f
C2598 FILLER_0_18_76/a_36_472# vdd 0.014249f
C2599 FILLER_0_9_223/a_36_472# _055_ 0.014713f
C2600 ctlp[7] net54 0.004355f
C2601 _079_ _074_ 0.025058f
C2602 net31 _047_ 0.029502f
C2603 _134_ FILLER_0_9_105/a_36_472# 0.004375f
C2604 net33 _434_/a_2665_112# 0.001043f
C2605 _144_ _132_ 0.185339f
C2606 _076_ FILLER_0_3_221/a_484_472# 0.001225f
C2607 _392_/a_36_68# _039_ 0.001522f
C2608 _411_/a_2665_112# net75 0.005223f
C2609 _372_/a_170_472# _152_ 0.037088f
C2610 _077_ cal_itt\[3\] 0.009816f
C2611 net27 FILLER_0_10_247/a_124_375# 0.015466f
C2612 _432_/a_1308_423# net80 0.030835f
C2613 result[9] _421_/a_1204_472# 0.014964f
C2614 net34 net35 2.497277f
C2615 FILLER_0_10_37/a_124_375# _453_/a_36_151# 0.017882f
C2616 cal_count\[3\] _095_ 0.06065f
C2617 FILLER_0_21_125/a_572_375# vdd -0.013698f
C2618 _137_ FILLER_0_17_104/a_1020_375# 0.001676f
C2619 output39/a_224_472# net39 0.129913f
C2620 _134_ vdd 0.482157f
C2621 _079_ _076_ 0.001575f
C2622 FILLER_0_15_142/a_36_472# vss 0.006166f
C2623 FILLER_0_9_28/a_572_375# net41 0.025588f
C2624 ctlp[2] _011_ 0.101324f
C2625 _448_/a_2665_112# trim_val\[4\] 0.004707f
C2626 net73 net70 0.040702f
C2627 output38/a_224_472# _064_ 0.017666f
C2628 _159_ _081_ 0.003646f
C2629 _104_ vdd 0.662413f
C2630 _339_/a_36_160# FILLER_0_19_171/a_36_472# 0.195478f
C2631 _337_/a_665_69# mask\[1\] 0.002125f
C2632 FILLER_0_8_138/a_124_375# _070_ 0.002997f
C2633 _444_/a_36_151# net49 0.007102f
C2634 _142_ mask\[2\] 0.093231f
C2635 _131_ _451_/a_2225_156# 0.008232f
C2636 net59 rstn 0.039664f
C2637 _128_ _426_/a_2665_112# 0.025626f
C2638 _442_/a_36_151# net69 0.048683f
C2639 FILLER_0_21_28/a_3260_375# vdd -0.001166f
C2640 FILLER_0_18_209/a_572_375# vdd 0.021356f
C2641 FILLER_0_18_209/a_124_375# vss 0.004598f
C2642 FILLER_0_5_109/a_572_375# _160_ 0.004207f
C2643 _320_/a_1568_472# _043_ 0.00177f
C2644 net52 FILLER_0_2_93/a_124_375# 0.007787f
C2645 output19/a_224_472# _009_ 0.003174f
C2646 _077_ _039_ 0.104126f
C2647 _410_/a_36_68# _453_/a_36_151# 0.002326f
C2648 output34/a_224_472# net61 0.008309f
C2649 _104_ net20 0.482229f
C2650 output12/a_224_472# net22 0.002662f
C2651 net7 net68 0.032489f
C2652 FILLER_0_8_127/a_124_375# _058_ 0.007791f
C2653 _126_ _320_/a_224_472# 0.003754f
C2654 net36 FILLER_0_20_87/a_36_472# 0.074773f
C2655 net57 FILLER_0_5_164/a_36_472# 0.032208f
C2656 _162_ FILLER_0_6_177/a_124_375# 0.031168f
C2657 FILLER_0_2_93/a_572_375# _030_ 0.001718f
C2658 net63 _435_/a_2248_156# 0.045342f
C2659 _074_ cal_itt\[1\] 0.120296f
C2660 net36 _451_/a_1353_112# 0.01266f
C2661 _093_ FILLER_0_17_104/a_1380_472# 0.014431f
C2662 _427_/a_36_151# net23 0.006844f
C2663 _447_/a_1308_423# _164_ 0.001422f
C2664 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_36_472# 0.003468f
C2665 _144_ _143_ 0.001774f
C2666 FILLER_0_4_107/a_932_472# net47 0.008252f
C2667 _086_ _154_ 0.102849f
C2668 _413_/a_1000_472# net21 0.041643f
C2669 net62 output30/a_224_472# 0.074425f
C2670 _186_ cal_count\[2\] 0.001605f
C2671 FILLER_0_7_72/a_1020_375# FILLER_0_6_79/a_124_375# 0.026339f
C2672 _132_ FILLER_0_11_109/a_124_375# 0.008627f
C2673 _106_ FILLER_0_17_226/a_124_375# 0.061857f
C2674 _115_ _322_/a_124_24# 0.019655f
C2675 FILLER_0_20_107/a_124_375# vdd 0.04384f
C2676 _083_ _084_ 0.016693f
C2677 _029_ net47 2.210804f
C2678 FILLER_0_12_20/a_124_375# net17 0.002167f
C2679 mask\[5\] FILLER_0_20_177/a_484_472# 0.016114f
C2680 _321_/a_170_472# net23 0.025371f
C2681 _449_/a_448_472# cal_count\[3\] 0.007511f
C2682 result[1] _416_/a_36_151# 0.007739f
C2683 _009_ FILLER_0_23_282/a_124_375# 0.012402f
C2684 FILLER_0_3_172/a_3172_472# net21 0.037958f
C2685 net14 FILLER_0_10_94/a_36_472# 0.003391f
C2686 _114_ _136_ 0.003405f
C2687 ctln[7] _442_/a_36_151# 0.007057f
C2688 mask\[5\] vdd 0.79138f
C2689 net72 cal_count\[1\] 0.13509f
C2690 _066_ net59 0.002935f
C2691 FILLER_0_18_107/a_124_375# FILLER_0_20_107/a_36_472# 0.00108f
C2692 net53 _451_/a_36_151# 0.030715f
C2693 net70 _451_/a_1040_527# 0.002679f
C2694 FILLER_0_21_133/a_36_472# vss 0.004298f
C2695 result[6] _421_/a_448_472# 0.038671f
C2696 FILLER_0_13_142/a_1380_472# net23 0.026285f
C2697 _120_ _039_ 0.148356f
C2698 _379_/a_36_472# vdd 0.004183f
C2699 _114_ FILLER_0_13_142/a_124_375# 0.00191f
C2700 _408_/a_56_524# net47 0.040511f
C2701 _425_/a_1204_472# net37 0.001403f
C2702 _075_ _414_/a_448_472# 0.020304f
C2703 net34 net22 0.031404f
C2704 _135_ _134_ 0.038135f
C2705 _144_ _146_ 0.333799f
C2706 net31 _291_/a_36_160# 0.005683f
C2707 _165_ _033_ 0.022734f
C2708 FILLER_0_4_123/a_36_472# FILLER_0_2_111/a_1468_375# 0.00189f
C2709 _415_/a_1308_423# result[1] 0.00761f
C2710 net41 _408_/a_728_93# 0.058816f
C2711 net70 _131_ 0.57653f
C2712 _176_ _055_ 0.001694f
C2713 _431_/a_1308_423# _137_ 0.008805f
C2714 net48 _123_ 0.153061f
C2715 net61 _418_/a_36_151# 0.042401f
C2716 net29 vdd 0.611195f
C2717 net29 _192_/a_67_603# 0.017997f
C2718 _079_ _081_ 1.441057f
C2719 output23/a_224_472# FILLER_0_24_130/a_124_375# 0.006051f
C2720 output36/a_224_472# net36 0.009109f
C2721 net82 FILLER_0_3_221/a_1380_472# 0.008049f
C2722 _426_/a_1308_423# vdd 0.008509f
C2723 output46/a_224_472# FILLER_0_21_28/a_36_472# 0.010684f
C2724 FILLER_0_3_204/a_124_375# net82 0.014222f
C2725 FILLER_0_8_247/a_932_472# calibrate 0.008694f
C2726 _065_ _447_/a_1204_472# 0.017675f
C2727 fanout77/a_36_113# net77 0.031558f
C2728 trim_mask\[2\] FILLER_0_3_54/a_36_472# 0.004063f
C2729 net71 FILLER_0_19_111/a_484_472# 0.004544f
C2730 _132_ FILLER_0_17_104/a_124_375# 0.001918f
C2731 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_572_375# 0.026339f
C2732 _233_/a_36_160# vss 0.01649f
C2733 FILLER_0_5_128/a_124_375# _152_ 0.017496f
C2734 _175_ FILLER_0_15_72/a_484_472# 0.020589f
C2735 _427_/a_448_472# net74 0.051943f
C2736 FILLER_0_2_93/a_36_472# net14 0.005108f
C2737 net72 FILLER_0_17_38/a_36_472# 0.123542f
C2738 _122_ _066_ 0.001217f
C2739 FILLER_0_13_228/a_124_375# net79 0.008554f
C2740 FILLER_0_21_142/a_572_375# FILLER_0_22_128/a_2276_472# 0.001543f
C2741 FILLER_0_17_64/a_36_472# vss 0.006428f
C2742 FILLER_0_18_107/a_2364_375# _022_ 0.001902f
C2743 FILLER_0_18_177/a_1380_472# _139_ 0.00195f
C2744 net23 _146_ 0.034955f
C2745 FILLER_0_17_142/a_36_472# vss 0.008239f
C2746 FILLER_0_17_142/a_484_472# vdd 0.004902f
C2747 net17 output40/a_224_472# 0.00187f
C2748 _335_/a_49_472# _137_ 0.03139f
C2749 output12/a_224_472# vdd 0.106635f
C2750 _151_ _365_/a_36_68# 0.001944f
C2751 FILLER_0_6_47/a_1020_375# vdd 0.016637f
C2752 FILLER_0_14_107/a_124_375# _451_/a_36_151# 0.059049f
C2753 net57 _121_ 0.004182f
C2754 _093_ FILLER_0_18_177/a_2812_375# 0.001989f
C2755 FILLER_0_18_107/a_3172_472# FILLER_0_17_133/a_124_375# 0.001543f
C2756 _427_/a_2665_112# _095_ 0.039612f
C2757 _126_ _176_ 0.057877f
C2758 _072_ FILLER_0_10_214/a_36_472# 0.015199f
C2759 FILLER_0_4_177/a_36_472# net22 0.006506f
C2760 _325_/a_224_472# _118_ 0.004845f
C2761 mask\[9\] FILLER_0_19_111/a_572_375# 0.027695f
C2762 _414_/a_448_472# net21 0.040301f
C2763 trim_mask\[2\] net14 0.060278f
C2764 FILLER_0_12_124/a_36_472# FILLER_0_11_124/a_36_472# 0.05841f
C2765 _186_ _043_ 0.045082f
C2766 _033_ net40 0.298492f
C2767 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1468_375# 0.086635f
C2768 _066_ _169_ 0.222791f
C2769 _256_/a_244_497# vss 0.001274f
C2770 FILLER_0_3_142/a_36_472# _443_/a_36_151# 0.001723f
C2771 _122_ net23 0.276617f
C2772 vdd FILLER_0_12_196/a_124_375# 0.015159f
C2773 _326_/a_36_160# _128_ 0.02761f
C2774 _428_/a_2248_156# net53 0.001188f
C2775 _339_/a_36_160# vss 0.027338f
C2776 trim_mask\[2\] _164_ 1.859062f
C2777 FILLER_0_10_78/a_36_472# cal_count\[3\] 0.266339f
C2778 _161_ _061_ 0.026347f
C2779 FILLER_0_5_128/a_484_472# net47 0.009309f
C2780 _050_ _436_/a_1308_423# 0.022688f
C2781 _081_ cal_itt\[1\] 0.009747f
C2782 _412_/a_2560_156# net1 0.005618f
C2783 net80 vdd 1.045288f
C2784 _444_/a_1000_472# net47 0.036015f
C2785 _161_ _311_/a_66_473# 0.021817f
C2786 _227_/a_36_160# net23 0.055152f
C2787 vdd FILLER_0_6_231/a_124_375# 0.024542f
C2788 net52 vss 1.608047f
C2789 net74 _318_/a_224_472# 0.001513f
C2790 net51 net6 0.142515f
C2791 _114_ net53 0.001275f
C2792 _068_ _313_/a_67_603# 0.012208f
C2793 net57 _443_/a_36_151# 0.003322f
C2794 FILLER_0_8_24/a_484_472# net47 0.042018f
C2795 net67 _450_/a_36_151# 0.067819f
C2796 FILLER_0_18_107/a_2276_472# vdd 0.004405f
C2797 net23 _169_ 0.00151f
C2798 _126_ _124_ 0.012466f
C2799 _434_/a_2560_156# mask\[6\] 0.010913f
C2800 trim_mask\[4\] _163_ 0.003686f
C2801 _273_/a_36_68# vss 0.095582f
C2802 net35 _434_/a_2665_112# 0.024254f
C2803 result[7] FILLER_0_24_290/a_124_375# 0.005026f
C2804 _132_ FILLER_0_19_134/a_124_375# 0.00141f
C2805 result[2] net19 0.065763f
C2806 _128_ _223_/a_36_160# 0.012824f
C2807 _102_ vss 0.068703f
C2808 _394_/a_1336_472# _175_ 0.002792f
C2809 _424_/a_1000_472# vdd 0.002952f
C2810 _413_/a_2248_156# cal_itt\[2\] 0.002527f
C2811 _093_ _137_ 0.201779f
C2812 _024_ net33 0.001047f
C2813 net41 FILLER_0_16_37/a_36_472# 0.009425f
C2814 FILLER_0_15_150/a_124_375# _427_/a_36_151# 0.001822f
C2815 net49 vss 0.689397f
C2816 net47 _163_ 0.64626f
C2817 _003_ cal_itt\[3\] 0.054183f
C2818 net20 FILLER_0_6_231/a_124_375# 0.060499f
C2819 output29/a_224_472# _416_/a_2665_112# 0.011048f
C2820 net34 vdd 1.161282f
C2821 net65 cal_itt\[1\] 0.049124f
C2822 _027_ FILLER_0_18_76/a_572_375# 0.08501f
C2823 _150_ FILLER_0_18_76/a_484_472# 0.003548f
C2824 _122_ FILLER_0_5_172/a_36_472# 0.003007f
C2825 FILLER_0_19_55/a_36_472# _052_ 0.019665f
C2826 net50 _441_/a_1000_472# 0.02354f
C2827 net52 _441_/a_2248_156# 0.023959f
C2828 FILLER_0_4_107/a_36_472# _153_ 0.042459f
C2829 FILLER_0_4_107/a_932_472# _154_ 0.017867f
C2830 _447_/a_2665_112# trim_val\[3\] 0.002721f
C2831 FILLER_0_23_290/a_124_375# FILLER_0_23_282/a_572_375# 0.012001f
C2832 FILLER_0_7_72/a_36_472# net52 0.014911f
C2833 net54 FILLER_0_19_111/a_36_472# 0.003467f
C2834 output36/a_224_472# _417_/a_2248_156# 0.023576f
C2835 net60 vdd 0.575502f
C2836 fanout73/a_36_113# _427_/a_36_151# 0.032681f
C2837 net27 _425_/a_2665_112# 0.001323f
C2838 net20 net34 0.003775f
C2839 net18 _417_/a_1204_472# 0.01349f
C2840 FILLER_0_16_57/a_572_375# net15 0.013085f
C2841 _029_ _154_ 0.116532f
C2842 _417_/a_2248_156# net30 0.048831f
C2843 _411_/a_2665_112# net19 0.00934f
C2844 _072_ _161_ 0.048567f
C2845 FILLER_0_12_136/a_1468_375# vdd 0.026145f
C2846 FILLER_0_12_136/a_1020_375# vss 0.018233f
C2847 _441_/a_2248_156# net49 0.048164f
C2848 FILLER_0_21_206/a_124_375# _204_/a_67_603# 0.003591f
C2849 _132_ net57 0.029479f
C2850 FILLER_0_5_172/a_124_375# _163_ 0.006403f
C2851 _074_ FILLER_0_6_177/a_124_375# 0.003608f
C2852 FILLER_0_8_239/a_124_375# vss 0.017196f
C2853 FILLER_0_8_239/a_36_472# vdd 0.079402f
C2854 FILLER_0_5_72/a_124_375# vdd -0.005497f
C2855 result[7] FILLER_0_24_274/a_1380_472# 0.006454f
C2856 net15 _183_ 0.007353f
C2857 _031_ FILLER_0_2_111/a_572_375# 0.023633f
C2858 net69 FILLER_0_2_111/a_1468_375# 0.021524f
C2859 net14 FILLER_0_4_91/a_124_375# 0.009573f
C2860 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_572_375# 0.086635f
C2861 net72 _038_ 0.013821f
C2862 net20 net60 0.033919f
C2863 _431_/a_2665_112# vdd 0.015335f
C2864 _050_ _208_/a_36_160# 0.001038f
C2865 FILLER_0_5_109/a_124_375# vdd 0.060786f
C2866 _053_ _059_ 0.042128f
C2867 _245_/a_234_472# _067_ 0.005071f
C2868 output20/a_224_472# _104_ 0.019295f
C2869 FILLER_0_5_128/a_484_472# net74 0.025425f
C2870 _292_/a_36_160# _204_/a_67_603# 0.003478f
C2871 trim_val\[0\] trim_mask\[1\] 0.003033f
C2872 _174_ _067_ 0.002678f
C2873 _065_ _064_ 0.007356f
C2874 FILLER_0_9_28/a_2276_472# vdd 0.003276f
C2875 FILLER_0_9_223/a_124_375# vss 0.009569f
C2876 _367_/a_36_68# _157_ 0.013352f
C2877 net20 FILLER_0_8_239/a_36_472# 0.004483f
C2878 FILLER_0_10_78/a_1468_375# FILLER_0_10_94/a_36_472# 0.086743f
C2879 _446_/a_36_151# net40 0.015376f
C2880 _012_ FILLER_0_23_44/a_484_472# 0.001572f
C2881 _096_ _113_ 0.650985f
C2882 net16 _402_/a_728_93# 0.040925f
C2883 net41 FILLER_0_23_44/a_36_472# 0.001116f
C2884 FILLER_0_4_177/a_572_375# vss 0.054783f
C2885 FILLER_0_4_177/a_36_472# vdd 0.114788f
C2886 _081_ FILLER_0_5_148/a_124_375# 0.021583f
C2887 _421_/a_36_151# net19 0.016842f
C2888 _011_ mask\[7\] 0.043474f
C2889 FILLER_0_7_72/a_3260_375# _053_ 0.071059f
C2890 fanout63/a_36_160# _098_ 0.003627f
C2891 net15 FILLER_0_15_59/a_572_375# 0.033245f
C2892 _008_ _418_/a_448_472# 0.052899f
C2893 net36 FILLER_0_15_180/a_572_375# 0.002531f
C2894 net74 _163_ 0.042013f
C2895 _432_/a_2665_112# _019_ 0.002852f
C2896 _114_ _311_/a_1660_473# 0.003304f
C2897 FILLER_0_4_197/a_932_472# net82 0.001826f
C2898 _116_ FILLER_0_13_206/a_124_375# 0.003926f
C2899 _267_/a_36_472# _055_ 0.035376f
C2900 FILLER_0_14_91/a_484_472# _176_ 0.003624f
C2901 FILLER_0_19_155/a_36_472# _145_ 0.005521f
C2902 fanout70/a_36_113# _095_ 0.003087f
C2903 FILLER_0_15_142/a_36_472# _095_ 0.001526f
C2904 _035_ _446_/a_448_472# 0.018273f
C2905 net51 _450_/a_2225_156# 0.009822f
C2906 _276_/a_36_160# vdd 0.010213f
C2907 _441_/a_36_151# _160_ 0.030777f
C2908 net57 FILLER_0_13_142/a_1380_472# 0.011768f
C2909 FILLER_0_15_72/a_572_375# vss 0.007579f
C2910 FILLER_0_15_72/a_36_472# vdd 0.108844f
C2911 FILLER_0_20_193/a_572_375# net35 0.002196f
C2912 FILLER_0_17_200/a_484_472# _093_ 0.007492f
C2913 _419_/a_36_151# net77 0.163616f
C2914 _427_/a_2248_156# state\[1\] 0.001849f
C2915 net52 FILLER_0_2_165/a_36_472# 0.002601f
C2916 net81 FILLER_0_15_212/a_1020_375# 0.006974f
C2917 net64 FILLER_0_12_220/a_1380_472# 0.011079f
C2918 FILLER_0_10_78/a_484_472# FILLER_0_9_72/a_1020_375# 0.001543f
C2919 net47 FILLER_0_4_91/a_36_472# 0.005186f
C2920 FILLER_0_3_2/a_124_375# vdd 0.021963f
C2921 _413_/a_2665_112# net59 0.066623f
C2922 _176_ state\[1\] 0.001641f
C2923 net27 FILLER_0_14_235/a_36_472# 0.003401f
C2924 _307_/a_234_472# _085_ 0.001966f
C2925 _432_/a_36_151# _098_ 0.00957f
C2926 _269_/a_36_472# _080_ 0.003981f
C2927 _083_ _260_/a_36_68# 0.047191f
C2928 _411_/a_796_472# vss 0.00159f
C2929 net55 FILLER_0_18_37/a_1380_472# 0.007432f
C2930 _136_ _137_ 0.417639f
C2931 FILLER_0_12_136/a_1380_472# cal_count\[3\] 0.00383f
C2932 FILLER_0_2_111/a_1380_472# FILLER_0_2_127/a_36_472# 0.013276f
C2933 _322_/a_1084_68# _128_ 0.002629f
C2934 net55 FILLER_0_17_56/a_124_375# 0.014472f
C2935 net72 FILLER_0_17_56/a_484_472# 0.003359f
C2936 _070_ FILLER_0_10_107/a_36_472# 0.013252f
C2937 net78 _421_/a_1204_472# 0.006482f
C2938 _144_ FILLER_0_18_107/a_2364_375# 0.002388f
C2939 _396_/a_224_472# _176_ 0.008359f
C2940 output19/a_224_472# net33 0.126671f
C2941 _441_/a_2560_156# _164_ 0.049213f
C2942 _056_ _061_ 0.445098f
C2943 result[7] _010_ 0.054533f
C2944 _093_ FILLER_0_17_72/a_1468_375# 0.005785f
C2945 FILLER_0_9_223/a_572_375# vdd 0.007158f
C2946 _428_/a_796_472# vdd 0.003502f
C2947 _056_ _311_/a_66_473# 0.026074f
C2948 _098_ _433_/a_796_472# 0.002825f
C2949 _130_ net53 0.00399f
C2950 FILLER_0_16_255/a_124_375# net19 0.008033f
C2951 net4 _083_ 0.135165f
C2952 net31 _104_ 0.102776f
C2953 _437_/a_448_472# net14 0.090442f
C2954 _127_ FILLER_0_11_135/a_36_472# 0.044488f
C2955 _088_ net59 0.270902f
C2956 _076_ FILLER_0_9_142/a_124_375# 0.001774f
C2957 FILLER_0_10_78/a_1380_472# _115_ 0.051132f
C2958 _431_/a_448_472# net36 0.010914f
C2959 net1 _265_/a_244_68# 0.023821f
C2960 _070_ _248_/a_36_68# 0.007095f
C2961 net31 FILLER_0_18_209/a_572_375# 0.001813f
C2962 _163_ _154_ 0.190662f
C2963 net20 FILLER_0_9_223/a_572_375# 0.03118f
C2964 output42/a_224_472# _444_/a_36_151# 0.002701f
C2965 FILLER_0_11_142/a_572_375# net23 0.010863f
C2966 _444_/a_2665_112# trim_val\[0\] 0.007249f
C2967 _081_ FILLER_0_6_177/a_124_375# 0.005524f
C2968 net6 clkc 0.036083f
C2969 _422_/a_1308_423# _009_ 0.008875f
C2970 _431_/a_36_151# _137_ 0.011412f
C2971 FILLER_0_16_57/a_1380_472# vss 0.011192f
C2972 ctln[6] vss 0.45431f
C2973 _077_ _115_ 0.131611f
C2974 net57 _122_ 0.034045f
C2975 state\[0\] calibrate 0.001061f
C2976 cal_count\[3\] FILLER_0_11_124/a_36_472# 0.00702f
C2977 _131_ _331_/a_448_472# 0.007271f
C2978 net15 _449_/a_1204_472# 0.01349f
C2979 output23/a_224_472# mask\[7\] 0.046766f
C2980 _086_ FILLER_0_6_177/a_124_375# 0.043788f
C2981 FILLER_0_20_177/a_572_375# _098_ 0.015373f
C2982 _061_ _068_ 1.857322f
C2983 FILLER_0_15_212/a_932_472# mask\[1\] 0.014799f
C2984 net81 FILLER_0_15_205/a_36_472# 0.081574f
C2985 net55 _452_/a_448_472# 0.05323f
C2986 trim_mask\[2\] _153_ 0.007934f
C2987 _123_ net37 0.002942f
C2988 _072_ _056_ 0.061377f
C2989 _068_ _311_/a_66_473# 0.071325f
C2990 result[7] FILLER_0_23_282/a_36_472# 0.014869f
C2991 _425_/a_36_151# _316_/a_848_380# 0.035903f
C2992 _187_ _408_/a_728_93# 0.002598f
C2993 net25 FILLER_0_23_88/a_124_375# 0.010782f
C2994 _093_ FILLER_0_19_142/a_36_472# 0.002415f
C2995 net76 FILLER_0_1_192/a_124_375# 0.00275f
C2996 _425_/a_2665_112# net18 0.003301f
C2997 _073_ net37 0.013152f
C2998 net57 _169_ 0.033365f
C2999 trim_mask\[1\] FILLER_0_6_47/a_484_472# 0.022211f
C3000 _414_/a_36_151# _079_ 0.037562f
C3001 _434_/a_2665_112# vdd 0.030225f
C3002 _073_ FILLER_0_3_221/a_1468_375# 0.006377f
C3003 FILLER_0_18_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001684f
C3004 _171_ net14 0.020479f
C3005 _043_ _225_/a_36_160# 0.007958f
C3006 _148_ mask\[7\] 0.010238f
C3007 net35 _024_ 0.001335f
C3008 net27 _415_/a_2560_156# 0.008433f
C3009 _114_ _058_ 0.013316f
C3010 net31 mask\[5\] 0.017182f
C3011 output33/a_224_472# result[6] 0.035032f
C3012 _105_ _011_ 0.003998f
C3013 _431_/a_1000_472# net36 0.001771f
C3014 _091_ FILLER_0_19_171/a_1020_375# 0.005708f
C3015 FILLER_0_19_125/a_36_472# _022_ 0.013011f
C3016 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_36_472# 0.002296f
C3017 FILLER_0_3_204/a_124_375# net21 0.010054f
C3018 _322_/a_124_24# vdd 0.01572f
C3019 fanout66/a_36_113# net69 0.001345f
C3020 _421_/a_36_151# _419_/a_448_472# 0.002098f
C3021 _043_ FILLER_0_12_196/a_36_472# 0.001526f
C3022 _115_ _120_ 0.076035f
C3023 FILLER_0_8_138/a_124_375# calibrate 0.013177f
C3024 FILLER_0_15_290/a_36_472# vss 0.010015f
C3025 FILLER_0_2_101/a_124_375# vdd 0.044073f
C3026 _446_/a_2665_112# _034_ 0.002484f
C3027 FILLER_0_4_144/a_124_375# vdd 0.005512f
C3028 vss FILLER_0_8_156/a_36_472# 0.00168f
C3029 vdd FILLER_0_8_156/a_484_472# 0.007249f
C3030 _412_/a_2665_112# vdd 0.014403f
C3031 net35 FILLER_0_22_128/a_2812_375# 0.010399f
C3032 net17 _452_/a_448_472# 0.043154f
C3033 _188_ FILLER_0_12_50/a_124_375# 0.00157f
C3034 net53 _137_ 0.008376f
C3035 _072_ _068_ 0.185471f
C3036 net33 mask\[6\] 0.881813f
C3037 net75 _263_/a_224_472# 0.004396f
C3038 FILLER_0_13_100/a_36_472# net14 0.046864f
C3039 net68 FILLER_0_6_47/a_1468_375# 0.022624f
C3040 net31 net29 0.009564f
C3041 output10/a_224_472# vdd 0.107357f
C3042 _064_ _445_/a_2560_156# 0.005361f
C3043 net15 _439_/a_796_472# 0.001822f
C3044 _185_ _405_/a_255_603# 0.002565f
C3045 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_572_375# 0.001597f
C3046 FILLER_0_18_139/a_484_472# FILLER_0_17_142/a_36_472# 0.026657f
C3047 FILLER_0_18_100/a_124_375# _438_/a_2248_156# 0.001068f
C3048 _052_ vss 0.077815f
C3049 vss _202_/a_36_160# 0.010418f
C3050 net60 _419_/a_796_472# 0.003097f
C3051 net61 _419_/a_1204_472# 0.012025f
C3052 output12/a_224_472# _413_/a_448_472# 0.001495f
C3053 FILLER_0_4_177/a_484_472# net76 0.006746f
C3054 output24/a_224_472# _025_ 0.010601f
C3055 FILLER_0_17_104/a_1468_375# vss 0.001786f
C3056 FILLER_0_17_104/a_36_472# vdd 0.095484f
C3057 _444_/a_36_151# net40 0.032012f
C3058 net47 net6 0.23883f
C3059 mask\[2\] net23 0.431197f
C3060 net62 FILLER_0_14_263/a_36_472# 0.019591f
C3061 _025_ vss 0.016676f
C3062 cal_count\[3\] cal_count\[0\] 0.098735f
C3063 ctlp[1] FILLER_0_21_286/a_484_472# 0.045536f
C3064 _322_/a_848_380# _125_ 0.013667f
C3065 net28 net29 0.178557f
C3066 _440_/a_1000_472# _029_ 0.004334f
C3067 output34/a_224_472# _093_ 0.012298f
C3068 fanout80/a_36_113# _098_ 0.011559f
C3069 _269_/a_36_472# vss 0.014227f
C3070 FILLER_0_18_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001597f
C3071 _114_ _389_/a_36_148# 0.009465f
C3072 _140_ _149_ 0.0088f
C3073 mask\[4\] FILLER_0_19_187/a_124_375# 0.006236f
C3074 FILLER_0_7_72/a_1828_472# _053_ 0.013271f
C3075 net55 FILLER_0_18_53/a_124_375# 0.011674f
C3076 net72 FILLER_0_18_53/a_484_472# 0.001067f
C3077 net52 _036_ 0.013473f
C3078 net50 net68 0.224698f
C3079 net16 FILLER_0_8_37/a_36_472# 0.012905f
C3080 FILLER_0_22_86/a_1468_375# FILLER_0_22_107/a_36_472# 0.007947f
C3081 ctln[3] output11/a_224_472# 0.068614f
C3082 _267_/a_36_472# state\[1\] 0.001647f
C3083 ctlp[8] _051_ 0.010337f
C3084 FILLER_0_23_290/a_124_375# vdd 0.030435f
C3085 net39 _445_/a_2665_112# 0.002831f
C3086 FILLER_0_15_116/a_36_472# net36 0.013546f
C3087 _413_/a_796_472# _002_ 0.009261f
C3088 mask\[2\] FILLER_0_15_212/a_484_472# 0.001641f
C3089 FILLER_0_5_72/a_1380_472# trim_mask\[1\] 0.01221f
C3090 _139_ _337_/a_49_472# 0.024331f
C3091 FILLER_0_16_89/a_124_375# _131_ 0.017319f
C3092 cal net2 0.081236f
C3093 FILLER_0_12_136/a_572_375# _126_ 0.01289f
C3094 _428_/a_36_151# FILLER_0_13_100/a_36_472# 0.004032f
C3095 _036_ net49 0.005235f
C3096 net80 FILLER_0_22_177/a_124_375# 0.013214f
C3097 FILLER_0_4_197/a_1380_472# _088_ 0.017451f
C3098 net81 net37 0.18149f
C3099 _414_/a_2248_156# FILLER_0_5_212/a_36_472# 0.035805f
C3100 _404_/a_36_472# _179_ 0.00141f
C3101 _063_ net67 0.039144f
C3102 _415_/a_2248_156# fanout62/a_36_160# 0.007753f
C3103 FILLER_0_4_99/a_36_472# net14 0.022408f
C3104 output42/a_224_472# _054_ 0.013225f
C3105 net50 _156_ 0.020099f
C3106 _050_ FILLER_0_22_107/a_124_375# 0.002634f
C3107 FILLER_0_20_193/a_572_375# vdd 0.029393f
C3108 _293_/a_36_472# vdd 0.087136f
C3109 FILLER_0_17_72/a_932_472# _131_ 0.002672f
C3110 _143_ _340_/a_36_160# 0.001064f
C3111 _065_ _383_/a_36_472# 0.02518f
C3112 trim_val\[4\] _066_ 0.015621f
C3113 _088_ FILLER_0_5_206/a_124_375# 0.001374f
C3114 _079_ FILLER_0_5_206/a_36_472# 0.008243f
C3115 net16 _160_ 0.354736f
C3116 _420_/a_448_472# _009_ 0.061681f
C3117 FILLER_0_19_111/a_124_375# net14 0.001837f
C3118 _136_ _040_ 0.788826f
C3119 mask\[7\] _436_/a_2665_112# 0.004274f
C3120 net34 FILLER_0_22_177/a_124_375# 0.006974f
C3121 FILLER_0_15_116/a_484_472# net70 0.049569f
C3122 FILLER_0_15_116/a_124_375# net53 0.009286f
C3123 _413_/a_36_151# FILLER_0_3_172/a_1916_375# 0.059049f
C3124 cal_itt\[3\] net76 0.017174f
C3125 _438_/a_36_151# net71 0.053065f
C3126 fanout61/a_36_113# vss 0.05514f
C3127 output10/a_224_472# net9 0.003212f
C3128 _421_/a_2248_156# _109_ 0.001349f
C3129 _432_/a_2665_112# FILLER_0_17_200/a_124_375# 0.006271f
C3130 FILLER_0_5_212/a_36_472# net37 0.007858f
C3131 FILLER_0_18_2/a_36_472# trimb[4] 0.001673f
C3132 _032_ net23 0.019676f
C3133 net52 _449_/a_448_472# 0.001042f
C3134 _286_/a_224_472# _094_ 0.008468f
C3135 _132_ net36 0.029615f
C3136 net31 net34 0.080525f
C3137 FILLER_0_5_54/a_36_472# vdd 0.006056f
C3138 FILLER_0_5_54/a_1468_375# vss 0.053407f
C3139 net32 ctlp[1] 0.032275f
C3140 FILLER_0_17_72/a_2364_375# net36 0.005483f
C3141 FILLER_0_16_241/a_36_472# FILLER_0_15_235/a_572_375# 0.001543f
C3142 output42/a_224_472# vss 0.00418f
C3143 FILLER_0_7_104/a_124_375# _153_ 0.001205f
C3144 FILLER_0_7_104/a_1020_375# _154_ 0.005051f
C3145 _442_/a_2248_156# vdd 0.038702f
C3146 trim_val\[4\] net23 0.014503f
C3147 FILLER_0_21_125/a_572_375# _140_ 0.01659f
C3148 _213_/a_67_603# _098_ 0.018092f
C3149 FILLER_0_18_177/a_1020_375# FILLER_0_20_177/a_932_472# 0.0027f
C3150 FILLER_0_10_37/a_124_375# _042_ 0.002437f
C3151 net34 _435_/a_2665_112# 0.009214f
C3152 net31 net60 0.012623f
C3153 net74 _172_ 0.006643f
C3154 FILLER_0_16_107/a_484_472# _132_ 0.005391f
C3155 _165_ _054_ 0.001337f
C3156 net38 _445_/a_2248_156# 0.029721f
C3157 net50 net67 0.518421f
C3158 FILLER_0_16_241/a_124_375# vss 0.04897f
C3159 FILLER_0_16_241/a_36_472# vdd 0.012388f
C3160 FILLER_0_18_177/a_1468_375# vdd 0.024167f
C3161 net47 _450_/a_2225_156# 0.057106f
C3162 _449_/a_1000_472# _067_ 0.021759f
C3163 _128_ _121_ 0.051501f
C3164 FILLER_0_12_20/a_484_472# vdd 0.003108f
C3165 _112_ vdd 0.086153f
C3166 cal_itt\[3\] FILLER_0_5_198/a_124_375# 0.01268f
C3167 _450_/a_448_472# _039_ 0.047559f
C3168 FILLER_0_18_2/a_2364_375# net40 0.002024f
C3169 output8/a_224_472# _000_ 0.182377f
C3170 cal_count\[3\] _070_ 0.059233f
C3171 net16 FILLER_0_18_37/a_124_375# 0.017482f
C3172 FILLER_0_18_2/a_932_472# trimb[1] 0.011513f
C3173 _095_ FILLER_0_15_72/a_572_375# 0.00352f
C3174 net81 _139_ 0.001762f
C3175 net23 FILLER_0_16_154/a_484_472# 0.001369f
C3176 cal valid 0.06045f
C3177 output9/a_224_472# net76 0.002042f
C3178 FILLER_0_4_197/a_932_472# net21 0.00663f
C3179 _341_/a_665_69# net23 0.001508f
C3180 FILLER_0_5_109/a_484_472# _163_ 0.005054f
C3181 net20 FILLER_0_16_241/a_36_472# 0.001528f
C3182 net69 _031_ 0.450281f
C3183 _070_ _059_ 0.041498f
C3184 net41 _450_/a_3129_107# 0.059083f
C3185 _104_ _421_/a_448_472# 0.001106f
C3186 output47/a_224_472# net38 0.082174f
C3187 _415_/a_2560_156# net18 0.010318f
C3188 _410_/a_36_68# _042_ 0.041079f
C3189 net17 FILLER_0_20_15/a_572_375# 0.018398f
C3190 _370_/a_124_24# vss 0.005764f
C3191 _370_/a_848_380# vdd -0.001256f
C3192 _163_ FILLER_0_5_148/a_124_375# 0.001706f
C3193 _165_ vss 0.048027f
C3194 FILLER_0_7_146/a_36_472# _059_ 0.073041f
C3195 mask\[7\] FILLER_0_22_128/a_1468_375# 0.0178f
C3196 FILLER_0_10_78/a_1468_375# _171_ 0.034647f
C3197 result[8] _011_ 0.001294f
C3198 _008_ _099_ 0.006163f
C3199 _239_/a_36_160# net41 0.006002f
C3200 FILLER_0_7_162/a_124_375# net57 0.033245f
C3201 net63 FILLER_0_20_193/a_484_472# 0.015851f
C3202 fanout53/a_36_160# _427_/a_2665_112# 0.00285f
C3203 _093_ _334_/a_36_160# 0.014676f
C3204 _414_/a_1204_472# _074_ 0.003142f
C3205 _343_/a_49_472# _137_ 0.001419f
C3206 FILLER_0_14_50/a_124_375# cal_count\[3\] 0.002524f
C3207 _428_/a_1000_472# _043_ 0.020031f
C3208 FILLER_0_21_28/a_2724_472# _424_/a_36_151# 0.001723f
C3209 _115_ FILLER_0_9_72/a_932_472# 0.001837f
C3210 net15 FILLER_0_21_60/a_484_472# 0.001552f
C3211 FILLER_0_19_125/a_36_472# _144_ 0.153815f
C3212 _430_/a_1000_472# net21 0.053061f
C3213 _054_ net40 0.072879f
C3214 _247_/a_36_160# vss 0.009308f
C3215 FILLER_0_15_150/a_124_375# mask\[2\] 0.002588f
C3216 _246_/a_36_68# _055_ 0.028938f
C3217 _356_/a_36_472# net36 0.004539f
C3218 FILLER_0_16_57/a_572_375# FILLER_0_15_59/a_484_472# 0.001543f
C3219 fanout69/a_36_113# trim_mask\[4\] 0.027938f
C3220 _024_ vdd 0.091532f
C3221 _176_ _394_/a_718_524# 0.00141f
C3222 _360_/a_36_160# _153_ 0.006561f
C3223 _077_ net22 0.049592f
C3224 _141_ FILLER_0_16_154/a_36_472# 0.00126f
C3225 net55 cal_count\[3\] 0.005157f
C3226 net57 _097_ 0.100409f
C3227 net63 _430_/a_2560_156# 0.009628f
C3228 cal_count\[1\] vdd 0.516859f
C3229 _428_/a_1308_423# _095_ 0.001504f
C3230 _411_/a_2248_156# _084_ 0.002258f
C3231 _002_ FILLER_0_3_172/a_2724_472# 0.006713f
C3232 _443_/a_1204_472# _170_ 0.002808f
C3233 net15 _440_/a_1308_423# 0.015192f
C3234 net2 net37 0.05083f
C3235 _077_ FILLER_0_9_72/a_1380_472# 0.006408f
C3236 _119_ FILLER_0_8_156/a_36_472# 0.010504f
C3237 _061_ _113_ 0.012561f
C3238 state\[2\] FILLER_0_13_142/a_1468_375# 0.018691f
C3239 net53 FILLER_0_13_142/a_484_472# 0.059444f
C3240 mask\[5\] _140_ 0.103728f
C3241 _043_ _039_ 0.001161f
C3242 result[5] _010_ 0.00244f
C3243 _016_ _327_/a_36_472# 0.04536f
C3244 net53 _040_ 0.035628f
C3245 FILLER_0_24_274/a_36_472# vss 0.001013f
C3246 FILLER_0_24_274/a_484_472# vdd 0.004641f
C3247 _367_/a_692_472# net14 0.00423f
C3248 _448_/a_2248_156# _037_ 0.027079f
C3249 net63 FILLER_0_18_177/a_2364_375# 0.009893f
C3250 FILLER_0_12_28/a_36_472# vss 0.003004f
C3251 _162_ _062_ 0.033583f
C3252 FILLER_0_10_78/a_36_472# net52 0.014225f
C3253 _449_/a_2665_112# _172_ 0.003296f
C3254 vss net40 0.898805f
C3255 FILLER_0_2_93/a_484_472# FILLER_0_0_96/a_124_375# 0.001338f
C3256 _178_ net40 0.029542f
C3257 _348_/a_49_472# _146_ 0.001552f
C3258 FILLER_0_22_128/a_2364_375# vss 0.017496f
C3259 FILLER_0_22_128/a_2812_375# vdd 0.003766f
C3260 output22/a_224_472# _435_/a_448_472# 0.010723f
C3261 fanout56/a_36_113# _136_ 0.002316f
C3262 FILLER_0_16_73/a_572_375# _131_ 0.011479f
C3263 net71 FILLER_0_22_107/a_36_472# 0.034505f
C3264 net35 mask\[6\] 0.041818f
C3265 mask\[8\] net35 2.631701f
C3266 FILLER_0_20_15/a_932_472# net40 0.002705f
C3267 FILLER_0_6_79/a_124_375# vss 0.007008f
C3268 FILLER_0_6_79/a_36_472# vdd 0.087807f
C3269 _028_ net50 0.087995f
C3270 _131_ _062_ 0.120189f
C3271 _087_ FILLER_0_3_172/a_1828_472# 0.027954f
C3272 net60 net77 0.046792f
C3273 _053_ FILLER_0_6_47/a_572_375# 0.008213f
C3274 _232_/a_67_603# trim_mask\[1\] 0.022808f
C3275 _308_/a_848_380# _115_ 0.00763f
C3276 result[7] vss 0.49466f
C3277 cal_count\[3\] net17 0.068527f
C3278 net57 mask\[2\] 0.022012f
C3279 net82 FILLER_0_3_172/a_1020_375# 0.010679f
C3280 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_36_472# 0.002765f
C3281 _095_ _281_/a_672_472# 0.00134f
C3282 FILLER_0_10_78/a_484_472# _176_ 0.001731f
C3283 net16 FILLER_0_19_47/a_36_472# 0.009509f
C3284 FILLER_0_15_282/a_36_472# vss 0.004616f
C3285 _120_ FILLER_0_9_72/a_1380_472# 0.001723f
C3286 FILLER_0_17_38/a_572_375# vss 0.007503f
C3287 FILLER_0_17_38/a_36_472# vdd 0.01637f
C3288 trim_mask\[4\] _371_/a_36_113# 0.007529f
C3289 _178_ FILLER_0_17_38/a_572_375# 0.031538f
C3290 net79 _018_ 0.069992f
C3291 FILLER_0_3_172/a_124_375# net65 0.021073f
C3292 net65 _425_/a_2665_112# 0.00628f
C3293 _392_/a_36_68# vdd 0.036386f
C3294 net72 cal_count\[2\] 0.073818f
C3295 vdd FILLER_0_3_212/a_124_375# 0.025095f
C3296 FILLER_0_6_177/a_124_375# _163_ 0.025831f
C3297 net62 _418_/a_36_151# 0.029844f
C3298 _198_/a_67_603# vss 0.003647f
C3299 _081_ _261_/a_36_160# 0.049069f
C3300 _316_/a_124_24# calibrate 0.016936f
C3301 net64 net36 0.037523f
C3302 output43/a_224_472# net40 0.014984f
C3303 fanout69/a_36_113# net74 0.034782f
C3304 valid sample 0.103192f
C3305 _086_ _331_/a_448_472# 0.004356f
C3306 _115_ FILLER_0_9_105/a_572_375# 0.003191f
C3307 en net59 0.490893f
C3308 FILLER_0_14_107/a_124_375# _040_ 0.001861f
C3309 _236_/a_36_160# _064_ 0.039922f
C3310 _028_ FILLER_0_7_72/a_3172_472# 0.001873f
C3311 valid net37 0.051518f
C3312 _053_ net52 0.042556f
C3313 _073_ net8 0.206839f
C3314 _187_ _174_ 0.001321f
C3315 _141_ FILLER_0_18_139/a_1380_472# 0.016119f
C3316 net73 FILLER_0_17_142/a_124_375# 0.003021f
C3317 net52 FILLER_0_6_47/a_2812_375# 0.018463f
C3318 FILLER_0_17_200/a_36_472# mask\[3\] 0.27914f
C3319 _028_ FILLER_0_5_72/a_572_375# 0.00123f
C3320 result[4] _417_/a_2248_156# 0.001436f
C3321 net72 FILLER_0_19_28/a_484_472# 0.004312f
C3322 net55 FILLER_0_19_28/a_124_375# 0.002644f
C3323 _077_ FILLER_0_9_105/a_36_472# 0.003177f
C3324 _077_ FILLER_0_8_138/a_36_472# 0.005953f
C3325 FILLER_0_7_104/a_932_472# _151_ 0.002092f
C3326 net32 _421_/a_2560_156# 0.049213f
C3327 _136_ _334_/a_36_160# 0.005574f
C3328 _402_/a_1948_68# _179_ 0.005403f
C3329 _093_ _437_/a_36_151# 0.056554f
C3330 net48 _079_ 0.012855f
C3331 FILLER_0_12_2/a_484_472# net6 0.005586f
C3332 net75 _316_/a_1084_68# 0.001531f
C3333 _127_ _118_ 0.141388f
C3334 _096_ FILLER_0_14_181/a_124_375# 0.002455f
C3335 _443_/a_1000_472# net69 0.008276f
C3336 FILLER_0_10_256/a_36_472# FILLER_0_10_247/a_36_472# 0.001963f
C3337 net80 _140_ 0.188514f
C3338 _077_ vdd 1.61568f
C3339 net54 FILLER_0_22_107/a_572_375# 0.002239f
C3340 _426_/a_2248_156# FILLER_0_8_239/a_124_375# 0.001068f
C3341 _433_/a_448_472# _145_ 0.045046f
C3342 FILLER_0_10_247/a_36_472# net64 0.059367f
C3343 net46 net40 0.254778f
C3344 _114_ _134_ 0.015298f
C3345 _432_/a_2665_112# FILLER_0_18_177/a_2276_472# 0.021761f
C3346 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_124_375# 0.004426f
C3347 net67 _039_ 0.302826f
C3348 FILLER_0_4_99/a_36_472# _153_ 0.066147f
C3349 _412_/a_2248_156# en 0.022108f
C3350 _328_/a_36_113# vdd 0.136098f
C3351 net22 mask\[6\] 0.612004f
C3352 net71 _433_/a_36_151# 0.014126f
C3353 FILLER_0_17_72/a_124_375# vdd 0.0132f
C3354 _077_ net20 0.094476f
C3355 FILLER_0_11_135/a_36_472# _118_ 0.002496f
C3356 trimb[0] output46/a_224_472# 0.048191f
C3357 output19/a_224_472# vdd 0.063651f
C3358 _430_/a_36_151# vss 0.011779f
C3359 net34 _140_ 0.033459f
C3360 net57 trim_val\[4\] 0.295336f
C3361 _091_ _432_/a_796_472# 0.018082f
C3362 net73 FILLER_0_18_107/a_932_472# 0.016711f
C3363 net55 FILLER_0_17_72/a_1828_472# 0.001217f
C3364 net29 FILLER_0_16_255/a_36_472# 0.086886f
C3365 FILLER_0_2_101/a_36_472# _156_ 0.001487f
C3366 net36 _006_ 0.001331f
C3367 FILLER_0_2_111/a_572_375# _158_ 0.031641f
C3368 FILLER_0_4_107/a_124_375# vdd 0.036972f
C3369 net74 _371_/a_36_113# 0.027966f
C3370 fanout69/a_36_113# _159_ 0.005623f
C3371 _115_ _125_ 0.049021f
C3372 net16 FILLER_0_14_50/a_36_472# 0.001377f
C3373 FILLER_0_19_28/a_124_375# net17 0.007234f
C3374 net47 net37 0.057409f
C3375 FILLER_0_18_171/a_124_375# FILLER_0_19_171/a_124_375# 0.05841f
C3376 _431_/a_36_151# _334_/a_36_160# 0.032942f
C3377 _445_/a_2665_112# net47 0.041188f
C3378 FILLER_0_21_125/a_124_375# _098_ 0.006462f
C3379 _440_/a_2560_156# vss 0.002793f
C3380 FILLER_0_8_138/a_36_472# _120_ 0.006759f
C3381 en net64 0.01789f
C3382 _029_ _365_/a_36_68# 0.013994f
C3383 net54 FILLER_0_20_98/a_124_375# 0.001639f
C3384 net57 FILLER_0_16_154/a_484_472# 0.001532f
C3385 _120_ vdd 0.750809f
C3386 net60 _421_/a_448_472# 0.052759f
C3387 FILLER_0_19_55/a_124_375# FILLER_0_18_53/a_484_472# 0.001684f
C3388 FILLER_0_7_72/a_2812_375# net14 0.025092f
C3389 net72 _043_ 0.05655f
C3390 _038_ vdd 0.043998f
C3391 _128_ _122_ 0.019207f
C3392 FILLER_0_21_28/a_3172_472# _012_ 0.018785f
C3393 net41 _445_/a_2248_156# 0.065247f
C3394 _144_ _208_/a_36_160# 0.00717f
C3395 net38 _034_ 0.025823f
C3396 _017_ FILLER_0_14_107/a_932_472# 0.001941f
C3397 _114_ _267_/a_672_472# 0.001566f
C3398 net79 vss 0.770834f
C3399 net81 _429_/a_1308_423# 0.008913f
C3400 FILLER_0_23_282/a_124_375# vdd -0.003896f
C3401 _303_/a_36_472# vss 0.011549f
C3402 FILLER_0_1_266/a_484_472# net8 0.016327f
C3403 _438_/a_2248_156# vdd 0.024595f
C3404 FILLER_0_13_142/a_1020_375# vdd 0.018221f
C3405 ctlp[1] _419_/a_2560_156# 0.002551f
C3406 FILLER_0_13_142/a_572_375# vss 0.04084f
C3407 net66 _440_/a_448_472# 0.023934f
C3408 FILLER_0_5_172/a_124_375# net37 0.014083f
C3409 net7 _446_/a_36_151# 0.001237f
C3410 net52 FILLER_0_5_72/a_36_472# 0.014911f
C3411 _053_ _359_/a_1044_488# 0.001474f
C3412 _184_ net40 0.122833f
C3413 _128_ net64 0.291788f
C3414 FILLER_0_9_28/a_3172_472# net51 0.047897f
C3415 _211_/a_36_160# _050_ 0.010927f
C3416 _258_/a_36_160# net37 0.006865f
C3417 _151_ net14 0.009212f
C3418 _010_ _108_ 0.002048f
C3419 FILLER_0_18_107/a_124_375# _438_/a_2665_112# 0.029834f
C3420 _106_ FILLER_0_17_226/a_36_472# 0.050907f
C3421 output36/a_224_472# output29/a_224_472# 0.007726f
C3422 _010_ net19 0.408364f
C3423 net19 FILLER_0_14_263/a_124_375# 0.032085f
C3424 output29/a_224_472# net30 0.044542f
C3425 net44 FILLER_0_15_2/a_36_472# 0.007808f
C3426 _371_/a_36_113# _159_ 0.021612f
C3427 FILLER_0_15_2/a_484_472# vss 0.003267f
C3428 _057_ net57 0.873864f
C3429 _081_ FILLER_0_5_136/a_124_375# 0.025819f
C3430 mask\[4\] _201_/a_67_603# 0.029139f
C3431 net23 _208_/a_36_160# 0.112626f
C3432 _091_ _043_ 0.041409f
C3433 net69 _157_ 0.112249f
C3434 _432_/a_36_151# _333_/a_36_160# 0.032942f
C3435 _164_ FILLER_0_6_47/a_36_472# 0.047981f
C3436 _074_ _062_ 0.005012f
C3437 net68 FILLER_0_5_54/a_484_472# 0.047601f
C3438 FILLER_0_11_282/a_124_375# vdd 0.026044f
C3439 mask\[4\] FILLER_0_18_177/a_932_472# 0.016924f
C3440 _326_/a_36_160# FILLER_0_7_104/a_1380_472# 0.002051f
C3441 net15 _453_/a_448_472# 0.040851f
C3442 _328_/a_36_113# _135_ 0.005635f
C3443 _030_ _160_ 0.063581f
C3444 net66 _034_ 0.139638f
C3445 net49 _166_ 0.007445f
C3446 _447_/a_2665_112# net69 0.002067f
C3447 net31 _293_/a_36_472# 0.005692f
C3448 _430_/a_1308_423# net36 0.003317f
C3449 _076_ _062_ 0.978627f
C3450 _000_ _411_/a_1000_472# 0.023042f
C3451 FILLER_0_5_109/a_36_472# FILLER_0_4_107/a_124_375# 0.001684f
C3452 FILLER_0_21_133/a_36_472# _098_ 0.002964f
C3453 mask\[6\] vdd 0.573103f
C3454 _417_/a_2248_156# _006_ 0.039121f
C3455 FILLER_0_7_104/a_932_472# _131_ 0.011713f
C3456 mask\[8\] vdd 0.423606f
C3457 _077_ fanout67/a_36_160# 0.017322f
C3458 _086_ _085_ 0.374127f
C3459 _320_/a_36_472# _090_ 0.001941f
C3460 net56 FILLER_0_17_142/a_124_375# 0.004803f
C3461 _253_/a_36_68# FILLER_0_3_221/a_1468_375# 0.014131f
C3462 _187_ _450_/a_3129_107# 0.00126f
C3463 _256_/a_716_497# _128_ 0.001035f
C3464 _429_/a_2560_156# vss 0.005255f
C3465 FILLER_0_17_56/a_36_472# vss 0.00167f
C3466 FILLER_0_17_56/a_484_472# vdd 0.002789f
C3467 FILLER_0_16_107/a_572_375# FILLER_0_18_107/a_484_472# 0.001512f
C3468 result[6] FILLER_0_21_286/a_124_375# 0.019179f
C3469 FILLER_0_13_212/a_1380_472# mask\[0\] 0.002361f
C3470 fanout52/a_36_160# vdd 0.026513f
C3471 _135_ _120_ 0.017522f
C3472 net10 ctln[4] 0.1323f
C3473 net79 _416_/a_2248_156# 0.026136f
C3474 net55 FILLER_0_18_76/a_572_375# 0.002278f
C3475 output27/a_224_472# net64 0.04953f
C3476 net62 _416_/a_2665_112# 0.037195f
C3477 vdd FILLER_0_13_290/a_36_472# 0.027484f
C3478 vss FILLER_0_13_290/a_124_375# 0.031844f
C3479 cal_count\[3\] _408_/a_1336_472# 0.010351f
C3480 state\[2\] vdd 0.392508f
C3481 FILLER_0_21_142/a_124_375# _433_/a_448_472# 0.006782f
C3482 FILLER_0_7_72/a_484_472# net50 0.059395f
C3483 net26 _424_/a_1204_472# 0.00194f
C3484 _186_ _180_ 0.003034f
C3485 _453_/a_1308_423# _042_ 0.001778f
C3486 _453_/a_448_472# net51 0.006397f
C3487 result[8] FILLER_0_24_274/a_1020_375# 0.00726f
C3488 FILLER_0_20_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001543f
C3489 _440_/a_36_151# _164_ 0.003699f
C3490 net4 net5 0.104296f
C3491 _386_/a_848_380# vss 0.012638f
C3492 FILLER_0_8_127/a_36_472# net74 0.063481f
C3493 result[7] _419_/a_1000_472# 0.015362f
C3494 _104_ output33/a_224_472# 0.032929f
C3495 _175_ vdd 0.147794f
C3496 net75 vss 0.662689f
C3497 _010_ _420_/a_36_151# 0.001838f
C3498 _421_/a_36_151# _009_ 0.00246f
C3499 _163_ _365_/a_36_68# 0.004035f
C3500 FILLER_0_19_171/a_1020_375# vdd 0.025918f
C3501 output35/a_224_472# net33 0.170613f
C3502 output14/a_224_472# FILLER_0_0_130/a_36_472# 0.023414f
C3503 _176_ _121_ 0.035608f
C3504 FILLER_0_22_86/a_484_472# net71 0.00583f
C3505 _377_/a_36_472# trim_mask\[1\] 0.001763f
C3506 FILLER_0_9_28/a_2724_472# trim_val\[0\] 0.001183f
C3507 net15 FILLER_0_13_72/a_36_472# 0.006713f
C3508 _095_ net40 0.674445f
C3509 net10 _000_ 0.001954f
C3510 net36 _097_ 0.022089f
C3511 _451_/a_1040_527# net14 0.029964f
C3512 FILLER_0_5_72/a_932_472# _164_ 0.011079f
C3513 _088_ FILLER_0_4_213/a_572_375# 0.022684f
C3514 fanout60/a_36_160# result[3] 0.00188f
C3515 net7 _447_/a_36_151# 0.002494f
C3516 net55 FILLER_0_21_28/a_2812_375# 0.004005f
C3517 _452_/a_836_156# vdd 0.002533f
C3518 cal cal_itt\[1\] 0.036277f
C3519 FILLER_0_23_290/a_124_375# net77 0.001783f
C3520 FILLER_0_13_65/a_124_375# net72 0.002341f
C3521 _024_ FILLER_0_22_177/a_124_375# 0.005166f
C3522 _036_ net40 0.599505f
C3523 FILLER_0_7_72/a_572_375# net50 0.012932f
C3524 _363_/a_36_68# vdd 0.04306f
C3525 _346_/a_49_472# vss 0.0031f
C3526 trim_mask\[4\] FILLER_0_2_111/a_1020_375# 0.02806f
C3527 _089_ vss 0.018272f
C3528 _003_ vdd 0.032367f
C3529 _050_ net71 0.033192f
C3530 FILLER_0_18_177/a_3172_472# net21 0.010321f
C3531 fanout63/a_36_160# mask\[1\] 0.009907f
C3532 _430_/a_448_472# net36 0.011598f
C3533 _077_ FILLER_0_7_72/a_1380_472# 0.001315f
C3534 FILLER_0_9_28/a_572_375# net16 0.042681f
C3535 _131_ net14 0.037705f
C3536 _004_ vss 0.115789f
C3537 _012_ FILLER_0_21_60/a_484_472# 0.01517f
C3538 FILLER_0_16_89/a_572_375# FILLER_0_17_72/a_2364_375# 0.026339f
C3539 _440_/a_1308_423# net47 0.009738f
C3540 _306_/a_36_68# _043_ 0.001086f
C3541 result[5] vss 0.307366f
C3542 FILLER_0_14_107/a_1020_375# vdd 0.008956f
C3543 FILLER_0_9_72/a_484_472# vss 0.008087f
C3544 FILLER_0_9_72/a_932_472# vdd 0.00604f
C3545 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_124_375# 0.012222f
C3546 _114_ FILLER_0_12_136/a_1468_375# 0.006974f
C3547 _420_/a_36_151# FILLER_0_23_282/a_36_472# 0.001723f
C3548 _013_ mask\[9\] 0.011224f
C3549 mask\[5\] output33/a_224_472# 0.0238f
C3550 net36 mask\[2\] 0.871463f
C3551 net15 FILLER_0_9_60/a_124_375# 0.003602f
C3552 net1 vdd 0.63891f
C3553 _010_ _419_/a_448_472# 0.003295f
C3554 _085_ _090_ 0.001012f
C3555 _116_ _060_ 0.020653f
C3556 _091_ FILLER_0_18_209/a_484_472# 0.001212f
C3557 _002_ _088_ 0.003969f
C3558 _086_ _062_ 0.066419f
C3559 fanout80/a_36_113# net21 0.021603f
C3560 _256_/a_2552_68# _076_ 0.00144f
C3561 _453_/a_2665_112# vss 0.037567f
C3562 _311_/a_2180_473# vdd 0.001974f
C3563 calibrate _059_ 0.506928f
C3564 _015_ _426_/a_2665_112# 0.018623f
C3565 net64 _416_/a_36_151# 0.013586f
C3566 _232_/a_67_603# net66 0.001758f
C3567 FILLER_0_19_47/a_36_472# _424_/a_1308_423# 0.010224f
C3568 FILLER_0_18_2/a_572_375# net44 0.072627f
C3569 _432_/a_36_151# mask\[1\] 0.003001f
C3570 _238_/a_67_603# net14 0.004718f
C3571 _131_ _404_/a_36_472# 0.031567f
C3572 _079_ net37 0.408392f
C3573 _426_/a_36_151# _317_/a_36_113# 0.001082f
C3574 output8/a_224_472# _078_ 0.001267f
C3575 FILLER_0_18_2/a_3172_472# net55 0.00602f
C3576 _136_ FILLER_0_16_154/a_1468_375# 0.0028f
C3577 _428_/a_36_151# _131_ 0.00821f
C3578 net3 FILLER_0_15_2/a_572_375# 0.004377f
C3579 _443_/a_2248_156# net59 0.002471f
C3580 net52 _387_/a_36_113# 0.02405f
C3581 fanout49/a_36_160# net49 0.032999f
C3582 FILLER_0_9_28/a_3260_375# vss 0.05542f
C3583 net40 output41/a_224_472# 0.081551f
C3584 _308_/a_848_380# FILLER_0_9_105/a_36_472# 0.15783f
C3585 _261_/a_36_160# _163_ 0.002002f
C3586 FILLER_0_16_89/a_1468_375# _040_ 0.004985f
C3587 _118_ _060_ 0.002868f
C3588 vdd _433_/a_2248_156# 0.008127f
C3589 mask\[0\] _429_/a_2248_156# 0.016246f
C3590 _294_/a_224_472# mask\[3\] 0.00233f
C3591 fanout77/a_36_113# _418_/a_36_151# 0.001082f
C3592 _005_ mask\[1\] 0.246517f
C3593 net41 _034_ 0.026084f
C3594 _308_/a_848_380# vdd 0.013895f
C3595 _288_/a_224_472# vdd 0.002071f
C3596 FILLER_0_3_172/a_2364_375# net22 0.013028f
C3597 FILLER_0_18_53/a_484_472# vdd 0.002358f
C3598 FILLER_0_18_53/a_36_472# vss 0.001471f
C3599 _094_ _418_/a_1000_472# 0.053462f
C3600 FILLER_0_17_133/a_124_375# vss 0.015434f
C3601 FILLER_0_17_133/a_36_472# vdd 0.097394f
C3602 net10 _411_/a_2665_112# 0.007912f
C3603 _189_/a_67_603# vdd 0.01494f
C3604 input5/a_36_113# vss 0.005833f
C3605 _052_ _424_/a_2560_156# 0.003401f
C3606 FILLER_0_16_57/a_484_472# _131_ 0.008223f
C3607 FILLER_0_5_109/a_36_472# _363_/a_36_68# 0.001024f
C3608 FILLER_0_7_72/a_1020_375# net50 0.014749f
C3609 _221_/a_36_160# vdd 0.073414f
C3610 FILLER_0_9_60/a_124_375# net51 0.002346f
C3611 output47/a_224_472# trimb[4] 0.044883f
C3612 FILLER_0_3_204/a_36_472# net59 0.001606f
C3613 fanout55/a_36_160# FILLER_0_13_80/a_36_472# 0.003699f
C3614 net55 FILLER_0_17_64/a_36_472# 0.034504f
C3615 _004_ _416_/a_2248_156# 0.001078f
C3616 _151_ _153_ 0.027868f
C3617 net20 _288_/a_224_472# 0.003019f
C3618 net36 FILLER_0_16_115/a_124_375# 0.001706f
C3619 _132_ _124_ 0.005668f
C3620 _321_/a_170_472# _176_ 0.059301f
C3621 net74 _390_/a_36_68# 0.008011f
C3622 ctlp[3] vss 0.037106f
C3623 _273_/a_36_68# _070_ 0.013247f
C3624 _189_/a_67_603# net20 0.011939f
C3625 FILLER_0_7_104/a_1380_472# _133_ 0.004838f
C3626 result[9] _420_/a_2560_156# 0.002295f
C3627 FILLER_0_10_28/a_124_375# vss 0.013087f
C3628 FILLER_0_10_28/a_36_472# vdd 0.092132f
C3629 _069_ _120_ 0.030804f
C3630 net16 _408_/a_728_93# 0.107634f
C3631 _126_ _136_ 0.086459f
C3632 FILLER_0_18_2/a_3172_472# net17 0.002402f
C3633 FILLER_0_15_235/a_124_375# vdd -0.006807f
C3634 result[0] vdd 0.193436f
C3635 net54 _210_/a_67_603# 0.001108f
C3636 FILLER_0_9_105/a_572_375# vdd 0.074717f
C3637 FILLER_0_13_142/a_1468_375# _043_ 0.009636f
C3638 FILLER_0_20_177/a_1468_375# vss 0.053913f
C3639 FILLER_0_20_177/a_36_472# vdd 0.114932f
C3640 net81 _100_ 0.24831f
C3641 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_572_375# 0.086635f
C3642 net64 FILLER_0_14_235/a_484_472# 0.012355f
C3643 net35 _423_/a_2665_112# 0.019085f
C3644 mask\[5\] _137_ 0.002972f
C3645 _132_ fanout71/a_36_113# 0.055078f
C3646 cal_itt\[1\] FILLER_0_3_221/a_1468_375# 0.020427f
C3647 _398_/a_36_113# net44 0.011803f
C3648 ctln[9] _447_/a_448_472# 0.003564f
C3649 net16 _447_/a_796_472# 0.003278f
C3650 net36 FILLER_0_15_212/a_572_375# 0.004606f
C3651 net20 FILLER_0_15_235/a_124_375# 0.001278f
C3652 net70 FILLER_0_16_115/a_36_472# 0.003407f
C3653 _077_ _449_/a_36_151# 0.002475f
C3654 _429_/a_36_151# FILLER_0_15_212/a_932_472# 0.001723f
C3655 _426_/a_36_151# _425_/a_1308_423# 0.001518f
C3656 _116_ _118_ 0.054068f
C3657 FILLER_0_20_15/a_1468_375# vss 0.055156f
C3658 FILLER_0_20_15/a_36_472# vdd 0.086947f
C3659 fanout70/a_36_113# FILLER_0_15_116/a_572_375# 0.003553f
C3660 _233_/a_36_160# net17 0.003831f
C3661 FILLER_0_18_107/a_124_375# vdd 0.030961f
C3662 _321_/a_3126_472# _118_ 0.002754f
C3663 net52 net55 0.016401f
C3664 _267_/a_36_472# _121_ 0.041237f
C3665 _422_/a_1308_423# vdd 0.004083f
C3666 _008_ net18 0.113775f
C3667 _168_ vss 0.171346f
C3668 _062_ _090_ 0.010805f
C3669 _106_ FILLER_0_17_218/a_124_375# 0.004655f
C3670 net79 FILLER_0_12_220/a_124_375# 0.010895f
C3671 _441_/a_796_472# vss 0.001231f
C3672 net34 output33/a_224_472# 0.077682f
C3673 FILLER_0_8_127/a_124_375# _077_ 0.005095f
C3674 _415_/a_36_151# result[1] 0.012965f
C3675 _063_ _033_ 0.250192f
C3676 _067_ FILLER_0_13_72/a_572_375# 0.001874f
C3677 net69 _158_ 0.033459f
C3678 _031_ _369_/a_36_68# 0.050502f
C3679 mask\[9\] net71 0.344312f
C3680 ctlp[3] _107_ 0.132316f
C3681 _064_ _446_/a_2665_112# 0.039211f
C3682 _053_ _165_ 0.123461f
C3683 FILLER_0_9_223/a_124_375# _070_ 0.002989f
C3684 mask\[5\] _049_ 0.008296f
C3685 FILLER_0_16_241/a_36_472# _282_/a_36_160# 0.006647f
C3686 output33/a_224_472# net60 0.002526f
C3687 FILLER_0_14_81/a_36_472# cal_count\[1\] 0.034486f
C3688 _432_/a_1000_472# _093_ 0.007509f
C3689 _005_ _416_/a_2560_156# 0.004273f
C3690 _176_ FILLER_0_10_94/a_484_472# 0.009483f
C3691 _125_ vdd 0.218505f
C3692 FILLER_0_5_117/a_124_375# vss 0.001764f
C3693 _141_ net56 0.012364f
C3694 _131_ FILLER_0_17_104/a_572_375# 0.003214f
C3695 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_36_472# 0.003468f
C3696 FILLER_0_6_239/a_36_472# vdd 0.092399f
C3697 FILLER_0_6_239/a_124_375# vss 0.017355f
C3698 output35/a_224_472# net35 0.007217f
C3699 ctlp[1] _421_/a_2248_156# 0.012937f
C3700 _139_ _019_ 0.094494f
C3701 net69 net66 0.09789f
C3702 net15 _423_/a_36_151# 0.003422f
C3703 FILLER_0_17_142/a_484_472# _137_ 0.003953f
C3704 FILLER_0_20_31/a_36_472# vss 0.004923f
C3705 _444_/a_2665_112# FILLER_0_6_37/a_124_375# 0.005477f
C3706 _449_/a_36_151# _038_ 0.019666f
C3707 FILLER_0_3_172/a_2364_375# vdd -0.010717f
C3708 _359_/a_36_488# _133_ 0.04287f
C3709 FILLER_0_5_54/a_572_375# _440_/a_36_151# 0.026916f
C3710 FILLER_0_11_101/a_124_375# net14 0.011983f
C3711 result[6] _420_/a_1000_472# 0.007761f
C3712 net63 FILLER_0_20_177/a_932_472# 0.004375f
C3713 FILLER_0_9_28/a_124_375# output42/a_224_472# 0.003337f
C3714 _108_ vss 0.160825f
C3715 net20 FILLER_0_6_239/a_36_472# 0.005138f
C3716 net16 FILLER_0_16_37/a_36_472# 0.015199f
C3717 FILLER_0_16_73/a_36_472# FILLER_0_16_57/a_1380_472# 0.013276f
C3718 _163_ FILLER_0_5_136/a_124_375# 0.009765f
C3719 _251_/a_468_472# vss 0.001679f
C3720 net81 FILLER_0_8_263/a_124_375# 0.026195f
C3721 output11/a_224_472# FILLER_0_0_232/a_36_472# 0.023414f
C3722 net63 vss 0.566021f
C3723 net19 vss 1.140787f
C3724 fanout80/a_36_113# mask\[1\] 0.020046f
C3725 net50 _033_ 0.003088f
C3726 net36 FILLER_0_15_205/a_124_375# 0.004337f
C3727 _232_/a_255_603# net47 0.001241f
C3728 _423_/a_36_151# FILLER_0_23_44/a_1380_472# 0.001723f
C3729 net76 net22 0.118787f
C3730 net49 net17 0.029142f
C3731 net62 result[1] 0.061866f
C3732 net81 FILLER_0_14_235/a_124_375# 0.01391f
C3733 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1468_375# 0.016748f
C3734 FILLER_0_9_28/a_1380_472# _120_ 0.00154f
C3735 net15 FILLER_0_17_72/a_36_472# 0.006905f
C3736 _414_/a_448_472# _074_ 0.008725f
C3737 vss _416_/a_796_472# 0.001468f
C3738 output46/a_224_472# vdd 0.043652f
C3739 _422_/a_1000_472# _108_ 0.027806f
C3740 _188_ vss 0.032923f
C3741 _069_ state\[2\] 0.023375f
C3742 net80 _137_ 0.260786f
C3743 _281_/a_672_472# _098_ 0.002084f
C3744 net65 FILLER_0_2_171/a_36_472# 0.023858f
C3745 FILLER_0_21_206/a_36_472# net21 0.132984f
C3746 net52 net82 0.108202f
C3747 FILLER_0_8_107/a_36_472# _062_ 0.001832f
C3748 _140_ _024_ 0.00287f
C3749 net4 _055_ 0.216844f
C3750 _086_ FILLER_0_7_104/a_932_472# 0.001786f
C3751 FILLER_0_11_142/a_124_375# cal_count\[3\] 0.010782f
C3752 FILLER_0_22_177/a_124_375# mask\[6\] 0.002672f
C3753 _098_ _434_/a_2248_156# 0.016991f
C3754 FILLER_0_18_107/a_2276_472# _137_ 0.001752f
C3755 _089_ FILLER_0_5_198/a_36_472# 0.001314f
C3756 _053_ FILLER_0_6_79/a_124_375# 0.003818f
C3757 cal_itt\[3\] _078_ 0.024443f
C3758 FILLER_0_14_91/a_484_472# _136_ 0.038919f
C3759 net7 vss 0.117948f
C3760 net79 FILLER_0_12_236/a_36_472# 0.009225f
C3761 output31/a_224_472# _289_/a_36_472# 0.00101f
C3762 net69 FILLER_0_3_54/a_124_375# 0.004245f
C3763 FILLER_0_15_142/a_572_375# net53 0.021481f
C3764 net81 _060_ 0.019654f
C3765 net16 trim_val\[2\] 0.124462f
C3766 FILLER_0_4_49/a_36_472# net66 0.012791f
C3767 output13/a_224_472# _037_ 0.019694f
C3768 ctln[6] _387_/a_36_113# 0.007687f
C3769 _140_ FILLER_0_22_128/a_2812_375# 0.003154f
C3770 net52 FILLER_0_3_78/a_484_472# 0.003143f
C3771 _108_ _107_ 0.018045f
C3772 en_co_clk fanout55/a_36_160# 0.041263f
C3773 net35 _435_/a_2248_156# 0.001854f
C3774 _068_ net23 0.432092f
C3775 net68 _167_ 0.001302f
C3776 _257_/a_36_472# _122_ 0.007741f
C3777 FILLER_0_2_177/a_124_375# net22 0.001318f
C3778 net49 FILLER_0_3_78/a_484_472# 0.048729f
C3779 FILLER_0_17_161/a_124_375# vss 0.00824f
C3780 FILLER_0_17_161/a_36_472# vdd 0.006972f
C3781 _125_ _135_ 0.001926f
C3782 _043_ net22 0.041447f
C3783 _413_/a_1000_472# net65 0.02866f
C3784 _320_/a_1792_472# vdd 0.001113f
C3785 net15 _447_/a_2248_156# 0.01843f
C3786 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_124_375# 0.012552f
C3787 output35/a_224_472# net22 0.028095f
C3788 net26 net72 0.868238f
C3789 _431_/a_2665_112# _137_ 0.010924f
C3790 _098_ _202_/a_36_160# 0.006831f
C3791 cal_count\[2\] vdd 0.932907f
C3792 _235_/a_67_603# net68 0.027525f
C3793 result[7] _421_/a_1308_423# 0.022204f
C3794 net34 _049_ 0.048403f
C3795 FILLER_0_3_172/a_3172_472# net65 0.001777f
C3796 _005_ _099_ 0.001603f
C3797 _127_ net74 0.0588f
C3798 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_124_375# 0.012001f
C3799 _057_ _128_ 0.036548f
C3800 FILLER_0_9_28/a_124_375# net40 0.047331f
C3801 _013_ _424_/a_36_151# 0.012928f
C3802 _095_ FILLER_0_14_107/a_572_375# 0.01418f
C3803 net72 FILLER_0_12_50/a_124_375# 0.011077f
C3804 net19 _416_/a_2248_156# 0.024466f
C3805 _420_/a_448_472# vdd 0.010071f
C3806 _420_/a_36_151# vss 0.043027f
C3807 net4 FILLER_0_12_220/a_572_375# 0.019052f
C3808 input3/a_36_113# vdd 0.117445f
C3809 _057_ _311_/a_692_473# 0.002083f
C3810 FILLER_0_19_47/a_572_375# _052_ 0.020156f
C3811 FILLER_0_21_133/a_124_375# _433_/a_36_151# 0.059049f
C3812 FILLER_0_4_49/a_572_375# FILLER_0_3_54/a_36_472# 0.001597f
C3813 _228_/a_36_68# _060_ 0.016962f
C3814 net61 fanout78/a_36_113# 0.056484f
C3815 FILLER_0_19_28/a_484_472# vdd 0.010504f
C3816 ctln[1] _411_/a_36_151# 0.018351f
C3817 net47 _365_/a_244_472# 0.001431f
C3818 trimb[1] FILLER_0_20_2/a_36_472# 0.003628f
C3819 _446_/a_1204_472# net66 0.001885f
C3820 net76 vdd 1.272072f
C3821 FILLER_0_24_130/a_36_472# ctlp[7] 0.012298f
C3822 vss _450_/a_36_151# 0.02803f
C3823 vdd _450_/a_448_472# 0.011591f
C3824 cal_count\[3\] _373_/a_1060_68# 0.00165f
C3825 _431_/a_2560_156# net36 0.001858f
C3826 ctln[3] cal_itt\[0\] 0.002081f
C3827 trim_mask\[1\] FILLER_0_4_91/a_484_472# 0.002806f
C3828 _423_/a_2248_156# vss 0.010039f
C3829 _423_/a_2665_112# vdd 0.022696f
C3830 FILLER_0_16_57/a_1380_472# net55 0.002219f
C3831 net69 net23 0.064573f
C3832 _104_ output34/a_224_472# 0.112239f
C3833 FILLER_0_16_89/a_36_472# vss 0.001289f
C3834 FILLER_0_24_96/a_36_472# net24 0.028193f
C3835 cal_count\[3\] _171_ 0.00961f
C3836 net20 net76 0.021613f
C3837 _076_ FILLER_0_8_156/a_124_375# 0.0062f
C3838 _070_ FILLER_0_8_156/a_36_472# 0.001338f
C3839 FILLER_0_4_197/a_1468_375# FILLER_0_4_213/a_36_472# 0.086743f
C3840 FILLER_0_20_193/a_124_375# _098_ 0.009717f
C3841 _062_ _163_ 0.001206f
C3842 _414_/a_448_472# _081_ 0.024533f
C3843 FILLER_0_16_154/a_124_375# vdd 0.00439f
C3844 _253_/a_672_68# _074_ 0.001857f
C3845 FILLER_0_14_91/a_484_472# net53 0.00544f
C3846 _150_ vdd 0.05295f
C3847 FILLER_0_4_49/a_572_375# _164_ 0.005532f
C3848 _440_/a_36_151# FILLER_0_6_47/a_2724_472# 0.001653f
C3849 fanout80/a_36_113# mask\[0\] 0.002212f
C3850 FILLER_0_17_72/a_3172_472# vdd 0.002712f
C3851 net22 _435_/a_2248_156# 0.003453f
C3852 _431_/a_2248_156# vdd 0.00968f
C3853 _079_ net8 0.001928f
C3854 FILLER_0_5_198/a_124_375# vdd 0.010749f
C3855 FILLER_0_22_86/a_1020_375# net14 0.047331f
C3856 _419_/a_1308_423# vdd 0.007543f
C3857 _185_ net40 0.048742f
C3858 _132_ FILLER_0_18_107/a_1380_472# 0.034976f
C3859 _035_ _160_ 0.120469f
C3860 mask\[0\] cal_count\[3\] 0.002612f
C3861 FILLER_0_5_117/a_124_375# _119_ 0.002747f
C3862 _116_ _228_/a_36_68# 0.013091f
C3863 ctln[5] _448_/a_1000_472# 0.007584f
C3864 _152_ net23 0.001895f
C3865 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3172_472# 0.026657f
C3866 output20/a_224_472# _422_/a_1308_423# 0.005632f
C3867 FILLER_0_2_177/a_124_375# vdd 0.019296f
C3868 _372_/a_358_69# _070_ 0.001293f
C3869 net74 FILLER_0_13_72/a_36_472# 0.007448f
C3870 net44 _190_/a_36_160# 0.015628f
C3871 net20 _419_/a_1308_423# 0.022245f
C3872 _043_ vdd 0.827689f
C3873 net53 state\[1\] 0.00554f
C3874 output15/a_224_472# ctln[8] 0.079231f
C3875 trim_val\[4\] FILLER_0_3_172/a_572_375# 0.001076f
C3876 output35/a_224_472# vdd 0.064053f
C3877 mask\[3\] FILLER_0_18_177/a_1828_472# 0.004274f
C3878 _072_ FILLER_0_12_220/a_484_472# 0.028355f
C3879 net4 FILLER_0_12_236/a_484_472# 0.014212f
C3880 net70 FILLER_0_14_99/a_124_375# 0.002922f
C3881 _016_ _131_ 0.017461f
C3882 net62 FILLER_0_13_212/a_124_375# 0.001597f
C3883 FILLER_0_6_90/a_484_472# _163_ 0.011711f
C3884 _058_ _055_ 0.070216f
C3885 _186_ vss 0.0718f
C3886 net20 _043_ 0.094689f
C3887 _178_ _186_ 0.020123f
C3888 _020_ net73 0.057454f
C3889 _369_/a_36_68# _157_ 0.068266f
C3890 net4 FILLER_0_3_221/a_124_375# 0.015788f
C3891 FILLER_0_4_49/a_484_472# net47 0.002964f
C3892 mask\[7\] _435_/a_796_472# 0.009587f
C3893 _394_/a_56_524# cal_count\[1\] 0.022487f
C3894 net55 _052_ 0.095046f
C3895 FILLER_0_9_28/a_2724_472# _453_/a_36_151# 0.013806f
C3896 mask\[3\] _094_ 0.00554f
C3897 mask\[3\] FILLER_0_17_218/a_572_375# 0.015907f
C3898 output31/a_224_472# net19 0.072666f
C3899 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1468_375# 0.086635f
C3900 _131_ FILLER_0_14_123/a_124_375# 0.016964f
C3901 _272_/a_36_472# _087_ 0.048282f
C3902 _059_ _242_/a_36_160# 0.001942f
C3903 _062_ _117_ 0.042699f
C3904 _091_ FILLER_0_13_228/a_124_375# 0.001657f
C3905 net16 _174_ 0.022224f
C3906 net22 FILLER_0_18_209/a_484_472# 0.005297f
C3907 net68 vdd 1.026897f
C3908 cal_itt\[1\] net8 0.040042f
C3909 net63 _275_/a_224_472# 0.002538f
C3910 _176_ _174_ 0.00677f
C3911 mask\[5\] FILLER_0_19_171/a_484_472# 0.007647f
C3912 _093_ net30 0.001859f
C3913 _026_ vdd 0.15542f
C3914 net4 state\[1\] 0.010195f
C3915 net23 FILLER_0_22_128/a_2276_472# 0.011079f
C3916 FILLER_0_3_2/a_36_472# _446_/a_36_151# 0.004032f
C3917 _426_/a_448_472# calibrate 0.002745f
C3918 FILLER_0_18_139/a_1020_375# vss 0.032606f
C3919 FILLER_0_18_139/a_1468_375# vdd 0.015542f
C3920 _255_/a_224_552# _058_ 0.06267f
C3921 FILLER_0_9_72/a_36_472# _439_/a_36_151# 0.001723f
C3922 FILLER_0_21_125/a_124_375# mask\[7\] 0.00145f
C3923 FILLER_0_15_282/a_124_375# net18 0.048284f
C3924 _036_ _168_ 0.01699f
C3925 FILLER_0_15_282/a_484_472# output30/a_224_472# 0.001711f
C3926 net19 _419_/a_1000_472# 0.012949f
C3927 FILLER_0_10_256/a_36_472# _426_/a_36_151# 0.059238f
C3928 FILLER_0_12_28/a_36_472# cal_count\[0\] 0.001662f
C3929 net15 net51 0.191328f
C3930 FILLER_0_18_177/a_3260_375# _202_/a_36_160# 0.001948f
C3931 vdd _156_ 0.178622f
C3932 _426_/a_36_151# net64 0.022056f
C3933 _063_ _444_/a_36_151# 0.030369f
C3934 FILLER_0_14_81/a_36_472# _175_ 0.076977f
C3935 _392_/a_36_68# FILLER_0_12_50/a_36_472# 0.002811f
C3936 _439_/a_36_151# _453_/a_2248_156# 0.001082f
C3937 FILLER_0_12_136/a_1380_472# FILLER_0_13_142/a_572_375# 0.001684f
C3938 FILLER_0_17_200/a_572_375# FILLER_0_18_177/a_3172_472# 0.001597f
C3939 output25/a_224_472# _214_/a_36_160# 0.027335f
C3940 FILLER_0_1_204/a_36_472# net11 0.014707f
C3941 _140_ mask\[6\] 0.605898f
C3942 mask\[8\] _140_ 0.003375f
C3943 _440_/a_2665_112# _160_ 0.008418f
C3944 net71 _437_/a_2248_156# 0.025557f
C3945 net57 _068_ 0.029812f
C3946 _435_/a_2248_156# vdd 0.00571f
C3947 _112_ _083_ 0.003571f
C3948 _136_ _451_/a_1353_112# 0.058703f
C3949 net38 _444_/a_1204_472# 0.018432f
C3950 FILLER_0_17_72/a_2812_375# net14 0.018463f
C3951 _352_/a_49_472# _436_/a_36_151# 0.005127f
C3952 _074_ FILLER_0_3_221/a_1380_472# 0.001341f
C3953 result[4] net61 0.023257f
C3954 _256_/a_244_497# calibrate 0.002421f
C3955 _103_ _418_/a_2560_156# 0.002179f
C3956 fanout65/a_36_113# vdd 0.10473f
C3957 _443_/a_36_151# net13 0.001896f
C3958 _443_/a_1308_423# net23 0.034115f
C3959 FILLER_0_8_2/a_36_472# net40 0.002477f
C3960 output28/a_224_472# vss -0.0033f
C3961 FILLER_0_18_76/a_484_472# vss 0.005065f
C3962 _149_ _437_/a_36_151# 0.037766f
C3963 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_1020_375# 0.026339f
C3964 _392_/a_244_472# cal_count\[0\] 0.003287f
C3965 _070_ _370_/a_124_24# 0.00219f
C3966 _029_ net14 0.042032f
C3967 net67 vdd 0.638702f
C3968 ctln[5] FILLER_0_0_198/a_36_472# 0.012298f
C3969 FILLER_0_10_78/a_36_472# _453_/a_2665_112# 0.007491f
C3970 _426_/a_2665_112# net4 0.011288f
C3971 FILLER_0_11_124/a_124_375# _120_ 0.012164f
C3972 output8/a_224_472# _080_ 0.001971f
C3973 FILLER_0_21_125/a_484_472# vdd 0.002728f
C3974 FILLER_0_21_125/a_36_472# vss 0.00143f
C3975 ctln[4] vdd 0.210384f
C3976 trim_val\[4\] _443_/a_2248_156# 0.050943f
C3977 output39/a_224_472# trim[1] 0.061797f
C3978 _077_ FILLER_0_12_50/a_36_472# 0.177624f
C3979 _020_ _131_ 0.011012f
C3980 _114_ FILLER_0_10_78/a_1380_472# 0.011079f
C3981 net54 FILLER_0_18_107/a_36_472# 0.002116f
C3982 _126_ _389_/a_36_148# 0.007813f
C3983 _029_ _164_ 0.031781f
C3984 FILLER_0_8_107/a_36_472# net14 0.001596f
C3985 FILLER_0_11_64/a_36_472# vdd 0.015144f
C3986 FILLER_0_11_64/a_124_375# vss 0.021069f
C3987 _070_ _247_/a_36_160# 0.0169f
C3988 output13/a_224_472# _448_/a_2248_156# 0.009013f
C3989 FILLER_0_12_236/a_124_375# vdd 0.005169f
C3990 _010_ _009_ 0.030637f
C3991 net20 ctln[4] 0.00225f
C3992 net38 _064_ 0.02996f
C3993 net34 output34/a_224_472# 0.031833f
C3994 _132_ _428_/a_448_472# 0.034825f
C3995 _335_/a_49_472# FILLER_0_15_180/a_572_375# 0.001126f
C3996 FILLER_0_8_138/a_124_375# _076_ 0.031436f
C3997 _077_ _114_ 0.047702f
C3998 FILLER_0_14_91/a_124_375# vdd -0.010114f
C3999 FILLER_0_15_282/a_572_375# _417_/a_36_151# 0.001597f
C4000 FILLER_0_7_104/a_1020_375# _062_ 0.003073f
C4001 net63 FILLER_0_22_177/a_572_375# 0.001597f
C4002 FILLER_0_21_133/a_36_472# mask\[7\] 0.003404f
C4003 _442_/a_36_151# _031_ 0.013852f
C4004 _445_/a_36_151# vss 0.009726f
C4005 _445_/a_448_472# vdd 0.007946f
C4006 FILLER_0_18_209/a_484_472# vdd 0.00367f
C4007 FILLER_0_18_209/a_36_472# vss 0.005442f
C4008 FILLER_0_21_28/a_484_472# vdd 0.011209f
C4009 FILLER_0_18_171/a_124_375# net80 0.024341f
C4010 net50 FILLER_0_2_93/a_124_375# 0.007132f
C4011 net52 FILLER_0_2_93/a_36_472# 0.009026f
C4012 FILLER_0_7_162/a_36_472# _062_ 0.016683f
C4013 _187_ _453_/a_36_151# 0.001829f
C4014 _423_/a_36_151# _012_ 0.021631f
C4015 _104_ output21/a_224_472# 0.002459f
C4016 _052_ _216_/a_67_603# 0.006658f
C4017 FILLER_0_13_65/a_124_375# vdd 0.011301f
C4018 _328_/a_36_113# _114_ 0.058671f
C4019 output12/a_224_472# net12 0.007193f
C4020 _028_ FILLER_0_7_72/a_1468_375# 0.003785f
C4021 output15/a_224_472# fanout50/a_36_160# 0.003531f
C4022 _000_ vdd 0.215988f
C4023 FILLER_0_8_127/a_124_375# _125_ 0.003105f
C4024 _144_ net71 0.039862f
C4025 net38 net42 0.012245f
C4026 _161_ FILLER_0_6_177/a_572_375# 0.004064f
C4027 _162_ FILLER_0_6_177/a_36_472# 0.001723f
C4028 _091_ _430_/a_2560_156# 0.047345f
C4029 FILLER_0_2_93/a_36_472# net49 0.001451f
C4030 net63 _435_/a_2560_156# 0.023868f
C4031 net36 _451_/a_836_156# 0.007104f
C4032 FILLER_0_8_239/a_124_375# calibrate 0.008393f
C4033 output42/a_224_472# net17 0.047757f
C4034 output36/a_224_472# net62 0.317201f
C4035 _427_/a_1308_423# net23 0.004863f
C4036 net52 trim_mask\[2\] 0.036196f
C4037 net76 FILLER_0_5_198/a_572_375# 0.006974f
C4038 net68 fanout67/a_36_160# 0.02648f
C4039 FILLER_0_12_50/a_36_472# _120_ 0.005447f
C4040 _086_ _153_ 0.017325f
C4041 FILLER_0_13_212/a_572_375# _248_/a_36_68# 0.030745f
C4042 net47 FILLER_0_6_37/a_36_472# 0.001161f
C4043 net62 net30 0.339141f
C4044 ctln[5] net11 0.004569f
C4045 net20 _000_ 0.159624f
C4046 mask\[4\] _346_/a_665_69# 0.001125f
C4047 _068_ _315_/a_244_497# 0.004768f
C4048 _186_ _184_ 0.047995f
C4049 _115_ _322_/a_692_472# 0.00171f
C4050 mask\[5\] FILLER_0_20_177/a_1380_472# 0.016114f
C4051 FILLER_0_20_107/a_36_472# vss 0.004557f
C4052 output24/a_224_472# net24 0.005559f
C4053 trim_mask\[2\] net49 0.041781f
C4054 _064_ net66 0.304028f
C4055 net76 FILLER_0_2_177/a_572_375# 0.053951f
C4056 output28/a_224_472# _416_/a_2248_156# 0.023576f
C4057 result[1] _416_/a_1308_423# 0.002597f
C4058 _009_ FILLER_0_23_282/a_36_472# 0.005974f
C4059 _114_ _120_ 0.334426f
C4060 net24 vss 0.172755f
C4061 output14/a_224_472# _442_/a_2248_156# 0.001723f
C4062 _112_ _425_/a_36_151# 0.032941f
C4063 net16 _450_/a_3129_107# 0.064714f
C4064 FILLER_0_18_2/a_932_472# net38 0.020589f
C4065 net72 _180_ 0.040135f
C4066 FILLER_0_16_57/a_124_375# _176_ 0.015872f
C4067 _131_ FILLER_0_18_37/a_1380_472# 0.035078f
C4068 net53 _451_/a_1353_112# 0.028324f
C4069 result[6] _421_/a_796_472# 0.004697f
C4070 _091_ FILLER_0_18_171/a_36_472# 0.00395f
C4071 _131_ FILLER_0_17_56/a_124_375# 0.001609f
C4072 _065_ output16/a_224_472# 0.049052f
C4073 _239_/a_36_160# net16 0.003137f
C4074 _114_ FILLER_0_13_142/a_1020_375# 0.001964f
C4075 _425_/a_2665_112# net37 0.008519f
C4076 _128_ FILLER_0_10_214/a_36_472# 0.00186f
C4077 output21/a_224_472# mask\[5\] 0.009585f
C4078 FILLER_0_5_128/a_572_375# _081_ 0.023853f
C4079 _028_ vdd 0.626868f
C4080 net55 net40 0.043962f
C4081 FILLER_0_16_107/a_572_375# net36 0.001706f
C4082 trim[4] _221_/a_36_160# 0.002685f
C4083 net7 output41/a_224_472# 0.019483f
C4084 _182_ cal_count\[1\] 0.166348f
C4085 result[0] FILLER_0_9_290/a_36_472# 0.020103f
C4086 _017_ _131_ 0.005879f
C4087 FILLER_0_14_81/a_124_375# vdd 0.023163f
C4088 _140_ _352_/a_665_69# 0.001363f
C4089 net60 _418_/a_36_151# 0.016348f
C4090 _141_ _145_ 0.094128f
C4091 result[2] vdd 0.18482f
C4092 _432_/a_2248_156# _139_ 0.002904f
C4093 _426_/a_1000_472# vdd 0.007031f
C4094 _303_/a_36_472# _098_ 0.021192f
C4095 _140_ _433_/a_2248_156# 0.003337f
C4096 net46 FILLER_0_21_28/a_36_472# 0.051176f
C4097 net82 _370_/a_124_24# 0.001011f
C4098 FILLER_0_9_290/a_124_375# vdd 0.028723f
C4099 mask\[4\] mask\[3\] 1.118454f
C4100 FILLER_0_12_220/a_932_472# _060_ 0.002471f
C4101 _413_/a_448_472# net76 0.029504f
C4102 output38/a_224_472# net38 0.018882f
C4103 fanout67/a_36_160# net67 0.017633f
C4104 _176_ FILLER_0_15_59/a_124_375# 0.007169f
C4105 _065_ _447_/a_2665_112# 0.034757f
C4106 _163_ net14 0.040169f
C4107 _021_ _141_ 0.047816f
C4108 _132_ FILLER_0_17_104/a_1020_375# 0.009251f
C4109 _063_ vss 0.157186f
C4110 output27/a_224_472# FILLER_0_9_282/a_124_375# 0.029138f
C4111 _427_/a_796_472# net74 0.020124f
C4112 FILLER_0_3_204/a_124_375# net65 0.003831f
C4113 net55 FILLER_0_17_38/a_572_375# 0.007646f
C4114 net62 _417_/a_36_151# 0.044051f
C4115 _009_ _299_/a_36_472# 0.006927f
C4116 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_124_375# 0.012552f
C4117 _259_/a_455_68# net20 0.001427f
C4118 net64 FILLER_0_8_247/a_1380_472# 0.001021f
C4119 ctlp[5] ctlp[4] 0.001257f
C4120 output15/a_224_472# net14 0.003312f
C4121 net17 FILLER_0_12_28/a_36_472# 0.012286f
C4122 ctln[0] vss 0.125714f
C4123 _411_/a_2665_112# vdd 0.026095f
C4124 _163_ _164_ 0.021311f
C4125 net81 net2 1.204674f
C4126 net17 net40 1.095167f
C4127 _225_/a_36_160# vss 0.003244f
C4128 FILLER_0_6_47/a_1468_375# vss 0.003462f
C4129 FILLER_0_6_47/a_1916_375# vdd -0.014642f
C4130 _057_ _176_ 0.001304f
C4131 _069_ _043_ 0.04044f
C4132 output8/a_224_472# vss 0.076244f
C4133 net50 _054_ 0.131493f
C4134 _231_/a_244_68# _059_ 0.004384f
C4135 _431_/a_448_472# _093_ 0.002095f
C4136 FILLER_0_13_290/a_36_472# output30/a_224_472# 0.0323f
C4137 _076_ FILLER_0_5_148/a_36_472# 0.011563f
C4138 result[8] FILLER_0_21_206/a_36_472# 0.001292f
C4139 mask\[9\] FILLER_0_19_111/a_484_472# 0.041744f
C4140 _193_/a_36_160# result[3] 0.002218f
C4141 output15/a_224_472# _164_ 0.031363f
C4142 FILLER_0_12_124/a_36_472# _131_ 0.028609f
C4143 vss FILLER_0_12_196/a_36_472# 0.003551f
C4144 net4 _223_/a_36_160# 0.020711f
C4145 _412_/a_448_472# _001_ 0.01124f
C4146 FILLER_0_16_73/a_484_472# _176_ 0.010681f
C4147 _128_ _161_ 0.027657f
C4148 _428_/a_2560_156# net53 0.002265f
C4149 FILLER_0_16_73/a_124_375# net15 0.005202f
C4150 _369_/a_36_68# _158_ 0.042315f
C4151 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_572_375# 0.086635f
C4152 _050_ _436_/a_1000_472# 0.02064f
C4153 output38/a_224_472# net66 0.148811f
C4154 _186_ _095_ 0.042856f
C4155 vss FILLER_0_6_231/a_572_375# 0.057794f
C4156 vdd FILLER_0_6_231/a_36_472# 0.014642f
C4157 net50 vss 1.178736f
C4158 net74 _118_ 0.060991f
C4159 _421_/a_36_151# vdd -0.053849f
C4160 _114_ state\[2\] 0.528838f
C4161 _128_ _129_ 0.029628f
C4162 net67 _450_/a_1353_112# 0.025358f
C4163 FILLER_0_18_107/a_2724_472# vss 0.003148f
C4164 FILLER_0_18_107/a_3172_472# vdd 0.004296f
C4165 _136_ FILLER_0_15_180/a_572_375# 0.001571f
C4166 net79 _070_ 0.009715f
C4167 FILLER_0_7_195/a_36_472# cal_itt\[3\] 0.070665f
C4168 output33/a_224_472# output19/a_224_472# 0.115114f
C4169 _424_/a_2248_156# vdd -0.005751f
C4170 FILLER_0_1_192/a_124_375# vss 0.049811f
C4171 FILLER_0_1_192/a_36_472# vdd 0.011806f
C4172 net26 FILLER_0_23_44/a_124_375# 0.007775f
C4173 _320_/a_1120_472# state\[1\] 0.001998f
C4174 _265_/a_224_472# net59 0.001052f
C4175 net20 FILLER_0_6_231/a_36_472# 0.045553f
C4176 net57 _113_ 0.012056f
C4177 _432_/a_448_472# _093_ 0.048289f
C4178 _027_ FILLER_0_18_76/a_484_472# 0.00705f
C4179 state\[0\] _090_ 0.003121f
C4180 _274_/a_36_68# vss 0.052669f
C4181 net52 _441_/a_2560_156# 0.004721f
C4182 net50 _441_/a_2248_156# 0.027849f
C4183 mask\[4\] FILLER_0_17_200/a_36_472# 0.001242f
C4184 _035_ FILLER_0_4_49/a_124_375# 0.00215f
C4185 net15 net47 0.035839f
C4186 FILLER_0_7_72/a_36_472# net50 0.011974f
C4187 net81 valid 0.11798f
C4188 net34 _422_/a_1204_472# 0.001029f
C4189 FILLER_0_16_57/a_1468_375# net15 0.012909f
C4190 _029_ _153_ 0.023421f
C4191 FILLER_0_7_72/a_3172_472# vss 0.002425f
C4192 _417_/a_2560_156# net30 0.049334f
C4193 _049_ FILLER_0_22_128/a_2812_375# 0.001905f
C4194 FILLER_0_12_136/a_36_472# vss 0.003185f
C4195 FILLER_0_12_136/a_484_472# vdd 0.005304f
C4196 _258_/a_36_160# _073_ 0.079254f
C4197 _449_/a_36_151# _043_ 0.001572f
C4198 _340_/a_36_160# FILLER_0_20_169/a_124_375# 0.005494f
C4199 output35/a_224_472# _435_/a_2665_112# 0.008469f
C4200 output32/a_224_472# result[9] 0.047198f
C4201 _130_ _120_ 0.014675f
C4202 net15 _012_ 0.043755f
C4203 _074_ FILLER_0_6_177/a_36_472# 0.045576f
C4204 _256_/a_1612_497# net4 0.002497f
C4205 FILLER_0_19_134/a_36_472# _145_ 0.080913f
C4206 FILLER_0_5_72/a_1020_375# vdd 0.009501f
C4207 FILLER_0_5_72/a_572_375# vss 0.006023f
C4208 net21 _434_/a_2248_156# 0.001467f
C4209 net41 FILLER_0_21_28/a_572_375# 0.054443f
C4210 net69 FILLER_0_2_111/a_484_472# 0.010567f
C4211 _031_ FILLER_0_2_111/a_1468_375# 0.013595f
C4212 net14 FILLER_0_4_91/a_36_472# 0.005793f
C4213 FILLER_0_6_239/a_36_472# FILLER_0_6_231/a_484_472# 0.013277f
C4214 _420_/a_448_472# net77 0.001276f
C4215 _050_ FILLER_0_22_128/a_124_375# 0.002607f
C4216 net61 _422_/a_2665_112# 0.023601f
C4217 _098_ FILLER_0_19_171/a_572_375# 0.001946f
C4218 FILLER_0_5_54/a_572_375# _029_ 0.00494f
C4219 calibrate FILLER_0_8_156/a_36_472# 0.001283f
C4220 _315_/a_36_68# _121_ 0.031617f
C4221 _122_ FILLER_0_8_156/a_572_375# 0.002572f
C4222 _441_/a_36_151# _440_/a_448_472# 0.002538f
C4223 net16 trim_val\[0\] 0.00463f
C4224 net41 _064_ 0.301777f
C4225 _446_/a_1308_423# net40 0.038281f
C4226 _426_/a_36_151# FILLER_0_8_247/a_572_375# 0.059049f
C4227 _012_ FILLER_0_23_44/a_1380_472# 0.001572f
C4228 vdd _380_/a_224_472# 0.001733f
C4229 _412_/a_2665_112# fanout59/a_36_160# 0.016426f
C4230 FILLER_0_4_177/a_484_472# vss 0.002399f
C4231 _346_/a_49_472# _098_ 0.028579f
C4232 _081_ FILLER_0_5_148/a_36_472# 0.020403f
C4233 FILLER_0_21_150/a_124_375# _433_/a_2665_112# 0.029834f
C4234 FILLER_0_16_255/a_124_375# vdd 0.029925f
C4235 _421_/a_1308_423# net19 0.055838f
C4236 _308_/a_124_24# _439_/a_2248_156# 0.01963f
C4237 _074_ _316_/a_124_24# 0.018608f
C4238 _431_/a_1308_423# _427_/a_36_151# 0.001256f
C4239 net15 FILLER_0_15_59/a_484_472# 0.015199f
C4240 net36 FILLER_0_15_180/a_484_472# 0.00702f
C4241 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_124_375# 0.012001f
C4242 _431_/a_448_472# _136_ 0.064724f
C4243 net39 net47 0.13057f
C4244 _114_ _311_/a_2180_473# 0.00515f
C4245 _253_/a_36_68# _073_ 0.027664f
C4246 net47 net51 0.007412f
C4247 _093_ _046_ 0.061989f
C4248 FILLER_0_7_72/a_1916_375# FILLER_0_6_90/a_36_472# 0.001684f
C4249 _005_ net18 0.073455f
C4250 net16 _445_/a_2248_156# 0.003321f
C4251 net50 FILLER_0_5_88/a_124_375# 0.03181f
C4252 FILLER_0_22_177/a_932_472# _435_/a_36_151# 0.001723f
C4253 _372_/a_3662_472# _122_ 0.002653f
C4254 _035_ _446_/a_796_472# 0.013039f
C4255 net21 _202_/a_36_160# 0.09166f
C4256 FILLER_0_9_28/a_1380_472# net68 0.008573f
C4257 net15 net74 0.05717f
C4258 FILLER_0_15_72/a_484_472# vss 0.010761f
C4259 mask\[4\] FILLER_0_19_155/a_572_375# 0.020261f
C4260 _069_ FILLER_0_18_209/a_484_472# 0.013944f
C4261 _127_ FILLER_0_9_142/a_124_375# 0.005447f
C4262 net43 FILLER_0_20_15/a_36_472# 0.002803f
C4263 net81 FILLER_0_15_212/a_36_472# 0.003945f
C4264 _413_/a_448_472# ctln[4] 0.001072f
C4265 net32 _011_ 0.072502f
C4266 FILLER_0_17_226/a_124_375# _008_ 0.006576f
C4267 FILLER_0_21_150/a_124_375# vdd 0.020581f
C4268 FILLER_0_3_2/a_36_472# vss 0.004076f
C4269 _308_/a_848_380# _114_ 0.005266f
C4270 _326_/a_36_160# _058_ 0.003897f
C4271 _028_ FILLER_0_7_72/a_1380_472# 0.001777f
C4272 _057_ _267_/a_36_472# 0.038568f
C4273 _015_ net64 1.212892f
C4274 net26 vdd 0.487733f
C4275 ctln[7] FILLER_0_0_96/a_124_375# 0.025944f
C4276 net55 FILLER_0_17_56/a_36_472# 0.019193f
C4277 cal_itt\[3\] vss 0.15522f
C4278 _133_ FILLER_0_10_107/a_484_472# 0.001798f
C4279 _293_/a_36_472# output34/a_224_472# 0.001888f
C4280 _128_ _056_ 0.026612f
C4281 _432_/a_448_472# _136_ 0.001892f
C4282 FILLER_0_23_88/a_36_472# net14 0.003077f
C4283 _132_ _093_ 0.105039f
C4284 _431_/a_1000_472# _136_ 0.024253f
C4285 FILLER_0_12_50/a_124_375# vdd 0.039185f
C4286 _093_ FILLER_0_17_72/a_2364_375# 0.010888f
C4287 _061_ _311_/a_66_473# 0.030169f
C4288 _428_/a_1204_472# vdd 0.001231f
C4289 _098_ _433_/a_1204_472# 0.014374f
C4290 _071_ _225_/a_36_160# 0.002808f
C4291 _009_ vss 0.105833f
C4292 FILLER_0_24_96/a_124_375# net24 0.040364f
C4293 valid net2 0.062523f
C4294 _068_ FILLER_0_9_142/a_36_472# 0.009073f
C4295 _394_/a_728_93# vdd 0.006211f
C4296 _394_/a_1336_472# vss 0.040135f
C4297 FILLER_0_4_177/a_572_375# FILLER_0_5_181/a_124_375# 0.05841f
C4298 cal_count\[1\] _040_ 0.019478f
C4299 net41 output38/a_224_472# 0.017358f
C4300 _163_ _153_ 0.243815f
C4301 _449_/a_36_151# FILLER_0_11_64/a_36_472# 0.046516f
C4302 FILLER_0_24_274/a_932_472# FILLER_0_23_282/a_36_472# 0.05841f
C4303 FILLER_0_11_142/a_484_472# net23 0.006988f
C4304 _081_ FILLER_0_6_177/a_36_472# 0.00483f
C4305 _422_/a_1000_472# _009_ 0.007191f
C4306 _408_/a_1336_472# net40 0.020063f
C4307 vss _039_ 0.180364f
C4308 FILLER_0_14_81/a_36_472# _043_ 0.001714f
C4309 FILLER_0_9_28/a_1020_375# net50 0.001512f
C4310 FILLER_0_8_247/a_124_375# FILLER_0_8_239/a_124_375# 0.003732f
C4311 FILLER_0_19_47/a_572_375# FILLER_0_18_53/a_36_472# 0.001684f
C4312 _189_/a_67_603# FILLER_0_13_228/a_36_472# 0.005759f
C4313 FILLER_0_7_72/a_572_375# vdd 0.004039f
C4314 output9/a_224_472# vss 0.007544f
C4315 _128_ _068_ 0.863174f
C4316 _131_ cal_count\[3\] 0.035391f
C4317 _086_ FILLER_0_6_177/a_36_472# 0.064045f
C4318 _016_ _427_/a_448_472# 0.016416f
C4319 net1 _083_ 0.30074f
C4320 FILLER_0_20_177/a_1468_375# _098_ 0.012889f
C4321 output46/a_224_472# net43 0.10562f
C4322 FILLER_0_13_65/a_124_375# _449_/a_36_151# 0.059049f
C4323 net62 fanout78/a_36_113# 0.014177f
C4324 net55 _452_/a_1040_527# 0.021721f
C4325 _431_/a_448_472# net53 0.002087f
C4326 FILLER_0_5_164/a_572_375# _386_/a_848_380# 0.001121f
C4327 FILLER_0_9_28/a_3172_472# FILLER_0_9_60/a_36_472# 0.013276f
C4328 _052_ FILLER_0_18_61/a_124_375# 0.006877f
C4329 result[9] _094_ 0.03984f
C4330 _068_ _311_/a_692_473# 0.002377f
C4331 _072_ _061_ 0.448032f
C4332 _092_ FILLER_0_17_218/a_124_375# 0.020704f
C4333 mask\[5\] _346_/a_257_69# 0.001764f
C4334 _412_/a_2665_112# net5 0.042084f
C4335 _411_/a_36_151# net65 0.001415f
C4336 FILLER_0_9_28/a_36_472# FILLER_0_10_28/a_36_472# 0.05841f
C4337 _072_ _311_/a_66_473# 0.031716f
C4338 _427_/a_36_151# FILLER_0_14_123/a_36_472# 0.004032f
C4339 _081_ _316_/a_124_24# 0.011421f
C4340 _302_/a_224_472# _012_ 0.002675f
C4341 _143_ _093_ 0.003295f
C4342 net80 FILLER_0_16_154/a_1468_375# 0.013593f
C4343 _062_ net37 0.082701f
C4344 _173_ net51 0.016607f
C4345 _274_/a_716_497# net64 0.007904f
C4346 trim_mask\[1\] FILLER_0_6_47/a_1380_472# 0.006166f
C4347 _009_ _107_ 0.027726f
C4348 FILLER_0_18_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001684f
C4349 _432_/a_36_151# FILLER_0_15_180/a_36_472# 0.002018f
C4350 output10/a_224_472# _411_/a_2248_156# 0.019736f
C4351 _102_ _099_ 0.151018f
C4352 _093_ _356_/a_36_472# 0.009235f
C4353 _065_ net66 0.003956f
C4354 FILLER_0_15_116/a_36_472# _136_ 0.003818f
C4355 FILLER_0_13_228/a_124_375# vdd -0.007362f
C4356 _000_ cal_itt\[2\] 0.042235f
C4357 FILLER_0_5_128/a_572_375# _163_ 0.007391f
C4358 FILLER_0_10_247/a_124_375# _100_ 0.001804f
C4359 _079_ _073_ 0.234533f
C4360 _091_ FILLER_0_19_171/a_36_472# 0.029168f
C4361 _322_/a_848_380# vss 0.026127f
C4362 net18 _416_/a_448_472# 0.05521f
C4363 mask\[5\] _204_/a_67_603# 0.023791f
C4364 net75 _425_/a_448_472# 0.038993f
C4365 _095_ _225_/a_36_160# 0.001084f
C4366 FILLER_0_15_10/a_124_375# vdd 0.021578f
C4367 FILLER_0_2_101/a_36_472# vss 0.004743f
C4368 FILLER_0_4_144/a_36_472# vdd 0.004289f
C4369 FILLER_0_4_144/a_572_375# vss 0.072463f
C4370 fanout61/a_36_113# FILLER_0_21_286/a_572_375# 0.015816f
C4371 net20 FILLER_0_13_228/a_124_375# 0.047331f
C4372 _126_ FILLER_0_12_196/a_124_375# 0.001392f
C4373 net35 FILLER_0_22_128/a_36_472# 0.00784f
C4374 _102_ _419_/a_2248_156# 0.001679f
C4375 net17 _452_/a_1040_527# 0.034254f
C4376 _285_/a_36_472# _094_ 0.045394f
C4377 _411_/a_1000_472# vss 0.002964f
C4378 fanout79/a_36_160# _060_ 0.005814f
C4379 _247_/a_36_160# net21 0.002254f
C4380 net75 _082_ 0.417366f
C4381 net75 net82 0.214597f
C4382 _265_/a_244_68# vss 0.009604f
C4383 FILLER_0_18_2/a_1020_375# net55 0.003942f
C4384 _281_/a_234_472# _097_ 0.004169f
C4385 FILLER_0_18_139/a_932_472# FILLER_0_17_142/a_484_472# 0.026657f
C4386 net60 _419_/a_1204_472# 0.023544f
C4387 net61 _419_/a_2665_112# 0.022394f
C4388 _132_ _136_ 0.034253f
C4389 _413_/a_36_151# vdd 0.130213f
C4390 _013_ net36 0.032392f
C4391 net47 clkc 0.002956f
C4392 net54 FILLER_0_22_128/a_572_375# 0.048634f
C4393 FILLER_0_17_104/a_932_472# vdd 0.020019f
C4394 _444_/a_1308_423# net40 0.043396f
C4395 _070_ FILLER_0_9_105/a_124_375# 0.017687f
C4396 _013_ FILLER_0_18_37/a_932_472# 0.010651f
C4397 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_124_375# 0.003732f
C4398 FILLER_0_17_72/a_2364_375# _136_ 0.047331f
C4399 FILLER_0_16_89/a_36_472# _451_/a_448_472# 0.011974f
C4400 output9/a_224_472# fanout76/a_36_160# 0.016067f
C4401 result[9] net78 0.015761f
C4402 FILLER_0_8_24/a_572_375# net40 0.038492f
C4403 FILLER_0_7_72/a_1020_375# vdd 0.004039f
C4404 FILLER_0_8_127/a_36_472# _062_ 0.01783f
C4405 _078_ vdd 0.181583f
C4406 net63 _098_ 0.055686f
C4407 mask\[4\] FILLER_0_19_187/a_36_472# 0.004669f
C4408 FILLER_0_18_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001597f
C4409 _374_/a_36_68# _058_ 0.010442f
C4410 FILLER_0_4_197/a_572_375# net22 0.016547f
C4411 _073_ cal_itt\[1\] 0.058541f
C4412 net55 FILLER_0_18_53/a_36_472# 0.00953f
C4413 net50 _036_ 0.002727f
C4414 net63 _434_/a_3041_156# 0.001449f
C4415 FILLER_0_23_290/a_36_472# vss 0.0074f
C4416 output32/a_224_472# _094_ 0.005545f
C4417 _432_/a_1204_472# net80 0.009362f
C4418 mask\[2\] FILLER_0_15_212/a_1380_472# 0.001225f
C4419 net20 _078_ 0.105266f
C4420 FILLER_0_16_89/a_1020_375# _131_ 0.015706f
C4421 _115_ FILLER_0_10_94/a_124_375# 0.010311f
C4422 FILLER_0_12_136/a_1468_375# _126_ 0.012732f
C4423 net80 FILLER_0_22_177/a_1020_375# 0.00258f
C4424 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3172_472# 0.013277f
C4425 trim[4] net67 0.06366f
C4426 _431_/a_36_151# _132_ 0.051016f
C4427 net10 vss 0.324553f
C4428 output7/a_224_472# trim[3] 0.103375f
C4429 FILLER_0_8_107/a_124_375# _219_/a_36_160# 0.002515f
C4430 trim_mask\[2\] net40 0.401672f
C4431 _415_/a_2665_112# FILLER_0_9_290/a_124_375# 0.001597f
C4432 _413_/a_448_472# FILLER_0_1_192/a_36_472# 0.001462f
C4433 output25/a_224_472# net25 0.179738f
C4434 FILLER_0_20_177/a_124_375# FILLER_0_20_169/a_124_375# 0.003732f
C4435 _050_ FILLER_0_22_107/a_36_472# 0.001098f
C4436 FILLER_0_20_193/a_484_472# vdd 0.00749f
C4437 FILLER_0_20_193/a_36_472# vss 0.001978f
C4438 FILLER_0_16_73/a_124_375# FILLER_0_16_57/a_1468_375# 0.012222f
C4439 ctln[0] output41/a_224_472# 0.001583f
C4440 FILLER_0_17_72/a_1828_472# _131_ 0.004882f
C4441 net16 _034_ 0.096088f
C4442 _106_ ctlp[1] 0.002631f
C4443 _420_/a_796_472# _009_ 0.012395f
C4444 FILLER_0_19_111/a_36_472# net14 0.00143f
C4445 net34 FILLER_0_22_177/a_1020_375# 0.006974f
C4446 _119_ cal_itt\[3\] 0.010152f
C4447 net72 vss 0.472104f
C4448 FILLER_0_15_116/a_36_472# net53 0.005099f
C4449 _413_/a_36_151# FILLER_0_3_172/a_2812_375# 0.059049f
C4450 net68 FILLER_0_8_37/a_124_375# 0.004818f
C4451 _133_ _058_ 0.092697f
C4452 _178_ net72 0.007093f
C4453 _136_ _356_/a_36_472# 0.004667f
C4454 _101_ _094_ 0.304499f
C4455 FILLER_0_18_107/a_3260_375# FILLER_0_19_134/a_124_375# 0.026339f
C4456 FILLER_0_5_54/a_484_472# vss 0.001929f
C4457 FILLER_0_5_54/a_932_472# vdd 0.003166f
C4458 FILLER_0_17_161/a_124_375# _098_ 0.002013f
C4459 trim_mask\[4\] net47 0.264421f
C4460 _404_/a_36_472# _183_ 0.002637f
C4461 FILLER_0_7_104/a_1020_375# _153_ 0.026997f
C4462 _176_ _129_ 0.036112f
C4463 FILLER_0_21_125/a_484_472# _140_ 0.013936f
C4464 _144_ FILLER_0_21_133/a_124_375# 0.001885f
C4465 FILLER_0_18_177/a_1468_375# FILLER_0_20_177/a_1380_472# 0.0027f
C4466 result[4] net62 0.050684f
C4467 _442_/a_2665_112# vss 0.001727f
C4468 _442_/a_2560_156# vdd 0.006195f
C4469 _442_/a_36_151# _158_ 0.001257f
C4470 mask\[9\] _438_/a_36_151# 0.060632f
C4471 FILLER_0_10_37/a_36_472# net51 0.002346f
C4472 _030_ _367_/a_36_68# 0.015584f
C4473 _149_ FILLER_0_20_87/a_36_472# 0.001938f
C4474 _079_ FILLER_0_5_212/a_36_472# 0.005671f
C4475 net15 FILLER_0_6_47/a_1828_472# 0.014911f
C4476 FILLER_0_10_28/a_124_375# net17 0.00917f
C4477 FILLER_0_18_177/a_2364_375# vdd 0.020562f
C4478 _449_/a_2248_156# _067_ 0.040648f
C4479 _415_/a_36_151# FILLER_0_10_256/a_36_472# 0.004847f
C4480 cal_itt\[3\] FILLER_0_5_198/a_36_472# 0.07099f
C4481 FILLER_0_11_101/a_124_375# cal_count\[3\] 0.00419f
C4482 _450_/a_1040_527# _039_ 0.015478f
C4483 _415_/a_36_151# net64 0.001735f
C4484 _186_ _185_ 0.007962f
C4485 output32/a_224_472# net78 0.002901f
C4486 FILLER_0_17_133/a_36_472# _137_ 0.001963f
C4487 _130_ _125_ 0.002745f
C4488 _093_ _103_ 0.124026f
C4489 FILLER_0_18_2/a_3260_375# net40 0.035372f
C4490 _132_ net53 0.035348f
C4491 FILLER_0_9_223/a_572_375# _055_ 0.022619f
C4492 net16 FILLER_0_18_37/a_1020_375# 0.005406f
C4493 _091_ vss 0.56693f
C4494 FILLER_0_15_282/a_572_375# _006_ 0.001054f
C4495 _095_ FILLER_0_15_72/a_484_472# 0.002306f
C4496 net81 _019_ 0.004079f
C4497 FILLER_0_15_142/a_36_472# net73 0.001893f
C4498 fanout70/a_36_113# net73 0.21211f
C4499 _399_/a_224_472# net16 0.003817f
C4500 net69 _441_/a_36_151# 0.035817f
C4501 _076_ _059_ 1.03702f
C4502 FILLER_0_18_171/a_36_472# vdd 0.010704f
C4503 net81 cal_itt\[1\] 0.387207f
C4504 FILLER_0_15_142/a_484_472# _427_/a_36_151# 0.001723f
C4505 _430_/a_36_151# net21 0.019114f
C4506 _187_ _042_ 0.009526f
C4507 mask\[7\] FILLER_0_22_128/a_2364_375# 0.003632f
C4508 net17 FILLER_0_20_15/a_1468_375# 0.010099f
C4509 _163_ FILLER_0_5_148/a_36_472# 0.002454f
C4510 _033_ vdd 0.509957f
C4511 _129_ _124_ 0.010499f
C4512 FILLER_0_10_78/a_1020_375# _176_ 0.020379f
C4513 cal_count\[2\] FILLER_0_15_10/a_36_472# 0.015502f
C4514 _412_/a_36_151# net59 0.003938f
C4515 FILLER_0_15_116/a_124_375# FILLER_0_14_107/a_1020_375# 0.026339f
C4516 FILLER_0_4_197/a_572_375# vdd 0.002455f
C4517 net36 net71 0.148833f
C4518 _065_ net41 0.001765f
C4519 FILLER_0_24_290/a_124_375# vdd 0.026739f
C4520 _093_ FILLER_0_18_61/a_36_472# 0.004039f
C4521 net53 _427_/a_36_151# 0.13192f
C4522 net56 _427_/a_2665_112# 0.012193f
C4523 FILLER_0_14_123/a_36_472# FILLER_0_14_107/a_1380_472# 0.013276f
C4524 net31 FILLER_0_16_255/a_124_375# 0.029277f
C4525 state\[1\] FILLER_0_12_196/a_124_375# 0.063785f
C4526 _248_/a_36_68# _090_ 0.041161f
C4527 _448_/a_36_151# net22 0.027581f
C4528 _428_/a_2248_156# _043_ 0.011841f
C4529 trim_val\[3\] trim_mask\[3\] 0.48462f
C4530 fanout74/a_36_113# vdd 0.099021f
C4531 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_124_375# 0.012222f
C4532 net52 _439_/a_448_472# 0.042072f
C4533 FILLER_0_9_223/a_36_472# _068_ 0.076678f
C4534 FILLER_0_10_78/a_124_375# _176_ 0.002785f
C4535 _335_/a_257_69# mask\[1\] 0.001543f
C4536 _412_/a_1000_472# net1 0.027748f
C4537 _250_/a_36_68# vdd 0.014409f
C4538 net74 trim_mask\[4\] 0.548293f
C4539 FILLER_0_24_96/a_36_472# net35 0.002526f
C4540 _114_ _043_ 0.071339f
C4541 _176_ _394_/a_1936_472# 0.001255f
C4542 _128_ _113_ 0.002117f
C4543 en_co_clk cal_count\[3\] 0.001359f
C4544 trimb[1] net38 0.161478f
C4545 _180_ vdd 0.176915f
C4546 _428_/a_1000_472# _095_ 0.001101f
C4547 _028_ FILLER_0_6_47/a_2364_375# 0.016593f
C4548 net74 net47 0.030815f
C4549 net62 net64 0.078454f
C4550 net79 net21 0.645949f
C4551 _443_/a_2665_112# _170_ 0.019855f
C4552 net15 _440_/a_1000_472# 0.056791f
C4553 state\[2\] FILLER_0_13_142/a_484_472# 0.004186f
C4554 net53 FILLER_0_13_142/a_1380_472# 0.041222f
C4555 _053_ _414_/a_796_472# 0.008213f
C4556 _015_ FILLER_0_8_247/a_572_375# 0.00706f
C4557 _421_/a_36_151# net77 0.028951f
C4558 FILLER_0_3_78/a_124_375# vss 0.004739f
C4559 FILLER_0_3_78/a_572_375# vdd 0.014442f
C4560 _432_/a_1000_472# net80 0.033803f
C4561 FILLER_0_2_127/a_124_375# vdd 0.013496f
C4562 _394_/a_1336_472# _095_ 0.031869f
C4563 FILLER_0_24_274/a_932_472# vss 0.001001f
C4564 _132_ FILLER_0_14_107/a_124_375# 0.003315f
C4565 _448_/a_2560_156# _037_ 0.011661f
C4566 output42/a_224_472# output6/a_224_472# 0.292612f
C4567 vss trim[2] 0.026644f
C4568 _326_/a_36_160# _134_ 0.003299f
C4569 _348_/a_665_69# _146_ 0.001153f
C4570 FILLER_0_22_128/a_36_472# vdd 0.004601f
C4571 FILLER_0_22_128/a_3260_375# vss 0.006346f
C4572 _175_ _040_ 0.00133f
C4573 net33 vss 0.674927f
C4574 _372_/a_170_472# net23 0.025555f
C4575 net27 _426_/a_448_472# 0.023676f
C4576 output15/a_224_472# FILLER_0_0_96/a_36_472# 0.023414f
C4577 net56 FILLER_0_18_139/a_124_375# 0.00281f
C4578 trimb[0] vss 0.097724f
C4579 FILLER_0_12_20/a_124_375# net6 0.003726f
C4580 _079_ FILLER_0_3_172/a_2276_472# 0.00261f
C4581 _425_/a_448_472# net19 0.034226f
C4582 net60 _007_ 0.025806f
C4583 _053_ FILLER_0_6_47/a_1468_375# 0.008103f
C4584 fanout70/a_36_113# _131_ 0.003364f
C4585 net76 _083_ 0.002446f
C4586 net82 FILLER_0_3_172/a_1916_375# 0.010202f
C4587 _260_/a_36_68# net59 0.004346f
C4588 _411_/a_36_151# FILLER_0_0_232/a_124_375# 0.059049f
C4589 FILLER_0_13_228/a_36_472# _043_ 0.02119f
C4590 _235_/a_67_603# _447_/a_36_151# 0.038675f
C4591 FILLER_0_17_38/a_484_472# vss 0.001229f
C4592 trim_mask\[4\] _159_ 0.049552f
C4593 FILLER_0_3_172/a_1020_375# net65 0.006035f
C4594 net19 _082_ 0.029316f
C4595 _127_ _085_ 0.00179f
C4596 _446_/a_36_151# vdd 0.06703f
C4597 net79 _418_/a_448_472# 0.034736f
C4598 net82 net19 1.14585f
C4599 vss FILLER_0_3_212/a_36_472# 0.00838f
C4600 FILLER_0_6_177/a_36_472# _163_ 0.025039f
C4601 _159_ net47 0.01358f
C4602 _449_/a_36_151# FILLER_0_12_50/a_124_375# 0.017882f
C4603 net62 _006_ 0.136418f
C4604 _376_/a_36_160# _163_ 0.006811f
C4605 net16 _453_/a_36_151# 0.001634f
C4606 _322_/a_124_24# _126_ 0.019609f
C4607 net72 _401_/a_36_68# 0.006818f
C4608 net7 net17 0.050676f
C4609 FILLER_0_17_282/a_124_375# vss 0.024404f
C4610 FILLER_0_17_282/a_36_472# vdd 0.107351f
C4611 _081_ _059_ 0.04053f
C4612 _316_/a_848_380# _122_ 0.002234f
C4613 _316_/a_692_472# calibrate 0.006232f
C4614 _161_ _267_/a_36_472# 0.043279f
C4615 net58 net75 0.061787f
C4616 _086_ cal_count\[3\] 0.259095f
C4617 _115_ FILLER_0_9_105/a_484_472# 0.004075f
C4618 net79 FILLER_0_21_286/a_572_375# 0.001476f
C4619 net4 net59 0.102012f
C4620 FILLER_0_9_142/a_124_375# _118_ 0.06224f
C4621 _429_/a_2665_112# net64 0.013014f
C4622 _306_/a_36_68# vss 0.008326f
C4623 trim_mask\[4\] _154_ 0.014658f
C4624 _053_ net50 0.711279f
C4625 _449_/a_36_151# _394_/a_728_93# 0.002727f
C4626 net33 _107_ 0.001322f
C4627 net2 cal_itt\[1\] 0.284695f
C4628 _144_ FILLER_0_19_155/a_572_375# 0.003611f
C4629 net73 FILLER_0_17_142/a_36_472# 0.002925f
C4630 output43/a_224_472# trimb[0] 0.043402f
C4631 _448_/a_36_151# vdd 0.133302f
C4632 net47 _154_ 0.055128f
C4633 _115_ vss 0.372063f
C4634 _413_/a_36_151# FILLER_0_2_177/a_572_375# 0.073306f
C4635 _028_ FILLER_0_5_72/a_1468_375# 0.00123f
C4636 _310_/a_49_472# vdd 0.043164f
C4637 net81 fanout79/a_36_160# 0.057526f
C4638 FILLER_0_23_60/a_36_472# vdd 0.090554f
C4639 FILLER_0_23_60/a_124_375# vss 0.004081f
C4640 result[4] _417_/a_2560_156# 0.001076f
C4641 mask\[9\] FILLER_0_20_98/a_36_472# 0.005917f
C4642 cal_count\[2\] _182_ 0.044348f
C4643 net55 FILLER_0_19_28/a_36_472# 0.001572f
C4644 FILLER_0_3_142/a_124_375# trim_mask\[4\] 0.002514f
C4645 net75 calibrate 0.101912f
C4646 FILLER_0_18_100/a_36_472# vdd 0.012574f
C4647 FILLER_0_18_100/a_124_375# vss 0.025563f
C4648 net78 _094_ 0.050187f
C4649 _442_/a_36_151# net23 0.00157f
C4650 _104_ net30 0.001375f
C4651 _021_ _432_/a_36_151# 0.033849f
C4652 _379_/a_36_472# _160_ 0.023459f
C4653 ctlp[3] ctlp[2] 0.006764f
C4654 net55 _423_/a_2248_156# 0.001188f
C4655 _176_ FILLER_0_11_101/a_572_375# 0.00389f
C4656 net54 FILLER_0_22_107/a_484_472# 0.005897f
C4657 FILLER_0_14_99/a_124_375# net14 0.04852f
C4658 net75 FILLER_0_10_256/a_124_375# 0.027258f
C4659 _004_ net58 0.00116f
C4660 _010_ vdd 0.121474f
C4661 FILLER_0_14_263/a_124_375# vdd 0.026205f
C4662 FILLER_0_21_142/a_572_375# net23 0.007884f
C4663 _053_ FILLER_0_7_72/a_3172_472# 0.032946f
C4664 _386_/a_124_24# _169_ 0.02709f
C4665 FILLER_0_17_72/a_572_375# vss 0.008057f
C4666 FILLER_0_17_72/a_1020_375# vdd 0.002541f
C4667 _274_/a_1612_497# net4 0.00807f
C4668 FILLER_0_17_161/a_36_472# _137_ 0.013985f
C4669 net4 _122_ 0.03487f
C4670 net73 FILLER_0_18_107/a_1828_472# 0.01544f
C4671 FILLER_0_4_197/a_36_472# net22 0.003404f
C4672 net20 _010_ 0.016197f
C4673 FILLER_0_4_107/a_1020_375# vdd 0.025121f
C4674 _273_/a_36_68# FILLER_0_10_214/a_124_375# 0.003707f
C4675 net74 _159_ 0.129233f
C4676 FILLER_0_9_270/a_572_375# vdd 0.02345f
C4677 FILLER_0_19_28/a_36_472# net17 0.009277f
C4678 _415_/a_2248_156# output27/a_224_472# 0.001506f
C4679 output21/a_224_472# output19/a_224_472# 0.007877f
C4680 net38 FILLER_0_20_2/a_36_472# 0.002204f
C4681 _230_/a_244_68# _060_ 0.002039f
C4682 net17 _450_/a_36_151# 0.006157f
C4683 FILLER_0_21_125/a_36_472# _098_ 0.002923f
C4684 _093_ mask\[2\] 0.009354f
C4685 result[9] _418_/a_2248_156# 0.043716f
C4686 FILLER_0_16_241/a_124_375# _099_ 0.040547f
C4687 net52 FILLER_0_2_111/a_124_375# 0.00483f
C4688 ctlp[2] _422_/a_448_472# 0.011383f
C4689 _063_ _166_ 0.025402f
C4690 _089_ net21 0.006605f
C4691 net4 net64 0.060449f
C4692 mask\[4\] FILLER_0_19_195/a_124_375# 0.006236f
C4693 _004_ FILLER_0_10_256/a_124_375# 0.006989f
C4694 FILLER_0_21_142/a_484_472# vdd 0.004917f
C4695 net52 _440_/a_36_151# 0.01571f
C4696 net57 FILLER_0_16_154/a_1380_472# 0.041458f
C4697 net60 _421_/a_796_472# 0.002046f
C4698 net74 _154_ 0.002976f
C4699 valid cal_itt\[1\] 0.011576f
C4700 _449_/a_2665_112# net74 0.001185f
C4701 _401_/a_244_472# _180_ 0.001689f
C4702 ctlp[5] _435_/a_36_151# 0.003815f
C4703 net41 _445_/a_2560_156# 0.002221f
C4704 net53 FILLER_0_14_107/a_1380_472# 0.059367f
C4705 trim[0] _034_ 0.044322f
C4706 _091_ _275_/a_224_472# 0.003461f
C4707 net79 mask\[1\] 0.029512f
C4708 ctlp[6] output24/a_224_472# 0.004288f
C4709 net81 _429_/a_1000_472# 0.011018f
C4710 _415_/a_1000_472# _004_ 0.005004f
C4711 _141_ FILLER_0_19_155/a_124_375# 0.029562f
C4712 FILLER_0_23_282/a_36_472# vdd 0.106034f
C4713 FILLER_0_23_282/a_572_375# vss 0.058599f
C4714 _438_/a_2560_156# vdd 0.001166f
C4715 _438_/a_2665_112# vss 0.001389f
C4716 FILLER_0_13_142/a_36_472# vdd 0.104785f
C4717 ctlp[6] vss 0.115894f
C4718 FILLER_0_13_142/a_1468_375# vss 0.00614f
C4719 net66 _440_/a_796_472# 0.002718f
C4720 net49 _440_/a_36_151# 0.021133f
C4721 _127_ _062_ 0.020537f
C4722 _143_ _343_/a_49_472# 0.00918f
C4723 _131_ FILLER_0_17_64/a_36_472# 0.002638f
C4724 net52 FILLER_0_5_72/a_932_472# 0.008749f
C4725 _257_/a_36_472# _068_ 0.002986f
C4726 FILLER_0_19_142/a_124_375# vdd 0.022448f
C4727 net72 _095_ 0.136566f
C4728 net1 fanout59/a_36_160# 0.002325f
C4729 result[7] _298_/a_224_472# 0.007724f
C4730 FILLER_0_17_56/a_572_375# FILLER_0_18_61/a_36_472# 0.001597f
C4731 cal_count\[3\] _090_ 0.243462f
C4732 _447_/a_36_151# vdd 0.067176f
C4733 _048_ FILLER_0_18_209/a_124_375# 0.001615f
C4734 output36/a_224_472# net29 0.077505f
C4735 _087_ FILLER_0_5_172/a_36_472# 0.00443f
C4736 net29 net30 0.053996f
C4737 result[2] output30/a_224_472# 0.045862f
C4738 ctlp[2] _108_ 0.034027f
C4739 FILLER_0_19_55/a_124_375# vss 0.001882f
C4740 FILLER_0_19_55/a_36_472# vdd 0.085984f
C4741 _152_ FILLER_0_5_136/a_36_472# 0.049485f
C4742 FILLER_0_24_96/a_36_472# vdd 0.094828f
C4743 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_572_375# 0.026339f
C4744 net81 FILLER_0_10_247/a_124_375# 0.044906f
C4745 _137_ FILLER_0_16_154/a_124_375# 0.007998f
C4746 _292_/a_36_160# _201_/a_67_603# 0.003917f
C4747 _258_/a_36_160# _079_ 0.026618f
C4748 _031_ _157_ 0.104339f
C4749 ctlp[2] net19 0.017506f
C4750 net54 _433_/a_448_472# 0.008777f
C4751 _164_ FILLER_0_6_47/a_932_472# 0.004272f
C4752 FILLER_0_11_282/a_36_472# vss 0.007114f
C4753 _106_ _092_ 0.140596f
C4754 FILLER_0_20_107/a_36_472# _098_ 0.011046f
C4755 mask\[4\] FILLER_0_18_177/a_1828_472# 0.014226f
C4756 _256_/a_716_497# net4 0.001936f
C4757 FILLER_0_9_223/a_572_375# _426_/a_2665_112# 0.005202f
C4758 FILLER_0_8_107/a_124_375# _058_ 0.01823f
C4759 _093_ FILLER_0_16_115/a_124_375# 0.003988f
C4760 _431_/a_2248_156# _137_ 0.01617f
C4761 _136_ _097_ 0.002577f
C4762 FILLER_0_17_38/a_572_375# _179_ 0.002825f
C4763 _053_ cal_itt\[3\] 0.471909f
C4764 FILLER_0_14_81/a_36_472# _394_/a_728_93# 0.005826f
C4765 _018_ net22 0.141743f
C4766 _091_ _095_ 0.005006f
C4767 net81 FILLER_0_15_228/a_124_375# 0.006974f
C4768 _133_ _134_ 0.015205f
C4769 _186_ net17 0.001172f
C4770 vdd FILLER_0_10_94/a_124_375# 0.020076f
C4771 result[5] _418_/a_448_472# 0.007308f
C4772 _417_/a_2560_156# _006_ 0.007804f
C4773 net35 vss 0.434438f
C4774 _299_/a_36_472# vdd 0.098451f
C4775 _140_ FILLER_0_21_150/a_124_375# 0.019084f
C4776 _320_/a_224_472# _113_ 0.00871f
C4777 net56 FILLER_0_17_142/a_36_472# 0.003603f
C4778 _137_ _043_ 0.007284f
C4779 FILLER_0_4_197/a_36_472# vdd 0.042721f
C4780 output32/a_224_472# _418_/a_2248_156# 0.024448f
C4781 _415_/a_2248_156# _416_/a_36_151# 0.001495f
C4782 output21/a_224_472# mask\[6\] 0.013037f
C4783 result[6] FILLER_0_21_286/a_36_472# 0.015369f
C4784 _449_/a_448_472# net72 0.01383f
C4785 _091_ FILLER_0_12_220/a_124_375# 0.006907f
C4786 _025_ _436_/a_448_472# 0.044246f
C4787 FILLER_0_17_226/a_124_375# fanout63/a_36_160# 0.008215f
C4788 _079_ _253_/a_36_68# 0.002433f
C4789 _316_/a_1084_68# vdd 0.001166f
C4790 net79 _416_/a_2560_156# 0.013576f
C4791 net55 FILLER_0_18_76/a_484_472# 0.003745f
C4792 _444_/a_36_151# vdd 0.071209f
C4793 _093_ FILLER_0_19_111/a_572_375# 0.002743f
C4794 cal_count\[3\] _408_/a_56_524# 0.001685f
C4795 _238_/a_67_603# net52 0.006325f
C4796 _000_ _083_ 0.017601f
C4797 _136_ mask\[2\] 1.822289f
C4798 _193_/a_36_160# _044_ 0.025719f
C4799 output10/a_224_472# FILLER_0_0_266/a_124_375# 0.00515f
C4800 FILLER_0_4_197/a_1020_375# _088_ 0.013641f
C4801 _390_/a_36_68# net14 0.010844f
C4802 _198_/a_67_603# _099_ 0.0109f
C4803 _306_/a_36_68# _071_ 0.054312f
C4804 _453_/a_1000_472# _042_ 0.004985f
C4805 result[8] FILLER_0_24_274/a_36_472# 0.005458f
C4806 output31/a_224_472# FILLER_0_17_282/a_124_375# 0.002977f
C4807 _058_ FILLER_0_10_94/a_484_472# 0.002096f
C4808 _311_/a_1212_473# _117_ 0.001673f
C4809 FILLER_0_20_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001543f
C4810 _412_/a_1000_472# net76 0.024114f
C4811 _448_/a_448_472# net76 0.003937f
C4812 _119_ _115_ 0.06747f
C4813 result[7] _419_/a_2248_156# 0.001916f
C4814 FILLER_0_2_93/a_124_375# vdd 0.008901f
C4815 vss _167_ 0.043544f
C4816 _080_ vdd 0.123811f
C4817 _118_ _331_/a_448_472# 0.001166f
C4818 FILLER_0_19_171/a_36_472# vdd 0.004762f
C4819 FILLER_0_19_171/a_1468_375# vss 0.054352f
C4820 FILLER_0_22_86/a_1380_472# net71 0.011277f
C4821 mask\[8\] _437_/a_36_151# 0.005179f
C4822 FILLER_0_18_139/a_1468_375# _137_ 0.004111f
C4823 net16 _013_ 0.060401f
C4824 mask\[4\] FILLER_0_22_128/a_3172_472# 0.001484f
C4825 FILLER_0_5_109/a_484_472# net47 0.002299f
C4826 _036_ FILLER_0_3_78/a_124_375# 0.00215f
C4827 _088_ FILLER_0_4_213/a_484_472# 0.018066f
C4828 cal_count\[3\] _314_/a_224_472# 0.002143f
C4829 net60 net30 0.001168f
C4830 _452_/a_3129_107# vdd 0.016611f
C4831 input5/a_36_113# clk 0.01086f
C4832 net72 FILLER_0_21_28/a_1380_472# 0.048287f
C4833 _058_ _122_ 0.040376f
C4834 result[7] result[8] 0.201281f
C4835 net20 _080_ 0.093195f
C4836 _235_/a_67_603# vss 0.002019f
C4837 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2812_375# 0.001597f
C4838 FILLER_0_7_195/a_36_472# vdd 0.04565f
C4839 FILLER_0_7_195/a_124_375# vss 0.006314f
C4840 net47 FILLER_0_5_148/a_124_375# 0.008947f
C4841 net58 net19 0.044785f
C4842 net1 net5 0.266194f
C4843 mask\[0\] net79 0.243338f
C4844 _253_/a_36_68# cal_itt\[1\] 0.039692f
C4845 FILLER_0_6_177/a_484_472# FILLER_0_5_181/a_36_472# 0.05841f
C4846 _359_/a_36_488# _129_ 0.002527f
C4847 FILLER_0_23_44/a_572_375# vdd -0.011314f
C4848 FILLER_0_10_214/a_36_472# _246_/a_36_68# 0.001844f
C4849 _058_ _227_/a_36_160# 0.008511f
C4850 _004_ mask\[1\] 0.052788f
C4851 trim_mask\[2\] _168_ 0.00704f
C4852 FILLER_0_7_59/a_124_375# FILLER_0_6_47/a_1468_375# 0.05841f
C4853 _077_ _055_ 0.083808f
C4854 net22 vss 1.28233f
C4855 FILLER_0_16_89/a_36_472# FILLER_0_17_72/a_1916_375# 0.001723f
C4856 FILLER_0_16_89/a_1020_375# FILLER_0_17_72/a_2812_375# 0.026339f
C4857 _018_ vdd 0.048119f
C4858 _440_/a_1000_472# net47 0.011283f
C4859 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_572_375# 0.086635f
C4860 net19 calibrate 0.043159f
C4861 FILLER_0_14_107/a_1468_375# vss 0.055167f
C4862 FILLER_0_14_107/a_36_472# vdd 0.114495f
C4863 FILLER_0_9_72/a_1380_472# vss 0.007254f
C4864 _448_/a_36_151# FILLER_0_2_177/a_572_375# 0.001597f
C4865 FILLER_0_18_177/a_3260_375# FILLER_0_18_209/a_36_472# 0.086742f
C4866 _136_ FILLER_0_16_115/a_124_375# 0.006372f
C4867 _114_ FILLER_0_12_136/a_484_472# 0.003953f
C4868 _343_/a_257_69# _137_ 0.003494f
C4869 FILLER_0_22_177/a_572_375# net33 0.013337f
C4870 _433_/a_36_151# _022_ 0.017789f
C4871 fanout66/a_36_113# net66 0.032757f
C4872 cal_itt\[3\] _375_/a_36_68# 0.005168f
C4873 FILLER_0_10_256/a_124_375# net19 0.002884f
C4874 _395_/a_36_488# _071_ 0.00276f
C4875 FILLER_0_17_72/a_1468_375# _150_ 0.001076f
C4876 _010_ _419_/a_796_472# 0.001613f
C4877 _445_/a_36_151# net17 0.009838f
C4878 _437_/a_2665_112# FILLER_0_22_107/a_572_375# 0.001597f
C4879 FILLER_0_21_28/a_36_472# net17 0.00347f
C4880 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_124_375# 0.003732f
C4881 _306_/a_36_68# _095_ 0.001366f
C4882 FILLER_0_16_107/a_36_472# net14 0.004691f
C4883 net63 net21 0.278824f
C4884 _069_ _310_/a_49_472# 0.023925f
C4885 ctlp[3] mask\[7\] 0.103955f
C4886 net50 fanout49/a_36_160# 0.059373f
C4887 _415_/a_1000_472# net19 0.001125f
C4888 net50 FILLER_0_7_59/a_124_375# 0.002292f
C4889 _077_ _255_/a_224_552# 0.025141f
C4890 _071_ FILLER_0_13_142/a_1468_375# 0.007453f
C4891 FILLER_0_18_2/a_2364_375# vdd 0.002983f
C4892 net63 FILLER_0_19_171/a_932_472# 0.00128f
C4893 _096_ net57 0.05086f
C4894 _402_/a_728_93# cal_count\[1\] 0.057043f
C4895 net54 FILLER_0_22_86/a_932_472# 0.047897f
C4896 net79 _099_ 0.010543f
C4897 _136_ FILLER_0_16_154/a_484_472# 0.007583f
C4898 net3 FILLER_0_15_2/a_484_472# 0.002224f
C4899 net53 mask\[2\] 0.005907f
C4900 _428_/a_1308_423# _131_ 0.037599f
C4901 net48 _316_/a_124_24# 0.068708f
C4902 net52 _170_ 0.378738f
C4903 net60 _417_/a_36_151# 0.007446f
C4904 FILLER_0_7_72/a_1468_375# vss 0.003253f
C4905 trim[2] output41/a_224_472# 0.005452f
C4906 output40/a_224_472# trim[3] 0.122003f
C4907 FILLER_0_9_223/a_572_375# _223_/a_36_160# 0.001177f
C4908 _431_/a_36_151# FILLER_0_16_115/a_124_375# 0.035117f
C4909 _328_/a_36_113# _126_ 0.023932f
C4910 mask\[8\] _051_ 0.003475f
C4911 _059_ _163_ 0.038651f
C4912 mask\[5\] FILLER_0_18_177/a_36_472# 0.001063f
C4913 result[0] net5 0.001104f
C4914 FILLER_0_16_89/a_484_472# _040_ 0.009871f
C4915 _087_ _088_ 0.001219f
C4916 vss _433_/a_2665_112# 0.035903f
C4917 mask\[0\] _429_/a_2560_156# 0.010913f
C4918 net16 FILLER_0_6_37/a_124_375# 0.010358f
C4919 cal_count\[3\] FILLER_0_11_78/a_124_375# 0.019818f
C4920 _402_/a_56_567# net40 0.033835f
C4921 FILLER_0_3_172/a_3260_375# net22 0.015274f
C4922 _413_/a_2248_156# net59 0.05485f
C4923 net73 FILLER_0_17_104/a_1468_375# 0.002342f
C4924 _094_ _418_/a_2248_156# 0.028557f
C4925 FILLER_0_12_136/a_124_375# _127_ 0.004013f
C4926 _422_/a_448_472# mask\[7\] 0.048658f
C4927 FILLER_0_16_57/a_1380_472# _131_ 0.008223f
C4928 fanout66/a_36_113# FILLER_0_3_54/a_124_375# 0.002853f
C4929 _086_ _267_/a_224_472# 0.004041f
C4930 net44 _221_/a_36_160# 0.013363f
C4931 _430_/a_796_472# mask\[2\] 0.006305f
C4932 _054_ vdd 0.360345f
C4933 FILLER_0_9_60/a_36_472# net51 0.059421f
C4934 FILLER_0_6_177/a_124_375# net47 0.002925f
C4935 net75 output48/a_224_472# 0.070114f
C4936 _116_ _085_ 0.049304f
C4937 fanout77/a_36_113# _103_ 0.006045f
C4938 _321_/a_2590_472# _176_ 0.001932f
C4939 _069_ _395_/a_1044_488# 0.002244f
C4940 FILLER_0_17_200/a_572_375# _430_/a_36_151# 0.059049f
C4941 _445_/a_1204_472# net40 0.003916f
C4942 _273_/a_36_68# _076_ 0.001503f
C4943 _132_ _149_ 0.087289f
C4944 ctln[5] _037_ 0.19244f
C4945 net75 FILLER_0_8_247/a_124_375# 0.002085f
C4946 _126_ _120_ 0.055349f
C4947 _126_ _038_ 0.031198f
C4948 FILLER_0_15_235/a_572_375# vss 0.002683f
C4949 FILLER_0_15_235/a_36_472# vdd 0.019127f
C4950 vdd _278_/a_36_160# 0.016488f
C4951 FILLER_0_9_105/a_36_472# vss 0.002744f
C4952 FILLER_0_9_105/a_484_472# vdd 0.03152f
C4953 _053_ FILLER_0_5_54/a_484_472# 0.001135f
C4954 FILLER_0_8_138/a_36_472# vss 0.008189f
C4955 FILLER_0_13_142/a_484_472# _043_ 0.011974f
C4956 FILLER_0_20_177/a_484_472# vss 0.001256f
C4957 FILLER_0_20_177/a_932_472# vdd 0.035019f
C4958 FILLER_0_18_2/a_3260_375# FILLER_0_20_31/a_36_472# 0.001338f
C4959 net81 _425_/a_2665_112# 0.010188f
C4960 FILLER_0_4_185/a_36_472# FILLER_0_4_177/a_484_472# 0.013276f
C4961 output24/a_224_472# vdd 0.08781f
C4962 _008_ FILLER_0_17_226/a_36_472# 0.001842f
C4963 _326_/a_36_160# _322_/a_124_24# 0.004397f
C4964 _274_/a_36_68# _070_ 0.032424f
C4965 ctlp[3] _422_/a_2248_156# 0.001888f
C4966 vdd vss 15.42941f
C4967 FILLER_0_2_101/a_124_375# _160_ 0.001047f
C4968 _192_/a_67_603# vss 0.007021f
C4969 net16 _447_/a_1204_472# 0.00194f
C4970 output16/a_224_472# _447_/a_2665_112# 0.005471f
C4971 _178_ vdd 0.440802f
C4972 FILLER_0_13_65/a_36_472# net72 0.00272f
C4973 net36 FILLER_0_15_212/a_1468_375# 0.005276f
C4974 _408_/a_1336_472# _186_ 0.010089f
C4975 net20 FILLER_0_15_235/a_36_472# 0.002227f
C4976 net41 FILLER_0_18_37/a_36_472# 0.007459f
C4977 input2/a_36_113# input5/a_36_113# 0.01088f
C4978 _013_ _041_ 0.00271f
C4979 FILLER_0_17_56/a_124_375# _183_ 0.019253f
C4980 FILLER_0_2_165/a_36_472# net22 0.028367f
C4981 FILLER_0_20_98/a_124_375# net14 0.05242f
C4982 FILLER_0_20_15/a_932_472# vdd 0.002617f
C4983 cal_count\[3\] _117_ 0.00114f
C4984 mask\[7\] _108_ 0.785154f
C4985 _104_ _046_ 0.035267f
C4986 fanout70/a_36_113# FILLER_0_15_116/a_484_472# 0.002001f
C4987 _079_ cal_itt\[1\] 0.012324f
C4988 FILLER_0_24_130/a_36_472# net54 0.06125f
C4989 FILLER_0_18_107/a_1020_375# vdd -0.008765f
C4990 _411_/a_1204_472# net75 0.008304f
C4991 FILLER_0_5_109/a_484_472# _154_ 0.039428f
C4992 _076_ FILLER_0_8_239/a_124_375# 0.007237f
C4993 mask\[3\] net36 0.002974f
C4994 _422_/a_1000_472# vdd 0.005284f
C4995 net20 vss 1.402494f
C4996 _063_ trim_val\[1\] 0.038045f
C4997 net63 mask\[7\] 0.069252f
C4998 mask\[7\] net19 0.003605f
C4999 cal_count\[2\] _452_/a_2225_156# 0.003086f
C5000 _062_ _060_ 0.032472f
C5001 _106_ FILLER_0_17_218/a_36_472# 0.002777f
C5002 net79 FILLER_0_12_220/a_1020_375# 0.010818f
C5003 FILLER_0_18_139/a_124_375# _145_ 0.00346f
C5004 _441_/a_2248_156# vdd -0.003818f
C5005 _441_/a_1204_472# vss 0.011996f
C5006 FILLER_0_3_221/a_124_375# FILLER_0_3_212/a_124_375# 0.002036f
C5007 _232_/a_255_603# _164_ 0.001274f
C5008 _031_ _158_ 0.015116f
C5009 FILLER_0_7_72/a_36_472# vdd 0.106377f
C5010 trim_val\[4\] _386_/a_124_24# 0.001172f
C5011 FILLER_0_9_223/a_124_375# _076_ 0.004399f
C5012 _430_/a_2248_156# vss 0.030251f
C5013 _447_/a_448_472# net68 0.012962f
C5014 _165_ FILLER_0_6_47/a_36_472# 0.077573f
C5015 FILLER_0_8_239/a_36_472# _317_/a_36_113# 0.00191f
C5016 FILLER_0_19_47/a_124_375# net26 0.008432f
C5017 _039_ cal_count\[0\] 0.219667f
C5018 _132_ _134_ 0.029512f
C5019 output43/a_224_472# vdd -0.032713f
C5020 _131_ FILLER_0_17_104/a_1468_375# 0.006022f
C5021 ctlp[1] _421_/a_2560_156# 0.001062f
C5022 fanout71/a_36_113# net71 0.087994f
C5023 vdd _107_ 0.038236f
C5024 FILLER_0_21_28/a_1916_375# _423_/a_36_151# 0.001597f
C5025 net69 _030_ 0.49547f
C5026 _077_ _414_/a_2665_112# 0.001675f
C5027 net15 _423_/a_1308_423# 0.001999f
C5028 _226_/a_1044_68# net21 0.001903f
C5029 FILLER_0_16_73/a_36_472# _394_/a_1336_472# 0.00108f
C5030 _442_/a_1308_423# FILLER_0_2_111/a_1468_375# 0.001048f
C5031 _449_/a_1308_423# _038_ 0.021006f
C5032 FILLER_0_24_96/a_124_375# net35 0.001886f
C5033 FILLER_0_3_172/a_3260_375# vdd -0.013516f
C5034 output8/a_224_472# net82 0.002936f
C5035 _359_/a_1492_488# _133_ 0.003815f
C5036 FILLER_0_5_54/a_1468_375# _440_/a_36_151# 0.059049f
C5037 net50 net17 0.010654f
C5038 FILLER_0_15_290/a_36_472# net18 0.002452f
C5039 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_36_472# 0.086635f
C5040 FILLER_0_11_101/a_36_472# net14 0.04522f
C5041 result[6] _420_/a_2248_156# 0.003418f
C5042 FILLER_0_15_290/a_124_375# result[3] 0.020277f
C5043 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_1020_375# 0.026339f
C5044 net50 trim_val\[1\] 0.002079f
C5045 FILLER_0_7_104/a_572_375# _058_ 0.006125f
C5046 _127_ _428_/a_36_151# 0.030717f
C5047 _052_ FILLER_0_18_37/a_572_375# 0.00706f
C5048 _251_/a_1130_472# vss 0.001211f
C5049 _267_/a_36_472# _113_ 0.014178f
C5050 FILLER_0_10_28/a_124_375# output6/a_224_472# 0.002633f
C5051 net9 vss 0.086497f
C5052 _077_ _439_/a_36_151# 0.035432f
C5053 _147_ net33 0.001686f
C5054 net63 mask\[1\] 0.120872f
C5055 _106_ _199_/a_36_160# 0.003376f
C5056 fanout76/a_36_160# vdd 0.108854f
C5057 net81 FILLER_0_14_235/a_36_472# 0.002571f
C5058 net15 FILLER_0_17_72/a_932_472# 0.001122f
C5059 output17/a_224_472# vss 0.009426f
C5060 _144_ _433_/a_36_151# 0.086558f
C5061 FILLER_0_18_76/a_124_375# net71 0.008427f
C5062 net70 net74 0.017928f
C5063 vdd _416_/a_2248_156# 0.004325f
C5064 output46/a_224_472# net44 0.003804f
C5065 _044_ _416_/a_36_151# 0.032206f
C5066 net46 vdd 0.255965f
C5067 _422_/a_2248_156# _108_ 0.019477f
C5068 _135_ vss 0.097337f
C5069 _410_/a_36_68# _187_ 0.038745f
C5070 _126_ state\[2\] 0.030985f
C5071 FILLER_0_5_88/a_124_375# vdd 0.020896f
C5072 _115_ FILLER_0_10_78/a_36_472# 0.002611f
C5073 FILLER_0_8_107/a_124_375# _134_ 0.007753f
C5074 _422_/a_2248_156# net19 0.003451f
C5075 ctlp[5] net23 0.025206f
C5076 FILLER_0_10_214/a_124_375# _247_/a_36_160# 0.005732f
C5077 _432_/a_448_472# net80 0.045963f
C5078 FILLER_0_11_142/a_36_472# cal_count\[3\] 0.008454f
C5079 FILLER_0_22_177/a_1020_375# mask\[6\] 0.002657f
C5080 _098_ _434_/a_2560_156# 0.003888f
C5081 net35 FILLER_0_22_177/a_572_375# 0.007797f
C5082 _195_/a_67_603# vdd 0.022493f
C5083 _010_ net77 0.009534f
C5084 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3260_375# 0.086635f
C5085 _176_ FILLER_0_11_78/a_572_375# 0.013887f
C5086 _431_/a_2560_156# _136_ 0.013111f
C5087 _365_/a_244_472# net14 0.001257f
C5088 _056_ _246_/a_36_68# 0.017953f
C5089 _289_/a_36_472# _099_ 0.035055f
C5090 FILLER_0_2_165/a_36_472# vdd -0.003333f
C5091 FILLER_0_2_165/a_124_375# vss 0.008386f
C5092 net16 _064_ 0.121797f
C5093 FILLER_0_4_49/a_572_375# net49 0.004345f
C5094 fanout54/a_36_160# FILLER_0_18_139/a_1020_375# 0.031033f
C5095 ctln[6] _170_ 0.005146f
C5096 _140_ FILLER_0_22_128/a_36_472# 0.050084f
C5097 _118_ _062_ 0.029651f
C5098 result[1] FILLER_0_11_282/a_124_375# 0.018322f
C5099 fanout67/a_36_160# vss 0.005344f
C5100 result[6] _419_/a_2665_112# 0.001225f
C5101 _256_/a_1164_497# _076_ 0.001871f
C5102 _148_ FILLER_0_22_107/a_572_375# 0.00652f
C5103 _036_ _167_ 0.003223f
C5104 trim_mask\[1\] FILLER_0_6_90/a_36_472# 0.001162f
C5105 _072_ net23 0.006278f
C5106 FILLER_0_2_177/a_36_472# net22 0.002517f
C5107 FILLER_0_5_117/a_124_375# _360_/a_36_160# 0.004736f
C5108 net15 _447_/a_2560_156# 0.001586f
C5109 _323_/a_36_113# FILLER_0_10_247/a_36_472# 0.00136f
C5110 FILLER_0_14_107/a_484_472# _043_ 0.001641f
C5111 _105_ _108_ 0.548284f
C5112 _069_ _018_ 0.002777f
C5113 _077_ _426_/a_2665_112# 0.001392f
C5114 net34 FILLER_0_22_128/a_1380_472# 0.001011f
C5115 net44 cal_count\[2\] 0.191151f
C5116 result[2] FILLER_0_14_263/a_36_472# 0.001134f
C5117 _184_ vdd 0.202732f
C5118 _235_/a_67_603# _036_ 0.043345f
C5119 result[7] _421_/a_1000_472# 0.015328f
C5120 _401_/a_36_68# vdd 0.003745f
C5121 net69 trim_mask\[3\] 0.017779f
C5122 _279_/a_652_68# vdd 0.001562f
C5123 _105_ net19 0.049611f
C5124 fanout61/a_36_113# net18 0.001668f
C5125 _183_ FILLER_0_18_53/a_124_375# 0.001032f
C5126 _374_/a_36_68# FILLER_0_8_156/a_484_472# 0.002559f
C5127 _068_ _246_/a_36_68# 0.059106f
C5128 _013_ _424_/a_1308_423# 0.007751f
C5129 _095_ FILLER_0_14_107/a_1468_375# 0.010523f
C5130 net16 _042_ 0.012486f
C5131 _420_/a_1308_423# vss 0.001461f
C5132 FILLER_0_7_72/a_1828_472# _163_ 0.002095f
C5133 _359_/a_36_488# _152_ 0.032195f
C5134 net44 input3/a_36_113# 0.016865f
C5135 _057_ _311_/a_1660_473# 0.004637f
C5136 FILLER_0_19_47/a_484_472# _052_ 0.01589f
C5137 _119_ FILLER_0_8_138/a_36_472# 0.003894f
C5138 FILLER_0_5_128/a_36_472# _070_ 0.036f
C5139 FILLER_0_4_49/a_484_472# FILLER_0_3_54/a_36_472# 0.026657f
C5140 FILLER_0_12_220/a_36_472# _248_/a_36_68# 0.006596f
C5141 output47/a_224_472# FILLER_0_15_2/a_36_472# 0.035046f
C5142 FILLER_0_9_28/a_1020_375# vdd 0.033815f
C5143 _444_/a_448_472# net67 0.046278f
C5144 _177_ _451_/a_2225_156# 0.031347f
C5145 net72 _394_/a_244_524# 0.001083f
C5146 net52 _443_/a_448_472# 0.050192f
C5147 net47 _365_/a_36_68# 0.020511f
C5148 valid _425_/a_2665_112# 0.001839f
C5149 trim_mask\[0\] net14 0.499565f
C5150 _119_ vdd 0.38257f
C5151 net44 _450_/a_448_472# 0.050752f
C5152 mask\[5\] _143_ 0.032539f
C5153 _446_/a_2665_112# net66 0.00195f
C5154 vdd _450_/a_1040_527# 0.005529f
C5155 _071_ vdd 0.074299f
C5156 mask\[8\] _436_/a_36_151# 0.032521f
C5157 FILLER_0_16_241/a_36_472# net30 0.001025f
C5158 _322_/a_848_380# _070_ 0.006182f
C5159 _423_/a_2560_156# vss 0.002241f
C5160 FILLER_0_4_152/a_36_472# vss 0.009467f
C5161 net4 FILLER_0_4_213/a_572_375# 0.001015f
C5162 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001597f
C5163 output48/a_224_472# net19 0.054227f
C5164 net69 net13 0.005834f
C5165 output31/a_224_472# vdd 0.083516f
C5166 FILLER_0_16_89/a_1380_472# vdd 0.010554f
C5167 FILLER_0_9_28/a_1916_375# _453_/a_36_151# 0.001543f
C5168 ctln[7] trim_mask\[3\] 0.059414f
C5169 cal_count\[3\] _172_ 0.03048f
C5170 _316_/a_124_24# net37 0.011141f
C5171 _076_ FILLER_0_8_156/a_36_472# 0.006989f
C5172 _068_ FILLER_0_8_156/a_572_375# 0.00185f
C5173 FILLER_0_20_193/a_36_472# _098_ 0.006652f
C5174 FILLER_0_16_73/a_572_375# net15 0.002076f
C5175 FILLER_0_20_177/a_572_375# _434_/a_36_151# 0.059049f
C5176 FILLER_0_7_72/a_1380_472# vss 0.001117f
C5177 _273_/a_36_68# _090_ 0.034955f
C5178 FILLER_0_16_154/a_1020_375# vdd 0.004279f
C5179 FILLER_0_16_154/a_572_375# vss 0.003976f
C5180 cal_itt\[2\] _080_ 0.062471f
C5181 _323_/a_36_113# _128_ 0.014377f
C5182 _431_/a_1456_156# net73 0.001304f
C5183 _027_ vdd 0.146607f
C5184 FILLER_0_4_49/a_484_472# _164_ 0.003258f
C5185 output20/a_224_472# vss -0.004787f
C5186 output31/a_224_472# net20 0.004424f
C5187 _431_/a_2560_156# net53 0.002265f
C5188 _421_/a_448_472# _010_ 0.039422f
C5189 _181_ _402_/a_1948_68# 0.001223f
C5190 _274_/a_2124_68# net4 0.00137f
C5191 net22 _435_/a_2560_156# 0.002281f
C5192 FILLER_0_5_198/a_36_472# vdd 0.088893f
C5193 FILLER_0_5_198/a_572_375# vss 0.055087f
C5194 FILLER_0_22_86/a_36_472# net14 0.003007f
C5195 _065_ _441_/a_36_151# 0.00701f
C5196 _419_/a_1000_472# vdd 0.004107f
C5197 ctlp[3] result[8] 0.278543f
C5198 _132_ FILLER_0_18_107/a_2276_472# 0.006713f
C5199 _035_ _034_ 1.26804f
C5200 mask\[5\] _146_ 0.051687f
C5201 ctln[5] _448_/a_2248_156# 0.004396f
C5202 net17 _039_ 0.079171f
C5203 FILLER_0_2_177/a_36_472# vdd 0.110255f
C5204 FILLER_0_2_177/a_572_375# vss 0.008507f
C5205 ctln[1] net75 0.159105f
C5206 net27 net79 0.059863f
C5207 net19 _420_/a_1204_472# 0.001828f
C5208 _076_ _269_/a_36_472# 0.001618f
C5209 net20 _419_/a_1000_472# 0.022734f
C5210 _078_ _083_ 0.01015f
C5211 FILLER_0_21_142/a_484_472# _140_ 0.011035f
C5212 state\[2\] state\[1\] 0.229832f
C5213 net15 ctln[8] 0.205163f
C5214 net52 _029_ 0.03261f
C5215 _144_ FILLER_0_22_128/a_3172_472# 0.001287f
C5216 _069_ vss 0.323941f
C5217 result[9] FILLER_0_24_274/a_572_375# 0.003576f
C5218 FILLER_0_13_212/a_572_375# net79 0.009626f
C5219 _091_ _098_ 1.501073f
C5220 FILLER_0_16_107/a_572_375# _093_ 0.002827f
C5221 FILLER_0_24_96/a_124_375# vdd 0.029269f
C5222 net62 FILLER_0_13_212/a_1020_375# 0.001597f
C5223 _095_ vdd 1.051346f
C5224 output21/a_224_472# output35/a_224_472# 0.001374f
C5225 output12/a_224_472# net59 0.015069f
C5226 net49 _029_ 0.004408f
C5227 _158_ _157_ 0.001663f
C5228 _114_ _250_/a_36_68# 0.017773f
C5229 net4 FILLER_0_3_221/a_1020_375# 0.006974f
C5230 mask\[7\] _435_/a_1204_472# 0.007888f
C5231 result[8] _422_/a_448_472# 0.002989f
C5232 _394_/a_718_524# cal_count\[1\] 0.009499f
C5233 mask\[3\] FILLER_0_17_218/a_484_472# 0.017442f
C5234 net63 FILLER_0_15_212/a_124_375# 0.001597f
C5235 output12/a_224_472# FILLER_0_0_198/a_124_375# 0.00515f
C5236 output9/a_224_472# net82 0.003636f
C5237 _450_/a_36_151# output6/a_224_472# 0.134892f
C5238 _261_/a_36_160# net47 0.010976f
C5239 _089_ _270_/a_36_472# 0.00437f
C5240 _036_ vdd 0.364747f
C5241 net57 _061_ 0.127011f
C5242 _143_ net80 0.023487f
C5243 FILLER_0_7_72/a_2276_472# _077_ 0.00475f
C5244 output26/a_224_472# vdd 0.047141f
C5245 mask\[5\] FILLER_0_19_171/a_1380_472# 0.007596f
C5246 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_124_375# 0.001597f
C5247 _326_/a_36_160# _077_ 0.00419f
C5248 net57 _311_/a_66_473# 0.013777f
C5249 FILLER_0_12_220/a_124_375# vdd -0.008946f
C5250 FILLER_0_12_136/a_572_375# _427_/a_1308_423# 0.001238f
C5251 net23 FILLER_0_22_128/a_3172_472# 0.015058f
C5252 result[7] net18 0.098317f
C5253 FILLER_0_18_139/a_36_472# vss 0.007877f
C5254 FILLER_0_18_139/a_484_472# vdd 0.003106f
C5255 FILLER_0_4_123/a_124_375# _370_/a_124_24# 0.007188f
C5256 FILLER_0_5_109/a_124_375# FILLER_0_4_107/a_484_472# 0.001684f
C5257 output8/a_224_472# net58 0.018549f
C5258 _165_ _220_/a_67_603# 0.004199f
C5259 _057_ _058_ 0.098076f
C5260 FILLER_0_9_72/a_932_472# _439_/a_36_151# 0.001723f
C5261 FILLER_0_21_125/a_36_472# mask\[7\] 0.00344f
C5262 FILLER_0_15_282/a_36_472# net18 0.036858f
C5263 fanout65/a_36_113# net5 0.027955f
C5264 _126_ _125_ 0.032402f
C5265 FILLER_0_22_177/a_124_375# vss 0.002674f
C5266 FILLER_0_22_177/a_572_375# vdd -0.003694f
C5267 FILLER_0_18_107/a_484_472# mask\[9\] 0.001955f
C5268 FILLER_0_15_282/a_572_375# result[3] 0.038939f
C5269 net19 _419_/a_2248_156# 0.012726f
C5270 _390_/a_692_472# _136_ 0.004782f
C5271 net20 FILLER_0_12_220/a_124_375# 0.003161f
C5272 trim_val\[3\] _441_/a_1308_423# 0.001312f
C5273 _050_ net23 0.003752f
C5274 _426_/a_1308_423# net64 0.021119f
C5275 FILLER_0_4_107/a_124_375# _160_ 0.005906f
C5276 net31 vss 0.562041f
C5277 FILLER_0_9_28/a_1380_472# _054_ 0.004017f
C5278 result[8] _108_ 0.007884f
C5279 net71 _437_/a_2560_156# 0.037081f
C5280 _081_ _265_/a_468_472# 0.005156f
C5281 _435_/a_2560_156# vdd 0.001372f
C5282 _435_/a_2665_112# vss 0.002665f
C5283 result[0] result[1] 0.06045f
C5284 net80 _146_ 0.021227f
C5285 net63 result[8] 0.013631f
C5286 result[4] net60 0.244453f
C5287 _449_/a_448_472# vdd 0.007757f
C5288 _449_/a_36_151# vss 0.014774f
C5289 FILLER_0_5_109/a_572_375# FILLER_0_5_117/a_36_472# 0.086635f
C5290 net57 _072_ 0.108982f
C5291 _154_ _365_/a_36_68# 0.02267f
C5292 _091_ _070_ 0.162632f
C5293 net25 _214_/a_36_160# 0.019894f
C5294 FILLER_0_17_200/a_36_472# FILLER_0_18_177/a_2724_472# 0.026657f
C5295 _265_/a_244_68# _082_ 0.031951f
C5296 _443_/a_1308_423# net13 0.004098f
C5297 _443_/a_1000_472# net23 0.034596f
C5298 net72 net55 0.233515f
C5299 net28 vss 0.185012f
C5300 net28 _192_/a_255_603# 0.003166f
C5301 _091_ FILLER_0_15_180/a_124_375# 0.001415f
C5302 _149_ _437_/a_1308_423# 0.015677f
C5303 _026_ _437_/a_36_151# 0.012193f
C5304 FILLER_0_8_127/a_124_375# vss 0.019066f
C5305 vdd output41/a_224_472# 0.003282f
C5306 net44 net67 0.08001f
C5307 fanout80/a_36_113# FILLER_0_15_205/a_36_472# 0.010419f
C5308 _341_/a_49_472# FILLER_0_17_161/a_36_472# 0.079018f
C5309 net34 _146_ 0.004718f
C5310 ctln[1] input5/a_36_113# 0.01908f
C5311 _122_ FILLER_0_6_231/a_124_375# 0.013183f
C5312 net27 net75 0.037524f
C5313 FILLER_0_17_200/a_572_375# net63 0.007512f
C5314 trim_val\[4\] _443_/a_2560_156# 0.049334f
C5315 _448_/a_2560_156# trim_mask\[4\] 0.001306f
C5316 net41 _446_/a_2665_112# 0.004501f
C5317 cal_itt\[2\] vss 0.249871f
C5318 net39 trim[1] 0.115976f
C5319 net21 FILLER_0_12_196/a_36_472# 0.001298f
C5320 FILLER_0_14_263/a_124_375# output30/a_224_472# 0.011584f
C5321 _164_ FILLER_0_6_37/a_36_472# 0.001049f
C5322 _402_/a_1296_93# vdd 0.017239f
C5323 _077_ FILLER_0_7_72/a_932_472# 0.001315f
C5324 _083_ _263_/a_224_472# 0.003191f
C5325 _415_/a_2665_112# vss 0.015461f
C5326 net29 _006_ 0.135646f
C5327 net75 fanout75/a_36_113# 0.035159f
C5328 net50 FILLER_0_8_24/a_572_375# 0.001597f
C5329 FILLER_0_12_236/a_36_472# vdd 0.086431f
C5330 FILLER_0_12_236/a_572_375# vss 0.025768f
C5331 trim[0] _064_ 0.014422f
C5332 _132_ _428_/a_796_472# 0.001472f
C5333 output37/a_224_472# vdd 0.082206f
C5334 FILLER_0_16_107/a_572_375# _136_ 0.006445f
C5335 FILLER_0_14_91/a_572_375# vss 0.054783f
C5336 FILLER_0_14_91/a_36_472# vdd 0.08739f
C5337 FILLER_0_15_282/a_484_472# _417_/a_36_151# 0.059367f
C5338 FILLER_0_15_282/a_36_472# _417_/a_448_472# 0.011962f
C5339 _077_ _256_/a_1612_497# 0.002724f
C5340 fanout82/a_36_113# _316_/a_848_380# 0.001292f
C5341 net63 FILLER_0_22_177/a_1468_375# 0.005028f
C5342 _385_/a_36_68# vdd 0.01625f
C5343 net52 _163_ 0.00157f
C5344 FILLER_0_21_142/a_484_472# FILLER_0_21_150/a_36_472# 0.013277f
C5345 _442_/a_1308_423# _031_ 0.003679f
C5346 FILLER_0_21_28/a_1380_472# vdd 0.007073f
C5347 _053_ net22 0.039386f
C5348 net72 net17 0.004503f
C5349 ctlp[2] _009_ 0.220631f
C5350 net50 FILLER_0_2_93/a_36_472# 0.008147f
C5351 FILLER_0_9_28/a_932_472# net16 0.017841f
C5352 _423_/a_1308_423# _012_ 0.01389f
C5353 FILLER_0_1_192/a_124_375# net21 0.067765f
C5354 FILLER_0_13_100/a_124_375# _043_ 0.010818f
C5355 _016_ _127_ 0.01898f
C5356 net20 FILLER_0_12_236/a_36_472# 0.003143f
C5357 net27 _004_ 0.080285f
C5358 _104_ _422_/a_2665_112# 0.040586f
C5359 _144_ mask\[4\] 0.268823f
C5360 net36 _438_/a_36_151# 0.076525f
C5361 output15/a_224_472# net52 0.007862f
C5362 net15 fanout50/a_36_160# 0.029852f
C5363 _001_ cal_itt\[0\] 0.004843f
C5364 _429_/a_36_151# net79 0.02414f
C5365 net52 FILLER_0_11_78/a_124_375# 0.006273f
C5366 net62 _429_/a_448_472# 0.002713f
C5367 _161_ FILLER_0_6_177/a_484_472# 0.001723f
C5368 net36 _451_/a_3129_107# 0.013154f
C5369 net15 _110_ 0.016359f
C5370 net54 _437_/a_2665_112# 0.061157f
C5371 _427_/a_1000_472# net23 0.003046f
C5372 net47 FILLER_0_5_136/a_124_375# 0.010674f
C5373 FILLER_0_21_28/a_1468_375# _424_/a_36_151# 0.059049f
C5374 net50 trim_mask\[2\] 0.267074f
C5375 net76 FILLER_0_5_198/a_484_472# 0.00169f
C5376 net79 net18 0.222939f
C5377 output47/a_224_472# _398_/a_36_113# 0.001605f
C5378 output15/a_224_472# net49 0.005626f
C5379 net58 _412_/a_2560_156# 0.005111f
C5380 _332_/a_36_472# vdd 0.017097f
C5381 output23/a_224_472# _210_/a_67_603# 0.021084f
C5382 net62 result[3] 0.451989f
C5383 FILLER_0_14_50/a_36_472# cal_count\[1\] 0.030015f
C5384 _068_ _315_/a_36_68# 0.003516f
C5385 _144_ mask\[9\] 0.001909f
C5386 _430_/a_2665_112# mask\[2\] 0.028551f
C5387 net64 FILLER_0_8_239/a_36_472# 0.002666f
C5388 net77 vss 0.327705f
C5389 net76 FILLER_0_2_177/a_484_472# 0.012872f
C5390 result[1] _416_/a_1000_472# 0.001529f
C5391 net28 _416_/a_2248_156# 0.001082f
C5392 FILLER_0_10_247/a_124_375# fanout79/a_36_160# 0.010334f
C5393 _077_ FILLER_0_10_78/a_484_472# 0.002486f
C5394 FILLER_0_10_78/a_36_472# vdd 0.001865f
C5395 FILLER_0_18_2/a_1828_472# net38 0.006713f
C5396 mask\[4\] net23 0.111873f
C5397 FILLER_0_16_57/a_1020_375# _176_ 0.006334f
C5398 _053_ FILLER_0_7_72/a_1468_375# 0.014569f
C5399 ctln[2] net19 0.073057f
C5400 net53 _451_/a_836_156# 0.006521f
C5401 result[6] _421_/a_1204_472# 0.005361f
C5402 _119_ _069_ 0.00226f
C5403 _077_ _374_/a_36_68# 0.012411f
C5404 _131_ FILLER_0_17_56/a_36_472# 0.001491f
C5405 _065_ net16 0.068602f
C5406 _142_ net23 0.037306f
C5407 net28 _195_/a_67_603# 0.012984f
C5408 trim[4] _054_ 0.005511f
C5409 _075_ cal_itt\[3\] 0.731221f
C5410 _370_/a_124_24# _081_ 0.015048f
C5411 net54 net14 0.121719f
C5412 _182_ _180_ 0.090106f
C5413 _412_/a_448_472# en 0.011052f
C5414 _275_/a_224_472# _069_ 0.004466f
C5415 _411_/a_36_151# net8 0.012319f
C5416 FILLER_0_14_81/a_36_472# vss 0.007047f
C5417 net60 _418_/a_1308_423# 0.016365f
C5418 ctln[1] net19 0.001327f
C5419 output39/a_224_472# net49 0.039256f
C5420 output29/a_224_472# _044_ 0.087528f
C5421 net60 _006_ 0.006254f
C5422 _115_ _070_ 0.890903f
C5423 _011_ _109_ 0.055905f
C5424 FILLER_0_4_152/a_124_375# vss 0.019426f
C5425 _426_/a_2248_156# vdd 0.003943f
C5426 _439_/a_2665_112# trim_mask\[0\] 0.020363f
C5427 _147_ vdd 0.09215f
C5428 _098_ _438_/a_2665_112# 0.004321f
C5429 FILLER_0_9_290/a_36_472# vss 0.011755f
C5430 _104_ mask\[2\] 0.002737f
C5431 output38/a_224_472# trim[0] 0.026911f
C5432 _176_ FILLER_0_15_59/a_36_472# 0.00622f
C5433 FILLER_0_10_78/a_484_472# _120_ 0.004669f
C5434 net60 _103_ 0.066266f
C5435 _059_ net37 0.011845f
C5436 trim[4] vss 0.033925f
C5437 net79 _417_/a_448_472# 0.028398f
C5438 FILLER_0_16_107/a_124_375# FILLER_0_17_104/a_484_472# 0.001723f
C5439 _077_ _133_ 0.003921f
C5440 output27/a_224_472# FILLER_0_9_282/a_36_472# 0.001711f
C5441 _427_/a_1204_472# net74 0.003057f
C5442 net50 FILLER_0_4_91/a_124_375# 0.022557f
C5443 net55 FILLER_0_17_38/a_484_472# 0.013624f
C5444 net62 _417_/a_1308_423# 0.006676f
C5445 _053_ vdd 1.467835f
C5446 net20 _426_/a_2248_156# 0.007902f
C5447 cal_itt\[3\] calibrate 1.141592f
C5448 _114_ FILLER_0_10_94/a_124_375# 0.040691f
C5449 FILLER_0_4_197/a_124_375# net22 0.00145f
C5450 FILLER_0_7_72/a_2724_472# trim_mask\[0\] 0.006975f
C5451 _335_/a_49_472# _138_ 0.005957f
C5452 FILLER_0_14_107/a_36_472# _451_/a_36_151# 0.001723f
C5453 FILLER_0_6_47/a_2364_375# vss 0.008275f
C5454 FILLER_0_6_47/a_2812_375# vdd 0.002455f
C5455 net73 FILLER_0_17_133/a_124_375# 0.022541f
C5456 _126_ _043_ 0.128227f
C5457 net18 FILLER_0_13_290/a_124_375# 0.007717f
C5458 FILLER_0_15_142/a_572_375# _431_/a_2248_156# 0.001374f
C5459 _068_ FILLER_0_5_148/a_484_472# 0.016952f
C5460 net15 _164_ 0.026132f
C5461 cal_itt\[3\] net21 0.175781f
C5462 trimb[0] net17 0.006176f
C5463 FILLER_0_24_290/a_36_472# FILLER_0_24_274/a_1380_472# 0.013277f
C5464 _285_/a_36_472# net36 0.003032f
C5465 cal_count\[2\] _402_/a_728_93# 0.036871f
C5466 output9/a_224_472# net58 0.050634f
C5467 net31 output31/a_224_472# 0.002146f
C5468 _431_/a_2248_156# FILLER_0_18_139/a_932_472# 0.001148f
C5469 FILLER_0_13_65/a_36_472# vdd 0.005885f
C5470 FILLER_0_4_99/a_124_375# _156_ 0.081915f
C5471 _140_ vss 0.53195f
C5472 _282_/a_36_160# vss 0.005221f
C5473 _415_/a_448_472# FILLER_0_11_282/a_124_375# 0.008952f
C5474 FILLER_0_19_55/a_124_375# FILLER_0_19_47/a_572_375# 0.012001f
C5475 FILLER_0_19_195/a_36_472# FILLER_0_19_187/a_484_472# 0.013276f
C5476 FILLER_0_6_90/a_572_375# net14 0.031929f
C5477 _050_ _436_/a_2248_156# 0.023725f
C5478 fanout71/a_36_113# FILLER_0_19_111/a_484_472# 0.007864f
C5479 net38 net66 0.040578f
C5480 net32 _102_ 0.038622f
C5481 fanout80/a_36_113# _139_ 0.009968f
C5482 _327_/a_36_472# FILLER_0_12_136/a_36_472# 0.096379f
C5483 _395_/a_36_488# _070_ 0.005165f
C5484 _119_ FILLER_0_8_127/a_124_375# 0.013315f
C5485 net35 _098_ 0.017288f
C5486 vss FILLER_0_6_231/a_484_472# 0.005629f
C5487 _421_/a_448_472# vss -0.001027f
C5488 _421_/a_1308_423# vdd 0.021664f
C5489 net38 _067_ 0.062447f
C5490 _411_/a_448_472# net75 0.072712f
C5491 _412_/a_2665_112# net59 0.055415f
C5492 _133_ _120_ 0.003762f
C5493 net67 _450_/a_836_156# 0.008805f
C5494 _104_ _420_/a_2248_156# 0.027923f
C5495 FILLER_0_8_37/a_124_375# _054_ 0.014206f
C5496 _136_ FILLER_0_15_180/a_484_472# 0.002128f
C5497 _424_/a_2665_112# vss 0.013462f
C5498 net26 FILLER_0_23_44/a_1020_375# 0.001646f
C5499 _320_/a_1792_472# state\[1\] 0.001901f
C5500 _210_/a_67_603# _436_/a_2665_112# 0.007103f
C5501 net20 _421_/a_1308_423# 0.012036f
C5502 net55 FILLER_0_17_72/a_572_375# 0.023585f
C5503 _096_ _320_/a_224_472# 0.001285f
C5504 state\[0\] _060_ 0.047136f
C5505 net50 _441_/a_2560_156# 0.008865f
C5506 _443_/a_36_151# _370_/a_848_380# 0.001568f
C5507 _287_/a_36_472# _102_ 0.028733f
C5508 result[9] _417_/a_2248_156# 0.046399f
C5509 FILLER_0_9_28/a_124_375# vdd -0.004893f
C5510 net29 mask\[2\] 0.122202f
C5511 result[5] net18 0.173673f
C5512 net82 FILLER_0_3_212/a_36_472# 0.011542f
C5513 net34 _422_/a_2665_112# 0.006103f
C5514 FILLER_0_16_57/a_484_472# net15 0.008573f
C5515 FILLER_0_1_98/a_124_375# net14 0.049552f
C5516 FILLER_0_8_37/a_124_375# vss 0.00252f
C5517 FILLER_0_8_37/a_572_375# vdd 0.013575f
C5518 FILLER_0_12_136/a_932_472# vss 0.008682f
C5519 FILLER_0_12_136/a_1380_472# vdd 0.006419f
C5520 output35/a_224_472# _204_/a_67_603# 0.012678f
C5521 _449_/a_2248_156# _176_ 0.013753f
C5522 FILLER_0_21_28/a_1916_375# _012_ 0.023886f
C5523 net27 net19 0.036883f
C5524 FILLER_0_5_72/a_36_472# vdd 0.107678f
C5525 FILLER_0_5_72/a_1468_375# vss 0.057097f
C5526 _031_ FILLER_0_2_111/a_484_472# 0.027347f
C5527 net69 FILLER_0_2_111/a_1380_472# 0.021896f
C5528 _050_ FILLER_0_22_128/a_1020_375# 0.002647f
C5529 FILLER_0_5_54/a_124_375# trim_mask\[1\] 0.024065f
C5530 FILLER_0_5_54/a_1468_375# _029_ 0.008339f
C5531 _122_ FILLER_0_8_156/a_484_472# 0.007378f
C5532 FILLER_0_20_87/a_124_375# vdd 0.008846f
C5533 _127_ _017_ 0.005836f
C5534 _449_/a_36_151# _095_ 0.003412f
C5535 _326_/a_36_160# FILLER_0_9_105/a_572_375# 0.005489f
C5536 _114_ FILLER_0_14_107/a_36_472# 0.00191f
C5537 _451_/a_36_151# vss 0.028073f
C5538 _451_/a_448_472# vdd 0.04463f
C5539 FILLER_0_4_197/a_124_375# vdd 0.011327f
C5540 _093_ _013_ 0.064462f
C5541 _446_/a_1000_472# net40 0.0368f
C5542 _426_/a_36_151# FILLER_0_8_247/a_1468_375# 0.059049f
C5543 _247_/a_36_160# _090_ 0.010285f
C5544 vdd _166_ 0.108744f
C5545 net74 _062_ 0.062376f
C5546 output11/a_224_472# _413_/a_2665_112# 0.001492f
C5547 _375_/a_36_68# vdd 0.010344f
C5548 _144_ _022_ 0.139742f
C5549 _430_/a_448_472# net80 0.00896f
C5550 FILLER_0_16_255/a_36_472# vss 0.00184f
C5551 input4/a_36_68# en 0.064323f
C5552 _421_/a_1000_472# net19 0.03394f
C5553 FILLER_0_15_150/a_36_472# vdd 0.088307f
C5554 FILLER_0_18_53/a_124_375# FILLER_0_18_37/a_1468_375# 0.012222f
C5555 _053_ fanout67/a_36_160# 0.05724f
C5556 _008_ _418_/a_1204_472# 0.002933f
C5557 _114_ _311_/a_3220_473# 0.003283f
C5558 FILLER_0_14_91/a_484_472# _043_ 0.00134f
C5559 net54 _148_ 0.098648f
C5560 FILLER_0_11_124/a_124_375# vss 0.017354f
C5561 FILLER_0_11_124/a_36_472# vdd 0.005222f
C5562 _267_/a_1568_472# _055_ 0.001681f
C5563 _098_ net22 0.157058f
C5564 FILLER_0_19_55/a_124_375# net55 0.005311f
C5565 FILLER_0_16_89/a_124_375# _177_ 0.008257f
C5566 mask\[7\] _009_ 0.078131f
C5567 net80 mask\[2\] 0.048734f
C5568 _185_ vdd 0.325358f
C5569 ctln[4] FILLER_0_1_212/a_124_375# 0.008197f
C5570 net43 vss 0.132286f
C5571 FILLER_0_18_2/a_2276_472# net47 0.001369f
C5572 net66 FILLER_0_3_54/a_124_375# 0.038548f
C5573 _345_/a_36_160# vdd 0.100094f
C5574 net22 _205_/a_36_160# 0.109939f
C5575 mask\[4\] FILLER_0_19_155/a_484_472# 0.024522f
C5576 input1/a_36_113# input4/a_36_68# 0.015796f
C5577 FILLER_0_14_91/a_572_375# _095_ 0.011885f
C5578 net75 _074_ 1.343862f
C5579 FILLER_0_12_124/a_36_472# _127_ 0.01468f
C5580 _350_/a_257_69# net23 0.003052f
C5581 _261_/a_36_160# FILLER_0_5_148/a_124_375# 0.005705f
C5582 _056_ net4 0.002408f
C5583 output9/a_224_472# fanout81/a_36_160# 0.012218f
C5584 net79 _284_/a_224_472# 0.009327f
C5585 _431_/a_1204_472# net73 0.026905f
C5586 _419_/a_1000_472# net77 0.001113f
C5587 FILLER_0_18_107/a_36_472# net14 0.005297f
C5588 FILLER_0_4_185/a_36_472# net22 0.006506f
C5589 net81 FILLER_0_15_212/a_932_472# 0.003953f
C5590 FILLER_0_9_223/a_484_472# vdd 0.004285f
C5591 _372_/a_358_69# _163_ 0.001427f
C5592 state\[1\] _043_ 0.1587f
C5593 FILLER_0_21_150/a_36_472# vss 0.012815f
C5594 _326_/a_36_160# _125_ 0.050008f
C5595 _161_ _058_ 0.101968f
C5596 _112_ net59 0.002846f
C5597 _083_ _080_ 0.043927f
C5598 _136_ _138_ 0.186242f
C5599 cal_count\[3\] _390_/a_36_68# 0.003074f
C5600 FILLER_0_9_223/a_484_472# net20 0.002601f
C5601 _128_ _061_ 0.76584f
C5602 vss output30/a_224_472# 0.030732f
C5603 fanout62/a_36_160# _416_/a_36_151# 0.016215f
C5604 _129_ _058_ 0.050726f
C5605 ctlp[2] net33 0.004972f
C5606 FILLER_0_24_63/a_124_375# vss 0.03143f
C5607 net54 FILLER_0_19_134/a_36_472# 0.061344f
C5608 FILLER_0_16_57/a_1020_375# FILLER_0_17_64/a_124_375# 0.026339f
C5609 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_124_375# 0.012001f
C5610 FILLER_0_10_37/a_124_375# net16 0.010358f
C5611 FILLER_0_12_50/a_36_472# vss 0.0027f
C5612 _106_ _008_ 0.034748f
C5613 _093_ FILLER_0_17_72/a_3260_375# 0.011936f
C5614 FILLER_0_16_37/a_124_375# net72 0.013591f
C5615 _428_/a_2665_112# vdd 0.004735f
C5616 output43/a_224_472# net43 0.11662f
C5617 _098_ _433_/a_2665_112# 0.01601f
C5618 fanout53/a_36_160# vdd 0.016868f
C5619 FILLER_0_20_193/a_36_472# net21 0.001099f
C5620 net4 _068_ 0.040977f
C5621 _437_/a_1204_472# net14 0.004949f
C5622 _119_ _324_/a_224_472# 0.00368f
C5623 _394_/a_56_524# vss 0.003797f
C5624 _053_ FILLER_0_7_72/a_1380_472# 0.01339f
C5625 _114_ vss 0.365613f
C5626 net41 net38 0.059214f
C5627 FILLER_0_24_274/a_1380_472# FILLER_0_23_282/a_484_472# 0.058411f
C5628 _070_ net22 0.032551f
C5629 _422_/a_2248_156# _009_ 0.061786f
C5630 _408_/a_56_524# net40 0.001367f
C5631 _407_/a_36_472# vdd 0.095308f
C5632 _121_ _120_ 0.069685f
C5633 vdd cal_count\[0\] 0.491891f
C5634 FILLER_0_8_2/a_124_375# _054_ 0.001055f
C5635 _112_ _122_ 0.120159f
C5636 net36 _094_ 0.086414f
C5637 FILLER_0_11_124/a_36_472# _135_ 0.110114f
C5638 _432_/a_2665_112# _430_/a_36_151# 0.030053f
C5639 _098_ FILLER_0_15_235/a_572_375# 0.001343f
C5640 _016_ _427_/a_796_472# 0.001666f
C5641 output22/a_224_472# net63 0.017997f
C5642 FILLER_0_20_177/a_484_472# _098_ 0.009817f
C5643 net46 net43 0.215092f
C5644 _155_ FILLER_0_4_107/a_124_375# 0.00162f
C5645 FILLER_0_9_28/a_1916_375# _042_ 0.002352f
C5646 _072_ _128_ 0.072191f
C5647 _093_ net71 0.133323f
C5648 _068_ _311_/a_1660_473# 0.003542f
C5649 FILLER_0_14_81/a_36_472# _095_ 0.014706f
C5650 _092_ FILLER_0_17_218/a_36_472# 0.033277f
C5651 FILLER_0_18_177/a_1916_375# net21 0.004339f
C5652 net60 _420_/a_2248_156# 0.035104f
C5653 net15 FILLER_0_5_54/a_572_375# 0.002259f
C5654 _098_ vdd 2.272938f
C5655 FILLER_0_16_73/a_36_472# vdd 0.08735f
C5656 net54 _436_/a_2665_112# 0.042428f
C5657 FILLER_0_5_128/a_484_472# _370_/a_124_24# 0.00171f
C5658 net63 _429_/a_36_151# 0.0144f
C5659 _110_ _012_ 0.046196f
C5660 trim_mask\[1\] FILLER_0_6_47/a_2276_472# 0.006166f
C5661 _424_/a_448_472# _012_ 0.007299f
C5662 FILLER_0_19_55/a_124_375# _216_/a_67_603# 0.003017f
C5663 _091_ net21 0.030022f
C5664 _073_ FILLER_0_3_221/a_1380_472# 0.045839f
C5665 _033_ _444_/a_448_472# 0.047424f
C5666 _205_/a_36_160# vdd 0.016131f
C5667 FILLER_0_8_2/a_124_375# vss 0.003001f
C5668 FILLER_0_8_2/a_36_472# vdd 0.104141f
C5669 _118_ _315_/a_716_497# 0.001968f
C5670 net41 _424_/a_36_151# 0.00413f
C5671 fanout51/a_36_113# FILLER_0_9_72/a_36_472# 0.001391f
C5672 _091_ _333_/a_36_160# 0.031262f
C5673 net19 net18 0.028285f
C5674 _065_ _030_ 0.001499f
C5675 net41 net66 0.08664f
C5676 net67 _439_/a_36_151# 0.136402f
C5677 net20 _098_ 0.087341f
C5678 FILLER_0_9_28/a_36_472# vss -0.001119f
C5679 FILLER_0_13_228/a_36_472# vss 0.006491f
C5680 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_124_375# 0.026339f
C5681 _328_/a_36_113# _132_ 0.006002f
C5682 FILLER_0_19_47/a_572_375# vdd 0.019566f
C5683 FILLER_0_19_47/a_124_375# vss 0.002211f
C5684 FILLER_0_4_185/a_36_472# vdd 0.122463f
C5685 _091_ FILLER_0_19_171/a_932_472# 0.002509f
C5686 net41 _067_ 0.033696f
C5687 fanout66/a_36_113# _441_/a_36_151# 0.032681f
C5688 net18 _416_/a_796_472# 0.007144f
C5689 net19 _196_/a_36_160# 0.027835f
C5690 ctln[5] output13/a_224_472# 0.023159f
C5691 net75 _425_/a_796_472# 0.001146f
C5692 net35 FILLER_0_22_86/a_124_375# 0.01209f
C5693 mask\[8\] FILLER_0_22_86/a_572_375# 0.013048f
C5694 net44 FILLER_0_15_10/a_124_375# 0.009108f
C5695 fanout49/a_36_160# vdd 0.099887f
C5696 FILLER_0_15_10/a_36_472# vss 0.002605f
C5697 FILLER_0_4_144/a_484_472# vss 0.033414f
C5698 net75 _081_ 0.060976f
C5699 _178_ FILLER_0_15_10/a_36_472# 0.001356f
C5700 FILLER_0_7_59/a_124_375# vdd -0.006113f
C5701 FILLER_0_13_212/a_124_375# _043_ 0.011912f
C5702 _105_ _009_ 0.01731f
C5703 _016_ _118_ 0.001549f
C5704 FILLER_0_22_128/a_2812_375# _146_ 0.001336f
C5705 net35 FILLER_0_22_128/a_932_472# 0.007806f
C5706 net17 _452_/a_1293_527# 0.001011f
C5707 _235_/a_67_603# net17 0.018056f
C5708 FILLER_0_5_164/a_572_375# net22 0.002238f
C5709 fanout64/a_36_160# vdd 0.010802f
C5710 _383_/a_36_472# trim_mask\[3\] 0.003193f
C5711 FILLER_0_10_78/a_1020_375# _389_/a_36_148# 0.001335f
C5712 net34 _419_/a_2665_112# 0.001468f
C5713 _387_/a_36_113# vdd 0.041853f
C5714 net59 FILLER_0_3_212/a_124_375# 0.057221f
C5715 FILLER_0_18_177/a_3260_375# net22 0.049279f
C5716 net17 FILLER_0_23_44/a_124_375# 0.007634f
C5717 FILLER_0_18_2/a_1916_375# net55 0.008235f
C5718 _077_ FILLER_0_8_107/a_124_375# 0.010439f
C5719 net65 _386_/a_848_380# 0.00123f
C5720 _412_/a_1308_423# output9/a_224_472# 0.001352f
C5721 _132_ _120_ 0.034714f
C5722 net60 _419_/a_2665_112# 0.059916f
C5723 net75 net65 0.135447f
C5724 _089_ _081_ 0.002206f
C5725 FILLER_0_4_177/a_36_472# trim_val\[4\] 0.001889f
C5726 _444_/a_1000_472# net40 0.038229f
C5727 net54 FILLER_0_22_128/a_1468_375# 0.004731f
C5728 ctlp[7] _025_ 0.007483f
C5729 FILLER_0_17_104/a_1380_472# vss 0.001141f
C5730 _070_ FILLER_0_9_105/a_36_472# 0.023853f
C5731 FILLER_0_8_138/a_36_472# _070_ 0.001342f
C5732 FILLER_0_8_24/a_484_472# net40 0.004383f
C5733 _039_ output6/a_224_472# 0.012051f
C5734 _013_ FILLER_0_17_56/a_572_375# 0.001047f
C5735 result[1] result[2] 0.072492f
C5736 _083_ vss 0.0284f
C5737 _070_ vdd 1.546772f
C5738 FILLER_0_21_125/a_36_472# _354_/a_49_472# 0.063744f
C5739 FILLER_0_18_107/a_1020_375# FILLER_0_17_104/a_1380_472# 0.001597f
C5740 _056_ _058_ 0.988919f
C5741 ctlp[6] FILLER_0_24_130/a_124_375# 0.021926f
C5742 FILLER_0_17_72/a_1380_472# _438_/a_36_151# 0.001221f
C5743 net47 net14 0.033547f
C5744 FILLER_0_7_146/a_36_472# vdd 0.072981f
C5745 FILLER_0_7_146/a_124_375# vss 0.050543f
C5746 FILLER_0_15_180/a_124_375# vdd 0.016985f
C5747 FILLER_0_6_90/a_572_375# _439_/a_2665_112# 0.001646f
C5748 net33 net21 0.052426f
C5749 _009_ _298_/a_224_472# 0.002441f
C5750 FILLER_0_22_86/a_1380_472# FILLER_0_22_107/a_36_472# 0.001963f
C5751 net56 FILLER_0_17_161/a_124_375# 0.001108f
C5752 _144_ net23 0.091811f
C5753 FILLER_0_16_89/a_36_472# _131_ 0.013616f
C5754 net82 net22 1.960347f
C5755 net20 _070_ 0.075448f
C5756 output25/a_224_472# ctlp[8] 0.018544f
C5757 _115_ FILLER_0_10_94/a_36_472# 0.014605f
C5758 net47 _164_ 0.118311f
C5759 FILLER_0_21_28/a_124_375# net40 0.060428f
C5760 FILLER_0_5_128/a_36_472# _360_/a_36_160# 0.195479f
C5761 FILLER_0_12_136/a_484_472# _126_ 0.014541f
C5762 trim_mask\[2\] FILLER_0_3_78/a_124_375# 0.010185f
C5763 _321_/a_170_472# _120_ 0.040613f
C5764 net80 FILLER_0_22_177/a_36_472# 0.018848f
C5765 FILLER_0_18_2/a_1916_375# net17 0.013121f
C5766 net23 _066_ 0.031928f
C5767 _420_/a_36_151# net18 0.001426f
C5768 fanout57/a_36_113# net22 0.024465f
C5769 FILLER_0_14_50/a_124_375# vdd 0.026996f
C5770 FILLER_0_7_72/a_2724_472# FILLER_0_6_90/a_572_375# 0.001684f
C5771 FILLER_0_6_239/a_124_375# _074_ 0.010359f
C5772 output33/a_224_472# vss 0.05089f
C5773 _077_ FILLER_0_10_94/a_484_472# 0.001548f
C5774 net27 output28/a_224_472# 0.011692f
C5775 FILLER_0_17_72/a_2724_472# _131_ 0.004095f
C5776 _176_ _451_/a_3129_107# 0.021559f
C5777 _065_ trim_mask\[3\] 0.020092f
C5778 _028_ _439_/a_36_151# 0.009268f
C5779 _127_ cal_count\[3\] 0.306114f
C5780 FILLER_0_13_65/a_36_472# _449_/a_36_151# 0.001723f
C5781 _130_ vss 0.090346f
C5782 _420_/a_1204_472# _009_ 0.009314f
C5783 net34 FILLER_0_22_177/a_36_472# 0.003953f
C5784 _133_ _125_ 0.014858f
C5785 _068_ _058_ 0.092852f
C5786 net55 vdd 1.248648f
C5787 net68 FILLER_0_8_37/a_36_472# 0.001088f
C5788 _127_ _059_ 0.002878f
C5789 cal_count\[3\] _453_/a_448_472# 0.001494f
C5790 _132_ mask\[8\] 0.029292f
C5791 _095_ _451_/a_36_151# 0.008311f
C5792 _005_ _100_ 0.004305f
C5793 _074_ _251_/a_468_472# 0.001217f
C5794 _035_ _064_ 0.02225f
C5795 _074_ net19 0.035973f
C5796 FILLER_0_5_54/a_1380_472# vss 0.007301f
C5797 _053_ _385_/a_244_472# 0.00134f
C5798 _077_ _122_ 0.144611f
C5799 cal_count\[3\] FILLER_0_11_135/a_36_472# 0.005101f
C5800 FILLER_0_17_72/a_484_472# net36 0.001629f
C5801 FILLER_0_7_104/a_932_472# _154_ 0.002023f
C5802 FILLER_0_9_28/a_484_472# net41 0.042989f
C5803 mask\[9\] _438_/a_1308_423# 0.044336f
C5804 FILLER_0_5_164/a_572_375# vdd 0.0042f
C5805 net74 net14 0.034568f
C5806 _026_ FILLER_0_20_87/a_36_472# 0.004568f
C5807 output39/a_224_472# net40 0.087367f
C5808 _119_ _114_ 0.001581f
C5809 _182_ vss 0.068928f
C5810 net15 FILLER_0_6_47/a_2724_472# 0.006158f
C5811 _114_ _071_ 0.040513f
C5812 _178_ _182_ 0.067534f
C5813 net68 _160_ 0.072339f
C5814 fanout55/a_36_160# net74 0.016856f
C5815 FILLER_0_18_177/a_3260_375# vdd 0.003399f
C5816 output8/a_224_472# FILLER_0_3_221/a_572_375# 0.03228f
C5817 _077_ _227_/a_36_160# 0.012587f
C5818 _449_/a_2560_156# _067_ 0.007511f
C5819 output8/a_224_472# ctln[1] 0.020259f
C5820 _155_ _363_/a_36_68# 0.013915f
C5821 FILLER_0_7_59/a_124_375# fanout67/a_36_160# 0.001597f
C5822 net66 FILLER_0_5_54/a_124_375# 0.002093f
C5823 FILLER_0_11_101/a_36_472# cal_count\[3\] 0.005101f
C5824 FILLER_0_24_63/a_36_472# _423_/a_2665_112# 0.001873f
C5825 net18 _419_/a_448_472# 0.037373f
C5826 net16 FILLER_0_18_37/a_36_472# 0.001132f
C5827 FILLER_0_15_282/a_484_472# _006_ 0.00444f
C5828 _091_ mask\[1\] 0.064614f
C5829 net17 vdd 2.139315f
C5830 net69 _441_/a_1308_423# 0.016223f
C5831 calibrate FILLER_0_9_270/a_124_375# 0.002292f
C5832 trim_val\[1\] vdd 0.173304f
C5833 _201_/a_67_603# _047_ 0.013357f
C5834 trimb[4] net38 0.124219f
C5835 _425_/a_36_151# vss 0.00158f
C5836 _425_/a_448_472# vdd 0.029071f
C5837 mask\[4\] _348_/a_49_472# 0.001241f
C5838 mask\[7\] FILLER_0_22_128/a_3260_375# 0.00186f
C5839 net17 FILLER_0_20_15/a_484_472# 0.011079f
C5840 _156_ _160_ 0.299745f
C5841 FILLER_0_15_116/a_572_375# FILLER_0_14_107/a_1468_375# 0.026339f
C5842 FILLER_0_15_116/a_36_472# FILLER_0_14_107/a_1020_375# 0.001723f
C5843 mask\[7\] net33 0.02491f
C5844 FILLER_0_23_60/a_124_375# FILLER_0_23_44/a_1468_375# 0.012001f
C5845 FILLER_0_24_290/a_36_472# vss 0.007621f
C5846 net53 _427_/a_1308_423# 0.007426f
C5847 output14/a_224_472# vss 0.012129f
C5848 _122_ _120_ 0.143427f
C5849 net57 _067_ 0.018966f
C5850 _248_/a_36_68# _060_ 0.004581f
C5851 net67 FILLER_0_8_37/a_36_472# 0.001479f
C5852 _448_/a_36_151# net12 0.133216f
C5853 _448_/a_1308_423# net22 0.045644f
C5854 _413_/a_2560_156# net59 0.016463f
C5855 _082_ vdd 0.191411f
C5856 _428_/a_2560_156# _043_ 0.009909f
C5857 net82 vdd 1.014512f
C5858 FILLER_0_18_76/a_124_375# _438_/a_36_151# 0.001252f
C5859 _428_/a_36_151# net74 0.020444f
C5860 net50 _439_/a_448_472# 0.020872f
C5861 net52 _439_/a_796_472# 0.003099f
C5862 FILLER_0_21_28/a_3260_375# FILLER_0_21_60/a_36_472# 0.086742f
C5863 _445_/a_2665_112# net49 0.03968f
C5864 _137_ vss 0.343959f
C5865 mask\[9\] net36 1.116767f
C5866 _098_ FILLER_0_16_154/a_572_375# 0.001791f
C5867 fanout57/a_36_113# vdd 0.005473f
C5868 _013_ FILLER_0_18_53/a_572_375# 0.015534f
C5869 _028_ FILLER_0_6_47/a_3260_375# 0.013006f
C5870 net20 net82 0.026007f
C5871 _443_/a_2665_112# _037_ 0.004052f
C5872 _043_ FILLER_0_13_80/a_124_375# 0.013485f
C5873 state\[2\] FILLER_0_13_142/a_1380_472# 0.019965f
C5874 FILLER_0_3_78/a_36_472# vss 0.004461f
C5875 net67 _160_ 0.003659f
C5876 FILLER_0_2_127/a_36_472# vss 0.002567f
C5877 _394_/a_56_524# _095_ 0.10007f
C5878 FILLER_0_22_86/a_124_375# vdd 0.024158f
C5879 FILLER_0_24_63/a_124_375# output26/a_224_472# 0.00515f
C5880 _132_ FILLER_0_14_107/a_1020_375# 0.029702f
C5881 _152_ _058_ 0.00259f
C5882 _114_ _095_ 0.001338f
C5883 _154_ net14 0.02512f
C5884 net63 FILLER_0_18_177/a_484_472# 0.061539f
C5885 output42/a_224_472# net6 0.010571f
C5886 FILLER_0_22_128/a_932_472# vdd 0.004405f
C5887 FILLER_0_22_128/a_484_472# vss 0.002338f
C5888 mask\[6\] _146_ 0.181681f
C5889 _216_/a_67_603# vdd 0.030831f
C5890 _035_ output38/a_224_472# 0.091395f
C5891 net32 result[7] 0.103491f
C5892 _049_ vss 0.026036f
C5893 net27 _426_/a_796_472# 0.001678f
C5894 net15 fanout72/a_36_113# 0.010284f
C5895 mask\[5\] FILLER_0_19_187/a_124_375# 0.007169f
C5896 FILLER_0_5_117/a_124_375# _086_ 0.003725f
C5897 _346_/a_49_472# _145_ 0.001141f
C5898 net56 FILLER_0_18_139/a_1020_375# 0.018398f
C5899 output27/a_224_472# FILLER_0_8_263/a_36_472# 0.002002f
C5900 FILLER_0_12_20/a_36_472# net6 0.007073f
C5901 _441_/a_2665_112# FILLER_0_3_78/a_572_375# 0.010688f
C5902 _063_ FILLER_0_6_47/a_36_472# 0.007244f
C5903 _116_ _248_/a_36_68# 0.007314f
C5904 _174_ cal_count\[1\] 0.081252f
C5905 output17/a_224_472# net17 0.09023f
C5906 _069_ _098_ 0.029447f
C5907 _088_ FILLER_0_3_172/a_2724_472# 0.005827f
C5908 _111_ vdd 0.3227f
C5909 _053_ FILLER_0_6_47/a_2364_375# 0.007053f
C5910 FILLER_0_16_241/a_36_472# mask\[2\] 0.025337f
C5911 net64 FILLER_0_11_282/a_124_375# 0.023042f
C5912 _411_/a_36_151# _073_ 0.00135f
C5913 net82 FILLER_0_3_172/a_2812_375# 0.010439f
C5914 _140_ _147_ 0.08953f
C5915 _093_ FILLER_0_18_107/a_3260_375# 0.008393f
C5916 FILLER_0_7_72/a_2812_375# net50 0.006598f
C5917 net34 _208_/a_36_160# 0.002666f
C5918 FILLER_0_15_150/a_124_375# net23 0.03361f
C5919 FILLER_0_3_172/a_1916_375# net65 0.003745f
C5920 net9 _082_ 0.001006f
C5921 _446_/a_1308_423# vdd 0.002346f
C5922 net82 net9 0.004599f
C5923 FILLER_0_4_177/a_124_375# _087_ 0.002288f
C5924 output28/a_224_472# net18 0.015144f
C5925 net72 _179_ 0.083699f
C5926 net35 net21 0.001845f
C5927 _316_/a_124_24# _123_ 0.009391f
C5928 FILLER_0_15_116/a_572_375# vdd 0.017636f
C5929 net65 net19 0.044106f
C5930 _076_ _226_/a_1044_68# 0.0023f
C5931 _075_ FILLER_0_7_195/a_124_375# 0.008178f
C5932 _187_ _067_ 0.035532f
C5933 _095_ FILLER_0_15_10/a_36_472# 0.00335f
C5934 _144_ FILLER_0_19_155/a_484_472# 0.006137f
C5935 net57 _066_ 0.069098f
C5936 _448_/a_1308_423# vdd 0.006042f
C5937 net47 _153_ 0.755476f
C5938 _431_/a_1288_156# net73 0.001033f
C5939 _413_/a_36_151# FILLER_0_2_177/a_484_472# 0.006095f
C5940 _028_ FILLER_0_5_72/a_484_472# 0.003042f
C5941 FILLER_0_17_200/a_484_472# vss 0.003134f
C5942 FILLER_0_3_142/a_36_472# net23 0.043034f
C5943 _432_/a_2560_156# _139_ 0.002737f
C5944 _182_ _401_/a_36_68# 0.088487f
C5945 _091_ mask\[0\] 0.04171f
C5946 _442_/a_36_151# net13 0.009343f
C5947 net15 FILLER_0_17_56/a_124_375# 0.001854f
C5948 FILLER_0_5_54/a_572_375# net47 0.009717f
C5949 FILLER_0_7_59/a_572_375# net68 0.005738f
C5950 _075_ net22 0.180274f
C5951 net26 FILLER_0_21_28/a_1828_472# 0.010367f
C5952 net55 _423_/a_2560_156# 0.002265f
C5953 net1 net59 0.920133f
C5954 _176_ FILLER_0_11_101/a_484_472# 0.001777f
C5955 _105_ net33 0.202272f
C5956 net75 FILLER_0_0_232/a_124_375# 0.00217f
C5957 FILLER_0_7_72/a_2276_472# _028_ 0.001777f
C5958 FILLER_0_14_263/a_36_472# vss 0.003195f
C5959 FILLER_0_1_98/a_36_472# FILLER_0_0_96/a_124_375# 0.001684f
C5960 fanout57/a_36_113# FILLER_0_2_165/a_124_375# 0.008057f
C5961 net40 net6 0.00772f
C5962 ctlp[6] mask\[7\] 0.011418f
C5963 net57 net23 0.324262f
C5964 _069_ _070_ 0.257147f
C5965 FILLER_0_16_107/a_124_375# vdd 0.026251f
C5966 _072_ _176_ 0.298077f
C5967 net27 _274_/a_36_68# 0.027359f
C5968 FILLER_0_24_130/a_124_375# vdd 0.027763f
C5969 _386_/a_692_472# _169_ 0.004014f
C5970 _386_/a_848_380# _163_ 0.026484f
C5971 _089_ _414_/a_36_151# 0.039611f
C5972 FILLER_0_7_195/a_124_375# calibrate 0.00576f
C5973 _177_ fanout55/a_36_160# 0.002687f
C5974 FILLER_0_17_72/a_1916_375# vdd 0.002595f
C5975 FILLER_0_17_72/a_1468_375# vss 0.003461f
C5976 trimb[0] trimb[3] 0.549457f
C5977 FILLER_0_12_20/a_124_375# net47 0.047331f
C5978 ctlp[2] vdd 0.617599f
C5979 _003_ _122_ 0.033778f
C5980 result[8] FILLER_0_23_290/a_36_472# 0.001414f
C5981 output9/a_224_472# ctln[2] 0.080206f
C5982 net73 FILLER_0_18_107/a_2724_472# 0.02814f
C5983 FILLER_0_4_107/a_36_472# vdd 0.119007f
C5984 FILLER_0_4_107/a_1468_375# vss 0.055184f
C5985 FILLER_0_2_111/a_484_472# _158_ 0.003604f
C5986 FILLER_0_9_270/a_36_472# vss 0.001642f
C5987 FILLER_0_9_270/a_484_472# vdd 0.006354f
C5988 FILLER_0_5_128/a_572_375# net47 0.010055f
C5989 _008_ ctlp[1] 0.002566f
C5990 FILLER_0_7_195/a_124_375# net21 0.007906f
C5991 calibrate net22 0.036525f
C5992 net52 FILLER_0_2_111/a_1020_375# 0.00245f
C5993 output19/a_224_472# _422_/a_2665_112# 0.024396f
C5994 net20 ctlp[2] 0.254928f
C5995 _412_/a_2248_156# net1 0.044934f
C5996 _424_/a_2248_156# FILLER_0_21_60/a_124_375# 0.001068f
C5997 _432_/a_2665_112# net63 0.067487f
C5998 FILLER_0_2_101/a_124_375# _367_/a_36_68# 0.001176f
C5999 FILLER_0_8_107/a_36_472# FILLER_0_9_105/a_124_375# 0.001684f
C6000 trim_mask\[2\] _167_ 0.027204f
C6001 _091_ FILLER_0_15_212/a_124_375# 0.025529f
C6002 net52 _440_/a_1308_423# 0.047012f
C6003 net61 _421_/a_2665_112# 0.001339f
C6004 net60 _421_/a_1204_472# 0.021679f
C6005 mask\[3\] FILLER_0_18_177/a_572_375# 0.002924f
C6006 net22 net21 1.937266f
C6007 net50 FILLER_0_8_37/a_484_472# 0.003311f
C6008 fanout71/a_36_113# _433_/a_36_151# 0.138322f
C6009 net81 _429_/a_2248_156# 0.017036f
C6010 FILLER_0_11_142/a_572_375# _120_ 0.009014f
C6011 _408_/a_1336_472# vdd 0.040992f
C6012 FILLER_0_23_282/a_484_472# vss 0.005378f
C6013 _141_ FILLER_0_19_155/a_36_472# 0.05777f
C6014 _413_/a_1204_472# vdd 0.001027f
C6015 _114_ _332_/a_36_472# 0.021351f
C6016 net62 _044_ 0.101165f
C6017 FILLER_0_13_142/a_484_472# vss 0.024835f
C6018 net49 _440_/a_1308_423# 0.022006f
C6019 net35 mask\[7\] 0.954332f
C6020 _308_/a_1152_472# trim_mask\[0\] 0.004076f
C6021 _235_/a_67_603# trim_mask\[2\] 0.022726f
C6022 FILLER_0_7_59/a_572_375# net67 0.007538f
C6023 FILLER_0_19_142/a_36_472# vss 0.011026f
C6024 FILLER_0_17_56/a_484_472# FILLER_0_18_61/a_36_472# 0.026657f
C6025 _323_/a_36_113# _015_ 0.003795f
C6026 _040_ vss 0.216709f
C6027 _308_/a_848_380# FILLER_0_10_94/a_484_472# 0.019491f
C6028 cal_count\[3\] _060_ 0.007037f
C6029 _447_/a_1308_423# vdd 0.004739f
C6030 output36/a_224_472# result[2] 0.002356f
C6031 _028_ FILLER_0_7_72/a_932_472# 0.001777f
C6032 _174_ _120_ 0.002521f
C6033 result[2] net30 0.019568f
C6034 FILLER_0_4_197/a_572_375# FILLER_0_5_198/a_484_472# 0.001723f
C6035 _115_ _171_ 0.033359f
C6036 _137_ FILLER_0_16_154/a_1020_375# 0.010692f
C6037 FILLER_0_5_72/a_572_375# _440_/a_36_151# 0.035849f
C6038 _321_/a_170_472# _125_ 0.008492f
C6039 mask\[4\] FILLER_0_18_177/a_2724_472# 0.014625f
C6040 FILLER_0_5_128/a_572_375# net74 0.050735f
C6041 _075_ vdd 0.190898f
C6042 _450_/a_2225_156# net40 0.04513f
C6043 _432_/a_36_151# _337_/a_49_472# 0.002462f
C6044 _447_/a_2665_112# _441_/a_36_151# 0.028591f
C6045 FILLER_0_8_127/a_124_375# _070_ 0.003265f
C6046 result[7] _420_/a_2665_112# 0.039448f
C6047 ctln[1] _411_/a_1000_472# 0.040782f
C6048 FILLER_0_11_101/a_572_375# _134_ 0.0024f
C6049 vss FILLER_0_10_94/a_572_375# 0.013232f
C6050 vdd FILLER_0_10_94/a_36_472# 0.086035f
C6051 _444_/a_448_472# _054_ 0.017318f
C6052 net58 vdd 0.929215f
C6053 result[5] _418_/a_796_472# 0.001983f
C6054 FILLER_0_18_2/a_1380_472# _452_/a_448_472# 0.059367f
C6055 net82 FILLER_0_2_177/a_572_375# 0.003837f
C6056 FILLER_0_7_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001723f
C6057 _189_/a_67_603# net64 0.064691f
C6058 FILLER_0_8_24/a_124_375# _054_ 0.008177f
C6059 mask\[4\] FILLER_0_17_218/a_484_472# 0.001232f
C6060 _261_/a_36_160# FILLER_0_5_136/a_124_375# 0.003477f
C6061 cal_count\[1\] FILLER_0_15_59/a_124_375# 0.010034f
C6062 _256_/a_36_68# net22 0.019035f
C6063 state\[0\] FILLER_0_12_220/a_932_472# 0.001003f
C6064 FILLER_0_8_138/a_36_472# calibrate 0.047835f
C6065 _154_ _153_ 0.719561f
C6066 output8/a_224_472# _411_/a_448_472# 0.010723f
C6067 _116_ cal_count\[3\] 0.384121f
C6068 _449_/a_796_472# net72 0.00138f
C6069 _449_/a_36_151# net55 0.003388f
C6070 _091_ FILLER_0_12_220/a_1020_375# 0.001598f
C6071 _025_ _436_/a_796_472# 0.026852f
C6072 _187_ net41 0.002046f
C6073 calibrate vdd 0.857987f
C6074 output34/a_224_472# vss 0.011966f
C6075 fanout54/a_36_160# vdd 0.008482f
C6076 _078_ FILLER_0_3_221/a_124_375# 0.002694f
C6077 _126_ _250_/a_36_68# 0.022134f
C6078 net64 FILLER_0_15_235/a_124_375# 0.025203f
C6079 mask\[3\] _093_ 2.443356f
C6080 FILLER_0_16_37/a_124_375# vdd 0.038329f
C6081 _444_/a_1308_423# vdd 0.005677f
C6082 result[0] net64 0.09782f
C6083 _289_/a_244_68# _103_ 0.001153f
C6084 _093_ FILLER_0_19_111/a_484_472# 0.001009f
C6085 cal_count\[3\] _408_/a_718_524# 0.005968f
C6086 _238_/a_67_603# net50 0.002229f
C6087 FILLER_0_10_256/a_124_375# vdd 0.041848f
C6088 FILLER_0_8_24/a_572_375# vdd 0.011353f
C6089 fanout59/a_36_160# vss 0.010949f
C6090 mask\[7\] net22 0.275179f
C6091 net20 calibrate 0.044792f
C6092 net21 vdd 1.653552f
C6093 result[8] FILLER_0_24_274/a_932_472# 0.005458f
C6094 FILLER_0_7_72/a_572_375# FILLER_0_6_47/a_3260_375# 0.026339f
C6095 _106_ fanout63/a_36_160# 0.00715f
C6096 _028_ FILLER_0_7_59/a_572_375# 0.00133f
C6097 _333_/a_36_160# vdd 0.107883f
C6098 FILLER_0_16_73/a_484_472# cal_count\[1\] 0.001135f
C6099 net50 fanout68/a_36_113# 0.020067f
C6100 net38 _452_/a_36_151# 0.010095f
C6101 FILLER_0_4_49/a_124_375# net68 0.008422f
C6102 _371_/a_36_113# _370_/a_124_24# 0.008354f
C6103 _415_/a_1000_472# vdd 0.002497f
C6104 _438_/a_448_472# net14 0.020612f
C6105 FILLER_0_2_93/a_572_375# vss 0.055237f
C6106 _072_ _267_/a_36_472# 0.024239f
C6107 net10 ctln[1] 0.029592f
C6108 _413_/a_448_472# net82 0.004927f
C6109 cal_count\[3\] _118_ 0.009058f
C6110 FILLER_0_19_171/a_932_472# vdd 0.011399f
C6111 FILLER_0_19_171/a_484_472# vss 0.001913f
C6112 _144_ _340_/a_36_160# 0.008886f
C6113 result[8] net33 0.474056f
C6114 ctln[7] FILLER_0_0_130/a_36_472# 0.012298f
C6115 trim[4] FILLER_0_8_2/a_36_472# 0.019134f
C6116 mask\[8\] _437_/a_1308_423# 0.001928f
C6117 _288_/a_224_472# _006_ 0.001278f
C6118 FILLER_0_18_171/a_124_375# vss 0.048769f
C6119 result[9] net61 0.014374f
C6120 net57 FILLER_0_3_142/a_36_472# 0.002298f
C6121 _118_ _059_ 0.022651f
C6122 net23 FILLER_0_5_148/a_572_375# 0.039975f
C6123 net44 _452_/a_3129_107# 0.067848f
C6124 net60 result[3] 0.001124f
C6125 fanout56/a_36_113# vss 0.03072f
C6126 _103_ _288_/a_224_472# 0.002992f
C6127 net58 net9 0.018829f
C6128 trim_mask\[2\] vdd 0.376424f
C6129 FILLER_0_21_28/a_124_375# FILLER_0_20_15/a_1468_375# 0.026339f
C6130 net47 FILLER_0_5_148/a_36_472# 0.004409f
C6131 FILLER_0_6_239/a_36_472# _122_ 0.01785f
C6132 _024_ FILLER_0_22_177/a_36_472# 0.003242f
C6133 FILLER_0_2_93/a_124_375# _441_/a_2665_112# 0.006271f
C6134 net16 _446_/a_2665_112# 0.045966f
C6135 _140_ _098_ 0.647503f
C6136 _282_/a_36_160# _098_ 0.00388f
C6137 _055_ _310_/a_49_472# 0.00384f
C6138 _016_ net74 0.568682f
C6139 net81 _005_ 0.003646f
C6140 FILLER_0_23_44/a_1468_375# vdd -0.013698f
C6141 _028_ _133_ 0.007084f
C6142 net15 _441_/a_448_472# 0.049213f
C6143 _143_ FILLER_0_17_161/a_36_472# 0.00363f
C6144 _119_ FILLER_0_4_107/a_1468_375# 0.001695f
C6145 FILLER_0_18_209/a_572_375# _201_/a_67_603# 0.008812f
C6146 _408_/a_728_93# cal_count\[2\] 0.001568f
C6147 FILLER_0_7_59/a_572_375# FILLER_0_6_47/a_1916_375# 0.05841f
C6148 net12 vss 0.043754f
C6149 FILLER_0_16_89/a_1468_375# FILLER_0_17_72/a_3260_375# 0.026339f
C6150 FILLER_0_16_89/a_484_472# FILLER_0_17_72/a_2364_375# 0.001723f
C6151 mask\[1\] net22 0.029526f
C6152 _440_/a_2248_156# net47 0.017063f
C6153 FILLER_0_5_117/a_124_375# _163_ 0.003096f
C6154 FILLER_0_18_61/a_36_472# FILLER_0_18_53/a_484_472# 0.013276f
C6155 _363_/a_36_68# FILLER_0_7_104/a_572_375# 0.002308f
C6156 _418_/a_36_151# vss 0.041728f
C6157 FILLER_0_14_107/a_932_472# vdd 0.006908f
C6158 FILLER_0_14_107/a_484_472# vss -0.001894f
C6159 _448_/a_448_472# FILLER_0_2_177/a_36_472# 0.001927f
C6160 _448_/a_36_151# FILLER_0_2_177/a_484_472# 0.059367f
C6161 _114_ FILLER_0_12_136/a_1380_472# 0.003953f
C6162 FILLER_0_3_172/a_2812_375# net21 0.015743f
C6163 clk vdd 0.053789f
C6164 _056_ FILLER_0_12_196/a_124_375# 0.027077f
C6165 FILLER_0_22_177/a_1468_375# net33 0.017455f
C6166 _433_/a_1308_423# _022_ 0.015376f
C6167 fanout66/a_36_113# _030_ 0.038252f
C6168 cal_itt\[3\] _162_ 0.141474f
C6169 FILLER_0_16_255/a_124_375# net30 0.001055f
C6170 FILLER_0_17_200/a_36_472# _093_ 0.005101f
C6171 FILLER_0_21_286/a_124_375# vss 0.005049f
C6172 FILLER_0_21_286/a_572_375# vdd 0.03062f
C6173 FILLER_0_17_72/a_2364_375# _150_ 0.001083f
C6174 FILLER_0_15_116/a_124_375# _095_ 0.002659f
C6175 cal_itt\[2\] _082_ 0.032565f
C6176 _445_/a_1308_423# net17 0.002172f
C6177 mask\[5\] FILLER_0_20_169/a_124_375# 0.011078f
C6178 _412_/a_2560_156# net18 0.015371f
C6179 _437_/a_2665_112# FILLER_0_22_107/a_484_472# 0.007376f
C6180 _290_/a_224_472# net18 0.00868f
C6181 _120_ _450_/a_3129_107# 0.001598f
C6182 cal_itt\[2\] net82 0.663246f
C6183 output20/a_224_472# ctlp[2] 0.085373f
C6184 net50 _220_/a_67_603# 0.005566f
C6185 FILLER_0_21_28/a_572_375# FILLER_0_20_31/a_124_375# 0.026339f
C6186 fanout81/a_36_160# vdd 0.095319f
C6187 FILLER_0_7_72/a_572_375# FILLER_0_5_72/a_484_472# 0.001512f
C6188 net50 FILLER_0_7_59/a_36_472# 0.01018f
C6189 _077_ _057_ 0.584179f
C6190 _144_ _348_/a_49_472# 0.037768f
C6191 FILLER_0_18_2/a_3260_375# vdd 0.046682f
C6192 _053_ FILLER_0_7_146/a_124_375# 0.005844f
C6193 net20 _256_/a_36_68# 0.02797f
C6194 _132_ _043_ 0.038747f
C6195 _431_/a_2248_156# _427_/a_36_151# 0.001081f
C6196 _402_/a_728_93# _180_ 0.008035f
C6197 FILLER_0_3_54/a_36_472# _381_/a_36_472# 0.010679f
C6198 mask\[5\] _201_/a_67_603# 0.001222f
C6199 FILLER_0_18_61/a_124_375# vdd 0.022663f
C6200 _136_ FILLER_0_16_154/a_1380_472# 0.006517f
C6201 net62 FILLER_0_15_212/a_1468_375# 0.001106f
C6202 _334_/a_36_160# vss 0.002713f
C6203 _428_/a_1000_472# _131_ 0.035998f
C6204 net52 _037_ 0.103749f
C6205 _324_/a_224_472# _070_ 0.00142f
C6206 mask\[7\] vdd 1.098711f
C6207 net40 trim[3] 0.084824f
C6208 net70 net14 0.106631f
C6209 FILLER_0_14_81/a_36_472# net55 0.015878f
C6210 FILLER_0_16_89/a_1380_472# _040_ 0.008446f
C6211 vdd FILLER_0_4_91/a_124_375# 0.019812f
C6212 _074_ FILLER_0_6_231/a_572_375# 0.009029f
C6213 FILLER_0_8_247/a_36_472# _316_/a_124_24# 0.001386f
C6214 net15 cal_count\[3\] 0.045013f
C6215 _327_/a_36_472# vdd 0.00142f
C6216 _155_ _156_ 0.037229f
C6217 net76 net59 3.439686f
C6218 cal_count\[3\] FILLER_0_11_78/a_36_472# 0.031399f
C6219 ctlp[1] FILLER_0_24_274/a_1020_375# 0.004803f
C6220 FILLER_0_3_172/a_484_472# net22 0.012284f
C6221 _427_/a_36_151# _043_ 0.002267f
C6222 _438_/a_2665_112# FILLER_0_19_111/a_124_375# 0.006271f
C6223 _094_ _418_/a_2560_156# 0.011088f
C6224 net16 trim_mask\[1\] 0.007065f
C6225 _422_/a_796_472# mask\[7\] 0.001755f
C6226 output16/a_224_472# net16 0.054603f
C6227 net5 vss 0.326032f
C6228 _086_ _267_/a_1120_472# 0.004245f
C6229 net44 _054_ 0.003562f
C6230 _301_/a_36_472# net25 0.003165f
C6231 _003_ FILLER_0_5_181/a_36_472# 0.003545f
C6232 _076_ FILLER_0_6_231/a_572_375# 0.001647f
C6233 net23 _348_/a_49_472# 0.0037f
C6234 FILLER_0_6_177/a_36_472# net47 0.011891f
C6235 net75 net48 0.10167f
C6236 output18/a_224_472# net33 0.135766f
C6237 net36 net23 0.028202f
C6238 FILLER_0_11_78/a_572_375# _389_/a_36_148# 0.021545f
C6239 _105_ net22 0.01308f
C6240 _096_ _335_/a_49_472# 0.00151f
C6241 _077_ FILLER_0_9_28/a_2364_375# 0.00397f
C6242 _321_/a_3662_472# _176_ 0.002006f
C6243 _150_ _356_/a_36_472# 0.007271f
C6244 _164_ _381_/a_36_472# 0.007224f
C6245 FILLER_0_16_37/a_36_472# cal_count\[2\] 0.008691f
C6246 _250_/a_36_68# state\[1\] 0.103037f
C6247 net75 FILLER_0_8_247/a_1020_375# 0.009573f
C6248 FILLER_0_5_181/a_124_375# net22 0.00205f
C6249 _408_/a_728_93# _043_ 0.029183f
C6250 _436_/a_2665_112# FILLER_0_22_128/a_572_375# 0.001092f
C6251 _436_/a_2560_156# FILLER_0_22_128/a_124_375# 0.001178f
C6252 FILLER_0_15_235/a_484_472# vss 0.003614f
C6253 ctln[3] output10/a_224_472# 0.064347f
C6254 FILLER_0_15_235/a_572_375# mask\[1\] 0.013718f
C6255 _053_ FILLER_0_5_54/a_1380_472# 0.00114f
C6256 FILLER_0_13_142/a_1380_472# _043_ 0.011974f
C6257 FILLER_0_20_177/a_1380_472# vss 0.004504f
C6258 net38 FILLER_0_20_15/a_124_375# 0.012947f
C6259 fanout72/a_36_113# net74 0.02894f
C6260 FILLER_0_5_198/a_124_375# net59 0.00174f
C6261 FILLER_0_9_28/a_2276_472# _453_/a_36_151# 0.059367f
C6262 _428_/a_36_151# net70 0.040167f
C6263 ctlp[3] _422_/a_2560_156# 0.001006f
C6264 net44 vss 0.477283f
C6265 cal_itt\[1\] FILLER_0_3_221/a_1380_472# 0.004939f
C6266 _192_/a_67_603# mask\[1\] 0.020097f
C6267 mask\[1\] vdd 0.741266f
C6268 fanout52/a_36_160# trim_val\[4\] 0.019286f
C6269 output29/a_224_472# _094_ 0.006731f
C6270 FILLER_0_20_169/a_36_472# _339_/a_36_160# 0.001448f
C6271 net36 FILLER_0_15_212/a_484_472# 0.007742f
C6272 fanout80/a_36_113# net81 0.097873f
C6273 fanout81/a_36_160# net9 0.002274f
C6274 _414_/a_796_472# _081_ 0.003538f
C6275 net76 _122_ 0.028025f
C6276 _412_/a_1204_472# net59 0.001824f
C6277 FILLER_0_2_177/a_124_375# net59 0.005212f
C6278 FILLER_0_11_142/a_124_375# vdd 0.010672f
C6279 FILLER_0_17_56/a_36_472# _183_ 0.056523f
C6280 FILLER_0_17_226/a_124_375# net63 0.00507f
C6281 _429_/a_2665_112# FILLER_0_15_212/a_1468_375# 0.010688f
C6282 cal_count\[3\] net51 0.042416f
C6283 _114_ _428_/a_2665_112# 0.002329f
C6284 net80 FILLER_0_20_169/a_124_375# 0.054969f
C6285 FILLER_0_20_15/a_1380_472# vss 0.003678f
C6286 _322_/a_124_24# _129_ 0.017754f
C6287 output21/a_224_472# vss 0.082781f
C6288 FILLER_0_18_107/a_1916_375# vdd 0.018831f
C6289 _098_ FILLER_0_21_150/a_36_472# 0.002964f
C6290 output9/a_224_472# net18 0.114757f
C6291 FILLER_0_5_109/a_484_472# _153_ 0.071582f
C6292 FILLER_0_12_50/a_36_472# cal_count\[0\] 0.001857f
C6293 net24 FILLER_0_22_86/a_1020_375# 0.022658f
C6294 _422_/a_2248_156# vdd 0.005833f
C6295 net20 mask\[1\] 0.09671f
C6296 FILLER_0_7_104/a_124_375# vdd 0.031505f
C6297 net79 FILLER_0_12_220/a_36_472# 0.005464f
C6298 _441_/a_2665_112# vss 0.005169f
C6299 _074_ _375_/a_960_497# 0.004175f
C6300 net55 _424_/a_2665_112# 0.056555f
C6301 _149_ net71 0.827628f
C6302 net27 _091_ 0.023019f
C6303 _430_/a_2248_156# mask\[1\] 0.001498f
C6304 mask\[0\] net22 0.054097f
C6305 _447_/a_796_472# net68 0.001593f
C6306 _447_/a_448_472# _036_ 0.015378f
C6307 FILLER_0_21_28/a_124_375# FILLER_0_19_28/a_36_472# 0.001512f
C6308 FILLER_0_17_56/a_572_375# FILLER_0_15_59/a_36_472# 0.001188f
C6309 input2/a_36_113# vdd 0.096633f
C6310 _122_ FILLER_0_5_198/a_124_375# 0.001352f
C6311 FILLER_0_19_47/a_36_472# net26 0.050805f
C6312 _143_ FILLER_0_18_139/a_1468_375# 0.001097f
C6313 net47 _452_/a_448_472# 0.005335f
C6314 _208_/a_36_160# FILLER_0_22_128/a_2812_375# 0.026361f
C6315 _131_ FILLER_0_17_104/a_484_472# 0.003483f
C6316 _091_ FILLER_0_13_212/a_572_375# 0.022882f
C6317 _441_/a_36_151# net66 0.057618f
C6318 result[8] net35 0.001362f
C6319 net32 _108_ 0.035815f
C6320 FILLER_0_9_142/a_36_472# net23 0.001099f
C6321 net15 _423_/a_1000_472# 0.001786f
C6322 _437_/a_36_151# vss 0.006865f
C6323 _437_/a_448_472# vdd 0.010432f
C6324 net32 net19 0.65591f
C6325 _449_/a_1000_472# _038_ 0.021492f
C6326 FILLER_0_3_172/a_36_472# vss 0.001848f
C6327 FILLER_0_3_172/a_484_472# vdd 0.007258f
C6328 _091_ FILLER_0_10_214/a_124_375# 0.006331f
C6329 FILLER_0_5_198/a_572_375# net21 0.023563f
C6330 FILLER_0_11_109/a_36_472# FILLER_0_10_107/a_124_375# 0.001684f
C6331 output21/a_224_472# _107_ 0.086601f
C6332 net41 _452_/a_36_151# 0.036301f
C6333 output8/a_224_472# net65 0.084944f
C6334 _412_/a_1308_423# vdd 0.003842f
C6335 net16 _444_/a_2665_112# 0.011295f
C6336 fanout71/a_36_113# mask\[9\] 0.044939f
C6337 _052_ FILLER_0_18_37/a_1468_375# 0.001585f
C6338 FILLER_0_21_286/a_484_472# _420_/a_36_151# 0.027236f
C6339 FILLER_0_10_28/a_124_375# net6 0.007948f
C6340 _077_ _439_/a_1308_423# 0.022235f
C6341 cal_count\[3\] _228_/a_36_68# 0.01871f
C6342 _147_ _049_ 0.001131f
C6343 _128_ net23 0.041791f
C6344 _105_ vdd 0.565719f
C6345 FILLER_0_5_72/a_36_472# FILLER_0_5_54/a_1380_472# 0.003468f
C6346 FILLER_0_18_2/a_36_472# cal_count\[2\] 0.001929f
C6347 _017_ net74 0.041246f
C6348 net64 _043_ 0.004021f
C6349 _144_ _433_/a_1308_423# 0.027969f
C6350 _057_ state\[2\] 0.054838f
C6351 vss _416_/a_2665_112# 0.002676f
C6352 vdd _416_/a_2560_156# 0.00165f
C6353 _422_/a_2560_156# _108_ 0.008253f
C6354 trimb[3] vdd 0.283005f
C6355 FILLER_0_5_181/a_124_375# vdd 0.009553f
C6356 FILLER_0_7_195/a_36_472# _055_ 0.03271f
C6357 _360_/a_36_160# vdd 0.006439f
C6358 cal_itt\[3\] _074_ 0.584958f
C6359 vdd output6/a_224_472# 0.009312f
C6360 net80 _138_ 0.002053f
C6361 FILLER_0_4_197/a_1380_472# net76 0.003767f
C6362 FILLER_0_5_88/a_36_472# vss 0.005793f
C6363 _028_ _155_ 0.049284f
C6364 _069_ net21 0.032615f
C6365 FILLER_0_22_177/a_36_472# mask\[6\] 0.006882f
C6366 _130_ FILLER_0_11_124/a_36_472# 0.003572f
C6367 net35 FILLER_0_22_177/a_1468_375# 0.048182f
C6368 mask\[9\] FILLER_0_18_76/a_124_375# 0.004592f
C6369 cal_itt\[3\] _076_ 0.002726f
C6370 _171_ vdd 0.038202f
C6371 net76 FILLER_0_5_206/a_124_375# 0.006974f
C6372 _176_ FILLER_0_11_78/a_484_472# 0.008724f
C6373 FILLER_0_13_206/a_124_375# net79 0.009649f
C6374 net72 _131_ 0.186396f
C6375 _280_/a_224_472# _097_ 0.007508f
C6376 _365_/a_36_68# net14 0.017522f
C6377 FILLER_0_15_150/a_124_375# net36 0.005687f
C6378 FILLER_0_4_49/a_484_472# net49 0.006499f
C6379 output48/a_224_472# vdd 0.038342f
C6380 net54 FILLER_0_18_139/a_124_375# 0.002807f
C6381 FILLER_0_16_73/a_484_472# _175_ 0.036868f
C6382 ctln[6] _037_ 0.031407f
C6383 ctln[4] net59 0.10527f
C6384 FILLER_0_12_124/a_36_472# net74 0.021369f
C6385 _025_ FILLER_0_22_107/a_572_375# 0.090334f
C6386 _148_ FILLER_0_22_107/a_484_472# 0.004761f
C6387 fanout56/a_36_113# _095_ 0.004331f
C6388 _114_ _070_ 0.507391f
C6389 ctln[4] FILLER_0_0_198/a_124_375# 0.015879f
C6390 _413_/a_448_472# net21 0.052657f
C6391 fanout73/a_36_113# net36 0.01199f
C6392 FILLER_0_7_72/a_124_375# net52 0.029774f
C6393 mask\[0\] vdd 0.181371f
C6394 _096_ _136_ 0.022182f
C6395 FILLER_0_14_107/a_1380_472# _043_ 0.001641f
C6396 FILLER_0_13_100/a_36_472# vdd 0.021826f
C6397 FILLER_0_16_57/a_124_375# FILLER_0_18_53/a_484_472# 0.001512f
C6398 FILLER_0_13_100/a_124_375# vss 0.00513f
C6399 FILLER_0_7_72/a_3260_375# FILLER_0_7_104/a_36_472# 0.086905f
C6400 FILLER_0_14_50/a_36_472# FILLER_0_12_50/a_124_375# 0.0027f
C6401 _051_ vss 0.050185f
C6402 result[8] net22 0.278936f
C6403 net10 _411_/a_448_472# 0.010544f
C6404 net20 _298_/a_224_472# 0.001861f
C6405 _033_ _160_ 0.020281f
C6406 _136_ FILLER_0_14_99/a_36_472# 0.01535f
C6407 _430_/a_36_151# _139_ 0.012035f
C6408 _126_ _018_ 0.001243f
C6409 net34 FILLER_0_22_128/a_2276_472# 0.005532f
C6410 result[9] FILLER_0_23_274/a_36_472# 0.0064f
C6411 net58 cal_itt\[2\] 0.003431f
C6412 trim_val\[2\] net68 0.010894f
C6413 _031_ trim_mask\[3\] 0.016747f
C6414 _183_ FILLER_0_18_53/a_36_472# 0.007412f
C6415 _179_ vdd 0.049022f
C6416 _061_ FILLER_0_8_156/a_572_375# 0.023346f
C6417 net20 mask\[0\] 0.103301f
C6418 net58 _415_/a_2665_112# 0.005219f
C6419 output20/a_224_472# mask\[7\] 0.024731f
C6420 _130_ _428_/a_2665_112# 0.001241f
C6421 _420_/a_1000_472# vss 0.002146f
C6422 FILLER_0_20_107/a_124_375# net71 0.03452f
C6423 _013_ _424_/a_1000_472# 0.037585f
C6424 _095_ FILLER_0_14_107/a_484_472# 0.014431f
C6425 net17 net43 0.144179f
C6426 _000_ net59 0.004356f
C6427 _086_ _375_/a_960_497# 0.001454f
C6428 _072_ _246_/a_36_68# 0.064797f
C6429 _435_/a_2665_112# net21 0.067461f
C6430 _394_/a_1336_472# FILLER_0_13_72/a_124_375# 0.001597f
C6431 net4 FILLER_0_12_220/a_484_472# 0.022264f
C6432 net3 vdd 0.118499f
C6433 trimb[3] output17/a_224_472# 0.047604f
C6434 net57 net36 0.087967f
C6435 FILLER_0_10_256/a_124_375# net28 0.034928f
C6436 FILLER_0_17_200/a_572_375# net22 0.047331f
C6437 FILLER_0_10_78/a_572_375# cal_count\[3\] 0.002314f
C6438 fanout65/a_36_113# net64 0.002858f
C6439 trimb[4] FILLER_0_15_2/a_124_375# 0.003305f
C6440 _242_/a_36_160# vdd 0.007995f
C6441 net61 net78 1.588656f
C6442 _444_/a_796_472# net67 0.006859f
C6443 cal_itt\[3\] FILLER_0_5_164/a_484_472# 0.001518f
C6444 FILLER_0_21_125/a_124_375# net54 0.008377f
C6445 _113_ FILLER_0_12_196/a_124_375# 0.001597f
C6446 _090_ FILLER_0_12_196/a_36_472# 0.002321f
C6447 net52 _443_/a_796_472# 0.004334f
C6448 _323_/a_36_113# net4 0.005657f
C6449 net44 _450_/a_1040_527# 0.002267f
C6450 _446_/a_2248_156# net49 0.006196f
C6451 net67 FILLER_0_8_24/a_36_472# 0.001252f
C6452 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_36_472# 0.002296f
C6453 _099_ FILLER_0_15_235/a_572_375# 0.001327f
C6454 net35 _436_/a_448_472# 0.012374f
C6455 _091_ _429_/a_36_151# 0.006557f
C6456 _174_ cal_count\[2\] 0.004821f
C6457 FILLER_0_3_78/a_572_375# _160_ 0.003506f
C6458 net48 _251_/a_468_472# 0.002731f
C6459 _322_/a_848_380# _076_ 0.006699f
C6460 net52 _448_/a_2248_156# 0.002555f
C6461 _233_/a_36_160# FILLER_0_6_37/a_36_472# 0.012692f
C6462 FILLER_0_15_212/a_124_375# vdd -0.004549f
C6463 _099_ vdd 0.326559f
C6464 FILLER_0_4_107/a_572_375# _151_ 0.00162f
C6465 _093_ _438_/a_36_151# 0.088469f
C6466 FILLER_0_20_177/a_1468_375# _434_/a_36_151# 0.001822f
C6467 _273_/a_36_68# _060_ 0.010339f
C6468 net32 _419_/a_448_472# 0.011757f
C6469 FILLER_0_16_154/a_1468_375# vss 0.002071f
C6470 FILLER_0_16_154/a_36_472# vdd 0.00225f
C6471 FILLER_0_4_99/a_36_472# vdd 0.094733f
C6472 FILLER_0_4_99/a_124_375# vss 0.017518f
C6473 _341_/a_49_472# vss 0.003485f
C6474 cal_itt\[3\] _081_ 0.03503f
C6475 net64 FILLER_0_12_236/a_124_375# 0.043517f
C6476 output37/a_224_472# fanout59/a_36_160# 0.021845f
C6477 net27 FILLER_0_9_270/a_124_375# 0.079454f
C6478 trim_mask\[1\] FILLER_0_6_47/a_124_375# 0.005902f
C6479 _055_ vss 0.365503f
C6480 FILLER_0_19_111/a_124_375# vdd 0.005128f
C6481 net20 _099_ 0.011124f
C6482 _421_/a_796_472# _010_ 0.037434f
C6483 FILLER_0_5_198/a_484_472# vss 0.001338f
C6484 FILLER_0_22_86/a_932_472# net14 0.020589f
C6485 _419_/a_2248_156# vdd 0.040646f
C6486 _086_ cal_itt\[3\] 0.046874f
C6487 _386_/a_848_380# net37 0.006086f
C6488 net75 net37 0.07785f
C6489 FILLER_0_18_107/a_572_375# FILLER_0_19_111/a_124_375# 0.058411f
C6490 net19 _420_/a_2665_112# 0.012322f
C6491 _142_ FILLER_0_17_142/a_572_375# 0.012321f
C6492 _232_/a_67_603# FILLER_0_5_54/a_36_472# 0.025312f
C6493 mask\[7\] FILLER_0_22_177/a_124_375# 0.001315f
C6494 net76 FILLER_0_3_172/a_932_472# 0.005391f
C6495 fanout53/a_36_160# _137_ 0.001852f
C6496 _189_/a_67_603# FILLER_0_12_220/a_1468_375# 0.029786f
C6497 _255_/a_224_552# vss 0.001019f
C6498 result[8] vdd 0.590386f
C6499 net50 _029_ 0.025102f
C6500 mask\[8\] _354_/a_257_69# 0.003809f
C6501 _079_ _260_/a_244_472# 0.00325f
C6502 _069_ mask\[1\] 0.029447f
C6503 _126_ vss 0.399848f
C6504 net53 FILLER_0_14_99/a_36_472# 0.004153f
C6505 _414_/a_1000_472# _003_ 0.002053f
C6506 FILLER_0_13_212/a_1468_375# net79 0.009597f
C6507 _089_ net37 0.0326f
C6508 FILLER_0_21_133/a_36_472# net54 0.02286f
C6509 net62 FILLER_0_13_212/a_36_472# 0.015187f
C6510 FILLER_0_4_91/a_572_375# _156_ 0.004958f
C6511 _069_ FILLER_0_11_142/a_124_375# 0.030279f
C6512 net16 _424_/a_36_151# 0.002969f
C6513 net4 FILLER_0_3_221/a_36_472# 0.010517f
C6514 net16 net66 0.030521f
C6515 cal_count\[3\] net47 0.043032f
C6516 mask\[7\] _435_/a_2665_112# 0.030393f
C6517 net20 result[8] 0.014571f
C6518 net69 FILLER_0_2_101/a_124_375# 0.015032f
C6519 FILLER_0_15_142/a_124_375# vdd -0.003809f
C6520 net58 FILLER_0_9_290/a_36_472# 0.005553f
C6521 _394_/a_1936_472# cal_count\[1\] 0.008364f
C6522 net76 FILLER_0_5_181/a_36_472# 0.014784f
C6523 net18 net33 0.001671f
C6524 net57 _128_ 0.040656f
C6525 net63 FILLER_0_15_212/a_1020_375# 0.001012f
C6526 net16 _067_ 0.039705f
C6527 FILLER_0_1_212/a_124_375# vss 0.011796f
C6528 FILLER_0_1_212/a_36_472# vdd 0.10765f
C6529 FILLER_0_8_263/a_36_472# FILLER_0_8_247/a_1380_472# 0.013277f
C6530 _450_/a_1353_112# output6/a_224_472# 0.008732f
C6531 _450_/a_36_151# net6 0.035997f
C6532 FILLER_0_17_200/a_572_375# vdd 0.006861f
C6533 FILLER_0_15_142/a_572_375# vss 0.095176f
C6534 _059_ net47 0.00606f
C6535 net73 _438_/a_2665_112# 0.001708f
C6536 _174_ _043_ 0.964645f
C6537 _176_ _067_ 0.046599f
C6538 FILLER_0_9_28/a_36_472# net17 0.012954f
C6539 net27 FILLER_0_11_282/a_36_472# 0.001526f
C6540 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_572_375# 0.001597f
C6541 output9/a_224_472# net65 0.095296f
C6542 _077_ _161_ 0.023053f
C6543 _115_ _131_ 0.410424f
C6544 FILLER_0_12_220/a_572_375# vss 0.007775f
C6545 FILLER_0_12_220/a_1020_375# vdd -0.014642f
C6546 FILLER_0_16_107/a_124_375# _451_/a_36_151# 0.001597f
C6547 _426_/a_1204_472# calibrate 0.00182f
C6548 FILLER_0_18_139/a_932_472# vss 0.041568f
C6549 _137_ _098_ 0.07262f
C6550 FILLER_0_18_139/a_1380_472# vdd 0.005855f
C6551 net20 FILLER_0_1_212/a_36_472# 0.013846f
C6552 net63 _434_/a_36_151# 0.005153f
C6553 _030_ _157_ 0.011014f
C6554 _270_/a_36_472# net22 0.002857f
C6555 output39/a_224_472# _445_/a_36_151# 0.11862f
C6556 FILLER_0_5_72/a_572_375# _029_ 0.010208f
C6557 FILLER_0_22_177/a_1468_375# vdd -0.007187f
C6558 FILLER_0_15_282/a_484_472# result[3] 0.026996f
C6559 net19 _419_/a_2560_156# 0.003213f
C6560 _077_ _129_ 0.08682f
C6561 net20 FILLER_0_12_220/a_1020_375# 0.047331f
C6562 _447_/a_2665_112# _030_ 0.001226f
C6563 FILLER_0_4_144/a_572_375# _081_ 0.002236f
C6564 FILLER_0_4_144/a_124_375# _152_ 0.007333f
C6565 _426_/a_1000_472# net64 0.008796f
C6566 mask\[2\] FILLER_0_16_154/a_124_375# 0.087247f
C6567 FILLER_0_4_107/a_1020_375# _160_ 0.015684f
C6568 net18 FILLER_0_17_282/a_124_375# 0.048177f
C6569 FILLER_0_4_213/a_124_375# vdd 0.009037f
C6570 _008_ _199_/a_36_160# 0.002015f
C6571 FILLER_0_17_282/a_36_472# net30 0.001189f
C6572 FILLER_0_1_192/a_36_472# net59 0.082738f
C6573 _136_ _438_/a_36_151# 0.030558f
C6574 FILLER_0_17_72/a_572_375# _131_ 0.006224f
C6575 _081_ _265_/a_244_68# 0.03338f
C6576 _204_/a_67_603# vss 0.010366f
C6577 fanout62/a_36_160# net62 0.02201f
C6578 net38 _444_/a_1288_156# 0.001147f
C6579 _449_/a_1308_423# vss 0.027539f
C6580 FILLER_0_21_286/a_572_375# net77 0.044323f
C6581 _153_ _365_/a_36_68# 0.056496f
C6582 net70 FILLER_0_14_123/a_124_375# 0.032077f
C6583 net74 cal_count\[3\] 0.040777f
C6584 output37/a_224_472# net5 0.072504f
C6585 result[1] vss 0.311464f
C6586 mask\[0\] _283_/a_36_472# 0.004645f
C6587 _091_ FILLER_0_15_180/a_36_472# 0.00375f
C6588 net28 mask\[1\] 0.572459f
C6589 _411_/a_1000_472# net65 0.001916f
C6590 _443_/a_2665_112# trim_mask\[4\] 0.013708f
C6591 _077_ FILLER_0_10_78/a_1020_375# 0.001131f
C6592 _026_ _437_/a_1308_423# 0.018479f
C6593 _149_ _437_/a_1000_472# 0.019115f
C6594 FILLER_0_17_161/a_124_375# FILLER_0_16_154/a_932_472# 0.001723f
C6595 net33 _048_ 0.017633f
C6596 net74 _059_ 0.004133f
C6597 net63 FILLER_0_15_205/a_36_472# 0.047903f
C6598 _451_/a_448_472# _040_ 0.026819f
C6599 output36/a_224_472# FILLER_0_14_263/a_124_375# 0.029138f
C6600 net15 FILLER_0_17_64/a_36_472# 0.015524f
C6601 _122_ FILLER_0_6_231/a_36_472# 0.015997f
C6602 ctln[2] vdd 0.245598f
C6603 _129_ _120_ 0.017802f
C6604 FILLER_0_14_263/a_124_375# net30 0.016642f
C6605 _402_/a_56_567# vdd 0.014708f
C6606 _178_ _402_/a_728_93# 0.050963f
C6607 _083_ _082_ 0.018442f
C6608 _077_ FILLER_0_10_78/a_124_375# 0.001886f
C6609 output18/a_224_472# vdd -0.01545f
C6610 net82 _083_ 0.010347f
C6611 net55 _182_ 0.012838f
C6612 net50 FILLER_0_8_24/a_484_472# 0.059367f
C6613 _340_/a_36_160# _348_/a_49_472# 0.001528f
C6614 _132_ _428_/a_1204_472# 0.025555f
C6615 FILLER_0_12_236/a_484_472# vss 0.002739f
C6616 FILLER_0_18_2/a_572_375# trimb[1] 0.010125f
C6617 _137_ FILLER_0_15_180/a_124_375# 0.003108f
C6618 _414_/a_2665_112# vss 0.010021f
C6619 FILLER_0_14_91/a_484_472# vss 0.003257f
C6620 FILLER_0_7_104/a_932_472# _062_ 0.001184f
C6621 net63 FILLER_0_22_177/a_484_472# 0.059367f
C6622 net50 _163_ 0.068547f
C6623 output24/a_224_472# _436_/a_36_151# 0.053592f
C6624 _442_/a_1000_472# _031_ 0.004174f
C6625 FILLER_0_21_28/a_2276_472# vdd 0.002733f
C6626 FILLER_0_21_28/a_1828_472# vss -0.001894f
C6627 _436_/a_448_472# vdd 0.038494f
C6628 FILLER_0_3_221/a_124_375# vss 0.034009f
C6629 _423_/a_1000_472# _012_ 0.013415f
C6630 ctln[1] vdd 0.825166f
C6631 FILLER_0_17_282/a_36_472# _417_/a_36_151# 0.001723f
C6632 FILLER_0_1_192/a_124_375# net11 0.003537f
C6633 net31 _105_ 0.054065f
C6634 trim_mask\[3\] _157_ 0.052956f
C6635 net36 _438_/a_1308_423# 0.012976f
C6636 _069_ mask\[0\] 0.040599f
C6637 output15/a_224_472# net50 0.00515f
C6638 ctln[8] fanout50/a_36_160# 0.004838f
C6639 net15 net52 0.166073f
C6640 FILLER_0_10_78/a_1020_375# _120_ 0.003403f
C6641 net52 FILLER_0_11_78/a_36_472# 0.005678f
C6642 _439_/a_36_151# vss 0.032466f
C6643 _439_/a_448_472# vdd 0.006996f
C6644 net81 _426_/a_448_472# 0.003907f
C6645 _270_/a_36_472# vdd 0.09815f
C6646 FILLER_0_9_28/a_484_472# net16 0.021584f
C6647 _283_/a_36_472# _099_ 0.004667f
C6648 output39/a_224_472# _063_ 0.001019f
C6649 net39 _233_/a_36_160# 0.017979f
C6650 FILLER_0_8_239/a_124_375# _123_ 0.001286f
C6651 _071_ _055_ 0.002641f
C6652 net36 _451_/a_2449_156# 0.016229f
C6653 net20 FILLER_0_3_221/a_572_375# 0.004331f
C6654 result[9] net62 0.339372f
C6655 _427_/a_2248_156# net23 0.033973f
C6656 FILLER_0_21_28/a_2364_375# _424_/a_36_151# 0.059049f
C6657 ctln[1] net20 0.135151f
C6658 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_124_375# 0.003228f
C6659 _095_ FILLER_0_13_100/a_124_375# 0.001989f
C6660 state\[1\] vss 0.294171f
C6661 net15 net49 0.057277f
C6662 _307_/a_234_472# vdd 0.001209f
C6663 FILLER_0_4_144/a_36_472# _443_/a_36_151# 0.00271f
C6664 FILLER_0_14_50/a_36_472# _180_ 0.153222f
C6665 _020_ net70 0.014391f
C6666 FILLER_0_10_78/a_124_375# _120_ 0.006134f
C6667 _176_ net23 0.036283f
C6668 _091_ FILLER_0_18_177/a_484_472# 0.004272f
C6669 _007_ vss 0.017377f
C6670 _321_/a_786_69# net23 0.001073f
C6671 _449_/a_2665_112# cal_count\[3\] 0.001422f
C6672 ctlp[7] net24 0.078667f
C6673 _002_ FILLER_0_3_172/a_2364_375# 0.016984f
C6674 FILLER_0_18_171/a_36_472# FILLER_0_18_177/a_36_472# 0.003468f
C6675 result[1] _416_/a_2248_156# 0.001888f
C6676 FILLER_0_0_266/a_36_472# vdd 0.05043f
C6677 FILLER_0_0_266/a_124_375# vss 0.007654f
C6678 ctln[7] _442_/a_2248_156# 0.006094f
C6679 FILLER_0_7_72/a_36_472# _439_/a_36_151# 0.013806f
C6680 _112_ _425_/a_1000_472# 0.001973f
C6681 FILLER_0_6_239/a_124_375# net37 0.001989f
C6682 FILLER_0_16_57/a_36_472# _176_ 0.075537f
C6683 ctln[2] net9 0.022757f
C6684 net53 _451_/a_3129_107# 0.002806f
C6685 result[6] _421_/a_2665_112# 0.034452f
C6686 _077_ _056_ 1.777574f
C6687 output23/a_224_472# FILLER_0_24_130/a_36_472# 0.001994f
C6688 _126_ _071_ 0.090032f
C6689 _065_ ctln[9] 0.123393f
C6690 net41 net16 2.918931f
C6691 _077_ FILLER_0_7_59/a_484_472# 0.001371f
C6692 _077_ _453_/a_36_151# 0.042928f
C6693 net62 _285_/a_36_472# 0.001288f
C6694 net18 FILLER_0_11_282/a_36_472# 0.048657f
C6695 _354_/a_49_472# vdd -0.001073f
C6696 _069_ FILLER_0_15_212/a_124_375# 0.039975f
C6697 net52 net51 0.091698f
C6698 _370_/a_692_472# _081_ 0.00129f
C6699 _370_/a_848_380# _152_ 0.031499f
C6700 net19 net37 0.030961f
C6701 net7 trim[3] 0.044017f
C6702 _140_ mask\[7\] 0.064343f
C6703 net60 _418_/a_1000_472# 0.007557f
C6704 net39 net49 0.158007f
C6705 net29 _044_ 0.01495f
C6706 FILLER_0_7_72/a_2812_375# vdd 0.02125f
C6707 _062_ net14 0.003317f
C6708 _115_ _076_ 0.051404f
C6709 output20/a_224_472# result[8] 0.038114f
C6710 net24 FILLER_0_23_88/a_36_472# 0.006289f
C6711 _028_ FILLER_0_7_104/a_572_375# 0.003664f
C6712 net82 _425_/a_36_151# 0.002959f
C6713 _426_/a_2665_112# vss 0.006288f
C6714 FILLER_0_16_107/a_484_472# net36 0.003765f
C6715 FILLER_0_1_98/a_124_375# net52 0.001167f
C6716 FILLER_0_9_28/a_1828_472# vdd 0.006263f
C6717 _239_/a_36_160# net68 0.043367f
C6718 _095_ _055_ 0.002933f
C6719 result[0] FILLER_0_9_282/a_124_375# 0.00283f
C6720 _132_ FILLER_0_17_104/a_932_472# 0.006091f
C6721 net79 _417_/a_796_472# 0.001042f
C6722 _077_ _068_ 0.601166f
C6723 net29 _287_/a_244_68# 0.001262f
C6724 net50 FILLER_0_4_91/a_36_472# 0.058499f
C6725 net62 _417_/a_1000_472# 0.005762f
C6726 _003_ _161_ 0.004981f
C6727 _414_/a_36_151# cal_itt\[3\] 0.049033f
C6728 net27 FILLER_0_15_235/a_572_375# 0.001554f
C6729 FILLER_0_17_72/a_3260_375# FILLER_0_17_104/a_36_472# 0.086904f
C6730 output13/a_224_472# FILLER_0_0_130/a_124_375# 0.00363f
C6731 _151_ vdd 0.157764f
C6732 _114_ FILLER_0_10_94/a_36_472# 0.08191f
C6733 ctln[8] net14 0.001447f
C6734 _057_ _043_ 0.02152f
C6735 _120_ _453_/a_36_151# 0.001848f
C6736 FILLER_0_6_47/a_36_472# vdd 0.090192f
C6737 FILLER_0_6_47/a_3260_375# vss 0.061766f
C6738 net15 FILLER_0_15_72/a_572_375# 0.002741f
C6739 FILLER_0_13_290/a_36_472# result[3] 0.001069f
C6740 fanout58/a_36_160# vdd 0.101571f
C6741 net27 vdd 0.88294f
C6742 mask\[8\] FILLER_0_22_107/a_124_375# 0.015331f
C6743 FILLER_0_16_255/a_124_375# _006_ 0.02007f
C6744 FILLER_0_11_135/a_124_375# _120_ 0.017316f
C6745 cal_count\[2\] _402_/a_244_567# 0.004411f
C6746 net31 _099_ 0.01086f
C6747 net36 FILLER_0_15_228/a_36_472# 0.008225f
C6748 _402_/a_728_93# _401_/a_36_68# 0.002178f
C6749 fanout75/a_36_113# vdd 0.028614f
C6750 cal_itt\[3\] _163_ 0.021146f
C6751 FILLER_0_9_28/a_2276_472# _042_ 0.002496f
C6752 net70 _017_ 0.015488f
C6753 net75 net8 0.553872f
C6754 FILLER_0_13_212/a_572_375# vdd 0.001551f
C6755 FILLER_0_13_212/a_124_375# vss 0.007116f
C6756 _093_ _094_ 0.003586f
C6757 _093_ FILLER_0_17_218/a_572_375# 0.0029f
C6758 _429_/a_2248_156# FILLER_0_15_228/a_124_375# 0.030666f
C6759 FILLER_0_6_90/a_484_472# net14 0.014785f
C6760 _050_ _436_/a_2560_156# 0.01099f
C6761 _131_ FILLER_0_14_107/a_1468_375# 0.051201f
C6762 trim[0] net66 0.376153f
C6763 net63 _139_ 0.003073f
C6764 fanout80/a_36_113# _019_ 0.003644f
C6765 _430_/a_2665_112# mask\[3\] 0.002697f
C6766 FILLER_0_11_101/a_572_375# _120_ 0.006382f
C6767 FILLER_0_12_220/a_1468_375# _043_ 0.002509f
C6768 _421_/a_1000_472# vdd 0.006281f
C6769 FILLER_0_20_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001543f
C6770 FILLER_0_17_200/a_572_375# _069_ 0.011239f
C6771 FILLER_0_10_214/a_124_375# vdd 0.018944f
C6772 _446_/a_448_472# net17 0.026011f
C6773 net73 vdd 0.44835f
C6774 net20 fanout75/a_36_113# 0.001027f
C6775 _068_ _120_ 0.447243f
C6776 net57 _443_/a_2248_156# 0.001117f
C6777 _104_ _420_/a_2560_156# 0.002734f
C6778 output22/a_224_472# net22 0.032714f
C6779 _114_ net21 0.022033f
C6780 net31 _419_/a_2248_156# 0.001521f
C6781 net20 FILLER_0_13_212/a_572_375# 0.002085f
C6782 FILLER_0_8_37/a_36_472# _054_ 0.015053f
C6783 net62 _101_ 0.023932f
C6784 FILLER_0_15_142/a_572_375# _095_ 0.003935f
C6785 output33/a_224_472# ctlp[2] 0.00175f
C6786 _091_ _432_/a_2665_112# 0.002978f
C6787 _394_/a_1936_472# _175_ 0.017848f
C6788 _002_ net76 0.213703f
C6789 vdd FILLER_0_21_60/a_572_375# 0.022291f
C6790 vss FILLER_0_21_60/a_124_375# 0.003723f
C6791 net26 FILLER_0_23_44/a_36_472# 0.013977f
C6792 FILLER_0_15_150/a_124_375# _427_/a_2248_156# 0.001221f
C6793 net73 FILLER_0_18_107/a_572_375# 0.008889f
C6794 net55 FILLER_0_17_72/a_1468_375# 0.014449f
C6795 net20 _421_/a_1000_472# 0.012469f
C6796 _422_/a_36_151# _421_/a_2665_112# 0.001725f
C6797 _096_ _320_/a_1120_472# 0.004315f
C6798 fanout53/a_36_160# fanout56/a_36_113# 0.001636f
C6799 FILLER_0_2_111/a_124_375# vdd 0.024756f
C6800 _429_/a_36_151# net22 0.020582f
C6801 _412_/a_36_151# _001_ 0.006762f
C6802 output47/a_224_472# cal_count\[2\] 0.080405f
C6803 _413_/a_36_151# net59 0.02781f
C6804 output44/a_224_472# _452_/a_448_472# 0.004683f
C6805 _440_/a_36_151# vdd 0.117768f
C6806 _091_ _090_ 0.117348f
C6807 result[9] _417_/a_2560_156# 0.00263f
C6808 result[6] result[9] 0.026511f
C6809 _277_/a_36_160# _102_ 0.061995f
C6810 FILLER_0_16_57/a_1380_472# net15 0.017841f
C6811 fanout51/a_36_113# _120_ 0.014349f
C6812 FILLER_0_8_37/a_484_472# vdd 0.009603f
C6813 trim[4] output6/a_224_472# 0.004337f
C6814 net66 _030_ 0.087608f
C6815 _078_ net59 0.168928f
C6816 FILLER_0_21_133/a_124_375# FILLER_0_21_125/a_572_375# 0.012001f
C6817 result[8] _435_/a_2665_112# 0.001855f
C6818 _267_/a_36_472# net23 0.001178f
C6819 fanout74/a_36_113# _443_/a_36_151# 0.032681f
C6820 FILLER_0_21_28/a_2812_375# _012_ 0.016736f
C6821 output47/a_224_472# input3/a_36_113# 0.001371f
C6822 FILLER_0_9_28/a_2364_375# net68 0.019969f
C6823 FILLER_0_5_72/a_484_472# vss 0.003738f
C6824 FILLER_0_5_72/a_932_472# vdd 0.002735f
C6825 _031_ FILLER_0_2_111/a_1380_472# 0.01562f
C6826 FILLER_0_5_128/a_36_472# _163_ 0.009857f
C6827 FILLER_0_12_136/a_932_472# FILLER_0_11_142/a_124_375# 0.001543f
C6828 _098_ FILLER_0_19_171/a_484_472# 0.010731f
C6829 FILLER_0_5_54/a_1020_375# trim_mask\[1\] 0.010745f
C6830 FILLER_0_10_78/a_124_375# FILLER_0_9_72/a_932_472# 0.001543f
C6831 _104_ mask\[3\] 0.078406f
C6832 _086_ _115_ 0.4112f
C6833 FILLER_0_18_171/a_124_375# _098_ 0.032114f
C6834 FILLER_0_1_98/a_36_472# trim_mask\[3\] 0.106084f
C6835 FILLER_0_20_87/a_36_472# vss 0.006244f
C6836 net41 _041_ 0.076779f
C6837 _326_/a_36_160# FILLER_0_9_105/a_484_472# 0.002647f
C6838 state\[1\] _071_ 0.196063f
C6839 fanout63/a_36_160# FILLER_0_15_228/a_124_375# 0.001177f
C6840 _451_/a_1040_527# vdd 0.004038f
C6841 fanout56/a_36_113# _098_ 0.019463f
C6842 _446_/a_2248_156# net40 0.037373f
C6843 _062_ FILLER_0_8_156/a_124_375# 0.008116f
C6844 _247_/a_36_160# _060_ 0.055366f
C6845 FILLER_0_3_204/a_36_472# _088_ 0.004381f
C6846 _426_/a_36_151# FILLER_0_8_247/a_484_472# 0.001723f
C6847 _070_ FILLER_0_10_94/a_572_375# 0.009837f
C6848 net57 _427_/a_2248_156# 0.002706f
C6849 vss _160_ 1.119894f
C6850 _443_/a_36_151# FILLER_0_2_127/a_124_375# 0.073306f
C6851 _412_/a_796_472# net1 0.002922f
C6852 net55 _040_ 0.107198f
C6853 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_124_375# 0.012001f
C6854 _326_/a_36_160# vss 0.002357f
C6855 _162_ vdd 0.073371f
C6856 fanout60/a_36_160# net61 0.001167f
C6857 input4/a_36_68# net4 0.004679f
C6858 _421_/a_2248_156# net19 0.016721f
C6859 fanout70/a_36_113# net74 0.002663f
C6860 FILLER_0_12_2/a_572_375# _450_/a_36_151# 0.001597f
C6861 FILLER_0_15_142/a_36_472# net74 0.003166f
C6862 net57 _176_ 0.192223f
C6863 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1468_375# 0.086742f
C6864 FILLER_0_10_78/a_572_375# net52 0.003311f
C6865 _008_ _418_/a_2665_112# 0.010862f
C6866 net63 FILLER_0_19_187/a_572_375# 0.049706f
C6867 net54 _025_ 0.00573f
C6868 _058_ _313_/a_67_603# 0.010094f
C6869 FILLER_0_18_2/a_124_375# output44/a_224_472# 0.001168f
C6870 _131_ vdd 1.344823f
C6871 mask\[4\] FILLER_0_18_177/a_572_375# 0.015941f
C6872 _078_ _122_ 0.185069f
C6873 _083_ calibrate 0.001446f
C6874 net68 trim_val\[0\] 0.052045f
C6875 _223_/a_36_160# vss 0.007187f
C6876 FILLER_0_7_146/a_124_375# calibrate 0.014163f
C6877 _327_/a_36_472# _428_/a_2248_156# 0.001757f
C6878 _423_/a_36_151# net40 0.004045f
C6879 net56 _433_/a_2665_112# 0.003434f
C6880 net22 _048_ 0.268142f
C6881 input1/a_36_113# en 0.036849f
C6882 _367_/a_36_68# _156_ 0.096366f
C6883 FILLER_0_14_91/a_484_472# _095_ 0.011772f
C6884 output22/a_224_472# vdd 0.111234f
C6885 _059_ FILLER_0_5_148/a_124_375# 0.007657f
C6886 _261_/a_36_160# FILLER_0_5_148/a_36_472# 0.195478f
C6887 _128_ FILLER_0_9_142/a_36_472# 0.005101f
C6888 _091_ _021_ 0.016024f
C6889 net79 _100_ 0.170973f
C6890 net62 _094_ 0.04063f
C6891 FILLER_0_20_87/a_124_375# _437_/a_36_151# 0.059049f
C6892 net15 _052_ 0.001074f
C6893 _086_ _395_/a_36_488# 0.00825f
C6894 _327_/a_36_472# _114_ 0.019746f
C6895 FILLER_0_20_169/a_124_375# mask\[6\] 0.001178f
C6896 _372_/a_1194_69# _163_ 0.001328f
C6897 FILLER_0_18_37/a_124_375# vss 0.002958f
C6898 FILLER_0_18_37/a_572_375# vdd 0.02259f
C6899 FILLER_0_0_130/a_36_472# _442_/a_36_151# 0.001723f
C6900 _429_/a_36_151# vdd 0.076815f
C6901 fanout50/a_36_160# _164_ 0.08721f
C6902 _057_ _267_/a_1568_472# 0.002083f
C6903 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_124_375# 0.012222f
C6904 FILLER_0_18_171/a_36_472# _143_ 0.005167f
C6905 _233_/a_36_160# net47 0.054273f
C6906 FILLER_0_7_195/a_124_375# _074_ 0.019559f
C6907 output36/a_224_472# vss -0.002521f
C6908 _363_/a_244_472# vdd 0.002075f
C6909 _126_ _332_/a_36_472# 0.009299f
C6910 net10 FILLER_0_0_232/a_124_375# 0.022977f
C6911 _238_/a_67_603# vdd 0.004498f
C6912 net18 vdd 1.496006f
C6913 net32 _009_ 0.003756f
C6914 output46/a_224_472# FILLER_0_20_2/a_124_375# 0.030009f
C6915 vss net30 0.17209f
C6916 _095_ state\[1\] 0.069906f
C6917 _129_ _125_ 0.069221f
C6918 net10 net11 0.007522f
C6919 net20 _429_/a_36_151# 0.002103f
C6920 net31 output18/a_224_472# 0.04975f
C6921 _093_ FILLER_0_17_72/a_484_472# 0.008637f
C6922 _196_/a_36_160# vdd 0.106963f
C6923 FILLER_0_7_72/a_932_472# vss 0.002763f
C6924 fanout68/a_36_113# vdd 0.012621f
C6925 net56 vdd 0.277166f
C6926 _074_ net22 0.079421f
C6927 FILLER_0_4_197/a_572_375# net59 0.001512f
C6928 net20 net18 0.025322f
C6929 _396_/a_224_472# _095_ 0.001351f
C6930 _437_/a_2665_112# net14 0.002936f
C6931 _072_ net4 0.097916f
C6932 _263_/a_224_472# net59 0.002558f
C6933 _394_/a_718_524# vss 0.002666f
C6934 _256_/a_1612_497# vss 0.004265f
C6935 FILLER_0_24_63/a_36_472# vss 0.008178f
C6936 _076_ net22 0.03249f
C6937 net20 _411_/a_448_472# 0.002167f
C6938 net67 trim_val\[0\] 0.382079f
C6939 net27 _283_/a_36_472# 0.023243f
C6940 net52 trim_mask\[4\] 0.034276f
C6941 FILLER_0_13_80/a_124_375# vss 0.042254f
C6942 FILLER_0_13_80/a_36_472# vdd 0.087291f
C6943 _422_/a_2560_156# _009_ 0.002551f
C6944 _408_/a_718_524# net40 0.011463f
C6945 _254_/a_448_472# net22 0.009088f
C6946 _077_ FILLER_0_9_28/a_2812_375# 0.006629f
C6947 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_124_375# 0.009654f
C6948 net52 net47 0.039912f
C6949 _187_ net16 0.161791f
C6950 _131_ _135_ 0.068855f
C6951 _098_ FILLER_0_15_235/a_484_472# 0.004898f
C6952 FILLER_0_20_177/a_1380_472# _098_ 0.00679f
C6953 output13/a_224_472# net52 0.018089f
C6954 trimb[3] net43 0.221036f
C6955 _099_ _282_/a_36_160# 0.005808f
C6956 FILLER_0_10_78/a_1380_472# _308_/a_124_24# 0.037778f
C6957 net62 net78 0.001947f
C6958 mask\[4\] _093_ 0.469687f
C6959 net63 FILLER_0_17_226/a_36_472# 0.001822f
C6960 net55 _452_/a_2225_156# 0.022788f
C6961 net49 net47 0.53353f
C6962 _444_/a_448_472# net17 0.022222f
C6963 _068_ _311_/a_2180_473# 0.001454f
C6964 FILLER_0_18_177/a_2812_375# net21 0.048071f
C6965 net60 _420_/a_2560_156# 0.001358f
C6966 net15 FILLER_0_5_54/a_1468_375# 0.039975f
C6967 _394_/a_728_93# _174_ 0.012471f
C6968 _425_/a_36_151# calibrate 0.071513f
C6969 FILLER_0_3_54/a_36_472# _164_ 0.012512f
C6970 FILLER_0_8_24/a_124_375# net17 0.039695f
C6971 _142_ _093_ 0.492191f
C6972 trim_mask\[1\] FILLER_0_6_47/a_3172_472# 0.004605f
C6973 _077_ _308_/a_124_24# 0.018118f
C6974 mask\[3\] net80 0.02972f
C6975 net62 FILLER_0_14_235/a_572_375# 0.017549f
C6976 _033_ _444_/a_796_472# 0.0099f
C6977 _165_ _444_/a_2248_156# 0.006027f
C6978 net44 FILLER_0_8_2/a_36_472# 0.005851f
C6979 _245_/a_672_472# _039_ 0.001025f
C6980 _048_ vdd 0.270091f
C6981 cal_itt\[2\] FILLER_0_3_221/a_572_375# 0.060779f
C6982 FILLER_0_12_136/a_572_375# net23 0.00281f
C6983 ctln[1] cal_itt\[2\] 0.053339f
C6984 net80 _434_/a_448_472# 0.113898f
C6985 _417_/a_36_151# vss 0.040392f
C6986 net19 net8 0.056454f
C6987 _093_ mask\[9\] 0.460108f
C6988 FILLER_0_10_78/a_484_472# vss 0.005854f
C6989 net45 net26 0.002978f
C6990 FILLER_0_4_123/a_124_375# vdd 0.027816f
C6991 FILLER_0_9_28/a_1020_375# FILLER_0_8_37/a_36_472# 0.001723f
C6992 FILLER_0_19_47/a_484_472# vdd 0.001133f
C6993 FILLER_0_19_47/a_36_472# vss 0.001559f
C6994 _220_/a_67_603# vdd 0.020078f
C6995 net18 _416_/a_1204_472# 0.027218f
C6996 _374_/a_36_68# vss 0.047832f
C6997 net75 _425_/a_1204_472# 0.015778f
C6998 mask\[8\] FILLER_0_22_86/a_1468_375# 0.015339f
C6999 net35 FILLER_0_22_86/a_1020_375# 0.010202f
C7000 FILLER_0_7_59/a_36_472# vdd 0.016778f
C7001 FILLER_0_7_59/a_572_375# vss 0.017487f
C7002 FILLER_0_13_212/a_1020_375# _043_ 0.01418f
C7003 _193_/a_36_160# _416_/a_36_151# 0.065269f
C7004 net35 FILLER_0_22_128/a_1828_472# 0.016187f
C7005 net17 _452_/a_2225_156# 0.001943f
C7006 net79 _060_ 0.019511f
C7007 net57 _267_/a_36_472# 0.032037f
C7008 FILLER_0_19_125/a_124_375# vdd 0.032954f
C7009 _170_ vdd 0.18848f
C7010 net82 _386_/a_1084_68# 0.001068f
C7011 FILLER_0_12_2/a_124_375# net67 0.003339f
C7012 result[4] FILLER_0_17_282/a_36_472# 0.017375f
C7013 net68 FILLER_0_6_47/a_484_472# 0.005391f
C7014 _137_ _333_/a_36_160# 0.022811f
C7015 _000_ FILLER_0_3_221/a_1020_375# 0.016709f
C7016 FILLER_0_18_2/a_2812_375# net55 0.007169f
C7017 _098_ _437_/a_36_151# 0.092841f
C7018 FILLER_0_10_214/a_124_375# _069_ 0.014379f
C7019 _119_ _160_ 0.037232f
C7020 output42/a_224_472# net39 0.027208f
C7021 _074_ vdd 1.221102f
C7022 _119_ _326_/a_36_160# 0.003944f
C7023 _428_/a_36_151# net14 0.004485f
C7024 FILLER_0_8_138/a_36_472# _076_ 0.016628f
C7025 FILLER_0_9_60/a_572_375# FILLER_0_9_72/a_36_472# 0.009654f
C7026 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_572_375# 0.007947f
C7027 FILLER_0_16_89/a_1380_472# _451_/a_1353_112# 0.010457f
C7028 _013_ FILLER_0_17_56/a_484_472# 0.002659f
C7029 _448_/a_36_151# net59 0.062656f
C7030 _039_ net6 0.104745f
C7031 FILLER_0_11_101/a_124_375# vdd 0.024363f
C7032 _327_/a_36_472# _130_ 0.001474f
C7033 mask\[5\] FILLER_0_19_155/a_572_375# 0.007026f
C7034 _440_/a_2665_112# trim_mask\[1\] 0.007959f
C7035 _133_ vss 0.18326f
C7036 _076_ vdd 0.806117f
C7037 FILLER_0_18_100/a_36_472# _356_/a_36_472# 0.010679f
C7038 _081_ net22 0.103561f
C7039 net20 _074_ 0.038279f
C7040 _061_ _058_ 0.02828f
C7041 _114_ _171_ 0.203692f
C7042 FILLER_0_15_180/a_572_375# vss 0.010974f
C7043 FILLER_0_15_180/a_36_472# vdd 0.017678f
C7044 FILLER_0_16_107/a_124_375# _040_ 0.008721f
C7045 _189_/a_255_603# net64 0.002455f
C7046 _086_ net22 0.00117f
C7047 _131_ _403_/a_224_472# 0.003274f
C7048 net20 _076_ 0.228128f
C7049 FILLER_0_16_89/a_932_472# _131_ 0.008223f
C7050 _412_/a_1000_472# net58 0.030238f
C7051 FILLER_0_12_136/a_1380_472# _126_ 0.014722f
C7052 trim_mask\[2\] FILLER_0_3_78/a_36_472# 0.005209f
C7053 FILLER_0_10_78/a_36_472# _439_/a_36_151# 0.00271f
C7054 net80 FILLER_0_22_177/a_932_472# 0.002472f
C7055 net73 FILLER_0_18_139/a_36_472# 0.002491f
C7056 _116_ net79 0.081785f
C7057 FILLER_0_18_2/a_2812_375# net17 0.012909f
C7058 net65 net22 0.374917f
C7059 FILLER_0_14_50/a_36_472# vss 0.002954f
C7060 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_124_375# 0.012222f
C7061 _178_ FILLER_0_14_50/a_36_472# 0.001492f
C7062 ctlp[8] net25 0.055914f
C7063 vdd FILLER_0_13_72/a_124_375# -0.004549f
C7064 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_124_375# 0.009654f
C7065 ctln[0] trim[3] 0.216084f
C7066 net68 _440_/a_448_472# 0.02254f
C7067 net75 FILLER_0_8_263/a_124_375# 0.001386f
C7068 _176_ _451_/a_2449_156# 0.038547f
C7069 _086_ _311_/a_2700_473# 0.00176f
C7070 _420_/a_2665_112# _009_ 0.001752f
C7071 FILLER_0_16_89/a_572_375# net36 0.003629f
C7072 net34 FILLER_0_22_177/a_932_472# 0.003953f
C7073 net55 net44 0.018961f
C7074 en_co_clk vdd 0.245319f
C7075 _255_/a_224_552# _375_/a_36_68# 0.00229f
C7076 net23 net13 0.018808f
C7077 _072_ _058_ 0.029688f
C7078 _095_ _451_/a_1353_112# 0.00475f
C7079 net52 _154_ 0.001512f
C7080 _136_ mask\[9\] 0.015204f
C7081 output31/a_224_472# output36/a_224_472# 0.00289f
C7082 _074_ _251_/a_1130_472# 0.00237f
C7083 _074_ net9 0.002862f
C7084 _063_ _445_/a_2665_112# 0.009759f
C7085 _053_ _414_/a_2665_112# 0.032254f
C7086 FILLER_0_9_223/a_484_472# _055_ 0.026026f
C7087 net27 _415_/a_2665_112# 0.030051f
C7088 FILLER_0_17_72/a_1380_472# net36 0.021039f
C7089 output31/a_224_472# net30 0.149277f
C7090 _359_/a_1044_488# net74 0.005311f
C7091 FILLER_0_17_200/a_484_472# net21 0.017997f
C7092 output44/a_224_472# FILLER_0_19_28/a_124_375# 0.005166f
C7093 net52 FILLER_0_3_142/a_124_375# 0.002239f
C7094 _051_ _098_ 0.006332f
C7095 mask\[9\] _438_/a_1000_472# 0.056239f
C7096 FILLER_0_5_164/a_36_472# vss 0.001809f
C7097 FILLER_0_5_164/a_484_472# vdd 0.005235f
C7098 _415_/a_2248_156# FILLER_0_11_282/a_124_375# 0.001221f
C7099 net27 FILLER_0_12_236/a_572_375# 0.083731f
C7100 _251_/a_906_472# _068_ 0.001762f
C7101 fanout67/a_36_160# _220_/a_67_603# 0.005474f
C7102 net39 net40 0.279259f
C7103 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_572_375# 0.001597f
C7104 FILLER_0_9_223/a_36_472# _128_ 0.00702f
C7105 net51 FILLER_0_12_28/a_36_472# 0.005661f
C7106 result[6] net78 0.027123f
C7107 net52 _442_/a_448_472# 0.044149f
C7108 _036_ _160_ 0.034434f
C7109 _257_/a_244_68# _053_ 0.001138f
C7110 net51 net40 0.060626f
C7111 _428_/a_36_151# FILLER_0_11_109/a_36_472# 0.001221f
C7112 FILLER_0_18_177/a_484_472# vdd 0.006177f
C7113 FILLER_0_18_177/a_36_472# vss 0.002187f
C7114 _431_/a_448_472# vss 0.005583f
C7115 output8/a_224_472# FILLER_0_3_221/a_1468_375# 0.032044f
C7116 _427_/a_2248_156# net36 0.004462f
C7117 FILLER_0_15_142/a_572_375# FILLER_0_15_150/a_36_472# 0.086635f
C7118 mask\[0\] FILLER_0_13_228/a_36_472# 0.002986f
C7119 FILLER_0_7_59/a_36_472# fanout67/a_36_160# 0.013068f
C7120 net56 FILLER_0_16_154/a_572_375# 0.002321f
C7121 _450_/a_2225_156# _039_ 0.034731f
C7122 net18 _419_/a_796_472# 0.006586f
C7123 _431_/a_36_151# _142_ 0.030496f
C7124 _439_/a_36_151# FILLER_0_6_47/a_2812_375# 0.001512f
C7125 net16 FILLER_0_18_37/a_932_472# 0.008749f
C7126 output13/a_224_472# ctln[6] 0.080817f
C7127 net44 net17 0.046636f
C7128 _176_ net36 0.336675f
C7129 net48 _265_/a_244_68# 0.00365f
C7130 net69 _441_/a_1000_472# 0.018209f
C7131 FILLER_0_21_142/a_36_472# vss 0.009084f
C7132 FILLER_0_17_104/a_572_375# net14 0.004285f
C7133 _429_/a_448_472# _043_ 0.003615f
C7134 calibrate FILLER_0_9_270/a_36_472# 0.00119f
C7135 _425_/a_796_472# vdd 0.002206f
C7136 FILLER_0_17_282/a_36_472# _418_/a_1308_423# 0.001295f
C7137 _081_ vdd 0.729534f
C7138 mask\[7\] FILLER_0_22_128/a_484_472# 0.010605f
C7139 net17 FILLER_0_20_15/a_1380_472# 0.012286f
C7140 FILLER_0_17_282/a_36_472# _006_ 0.002964f
C7141 _069_ _429_/a_36_151# 0.010076f
C7142 net37 FILLER_0_6_231/a_572_375# 0.001989f
C7143 mask\[8\] net71 0.424276f
C7144 FILLER_0_15_116/a_484_472# FILLER_0_14_107/a_1468_375# 0.001723f
C7145 mask\[7\] _049_ 0.234746f
C7146 net64 FILLER_0_9_270/a_572_375# 0.017924f
C7147 _430_/a_36_151# _337_/a_49_472# 0.023882f
C7148 net53 _427_/a_1000_472# 0.008132f
C7149 _247_/a_36_160# _228_/a_36_68# 0.001919f
C7150 _067_ FILLER_0_12_20/a_572_375# 0.01186f
C7151 _105_ output33/a_224_472# 0.099107f
C7152 _448_/a_1000_472# net22 0.011389f
C7153 _086_ vdd 1.212255f
C7154 _096_ FILLER_0_12_196/a_124_375# 0.002309f
C7155 _050_ _352_/a_49_472# 0.005393f
C7156 _090_ net22 0.032492f
C7157 _428_/a_1308_423# net74 0.0098f
C7158 net20 _081_ 0.024512f
C7159 output7/a_224_472# output40/a_224_472# 0.038066f
C7160 net50 _439_/a_796_472# 0.002389f
C7161 net52 _439_/a_1204_472# 0.027632f
C7162 ctln[3] ctln[4] 0.073214f
C7163 net3 FILLER_0_15_10/a_36_472# 0.002825f
C7164 _137_ mask\[1\] 0.782055f
C7165 FILLER_0_4_49/a_572_375# vdd 0.005972f
C7166 _098_ FILLER_0_16_154/a_1468_375# 0.009042f
C7167 net65 vdd 1.430654f
C7168 fanout54/a_36_160# FILLER_0_19_142/a_36_472# 0.002647f
C7169 _119_ _374_/a_36_68# 0.001756f
C7170 output31/a_224_472# _417_/a_36_151# 0.07368f
C7171 _013_ FILLER_0_18_53/a_484_472# 0.012916f
C7172 _431_/a_1000_472# vss 0.002491f
C7173 _136_ _337_/a_257_69# 0.002933f
C7174 _015_ FILLER_0_8_247/a_484_472# 0.005458f
C7175 net32 net33 0.467071f
C7176 _176_ FILLER_0_10_107/a_572_375# 0.012296f
C7177 net20 net65 0.335083f
C7178 _142_ net53 0.001961f
C7179 FILLER_0_22_86/a_1020_375# vdd 0.008761f
C7180 _132_ FILLER_0_14_107/a_36_472# 0.002187f
C7181 _153_ net14 0.260217f
C7182 _104_ _294_/a_224_472# 0.003008f
C7183 FILLER_0_11_78/a_572_375# _120_ 0.01683f
C7184 net63 FILLER_0_18_177/a_1380_472# 0.070445f
C7185 output42/a_224_472# clkc 0.004924f
C7186 mask\[4\] FILLER_0_19_171/a_124_375# 0.001988f
C7187 fanout77/a_36_113# _094_ 0.002244f
C7188 _095_ FILLER_0_13_80/a_124_375# 0.001989f
C7189 FILLER_0_22_128/a_1828_472# vdd 0.005724f
C7190 FILLER_0_22_128/a_1380_472# vss 0.007305f
C7191 _077_ _042_ 0.045685f
C7192 _140_ _354_/a_49_472# 0.004731f
C7193 _186_ _181_ 0.018817f
C7194 ctln[3] _000_ 0.008418f
C7195 _035_ net38 0.02987f
C7196 _430_/a_2560_156# mask\[2\] 0.010268f
C7197 FILLER_0_4_152/a_36_472# _170_ 0.005476f
C7198 _372_/a_3662_472# net23 0.002864f
C7199 mask\[5\] FILLER_0_19_187/a_36_472# 0.007596f
C7200 ctln[8] FILLER_0_0_96/a_36_472# 0.012298f
C7201 output9/a_224_472# cal 0.011495f
C7202 FILLER_0_16_89/a_36_472# _397_/a_36_472# 0.004546f
C7203 state\[0\] _274_/a_1164_497# 0.002914f
C7204 net56 FILLER_0_18_139/a_36_472# 0.002172f
C7205 net27 FILLER_0_9_290/a_36_472# 0.006729f
C7206 _121_ vss 0.082882f
C7207 FILLER_0_9_28/a_572_375# _054_ 0.002983f
C7208 fanout78/a_36_113# vss 0.031944f
C7209 _174_ _180_ 0.102241f
C7210 net31 net18 0.114197f
C7211 _297_/a_36_472# _108_ 0.011437f
C7212 FILLER_0_24_63/a_36_472# output26/a_224_472# 0.023414f
C7213 output32/a_224_472# _419_/a_36_151# 0.129117f
C7214 net63 FILLER_0_17_218/a_124_375# 0.040329f
C7215 _445_/a_448_472# _034_ 0.03826f
C7216 _053_ FILLER_0_6_47/a_3260_375# 0.002746f
C7217 _119_ _133_ 0.038875f
C7218 _185_ _402_/a_728_93# 0.007151f
C7219 net36 FILLER_0_18_76/a_124_375# 0.001741f
C7220 net82 FILLER_0_3_172/a_36_472# 0.007612f
C7221 _080_ net59 0.038227f
C7222 mask\[5\] ctlp[4] 0.001643f
C7223 _124_ FILLER_0_10_107/a_572_375# 0.002135f
C7224 _430_/a_36_151# net81 0.017255f
C7225 _067_ FILLER_0_12_28/a_124_375# 0.012779f
C7226 _093_ FILLER_0_18_107/a_484_472# 0.008683f
C7227 trim_mask\[2\] _447_/a_448_472# 0.002533f
C7228 trim_val\[2\] _447_/a_36_151# 0.022122f
C7229 net78 _422_/a_36_151# 0.023285f
C7230 FILLER_0_3_172/a_2812_375# net65 0.003745f
C7231 FILLER_0_3_172/a_36_472# fanout57/a_36_113# 0.19419f
C7232 _128_ _176_ 0.180252f
C7233 _391_/a_245_68# cal_count\[0\] 0.001201f
C7234 _446_/a_1000_472# vdd 0.001598f
C7235 _046_ vss 0.088886f
C7236 _155_ vss 0.13648f
C7237 _432_/a_2665_112# vdd 0.009104f
C7238 FILLER_0_4_197/a_484_472# _088_ 0.014756f
C7239 _086_ _135_ 0.005637f
C7240 FILLER_0_15_116/a_484_472# vdd 0.006111f
C7241 _443_/a_448_472# vdd 0.007773f
C7242 net65 net9 0.061456f
C7243 _443_/a_36_151# vss 0.019802f
C7244 FILLER_0_22_86/a_124_375# _437_/a_36_151# 0.001597f
C7245 _120_ _042_ 0.031451f
C7246 _035_ net66 1.624557f
C7247 _414_/a_2248_156# cal_itt\[3\] 0.032294f
C7248 _070_ _055_ 0.516713f
C7249 net28 _196_/a_36_160# 0.060575f
C7250 net68 _232_/a_67_603# 0.00184f
C7251 output48/a_224_472# _425_/a_36_151# 0.004037f
C7252 _439_/a_2665_112# net14 0.004943f
C7253 _448_/a_1000_472# vdd 0.004267f
C7254 _028_ FILLER_0_5_72/a_1380_472# 0.002164f
C7255 _415_/a_2665_112# net18 0.004988f
C7256 net81 net79 0.178225f
C7257 net68 _220_/a_255_603# 0.001908f
C7258 _090_ vdd 0.751973f
C7259 _149_ FILLER_0_20_98/a_36_472# 0.067283f
C7260 _104_ result[9] 0.169685f
C7261 _182_ _179_ 0.109377f
C7262 FILLER_0_16_57/a_572_375# net72 0.012909f
C7263 _425_/a_36_151# FILLER_0_8_247/a_124_375# 0.001597f
C7264 fanout77/a_36_113# net78 0.019286f
C7265 net75 _123_ 0.173358f
C7266 _128_ _124_ 0.111918f
C7267 FILLER_0_5_54/a_1468_375# net47 0.005049f
C7268 FILLER_0_7_59/a_484_472# net68 0.002785f
C7269 fanout70/a_36_113# net70 0.073707f
C7270 _261_/a_36_160# _059_ 0.004993f
C7271 net68 _453_/a_36_151# 0.039234f
C7272 net57 _428_/a_448_472# 0.032029f
C7273 cal_itt\[3\] net37 0.03677f
C7274 net75 _073_ 0.34505f
C7275 output42/a_224_472# net47 0.083794f
C7276 net72 _183_ 0.093818f
C7277 _433_/a_2665_112# _145_ 0.018359f
C7278 FILLER_0_21_142/a_124_375# net35 0.00123f
C7279 FILLER_0_7_72/a_2724_472# net14 0.012436f
C7280 _016_ FILLER_0_12_136/a_124_375# 0.008914f
C7281 _098_ _204_/a_67_603# 0.00539f
C7282 net65 FILLER_0_2_165/a_124_375# 0.001177f
C7283 _255_/a_224_552# _070_ 0.001333f
C7284 _242_/a_36_160# FILLER_0_5_164/a_124_375# 0.005705f
C7285 _069_ _076_ 0.033276f
C7286 _126_ _070_ 0.089475f
C7287 _132_ vss 0.492496f
C7288 FILLER_0_7_195/a_124_375# _414_/a_36_151# 0.059049f
C7289 ctln[6] _442_/a_448_472# 0.003039f
C7290 _386_/a_1152_472# _163_ 0.004076f
C7291 _053_ FILLER_0_8_37/a_36_472# 0.001011f
C7292 _126_ FILLER_0_15_180/a_124_375# 0.001238f
C7293 FILLER_0_17_72/a_2812_375# vdd 0.005986f
C7294 FILLER_0_12_20/a_36_472# net47 0.020589f
C7295 FILLER_0_8_263/a_124_375# net19 0.039576f
C7296 ctln[3] _411_/a_2665_112# 0.003037f
C7297 mask\[0\] _137_ 0.009052f
C7298 FILLER_0_4_107/a_932_472# vdd 0.00987f
C7299 _414_/a_36_151# net22 0.014398f
C7300 trim_mask\[4\] _370_/a_124_24# 0.015021f
C7301 _427_/a_36_151# vss 0.019281f
C7302 net34 _421_/a_2665_112# 0.001056f
C7303 net72 FILLER_0_15_59/a_572_375# 0.00799f
C7304 _029_ vdd 0.223076f
C7305 _043_ FILLER_0_13_72/a_572_375# 0.013294f
C7306 net52 FILLER_0_2_111/a_36_472# 0.0659f
C7307 _370_/a_124_24# net47 0.017609f
C7308 FILLER_0_7_195/a_124_375# _163_ 0.001308f
C7309 net18 net77 0.378783f
C7310 _424_/a_2665_112# FILLER_0_21_60/a_572_375# 0.001077f
C7311 _053_ _160_ 0.0539f
C7312 FILLER_0_7_72/a_2276_472# _053_ 0.016004f
C7313 FILLER_0_8_107/a_124_375# FILLER_0_9_105/a_484_472# 0.001684f
C7314 trim_mask\[2\] FILLER_0_2_93/a_572_375# 0.002818f
C7315 _091_ FILLER_0_15_212/a_1020_375# 0.00799f
C7316 net52 _440_/a_1000_472# 0.013793f
C7317 mask\[3\] FILLER_0_16_241/a_36_472# 0.00209f
C7318 mask\[3\] FILLER_0_18_177/a_1468_375# 0.002924f
C7319 net60 _421_/a_2665_112# 0.044114f
C7320 vdd _145_ 0.082579f
C7321 _321_/a_170_472# vss 0.024882f
C7322 FILLER_0_14_50/a_36_472# _095_ 0.013704f
C7323 fanout74/a_36_113# _032_ 0.012909f
C7324 mask\[4\] _343_/a_49_472# 0.036987f
C7325 FILLER_0_8_107/a_36_472# vdd 0.117254f
C7326 FILLER_0_8_107/a_124_375# vss 0.031335f
C7327 _452_/a_36_151# _041_ 0.013289f
C7328 ctlp[6] ctlp[7] 0.002504f
C7329 net81 _429_/a_2560_156# 0.003888f
C7330 FILLER_0_11_142/a_484_472# _120_ 0.007893f
C7331 _408_/a_56_524# vdd 0.003158f
C7332 _408_/a_728_93# vss 0.001345f
C7333 _163_ net22 0.005017f
C7334 FILLER_0_13_142/a_1380_472# vss 0.004953f
C7335 net49 _440_/a_1000_472# 0.020434f
C7336 _021_ vdd 0.022473f
C7337 net7 _446_/a_2248_156# 0.001166f
C7338 _235_/a_255_603# trim_val\[2\] 0.002471f
C7339 FILLER_0_7_59/a_484_472# net67 0.03109f
C7340 _078_ FILLER_0_4_213/a_572_375# 0.02957f
C7341 _143_ vss 0.02001f
C7342 FILLER_0_9_223/a_484_472# _426_/a_2665_112# 0.004209f
C7343 _447_/a_1000_472# vdd 0.003392f
C7344 _032_ FILLER_0_2_127/a_124_375# 0.002221f
C7345 net58 _411_/a_2248_156# 0.014884f
C7346 net58 net5 0.387314f
C7347 result[9] net29 0.001272f
C7348 net57 FILLER_0_8_156/a_572_375# 0.014948f
C7349 _318_/a_224_472# vdd 0.001873f
C7350 _136_ _067_ 0.051914f
C7351 result[4] vss 0.306116f
C7352 _081_ FILLER_0_5_198/a_572_375# 0.001285f
C7353 FILLER_0_12_2/a_572_375# _039_ 0.005407f
C7354 FILLER_0_11_64/a_36_472# _453_/a_36_151# 0.001723f
C7355 result[2] result[3] 0.09741f
C7356 net23 FILLER_0_22_128/a_1916_375# 0.004205f
C7357 net59 vss 1.191297f
C7358 mask\[4\] _047_ 0.080091f
C7359 _137_ FILLER_0_16_154/a_36_472# 0.005011f
C7360 output29/a_224_472# _193_/a_36_160# 0.006363f
C7361 net47 net40 0.635497f
C7362 _341_/a_257_69# _137_ 0.004351f
C7363 cal_itt\[2\] _074_ 0.082824f
C7364 FILLER_0_0_198/a_124_375# vss 0.017602f
C7365 FILLER_0_0_198/a_36_472# vdd 0.052226f
C7366 _315_/a_36_68# net23 0.030384f
C7367 net75 net81 0.420021f
C7368 ctlp[3] _109_ 0.001371f
C7369 _093_ net23 0.042838f
C7370 _308_/a_692_472# trim_mask\[0\] 0.004377f
C7371 net15 _453_/a_2665_112# 0.011775f
C7372 _002_ _413_/a_36_151# 0.0076f
C7373 fanout60/a_36_160# net62 0.049222f
C7374 FILLER_0_21_125/a_572_375# _433_/a_36_151# 0.059049f
C7375 net68 net69 0.053856f
C7376 net74 _370_/a_124_24# 0.083426f
C7377 _119_ _121_ 0.007336f
C7378 net41 FILLER_0_12_28/a_124_375# 0.003909f
C7379 _016_ _428_/a_36_151# 0.001824f
C7380 vss FILLER_0_10_94/a_484_472# 0.001244f
C7381 _444_/a_796_472# _054_ 0.001838f
C7382 _071_ _121_ 0.007734f
C7383 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_124_375# 0.007947f
C7384 _418_/a_2665_112# _417_/a_2665_112# 0.00131f
C7385 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_36_472# 0.026657f
C7386 _146_ vss 0.078821f
C7387 FILLER_0_18_2/a_2724_472# _452_/a_36_151# 0.011733f
C7388 FILLER_0_18_2/a_1828_472# _452_/a_1353_112# 0.001313f
C7389 FILLER_0_18_2/a_36_472# _452_/a_3129_107# 0.035307f
C7390 net82 FILLER_0_2_177/a_484_472# 0.001777f
C7391 output8/a_224_472# net8 0.034396f
C7392 result[8] FILLER_0_24_290/a_36_472# 0.004676f
C7393 _053_ FILLER_0_7_72/a_932_472# 0.01339f
C7394 FILLER_0_8_24/a_36_472# _054_ 0.007348f
C7395 _449_/a_36_151# FILLER_0_13_72/a_124_375# 0.059049f
C7396 cal_count\[1\] FILLER_0_15_59/a_36_472# 0.00544f
C7397 _180_ FILLER_0_15_59/a_124_375# 0.009926f
C7398 _138_ _043_ 0.005826f
C7399 _412_/a_2248_156# vss 0.005692f
C7400 net65 FILLER_0_2_177/a_572_375# 0.017058f
C7401 _086_ _069_ 0.580351f
C7402 FILLER_0_14_91/a_484_472# _070_ 0.001773f
C7403 _085_ cal_count\[3\] 0.653405f
C7404 net69 _156_ 0.008057f
C7405 _414_/a_36_151# vdd 0.166006f
C7406 _449_/a_1308_423# net55 0.001985f
C7407 _091_ FILLER_0_12_220/a_36_472# 0.003655f
C7408 _004_ net81 0.993594f
C7409 _025_ _436_/a_1204_472# 0.01349f
C7410 _422_/a_448_472# _109_ 0.006344f
C7411 FILLER_0_5_206/a_36_472# net22 0.049294f
C7412 _057_ _250_/a_36_68# 0.014333f
C7413 _122_ vss 0.750387f
C7414 _090_ _279_/a_244_68# 0.001986f
C7415 net33 _434_/a_36_151# 0.002776f
C7416 _035_ net41 0.048883f
C7417 _083_ FILLER_0_3_221/a_572_375# 0.001072f
C7418 _119_ _312_/a_672_472# 0.00145f
C7419 net64 FILLER_0_15_235/a_36_472# 0.046292f
C7420 FILLER_0_16_37/a_36_472# vss 0.005874f
C7421 _444_/a_1000_472# vdd 0.004148f
C7422 _178_ FILLER_0_16_37/a_36_472# 0.007425f
C7423 FILLER_0_7_233/a_36_472# vdd 0.016804f
C7424 FILLER_0_7_233/a_124_375# vss 0.003952f
C7425 net41 FILLER_0_17_38/a_124_375# 0.001109f
C7426 _044_ FILLER_0_13_290/a_36_472# 0.001194f
C7427 cal_count\[3\] _408_/a_1936_472# 0.007046f
C7428 FILLER_0_0_232/a_124_375# vdd 0.012494f
C7429 FILLER_0_10_256/a_36_472# vss 0.001792f
C7430 FILLER_0_8_24/a_36_472# vss 0.001239f
C7431 FILLER_0_8_24/a_484_472# vdd 0.009032f
C7432 FILLER_0_21_142/a_124_375# _433_/a_2665_112# 0.004834f
C7433 net78 _419_/a_36_151# 0.007437f
C7434 _227_/a_36_160# vss 0.010455f
C7435 output33/a_224_472# output18/a_224_472# 0.111946f
C7436 net64 vss 0.636644f
C7437 _453_/a_2665_112# net51 0.046426f
C7438 net11 vdd 0.330644f
C7439 _166_ _160_ 0.492224f
C7440 net35 FILLER_0_23_88/a_36_472# 0.00675f
C7441 _440_/a_2248_156# _164_ 0.054298f
C7442 fanout51/a_36_113# FILLER_0_11_64/a_36_472# 0.001396f
C7443 _070_ state\[1\] 0.032046f
C7444 net38 _452_/a_1353_112# 0.005918f
C7445 _169_ vss 0.037006f
C7446 net20 FILLER_0_7_233/a_36_472# 0.035074f
C7447 _163_ vdd 0.418075f
C7448 FILLER_0_4_49/a_36_472# net68 0.00894f
C7449 output23/a_224_472# FILLER_0_22_128/a_1468_375# 0.00242f
C7450 _010_ _420_/a_2248_156# 0.047408f
C7451 _159_ _370_/a_124_24# 0.021983f
C7452 fanout61/a_36_113# ctlp[1] 0.019606f
C7453 FILLER_0_0_96/a_36_472# net14 0.009584f
C7454 FILLER_0_2_93/a_484_472# vss 0.003689f
C7455 FILLER_0_19_171/a_1380_472# vss 0.004488f
C7456 _430_/a_2665_112# FILLER_0_17_218/a_572_375# 0.002362f
C7457 output21/a_224_472# net21 0.011791f
C7458 mask\[8\] _437_/a_1000_472# 0.00112f
C7459 result[9] net60 0.251903f
C7460 output15/a_224_472# vdd 0.025731f
C7461 FILLER_0_21_28/a_124_375# vdd 0.014155f
C7462 FILLER_0_11_78/a_124_375# vdd -0.011022f
C7463 _413_/a_448_472# net65 0.044062f
C7464 FILLER_0_9_28/a_3260_375# net51 0.001597f
C7465 net23 FILLER_0_5_148/a_484_472# 0.047258f
C7466 net44 _452_/a_2449_156# 0.0059f
C7467 _109_ _108_ 0.001806f
C7468 net5 clk 0.042578f
C7469 FILLER_0_0_96/a_124_375# trim_mask\[3\] 0.006277f
C7470 trim_val\[2\] vss 0.027243f
C7471 FILLER_0_6_239/a_124_375# _123_ 0.044771f
C7472 _327_/a_244_68# _130_ 0.00117f
C7473 net32 net22 0.042885f
C7474 net19 _109_ 0.005991f
C7475 FILLER_0_2_93/a_36_472# _441_/a_2665_112# 0.007491f
C7476 FILLER_0_4_152/a_124_375# _170_ 0.029927f
C7477 _253_/a_1528_68# cal_itt\[1\] 0.002251f
C7478 _131_ FILLER_0_11_124/a_124_375# 0.008946f
C7479 mask\[4\] _291_/a_36_160# 0.00591f
C7480 net15 _168_ 0.04897f
C7481 FILLER_0_21_142/a_124_375# vdd 0.020936f
C7482 _093_ FILLER_0_17_104/a_124_375# 0.01418f
C7483 FILLER_0_23_44/a_36_472# vss 0.002194f
C7484 FILLER_0_23_44/a_484_472# vdd 0.003276f
C7485 FILLER_0_2_165/a_36_472# net59 0.067972f
C7486 _053_ FILLER_0_7_59/a_572_375# 0.014569f
C7487 _305_/a_36_159# _112_ 0.001664f
C7488 mask\[5\] FILLER_0_19_195/a_124_375# 0.007169f
C7489 net15 _441_/a_796_472# 0.021664f
C7490 FILLER_0_5_164/a_36_472# _385_/a_36_68# 0.001674f
C7491 _173_ FILLER_0_12_28/a_36_472# 0.001633f
C7492 FILLER_0_18_209/a_484_472# _201_/a_67_603# 0.001605f
C7493 _408_/a_728_93# _184_ 0.001389f
C7494 FILLER_0_16_89/a_932_472# FILLER_0_17_72/a_2812_375# 0.001723f
C7495 _377_/a_36_472# net68 0.001305f
C7496 _440_/a_2560_156# net47 0.003888f
C7497 net29 _101_ 0.007132f
C7498 _136_ net23 0.031512f
C7499 _418_/a_1308_423# vss 0.001913f
C7500 FILLER_0_14_107/a_1380_472# vss 0.001338f
C7501 cal_itt\[2\] _081_ 0.003204f
C7502 _006_ vss 0.111492f
C7503 _105_ output34/a_224_472# 0.007506f
C7504 FILLER_0_10_28/a_124_375# net51 0.00979f
C7505 _433_/a_1000_472# _022_ 0.05526f
C7506 FILLER_0_4_197/a_1380_472# vss 0.007979f
C7507 FILLER_0_22_177/a_484_472# net33 0.013149f
C7508 FILLER_0_18_2/a_572_375# net38 0.007477f
C7509 _043_ _113_ 0.048005f
C7510 FILLER_0_15_116/a_36_472# _095_ 0.001098f
C7511 net52 FILLER_0_9_72/a_572_375# 0.022582f
C7512 FILLER_0_21_286/a_484_472# vdd 0.007903f
C7513 FILLER_0_21_286/a_36_472# vss 0.004123f
C7514 FILLER_0_13_142/a_124_375# net23 0.003962f
C7515 _103_ vss 0.098913f
C7516 FILLER_0_9_223/a_484_472# _223_/a_36_160# 0.004695f
C7517 FILLER_0_4_99/a_124_375# FILLER_0_4_107/a_36_472# 0.009654f
C7518 output39/a_224_472# vdd 0.022593f
C7519 _057_ _310_/a_49_472# 0.015839f
C7520 FILLER_0_1_266/a_572_375# vdd 0.030477f
C7521 _376_/a_36_160# _164_ 0.004503f
C7522 _069_ _090_ 1.067281f
C7523 _117_ vdd 0.050188f
C7524 FILLER_0_5_206/a_36_472# vdd 0.090007f
C7525 FILLER_0_5_206/a_124_375# vss 0.050652f
C7526 cal_count\[3\] _062_ 0.004405f
C7527 cal_itt\[2\] net65 0.514538f
C7528 _053_ _133_ 0.288819f
C7529 net63 _337_/a_49_472# 0.001801f
C7530 _071_ FILLER_0_13_142/a_1380_472# 0.001617f
C7531 FILLER_0_18_2/a_484_472# vdd 0.003495f
C7532 FILLER_0_18_2/a_36_472# vss 0.001872f
C7533 FILLER_0_17_226/a_124_375# vdd 0.026497f
C7534 _059_ _062_ 0.161331f
C7535 _303_/a_36_472# _012_ 0.001735f
C7536 _402_/a_2172_497# cal_count\[1\] 0.008211f
C7537 FILLER_0_5_109/a_36_472# _163_ 0.00319f
C7538 FILLER_0_18_61/a_36_472# vss 0.00605f
C7539 _428_/a_2248_156# _131_ 0.005621f
C7540 _089_ FILLER_0_3_172/a_2276_472# 0.001522f
C7541 FILLER_0_9_28/a_2812_375# net68 0.012462f
C7542 _093_ FILLER_0_19_134/a_124_375# 0.003473f
C7543 trim[2] trim[3] 0.056575f
C7544 _017_ net14 0.014743f
C7545 mask\[5\] FILLER_0_18_177/a_1828_472# 0.001038f
C7546 net82 FILLER_0_3_221/a_124_375# 0.015932f
C7547 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_36_472# 0.026657f
C7548 vss FILLER_0_4_91/a_572_375# 0.055113f
C7549 output25/a_224_472# mask\[8\] 0.015742f
C7550 _098_ FILLER_0_20_87/a_36_472# 0.016138f
C7551 FILLER_0_17_226/a_124_375# net20 0.001895f
C7552 _074_ FILLER_0_6_231/a_484_472# 0.004409f
C7553 vss _433_/a_3041_156# 0.001287f
C7554 _132_ _095_ 0.042874f
C7555 fanout75/a_36_113# _083_ 0.002133f
C7556 _114_ _131_ 0.036548f
C7557 output32/a_224_472# net60 0.191561f
C7558 _239_/a_36_160# _447_/a_36_151# 0.137659f
C7559 FILLER_0_3_172/a_1380_472# net22 0.012284f
C7560 output21/a_224_472# mask\[7\] 0.032297f
C7561 net73 FILLER_0_17_104/a_1380_472# 0.003206f
C7562 _438_/a_2665_112# FILLER_0_19_111/a_36_472# 0.007491f
C7563 FILLER_0_12_136/a_36_472# _127_ 0.023927f
C7564 _422_/a_1204_472# mask\[7\] 0.025592f
C7565 output16/a_224_472# ctln[9] 0.08624f
C7566 output31/a_224_472# result[4] 0.049147f
C7567 _377_/a_36_472# net67 0.005639f
C7568 _086_ _267_/a_1792_472# 0.002715f
C7569 net75 valid 0.002077f
C7570 net18 output30/a_224_472# 0.08667f
C7571 net57 _315_/a_36_68# 0.0036f
C7572 FILLER_0_11_78/a_484_472# _389_/a_36_148# 0.001043f
C7573 _427_/a_36_151# _095_ 0.029048f
C7574 FILLER_0_16_37/a_36_472# _184_ 0.001522f
C7575 net38 _398_/a_36_113# 0.061273f
C7576 _091_ _139_ 0.05535f
C7577 net75 FILLER_0_8_247/a_36_472# 0.002992f
C7578 net32 vdd 0.50705f
C7579 FILLER_0_17_72/a_2276_472# mask\[9\] 0.006767f
C7580 _430_/a_1308_423# vss 0.003054f
C7581 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_36_472# 0.026657f
C7582 FILLER_0_15_235/a_484_472# mask\[1\] 0.014415f
C7583 result[7] ctlp[1] 0.07619f
C7584 _104_ net78 0.049954f
C7585 _093_ FILLER_0_19_155/a_484_472# 0.001236f
C7586 _066_ _386_/a_124_24# 0.059053f
C7587 result[8] FILLER_0_23_282/a_484_472# 0.001908f
C7588 net74 FILLER_0_13_142/a_572_375# 0.001412f
C7589 FILLER_0_5_198/a_36_472# net59 0.059378f
C7590 ctlp[7] vdd 0.481613f
C7591 FILLER_0_15_142/a_484_472# net23 0.002884f
C7592 _428_/a_36_151# _017_ 0.021229f
C7593 fanout49/a_36_160# _160_ 0.009662f
C7594 _369_/a_692_472# vdd 0.003899f
C7595 net32 net20 0.006161f
C7596 comp vdd 0.108153f
C7597 net29 _094_ 0.313846f
C7598 net36 FILLER_0_15_212/a_1380_472# 0.006416f
C7599 _408_/a_728_93# _095_ 0.040366f
C7600 net81 net19 0.786284f
C7601 net53 net23 0.501857f
C7602 _119_ _122_ 0.155432f
C7603 _095_ FILLER_0_13_142/a_1380_472# 0.001782f
C7604 net2 input5/a_36_113# 0.007518f
C7605 input2/a_36_113# net5 0.001761f
C7606 FILLER_0_7_104/a_36_472# FILLER_0_9_105/a_124_375# 0.001188f
C7607 FILLER_0_2_177/a_36_472# net59 0.007582f
C7608 _176_ _124_ 0.036117f
C7609 FILLER_0_11_142/a_36_472# vdd 0.110248f
C7610 FILLER_0_11_142/a_572_375# vss 0.052505f
C7611 _188_ net51 0.044278f
C7612 _322_/a_692_472# _129_ 0.004891f
C7613 FILLER_0_18_107/a_2812_375# vdd 0.004212f
C7614 net23 _386_/a_124_24# 0.010805f
C7615 output9/a_224_472# net8 0.020421f
C7616 _434_/a_448_472# mask\[6\] 0.060756f
C7617 FILLER_0_20_193/a_36_472# FILLER_0_19_187/a_572_375# 0.001543f
C7618 trim_mask\[4\] _386_/a_848_380# 0.001657f
C7619 _422_/a_2665_112# vss 0.006352f
C7620 _287_/a_36_472# vdd 0.072871f
C7621 FILLER_0_7_104/a_1020_375# vdd 0.010571f
C7622 _119_ _227_/a_36_160# 0.01123f
C7623 FILLER_0_18_139/a_36_472# _145_ 0.002415f
C7624 net79 FILLER_0_12_220/a_932_472# 0.005532f
C7625 output34/a_224_472# _099_ 0.001498f
C7626 net47 _386_/a_848_380# 0.003045f
C7627 _074_ _375_/a_1612_497# 0.004567f
C7628 output29/a_224_472# _416_/a_36_151# 0.07368f
C7629 FILLER_0_7_162/a_36_472# vdd 0.026981f
C7630 FILLER_0_7_162/a_124_375# vss 0.018732f
C7631 _069_ _314_/a_224_472# 0.003461f
C7632 _026_ net71 0.406369f
C7633 net55 FILLER_0_21_60/a_124_375# 0.015315f
C7634 _174_ vss 0.188373f
C7635 FILLER_0_17_72/a_484_472# FILLER_0_18_76/a_36_472# 0.05841f
C7636 _178_ _174_ 0.012157f
C7637 _106_ net63 0.034574f
C7638 _447_/a_796_472# _036_ 0.006511f
C7639 calibrate _055_ 0.006584f
C7640 FILLER_0_23_88/a_124_375# vss 0.014165f
C7641 FILLER_0_23_88/a_36_472# vdd 0.002576f
C7642 _070_ _160_ 0.065914f
C7643 FILLER_0_21_28/a_572_375# FILLER_0_19_28/a_484_472# 0.001512f
C7644 _326_/a_36_160# _070_ 0.018037f
C7645 FILLER_0_12_124/a_36_472# _428_/a_36_151# 0.001723f
C7646 net80 FILLER_0_18_177/a_1828_472# 0.00195f
C7647 _122_ FILLER_0_5_198/a_36_472# 0.00305f
C7648 net47 _452_/a_1040_527# 0.014695f
C7649 output34/a_224_472# _419_/a_2248_156# 0.022045f
C7650 _062_ _226_/a_452_68# 0.001697f
C7651 _131_ FILLER_0_17_104/a_1380_472# 0.004125f
C7652 _091_ FILLER_0_13_212/a_1468_375# 0.003576f
C7653 _072_ _375_/a_692_497# 0.001113f
C7654 _441_/a_36_151# _030_ 0.005324f
C7655 mask\[9\] _149_ 0.040342f
C7656 _097_ vss 0.00839f
C7657 _055_ net21 0.025995f
C7658 net15 _423_/a_2248_156# 0.048449f
C7659 net50 FILLER_0_9_60/a_124_375# 0.001715f
C7660 result[7] FILLER_0_24_274/a_124_375# 0.006125f
C7661 fanout73/a_36_113# _136_ 0.002661f
C7662 net67 FILLER_0_6_37/a_124_375# 0.002918f
C7663 _449_/a_2248_156# _038_ 0.016483f
C7664 FILLER_0_3_172/a_1380_472# vdd 0.043045f
C7665 FILLER_0_15_212/a_1380_472# FILLER_0_15_228/a_36_472# 0.013277f
C7666 FILLER_0_5_54/a_1380_472# _440_/a_36_151# 0.001723f
C7667 FILLER_0_5_198/a_484_472# net21 0.051161f
C7668 FILLER_0_11_109/a_124_375# FILLER_0_10_107/a_484_472# 0.001684f
C7669 FILLER_0_7_104/a_484_472# _058_ 0.006506f
C7670 FILLER_0_16_107/a_572_375# FILLER_0_17_104/a_932_472# 0.001723f
C7671 _411_/a_1000_472# net8 0.007241f
C7672 cal_itt\[0\] _084_ 0.061227f
C7673 _422_/a_2665_112# _107_ 0.005055f
C7674 _052_ FILLER_0_18_37/a_484_472# 0.003861f
C7675 _144_ _352_/a_49_472# 0.00176f
C7676 _077_ _439_/a_1000_472# 0.030609f
C7677 _430_/a_448_472# vss 0.003371f
C7678 _424_/a_36_151# FILLER_0_20_31/a_124_375# 0.012574f
C7679 FILLER_0_3_204/a_124_375# FILLER_0_4_197/a_932_472# 0.001597f
C7680 trimb[0] trimb[2] 0.00878f
C7681 ctlp[0] vss 0.005302f
C7682 _144_ _433_/a_1000_472# 0.029564f
C7683 net50 trim_mask\[0\] 0.002835f
C7684 net45 vss 0.028798f
C7685 FILLER_0_5_181/a_36_472# vss 0.001068f
C7686 net44 output6/a_224_472# 0.078248f
C7687 vdd net6 0.134918f
C7688 output21/a_224_472# _105_ 0.034631f
C7689 _126_ net21 0.024842f
C7690 net57 _136_ 0.168299f
C7691 output31/a_224_472# _006_ 0.090006f
C7692 net73 _137_ 0.047989f
C7693 FILLER_0_22_177/a_932_472# mask\[6\] 0.006573f
C7694 ctlp[1] net79 0.002676f
C7695 mask\[2\] vss 0.536426f
C7696 _132_ _332_/a_36_472# 0.055537f
C7697 net35 FILLER_0_22_177/a_484_472# 0.00632f
C7698 net60 _094_ 0.579872f
C7699 mask\[9\] FILLER_0_18_76/a_36_472# 0.002584f
C7700 _130_ _131_ 0.005955f
C7701 _128_ _246_/a_36_68# 0.01024f
C7702 net57 FILLER_0_13_142/a_124_375# 0.011369f
C7703 _172_ vdd 0.008764f
C7704 output31/a_224_472# _103_ 0.006731f
C7705 net16 _041_ 0.029736f
C7706 _104_ mask\[4\] 0.001621f
C7707 net75 _253_/a_36_68# 0.047906f
C7708 net48 vdd 0.35704f
C7709 net54 FILLER_0_18_139/a_1020_375# 0.003589f
C7710 net2 net19 0.031976f
C7711 FILLER_0_7_72/a_3172_472# trim_mask\[0\] 0.001438f
C7712 mask\[4\] FILLER_0_18_209/a_572_375# 0.032112f
C7713 _053_ _312_/a_672_472# 0.001065f
C7714 FILLER_0_8_247/a_1020_375# vdd -0.002559f
C7715 _114_ FILLER_0_11_101/a_124_375# 0.013348f
C7716 _176_ _267_/a_36_472# 0.001681f
C7717 _085_ _267_/a_224_472# 0.002907f
C7718 _025_ FILLER_0_22_107/a_484_472# 0.00892f
C7719 trim_val\[3\] FILLER_0_2_93/a_124_375# 0.001032f
C7720 _114_ _076_ 0.088609f
C7721 net10 net8 0.003331f
C7722 _155_ _053_ 0.122798f
C7723 net58 result[1] 0.004614f
C7724 net20 net48 0.035427f
C7725 FILLER_0_7_72/a_124_375# net50 0.009304f
C7726 net55 FILLER_0_18_37/a_124_375# 0.005899f
C7727 _131_ _182_ 0.113302f
C7728 _141_ _432_/a_36_151# 0.008193f
C7729 trim_val\[1\] _160_ 0.024279f
C7730 FILLER_0_12_136/a_124_375# cal_count\[3\] 0.005006f
C7731 net76 FILLER_0_5_212/a_124_375# 0.004635f
C7732 _322_/a_848_380# _127_ 0.018892f
C7733 _015_ FILLER_0_10_247/a_36_472# 0.007508f
C7734 _067_ _389_/a_36_148# 0.002789f
C7735 output33/a_224_472# net18 0.110644f
C7736 output37/a_224_472# net59 0.001014f
C7737 net58 _412_/a_1456_156# 0.001045f
C7738 FILLER_0_15_150/a_124_375# net53 0.041074f
C7739 _077_ _410_/a_36_68# 0.020334f
C7740 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_572_375# 0.086635f
C7741 _430_/a_36_151# _019_ 0.019296f
C7742 net34 FILLER_0_22_128/a_3172_472# 0.003953f
C7743 _441_/a_448_472# _164_ 0.016938f
C7744 _064_ net68 0.059889f
C7745 trim_val\[2\] _036_ 0.279133f
C7746 _061_ FILLER_0_8_156/a_484_472# 0.00255f
C7747 _075_ _414_/a_2665_112# 0.050503f
C7748 _379_/a_36_472# trim_mask\[1\] 0.003592f
C7749 _013_ _424_/a_2248_156# 0.001828f
C7750 _420_/a_2665_112# vdd 0.024431f
C7751 _420_/a_2248_156# vss -0.001f
C7752 _095_ FILLER_0_14_107/a_1380_472# 0.011439f
C7753 net34 _050_ 0.004662f
C7754 fanout73/a_36_113# net53 0.047141f
C7755 net4 FILLER_0_12_220/a_1380_472# 0.016375f
C7756 _394_/a_1336_472# FILLER_0_13_72/a_36_472# 0.008136f
C7757 _394_/a_728_93# FILLER_0_13_72/a_572_375# 0.001064f
C7758 FILLER_0_15_205/a_36_472# net22 0.037011f
C7759 _018_ FILLER_0_15_205/a_124_375# 0.002309f
C7760 net44 net3 0.195171f
C7761 output26/a_224_472# FILLER_0_23_44/a_36_472# 0.026108f
C7762 _032_ vss 0.02257f
C7763 mask\[4\] mask\[5\] 0.176881f
C7764 vss FILLER_0_16_115/a_124_375# 0.006358f
C7765 vdd FILLER_0_16_115/a_36_472# 0.093403f
C7766 _002_ FILLER_0_4_197/a_36_472# 0.006574f
C7767 _098_ FILLER_0_15_180/a_572_375# 0.01526f
C7768 cal_count\[1\] _451_/a_3129_107# 0.028519f
C7769 net46 net45 0.038161f
C7770 _069_ _117_ 0.041311f
C7771 trimb[4] FILLER_0_15_2/a_36_472# 0.006046f
C7772 net60 net78 0.030634f
C7773 FILLER_0_21_125/a_36_472# net54 0.016672f
C7774 net52 _443_/a_1204_472# 0.005165f
C7775 _086_ FILLER_0_11_124/a_124_375# 0.016039f
C7776 net20 _420_/a_2665_112# 0.030202f
C7777 _431_/a_1308_423# net36 0.002865f
C7778 mask\[9\] FILLER_0_20_107/a_124_375# 0.004716f
C7779 trim_val\[4\] vss 0.192567f
C7780 vdd _450_/a_2225_156# 0.020301f
C7781 _099_ FILLER_0_15_235/a_484_472# 0.002657f
C7782 FILLER_0_16_57/a_572_375# vdd 0.004039f
C7783 FILLER_0_16_57/a_124_375# vss 0.001678f
C7784 _412_/a_2248_156# output37/a_224_472# 0.001141f
C7785 FILLER_0_16_37/a_36_472# _402_/a_1296_93# 0.001477f
C7786 net35 _436_/a_796_472# 0.002146f
C7787 mask\[8\] _436_/a_1000_472# 0.001091f
C7788 _091_ _429_/a_1308_423# 0.031247f
C7789 ctln[4] FILLER_0_0_232/a_36_472# 0.012298f
C7790 output34/a_224_472# output18/a_224_472# 0.002121f
C7791 net55 FILLER_0_13_80/a_124_375# 0.069951f
C7792 _415_/a_1000_472# result[1] 0.005365f
C7793 _174_ _401_/a_36_68# 0.033989f
C7794 net34 _210_/a_255_603# 0.002153f
C7795 FILLER_0_3_78/a_484_472# _160_ 0.004988f
C7796 net72 _181_ 0.004503f
C7797 _265_/a_916_472# _001_ 0.001719f
C7798 _063_ FILLER_0_6_37/a_36_472# 0.014315f
C7799 valid net19 0.00646f
C7800 _183_ vdd 0.109252f
C7801 _239_/a_36_160# vss 0.001596f
C7802 _410_/a_36_68# _120_ 0.073688f
C7803 FILLER_0_19_195/a_36_472# _434_/a_2248_156# 0.001731f
C7804 FILLER_0_15_212/a_572_375# vss 0.005835f
C7805 FILLER_0_15_212/a_1020_375# vdd -0.00211f
C7806 cal_count\[3\] net14 0.028995f
C7807 net68 _042_ 0.037716f
C7808 net57 net53 0.053565f
C7809 _122_ _385_/a_36_68# 0.003549f
C7810 _093_ _438_/a_1308_423# 0.001057f
C7811 _195_/a_67_603# mask\[2\] 0.003161f
C7812 FILLER_0_20_177/a_484_472# _434_/a_36_151# 0.001723f
C7813 _327_/a_36_472# _126_ 0.011444f
C7814 FILLER_0_16_154/a_932_472# vdd 0.00549f
C7815 FILLER_0_16_154/a_484_472# vss 0.003464f
C7816 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_124_375# 0.003732f
C7817 _445_/a_2248_156# _444_/a_36_151# 0.001081f
C7818 net57 _386_/a_124_24# 0.037058f
C7819 net64 FILLER_0_12_236/a_36_472# 0.052381f
C7820 _119_ FILLER_0_7_162/a_124_375# 0.059009f
C7821 output37/a_224_472# net64 0.110037f
C7822 net27 FILLER_0_9_270/a_36_472# 0.041681f
C7823 trim_mask\[1\] FILLER_0_6_47/a_1020_375# 0.007169f
C7824 _058_ net23 0.075446f
C7825 net20 FILLER_0_15_212/a_1020_375# 0.001629f
C7826 _434_/a_36_151# vdd 0.104871f
C7827 FILLER_0_19_111/a_572_375# vss 0.003337f
C7828 FILLER_0_19_111/a_36_472# vdd 0.034386f
C7829 net38 _190_/a_36_160# 0.062343f
C7830 _064_ net67 0.006691f
C7831 _274_/a_36_68# _060_ 0.02117f
C7832 _419_/a_2665_112# vss 0.004064f
C7833 _419_/a_2560_156# vdd 0.003021f
C7834 _053_ FILLER_0_8_107/a_124_375# 0.002386f
C7835 _074_ _083_ 0.035769f
C7836 FILLER_0_5_117/a_124_375# net47 0.011773f
C7837 FILLER_0_15_59/a_572_375# vdd 0.03104f
C7838 FILLER_0_15_59/a_124_375# vss 0.003806f
C7839 net15 FILLER_0_11_64/a_124_375# 0.047331f
C7840 FILLER_0_18_107/a_1020_375# FILLER_0_19_111/a_572_375# 0.05841f
C7841 FILLER_0_7_72/a_3260_375# net14 0.025344f
C7842 _116_ FILLER_0_12_196/a_36_472# 0.010951f
C7843 _080_ FILLER_0_3_221/a_1020_375# 0.001414f
C7844 _070_ _133_ 0.436976f
C7845 _076_ _083_ 0.006023f
C7846 _068_ _078_ 0.002973f
C7847 net54 FILLER_0_20_107/a_36_472# 0.050184f
C7848 _142_ FILLER_0_17_142/a_484_472# 0.01467f
C7849 FILLER_0_19_195/a_36_472# _202_/a_36_160# 0.002647f
C7850 fanout69/a_36_113# vdd 0.00378f
C7851 net76 FILLER_0_3_172/a_1828_472# 0.051851f
C7852 _414_/a_2248_156# net22 0.062122f
C7853 net56 _137_ 0.0313f
C7854 _413_/a_1308_423# net82 0.003079f
C7855 net67 net42 0.101108f
C7856 FILLER_0_7_146/a_36_472# _133_ 0.009796f
C7857 FILLER_0_7_146/a_124_375# _076_ 0.00688f
C7858 _057_ vss 0.169369f
C7859 net75 _079_ 0.071974f
C7860 state\[1\] net21 0.210202f
C7861 _088_ _260_/a_36_68# 0.003476f
C7862 _077_ _313_/a_67_603# 0.007446f
C7863 _086_ _114_ 1.371271f
C7864 result[9] FILLER_0_24_274/a_484_472# 0.003507f
C7865 _064_ _445_/a_448_472# 0.080931f
C7866 net41 FILLER_0_20_31/a_124_375# 0.049106f
C7867 FILLER_0_13_212/a_484_472# net79 0.00402f
C7868 cal vdd 0.318671f
C7869 _053_ net59 0.145863f
C7870 net62 FILLER_0_13_212/a_932_472# 0.059367f
C7871 FILLER_0_4_91/a_484_472# _156_ 0.009828f
C7872 FILLER_0_21_142/a_36_472# _098_ 0.002964f
C7873 output21/a_224_472# result[8] 0.149245f
C7874 _093_ net36 0.214976f
C7875 net81 output28/a_224_472# 0.01335f
C7876 net4 FILLER_0_3_221/a_932_472# 0.002116f
C7877 mask\[4\] net80 0.034957f
C7878 FILLER_0_16_73/a_484_472# vss 0.007212f
C7879 FILLER_0_13_206/a_124_375# net22 0.024537f
C7880 _031_ FILLER_0_2_101/a_124_375# 0.00179f
C7881 FILLER_0_15_205/a_124_375# vss 0.026372f
C7882 FILLER_0_15_205/a_36_472# vdd 0.010089f
C7883 _161_ _310_/a_49_472# 0.022411f
C7884 _147_ _146_ 0.001164f
C7885 net22 net37 0.03068f
C7886 net63 FILLER_0_15_212/a_36_472# 0.059367f
C7887 _450_/a_36_151# clkc 0.033095f
C7888 _450_/a_1353_112# net6 0.054189f
C7889 output47/a_224_472# _452_/a_3129_107# 0.018181f
C7890 FILLER_0_19_125/a_36_472# vss 0.001056f
C7891 _089_ _079_ 0.126206f
C7892 _003_ _087_ 0.054908f
C7893 _305_/a_36_159# net1 0.013619f
C7894 trim_val\[3\] vss 0.249446f
C7895 _013_ net26 0.174966f
C7896 _088_ net4 0.096522f
C7897 ctlp[9] vdd 0.17413f
C7898 FILLER_0_17_38/a_36_472# FILLER_0_18_37/a_36_472# 0.026657f
C7899 FILLER_0_12_220/a_36_472# vdd 0.027911f
C7900 FILLER_0_12_220/a_1468_375# vss 0.057853f
C7901 _132_ _451_/a_448_472# 0.001197f
C7902 FILLER_0_11_64/a_124_375# net51 0.027848f
C7903 output44/a_224_472# net40 0.006489f
C7904 net50 _447_/a_2248_156# 0.007602f
C7905 mask\[4\] net34 0.001774f
C7906 _426_/a_2665_112# calibrate 0.004837f
C7907 cal_count\[3\] FILLER_0_11_109/a_36_472# 0.00702f
C7908 net63 _434_/a_1308_423# 0.003686f
C7909 FILLER_0_17_72/a_2364_375# _451_/a_448_472# 0.001512f
C7910 net40 _381_/a_36_472# 0.020876f
C7911 net31 net32 0.023293f
C7912 output39/a_224_472# _445_/a_1308_423# 0.010408f
C7913 net39 _445_/a_36_151# 0.006056f
C7914 _174_ _095_ 0.977766f
C7915 FILLER_0_20_193/a_124_375# FILLER_0_19_195/a_36_472# 0.001543f
C7916 trim_val\[4\] FILLER_0_2_165/a_36_472# 0.007765f
C7917 FILLER_0_5_72/a_1468_375# _029_ 0.007876f
C7918 FILLER_0_5_72/a_124_375# trim_mask\[1\] 0.010758f
C7919 FILLER_0_22_177/a_36_472# vss 0.002984f
C7920 FILLER_0_22_177/a_484_472# vdd 0.006974f
C7921 _432_/a_448_472# _098_ 0.032293f
C7922 _112_ _001_ 0.002527f
C7923 _099_ _195_/a_255_603# 0.002146f
C7924 trim_val\[3\] _441_/a_2248_156# 0.027464f
C7925 _313_/a_67_603# _120_ 0.005873f
C7926 _371_/a_36_113# vdd 0.007666f
C7927 FILLER_0_4_144/a_484_472# _081_ 0.001145f
C7928 FILLER_0_4_144/a_36_472# _152_ 0.008211f
C7929 FILLER_0_16_89/a_1020_375# net14 0.029702f
C7930 FILLER_0_21_125/a_572_375# _022_ 0.006025f
C7931 _369_/a_36_68# _156_ 0.001359f
C7932 _426_/a_2248_156# net64 0.01109f
C7933 net75 cal_itt\[1\] 0.704169f
C7934 mask\[2\] FILLER_0_16_154/a_1020_375# 0.020485f
C7935 FILLER_0_4_107/a_36_472# _160_ 0.009073f
C7936 _053_ _122_ 0.368823f
C7937 FILLER_0_4_213/a_36_472# vdd 0.087733f
C7938 FILLER_0_4_213/a_572_375# vss 0.017689f
C7939 trim_val\[0\] _054_ 0.010002f
C7940 _418_/a_448_472# _007_ 0.050316f
C7941 _095_ _097_ 0.030222f
C7942 ctln[2] net5 0.001249f
C7943 fanout79/a_36_160# net79 0.011193f
C7944 FILLER_0_21_142/a_572_375# _433_/a_2248_156# 0.006739f
C7945 FILLER_0_22_86/a_572_375# _098_ 0.001139f
C7946 FILLER_0_17_72/a_1468_375# _131_ 0.006871f
C7947 FILLER_0_9_223/a_36_472# _246_/a_36_68# 0.006596f
C7948 FILLER_0_9_28/a_1468_375# net16 0.005202f
C7949 _345_/a_36_160# _132_ 0.078243f
C7950 _136_ _451_/a_2449_156# 0.004653f
C7951 _367_/a_36_68# vss 0.001589f
C7952 mask\[7\] _436_/a_36_151# 0.030028f
C7953 net80 _435_/a_36_151# 0.035259f
C7954 _449_/a_1000_472# vss 0.029565f
C7955 output8/a_224_472# _073_ 0.043098f
C7956 FILLER_0_21_286/a_484_472# net77 0.02147f
C7957 _053_ _169_ 0.014161f
C7958 net4 cal_itt\[0\] 0.054266f
C7959 _028_ FILLER_0_6_90/a_124_375# 0.012573f
C7960 fanout58/a_36_160# fanout59/a_36_160# 0.001216f
C7961 _059_ FILLER_0_8_156/a_124_375# 0.00593f
C7962 _253_/a_36_68# net19 0.019615f
C7963 output25/a_224_472# _423_/a_2665_112# 0.001396f
C7964 net33 _023_ 0.015172f
C7965 _149_ _437_/a_2248_156# 0.031905f
C7966 _026_ _437_/a_1000_472# 0.042316f
C7967 FILLER_0_17_38/a_124_375# _452_/a_36_151# 0.006111f
C7968 vdd trim[3] 0.147228f
C7969 _372_/a_1602_69# _152_ 0.00262f
C7970 _083_ _081_ 0.03934f
C7971 ctlp[5] _024_ 0.022549f
C7972 mask\[3\] FILLER_0_17_161/a_36_472# 0.13873f
C7973 _451_/a_1040_527# _040_ 0.007154f
C7974 _414_/a_2248_156# vdd 0.00901f
C7975 trim_val\[0\] vss 0.11063f
C7976 ctln[1] net5 0.050549f
C7977 ctln[1] _411_/a_2248_156# 0.013381f
C7978 FILLER_0_14_181/a_124_375# _043_ 0.008393f
C7979 net34 _435_/a_36_151# 0.011954f
C7980 _123_ FILLER_0_6_231/a_572_375# 0.00487f
C7981 _402_/a_718_527# vdd 0.020893f
C7982 net15 FILLER_0_6_47/a_1468_375# 0.007439f
C7983 _002_ vss 0.08396f
C7984 net50 _444_/a_2248_156# 0.005539f
C7985 _114_ _090_ 0.001909f
C7986 ctlp[4] mask\[6\] 0.003054f
C7987 net47 _450_/a_36_151# 0.029201f
C7988 _126_ _171_ 0.01633f
C7989 _016_ FILLER_0_12_124/a_36_472# 0.002661f
C7990 _430_/a_36_151# _092_ 0.002363f
C7991 _128_ _315_/a_36_68# 0.04902f
C7992 _413_/a_3041_156# net59 0.001022f
C7993 fanout62/a_36_160# FILLER_0_11_282/a_124_375# 0.058702f
C7994 _196_/a_36_160# FILLER_0_14_263/a_36_472# 0.004828f
C7995 FILLER_0_4_197/a_124_375# net59 0.001026f
C7996 mask\[4\] _276_/a_36_160# 0.025336f
C7997 FILLER_0_19_155/a_124_375# vdd 0.019233f
C7998 FILLER_0_13_206/a_124_375# vdd 0.034528f
C7999 sample vdd 0.154389f
C8000 FILLER_0_18_2/a_1468_375# trimb[1] 0.002041f
C8001 _137_ FILLER_0_15_180/a_36_472# 0.004437f
C8002 _131_ _040_ 0.211618f
C8003 FILLER_0_5_117/a_124_375# _154_ 0.005866f
C8004 net63 FILLER_0_22_177/a_1380_472# 0.062289f
C8005 net41 FILLER_0_19_28/a_572_375# 0.040551f
C8006 net37 vdd 0.544653f
C8007 output24/a_224_472# _436_/a_1308_423# 0.005632f
C8008 _091_ FILLER_0_20_169/a_36_472# 0.007537f
C8009 _136_ net36 1.151311f
C8010 _431_/a_2560_156# vss 0.004767f
C8011 _445_/a_2665_112# vdd 0.055628f
C8012 FILLER_0_21_28/a_2724_472# vss -0.001553f
C8013 _436_/a_796_472# vdd 0.005009f
C8014 FILLER_0_3_221/a_1020_375# vss 0.003948f
C8015 FILLER_0_3_221/a_1468_375# vdd 0.008815f
C8016 _423_/a_2248_156# _012_ 0.011646f
C8017 FILLER_0_17_200/a_124_375# _430_/a_36_151# 0.059049f
C8018 net62 net36 0.034265f
C8019 cal_itt\[3\] _116_ 0.001364f
C8020 _403_/a_224_472# _183_ 0.007508f
C8021 net36 _438_/a_1000_472# 0.072117f
C8022 _126_ mask\[0\] 0.067513f
C8023 ctln[8] net52 0.005231f
C8024 net15 net50 0.177988f
C8025 FILLER_0_16_107/a_484_472# _136_ 0.013449f
C8026 _428_/a_2665_112# _427_/a_36_151# 0.028591f
C8027 _439_/a_1308_423# vss 0.009355f
C8028 net20 net37 0.039674f
C8029 net39 _063_ 0.004732f
C8030 FILLER_0_21_142/a_124_375# _140_ 0.016087f
C8031 _105_ _204_/a_67_603# 0.061486f
C8032 net20 FILLER_0_3_221/a_1468_375# 0.007234f
C8033 _427_/a_2560_156# net23 0.042069f
C8034 _086_ _130_ 0.008816f
C8035 FILLER_0_21_28/a_3260_375# _424_/a_36_151# 0.035849f
C8036 output47/a_224_472# vss 0.002843f
C8037 FILLER_0_8_24/a_572_375# FILLER_0_8_37/a_36_472# 0.007947f
C8038 net57 _058_ 0.028536f
C8039 _070_ _121_ 0.285424f
C8040 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_124_375# 0.007947f
C8041 _115_ _127_ 0.042389f
C8042 FILLER_0_14_99/a_124_375# vdd 0.040312f
C8043 _144_ _149_ 0.032178f
C8044 net62 _193_/a_36_160# 0.00227f
C8045 _132_ _098_ 0.038463f
C8046 _002_ FILLER_0_3_172/a_3260_375# 0.001683f
C8047 FILLER_0_9_28/a_932_472# net68 0.003603f
C8048 _431_/a_36_151# net36 0.006618f
C8049 net50 FILLER_0_6_90/a_572_375# 0.010099f
C8050 _077_ FILLER_0_9_72/a_124_375# 0.008103f
C8051 _056_ _310_/a_49_472# 0.003286f
C8052 FILLER_0_12_2/a_124_375# vss 0.002871f
C8053 FILLER_0_12_2/a_572_375# vdd 0.022401f
C8054 ctln[7] _442_/a_2560_156# 0.001742f
C8055 FILLER_0_10_247/a_124_375# net79 0.00498f
C8056 FILLER_0_16_57/a_932_472# _176_ 0.010635f
C8057 net53 _451_/a_2449_156# 0.015332f
C8058 fanout74/a_36_113# net69 0.006779f
C8059 _057_ _071_ 0.139904f
C8060 _091_ FILLER_0_17_218/a_124_375# 0.013726f
C8061 _077_ _061_ 0.031458f
C8062 ctlp[1] net19 0.029153f
C8063 FILLER_0_8_127/a_36_472# vdd 0.069117f
C8064 _077_ _453_/a_1308_423# 0.071515f
C8065 _077_ _311_/a_66_473# 0.002605f
C8066 _175_ _451_/a_3129_107# 0.021546f
C8067 _408_/a_728_93# cal_count\[0\] 0.007633f
C8068 _208_/a_36_160# vss 0.012188f
C8069 _139_ vdd 0.085044f
C8070 net62 FILLER_0_15_228/a_36_472# 0.002128f
C8071 net55 _216_/a_255_603# 0.001011f
C8072 _370_/a_1152_472# _152_ 0.001423f
C8073 trimb[1] FILLER_0_20_15/a_36_472# 0.001292f
C8074 cal_count\[3\] FILLER_0_12_20/a_124_375# 0.008038f
C8075 FILLER_0_4_123/a_124_375# FILLER_0_4_107/a_1468_375# 0.012001f
C8076 net69 FILLER_0_3_78/a_572_375# 0.002984f
C8077 net60 _418_/a_2248_156# 0.045472f
C8078 net69 FILLER_0_2_127/a_124_375# 0.08337f
C8079 result[2] _044_ 0.393081f
C8080 fanout58/a_36_160# net5 0.003758f
C8081 FILLER_0_4_197/a_1020_375# net76 0.006026f
C8082 trimb[2] vdd 0.084666f
C8083 fanout74/a_36_113# _152_ 0.017267f
C8084 FILLER_0_4_49/a_124_375# trim_val\[1\] 0.024557f
C8085 _004_ fanout79/a_36_160# 0.048599f
C8086 net73 _334_/a_36_160# 0.003275f
C8087 FILLER_0_15_142/a_484_472# net36 0.012033f
C8088 _065_ net68 0.194392f
C8089 trim_val\[2\] _166_ 0.014514f
C8090 trim_mask\[2\] _160_ 0.367302f
C8091 _127_ _395_/a_36_488# 0.00519f
C8092 FILLER_0_7_195/a_36_472# _161_ 0.015074f
C8093 _274_/a_36_68# net81 0.014689f
C8094 _144_ FILLER_0_21_125/a_572_375# 0.003787f
C8095 net62 _417_/a_2248_156# 0.005537f
C8096 _009_ _109_ 0.006736f
C8097 net53 net36 3.423337f
C8098 _412_/a_448_472# net1 0.035155f
C8099 _077_ _072_ 0.178678f
C8100 output34/a_224_472# net18 0.126175f
C8101 _328_/a_36_113# FILLER_0_11_101/a_484_472# 0.001826f
C8102 FILLER_0_9_282/a_124_375# vss 0.00451f
C8103 FILLER_0_9_282/a_572_375# vdd 0.002928f
C8104 FILLER_0_6_47/a_932_472# vdd 0.003435f
C8105 net15 FILLER_0_15_72/a_484_472# 0.002925f
C8106 _093_ FILLER_0_18_177/a_2724_472# 0.003036f
C8107 mask\[8\] FILLER_0_22_107/a_36_472# 0.017159f
C8108 net35 FILLER_0_22_107/a_572_375# 0.010438f
C8109 fanout59/a_36_160# net18 0.003981f
C8110 FILLER_0_2_101/a_124_375# _157_ 0.002818f
C8111 _053_ FILLER_0_7_104/a_572_375# 0.005239f
C8112 _057_ _095_ 0.001346f
C8113 _430_/a_796_472# net36 0.00117f
C8114 net32 _421_/a_448_472# 0.022214f
C8115 _402_/a_728_93# _179_ 0.011717f
C8116 FILLER_0_8_138/a_124_375# _059_ 0.007966f
C8117 _322_/a_848_380# _118_ 0.047787f
C8118 net33 _297_/a_36_472# 0.00521f
C8119 _053_ FILLER_0_7_162/a_124_375# 0.007494f
C8120 FILLER_0_13_212/a_1468_375# vdd -0.013698f
C8121 FILLER_0_13_212/a_1020_375# vss 0.041631f
C8122 _093_ FILLER_0_17_218/a_484_472# 0.004665f
C8123 FILLER_0_9_28/a_1916_375# net16 0.001431f
C8124 net72 _423_/a_36_151# 0.024965f
C8125 net63 _019_ 0.004471f
C8126 ctlp[1] _420_/a_36_151# 0.067975f
C8127 _413_/a_1308_423# net21 0.065716f
C8128 _098_ _146_ 0.004276f
C8129 FILLER_0_11_101/a_484_472# _120_ 0.011393f
C8130 _421_/a_2248_156# vdd 0.035239f
C8131 FILLER_0_20_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001543f
C8132 FILLER_0_10_214/a_36_472# vss 0.008006f
C8133 net19 cal_itt\[1\] 0.044717f
C8134 net20 FILLER_0_13_212/a_1468_375# 0.009573f
C8135 net35 _023_ 0.008361f
C8136 fanout50/a_36_160# net52 0.037383f
C8137 FILLER_0_8_107/a_124_375# _070_ 0.003069f
C8138 FILLER_0_19_187/a_572_375# vdd 0.023383f
C8139 vdd FILLER_0_21_60/a_484_472# 0.005181f
C8140 vss FILLER_0_21_60/a_36_472# 0.001384f
C8141 net26 FILLER_0_23_44/a_932_472# 0.001889f
C8142 net73 FILLER_0_18_107/a_1468_375# 0.024898f
C8143 mask\[0\] state\[1\] 0.064758f
C8144 _305_/a_36_159# net76 0.010842f
C8145 _096_ _320_/a_1792_472# 0.001419f
C8146 FILLER_0_13_65/a_36_472# _174_ 0.011724f
C8147 net56 fanout56/a_36_113# 0.015924f
C8148 FILLER_0_2_111/a_1020_375# vdd 0.007918f
C8149 trimb[2] output17/a_224_472# 0.008375f
C8150 _429_/a_1308_423# net22 0.001856f
C8151 _429_/a_448_472# _018_ 0.035489f
C8152 fanout82/a_36_113# vss 0.023533f
C8153 FILLER_0_4_91/a_124_375# _160_ 0.009765f
C8154 _173_ _186_ 0.002111f
C8155 net15 _394_/a_1336_472# 0.01144f
C8156 fanout50/a_36_160# net49 0.030626f
C8157 FILLER_0_11_109/a_124_375# _134_ 0.027704f
C8158 _445_/a_36_151# net47 0.002364f
C8159 _144_ mask\[5\] 0.38642f
C8160 _091_ _060_ 0.085764f
C8161 _440_/a_1308_423# vdd 0.00218f
C8162 _440_/a_448_472# vss 0.032037f
C8163 FILLER_0_12_124/a_36_472# _017_ 0.004641f
C8164 net18 _418_/a_36_151# 0.017941f
C8165 net64 _098_ 0.281888f
C8166 _016_ cal_count\[3\] 0.004588f
C8167 _077_ FILLER_0_9_60/a_572_375# 0.018665f
C8168 trim[4] net6 0.002404f
C8169 ctln[3] vss 0.133697f
C8170 _390_/a_36_68# vdd 0.012472f
C8171 net82 _443_/a_36_151# 0.03565f
C8172 _004_ FILLER_0_10_247/a_124_375# 0.004573f
C8173 FILLER_0_21_286/a_124_375# net18 0.015582f
C8174 net70 FILLER_0_14_107/a_572_375# 0.018214f
C8175 FILLER_0_5_72/a_1380_472# vss 0.004538f
C8176 _115_ trim_mask\[0\] 0.008966f
C8177 FILLER_0_20_2/a_572_375# vdd 0.010844f
C8178 FILLER_0_20_2/a_124_375# vss 0.002737f
C8179 _087_ net76 0.529571f
C8180 FILLER_0_12_136/a_1380_472# FILLER_0_11_142/a_572_375# 0.001543f
C8181 mask\[4\] _293_/a_36_472# 0.023203f
C8182 _098_ FILLER_0_19_171/a_1380_472# 0.001764f
C8183 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_124_375# 0.004426f
C8184 FILLER_0_5_54/a_36_472# trim_mask\[1\] 0.101342f
C8185 FILLER_0_5_54/a_1380_472# _029_ 0.01027f
C8186 _430_/a_36_151# FILLER_0_18_177/a_2276_472# 0.001793f
C8187 ctlp[1] _419_/a_448_472# 0.020153f
C8188 FILLER_0_7_72/a_3172_472# FILLER_0_7_104/a_36_472# 0.013276f
C8189 trimb[1] cal_count\[2\] 0.003178f
C8190 mask\[5\] net23 0.002188f
C8191 _446_/a_2560_156# net40 0.012204f
C8192 _412_/a_1000_472# net65 0.00929f
C8193 mask\[8\] _433_/a_36_151# 0.001402f
C8194 _448_/a_448_472# net65 0.001006f
C8195 _426_/a_36_151# FILLER_0_8_247/a_1380_472# 0.001723f
C8196 _070_ FILLER_0_10_94/a_484_472# 0.003573f
C8197 _304_/a_224_472# _013_ 0.002769f
C8198 _272_/a_36_472# _003_ 0.001634f
C8199 FILLER_0_5_198/a_572_375# net37 0.009149f
C8200 vss _034_ 0.008249f
C8201 _161_ vss 0.134214f
C8202 fanout60/a_36_160# net60 0.019034f
C8203 en net4 0.125535f
C8204 _421_/a_2560_156# net19 0.006572f
C8205 FILLER_0_12_2/a_484_472# _450_/a_36_151# 0.059367f
C8206 fanout64/a_36_160# net64 0.043709f
C8207 _114_ _117_ 0.008886f
C8208 FILLER_0_13_206/a_36_472# _043_ 0.011439f
C8209 net63 FILLER_0_19_187/a_484_472# 0.020823f
C8210 _442_/a_2248_156# _157_ 0.002731f
C8211 _033_ FILLER_0_6_37/a_124_375# 0.018812f
C8212 _164_ FILLER_0_6_47/a_572_375# 0.010099f
C8213 FILLER_0_18_2/a_1020_375# output44/a_224_472# 0.032639f
C8214 _129_ vss 0.141494f
C8215 FILLER_0_16_89/a_36_472# _177_ 0.048163f
C8216 mask\[4\] FILLER_0_18_177/a_1468_375# 0.01587f
C8217 _069_ FILLER_0_13_206/a_124_375# 0.009695f
C8218 _133_ calibrate 0.0188f
C8219 _070_ _122_ 0.153373f
C8220 net51 _039_ 0.398642f
C8221 FILLER_0_16_255/a_36_472# _287_/a_36_472# 0.004546f
C8222 net5 net18 0.015361f
C8223 _447_/a_36_151# net69 0.001216f
C8224 net49 FILLER_0_3_54/a_36_472# 0.00186f
C8225 _070_ FILLER_0_7_233/a_124_375# 0.004917f
C8226 output9/a_224_472# FILLER_0_1_266/a_484_472# 0.0323f
C8227 _128_ net4 0.039671f
C8228 net1 input4/a_36_68# 0.056389f
C8229 _408_/a_728_93# net17 0.005494f
C8230 net52 net14 0.072003f
C8231 output9/a_224_472# net81 0.02825f
C8232 _059_ FILLER_0_5_148/a_36_472# 0.010977f
C8233 FILLER_0_16_107/a_572_375# vss 0.055104f
C8234 _070_ _227_/a_36_160# 0.00254f
C8235 FILLER_0_17_226/a_36_472# vdd 0.087587f
C8236 _072_ state\[2\] 0.002629f
C8237 _052_ FILLER_0_21_28/a_1916_375# 0.002388f
C8238 _086_ _395_/a_1492_488# 0.001769f
C8239 _070_ _169_ 0.006335f
C8240 FILLER_0_18_37/a_1468_375# vdd 0.021186f
C8241 FILLER_0_16_107/a_36_472# vdd 0.110244f
C8242 _028_ FILLER_0_7_72/a_1916_375# 0.003862f
C8243 _317_/a_36_113# calibrate 0.011799f
C8244 net27 _415_/a_1204_472# 0.006198f
C8245 _096_ _043_ 0.842762f
C8246 _429_/a_448_472# vss 0.035246f
C8247 net49 net14 0.00344f
C8248 net52 _164_ 0.313379f
C8249 _093_ FILLER_0_16_89/a_572_375# 0.002889f
C8250 FILLER_0_12_220/a_1468_375# FILLER_0_12_236/a_36_472# 0.086742f
C8251 _063_ net47 0.142088f
C8252 FILLER_0_10_78/a_1020_375# vss 0.002352f
C8253 FILLER_0_14_99/a_36_472# _043_ 0.001242f
C8254 _307_/a_234_472# _126_ 0.00204f
C8255 net8 vdd 0.593788f
C8256 output47/a_224_472# _095_ 0.012266f
C8257 vss result[3] 0.28152f
C8258 net62 _416_/a_36_151# 0.054002f
C8259 _037_ net22 0.079675f
C8260 net49 _164_ 0.428468f
C8261 FILLER_0_16_57/a_932_472# FILLER_0_17_64/a_124_375# 0.001723f
C8262 net20 _429_/a_1308_423# 0.001186f
C8263 _021_ _137_ 0.002807f
C8264 _093_ FILLER_0_17_72/a_1380_472# 0.008517f
C8265 _144_ net34 0.029247f
C8266 FILLER_0_3_2/a_124_375# net66 0.027628f
C8267 FILLER_0_10_78/a_124_375# vss 0.006775f
C8268 net16 FILLER_0_12_28/a_124_375# 0.002225f
C8269 net1 _001_ 0.300335f
C8270 _394_/a_1936_472# vss 0.006085f
C8271 _238_/a_67_603# _441_/a_2665_112# 0.015187f
C8272 _082_ net59 0.004251f
C8273 _360_/a_36_160# _160_ 0.052885f
C8274 net82 net59 0.102279f
C8275 trim_mask\[1\] FILLER_0_6_79/a_36_472# 0.006265f
C8276 _122_ FILLER_0_5_164/a_572_375# 0.001352f
C8277 _310_/a_49_472# _113_ 0.020387f
C8278 _176_ _315_/a_36_68# 0.003811f
C8279 vss FILLER_0_22_107/a_124_375# 0.002881f
C8280 vdd FILLER_0_22_107/a_572_375# 0.005745f
C8281 _423_/a_36_151# FILLER_0_23_60/a_124_375# 0.005577f
C8282 _181_ vdd 0.209604f
C8283 FILLER_0_20_169/a_124_375# FILLER_0_19_171/a_36_472# 0.001543f
C8284 _132_ FILLER_0_15_116/a_572_375# 0.003964f
C8285 fanout57/a_36_113# net59 0.00178f
C8286 net50 net47 0.040157f
C8287 _035_ net16 0.034977f
C8288 FILLER_0_10_37/a_124_375# net68 0.012617f
C8289 FILLER_0_19_125/a_124_375# _334_/a_36_160# 0.001633f
C8290 net72 FILLER_0_21_28/a_1020_375# 0.040811f
C8291 net15 net72 0.157843f
C8292 net47 _382_/a_224_472# 0.001795f
C8293 net34 net23 0.058486f
C8294 net16 FILLER_0_17_38/a_124_375# 0.046435f
C8295 _320_/a_36_472# net79 0.029189f
C8296 FILLER_0_5_164/a_124_375# _163_ 0.048663f
C8297 _068_ _311_/a_3220_473# 0.004371f
C8298 FILLER_0_2_93/a_124_375# net69 0.015032f
C8299 net15 FILLER_0_5_54/a_484_472# 0.002186f
C8300 _141_ _339_/a_36_160# 0.011118f
C8301 _425_/a_448_472# _122_ 0.002863f
C8302 _425_/a_1308_423# calibrate 0.022697f
C8303 FILLER_0_8_24/a_36_472# net17 0.045619f
C8304 _140_ _434_/a_36_151# 0.025956f
C8305 _424_/a_1204_472# _012_ 0.003572f
C8306 _008_ _102_ 0.027578f
C8307 net62 FILLER_0_14_235/a_484_472# 0.017862f
C8308 _033_ _444_/a_1204_472# 0.002294f
C8309 _023_ vdd 0.062542f
C8310 FILLER_0_12_136/a_1468_375# net23 0.021046f
C8311 net63 _092_ 0.008819f
C8312 cal_itt\[2\] FILLER_0_3_221/a_1468_375# 0.016021f
C8313 _174_ cal_count\[0\] 0.009645f
C8314 net80 _434_/a_796_472# 0.039593f
C8315 _024_ _435_/a_36_151# 0.10993f
C8316 _417_/a_1308_423# vss 0.002064f
C8317 net9 net8 0.027272f
C8318 _232_/a_67_603# vss 0.00988f
C8319 _306_/a_36_68# _116_ 0.00183f
C8320 FILLER_0_20_98/a_124_375# vdd 0.0135f
C8321 FILLER_0_10_214/a_124_375# _055_ 0.001419f
C8322 _091_ _337_/a_49_472# 0.014992f
C8323 FILLER_0_16_107/a_124_375# _132_ 0.003315f
C8324 FILLER_0_4_123/a_36_472# vss 0.004542f
C8325 net82 _122_ 0.001375f
C8326 _127_ vdd 0.155954f
C8327 FILLER_0_19_55/a_36_472# _013_ 0.005889f
C8328 ctln[5] ctln[6] 0.017291f
C8329 FILLER_0_5_72/a_572_375# net47 0.006974f
C8330 _385_/a_244_472# net37 0.001593f
C8331 _056_ vss 0.193804f
C8332 net35 FILLER_0_22_86/a_36_472# 0.00797f
C8333 mask\[8\] FILLER_0_22_86/a_484_472# 0.012439f
C8334 output9/a_224_472# net2 0.003405f
C8335 _412_/a_448_472# net76 0.026446f
C8336 FILLER_0_5_212/a_124_375# _078_ 0.002018f
C8337 FILLER_0_7_59/a_484_472# vss 0.005804f
C8338 _453_/a_36_151# vss 0.007105f
C8339 _453_/a_448_472# vdd 0.010005f
C8340 FILLER_0_13_212/a_36_472# _043_ 0.011752f
C8341 FILLER_0_17_200/a_124_375# net63 0.008905f
C8342 _247_/a_36_160# _062_ 0.011327f
C8343 net35 FILLER_0_22_128/a_2724_472# 0.012359f
C8344 _015_ _426_/a_36_151# 0.01243f
C8345 trim_val\[2\] net17 0.019133f
C8346 _017_ cal_count\[3\] 0.003939f
C8347 net57 _267_/a_672_472# 0.004637f
C8348 FILLER_0_16_89/a_572_375# _136_ 0.069752f
C8349 ctln[1] FILLER_0_3_221/a_124_375# 0.001391f
C8350 _037_ vdd 0.158731f
C8351 FILLER_0_12_2/a_36_472# net67 0.013281f
C8352 _397_/a_36_472# vdd 0.094023f
C8353 net68 FILLER_0_6_47/a_1380_472# 0.049638f
C8354 FILLER_0_11_135/a_36_472# vdd 0.091206f
C8355 FILLER_0_11_135/a_124_375# vss 0.02843f
C8356 _308_/a_1084_68# trim_mask\[0\] 0.001592f
C8357 ctln[2] FILLER_0_0_266/a_124_375# 0.041898f
C8358 net17 FILLER_0_23_44/a_36_472# 0.071244f
C8359 mask\[8\] _050_ 0.001479f
C8360 _098_ _097_ 0.034041f
C8361 _064_ _033_ 0.001986f
C8362 _098_ _437_/a_1308_423# 0.005568f
C8363 _053_ FILLER_0_9_28/a_2364_375# 0.029866f
C8364 net60 _419_/a_3041_156# 0.001022f
C8365 net55 FILLER_0_18_61/a_36_472# 0.022296f
C8366 _115_ _118_ 1.045555f
C8367 FILLER_0_7_72/a_36_472# FILLER_0_7_59/a_484_472# 0.001963f
C8368 FILLER_0_9_60/a_484_472# FILLER_0_9_72/a_36_472# 0.002296f
C8369 FILLER_0_16_89/a_36_472# _451_/a_2225_156# 0.001329f
C8370 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_124_375# 0.012001f
C8371 _448_/a_1308_423# net59 0.014899f
C8372 _039_ clkc 0.003104f
C8373 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_124_375# 0.001597f
C8374 _093_ FILLER_0_18_76/a_124_375# 0.061549f
C8375 FILLER_0_11_101/a_36_472# vdd 0.093852f
C8376 FILLER_0_11_101/a_572_375# vss 0.055325f
C8377 _053_ FILLER_0_4_213/a_572_375# 0.003451f
C8378 _150_ _438_/a_36_151# 0.032532f
C8379 mask\[5\] FILLER_0_19_155/a_484_472# 0.043011f
C8380 _068_ vss 0.547532f
C8381 FILLER_0_18_107/a_36_472# FILLER_0_17_104/a_484_472# 0.026657f
C8382 _114_ _172_ 0.045798f
C8383 FILLER_0_13_212/a_1020_375# FILLER_0_12_220/a_124_375# 0.05841f
C8384 _033_ net42 0.002707f
C8385 _119_ _129_ 0.055585f
C8386 _052_ _424_/a_448_472# 0.017551f
C8387 FILLER_0_15_180/a_484_472# vss 0.001207f
C8388 mask\[1\] FILLER_0_15_180/a_572_375# 0.011186f
C8389 FILLER_0_4_99/a_36_472# _160_ 0.006222f
C8390 mask\[8\] _214_/a_36_160# 0.001264f
C8391 ctln[1] FILLER_0_0_266/a_124_375# 0.01186f
C8392 FILLER_0_1_98/a_124_375# _442_/a_2665_112# 0.003045f
C8393 _395_/a_36_488# _116_ 0.033784f
C8394 FILLER_0_12_124/a_36_472# cal_count\[3\] 0.004109f
C8395 FILLER_0_4_107/a_124_375# _157_ 0.001427f
C8396 _415_/a_1204_472# net18 0.001828f
C8397 _176_ _136_ 0.114837f
C8398 _091_ net81 0.03653f
C8399 net32 output33/a_224_472# 0.018183f
C8400 _018_ _138_ 0.008093f
C8401 _098_ mask\[2\] 0.06158f
C8402 FILLER_0_4_197/a_1380_472# net82 0.003084f
C8403 FILLER_0_9_28/a_3260_375# FILLER_0_9_60/a_36_472# 0.086742f
C8404 _053_ trim_val\[0\] 0.446477f
C8405 vdd FILLER_0_13_72/a_36_472# 0.108152f
C8406 vss FILLER_0_13_72/a_572_375# 0.061657f
C8407 fanout51/a_36_113# vss 0.0844f
C8408 net27 result[1] 0.187252f
C8409 net68 _440_/a_796_472# 0.021463f
C8410 _274_/a_36_68# FILLER_0_12_220/a_932_472# 0.001237f
C8411 _127_ _135_ 0.00622f
C8412 cal_itt\[3\] net47 0.00247f
C8413 _028_ _439_/a_1000_472# 0.003267f
C8414 FILLER_0_19_142/a_36_472# _145_ 0.010377f
C8415 FILLER_0_20_169/a_36_472# vdd 0.010522f
C8416 FILLER_0_20_169/a_124_375# vss 0.017635f
C8417 _345_/a_36_160# FILLER_0_19_111/a_572_375# 0.132282f
C8418 _413_/a_36_151# FILLER_0_3_172/a_1828_472# 0.001723f
C8419 FILLER_0_9_223/a_36_472# net4 0.014911f
C8420 _025_ _437_/a_2665_112# 0.001245f
C8421 _255_/a_224_552# _162_ 0.010564f
C8422 _057_ _375_/a_36_68# 0.003063f
C8423 _188_ _453_/a_796_472# 0.00103f
C8424 _106_ _091_ 0.001188f
C8425 output10/a_224_472# rstn 0.001656f
C8426 _443_/a_2248_156# _386_/a_124_24# 0.001257f
C8427 _414_/a_1000_472# _053_ 0.029433f
C8428 _097_ FILLER_0_15_180/a_124_375# 0.007065f
C8429 FILLER_0_17_72/a_2276_472# net36 0.004399f
C8430 FILLER_0_17_38/a_124_375# _041_ 0.009172f
C8431 _099_ net30 0.05959f
C8432 FILLER_0_14_50/a_124_375# _174_ 0.033245f
C8433 output44/a_224_472# FILLER_0_19_28/a_36_472# 0.023414f
C8434 net69 vss 0.34555f
C8435 vss _201_/a_67_603# 0.012925f
C8436 _442_/a_2248_156# _158_ 0.001288f
C8437 mask\[9\] _438_/a_2248_156# 0.036436f
C8438 net27 FILLER_0_12_236/a_484_472# 0.042937f
C8439 _064_ _446_/a_36_151# 0.006723f
C8440 _126_ _131_ 0.626666f
C8441 trim[1] net40 0.043114f
C8442 net52 _442_/a_796_472# 0.004871f
C8443 FILLER_0_18_177/a_1380_472# vdd 0.005692f
C8444 FILLER_0_18_177/a_932_472# vss -0.001894f
C8445 net47 _039_ 0.042757f
C8446 output8/a_224_472# FILLER_0_3_221/a_484_472# 0.001699f
C8447 _005_ _416_/a_448_472# 0.04044f
C8448 result[9] _419_/a_1308_423# 0.012036f
C8449 fanout53/a_36_160# FILLER_0_16_154/a_484_472# 0.014774f
C8450 net80 net57 0.002913f
C8451 FILLER_0_9_60/a_124_375# vdd 0.005798f
C8452 _450_/a_1284_156# _039_ 0.001226f
C8453 _450_/a_3129_107# cal_count\[0\] 0.020971f
C8454 _341_/a_49_472# net56 0.018486f
C8455 net15 FILLER_0_23_60/a_124_375# 0.038706f
C8456 FILLER_0_19_28/a_572_375# _452_/a_36_151# 0.0027f
C8457 _360_/a_36_160# _133_ 0.001878f
C8458 net69 _441_/a_2248_156# 0.036635f
C8459 net63 FILLER_0_19_195/a_36_472# 0.030832f
C8460 net65 net5 0.004409f
C8461 _100_ vdd 0.212037f
C8462 FILLER_0_17_218/a_124_375# vdd 0.00593f
C8463 _272_/a_36_472# net76 0.04597f
C8464 _425_/a_1204_472# vdd 0.015969f
C8465 state\[0\] _273_/a_36_68# 0.012187f
C8466 _152_ vss 0.140215f
C8467 mask\[7\] FILLER_0_22_128/a_1380_472# 0.015814f
C8468 _069_ _429_/a_1308_423# 0.027468f
C8469 net37 FILLER_0_6_231/a_484_472# 0.004323f
C8470 _297_/a_36_472# vdd 0.042391f
C8471 FILLER_0_19_125/a_36_472# _345_/a_36_160# 0.006647f
C8472 FILLER_0_5_128/a_36_472# net47 0.008459f
C8473 net53 _427_/a_2248_156# 0.038716f
C8474 _075_ net59 0.01129f
C8475 trim_mask\[0\] vdd 0.154098f
C8476 net64 FILLER_0_9_270/a_484_472# 0.017924f
C8477 ctln[7] vss 0.132613f
C8478 _067_ FILLER_0_12_20/a_484_472# 0.011046f
C8479 _147_ _208_/a_36_160# 0.006056f
C8480 output28/a_224_472# fanout79/a_36_160# 0.022393f
C8481 _394_/a_56_524# FILLER_0_15_59/a_572_375# 0.003413f
C8482 _423_/a_36_151# FILLER_0_23_44/a_124_375# 0.059049f
C8483 _448_/a_2248_156# net22 0.07925f
C8484 net15 FILLER_0_17_72/a_572_375# 0.003021f
C8485 _098_ FILLER_0_15_212/a_572_375# 0.009099f
C8486 _060_ net22 0.533421f
C8487 _428_/a_1000_472# net74 0.00735f
C8488 _176_ net53 0.083005f
C8489 output7/a_224_472# net40 0.009154f
C8490 fanout82/a_36_113# output37/a_224_472# 0.023409f
C8491 net52 _439_/a_2665_112# 0.00117f
C8492 FILLER_0_4_144/a_124_375# net23 0.011315f
C8493 _079_ FILLER_0_6_231/a_572_375# 0.002768f
C8494 _138_ vss 0.006962f
C8495 mask\[8\] mask\[9\] 0.078756f
C8496 net58 net59 0.066534f
C8497 _106_ net33 0.001049f
C8498 FILLER_0_4_49/a_36_472# vss 0.001931f
C8499 FILLER_0_4_49/a_484_472# vdd 0.003356f
C8500 FILLER_0_4_144/a_572_375# trim_mask\[4\] 0.014071f
C8501 net54 _438_/a_2665_112# 0.032855f
C8502 ctlp[6] net54 0.00409f
C8503 _432_/a_2248_156# net63 0.047337f
C8504 _020_ fanout70/a_36_113# 0.001266f
C8505 FILLER_0_4_144/a_572_375# net47 0.011686f
C8506 _119_ _056_ 0.008929f
C8507 _093_ FILLER_0_17_142/a_572_375# 0.009547f
C8508 _176_ FILLER_0_10_107/a_484_472# 0.009571f
C8509 FILLER_0_24_63/a_124_375# ctlp[9] 0.002726f
C8510 FILLER_0_22_86/a_36_472# vdd -0.001506f
C8511 FILLER_0_22_86/a_1468_375# vss 0.013146f
C8512 _132_ FILLER_0_14_107/a_932_472# 0.014911f
C8513 output8/a_224_472# cal_itt\[1\] 0.003894f
C8514 _002_ FILLER_0_4_197/a_124_375# 0.001406f
C8515 FILLER_0_11_78/a_484_472# _120_ 0.016839f
C8516 FILLER_0_15_142/a_572_375# net56 0.001809f
C8517 trim_val\[4\] _387_/a_36_113# 0.005339f
C8518 _038_ FILLER_0_11_78/a_484_472# 0.001782f
C8519 net63 FILLER_0_18_177/a_2276_472# 0.012025f
C8520 mask\[4\] FILLER_0_19_171/a_1020_375# 0.006236f
C8521 FILLER_0_9_223/a_124_375# state\[0\] 0.002912f
C8522 _430_/a_2665_112# net36 0.003477f
C8523 FILLER_0_22_128/a_2724_472# vdd 0.005923f
C8524 FILLER_0_22_128/a_2276_472# vss 0.02979f
C8525 _035_ trim[0] 0.171633f
C8526 _075_ _122_ 0.030339f
C8527 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_572_375# 0.086635f
C8528 _021_ FILLER_0_18_171/a_124_375# 0.004621f
C8529 _236_/a_36_160# net67 0.009332f
C8530 FILLER_0_7_72/a_124_375# vdd 0.01526f
C8531 _412_/a_2248_156# net58 0.010702f
C8532 net56 FILLER_0_18_139/a_932_472# 0.011079f
C8533 net59 net21 0.157689f
C8534 output38/a_224_472# _446_/a_36_151# 0.117966f
C8535 ctlp[0] net17 0.006778f
C8536 FILLER_0_5_128/a_36_472# net74 0.01163f
C8537 _211_/a_36_160# vss 0.002041f
C8538 output32/a_224_472# _419_/a_1308_423# 0.005111f
C8539 net63 FILLER_0_17_218/a_36_472# 0.003889f
C8540 net45 net17 0.192181f
C8541 _013_ vss 0.163674f
C8542 _445_/a_796_472# _034_ 0.009261f
C8543 _053_ FILLER_0_6_47/a_484_472# 0.006301f
C8544 FILLER_0_0_198/a_124_375# net21 0.004256f
C8545 _116_ net22 0.122052f
C8546 _119_ _068_ 0.040944f
C8547 net36 FILLER_0_18_76/a_36_472# 0.001728f
C8548 net82 FILLER_0_3_172/a_932_472# 0.007986f
C8549 FILLER_0_8_263/a_124_375# vdd 0.032664f
C8550 net54 net35 0.114666f
C8551 _124_ FILLER_0_10_107/a_484_472# 0.00438f
C8552 _093_ FILLER_0_18_107/a_1380_472# 0.001782f
C8553 en_co_clk FILLER_0_13_100/a_124_375# 0.002325f
C8554 vdd FILLER_0_14_235/a_124_375# -0.011193f
C8555 mask\[5\] _340_/a_36_160# 0.031249f
C8556 _064_ _447_/a_36_151# 0.004185f
C8557 FILLER_0_3_172/a_36_472# net65 0.014671f
C8558 _098_ FILLER_0_15_205/a_124_375# 0.009558f
C8559 _446_/a_2248_156# vdd 0.059236f
C8560 _322_/a_848_380# net74 0.00168f
C8561 _415_/a_36_151# _426_/a_36_151# 0.002121f
C8562 _173_ _039_ 0.0326f
C8563 net58 net64 0.590523f
C8564 fanout66/a_36_113# net68 0.01746f
C8565 net81 FILLER_0_9_270/a_124_375# 0.014206f
C8566 result[1] net18 0.056799f
C8567 _210_/a_67_603# vdd 0.028101f
C8568 _127_ _069_ 0.048146f
C8569 calibrate _122_ 0.074949f
C8570 _116_ _311_/a_2700_473# 0.001555f
C8571 _443_/a_1308_423# vss 0.031091f
C8572 FILLER_0_14_99/a_124_375# _451_/a_36_151# 0.001441f
C8573 _431_/a_796_472# _136_ 0.009889f
C8574 calibrate FILLER_0_7_233/a_124_375# 0.011958f
C8575 fanout67/a_36_160# FILLER_0_9_60/a_124_375# 0.02985f
C8576 _076_ _055_ 0.056585f
C8577 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_124_375# 0.012001f
C8578 cal_itt\[2\] net8 0.057335f
C8579 net48 _425_/a_36_151# 0.020568f
C8580 _448_/a_2248_156# vdd 0.008296f
C8581 net52 FILLER_0_6_47/a_2724_472# 0.011079f
C8582 net64 calibrate 0.096329f
C8583 _444_/a_1308_423# FILLER_0_8_24/a_36_472# 0.009119f
C8584 net15 net35 0.01797f
C8585 result[4] _418_/a_448_472# 0.004918f
C8586 _122_ net21 0.026632f
C8587 _060_ vdd 0.349556f
C8588 _113_ vss 0.147905f
C8589 _155_ FILLER_0_7_104/a_124_375# 0.007925f
C8590 _165_ _164_ 0.351097f
C8591 calibrate _169_ 0.001883f
C8592 output47/a_224_472# _185_ 0.001177f
C8593 _423_/a_36_151# vdd 0.088377f
C8594 _255_/a_224_552# _074_ 0.005907f
C8595 _392_/a_36_68# _067_ 0.020085f
C8596 FILLER_0_22_177/a_124_375# _023_ 0.001195f
C8597 clk net59 0.052607f
C8598 FILLER_0_5_54/a_484_472# net47 0.006652f
C8599 net68 _453_/a_1308_423# 0.002195f
C8600 net57 _428_/a_796_472# 0.003017f
C8601 net72 _012_ 0.002382f
C8602 _291_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C8603 FILLER_0_3_54/a_36_472# net40 0.069702f
C8604 ctlp[1] _009_ 0.085933f
C8605 net62 output29/a_224_472# 0.138536f
C8606 _217_/a_36_160# _052_ 0.016695f
C8607 net74 _372_/a_1194_69# 0.002006f
C8608 net20 _060_ 0.0426f
C8609 _016_ FILLER_0_12_136/a_1020_375# 0.001659f
C8610 _242_/a_36_160# FILLER_0_5_164/a_36_472# 0.193804f
C8611 _255_/a_224_552# _076_ 0.081663f
C8612 _057_ _070_ 0.033401f
C8613 _044_ FILLER_0_14_263/a_124_375# 0.001047f
C8614 _126_ FILLER_0_11_101/a_124_375# 0.011403f
C8615 FILLER_0_18_100/a_124_375# FILLER_0_18_107/a_36_472# 0.012267f
C8616 _126_ _076_ 0.005517f
C8617 FILLER_0_14_81/a_124_375# _451_/a_3129_107# 0.009542f
C8618 mask\[4\] _433_/a_2248_156# 0.001082f
C8619 _130_ _325_/a_224_472# 0.001685f
C8620 FILLER_0_17_72/a_3260_375# vss 0.052993f
C8621 FILLER_0_17_72/a_36_472# vdd 0.111688f
C8622 _134_ FILLER_0_10_107/a_572_375# 0.047331f
C8623 _048_ _204_/a_67_603# 0.004547f
C8624 _136_ FILLER_0_17_142/a_572_375# 0.001371f
C8625 cal_itt\[3\] _079_ 0.015743f
C8626 _064_ _444_/a_36_151# 0.001296f
C8627 _148_ _025_ 0.007252f
C8628 _412_/a_2560_156# cal_itt\[1\] 0.00454f
C8629 _132_ FILLER_0_18_107/a_1916_375# 0.019011f
C8630 FILLER_0_4_107/a_1380_472# vss 0.004455f
C8631 mask\[5\] _348_/a_49_472# 0.025962f
C8632 _075_ FILLER_0_5_206/a_124_375# 0.001024f
C8633 vss FILLER_0_6_37/a_124_375# 0.030885f
C8634 vdd FILLER_0_6_37/a_36_472# 0.138008f
C8635 _183_ _182_ 0.002134f
C8636 _370_/a_848_380# net23 0.001196f
C8637 _077_ _067_ 0.090648f
C8638 _142_ FILLER_0_17_133/a_36_472# 0.069383f
C8639 _427_/a_1308_423# vss 0.030292f
C8640 net72 FILLER_0_15_59/a_484_472# 0.008749f
C8641 net17 _450_/a_3129_107# 0.004255f
C8642 net52 FILLER_0_2_111/a_932_472# 0.061249f
C8643 _043_ FILLER_0_13_72/a_484_472# 0.016114f
C8644 _370_/a_692_472# net47 0.001021f
C8645 net18 _007_ 0.060872f
C8646 _164_ net40 0.048933f
C8647 _256_/a_716_497# calibrate 0.001066f
C8648 _116_ vdd 0.399137f
C8649 net56 state\[1\] 0.007364f
C8650 _444_/a_36_151# net42 0.006866f
C8651 trim_mask\[2\] FILLER_0_2_93/a_484_472# 0.001424f
C8652 _415_/a_2248_156# vss 0.00818f
C8653 _091_ FILLER_0_15_212/a_36_472# 0.007355f
C8654 net52 _440_/a_2248_156# 0.028463f
C8655 _053_ _161_ 0.001047f
C8656 net80 _340_/a_36_160# 0.004225f
C8657 mask\[3\] FILLER_0_18_177/a_2364_375# 0.002935f
C8658 _239_/a_36_160# net17 0.014703f
C8659 _144_ FILLER_0_22_128/a_2812_375# 0.001601f
C8660 net60 _421_/a_1288_156# 0.001147f
C8661 mask\[4\] FILLER_0_20_177/a_36_472# 0.001215f
C8662 net82 _032_ 0.014269f
C8663 net72 net74 0.035298f
C8664 FILLER_0_10_78/a_932_472# _176_ 0.0109f
C8665 trimb[2] net43 0.011999f
C8666 _095_ FILLER_0_13_72/a_572_375# 0.003559f
C8667 output24/a_224_472# net71 0.001495f
C8668 FILLER_0_6_79/a_124_375# _164_ 0.061565f
C8669 _100_ _283_/a_36_472# 0.033597f
C8670 _408_/a_718_524# vdd 0.002635f
C8671 net71 vss 0.335256f
C8672 _024_ net23 0.001994f
C8673 net49 _440_/a_2248_156# 0.025137f
C8674 net82 trim_val\[4\] 0.511271f
C8675 FILLER_0_10_78/a_572_375# _115_ 0.004573f
C8676 FILLER_0_4_185/a_36_472# _002_ 0.004231f
C8677 _053_ _129_ 0.003479f
C8678 FILLER_0_7_59/a_124_375# trim_val\[0\] 0.002169f
C8679 net29 net36 0.370099f
C8680 trim_mask\[2\] trim_val\[2\] 0.21814f
C8681 FILLER_0_18_171/a_36_472# mask\[3\] 0.00262f
C8682 _078_ FILLER_0_4_213/a_484_472# 0.003702f
C8683 FILLER_0_16_73/a_484_472# net55 0.004188f
C8684 trim_val\[4\] fanout57/a_36_113# 0.078297f
C8685 _447_/a_2248_156# vdd 0.009094f
C8686 _303_/a_36_472# _110_ 0.001606f
C8687 result[9] result[2] 0.001669f
C8688 net57 FILLER_0_8_156/a_484_472# 0.008895f
C8689 FILLER_0_16_57/a_36_472# cal_count\[1\] 0.002116f
C8690 _067_ _120_ 0.031156f
C8691 _118_ vdd 0.292155f
C8692 _038_ _067_ 0.503045f
C8693 FILLER_0_12_2/a_484_472# _039_ 0.003082f
C8694 net23 FILLER_0_22_128/a_2812_375# 0.050811f
C8695 _137_ FILLER_0_16_154/a_932_472# 0.004753f
C8696 _086_ _055_ 0.113385f
C8697 _292_/a_36_160# _047_ 0.001291f
C8698 net78 _420_/a_448_472# 0.001091f
C8699 net54 _433_/a_2665_112# 0.047439f
C8700 FILLER_0_5_72/a_484_472# _440_/a_36_151# 0.001723f
C8701 FILLER_0_18_107/a_124_375# mask\[9\] 0.006029f
C8702 FILLER_0_17_64/a_124_375# FILLER_0_17_56/a_572_375# 0.012001f
C8703 net61 net62 0.874859f
C8704 FILLER_0_21_125/a_484_472# _433_/a_36_151# 0.001723f
C8705 _036_ net69 0.353233f
C8706 _365_/a_692_472# _156_ 0.001127f
C8707 net74 _370_/a_692_472# 0.005066f
C8708 FILLER_0_17_218/a_124_375# _069_ 0.003162f
C8709 _016_ _428_/a_1308_423# 0.00107f
C8710 _414_/a_2665_112# _074_ 0.004912f
C8711 _109_ vdd 0.059259f
C8712 FILLER_0_18_2/a_2276_472# _452_/a_1040_527# 0.008652f
C8713 FILLER_0_18_2/a_484_472# _452_/a_2225_156# 0.019521f
C8714 _440_/a_36_151# _160_ 0.002966f
C8715 net52 _376_/a_36_160# 0.00267f
C8716 _449_/a_36_151# FILLER_0_13_72/a_36_472# 0.001723f
C8717 net32 output34/a_224_472# 0.027498f
C8718 net53 FILLER_0_17_142/a_572_375# 0.023771f
C8719 _180_ FILLER_0_15_59/a_36_472# 0.087308f
C8720 _086_ _255_/a_224_552# 0.073601f
C8721 FILLER_0_8_37/a_484_472# _160_ 0.001767f
C8722 net80 net36 0.036729f
C8723 net65 FILLER_0_2_177/a_484_472# 0.01675f
C8724 _029_ FILLER_0_5_88/a_36_472# 0.007596f
C8725 _086_ _126_ 0.063495f
C8726 _103_ _418_/a_448_472# 0.002678f
C8727 _079_ _265_/a_244_68# 0.021777f
C8728 _449_/a_1000_472# net55 0.001617f
C8729 _091_ FILLER_0_12_220/a_932_472# 0.001638f
C8730 ctlp[1] FILLER_0_23_290/a_36_472# 0.038596f
C8731 _116_ _373_/a_244_68# 0.001213f
C8732 _422_/a_796_472# _109_ 0.002086f
C8733 _123_ vdd 0.214703f
C8734 _113_ _279_/a_652_68# 0.001425f
C8735 net81 net22 0.064261f
C8736 FILLER_0_7_146/a_124_375# net37 0.005315f
C8737 net54 vdd 0.877573f
C8738 _430_/a_1308_423# net21 0.008506f
C8739 _444_/a_2248_156# vdd 0.041347f
C8740 net41 FILLER_0_17_38/a_36_472# 0.001308f
C8741 _073_ vdd 0.258125f
C8742 FILLER_0_0_232/a_36_472# vss 0.007185f
C8743 _330_/a_224_472# vdd 0.001701f
C8744 _008_ _198_/a_67_603# 0.012332f
C8745 _176_ _389_/a_36_148# 0.060256f
C8746 net78 _419_/a_1308_423# 0.018598f
C8747 _046_ _099_ 0.005245f
C8748 net64 mask\[1\] 0.038611f
C8749 _166_ _034_ 0.001936f
C8750 _412_/a_1308_423# net59 0.00291f
C8751 net20 _123_ 0.034801f
C8752 _430_/a_1204_472# net21 0.006991f
C8753 _440_/a_2560_156# _164_ 0.003934f
C8754 ctlp[2] _300_/a_224_472# 0.002954f
C8755 _375_/a_36_68# _161_ 0.028567f
C8756 _077_ net23 0.0245f
C8757 net65 FILLER_0_1_212/a_124_375# 0.005253f
C8758 FILLER_0_20_2/a_572_375# net43 0.051705f
C8759 net20 _073_ 0.437482f
C8760 output23/a_224_472# FILLER_0_22_128/a_2364_375# 0.002439f
C8761 _010_ _420_/a_2560_156# 0.070902f
C8762 _337_/a_49_472# vdd 0.028131f
C8763 FILLER_0_4_185/a_124_375# FILLER_0_4_177/a_572_375# 0.012001f
C8764 FILLER_0_5_212/a_36_472# net22 0.0015f
C8765 FILLER_0_7_162/a_124_375# calibrate 0.014255f
C8766 mask\[8\] _437_/a_2248_156# 0.004415f
C8767 _012_ FILLER_0_23_60/a_124_375# 0.002827f
C8768 _131_ _160_ 0.003984f
C8769 FILLER_0_21_28/a_1020_375# vdd 0.04353f
C8770 net15 vdd 2.073988f
C8771 FILLER_0_11_78/a_36_472# vdd -0.001328f
C8772 FILLER_0_11_78/a_572_375# vss 0.004808f
C8773 ctlp[2] _420_/a_2248_156# 0.001156f
C8774 _326_/a_36_160# _131_ 0.023688f
C8775 net42 _054_ 0.006314f
C8776 _431_/a_2665_112# net36 0.001523f
C8777 net55 FILLER_0_21_28/a_2724_472# 0.049771f
C8778 output10/a_224_472# cal_itt\[0\] 0.008003f
C8779 FILLER_0_15_290/a_124_375# FILLER_0_15_282/a_572_375# 0.012001f
C8780 _265_/a_244_68# cal_itt\[1\] 0.024108f
C8781 _064_ vss 0.228443f
C8782 net82 FILLER_0_4_213/a_572_375# 0.00123f
C8783 _053_ _220_/a_255_603# 0.001311f
C8784 net67 FILLER_0_9_60/a_572_375# 0.011073f
C8785 net27 _415_/a_448_472# 0.05785f
C8786 net63 _435_/a_448_472# 0.009878f
C8787 _253_/a_1100_68# _084_ 0.001651f
C8788 _116_ _279_/a_244_68# 0.001752f
C8789 ctln[8] _168_ 0.001145f
C8790 _228_/a_36_68# net22 0.052558f
C8791 _055_ _090_ 0.040233f
C8792 _093_ FILLER_0_17_104/a_1020_375# 0.01418f
C8793 FILLER_0_16_107/a_36_472# _451_/a_36_151# 0.059367f
C8794 FILLER_0_3_142/a_36_472# _370_/a_848_380# 0.001207f
C8795 FILLER_0_4_107/a_572_375# net47 0.006041f
C8796 _053_ FILLER_0_7_59/a_484_472# 0.013665f
C8797 net15 _441_/a_1204_472# 0.005939f
C8798 output48/a_224_472# net59 0.039277f
C8799 FILLER_0_5_164/a_124_375# net37 0.008158f
C8800 _142_ FILLER_0_17_161/a_36_472# 0.00657f
C8801 _140_ _023_ 0.079452f
C8802 FILLER_0_6_90/a_572_375# vdd 0.028324f
C8803 output47/a_224_472# net55 0.160037f
C8804 FILLER_0_16_89/a_1380_472# FILLER_0_17_72/a_3260_375# 0.001723f
C8805 net42 vss 0.017902f
C8806 mask\[5\] FILLER_0_20_177/a_124_375# 0.013531f
C8807 _120_ net23 0.147166f
C8808 _418_/a_1000_472# vss 0.001193f
C8809 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_36_472# 0.086635f
C8810 _333_/a_36_160# _097_ 0.001332f
C8811 _171_ FILLER_0_10_94/a_484_472# 0.001446f
C8812 FILLER_0_22_177/a_1380_472# net33 0.016037f
C8813 _073_ net9 0.005417f
C8814 FILLER_0_18_2/a_1468_375# net38 0.016983f
C8815 _115_ net74 0.033145f
C8816 _122_ FILLER_0_5_181/a_124_375# 0.001352f
C8817 net52 FILLER_0_9_72/a_1468_375# 0.003576f
C8818 _100_ FILLER_0_12_236/a_572_375# 0.015109f
C8819 FILLER_0_13_142/a_1020_375# net23 0.047331f
C8820 net81 FILLER_0_15_235/a_572_375# 0.009675f
C8821 _445_/a_2248_156# net17 0.06175f
C8822 net39 vdd 0.2282f
C8823 _255_/a_224_552# _090_ 0.001598f
C8824 FILLER_0_1_266/a_484_472# vdd 0.003622f
C8825 _414_/a_2665_112# _081_ 0.00247f
C8826 _042_ vss 0.008272f
C8827 net51 vdd 0.692054f
C8828 _069_ _060_ 0.538161f
C8829 _126_ _090_ 0.003538f
C8830 _425_/a_36_151# net37 0.003145f
C8831 _430_/a_448_472# net21 0.03842f
C8832 _002_ net82 0.034599f
C8833 FILLER_0_24_96/a_36_472# output25/a_224_472# 0.010475f
C8834 _040_ FILLER_0_16_115/a_36_472# 0.001876f
C8835 _053_ _068_ 0.066662f
C8836 net81 vdd 1.658963f
C8837 FILLER_0_18_2/a_484_472# net44 0.047503f
C8838 _095_ _113_ 0.004037f
C8839 _144_ mask\[6\] 0.230129f
C8840 FILLER_0_17_142/a_124_375# FILLER_0_17_133/a_124_375# 0.003228f
C8841 _144_ mask\[8\] 0.131592f
C8842 FILLER_0_11_109/a_124_375# _120_ 0.016902f
C8843 _378_/a_224_472# _165_ 0.00481f
C8844 _402_/a_2172_497# _180_ 0.001094f
C8845 FILLER_0_4_144/a_572_375# FILLER_0_5_148/a_124_375# 0.05841f
C8846 _137_ FILLER_0_19_155/a_124_375# 0.00129f
C8847 _428_/a_2560_156# _131_ 0.002853f
C8848 output47/a_224_472# net17 0.081437f
C8849 FILLER_0_1_98/a_124_375# vdd 0.036865f
C8850 FILLER_0_5_88/a_36_472# _163_ 0.006541f
C8851 _442_/a_36_151# FILLER_0_2_127/a_124_375# 0.001597f
C8852 mask\[2\] net21 0.033368f
C8853 net20 net81 0.036173f
C8854 result[6] net61 0.120359f
C8855 net38 _221_/a_36_160# 0.029767f
C8856 net82 FILLER_0_3_221/a_1020_375# 0.010208f
C8857 _333_/a_36_160# mask\[2\] 0.022517f
C8858 _350_/a_49_472# vdd 0.026837f
C8859 vss FILLER_0_4_91/a_484_472# 0.003328f
C8860 FILLER_0_8_247/a_572_375# calibrate 0.008498f
C8861 result[7] FILLER_0_23_274/a_124_375# 0.017938f
C8862 ctlp[1] FILLER_0_24_274/a_932_472# 0.003603f
C8863 _065_ _447_/a_36_151# 0.043351f
C8864 _027_ net71 0.057875f
C8865 FILLER_0_3_172/a_2276_472# net22 0.012151f
C8866 FILLER_0_5_212/a_124_375# vss 0.006344f
C8867 FILLER_0_5_212/a_36_472# vdd 0.107657f
C8868 output48/a_224_472# net64 0.002845f
C8869 mask\[9\] _423_/a_2665_112# 0.001735f
C8870 mask\[5\] _295_/a_36_472# 0.034027f
C8871 _106_ vdd 0.232973f
C8872 _142_ FILLER_0_16_154/a_124_375# 0.004001f
C8873 FILLER_0_12_20/a_572_375# FILLER_0_12_28/a_124_375# 0.012001f
C8874 FILLER_0_12_136/a_932_472# _127_ 0.002804f
C8875 _422_/a_2665_112# mask\[7\] 0.028271f
C8876 net16 ctln[9] 0.07797f
C8877 output36/a_224_472# net18 0.010751f
C8878 _086_ state\[1\] 0.043298f
C8879 FILLER_0_17_56/a_36_472# _404_/a_36_472# 0.004546f
C8880 mask\[8\] net25 0.035648f
C8881 net23 mask\[6\] 0.025699f
C8882 ctlp[1] net33 0.11288f
C8883 FILLER_0_10_214/a_36_472# _070_ 0.014734f
C8884 net18 net30 0.09055f
C8885 net19 _418_/a_2665_112# 0.040822f
C8886 output36/a_224_472# _196_/a_36_160# 0.001309f
C8887 _427_/a_1308_423# _095_ 0.022677f
C8888 _069_ _116_ 0.390834f
C8889 _150_ mask\[9\] 0.162185f
C8890 _106_ net20 0.050151f
C8891 _091_ _019_ 0.031681f
C8892 net62 FILLER_0_15_290/a_124_375# 0.034614f
C8893 mask\[0\] net64 0.45093f
C8894 fanout75/a_36_113# _317_/a_36_113# 0.001442f
C8895 net75 FILLER_0_8_247/a_932_472# 0.006746f
C8896 FILLER_0_15_142/a_124_375# _427_/a_36_151# 0.059049f
C8897 fanout52/a_36_160# net23 0.009496f
C8898 FILLER_0_10_78/a_572_375# FILLER_0_9_72/a_1380_472# 0.001543f
C8899 _228_/a_36_68# vdd 0.036391f
C8900 FILLER_0_4_123/a_124_375# _160_ 0.038272f
C8901 _066_ _386_/a_692_472# 0.001958f
C8902 net38 FILLER_0_20_15/a_36_472# 0.070475f
C8903 _115_ _449_/a_2665_112# 0.00947f
C8904 net80 FILLER_0_20_177/a_124_375# 0.001198f
C8905 net35 _012_ 0.007543f
C8906 _428_/a_1308_423# _017_ 0.005962f
C8907 _428_/a_448_472# net53 0.001959f
C8908 output21/a_224_472# net32 0.017976f
C8909 _369_/a_36_68# vss 0.002343f
C8910 net68 trim_mask\[1\] 0.054055f
C8911 _162_ _374_/a_36_68# 0.005729f
C8912 _044_ vss 0.038421f
C8913 _122_ _242_/a_36_160# 0.005377f
C8914 comp net44 0.079931f
C8915 _413_/a_2665_112# FILLER_0_3_212/a_124_375# 0.001077f
C8916 FILLER_0_20_169/a_36_472# _140_ 0.023696f
C8917 state\[2\] net23 0.331644f
C8918 FILLER_0_7_104/a_484_472# FILLER_0_9_105/a_572_375# 0.001188f
C8919 FILLER_0_11_142/a_484_472# vss 0.033416f
C8920 FILLER_0_18_107/a_3260_375# vss 0.056926f
C8921 FILLER_0_18_107/a_36_472# vdd 0.116746f
C8922 _139_ _137_ 0.093639f
C8923 _069_ _118_ 0.010986f
C8924 _434_/a_796_472# mask\[6\] 0.004416f
C8925 output20/a_224_472# _109_ 0.003452f
C8926 _414_/a_448_472# _089_ 0.003905f
C8927 FILLER_0_7_104/a_36_472# vdd 0.096343f
C8928 FILLER_0_7_104/a_1468_375# vss 0.003442f
C8929 _242_/a_36_160# _169_ 0.051038f
C8930 _277_/a_36_160# vdd 0.115507f
C8931 trim_mask\[1\] _156_ 0.007519f
C8932 fanout50/a_36_160# _168_ 0.033707f
C8933 net52 _384_/a_224_472# 0.001238f
C8934 net47 _167_ 0.003019f
C8935 net44 _245_/a_672_472# 0.001285f
C8936 net55 FILLER_0_21_60/a_36_472# 0.06794f
C8937 _053_ _152_ 0.032961f
C8938 _414_/a_36_151# _055_ 0.001987f
C8939 _077_ FILLER_0_9_28/a_2724_472# 0.006001f
C8940 mask\[4\] FILLER_0_18_139/a_1468_375# 0.023004f
C8941 net52 _441_/a_448_472# 0.04874f
C8942 FILLER_0_4_107/a_572_375# _154_ 0.052251f
C8943 FILLER_0_17_72/a_932_472# FILLER_0_18_76/a_484_472# 0.05841f
C8944 output40/a_224_472# net40 0.0374f
C8945 _088_ FILLER_0_3_212/a_124_375# 0.0042f
C8946 FILLER_0_12_236/a_572_375# _060_ 0.001597f
C8947 net64 _099_ 0.007017f
C8948 _076_ _160_ 0.006506f
C8949 _415_/a_448_472# net18 0.057688f
C8950 _077_ net57 0.025864f
C8951 _161_ _070_ 0.027757f
C8952 FILLER_0_1_212/a_36_472# net59 0.002567f
C8953 net2 vdd 0.434557f
C8954 _277_/a_36_160# net20 0.015569f
C8955 net18 _417_/a_36_151# 0.020548f
C8956 _143_ FILLER_0_18_139/a_1380_472# 0.002226f
C8957 _417_/a_448_472# net30 0.042386f
C8958 _062_ _226_/a_1044_68# 0.001944f
C8959 _091_ FILLER_0_13_212/a_484_472# 0.04953f
C8960 _072_ _375_/a_1388_497# 0.001138f
C8961 _441_/a_448_472# net49 0.001245f
C8962 mask\[9\] _026_ 0.002924f
C8963 output35/a_224_472# _435_/a_36_151# 0.001362f
C8964 _431_/a_448_472# net73 0.050964f
C8965 _157_ _156_ 0.005264f
C8966 net15 _423_/a_2560_156# 0.007083f
C8967 _097_ mask\[1\] 0.001232f
C8968 net50 FILLER_0_9_60/a_36_472# 0.001914f
C8969 result[7] FILLER_0_24_274/a_1020_375# 0.006125f
C8970 _428_/a_36_151# FILLER_0_14_107/a_572_375# 0.001597f
C8971 _449_/a_2560_156# _038_ 0.010532f
C8972 net61 _422_/a_36_151# 0.003736f
C8973 FILLER_0_3_172/a_2276_472# vdd 0.00806f
C8974 _131_ _133_ 0.20118f
C8975 _129_ _070_ 0.056776f
C8976 output46/a_224_472# net38 0.003296f
C8977 trim_mask\[4\] net22 0.027368f
C8978 net67 trim_mask\[1\] 0.01761f
C8979 FILLER_0_9_223/a_572_375# _128_ 0.006559f
C8980 _076_ _223_/a_36_160# 0.001756f
C8981 _057_ calibrate 0.002047f
C8982 FILLER_0_19_171/a_484_472# _434_/a_36_151# 0.002841f
C8983 fanout71/a_36_113# _149_ 0.001315f
C8984 state\[1\] _090_ 0.087906f
C8985 output11/a_224_472# ctln[4] 0.072677f
C8986 output7/a_224_472# net7 0.01565f
C8987 _077_ _439_/a_2248_156# 0.038814f
C8988 _012_ FILLER_0_23_44/a_124_375# 0.002474f
C8989 net4 _246_/a_36_68# 0.003771f
C8990 net34 _295_/a_36_472# 0.032003f
C8991 mask\[4\] _343_/a_257_69# 0.001786f
C8992 _176_ _134_ 0.035146f
C8993 output13/a_224_472# net22 0.022308f
C8994 FILLER_0_4_213/a_124_375# net59 0.039014f
C8995 FILLER_0_10_78/a_572_375# vdd -0.014642f
C8996 _114_ _127_ 0.006414f
C8997 _144_ _433_/a_2248_156# 0.021805f
C8998 _044_ _416_/a_2248_156# 0.005198f
C8999 _346_/a_49_472# _141_ 0.104653f
C9000 net44 net6 0.005889f
C9001 _057_ net21 0.143214f
C9002 vdd clkc 0.190259f
C9003 result[5] _008_ 0.165753f
C9004 FILLER_0_15_212/a_36_472# net22 0.003143f
C9005 net57 _120_ 0.012391f
C9006 _255_/a_224_552# _163_ 0.002169f
C9007 _105_ _422_/a_2665_112# 0.011125f
C9008 _408_/a_728_93# _402_/a_56_567# 0.001359f
C9009 net52 cal_count\[3\] 0.348542f
C9010 net61 fanout77/a_36_113# 0.080943f
C9011 _002_ _413_/a_1204_472# 0.003057f
C9012 _045_ vdd 0.246567f
C9013 net35 FILLER_0_22_177/a_1380_472# 0.01447f
C9014 mask\[2\] mask\[1\] 0.059794f
C9015 ctlp[1] FILLER_0_23_282/a_572_375# 0.009848f
C9016 FILLER_0_5_172/a_124_375# net22 0.002388f
C9017 _053_ _377_/a_36_472# 0.023504f
C9018 _187_ _392_/a_36_68# 0.058263f
C9019 _431_/a_1308_423# _136_ 0.027758f
C9020 FILLER_0_14_181/a_36_472# vdd 0.027265f
C9021 FILLER_0_14_181/a_124_375# vss 0.009291f
C9022 net57 FILLER_0_13_142/a_1020_375# 0.009442f
C9023 _431_/a_1000_472# net73 0.035816f
C9024 FILLER_0_18_2/a_3172_472# FILLER_0_19_28/a_124_375# 0.001684f
C9025 _103_ _099_ 0.025799f
C9026 FILLER_0_15_205/a_124_375# net21 0.002912f
C9027 output11/a_224_472# _000_ 0.006606f
C9028 fanout82/a_36_113# net82 0.003741f
C9029 FILLER_0_1_212/a_124_375# net11 0.029766f
C9030 net75 _253_/a_672_68# 0.003771f
C9031 valid vdd 0.148392f
C9032 _322_/a_848_380# FILLER_0_9_142/a_124_375# 0.001721f
C9033 _140_ FILLER_0_22_128/a_2724_472# 0.004196f
C9034 _124_ _134_ 0.002508f
C9035 net23 _433_/a_2248_156# 0.005588f
C9036 net2 net9 0.001033f
C9037 mask\[4\] FILLER_0_18_209/a_484_472# 0.021522f
C9038 _383_/a_36_472# vss 0.002794f
C9039 ctln[2] net59 0.009218f
C9040 _412_/a_2665_112# en 0.015256f
C9041 net81 _283_/a_36_472# 0.032292f
C9042 net38 cal_count\[2\] 0.047195f
C9043 FILLER_0_8_247/a_1468_375# vss 0.054783f
C9044 FILLER_0_8_247/a_36_472# vdd 0.112197f
C9045 _114_ FILLER_0_11_101/a_36_472# 0.00501f
C9046 trim_val\[3\] FILLER_0_2_93/a_36_472# 0.015653f
C9047 _256_/a_1612_497# _076_ 0.001111f
C9048 FILLER_0_16_73/a_124_375# vdd 0.008987f
C9049 net17 _034_ 0.020793f
C9050 _055_ _117_ 0.242156f
C9051 _155_ _151_ 0.10611f
C9052 net55 FILLER_0_18_37/a_1020_375# 0.005661f
C9053 _136_ _335_/a_49_472# 0.039074f
C9054 _132_ _354_/a_49_472# 0.034372f
C9055 trim_val\[1\] _034_ 0.001535f
C9056 FILLER_0_12_136/a_1020_375# cal_count\[3\] 0.002916f
C9057 FILLER_0_2_111/a_1468_375# FILLER_0_2_127/a_124_375# 0.012001f
C9058 _322_/a_124_24# _128_ 0.02077f
C9059 _431_/a_448_472# _131_ 0.006194f
C9060 _168_ _164_ 0.092012f
C9061 net78 _421_/a_36_151# 0.001368f
C9062 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_572_375# 0.001597f
C9063 _077_ _187_ 0.058967f
C9064 FILLER_0_16_255/a_124_375# _094_ 0.004398f
C9065 _081_ _160_ 0.00816f
C9066 FILLER_0_5_206/a_36_472# FILLER_0_5_198/a_484_472# 0.013276f
C9067 output25/a_224_472# vss 0.080847f
C9068 _064_ _036_ 0.003286f
C9069 trim_mask\[2\] trim_val\[3\] 0.003342f
C9070 result[7] _421_/a_1456_156# 0.001009f
C9071 ctln[1] net59 0.053978f
C9072 mask\[5\] FILLER_0_21_206/a_124_375# 0.011644f
C9073 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_572_375# 0.086635f
C9074 net16 _379_/a_36_472# 0.01109f
C9075 _086_ _160_ 0.007038f
C9076 net38 _450_/a_448_472# 0.031891f
C9077 _011_ _422_/a_448_472# 0.044695f
C9078 _326_/a_36_160# _086_ 0.063565f
C9079 _028_ trim_mask\[1\] 0.148182f
C9080 FILLER_0_16_241/a_36_472# net36 0.001988f
C9081 _394_/a_728_93# FILLER_0_13_72/a_484_472# 0.018997f
C9082 _276_/a_36_160# FILLER_0_17_218/a_484_472# 0.001448f
C9083 output26/a_224_472# FILLER_0_23_44/a_932_472# 0.0323f
C9084 trim_mask\[4\] vdd 0.20602f
C9085 trimb[3] ctlp[0] 0.384753f
C9086 _098_ FILLER_0_15_180/a_484_472# 0.014511f
C9087 trimb[3] net45 0.001109f
C9088 _292_/a_36_160# mask\[5\] 0.007486f
C9089 _444_/a_2665_112# net67 0.03521f
C9090 net47 vdd 2.422992f
C9091 _015_ net4 0.003985f
C9092 net81 _069_ 0.034401f
C9093 net52 _443_/a_2665_112# 0.05031f
C9094 _074_ _374_/a_36_68# 0.001447f
C9095 net57 fanout52/a_36_160# 0.122432f
C9096 _315_/a_244_497# _120_ 0.006419f
C9097 FILLER_0_16_57/a_1020_375# vss 0.004487f
C9098 FILLER_0_16_57/a_1468_375# vdd 0.020146f
C9099 cal_itt\[2\] _073_ 0.202415f
C9100 _091_ _429_/a_1000_472# 0.029742f
C9101 output13/a_224_472# vdd 0.045929f
C9102 net35 _436_/a_1204_472# 0.005186f
C9103 _093_ _136_ 0.226819f
C9104 _174_ _179_ 0.003183f
C9105 net15 _449_/a_36_151# 0.020788f
C9106 _012_ vdd 0.261844f
C9107 _091_ _092_ 0.028594f
C9108 _374_/a_36_68# _076_ 0.026674f
C9109 _056_ _070_ 0.045548f
C9110 _065_ vss 0.230397f
C9111 _187_ _120_ 0.144679f
C9112 FILLER_0_15_212/a_1468_375# vss 0.060206f
C9113 FILLER_0_15_212/a_572_375# mask\[1\] 0.012463f
C9114 FILLER_0_15_212/a_36_472# vdd 0.105575f
C9115 net57 state\[2\] 1.25275f
C9116 _431_/a_448_472# net56 0.001464f
C9117 trim_mask\[2\] _367_/a_36_68# 0.001302f
C9118 _002_ net21 0.056631f
C9119 _093_ _438_/a_1000_472# 0.001556f
C9120 fanout71/a_36_113# FILLER_0_20_107/a_124_375# 0.002853f
C9121 _119_ FILLER_0_7_104/a_1468_375# 0.022368f
C9122 FILLER_0_7_72/a_1916_375# vss 0.001259f
C9123 FILLER_0_16_154/a_1380_472# vss 0.003609f
C9124 FILLER_0_5_172/a_124_375# vdd 0.028449f
C9125 FILLER_0_9_270/a_572_375# FILLER_0_9_282/a_36_472# 0.009654f
C9126 _445_/a_2665_112# _444_/a_448_472# 0.001178f
C9127 mask\[3\] vss 0.664467f
C9128 net57 _386_/a_692_472# 0.00409f
C9129 _011_ _108_ 0.036521f
C9130 FILLER_0_20_169/a_124_375# _098_ 0.019219f
C9131 net79 FILLER_0_15_282/a_124_375# 0.001058f
C9132 sample fanout59/a_36_160# 0.001854f
C9133 _106_ _069_ 0.006716f
C9134 trim_mask\[1\] FILLER_0_6_47/a_1916_375# 0.007169f
C9135 net62 FILLER_0_15_282/a_572_375# 0.007699f
C9136 _434_/a_1308_423# vdd 0.033494f
C9137 FILLER_0_19_111/a_484_472# vss 0.003811f
C9138 _067_ _450_/a_448_472# 0.003113f
C9139 _414_/a_1000_472# net21 0.042244f
C9140 _148_ _352_/a_257_69# 0.001417f
C9141 _181_ _182_ 0.02735f
C9142 _258_/a_36_160# vdd 0.00617f
C9143 FILLER_0_21_133/a_124_375# vss 0.015693f
C9144 cal net5 0.039735f
C9145 net38 _043_ 0.117134f
C9146 _052_ FILLER_0_18_53/a_124_375# 0.001585f
C9147 _132_ net73 0.460325f
C9148 net36 cal_count\[1\] 0.011481f
C9149 FILLER_0_15_59/a_484_472# vdd 0.010447f
C9150 FILLER_0_15_59/a_36_472# vss 0.00459f
C9151 _431_/a_36_151# _093_ 0.004862f
C9152 _254_/a_244_472# _074_ 0.002716f
C9153 _130_ _127_ 0.195571f
C9154 _098_ _201_/a_67_603# 0.005932f
C9155 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_124_375# 0.005439f
C9156 _258_/a_36_160# net20 0.041584f
C9157 FILLER_0_11_101/a_572_375# _070_ 0.011557f
C9158 _069_ _228_/a_36_68# 0.001676f
C9159 FILLER_0_5_109/a_484_472# FILLER_0_4_107/a_572_375# 0.001684f
C9160 _133_ _076_ 0.11688f
C9161 _070_ _068_ 1.019801f
C9162 net35 FILLER_0_22_128/a_572_375# 0.010439f
C9163 trim_val\[4\] FILLER_0_3_172/a_484_472# 0.002633f
C9164 net74 vdd 1.451847f
C9165 FILLER_0_7_146/a_36_472# _068_ 0.012745f
C9166 _114_ trim_mask\[0\] 0.021887f
C9167 net73 _427_/a_36_151# 0.006328f
C9168 _376_/a_36_160# FILLER_0_6_79/a_124_375# 0.004736f
C9169 _074_ _317_/a_36_113# 0.003383f
C9170 _064_ _445_/a_796_472# 0.00673f
C9171 _413_/a_1308_423# net65 0.022097f
C9172 FILLER_0_13_212/a_1380_472# net79 0.006824f
C9173 net27 _274_/a_244_497# 0.010334f
C9174 FILLER_0_5_117/a_36_472# FILLER_0_4_107/a_1020_375# 0.001684f
C9175 FILLER_0_4_107/a_484_472# FILLER_0_2_111/a_124_375# 0.001404f
C9176 _126_ FILLER_0_11_142/a_36_472# 0.001428f
C9177 _253_/a_36_68# vdd 0.016219f
C9178 net61 _419_/a_36_151# 0.019141f
C9179 net81 net28 0.034606f
C9180 FILLER_0_5_109/a_36_472# net47 0.005565f
C9181 net69 fanout49/a_36_160# 0.005942f
C9182 FILLER_0_9_28/a_1380_472# net51 0.002012f
C9183 _008_ net19 0.027093f
C9184 fanout58/a_36_160# net59 0.048057f
C9185 _415_/a_36_151# net62 0.00514f
C9186 mask\[1\] FILLER_0_15_205/a_124_375# 0.007883f
C9187 _106_ net31 0.035117f
C9188 net63 FILLER_0_15_212/a_932_472# 0.002269f
C9189 ctln[2] FILLER_0_1_266/a_124_375# 0.047145f
C9190 _067_ _043_ 0.189767f
C9191 _414_/a_1204_472# cal_itt\[3\] 0.052432f
C9192 fanout78/a_36_113# net18 0.001419f
C9193 _372_/a_170_472# vss 0.027819f
C9194 _232_/a_67_603# trim_val\[1\] 0.009588f
C9195 FILLER_0_4_197/a_1020_375# vss 0.001981f
C9196 FILLER_0_17_38/a_484_472# FILLER_0_18_37/a_484_472# 0.026657f
C9197 fanout75/a_36_113# net59 0.00817f
C9198 trim_mask\[4\] FILLER_0_2_165/a_124_375# 0.011181f
C9199 FILLER_0_12_220/a_484_472# vss 0.006724f
C9200 FILLER_0_12_220/a_932_472# vdd 0.003359f
C9201 FILLER_0_17_133/a_36_472# FILLER_0_19_134/a_124_375# 0.001188f
C9202 _058_ FILLER_0_8_156/a_572_375# 0.007692f
C9203 FILLER_0_19_125/a_36_472# FILLER_0_18_107/a_1916_375# 0.001684f
C9204 net58 FILLER_0_9_282/a_124_375# 0.021949f
C9205 _079_ net22 0.039221f
C9206 _173_ vdd 0.080629f
C9207 net63 _434_/a_1000_472# 0.002404f
C9208 FILLER_0_17_72/a_1020_375# _451_/a_3129_107# 0.001202f
C9209 FILLER_0_17_200/a_36_472# vss 0.001182f
C9210 net39 _445_/a_1308_423# 0.008252f
C9211 trim[1] _445_/a_36_151# 0.008362f
C9212 FILLER_0_20_193/a_484_472# FILLER_0_19_195/a_124_375# 0.001543f
C9213 FILLER_0_5_72/a_484_472# _029_ 0.004625f
C9214 FILLER_0_5_72/a_1020_375# trim_mask\[1\] 0.010728f
C9215 net81 FILLER_0_12_236/a_572_375# 0.021025f
C9216 FILLER_0_22_177/a_932_472# vss -0.001894f
C9217 FILLER_0_22_177/a_1380_472# vdd 0.007188f
C9218 _099_ mask\[2\] 0.776725f
C9219 net20 FILLER_0_12_220/a_932_472# 0.007397f
C9220 net68 net66 0.81104f
C9221 ctln[1] FILLER_0_1_266/a_124_375# 0.002958f
C9222 _159_ vdd 0.025131f
C9223 net32 _204_/a_67_603# 0.037639f
C9224 FILLER_0_21_125/a_484_472# _022_ 0.004649f
C9225 _426_/a_2560_156# net64 0.00801f
C9226 mask\[2\] FILLER_0_16_154/a_36_472# 0.312123f
C9227 _452_/a_448_472# net40 0.047031f
C9228 ctln[4] FILLER_0_1_204/a_124_375# 0.008283f
C9229 FILLER_0_4_107/a_932_472# _160_ 0.014254f
C9230 FILLER_0_4_213/a_484_472# vss 0.007857f
C9231 trimb[1] _452_/a_3129_107# 0.007229f
C9232 net52 FILLER_0_0_130/a_124_375# 0.004055f
C9233 _412_/a_2248_156# fanout58/a_36_160# 0.005856f
C9234 _132_ _131_ 0.444097f
C9235 _086_ _374_/a_36_68# 0.009872f
C9236 FILLER_0_14_99/a_36_472# FILLER_0_14_107/a_36_472# 0.002296f
C9237 _418_/a_796_472# _007_ 0.012286f
C9238 FILLER_0_17_72/a_2364_375# _131_ 0.006037f
C9239 output38/a_224_472# output41/a_224_472# 0.00607f
C9240 trim_val\[4\] _241_/a_224_472# 0.003005f
C9241 net55 FILLER_0_13_72/a_572_375# 0.005919f
C9242 fanout51/a_36_113# net55 0.010147f
C9243 net38 net67 1.762405f
C9244 _136_ _451_/a_1697_156# 0.001053f
C9245 _154_ vdd 0.639978f
C9246 FILLER_0_17_72/a_2724_472# net14 0.007133f
C9247 _449_/a_2248_156# vss 0.008071f
C9248 _449_/a_2665_112# vdd 0.012848f
C9249 FILLER_0_7_72/a_1828_472# net52 0.00159f
C9250 net26 _423_/a_448_472# 0.011612f
C9251 FILLER_0_20_87/a_124_375# net71 0.003629f
C9252 net53 FILLER_0_14_123/a_36_472# 0.062713f
C9253 net27 FILLER_0_10_256/a_36_472# 0.008331f
C9254 net74 _135_ 0.002261f
C9255 FILLER_0_16_57/a_36_472# cal_count\[2\] 0.001952f
C9256 sample net5 0.359975f
C9257 mask\[0\] FILLER_0_15_212/a_572_375# 0.001158f
C9258 _443_/a_1456_156# net23 0.001009f
C9259 fanout75/a_36_113# _122_ 0.001035f
C9260 _131_ _427_/a_36_151# 0.0012f
C9261 net4 _084_ 0.029194f
C9262 _277_/a_36_160# net31 0.053915f
C9263 FILLER_0_3_142/a_124_375# vdd 0.00167f
C9264 _028_ FILLER_0_6_90/a_36_472# 0.013106f
C9265 _059_ FILLER_0_8_156/a_36_472# 0.18373f
C9266 FILLER_0_18_177/a_1916_375# FILLER_0_19_195/a_36_472# 0.001684f
C9267 net27 net64 1.364577f
C9268 net54 _140_ 1.37516f
C9269 _149_ _437_/a_2560_156# 0.008064f
C9270 FILLER_0_17_38/a_36_472# _452_/a_36_151# 0.096503f
C9271 _141_ FILLER_0_17_161/a_124_375# 0.040332f
C9272 _070_ _152_ 0.114651f
C9273 _133_ _081_ 0.002847f
C9274 _431_/a_36_151# _136_ 0.03371f
C9275 net41 cal_count\[2\] 0.079279f
C9276 result[9] FILLER_0_14_263/a_124_375# 0.003706f
C9277 result[9] _010_ 0.121471f
C9278 _442_/a_448_472# vdd 0.006758f
C9279 _442_/a_36_151# vss 0.021278f
C9280 _123_ FILLER_0_6_231/a_484_472# 0.001396f
C9281 net34 _435_/a_1308_423# 0.008652f
C9282 output34/a_224_472# _421_/a_2248_156# 0.001144f
C9283 net38 _445_/a_448_472# 0.023336f
C9284 net15 FILLER_0_6_47/a_2364_375# 0.022624f
C9285 _176_ FILLER_0_15_72/a_36_472# 0.002101f
C9286 net50 _444_/a_2560_156# 0.001479f
C9287 _178_ _402_/a_2172_497# 0.003871f
C9288 net25 _423_/a_2665_112# 0.007096f
C9289 _086_ _133_ 0.035637f
C9290 FILLER_0_8_107/a_124_375# _131_ 0.001624f
C9291 _114_ _060_ 0.003352f
C9292 net47 _450_/a_1353_112# 0.018879f
C9293 net68 FILLER_0_3_54/a_124_375# 0.022559f
C9294 _126_ _172_ 0.017618f
C9295 ctlp[1] vdd 0.942436f
C9296 _305_/a_36_159# vss 0.003366f
C9297 _128_ _315_/a_1657_68# 0.0013f
C9298 FILLER_0_4_152/a_36_472# trim_mask\[4\] 0.011746f
C9299 FILLER_0_21_142/a_572_375# vss 0.097474f
C9300 _340_/a_36_160# mask\[6\] 0.010151f
C9301 FILLER_0_19_47/a_572_375# _013_ 0.012993f
C9302 _115_ FILLER_0_10_107/a_124_375# 0.011098f
C9303 FILLER_0_14_181/a_124_375# _095_ 0.005538f
C9304 ctln[3] net58 0.00479f
C9305 FILLER_0_19_155/a_572_375# vss 0.004538f
C9306 FILLER_0_4_152/a_36_472# net47 0.007541f
C9307 FILLER_0_13_206/a_36_472# vss 0.003985f
C9308 FILLER_0_18_2/a_2364_375# trimb[1] 0.001523f
C9309 net23 FILLER_0_16_154/a_124_375# 0.002689f
C9310 fanout82/a_36_113# calibrate 0.004982f
C9311 FILLER_0_5_117/a_124_375# _153_ 0.079379f
C9312 net41 FILLER_0_19_28/a_484_472# 0.047447f
C9313 _345_/a_36_160# net71 0.002396f
C9314 ctlp[7] _436_/a_36_151# 0.002655f
C9315 _053_ FILLER_0_6_90/a_124_375# 0.003061f
C9316 net20 ctlp[1] 0.024556f
C9317 net67 _067_ 0.151887f
C9318 _072_ _250_/a_36_68# 0.007337f
C9319 FILLER_0_3_221/a_36_472# vss 0.046345f
C9320 FILLER_0_3_221/a_484_472# vdd 0.002974f
C9321 _401_/a_36_68# FILLER_0_15_59/a_36_472# 0.019798f
C9322 _436_/a_1204_472# vdd 0.003143f
C9323 FILLER_0_11_124/a_124_375# _118_ 0.030768f
C9324 _423_/a_2560_156# _012_ 0.004165f
C9325 mask\[7\] _208_/a_36_160# 0.105845f
C9326 _432_/a_2248_156# _091_ 0.007123f
C9327 _115_ FILLER_0_9_142/a_124_375# 0.010167f
C9328 ctln[8] net50 0.0032f
C9329 _098_ _113_ 0.001472f
C9330 _439_/a_1000_472# vss 0.032923f
C9331 FILLER_0_22_128/a_36_472# _433_/a_36_151# 0.001653f
C9332 net62 _429_/a_2665_112# 0.02887f
C9333 _087_ vss 0.09895f
C9334 _079_ vdd 0.476075f
C9335 trim[4] net39 0.004535f
C9336 result[9] FILLER_0_23_282/a_36_472# 0.001324f
C9337 net15 _424_/a_2665_112# 0.046592f
C9338 FILLER_0_16_107/a_36_472# _040_ 0.015026f
C9339 output29/a_224_472# net29 0.038602f
C9340 _445_/a_448_472# net66 0.010949f
C9341 FILLER_0_8_24/a_484_472# FILLER_0_8_37/a_36_472# 0.001963f
C9342 _053_ _042_ 0.00242f
C9343 net19 FILLER_0_23_274/a_124_375# 0.01233f
C9344 FILLER_0_24_96/a_124_375# output25/a_224_472# 0.002633f
C9345 _096_ vss 0.126096f
C9346 net53 _136_ 0.099584f
C9347 net23 _043_ 0.042095f
C9348 _076_ _121_ 0.013717f
C9349 _104_ net61 1.149805f
C9350 net20 _079_ 0.177911f
C9351 mask\[3\] _275_/a_224_472# 0.002528f
C9352 FILLER_0_5_109/a_36_472# _154_ 0.070958f
C9353 FILLER_0_14_99/a_36_472# vss 0.003598f
C9354 _008_ _419_/a_448_472# 0.01758f
C9355 mask\[3\] FILLER_0_16_154/a_1020_375# 0.001996f
C9356 _081_ FILLER_0_5_164/a_36_472# 0.001603f
C9357 _114_ _116_ 0.038641f
C9358 net57 _280_/a_224_472# 0.001032f
C9359 FILLER_0_13_65/a_124_375# _067_ 0.001283f
C9360 net50 FILLER_0_6_90/a_484_472# 0.012286f
C9361 net44 FILLER_0_12_2/a_572_375# 0.041552f
C9362 _443_/a_36_151# _170_ 0.014771f
C9363 FILLER_0_5_128/a_484_472# _160_ 0.003335f
C9364 _077_ FILLER_0_9_72/a_1020_375# 0.008103f
C9365 FILLER_0_12_2/a_36_472# vss 0.003757f
C9366 _177_ vdd 0.111636f
C9367 net53 FILLER_0_13_142/a_124_375# 0.001599f
C9368 mask\[0\] FILLER_0_12_220/a_1468_375# 0.001484f
C9369 _074_ _312_/a_672_472# 0.005399f
C9370 _161_ calibrate 0.044443f
C9371 FILLER_0_10_37/a_124_375# vss 0.006228f
C9372 FILLER_0_10_37/a_36_472# vdd 0.141896f
C9373 result[4] net18 0.048179f
C9374 net82 net69 0.005307f
C9375 _077_ _128_ 0.005311f
C9376 FILLER_0_24_274/a_124_375# vdd 0.012632f
C9377 _091_ FILLER_0_17_218/a_36_472# 0.066133f
C9378 net18 net59 0.695067f
C9379 _448_/a_448_472# _037_ 0.044085f
C9380 _120_ FILLER_0_10_107/a_572_375# 0.002214f
C9381 net63 FILLER_0_18_177/a_124_375# 0.001937f
C9382 FILLER_0_7_72/a_2364_375# _077_ 0.002969f
C9383 net28 _045_ 0.05144f
C9384 net41 _043_ 0.03188f
C9385 FILLER_0_22_128/a_572_375# vdd 0.001473f
C9386 trimb[1] vss 0.048527f
C9387 _077_ _453_/a_1000_472# 0.033726f
C9388 _348_/a_49_472# mask\[6\] 0.005525f
C9389 output32/a_224_472# _010_ 0.001508f
C9390 _053_ FILLER_0_5_212/a_124_375# 0.048501f
C9391 _129_ calibrate 0.04134f
C9392 _301_/a_36_472# mask\[8\] 0.016751f
C9393 _161_ net21 0.011799f
C9394 _019_ vdd 0.015401f
C9395 _236_/a_36_160# _444_/a_36_151# 0.034413f
C9396 _069_ FILLER_0_15_212/a_36_472# 0.046864f
C9397 _163_ _160_ 0.120564f
C9398 _343_/a_49_472# _093_ 0.001926f
C9399 net20 FILLER_0_24_274/a_124_375# 0.002751f
C9400 trimb[1] FILLER_0_20_15/a_932_472# 0.001069f
C9401 _431_/a_36_151# net53 0.001579f
C9402 cal_itt\[1\] vdd 0.410279f
C9403 _114_ _118_ 0.074399f
C9404 output7/a_224_472# ctln[0] 0.081823f
C9405 net69 FILLER_0_3_78/a_484_472# 0.002068f
C9406 _088_ FILLER_0_3_172/a_2364_375# 0.002377f
C9407 FILLER_0_9_28/a_124_375# net42 0.007403f
C9408 FILLER_0_9_142/a_36_472# _120_ 0.035902f
C9409 FILLER_0_18_139/a_1468_375# net23 0.04546f
C9410 net60 _418_/a_2560_156# 0.020147f
C9411 _031_ FILLER_0_2_127/a_124_375# 0.013811f
C9412 FILLER_0_19_125/a_124_375# _132_ 0.009167f
C9413 _119_ _372_/a_170_472# 0.003159f
C9414 _410_/a_36_68# vss 0.02717f
C9415 FILLER_0_21_206/a_124_375# _434_/a_2665_112# 0.002259f
C9416 _028_ FILLER_0_7_104/a_484_472# 0.00499f
C9417 _140_ _350_/a_49_472# 0.028997f
C9418 _013_ net55 0.239055f
C9419 FILLER_0_15_212/a_124_375# FILLER_0_15_205/a_124_375# 0.004426f
C9420 FILLER_0_0_130/a_36_472# net13 0.002757f
C9421 _070_ _113_ 0.01052f
C9422 net79 _248_/a_36_68# 0.018243f
C9423 net82 _152_ 0.001896f
C9424 _098_ net71 1.076897f
C9425 _397_/a_36_472# FILLER_0_17_72/a_1468_375# 0.001295f
C9426 _113_ FILLER_0_15_180/a_124_375# 0.001512f
C9427 _065_ _036_ 0.031728f
C9428 net41 net68 0.009755f
C9429 net54 FILLER_0_21_150/a_36_472# 0.005439f
C9430 _412_/a_2248_156# net18 0.05155f
C9431 _128_ _120_ 0.053476f
C9432 _144_ FILLER_0_21_125/a_484_472# 0.001616f
C9433 net62 _417_/a_2560_156# 0.003361f
C9434 _411_/a_36_151# net75 0.033786f
C9435 result[6] net62 0.005382f
C9436 _412_/a_796_472# net58 0.001182f
C9437 ctln[6] FILLER_0_0_130/a_124_375# 0.026786f
C9438 _420_/a_36_151# FILLER_0_23_274/a_124_375# 0.059049f
C9439 FILLER_0_9_282/a_36_472# vss 0.002224f
C9440 _308_/a_124_24# _070_ 0.001465f
C9441 FILLER_0_6_47/a_1828_472# vdd 0.002735f
C9442 FILLER_0_6_47/a_1380_472# vss 0.001431f
C9443 _429_/a_448_472# net21 0.014792f
C9444 cal_itt\[3\] _062_ 0.009718f
C9445 net35 FILLER_0_22_107/a_484_472# 0.008026f
C9446 net64 net18 1.557441f
C9447 _193_/a_36_160# FILLER_0_13_290/a_36_472# 0.004828f
C9448 FILLER_0_15_142/a_484_472# net53 0.044267f
C9449 _233_/a_36_160# net49 0.035342f
C9450 _053_ FILLER_0_7_104/a_1468_375# 0.001492f
C9451 result[4] _417_/a_448_472# 0.003485f
C9452 _430_/a_2665_112# FILLER_0_15_212/a_1380_472# 0.021761f
C9453 net75 _316_/a_124_24# 0.003078f
C9454 _322_/a_1152_472# _118_ 0.001235f
C9455 _322_/a_124_24# _124_ 0.041337f
C9456 FILLER_0_22_177/a_124_375# _434_/a_1308_423# 0.001064f
C9457 FILLER_0_13_212/a_36_472# vss 0.005259f
C9458 net26 FILLER_0_21_28/a_1468_375# 0.041169f
C9459 _131_ FILLER_0_14_107/a_1380_472# 0.01797f
C9460 ctlp[1] _420_/a_1308_423# 0.001418f
C9461 FILLER_0_20_107/a_36_472# net14 0.002543f
C9462 FILLER_0_5_109/a_484_472# vdd 0.007355f
C9463 _421_/a_2665_112# vss 0.002792f
C9464 _421_/a_2560_156# vdd 0.001862f
C9465 cal_count\[3\] net40 0.080767f
C9466 _446_/a_1204_472# net17 0.003628f
C9467 net9 cal_itt\[1\] 0.028339f
C9468 _086_ _121_ 0.049499f
C9469 net24 net14 0.172253f
C9470 net79 _005_ 1.006306f
C9471 net20 FILLER_0_13_212/a_484_472# 0.001273f
C9472 vdd FILLER_0_5_148/a_124_375# -0.011369f
C9473 _075_ _056_ 0.001957f
C9474 fanout50/a_36_160# net50 0.052685f
C9475 FILLER_0_8_107/a_36_472# _133_ 0.00589f
C9476 FILLER_0_19_187/a_484_472# vdd 0.011023f
C9477 FILLER_0_19_187/a_36_472# vss 0.001951f
C9478 _170_ net59 0.002301f
C9479 net41 net67 0.03408f
C9480 net73 FILLER_0_18_107/a_2364_375# 0.015484f
C9481 FILLER_0_5_117/a_36_472# vss 0.001215f
C9482 _429_/a_1000_472# net22 0.007429f
C9483 _429_/a_796_472# _018_ 0.002291f
C9484 net7 output40/a_224_472# 0.006944f
C9485 FILLER_0_2_111/a_36_472# vdd 0.033758f
C9486 FILLER_0_2_111/a_1468_375# vss 0.055168f
C9487 _431_/a_2665_112# FILLER_0_17_142/a_572_375# 0.001092f
C9488 FILLER_0_4_91/a_36_472# _160_ 0.007864f
C9489 net15 _394_/a_56_524# 0.006099f
C9490 net52 net49 0.092082f
C9491 _074_ net59 0.030221f
C9492 trimb[4] cal_count\[2\] 0.146942f
C9493 _443_/a_36_151# _081_ 0.001923f
C9494 _092_ net22 0.010937f
C9495 ctlp[4] vss 0.102044f
C9496 _440_/a_796_472# vss 0.001285f
C9497 net18 _418_/a_1308_423# 0.015651f
C9498 net18 _006_ 0.082256f
C9499 _077_ FILLER_0_9_60/a_484_472# 0.024249f
C9500 trim[4] clkc 0.005f
C9501 _076_ net59 0.005449f
C9502 _313_/a_67_603# vss 0.016047f
C9503 net82 _443_/a_1308_423# 0.006706f
C9504 _449_/a_36_151# net74 0.032989f
C9505 output47/a_224_472# net3 0.002186f
C9506 trimb[4] input3/a_36_113# 0.001221f
C9507 net41 _445_/a_448_472# 0.002211f
C9508 _017_ FILLER_0_14_107/a_572_375# 0.003679f
C9509 FILLER_0_21_286/a_36_472# net18 0.18097f
C9510 net70 FILLER_0_14_107/a_1468_375# 0.007955f
C9511 fanout79/a_36_160# vdd 0.099877f
C9512 net41 FILLER_0_21_28/a_484_472# 0.060027f
C9513 net44 FILLER_0_20_2/a_572_375# 0.002597f
C9514 mask\[4\] FILLER_0_20_193/a_484_472# 0.001215f
C9515 _088_ net76 0.214494f
C9516 _056_ calibrate 0.00931f
C9517 _050_ FILLER_0_22_128/a_36_472# 0.001098f
C9518 _103_ net18 0.11279f
C9519 FILLER_0_20_2/a_484_472# vdd 0.001049f
C9520 FILLER_0_17_200/a_124_375# net22 0.003602f
C9521 FILLER_0_5_54/a_932_472# trim_mask\[1\] 0.016187f
C9522 fanout62/a_36_160# vss 0.01343f
C9523 _430_/a_36_151# FILLER_0_18_177/a_3172_472# 0.001512f
C9524 _013_ _216_/a_67_603# 0.006454f
C9525 _075_ _068_ 0.006297f
C9526 _294_/a_224_472# vss 0.001022f
C9527 _438_/a_448_472# vdd 0.009409f
C9528 _438_/a_36_151# vss 0.014203f
C9529 ctlp[1] _419_/a_796_472# 0.001178f
C9530 _322_/a_848_380# _062_ 0.001872f
C9531 net34 net61 0.037731f
C9532 FILLER_0_8_127/a_124_375# net74 0.026604f
C9533 ctln[5] FILLER_0_1_192/a_124_375# 0.001391f
C9534 _451_/a_2225_156# vdd 0.012404f
C9535 _451_/a_3129_107# vss 0.01f
C9536 _000_ _411_/a_1308_423# 0.004012f
C9537 output19/a_224_472# _295_/a_36_472# 0.003896f
C9538 _291_/a_36_160# _093_ 0.017281f
C9539 _056_ net21 0.484506f
C9540 _111_ _013_ 0.024203f
C9541 FILLER_0_5_198/a_484_472# net37 0.009858f
C9542 net61 net60 0.059237f
C9543 _063_ _164_ 0.326812f
C9544 net57 _043_ 1.955053f
C9545 _074_ _122_ 0.300373f
C9546 _130_ _118_ 0.053869f
C9547 FILLER_0_18_53/a_36_472# FILLER_0_18_37/a_1380_472# 0.013276f
C9548 trim_val\[1\] FILLER_0_6_37/a_124_375# 0.007292f
C9549 ctlp[4] _107_ 0.080312f
C9550 _370_/a_848_380# FILLER_0_5_136/a_36_472# 0.001177f
C9551 _086_ _132_ 0.014693f
C9552 _074_ FILLER_0_7_233/a_124_375# 0.003081f
C9553 _415_/a_36_151# _416_/a_1308_423# 0.00119f
C9554 _430_/a_36_151# fanout80/a_36_113# 0.018169f
C9555 cal_itt\[2\] _253_/a_36_68# 0.010756f
C9556 _088_ FILLER_0_5_198/a_124_375# 0.001374f
C9557 _079_ FILLER_0_5_198/a_572_375# 0.011369f
C9558 FILLER_0_19_28/a_124_375# net40 0.047489f
C9559 _219_/a_36_160# _058_ 0.014194f
C9560 FILLER_0_18_2/a_1916_375# output44/a_224_472# 0.032639f
C9561 net68 FILLER_0_5_54/a_124_375# 0.018458f
C9562 mask\[4\] FILLER_0_18_177/a_2364_375# 0.01602f
C9563 FILLER_0_5_128/a_484_472# _133_ 0.037369f
C9564 _126_ FILLER_0_13_206/a_124_375# 0.002746f
C9565 _068_ calibrate 0.110297f
C9566 _076_ _122_ 0.097035f
C9567 _042_ cal_count\[0\] 0.006265f
C9568 FILLER_0_4_197/a_1468_375# net22 0.009108f
C9569 _033_ trim_mask\[1\] 0.001251f
C9570 net5 net8 0.001288f
C9571 _411_/a_2248_156# net8 0.06032f
C9572 trim[0] FILLER_0_3_2/a_124_375# 0.020708f
C9573 FILLER_0_9_28/a_2724_472# net68 0.010755f
C9574 FILLER_0_20_177/a_124_375# mask\[6\] 0.001158f
C9575 net36 FILLER_0_15_235/a_124_375# 0.007232f
C9576 _073_ _083_ 0.097365f
C9577 FILLER_0_6_177/a_124_375# vdd 0.017329f
C9578 net1 en 0.068102f
C9579 FILLER_0_4_152/a_124_375# trim_mask\[4\] 0.01182f
C9580 net50 net14 0.192231f
C9581 _430_/a_1308_423# _429_/a_36_151# 0.001722f
C9582 _430_/a_1000_472# net63 0.016386f
C9583 _076_ _227_/a_36_160# 0.004997f
C9584 _417_/a_448_472# _006_ 0.068545f
C9585 FILLER_0_7_104/a_572_375# _131_ 0.003031f
C9586 _068_ net21 0.030836f
C9587 FILLER_0_4_152/a_124_375# net47 0.009228f
C9588 FILLER_0_18_171/a_36_472# mask\[4\] 0.01222f
C9589 _052_ FILLER_0_21_28/a_2812_375# 0.002388f
C9590 _077_ FILLER_0_9_223/a_36_472# 0.005511f
C9591 _133_ _163_ 0.034905f
C9592 net32 net30 0.004658f
C9593 FILLER_0_18_37/a_484_472# vdd 0.008381f
C9594 FILLER_0_18_37/a_36_472# vss 0.003026f
C9595 _086_ _321_/a_170_472# 0.046783f
C9596 _093_ FILLER_0_16_89/a_1468_375# 0.003988f
C9597 net50 _164_ 0.080818f
C9598 net39 FILLER_0_8_2/a_124_375# 0.008405f
C9599 trim[4] net47 0.009333f
C9600 _174_ _131_ 0.002314f
C9601 _000_ _253_/a_244_68# 0.001243f
C9602 _372_/a_170_472# _385_/a_36_68# 0.009691f
C9603 _317_/a_36_113# FILLER_0_7_233/a_36_472# 0.003531f
C9604 result[9] vss 0.348416f
C9605 _092_ vdd 0.140213f
C9606 _164_ _382_/a_224_472# 0.011658f
C9607 net16 cal_count\[1\] 0.007291f
C9608 FILLER_0_9_72/a_36_472# _453_/a_2248_156# 0.013656f
C9609 input1/a_36_113# net1 0.003795f
C9610 net79 _416_/a_448_472# 0.078357f
C9611 FILLER_0_9_28/a_36_472# net51 0.002082f
C9612 _176_ cal_count\[1\] 0.297763f
C9613 _037_ net12 0.007817f
C9614 net62 _416_/a_1308_423# 0.002665f
C9615 fanout82/a_36_113# output48/a_224_472# 0.009784f
C9616 _256_/a_36_68# _056_ 0.008305f
C9617 _096_ _095_ 0.086147f
C9618 net31 ctlp[1] 0.050993f
C9619 _093_ FILLER_0_17_72/a_2276_472# 0.017114f
C9620 _081_ net59 0.185504f
C9621 FILLER_0_7_72/a_3172_472# net14 0.046751f
C9622 net70 vdd 0.858299f
C9623 FILLER_0_14_99/a_36_472# _095_ 0.011772f
C9624 net20 _092_ 0.001458f
C9625 net26 _424_/a_36_151# 0.062638f
C9626 FILLER_0_7_195/a_36_472# _072_ 0.008357f
C9627 _021_ _432_/a_448_472# 0.032563f
C9628 _431_/a_1204_472# _020_ 0.002176f
C9629 FILLER_0_17_200/a_124_375# vdd -0.010938f
C9630 FILLER_0_10_247/a_124_375# vdd 0.040502f
C9631 _004_ _005_ 0.004158f
C9632 _287_/a_36_472# net30 0.005402f
C9633 output44/a_224_472# vdd 0.043902f
C9634 FILLER_0_7_72/a_1916_375# _053_ 0.013335f
C9635 FILLER_0_9_105/a_124_375# FILLER_0_10_107/a_36_472# 0.001543f
C9636 vdd _381_/a_36_472# 0.014305f
C9637 _122_ FILLER_0_5_164/a_484_472# 0.002997f
C9638 _430_/a_2248_156# _092_ 0.003124f
C9639 vdd FILLER_0_22_107/a_484_472# 0.035591f
C9640 vss FILLER_0_22_107/a_36_472# 0.001514f
C9641 FILLER_0_22_86/a_124_375# net71 0.002239f
C9642 output44/a_224_472# FILLER_0_20_15/a_484_472# 0.0323f
C9643 _104_ FILLER_0_23_274/a_36_472# 0.001642f
C9644 _132_ FILLER_0_15_116/a_484_472# 0.010148f
C9645 net36 _280_/a_224_472# 0.001012f
C9646 FILLER_0_5_72/a_572_375# _164_ 0.005919f
C9647 FILLER_0_10_107/a_124_375# vdd 0.045066f
C9648 net65 net59 0.790496f
C9649 FILLER_0_12_50/a_124_375# _067_ 0.011869f
C9650 FILLER_0_16_255/a_36_472# _045_ 0.001653f
C9651 FILLER_0_15_228/a_124_375# vdd 0.013701f
C9652 _187_ _043_ 0.011995f
C9653 trim_mask\[0\] FILLER_0_10_94/a_572_375# 0.003359f
C9654 net55 FILLER_0_11_78/a_572_375# 0.002321f
C9655 _256_/a_36_68# _068_ 0.029112f
C9656 ctln[6] net52 0.1064f
C9657 _413_/a_2665_112# ctln[4] 0.001394f
C9658 FILLER_0_6_239/a_124_375# _316_/a_124_24# 0.003524f
C9659 net16 FILLER_0_17_38/a_36_472# 0.014381f
C9660 FILLER_0_5_164/a_36_472# _163_ 0.001777f
C9661 input4/a_36_68# vss 0.058179f
C9662 fanout66/a_36_113# vss 0.014789f
C9663 _444_/a_1204_472# net17 0.021952f
C9664 net16 _392_/a_36_68# 0.002191f
C9665 FILLER_0_2_93/a_36_472# net69 0.010977f
C9666 _111_ net71 0.002668f
C9667 net20 FILLER_0_15_228/a_124_375# 0.047331f
C9668 net15 FILLER_0_5_54/a_1380_472# 0.047774f
C9669 _155_ _029_ 0.174512f
C9670 _425_/a_796_472# _122_ 0.001701f
C9671 _425_/a_36_151# _123_ 0.006319f
C9672 _425_/a_1000_472# calibrate 0.027245f
C9673 FILLER_0_9_142/a_124_375# vdd 0.015952f
C9674 _081_ _122_ 2.557248f
C9675 _152_ calibrate 0.020369f
C9676 _072_ _311_/a_3220_473# 0.001995f
C9677 _119_ FILLER_0_5_117/a_36_472# 0.002628f
C9678 FILLER_0_4_197/a_1468_375# vdd 0.019672f
C9679 _424_/a_2665_112# _012_ 0.01024f
C9680 net38 FILLER_0_15_10/a_124_375# 0.047331f
C9681 ctln[3] _411_/a_1204_472# 0.00185f
C9682 _033_ _444_/a_2665_112# 0.004024f
C9683 FILLER_0_12_136/a_484_472# net23 0.002172f
C9684 cal_itt\[2\] FILLER_0_3_221/a_484_472# 0.016997f
C9685 net80 _434_/a_1204_472# 0.003997f
C9686 _024_ _435_/a_1308_423# 0.002661f
C9687 _417_/a_1000_472# vss 0.001822f
C9688 FILLER_0_9_72/a_572_375# vdd -0.014642f
C9689 FILLER_0_9_72/a_124_375# vss 0.047932f
C9690 _306_/a_36_68# _085_ 0.00755f
C9691 FILLER_0_20_98/a_36_472# vss 0.00206f
C9692 _086_ _122_ 0.033097f
C9693 trim_mask\[2\] net69 0.051795f
C9694 _412_/a_2248_156# net65 0.039861f
C9695 _304_/a_224_472# mask\[9\] 0.003125f
C9696 _155_ FILLER_0_8_107/a_36_472# 0.002068f
C9697 net73 FILLER_0_19_111/a_572_375# 0.04458f
C9698 _324_/a_224_472# net74 0.001704f
C9699 _093_ FILLER_0_18_139/a_572_375# 0.008393f
C9700 FILLER_0_10_78/a_1380_472# _176_ 0.009351f
C9701 _121_ _314_/a_224_472# 0.00323f
C9702 cal_itt\[2\] _079_ 0.017071f
C9703 net18 _416_/a_1288_156# 0.001147f
C9704 output32/a_224_472# vss -0.003023f
C9705 _081_ _169_ 0.260462f
C9706 _119_ _313_/a_67_603# 0.015457f
C9707 _061_ vss 0.046487f
C9708 FILLER_0_5_72/a_1468_375# net47 0.005049f
C9709 FILLER_0_21_28/a_572_375# net17 0.001455f
C9710 mask\[8\] FILLER_0_22_86/a_1380_472# 0.012151f
C9711 net35 FILLER_0_22_86/a_932_472# 0.007806f
C9712 FILLER_0_13_290/a_36_472# _416_/a_36_151# 0.001723f
C9713 _453_/a_1308_423# vss 0.003012f
C9714 FILLER_0_13_212/a_932_472# _043_ 0.014431f
C9715 _311_/a_254_473# vdd 0.001207f
C9716 cal_count\[2\] FILLER_0_15_2/a_124_375# 0.033559f
C9717 _323_/a_36_113# _426_/a_2248_156# 0.001661f
C9718 _015_ _426_/a_1308_423# 0.029444f
C9719 _077_ _176_ 0.00497f
C9720 _053_ _372_/a_170_472# 0.05895f
C9721 _064_ net17 0.108825f
C9722 FILLER_0_16_89/a_1468_375# _136_ 0.005791f
C9723 _138_ net21 0.003242f
C9724 ctlp[5] vss 0.032166f
C9725 ctln[1] FILLER_0_3_221/a_1020_375# 0.001554f
C9726 net65 net64 0.119915f
C9727 _001_ vss 0.004381f
C9728 ctlp[6] FILLER_0_24_130/a_36_472# 0.005932f
C9729 _000_ FILLER_0_3_221/a_932_472# 0.008308f
C9730 FILLER_0_18_2/a_932_472# net55 0.012117f
C9731 _337_/a_49_472# _137_ 0.046633f
C9732 ctlp[1] net77 0.716304f
C9733 net56 mask\[2\] 0.090254f
C9734 _098_ _437_/a_1000_472# 0.007963f
C9735 _132_ _145_ 0.010994f
C9736 FILLER_0_11_142/a_124_375# FILLER_0_11_135/a_124_375# 0.004426f
C9737 net54 FILLER_0_22_128/a_484_472# 0.055436f
C9738 mask\[5\] FILLER_0_18_177/a_572_375# 0.002653f
C9739 FILLER_0_17_72/a_2276_472# _136_ 0.055635f
C9740 net17 net42 0.056318f
C9741 _131_ FILLER_0_16_115/a_124_375# 0.016715f
C9742 vss _433_/a_36_151# 0.00618f
C9743 vdd _433_/a_448_472# 0.003821f
C9744 mask\[0\] _429_/a_448_472# 0.061449f
C9745 _448_/a_1000_472# net59 0.007647f
C9746 _093_ FILLER_0_18_76/a_36_472# 0.129892f
C9747 _101_ vss 0.05721f
C9748 _251_/a_244_472# net4 0.005273f
C9749 FILLER_0_11_101/a_484_472# vss 0.003923f
C9750 FILLER_0_3_172/a_124_375# net22 0.01308f
C9751 _128_ _125_ 0.017316f
C9752 _027_ _438_/a_36_151# 0.010763f
C9753 _150_ _438_/a_1308_423# 0.001472f
C9754 FILLER_0_20_98/a_124_375# _437_/a_36_151# 0.059049f
C9755 FILLER_0_18_100/a_36_472# mask\[9\] 0.005719f
C9756 result[6] fanout77/a_36_113# 0.001469f
C9757 FILLER_0_18_107/a_484_472# FILLER_0_17_104/a_932_472# 0.026657f
C9758 net63 fanout63/a_36_160# 0.011149f
C9759 FILLER_0_13_212/a_1468_375# FILLER_0_12_220/a_572_375# 0.05841f
C9760 _414_/a_448_472# cal_itt\[3\] 0.109704f
C9761 _052_ _424_/a_796_472# 0.002115f
C9762 FILLER_0_16_57/a_124_375# _131_ 0.012982f
C9763 _072_ vss 0.439154f
C9764 mask\[1\] FILLER_0_15_180/a_484_472# 0.003594f
C9765 _399_/a_224_472# _179_ 0.002288f
C9766 FILLER_0_19_125/a_36_472# net73 0.004017f
C9767 cal_itt\[2\] cal_itt\[1\] 0.057194f
C9768 FILLER_0_11_142/a_572_375# _076_ 0.031784f
C9769 _395_/a_36_488# _085_ 0.020572f
C9770 output27/a_224_472# result[0] 0.031252f
C9771 net16 _120_ 0.009918f
C9772 FILLER_0_4_197/a_1380_472# _081_ 0.001345f
C9773 FILLER_0_7_162/a_124_375# _074_ 0.007213f
C9774 net76 FILLER_0_6_177/a_572_375# 0.073022f
C9775 _132_ _318_/a_224_472# 0.001097f
C9776 _176_ _120_ 0.169846f
C9777 _176_ _038_ 0.039948f
C9778 net23 FILLER_0_21_150/a_124_375# 0.045928f
C9779 net19 _417_/a_2665_112# 0.042961f
C9780 FILLER_0_7_104/a_1020_375# _133_ 0.008772f
C9781 FILLER_0_19_195/a_124_375# vss 0.020433f
C9782 FILLER_0_19_195/a_36_472# vdd 0.094409f
C9783 _126_ _390_/a_36_68# 0.044675f
C9784 _011_ _009_ 0.035129f
C9785 _014_ vss 0.034646f
C9786 _104_ _093_ 0.109158f
C9787 _077_ _257_/a_36_472# 0.019883f
C9788 net81 _425_/a_36_151# 0.014663f
C9789 _085_ FILLER_0_13_142/a_1468_375# 0.001153f
C9790 FILLER_0_5_206/a_124_375# _081_ 0.031751f
C9791 cal_count\[3\] FILLER_0_9_72/a_484_472# 0.004129f
C9792 FILLER_0_14_181/a_124_375# _098_ 0.005696f
C9793 vss FILLER_0_13_72/a_484_472# 0.008682f
C9794 _360_/a_36_160# FILLER_0_4_123/a_36_472# 0.001165f
C9795 _093_ FILLER_0_18_209/a_572_375# 0.064723f
C9796 output16/a_224_472# _447_/a_36_151# 0.200384f
C9797 _365_/a_36_68# vdd 0.004308f
C9798 FILLER_0_16_89/a_484_472# net36 0.003595f
C9799 fanout69/a_36_113# _160_ 0.005933f
C9800 _345_/a_36_160# FILLER_0_19_111/a_484_472# 0.007907f
C9801 net63 _432_/a_36_151# 0.001392f
C9802 _413_/a_36_151# FILLER_0_3_172/a_2724_472# 0.001723f
C9803 _308_/a_124_24# FILLER_0_10_94/a_36_472# 0.001811f
C9804 _429_/a_36_151# FILLER_0_15_212/a_572_375# 0.059049f
C9805 net65 FILLER_0_1_266/a_124_375# 0.002654f
C9806 _155_ _163_ 0.296236f
C9807 net41 net26 0.057852f
C9808 output31/a_224_472# result[9] 0.082001f
C9809 _432_/a_2248_156# vdd 0.02369f
C9810 _150_ net36 0.108945f
C9811 FILLER_0_18_107/a_3172_472# FILLER_0_19_134/a_124_375# 0.001723f
C9812 _021_ _143_ 0.007778f
C9813 _097_ FILLER_0_15_180/a_36_472# 0.005242f
C9814 cal_count\[2\] _452_/a_36_151# 0.006982f
C9815 FILLER_0_17_38/a_36_472# _041_ 0.003805f
C9816 net74 FILLER_0_11_124/a_124_375# 0.047331f
C9817 FILLER_0_2_101/a_36_472# net14 0.051153f
C9818 _431_/a_2248_156# net36 0.001441f
C9819 _063_ _378_/a_224_472# 0.002323f
C9820 _343_/a_665_69# _141_ 0.002451f
C9821 _031_ vss 0.18315f
C9822 mask\[9\] _438_/a_2560_156# 0.008709f
C9823 net72 _424_/a_448_472# 0.011745f
C9824 _064_ _446_/a_1308_423# 0.001728f
C9825 output38/a_224_472# net17 0.04454f
C9826 net52 FILLER_0_5_54/a_1468_375# 0.003649f
C9827 _005_ net19 0.033451f
C9828 _074_ FILLER_0_5_181/a_36_472# 0.002385f
C9829 _015_ FILLER_0_8_239/a_36_472# 0.002627f
C9830 _320_/a_36_472# net22 0.005964f
C9831 FILLER_0_16_73/a_572_375# FILLER_0_17_72/a_572_375# 0.026339f
C9832 net52 _442_/a_1204_472# 0.005558f
C9833 _384_/a_224_472# _168_ 0.003461f
C9834 FILLER_0_18_177/a_1828_472# vss -0.001107f
C9835 FILLER_0_18_177/a_2276_472# vdd 0.005211f
C9836 output8/a_224_472# FILLER_0_3_221/a_1380_472# 0.001699f
C9837 _005_ _416_/a_796_472# 0.009162f
C9838 result[9] _419_/a_1000_472# 0.012469f
C9839 FILLER_0_2_101/a_124_375# trim_mask\[3\] 0.033692f
C9840 net38 _033_ 0.03598f
C9841 FILLER_0_14_81/a_36_472# _177_ 0.004294f
C9842 _441_/a_448_472# _168_ 0.033059f
C9843 _415_/a_2248_156# net58 0.001869f
C9844 net66 FILLER_0_5_54/a_932_472# 0.001419f
C9845 FILLER_0_9_60/a_36_472# vdd 0.08419f
C9846 FILLER_0_9_60/a_572_375# vss 0.022532f
C9847 net18 _419_/a_2665_112# 0.0371f
C9848 FILLER_0_13_212/a_124_375# FILLER_0_13_206/a_124_375# 0.005439f
C9849 mask\[3\] fanout53/a_36_160# 0.001205f
C9850 FILLER_0_16_73/a_484_472# _131_ 0.007761f
C9851 FILLER_0_18_2/a_3172_472# net40 0.046864f
C9852 FILLER_0_21_206/a_124_375# mask\[6\] 0.008881f
C9853 ctlp[1] _421_/a_448_472# 0.011026f
C9854 mask\[0\] _056_ 0.001878f
C9855 FILLER_0_17_104/a_484_472# net14 0.004272f
C9856 net69 _441_/a_2560_156# 0.002904f
C9857 _094_ vss 0.24519f
C9858 FILLER_0_17_218/a_572_375# vss 0.078608f
C9859 FILLER_0_17_218/a_36_472# vdd 0.084913f
C9860 FILLER_0_3_172/a_124_375# vdd 0.010886f
C9861 _425_/a_2665_112# vdd 0.012933f
C9862 _035_ _379_/a_36_472# 0.002226f
C9863 mask\[7\] FILLER_0_22_128/a_2276_472# 0.004398f
C9864 net63 FILLER_0_20_177/a_572_375# 0.00281f
C9865 _432_/a_36_151# FILLER_0_17_161/a_124_375# 0.035117f
C9866 _069_ _429_/a_1000_472# 0.029501f
C9867 _431_/a_2560_156# net73 0.001018f
C9868 _092_ _069_ 0.040267f
C9869 FILLER_0_14_181/a_124_375# FILLER_0_15_180/a_124_375# 0.026339f
C9870 net53 _427_/a_2560_156# 0.004594f
C9871 FILLER_0_22_128/a_36_472# _022_ 0.001541f
C9872 net28 fanout79/a_36_160# 0.036675f
C9873 _423_/a_36_151# FILLER_0_23_44/a_1020_375# 0.059049f
C9874 _350_/a_49_472# _049_ 0.025442f
C9875 _013_ FILLER_0_18_61/a_124_375# 0.016976f
C9876 _394_/a_718_524# FILLER_0_15_59/a_572_375# 0.001447f
C9877 _394_/a_56_524# FILLER_0_15_59/a_484_472# 0.001033f
C9878 _448_/a_2560_156# net22 0.00766f
C9879 _233_/a_36_160# net40 0.001875f
C9880 _274_/a_36_68# state\[0\] 0.001852f
C9881 FILLER_0_9_28/a_36_472# net47 0.006712f
C9882 _098_ FILLER_0_15_212/a_1468_375# 0.008327f
C9883 _429_/a_36_151# FILLER_0_15_205/a_124_375# 0.059049f
C9884 _428_/a_2248_156# net74 0.072805f
C9885 output7/a_224_472# trim[2] 0.008581f
C9886 net50 _439_/a_2665_112# 0.007973f
C9887 ctln[3] ctln[2] 0.012289f
C9888 FILLER_0_4_144/a_36_472# net23 0.016933f
C9889 _079_ FILLER_0_6_231/a_484_472# 0.008159f
C9890 _138_ mask\[1\] 0.085445f
C9891 _057_ net56 0.002158f
C9892 FILLER_0_4_144/a_484_472# trim_mask\[4\] 0.015778f
C9893 _331_/a_448_472# vdd 0.001343f
C9894 _086_ FILLER_0_11_142/a_572_375# 0.011726f
C9895 _098_ FILLER_0_16_154/a_1380_472# 0.00417f
C9896 ctln[0] output40/a_224_472# 0.017541f
C9897 FILLER_0_5_109/a_36_472# _365_/a_36_68# 0.07596f
C9898 _394_/a_56_524# net74 0.005616f
C9899 net54 FILLER_0_19_142/a_36_472# 0.07544f
C9900 mask\[3\] _098_ 0.026156f
C9901 _176_ _175_ 0.054439f
C9902 FILLER_0_4_144/a_484_472# net47 0.008338f
C9903 _119_ _061_ 0.132725f
C9904 _114_ net74 0.559239f
C9905 output46/a_224_472# FILLER_0_20_15/a_124_375# 0.029497f
C9906 _261_/a_36_160# vdd 0.0109f
C9907 _028_ FILLER_0_6_47/a_2276_472# 0.002066f
C9908 _086_ FILLER_0_7_104/a_572_375# 0.003137f
C9909 FILLER_0_11_101/a_36_472# FILLER_0_13_100/a_124_375# 0.001436f
C9910 _098_ _434_/a_448_472# 0.015893f
C9911 _238_/a_67_603# trim_val\[3\] 0.024283f
C9912 FILLER_0_21_133/a_124_375# _098_ 0.006462f
C9913 _093_ FILLER_0_17_142/a_484_472# 0.011974f
C9914 net48 _317_/a_36_113# 0.018494f
C9915 _412_/a_448_472# output37/a_224_472# 0.001155f
C9916 FILLER_0_7_72/a_2724_472# net50 0.007192f
C9917 net2 _425_/a_36_151# 0.012359f
C9918 _105_ _201_/a_67_603# 0.003335f
C9919 _411_/a_2665_112# cal_itt\[0\] 0.010667f
C9920 _412_/a_1000_472# net81 0.012828f
C9921 _394_/a_2215_68# _095_ 0.001134f
C9922 output31/a_224_472# output32/a_224_472# 0.00289f
C9923 FILLER_0_22_86/a_932_472# vdd 0.001826f
C9924 trim_val\[4\] _170_ 0.281942f
C9925 ctln[3] ctln[1] 0.926618f
C9926 _199_/a_36_160# vdd 0.036579f
C9927 mask\[4\] FILLER_0_19_171/a_36_472# 0.001776f
C9928 output45/a_224_472# vss 0.00543f
C9929 FILLER_0_22_128/a_3172_472# vss 0.006339f
C9930 FILLER_0_9_290/a_36_472# FILLER_0_9_282/a_484_472# 0.013276f
C9931 net35 _435_/a_448_472# 0.007865f
C9932 result[6] _419_/a_36_151# 0.001968f
C9933 output24/a_224_472# _050_ 0.061723f
C9934 net59 net11 0.016998f
C9935 net31 _092_ 0.04309f
C9936 net78 vss 0.167812f
C9937 net20 _199_/a_36_160# 0.05178f
C9938 _442_/a_2665_112# net14 0.011563f
C9939 _050_ vss 0.26237f
C9940 FILLER_0_24_63/a_36_472# ctlp[9] 0.012298f
C9941 net37 _160_ 0.003563f
C9942 _053_ FILLER_0_6_47/a_1380_472# 0.004472f
C9943 net80 _093_ 0.818824f
C9944 _320_/a_36_472# vdd 0.086964f
C9945 _445_/a_1204_472# _034_ 0.003057f
C9946 FILLER_0_0_198/a_124_375# net11 0.071885f
C9947 net15 _447_/a_448_472# 0.001766f
C9948 net49 net40 0.093233f
C9949 net52 FILLER_0_6_79/a_124_375# 0.010099f
C9950 net82 FILLER_0_3_172/a_1828_472# 0.004472f
C9951 FILLER_0_8_263/a_36_472# vss 0.001089f
C9952 _414_/a_1456_156# cal_itt\[3\] 0.001134f
C9953 _119_ _072_ 0.189217f
C9954 net34 FILLER_0_22_128/a_1916_375# 0.04185f
C9955 _093_ FILLER_0_18_107/a_2276_472# 0.001996f
C9956 _072_ _071_ 0.296543f
C9957 vss FILLER_0_14_235/a_572_375# 0.017196f
C9958 _442_/a_2248_156# trim_mask\[3\] 0.003039f
C9959 net27 FILLER_0_9_282/a_124_375# 0.003572f
C9960 FILLER_0_3_172/a_932_472# net65 0.002604f
C9961 ctln[3] FILLER_0_0_266/a_36_472# 0.012298f
C9962 _446_/a_2560_156# vdd 0.003959f
C9963 _446_/a_2665_112# vss 0.001781f
C9964 _360_/a_36_160# _152_ 0.040508f
C9965 FILLER_0_10_37/a_36_472# FILLER_0_8_37/a_124_375# 0.001512f
C9966 net81 FILLER_0_9_270/a_36_472# 0.084422f
C9967 net72 _404_/a_36_472# 0.019911f
C9968 fanout66/a_36_113# _036_ 0.014556f
C9969 _210_/a_255_603# vss 0.001246f
C9970 _127_ _126_ 0.398279f
C9971 net34 _093_ 0.005701f
C9972 result[7] _102_ 0.010818f
C9973 _094_ _195_/a_67_603# 0.043278f
C9974 _214_/a_36_160# vss 0.007045f
C9975 _086_ FILLER_0_5_181/a_36_472# 0.013437f
C9976 _443_/a_1000_472# vss 0.031435f
C9977 FILLER_0_22_86/a_36_472# _437_/a_36_151# 0.059367f
C9978 output43/a_224_472# output45/a_224_472# 0.246888f
C9979 _009_ FILLER_0_23_274/a_124_375# 0.010723f
C9980 cal_count\[3\] _188_ 0.048745f
C9981 _448_/a_2665_112# vss 0.009029f
C9982 _446_/a_36_151# net66 0.034846f
C9983 FILLER_0_17_72/a_124_375# FILLER_0_17_64/a_124_375# 0.003732f
C9984 _126_ FILLER_0_11_135/a_36_472# 0.002321f
C9985 mask\[1\] _113_ 0.032744f
C9986 FILLER_0_24_130/a_36_472# vdd 0.050082f
C9987 _122_ _163_ 0.156898f
C9988 _425_/a_36_151# FILLER_0_8_247/a_36_472# 0.02628f
C9989 _425_/a_1308_423# FILLER_0_8_247/a_1020_375# 0.001064f
C9990 _423_/a_1308_423# vdd 0.00335f
C9991 _423_/a_448_472# vss 0.002481f
C9992 FILLER_0_16_57/a_1020_375# net55 0.003303f
C9993 FILLER_0_16_57/a_484_472# net72 0.017841f
C9994 _057_ _074_ 0.013823f
C9995 FILLER_0_16_89/a_124_375# vdd 0.01011f
C9996 FILLER_0_5_54/a_1380_472# net47 0.003924f
C9997 net68 _453_/a_1000_472# 0.001816f
C9998 net57 _428_/a_1204_472# 0.015233f
C9999 net62 net29 0.082455f
C10000 FILLER_0_9_28/a_2364_375# _220_/a_67_603# 0.002082f
C10001 _118_ _311_/a_3740_473# 0.001244f
C10002 _016_ FILLER_0_12_136/a_36_472# 0.016227f
C10003 fanout60/a_36_160# FILLER_0_17_282/a_36_472# 0.002647f
C10004 net47 FILLER_0_5_164/a_124_375# 0.011983f
C10005 _057_ _076_ 0.041986f
C10006 net46 output45/a_224_472# 0.005906f
C10007 _126_ FILLER_0_11_101/a_36_472# 0.062336f
C10008 FILLER_0_15_72/a_124_375# cal_count\[1\] 0.00816f
C10009 trim_val\[4\] FILLER_0_5_164/a_484_472# 0.00172f
C10010 _169_ _163_ 0.013133f
C10011 FILLER_0_5_206/a_36_472# net59 0.060133f
C10012 FILLER_0_17_72/a_484_472# vss 0.005334f
C10013 _431_/a_2560_156# net56 0.001258f
C10014 _181_ _402_/a_728_93# 0.064373f
C10015 _134_ FILLER_0_10_107/a_484_472# 0.020725f
C10016 net22 _435_/a_448_472# 0.001929f
C10017 FILLER_0_5_136/a_124_375# vdd 0.035814f
C10018 _132_ FILLER_0_18_107/a_2812_375# 0.002706f
C10019 mask\[0\] _138_ 0.22533f
C10020 FILLER_0_12_20/a_124_375# _039_ 0.004669f
C10021 FILLER_0_4_107/a_36_472# _369_/a_36_68# 0.001709f
C10022 FILLER_0_4_107/a_1020_375# _158_ 0.003535f
C10023 FILLER_0_7_195/a_124_375# _062_ 0.001983f
C10024 _119_ _319_/a_234_472# 0.004559f
C10025 FILLER_0_3_78/a_124_375# _164_ 0.023555f
C10026 _427_/a_1000_472# vss 0.012657f
C10027 _091_ _274_/a_3368_68# 0.001328f
C10028 net17 _450_/a_2449_156# 0.05017f
C10029 trim_mask\[1\] vss 0.449335f
C10030 output11/a_224_472# vss 0.083244f
C10031 output16/a_224_472# vss 0.009875f
C10032 _372_/a_170_472# _070_ 0.024545f
C10033 _436_/a_36_151# FILLER_0_22_107/a_572_375# 0.059049f
C10034 _276_/a_36_160# _093_ 0.019339f
C10035 net76 FILLER_0_3_172/a_572_375# 0.003315f
C10036 _085_ vdd 0.227153f
C10037 FILLER_0_12_220/a_484_472# _070_ 0.004091f
C10038 _130_ net74 0.001655f
C10039 _091_ FILLER_0_15_212/a_932_472# 0.008749f
C10040 net8 FILLER_0_0_266/a_124_375# 0.001181f
C10041 net52 _440_/a_2560_156# 0.004924f
C10042 fanout74/a_36_113# net23 0.005294f
C10043 FILLER_0_21_142/a_572_375# _098_ 0.006558f
C10044 _065_ net17 0.035195f
C10045 net80 _136_ 0.034194f
C10046 trim_val\[0\] _220_/a_67_603# 0.005346f
C10047 _095_ FILLER_0_13_72/a_484_472# 0.027852f
C10048 output31/a_224_472# _094_ 0.004668f
C10049 _452_/a_836_156# _041_ 0.001052f
C10050 _250_/a_36_68# net23 0.002628f
C10051 _408_/a_1936_472# vdd 0.022538f
C10052 mask\[4\] vss 0.426009f
C10053 _091_ _141_ 0.010074f
C10054 net41 _033_ 0.033812f
C10055 net61 output19/a_224_472# 0.077658f
C10056 net49 _440_/a_2560_156# 0.011378f
C10057 net39 _444_/a_448_472# 0.002089f
C10058 _157_ vss 0.039512f
C10059 FILLER_0_7_59/a_36_472# trim_val\[0\] 0.003014f
C10060 FILLER_0_5_206/a_36_472# _122_ 0.003017f
C10061 net72 _217_/a_36_160# 0.068583f
C10062 _142_ vss 0.121933f
C10063 _104_ result[6] 0.096535f
C10064 trim_val\[4\] net65 0.015549f
C10065 _447_/a_2665_112# vss 0.012813f
C10066 fanout77/a_36_113# _419_/a_36_151# 0.002361f
C10067 _373_/a_1254_68# _090_ 0.001326f
C10068 mask\[5\] FILLER_0_19_171/a_124_375# 0.002206f
C10069 FILLER_0_16_57/a_932_472# cal_count\[1\] 0.002217f
C10070 mask\[9\] vss 0.649041f
C10071 _086_ _268_/a_245_68# 0.001044f
C10072 _115_ net14 0.037635f
C10073 output8/a_224_472# _411_/a_36_151# 0.12978f
C10074 FILLER_0_10_37/a_124_375# cal_count\[0\] 0.016543f
C10075 _176_ _125_ 0.089769f
C10076 _096_ _098_ 0.00638f
C10077 result[2] _193_/a_36_160# 0.040932f
C10078 FILLER_0_18_107/a_1020_375# mask\[9\] 0.005758f
C10079 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_124_375# 0.026339f
C10080 FILLER_0_12_136/a_572_375# _120_ 0.001584f
C10081 net60 net62 0.002144f
C10082 _405_/a_67_603# cal_count\[2\] 0.021962f
C10083 FILLER_0_18_100/a_124_375# net14 0.04037f
C10084 net68 _441_/a_36_151# 0.031891f
C10085 FILLER_0_4_185/a_36_472# _087_ 0.008805f
C10086 _106_ output34/a_224_472# 0.01606f
C10087 _431_/a_36_151# FILLER_0_18_107/a_2276_472# 0.002799f
C10088 FILLER_0_17_218/a_36_472# _069_ 0.001246f
C10089 _431_/a_2665_112# _136_ 0.035394f
C10090 _411_/a_2248_156# _073_ 0.003809f
C10091 _444_/a_2665_112# _054_ 0.003576f
C10092 net18 FILLER_0_9_282/a_124_375# 0.024657f
C10093 _414_/a_1000_472# _074_ 0.00222f
C10094 _440_/a_1308_423# _160_ 0.002554f
C10095 net75 _426_/a_448_472# 0.041705f
C10096 net71 _437_/a_448_472# 0.060858f
C10097 output27/a_224_472# fanout65/a_36_113# 0.011564f
C10098 _021_ _097_ 0.002219f
C10099 _435_/a_448_472# vdd 0.029967f
C10100 net50 _376_/a_36_160# 0.018407f
C10101 net38 _444_/a_36_151# 0.009033f
C10102 net53 FILLER_0_17_142/a_484_472# 0.001286f
C10103 mask\[0\] _113_ 0.01678f
C10104 _086_ _057_ 0.82902f
C10105 _410_/a_36_68# cal_count\[0\] 0.007618f
C10106 _141_ FILLER_0_22_128/a_3260_375# 0.003544f
C10107 trim_mask\[1\] FILLER_0_5_88/a_124_375# 0.072632f
C10108 _125_ _124_ 0.085897f
C10109 _449_/a_2248_156# net55 0.052445f
C10110 _422_/a_1204_472# _109_ 0.001807f
C10111 _110_ net35 0.053239f
C10112 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_36_472# 0.026657f
C10113 FILLER_0_16_73/a_572_375# vdd 0.005054f
C10114 _443_/a_448_472# _032_ 0.036717f
C10115 _413_/a_36_151# _088_ 0.001289f
C10116 FILLER_0_8_138/a_36_472# _062_ 0.001109f
C10117 _083_ FILLER_0_3_221/a_484_472# 0.02695f
C10118 trim_mask\[2\] FILLER_0_4_91/a_484_472# 0.0022f
C10119 _444_/a_2665_112# vss 0.002271f
C10120 _444_/a_2560_156# vdd 0.025035f
C10121 _424_/a_2248_156# net36 0.017101f
C10122 result[9] _421_/a_1308_423# 0.011854f
C10123 cal_count\[3\] _186_ 0.012453f
C10124 trim_val\[4\] _443_/a_448_472# 0.038063f
C10125 net41 _446_/a_36_151# 0.143017f
C10126 net25 FILLER_0_23_60/a_36_472# 0.005618f
C10127 _062_ vdd 0.393862f
C10128 net74 FILLER_0_2_127/a_36_472# 0.001261f
C10129 _088_ _078_ 0.047558f
C10130 _079_ _083_ 0.872842f
C10131 net78 _419_/a_1000_472# 0.040603f
C10132 output33/a_224_472# ctlp[1] 0.018552f
C10133 _028_ FILLER_0_7_72/a_2364_375# 0.003884f
C10134 FILLER_0_4_197/a_1020_375# net82 0.00123f
C10135 net38 _452_/a_3129_107# 0.005269f
C10136 FILLER_0_20_2/a_484_472# net43 0.005543f
C10137 _277_/a_36_160# output34/a_224_472# 0.014508f
C10138 _438_/a_2665_112# net14 0.026903f
C10139 mask\[8\] _437_/a_2560_156# 0.001171f
C10140 net80 FILLER_0_19_171/a_124_375# 0.024758f
C10141 FILLER_0_21_28/a_1916_375# vdd -0.009753f
C10142 ctln[8] vdd 0.125219f
C10143 _132_ FILLER_0_16_115/a_36_472# 0.015199f
C10144 FILLER_0_11_78/a_484_472# vss 0.004063f
C10145 _104_ _422_/a_36_151# 0.032235f
C10146 net16 cal_count\[2\] 0.041089f
C10147 FILLER_0_4_197/a_36_472# FILLER_0_3_172/a_2724_472# 0.026657f
C10148 net82 FILLER_0_4_213/a_484_472# 0.002255f
C10149 _232_/a_67_603# FILLER_0_6_47/a_36_472# 0.010206f
C10150 net67 FILLER_0_9_60/a_484_472# 0.001345f
C10151 _176_ cal_count\[2\] 0.005783f
C10152 FILLER_0_4_107/a_1468_375# trim_mask\[4\] 0.00157f
C10153 _077_ _246_/a_36_68# 0.006077f
C10154 ctlp[5] _147_ 0.001406f
C10155 _055_ _060_ 0.181186f
C10156 _058_ _134_ 0.034211f
C10157 _131_ _129_ 0.017222f
C10158 net54 _437_/a_36_151# 0.019307f
C10159 net32 _006_ 0.0012f
C10160 FILLER_0_8_127/a_36_472# _133_ 0.004423f
C10161 _093_ FILLER_0_17_104/a_36_472# 0.014431f
C10162 FILLER_0_4_107/a_1468_375# net47 0.012534f
C10163 net48 net59 0.015963f
C10164 FILLER_0_12_136/a_572_375# state\[2\] 0.001955f
C10165 FILLER_0_12_136/a_1468_375# net53 0.002709f
C10166 ctln[3] _411_/a_448_472# 0.00336f
C10167 FILLER_0_5_164/a_36_472# net37 0.008378f
C10168 net81 net5 0.006276f
C10169 net4 FILLER_0_6_231/a_124_375# 0.002212f
C10170 FILLER_0_2_171/a_36_472# net22 0.081357f
C10171 FILLER_0_6_90/a_36_472# vss 0.001409f
C10172 FILLER_0_6_90/a_484_472# vdd 0.003146f
C10173 _091_ FILLER_0_18_177/a_124_375# 0.010316f
C10174 _139_ FILLER_0_15_180/a_572_375# 0.022254f
C10175 FILLER_0_21_142/a_484_472# net23 0.005353f
C10176 _083_ cal_itt\[1\] 0.046464f
C10177 net32 _103_ 0.038496f
C10178 mask\[5\] FILLER_0_20_177/a_1020_375# 0.013294f
C10179 _418_/a_2665_112# vdd 0.028061f
C10180 _091_ state\[0\] 0.012343f
C10181 _431_/a_2665_112# net53 0.004057f
C10182 mask\[5\] _343_/a_49_472# 0.002228f
C10183 FILLER_0_18_177/a_3172_472# FILLER_0_18_209/a_36_472# 0.013276f
C10184 FILLER_0_16_107/a_572_375# _131_ 0.015859f
C10185 fanout74/a_36_113# FILLER_0_3_142/a_36_472# 0.016516f
C10186 output14/a_224_472# _442_/a_448_472# 0.008149f
C10187 FILLER_0_18_2/a_2364_375# net38 0.001683f
C10188 net35 net14 0.040959f
C10189 net31 _199_/a_36_160# 0.007888f
C10190 FILLER_0_17_72/a_1380_472# _150_ 0.014154f
C10191 net52 FILLER_0_9_72/a_484_472# 0.049391f
C10192 _100_ FILLER_0_12_236/a_484_472# 0.00195f
C10193 net70 _451_/a_36_151# 0.04524f
C10194 net81 FILLER_0_15_235/a_484_472# 0.0047f
C10195 FILLER_0_13_142/a_36_472# net23 0.003007f
C10196 _445_/a_2560_156# net17 0.010829f
C10197 net39 net44 0.0112f
C10198 _057_ _090_ 0.112325f
C10199 ctlp[1] FILLER_0_24_290/a_36_472# 0.037615f
C10200 trim[1] vdd 0.089624f
C10201 output37/a_224_472# _425_/a_2248_156# 0.00114f
C10202 net20 _418_/a_2665_112# 0.013517f
C10203 _287_/a_36_472# _006_ 0.00121f
C10204 _414_/a_1000_472# _081_ 0.006091f
C10205 _425_/a_1308_423# net37 0.002601f
C10206 _077_ FILLER_0_8_156/a_572_375# 0.007238f
C10207 FILLER_0_16_89/a_484_472# _176_ 0.004026f
C10208 _408_/a_728_93# _450_/a_2225_156# 0.00128f
C10209 net58 FILLER_0_8_247/a_1468_375# 0.001669f
C10210 trimb[1] net55 0.017528f
C10211 net52 _453_/a_2665_112# 0.073881f
C10212 net34 result[6] 0.072393f
C10213 FILLER_0_17_142/a_36_472# FILLER_0_17_133/a_124_375# 0.007947f
C10214 FILLER_0_18_2/a_2276_472# vdd 0.004679f
C10215 _002_ net65 0.042811f
C10216 _053_ _072_ 0.001774f
C10217 _289_/a_36_472# _102_ 0.046918f
C10218 _293_/a_36_472# _093_ 0.004121f
C10219 FILLER_0_11_64/a_124_375# cal_count\[3\] 0.002495f
C10220 net57 _250_/a_36_68# 0.001141f
C10221 FILLER_0_24_96/a_36_472# net25 0.040228f
C10222 net4 FILLER_0_8_239/a_36_472# 0.008503f
C10223 output27/a_224_472# FILLER_0_9_290/a_124_375# 0.02894f
C10224 _116_ _055_ 0.72331f
C10225 FILLER_0_1_98/a_36_472# vss 0.002275f
C10226 _442_/a_448_472# FILLER_0_2_127/a_36_472# 0.008634f
C10227 net48 _122_ 0.110769f
C10228 FILLER_0_10_78/a_1468_375# _115_ 0.032403f
C10229 ctln[5] net22 0.072969f
C10230 result[6] net60 0.094624f
C10231 net38 _054_ 0.640545f
C10232 output42/a_224_472# net40 0.003278f
C10233 net82 FILLER_0_3_221/a_36_472# 0.015923f
C10234 net48 FILLER_0_7_233/a_124_375# 0.013455f
C10235 net26 FILLER_0_18_37/a_932_472# 0.002613f
C10236 FILLER_0_4_197/a_572_375# _088_ 0.013597f
C10237 _098_ _438_/a_36_151# 0.009083f
C10238 ctlp[8] mask\[8\] 0.001554f
C10239 vss _022_ 0.067509f
C10240 FILLER_0_8_247/a_1468_375# calibrate 0.006404f
C10241 FILLER_0_12_220/a_572_375# _060_ 0.00145f
C10242 _065_ _447_/a_1308_423# 0.024822f
C10243 _443_/a_36_151# _371_/a_36_113# 0.001252f
C10244 FILLER_0_1_204/a_36_472# vdd 0.009339f
C10245 FILLER_0_1_204/a_124_375# vss 0.018397f
C10246 output44/a_224_472# net43 0.001041f
C10247 net65 FILLER_0_3_221/a_1020_375# 0.001641f
C10248 FILLER_0_3_172/a_3172_472# net22 0.010714f
C10249 valid fanout59/a_36_160# 0.029107f
C10250 _427_/a_2248_156# _043_ 0.001148f
C10251 _175_ FILLER_0_15_72/a_124_375# 0.009573f
C10252 net38 _278_/a_36_160# 0.010587f
C10253 net16 _043_ 0.049385f
C10254 output7/a_224_472# vdd 0.086699f
C10255 _176_ _043_ 0.04106f
C10256 FILLER_0_17_142/a_124_375# vdd 0.020936f
C10257 _308_/a_1084_68# net14 0.002892f
C10258 net18 result[3] 0.237732f
C10259 _120_ FILLER_0_8_156/a_572_375# 0.030218f
C10260 FILLER_0_11_78/a_572_375# _171_ 0.001028f
C10261 net20 FILLER_0_1_204/a_36_472# 0.001278f
C10262 _255_/a_224_552# _116_ 0.027303f
C10263 trimb[1] net17 0.084269f
C10264 net38 vss 0.633752f
C10265 FILLER_0_15_290/a_36_472# net79 0.04083f
C10266 _427_/a_1000_472# _095_ 0.021594f
C10267 _069_ _085_ 0.032519f
C10268 _027_ mask\[9\] 0.050723f
C10269 net38 _178_ 0.123812f
C10270 _164_ _167_ 0.311625f
C10271 _118_ _055_ 0.042556f
C10272 _321_/a_3126_472# _126_ 0.002939f
C10273 _321_/a_358_69# _069_ 0.001124f
C10274 FILLER_0_5_88/a_124_375# FILLER_0_6_90/a_36_472# 0.001543f
C10275 net42 output6/a_224_472# 0.009273f
C10276 _411_/a_796_472# net75 0.006358f
C10277 _104_ _291_/a_36_160# 0.006129f
C10278 net74 FILLER_0_13_142/a_484_472# 0.001771f
C10279 output23/a_224_472# ctlp[6] 0.024575f
C10280 _428_/a_1000_472# _017_ 0.012268f
C10281 FILLER_0_2_171/a_124_375# vss 0.049142f
C10282 FILLER_0_2_171/a_36_472# vdd 0.029996f
C10283 _236_/a_36_160# FILLER_0_8_2/a_36_472# 0.01395f
C10284 _343_/a_49_472# net80 0.001646f
C10285 _162_ _056_ 0.018616f
C10286 _158_ vss 0.007784f
C10287 net16 net68 0.275467f
C10288 FILLER_0_16_241/a_124_375# _198_/a_67_603# 0.002082f
C10289 _408_/a_2215_68# _186_ 0.001205f
C10290 _444_/a_448_472# net47 0.030563f
C10291 FILLER_0_19_125/a_36_472# _145_ 0.004858f
C10292 net2 net5 0.47659f
C10293 fanout50/a_36_160# vdd 0.009536f
C10294 FILLER_0_8_24/a_124_375# net47 0.025599f
C10295 _070_ _313_/a_67_603# 0.004265f
C10296 _141_ net35 0.003655f
C10297 _255_/a_224_552# _118_ 0.002405f
C10298 FILLER_0_18_107/a_932_472# vdd 0.009633f
C10299 _126_ _118_ 0.215385f
C10300 _434_/a_36_151# _146_ 0.003818f
C10301 _434_/a_1204_472# mask\[6\] 0.006692f
C10302 _110_ vdd 0.041979f
C10303 FILLER_0_7_146/a_36_472# _313_/a_67_603# 0.002287f
C10304 FILLER_0_7_104/a_932_472# vdd 0.020291f
C10305 _424_/a_36_151# vss 0.030774f
C10306 _424_/a_448_472# vdd 0.014219f
C10307 cal_count\[2\] _041_ 0.02197f
C10308 _432_/a_448_472# _139_ 0.001772f
C10309 net66 vss 0.265973f
C10310 net41 _444_/a_36_151# 0.013142f
C10311 cal net59 0.297816f
C10312 _074_ _161_ 0.191658f
C10313 result[2] _416_/a_36_151# 0.010509f
C10314 FILLER_0_3_204/a_124_375# FILLER_0_3_212/a_36_472# 0.009654f
C10315 net52 _168_ 0.726039f
C10316 trim_val\[4\] _163_ 0.03439f
C10317 _067_ vss 0.20904f
C10318 _414_/a_448_472# net22 0.047364f
C10319 net50 _441_/a_448_472# 0.074088f
C10320 FILLER_0_4_107/a_1468_375# _154_ 0.005202f
C10321 FILLER_0_4_107/a_572_375# _153_ 0.010165f
C10322 FILLER_0_12_28/a_36_472# net40 0.020589f
C10323 _114_ FILLER_0_10_107/a_124_375# 0.004825f
C10324 output40/a_224_472# trim[2] 0.025041f
C10325 FILLER_0_12_236/a_484_472# _060_ 0.002678f
C10326 FILLER_0_9_223/a_572_375# net4 0.02077f
C10327 fanout60/a_36_160# vss 0.035381f
C10328 _161_ _076_ 0.042123f
C10329 _413_/a_1000_472# vdd 0.002781f
C10330 net49 _168_ 0.031157f
C10331 net34 _422_/a_36_151# 0.032272f
C10332 net18 _417_/a_1308_423# 0.015651f
C10333 _417_/a_448_472# result[3] 0.003109f
C10334 ctln[5] vdd 0.256793f
C10335 _207_/a_67_603# FILLER_0_22_128/a_3260_375# 0.00744f
C10336 _091_ FILLER_0_13_212/a_1380_472# 0.003507f
C10337 FILLER_0_12_136/a_124_375# vdd 0.004378f
C10338 mask\[3\] net21 0.100738f
C10339 _207_/a_67_603# net33 0.005153f
C10340 FILLER_0_21_28/a_1828_472# _423_/a_36_151# 0.059367f
C10341 _437_/a_2665_112# vdd 0.050182f
C10342 result[7] FILLER_0_24_274/a_36_472# 0.006454f
C10343 _115_ _439_/a_2665_112# 0.003617f
C10344 net69 FILLER_0_2_111/a_124_375# 0.010762f
C10345 net61 _422_/a_1308_423# 0.002171f
C10346 net60 _422_/a_36_151# 0.008119f
C10347 FILLER_0_3_172/a_3172_472# vdd 0.003804f
C10348 _129_ _076_ 0.043637f
C10349 _345_/a_36_160# _433_/a_36_151# 0.015565f
C10350 _414_/a_36_151# _057_ 0.003902f
C10351 FILLER_0_7_104/a_1380_472# _125_ 0.001279f
C10352 FILLER_0_7_72/a_1468_375# _164_ 0.003223f
C10353 net16 net67 0.038448f
C10354 fanout61/a_36_113# net79 0.001865f
C10355 _065_ trim_mask\[2\] 0.002792f
C10356 FILLER_0_19_171/a_1380_472# _434_/a_36_151# 0.00271f
C10357 state\[1\] _060_ 0.003973f
C10358 fanout72/a_36_113# net72 0.02315f
C10359 net35 _148_ 0.114816f
C10360 _077_ _439_/a_2560_156# 0.012523f
C10361 FILLER_0_19_142/a_124_375# FILLER_0_19_134/a_124_375# 0.003732f
C10362 _307_/a_234_472# _113_ 0.007518f
C10363 _012_ FILLER_0_23_44/a_1020_375# 0.002827f
C10364 valid net5 0.044555f
C10365 output13/a_224_472# net12 0.002723f
C10366 FILLER_0_4_213/a_36_472# net59 0.044235f
C10367 cal_count\[3\] FILLER_0_12_196/a_36_472# 0.079338f
C10368 net55 _451_/a_3129_107# 0.098091f
C10369 FILLER_0_3_54/a_36_472# vdd 0.00827f
C10370 _144_ _433_/a_2560_156# 0.01064f
C10371 vss rstn 0.149553f
C10372 _069_ _062_ 0.029863f
C10373 net44 clkc 0.184915f
C10374 net57 _395_/a_1044_488# 0.002526f
C10375 output31/a_224_472# _418_/a_2248_156# 0.023576f
C10376 _102_ net19 0.011979f
C10377 _091_ _430_/a_1000_472# 0.025041f
C10378 FILLER_0_14_91/a_124_375# _176_ 0.019567f
C10379 net20 _274_/a_1164_497# 0.002879f
C10380 net10 _411_/a_36_151# 0.127193f
C10381 FILLER_0_22_177/a_572_375# _435_/a_36_151# 0.059049f
C10382 ctlp[1] FILLER_0_23_282/a_484_472# 0.007608f
C10383 FILLER_0_14_181/a_124_375# mask\[1\] 0.044784f
C10384 net57 FILLER_0_13_142/a_36_472# 0.011199f
C10385 vdd net14 2.23064f
C10386 _098_ FILLER_0_20_98/a_36_472# 0.0127f
C10387 FILLER_0_6_79/a_36_472# FILLER_0_6_47/a_3172_472# 0.013276f
C10388 fanout55/a_36_160# vdd 0.016488f
C10389 net54 FILLER_0_18_139/a_932_472# 0.003365f
C10390 _412_/a_1000_472# cal_itt\[1\] 0.012926f
C10391 _414_/a_2248_156# net59 0.004437f
C10392 FILLER_0_9_28/a_484_472# _054_ 0.002831f
C10393 FILLER_0_18_107/a_572_375# net14 0.00258f
C10394 FILLER_0_16_57/a_572_375# FILLER_0_18_61/a_36_472# 0.001512f
C10395 _287_/a_36_472# mask\[2\] 0.00492f
C10396 _177_ FILLER_0_17_72/a_1468_375# 0.026469f
C10397 _245_/a_234_472# net6 0.001301f
C10398 _164_ vdd 0.711488f
C10399 net71 _436_/a_448_472# 0.005274f
C10400 FILLER_0_8_247/a_484_472# vss -0.001894f
C10401 FILLER_0_8_247/a_932_472# vdd 0.008645f
C10402 _144_ vss 0.411237f
C10403 _116_ state\[1\] 0.693219f
C10404 _412_/a_448_472# _082_ 0.022743f
C10405 FILLER_0_17_200/a_36_472# net21 0.036768f
C10406 _432_/a_2560_156# net63 0.00227f
C10407 net55 FILLER_0_18_37/a_36_472# 0.006084f
C10408 _412_/a_448_472# net82 0.030379f
C10409 _414_/a_448_472# vdd 0.013377f
C10410 _066_ vss 0.08113f
C10411 output15/a_224_472# trim_val\[3\] 0.042209f
C10412 FILLER_0_12_136/a_36_472# cal_count\[3\] 0.006102f
C10413 _011_ vdd 0.182751f
C10414 net72 FILLER_0_17_56/a_124_375# 0.018942f
C10415 sample net59 0.001181f
C10416 net78 _421_/a_1308_423# 0.015694f
C10417 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_1020_375# 0.001597f
C10418 net37 net59 0.03883f
C10419 _430_/a_2560_156# net36 0.00164f
C10420 _404_/a_36_472# vdd 0.034854f
C10421 _428_/a_36_151# vdd 0.131612f
C10422 FILLER_0_4_99/a_36_472# FILLER_0_4_91/a_484_472# 0.013276f
C10423 _098_ _433_/a_36_151# 0.023263f
C10424 net38 _450_/a_1040_527# 0.027925f
C10425 _011_ _422_/a_796_472# 0.009261f
C10426 _086_ _161_ 0.077837f
C10427 FILLER_0_21_133/a_124_375# mask\[7\] 0.00145f
C10428 _141_ _433_/a_2665_112# 0.013144f
C10429 net41 _054_ 0.035503f
C10430 net25 vss 0.528437f
C10431 net23 vss 1.922425f
C10432 _131_ _152_ 0.002949f
C10433 net1 _265_/a_224_472# 0.005504f
C10434 FILLER_0_4_49/a_484_472# _160_ 0.001336f
C10435 _057_ _117_ 0.120323f
C10436 _414_/a_2248_156# _122_ 0.002838f
C10437 FILLER_0_14_50/a_36_472# _181_ 0.001514f
C10438 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_572_375# 0.086635f
C10439 _177_ _040_ 0.061289f
C10440 _074_ _056_ 0.002397f
C10441 FILLER_0_8_127/a_124_375# _062_ 0.046401f
C10442 _086_ _129_ 0.051553f
C10443 _149_ FILLER_0_20_107/a_124_375# 0.001244f
C10444 _315_/a_36_68# _120_ 0.00572f
C10445 FILLER_0_16_57/a_484_472# vdd 0.005894f
C10446 FILLER_0_16_57/a_36_472# vss 0.003789f
C10447 net35 _436_/a_2665_112# 0.012468f
C10448 _091_ _429_/a_2248_156# 0.006148f
C10449 output34/a_224_472# ctlp[1] 0.00277f
C10450 FILLER_0_14_81/a_124_375# _176_ 0.001549f
C10451 _112_ _316_/a_848_380# 0.022235f
C10452 _305_/a_36_159# calibrate 0.003505f
C10453 fanout68/a_36_113# net69 0.046009f
C10454 FILLER_0_11_109/a_124_375# FILLER_0_9_105/a_484_472# 0.0027f
C10455 _431_/a_2248_156# FILLER_0_17_142/a_572_375# 0.006739f
C10456 net15 _449_/a_1308_423# 0.015651f
C10457 _354_/a_49_472# net71 0.010421f
C10458 _008_ vdd 0.284571f
C10459 _056_ _076_ 0.938912f
C10460 _061_ _070_ 0.02813f
C10461 net41 vss 0.810444f
C10462 FILLER_0_15_212/a_1468_375# mask\[1\] 0.045287f
C10463 FILLER_0_15_212/a_932_472# vdd 0.001767f
C10464 FILLER_0_10_214/a_36_472# _090_ 0.011963f
C10465 net41 _178_ 0.019945f
C10466 net72 _452_/a_448_472# 0.001296f
C10467 FILLER_0_11_109/a_124_375# vss 0.006764f
C10468 FILLER_0_11_109/a_36_472# vdd 0.109453f
C10469 result[6] FILLER_0_23_290/a_124_375# 0.001492f
C10470 _093_ _438_/a_2248_156# 0.004221f
C10471 _411_/a_1308_423# vss 0.0013f
C10472 _359_/a_244_68# _059_ 0.002986f
C10473 _122_ net37 3.870625f
C10474 _072_ _374_/a_244_472# 0.001816f
C10475 _111_ _438_/a_36_151# 0.003619f
C10476 FILLER_0_20_177/a_1468_375# _434_/a_2248_156# 0.001221f
C10477 _053_ trim_mask\[1\] 0.110786f
C10478 net32 _419_/a_2665_112# 0.027035f
C10479 FILLER_0_5_172/a_36_472# vss 0.003406f
C10480 FILLER_0_9_270/a_484_472# FILLER_0_9_282/a_36_472# 0.002296f
C10481 FILLER_0_4_197/a_36_472# _088_ 0.067725f
C10482 net54 _436_/a_36_151# 0.004179f
C10483 _141_ vdd 0.439746f
C10484 _427_/a_2665_112# _225_/a_36_160# 0.001394f
C10485 _008_ net20 0.153014f
C10486 sample net64 0.209777f
C10487 FILLER_0_13_206/a_36_472# net21 0.00171f
C10488 net62 FILLER_0_15_282/a_484_472# 0.009524f
C10489 _434_/a_1000_472# vdd 0.032431f
C10490 _067_ _450_/a_1040_527# 0.007414f
C10491 ctln[1] FILLER_0_0_232/a_36_472# 0.005158f
C10492 FILLER_0_4_197/a_1380_472# FILLER_0_4_213/a_36_472# 0.013277f
C10493 _429_/a_36_151# _138_ 0.002064f
C10494 _074_ _068_ 0.011897f
C10495 _169_ net37 0.03934f
C10496 net27 _415_/a_2248_156# 0.022666f
C10497 _274_/a_2960_68# _070_ 0.001963f
C10498 result[5] fanout61/a_36_113# 0.001866f
C10499 _174_ _183_ 0.008231f
C10500 _430_/a_2248_156# FILLER_0_15_212/a_932_472# 0.035805f
C10501 FILLER_0_2_171/a_124_375# FILLER_0_2_177/a_36_472# 0.016748f
C10502 _446_/a_2248_156# _160_ 0.002464f
C10503 FILLER_0_11_101/a_484_472# _070_ 0.017841f
C10504 net38 _095_ 0.032393f
C10505 _080_ FILLER_0_3_221/a_932_472# 0.003217f
C10506 vdd FILLER_0_8_156/a_124_375# 0.005213f
C10507 _076_ _068_ 0.35956f
C10508 _013_ _131_ 0.001178f
C10509 net35 FILLER_0_22_128/a_1468_375# 0.015932f
C10510 _291_/a_36_160# _276_/a_36_160# 0.239422f
C10511 output23/a_224_472# vdd 0.033718f
C10512 _428_/a_36_151# _135_ 0.030608f
C10513 _072_ _070_ 2.141346f
C10514 _207_/a_255_603# mask\[6\] 0.003114f
C10515 net35 _207_/a_67_603# 0.005045f
C10516 _088_ _080_ 0.003418f
C10517 net68 FILLER_0_6_47/a_124_375# 0.002491f
C10518 _077_ _219_/a_36_160# 0.01438f
C10519 _064_ _445_/a_1204_472# 0.007445f
C10520 net15 _439_/a_36_151# 0.068183f
C10521 _093_ mask\[8\] 0.004026f
C10522 _406_/a_36_159# cal_count\[2\] 0.028829f
C10523 FILLER_0_4_107/a_932_472# FILLER_0_2_111/a_572_375# 0.001512f
C10524 _397_/a_244_68# net55 0.001173f
C10525 _091_ _248_/a_36_68# 0.071763f
C10526 _217_/a_36_160# vdd 0.092586f
C10527 _174_ FILLER_0_15_59/a_572_375# 0.007123f
C10528 net60 _419_/a_36_151# 0.016173f
C10529 net61 _419_/a_1308_423# 0.00793f
C10530 FILLER_0_4_177/a_124_375# net76 0.003962f
C10531 FILLER_0_17_104/a_572_375# vdd 0.03661f
C10532 _013_ FILLER_0_18_37/a_572_375# 0.003828f
C10533 FILLER_0_5_88/a_36_472# net47 0.003953f
C10534 FILLER_0_3_172/a_36_472# FILLER_0_5_172/a_124_375# 0.0027f
C10535 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_124_375# 0.026339f
C10536 _161_ _090_ 0.207838f
C10537 ctln[2] FILLER_0_1_266/a_36_472# 0.052489f
C10538 ctlp[1] FILLER_0_21_286/a_124_375# 0.025059f
C10539 _148_ vdd 0.01565f
C10540 _147_ _435_/a_36_151# 0.003096f
C10541 FILLER_0_4_197/a_484_472# net76 0.003719f
C10542 cal_count\[3\] _039_ 0.004827f
C10543 trimb[4] _452_/a_3129_107# 0.004943f
C10544 net73 net71 0.033964f
C10545 FILLER_0_10_78/a_1468_375# vdd 0.001778f
C10546 _440_/a_448_472# _029_ 0.043511f
C10547 _372_/a_2590_472# vss 0.00106f
C10548 net69 _170_ 0.006468f
C10549 FILLER_0_3_204/a_124_375# net22 0.031438f
C10550 FILLER_0_12_220/a_1380_472# vss 0.006172f
C10551 net46 net41 0.061224f
C10552 _058_ FILLER_0_8_156/a_484_472# 0.013955f
C10553 FILLER_0_11_109/a_36_472# _135_ 0.001891f
C10554 net58 FILLER_0_9_282/a_36_472# 0.062389f
C10555 FILLER_0_4_123/a_124_375# _152_ 0.039668f
C10556 net63 _434_/a_2248_156# 0.063346f
C10557 FILLER_0_17_72/a_3260_375# _451_/a_1040_527# 0.001117f
C10558 _095_ _067_ 0.00784f
C10559 _060_ _223_/a_36_160# 0.002922f
C10560 net39 _445_/a_1000_472# 0.007782f
C10561 FILLER_0_5_72/a_36_472# trim_mask\[1\] 0.015775f
C10562 FILLER_0_5_72/a_1380_472# _029_ 0.007385f
C10563 net81 FILLER_0_12_236/a_484_472# 0.001419f
C10564 _091_ _432_/a_36_151# 0.054497f
C10565 net68 _030_ 0.007737f
C10566 _036_ net66 0.04474f
C10567 FILLER_0_5_206/a_124_375# net37 0.005485f
C10568 _136_ _038_ 0.061274f
C10569 ctln[1] FILLER_0_1_266/a_36_472# 0.002068f
C10570 FILLER_0_20_193/a_124_375# FILLER_0_20_177/a_1468_375# 0.012222f
C10571 FILLER_0_16_89/a_932_472# net14 0.014714f
C10572 FILLER_0_15_150/a_124_375# vss 0.01957f
C10573 _452_/a_1040_527# net40 0.007832f
C10574 mask\[2\] FILLER_0_16_154/a_932_472# 0.021665f
C10575 _415_/a_36_151# FILLER_0_11_282/a_124_375# 0.001822f
C10576 trimb[1] _452_/a_2449_156# 0.001681f
C10577 FILLER_0_6_37/a_36_472# _160_ 0.008686f
C10578 _053_ _444_/a_2665_112# 0.001698f
C10579 _439_/a_36_151# net51 0.00711f
C10580 _086_ _056_ 0.043494f
C10581 FILLER_0_22_86/a_484_472# _098_ 0.003294f
C10582 FILLER_0_17_72/a_3260_375# _131_ 0.004986f
C10583 trim_mask\[1\] _166_ 0.124855f
C10584 net16 _380_/a_224_472# 0.008718f
C10585 net67 FILLER_0_6_47/a_124_375# 0.005516f
C10586 net55 FILLER_0_13_72/a_484_472# 0.004375f
C10587 vss FILLER_0_19_134/a_124_375# 0.021427f
C10588 vdd FILLER_0_19_134/a_36_472# 0.092128f
C10589 _153_ vdd 0.672318f
C10590 fanout73/a_36_113# vss 0.01873f
C10591 _070_ _319_/a_234_472# 0.004015f
C10592 _449_/a_2560_156# vss 0.002544f
C10593 net80 _435_/a_1000_472# 0.001079f
C10594 FILLER_0_15_116/a_124_375# net70 0.02416f
C10595 FILLER_0_7_72/a_1828_472# net50 0.094122f
C10596 FILLER_0_23_274/a_124_375# vdd 0.014998f
C10597 net26 _423_/a_796_472# 0.001077f
C10598 _030_ _156_ 0.153053f
C10599 net64 FILLER_0_9_282/a_572_375# 0.002322f
C10600 _086_ FILLER_0_11_135/a_124_375# 0.008238f
C10601 _001_ _082_ 0.46787f
C10602 FILLER_0_18_2/a_484_472# output47/a_224_472# 0.00175f
C10603 mask\[0\] FILLER_0_15_212/a_1468_375# 0.001182f
C10604 FILLER_0_3_142/a_36_472# vss 0.012379f
C10605 net82 _001_ 0.044461f
C10606 net63 _202_/a_36_160# 0.004414f
C10607 FILLER_0_5_54/a_572_375# vdd 0.004086f
C10608 FILLER_0_16_107/a_36_472# _132_ 0.001538f
C10609 FILLER_0_17_72/a_1020_375# net36 0.001777f
C10610 _076_ _152_ 0.063574f
C10611 _068_ _081_ 0.006663f
C10612 _451_/a_2225_156# _040_ 0.015815f
C10613 net41 _184_ 0.065857f
C10614 _119_ net23 0.0245f
C10615 net34 _435_/a_1000_472# 0.007444f
C10616 _071_ net23 0.027895f
C10617 mask\[9\] FILLER_0_20_87/a_124_375# 0.004793f
C10618 _402_/a_1948_68# vdd 0.001429f
C10619 _126_ FILLER_0_14_181/a_36_472# 0.008653f
C10620 FILLER_0_18_177/a_124_375# vdd 0.033102f
C10621 FILLER_0_9_28/a_1468_375# net68 0.013121f
C10622 _086_ _068_ 0.080666f
C10623 result[9] ctlp[2] 0.105977f
C10624 _413_/a_2665_112# vss 0.012213f
C10625 _036_ FILLER_0_3_54/a_124_375# 0.010221f
C10626 _449_/a_448_472# _067_ 0.0432f
C10627 net57 vss 0.818311f
C10628 net4 FILLER_0_3_212/a_124_375# 0.001739f
C10629 _127_ _121_ 0.023125f
C10630 FILLER_0_12_20/a_124_375# vdd 0.017452f
C10631 result[5] result[7] 0.016166f
C10632 state\[0\] vdd 0.120171f
C10633 FILLER_0_19_47/a_484_472# _013_ 0.009677f
C10634 net1 _084_ 0.008356f
C10635 FILLER_0_7_72/a_124_375# FILLER_0_7_59/a_572_375# 0.003228f
C10636 _115_ FILLER_0_10_107/a_36_472# 0.016715f
C10637 FILLER_0_19_155/a_484_472# vss 0.004002f
C10638 net66 output41/a_224_472# 0.015427f
C10639 _425_/a_448_472# _014_ 0.013561f
C10640 net58 _412_/a_448_472# 0.044616f
C10641 _214_/a_36_160# _098_ 0.001496f
C10642 mask\[2\] FILLER_0_15_205/a_36_472# 0.001204f
C10643 FILLER_0_5_128/a_572_375# vdd 0.008326f
C10644 FILLER_0_16_57/a_124_375# _183_ 0.005825f
C10645 _053_ FILLER_0_6_90/a_36_472# 0.002495f
C10646 net16 net26 0.273031f
C10647 FILLER_0_3_221/a_932_472# vss 0.002881f
C10648 FILLER_0_3_221/a_1380_472# vdd 0.003819f
C10649 _436_/a_2665_112# vdd 0.007946f
C10650 _436_/a_2248_156# vss 0.002799f
C10651 FILLER_0_4_99/a_124_375# net47 0.001409f
C10652 net20 state\[0\] 0.396139f
C10653 mask\[7\] FILLER_0_22_128/a_124_375# 0.01319f
C10654 _378_/a_224_472# vdd 0.002263f
C10655 FILLER_0_3_204/a_124_375# vdd 0.023302f
C10656 net74 FILLER_0_13_100/a_124_375# 0.005049f
C10657 FILLER_0_9_28/a_1828_472# _042_ 0.001809f
C10658 state\[1\] _228_/a_36_68# 0.024977f
C10659 net63 FILLER_0_20_193/a_124_375# 0.075841f
C10660 FILLER_0_14_123/a_124_375# FILLER_0_14_107/a_1468_375# 0.012001f
C10661 _415_/a_2248_156# net18 0.057604f
C10662 calibrate _313_/a_67_603# 0.021436f
C10663 _439_/a_2248_156# vss 0.003954f
C10664 _439_/a_2665_112# vdd 0.015979f
C10665 FILLER_0_22_128/a_932_472# _433_/a_36_151# 0.002841f
C10666 _289_/a_36_472# _198_/a_67_603# 0.027695f
C10667 _088_ vss 0.326434f
C10668 trim[4] trim[1] 0.001879f
C10669 _104_ net34 0.293336f
C10670 _428_/a_448_472# _043_ 0.063478f
C10671 ctlp[4] net21 0.04068f
C10672 net20 FILLER_0_3_221/a_1380_472# 0.008749f
C10673 _077_ net4 0.656292f
C10674 output29/a_224_472# result[2] 0.058798f
C10675 FILLER_0_21_28/a_1380_472# _424_/a_36_151# 0.001723f
C10676 trimb[4] vss 0.039934f
C10677 ctln[3] FILLER_0_0_232/a_124_375# 0.012394f
C10678 _115_ FILLER_0_9_72/a_1468_375# 0.025664f
C10679 FILLER_0_14_91/a_36_472# _067_ 0.004194f
C10680 FILLER_0_7_162/a_124_375# net37 0.011644f
C10681 mask\[3\] _099_ 0.10534f
C10682 _096_ mask\[1\] 0.010488f
C10683 net79 FILLER_0_13_290/a_124_375# 0.043673f
C10684 FILLER_0_8_138/a_124_375# vdd 0.024547f
C10685 _104_ net60 0.063407f
C10686 net62 FILLER_0_13_290/a_36_472# 0.003157f
C10687 fanout69/a_36_113# _032_ 0.003681f
C10688 FILLER_0_5_109/a_36_472# _153_ 0.034328f
C10689 _008_ _419_/a_796_472# 0.013039f
C10690 _176_ _394_/a_728_93# 0.002001f
C10691 FILLER_0_19_55/a_36_472# net36 0.001068f
C10692 _093_ FILLER_0_17_133/a_36_472# 0.010432f
C10693 FILLER_0_7_72/a_2724_472# vdd 0.007669f
C10694 net72 cal_count\[3\] 0.059493f
C10695 _114_ _085_ 0.056448f
C10696 net5 cal_itt\[1\] 0.057623f
C10697 _414_/a_36_151# _161_ 0.033054f
C10698 net44 FILLER_0_12_2/a_484_472# 0.046864f
C10699 _443_/a_1308_423# _170_ 0.043472f
C10700 _077_ FILLER_0_9_72/a_36_472# 0.006408f
C10701 FILLER_0_10_28/a_124_375# net40 0.047331f
C10702 state\[2\] FILLER_0_13_142/a_124_375# 0.010494f
C10703 _056_ _090_ 0.177189f
C10704 FILLER_0_24_96/a_124_375# net25 0.008342f
C10705 net53 FILLER_0_13_142/a_1020_375# 0.001597f
C10706 _432_/a_2248_156# _137_ 0.001775f
C10707 comp FILLER_0_12_2/a_124_375# 0.007468f
C10708 _095_ net23 0.053365f
C10709 FILLER_0_4_197/a_932_472# net22 0.0473f
C10710 net70 _040_ 0.018254f
C10711 trim_mask\[3\] _156_ 0.002638f
C10712 mask\[5\] net80 0.036014f
C10713 net8 net59 0.062623f
C10714 _448_/a_2665_112# _387_/a_36_113# 0.010064f
C10715 _448_/a_796_472# _037_ 0.009263f
C10716 net63 FILLER_0_18_177/a_1020_375# 0.007516f
C10717 _274_/a_3368_68# _069_ 0.001414f
C10718 vdd output40/a_224_472# 0.079607f
C10719 FILLER_0_22_128/a_1020_375# vss 0.003747f
C10720 FILLER_0_22_128/a_1468_375# vdd 0.016807f
C10721 _233_/a_36_160# _063_ 0.002771f
C10722 _077_ _453_/a_2248_156# 0.013877f
C10723 _077_ _311_/a_1660_473# 0.001653f
C10724 _132_ _127_ 0.112364f
C10725 _408_/a_728_93# _181_ 0.018292f
C10726 result[6] output19/a_224_472# 0.001526f
C10727 _207_/a_67_603# vdd 0.034688f
C10728 FILLER_0_20_15/a_1468_375# net40 0.030032f
C10729 _081_ _152_ 0.172002f
C10730 _161_ _163_ 0.024512f
C10731 _315_/a_244_497# vss 0.008724f
C10732 mask\[5\] net34 0.041303f
C10733 cal_itt\[0\] vss 0.11965f
C10734 net41 _095_ 0.641184f
C10735 _088_ FILLER_0_3_172/a_3260_375# 0.002239f
C10736 _430_/a_1000_472# net22 0.032221f
C10737 net15 _160_ 0.046497f
C10738 _187_ vss 0.080956f
C10739 FILLER_0_3_204/a_36_472# _413_/a_36_151# 0.001723f
C10740 FILLER_0_5_181/a_36_472# net37 0.010376f
C10741 mask\[4\] _098_ 0.041526f
C10742 _004_ net79 0.27387f
C10743 _093_ FILLER_0_18_107/a_124_375# 0.008393f
C10744 FILLER_0_15_282/a_124_375# vdd 0.011964f
C10745 _032_ _371_/a_36_113# 0.030245f
C10746 FILLER_0_16_37/a_124_375# FILLER_0_18_37/a_36_472# 0.001512f
C10747 _016_ vdd 0.114288f
C10748 fanout49/a_36_160# trim_mask\[1\] 0.00358f
C10749 net57 FILLER_0_2_165/a_36_472# 0.001562f
C10750 result[5] net79 0.036275f
C10751 FILLER_0_7_59/a_124_375# trim_mask\[1\] 0.001548f
C10752 FILLER_0_14_91/a_572_375# net14 0.005527f
C10753 _127_ _321_/a_170_472# 0.023836f
C10754 _087_ FILLER_0_5_181/a_124_375# 0.068f
C10755 FILLER_0_17_200/a_572_375# mask\[3\] 0.013879f
C10756 _276_/a_36_160# FILLER_0_18_209/a_572_375# 0.004736f
C10757 mask\[9\] _098_ 0.256513f
C10758 FILLER_0_6_47/a_2276_472# vss 0.004086f
C10759 FILLER_0_6_47/a_2724_472# vdd 0.002467f
C10760 FILLER_0_14_123/a_124_375# vdd 0.034436f
C10761 output45/a_224_472# net17 0.092967f
C10762 _126_ net74 1.001749f
C10763 FILLER_0_20_31/a_36_472# net40 0.045181f
C10764 FILLER_0_10_107/a_124_375# FILLER_0_10_94/a_572_375# 0.003228f
C10765 _412_/a_448_472# fanout81/a_36_160# 0.00998f
C10766 ctlp[4] mask\[7\] 0.080163f
C10767 FILLER_0_4_185/a_124_375# net22 0.004776f
C10768 FILLER_0_5_128/a_124_375# _360_/a_36_160# 0.005705f
C10769 net31 _008_ 0.292444f
C10770 _063_ net49 0.002854f
C10771 fanout52/a_36_160# _386_/a_124_24# 0.004695f
C10772 _053_ FILLER_0_7_104/a_484_472# 0.005353f
C10773 mask\[0\] FILLER_0_13_206/a_36_472# 0.012766f
C10774 FILLER_0_12_2/a_36_472# output6/a_224_472# 0.00108f
C10775 net75 _316_/a_692_472# 0.00138f
C10776 _322_/a_1084_68# _118_ 0.002515f
C10777 net53 state\[2\] 0.001982f
C10778 FILLER_0_13_212/a_932_472# vss 0.022933f
C10779 output39/a_224_472# _034_ 0.002236f
C10780 _066_ _385_/a_36_68# 0.001405f
C10781 _443_/a_448_472# net69 0.068491f
C10782 net26 FILLER_0_21_28/a_2364_375# 0.003691f
C10783 net55 _423_/a_448_472# 0.00206f
C10784 FILLER_0_15_142/a_572_375# net74 0.001652f
C10785 ctlp[1] _420_/a_1000_472# 0.001106f
C10786 _161_ _117_ 0.25528f
C10787 _114_ _062_ 0.028432f
C10788 _308_/a_848_380# _219_/a_36_160# 0.001045f
C10789 _446_/a_2665_112# net17 0.00149f
C10790 _077_ FILLER_0_10_78/a_932_472# 0.002503f
C10791 FILLER_0_4_197/a_932_472# vdd 0.003395f
C10792 _412_/a_36_151# net1 0.020184f
C10793 _072_ _395_/a_244_68# 0.001406f
C10794 result[7] _108_ 0.063624f
C10795 net20 FILLER_0_13_212/a_1380_472# 0.006746f
C10796 _446_/a_2665_112# trim_val\[1\] 0.001275f
C10797 _023_ _146_ 0.006636f
C10798 vdd FILLER_0_5_148/a_36_472# 0.001227f
C10799 vss FILLER_0_5_148/a_572_375# 0.042687f
C10800 FILLER_0_21_142/a_36_472# _210_/a_67_603# 0.001547f
C10801 net52 net50 0.702793f
C10802 output27/a_224_472# FILLER_0_9_270/a_572_375# 0.00135f
C10803 result[7] net19 0.087363f
C10804 net41 output41/a_224_472# 0.008587f
C10805 _037_ net59 0.799647f
C10806 FILLER_0_10_78/a_124_375# FILLER_0_11_78/a_124_375# 0.05841f
C10807 _189_/a_67_603# net62 0.001695f
C10808 _119_ net57 0.30462f
C10809 net73 FILLER_0_18_107/a_3260_375# 0.001629f
C10810 net55 FILLER_0_17_72/a_484_472# 0.019636f
C10811 net57 _071_ 0.12089f
C10812 _139_ mask\[2\] 0.035793f
C10813 _096_ mask\[0\] 0.052773f
C10814 FILLER_0_2_111/a_932_472# vdd 0.003808f
C10815 FILLER_0_2_111/a_124_375# _369_/a_36_68# 0.001176f
C10816 FILLER_0_2_111/a_484_472# vss -0.001894f
C10817 net7 net40 0.025164f
C10818 net34 net80 0.041846f
C10819 net15 _394_/a_718_524# 0.027444f
C10820 net41 _402_/a_1296_93# 0.001707f
C10821 net50 net49 0.238748f
C10822 FILLER_0_9_28/a_1916_375# net68 0.050307f
C10823 _440_/a_1204_472# vss 0.007007f
C10824 _440_/a_2248_156# vdd -0.003421f
C10825 FILLER_0_14_99/a_36_472# FILLER_0_13_100/a_36_472# 0.026657f
C10826 trim_val\[4\] net37 0.003661f
C10827 net18 _418_/a_1000_472# 0.050485f
C10828 _340_/a_36_160# vss 0.029871f
C10829 net62 FILLER_0_15_235/a_124_375# 0.001315f
C10830 _077_ _058_ 3.018054f
C10831 FILLER_0_15_150/a_124_375# _095_ 0.003939f
C10832 net57 FILLER_0_16_154/a_1020_375# 0.001902f
C10833 _020_ vdd 0.194776f
C10834 net82 _443_/a_1000_472# 0.008161f
C10835 _414_/a_36_151# _056_ 0.00356f
C10836 FILLER_0_21_28/a_1828_472# _012_ 0.021162f
C10837 _431_/a_36_151# FILLER_0_17_133/a_36_472# 0.001723f
C10838 net70 FILLER_0_14_107/a_484_472# 0.010987f
C10839 net44 FILLER_0_20_2/a_484_472# 0.039736f
C10840 FILLER_0_7_72/a_1468_375# _376_/a_36_160# 0.02985f
C10841 _050_ FILLER_0_22_128/a_932_472# 0.001098f
C10842 FILLER_0_10_78/a_932_472# _120_ 0.003672f
C10843 FILLER_0_18_2/a_3260_375# FILLER_0_18_37/a_36_472# 0.012267f
C10844 _004_ net75 0.003999f
C10845 FILLER_0_1_266/a_124_375# net8 0.012703f
C10846 FILLER_0_0_96/a_36_472# vdd 0.047982f
C10847 FILLER_0_0_96/a_124_375# vss 0.008342f
C10848 _306_/a_36_68# cal_count\[3\] 0.007663f
C10849 fanout72/a_36_113# vdd -0.002193f
C10850 ctlp[1] _419_/a_1204_472# 0.007338f
C10851 mask\[8\] _352_/a_49_472# 0.002573f
C10852 _086_ _113_ 0.072034f
C10853 net52 FILLER_0_5_72/a_572_375# 0.024148f
C10854 fanout73/a_36_113# _095_ 0.003989f
C10855 _075_ _072_ 0.024301f
C10856 _093_ FILLER_0_17_161/a_36_472# 0.006224f
C10857 _077_ _251_/a_244_472# 0.002492f
C10858 _115_ cal_count\[3\] 0.004426f
C10859 fanout66/a_36_113# trim_mask\[2\] 0.015961f
C10860 _061_ net21 0.049282f
C10861 _144_ _147_ 0.057955f
C10862 FILLER_0_5_72/a_572_375# net49 0.001158f
C10863 _311_/a_66_473# net21 0.02018f
C10864 FILLER_0_4_185/a_124_375# vdd 0.02924f
C10865 FILLER_0_15_2/a_572_375# vdd 0.017581f
C10866 FILLER_0_15_2/a_124_375# vss 0.002713f
C10867 _008_ net77 0.029049f
C10868 _189_/a_67_603# _429_/a_2665_112# 0.015187f
C10869 net63 _430_/a_36_151# 0.026607f
C10870 cal_itt\[2\] _253_/a_672_68# 0.0016f
C10871 _079_ FILLER_0_5_198/a_484_472# 0.008167f
C10872 FILLER_0_19_28/a_36_472# net40 0.020968f
C10873 trim_val\[1\] trim_mask\[1\] 0.519723f
C10874 _058_ _120_ 0.008566f
C10875 net68 FILLER_0_5_54/a_1020_375# 0.00648f
C10876 FILLER_0_5_109/a_572_375# vss 0.055343f
C10877 net15 FILLER_0_7_59/a_572_375# 0.033245f
C10878 mask\[4\] FILLER_0_18_177/a_3260_375# 0.013881f
C10879 net57 _095_ 0.07431f
C10880 _248_/a_36_68# net22 0.002193f
C10881 result[7] _420_/a_36_151# 0.006868f
C10882 net66 _166_ 0.011066f
C10883 net16 _033_ 0.042852f
C10884 _072_ calibrate 0.539702f
C10885 _432_/a_796_472# _093_ 0.002586f
C10886 net36 FILLER_0_15_235/a_36_472# 0.00664f
C10887 FILLER_0_6_177/a_36_472# vdd 0.109918f
C10888 FILLER_0_6_177/a_572_375# vss 0.008666f
C10889 _411_/a_36_151# vdd 0.077963f
C10890 net1 net4 0.03357f
C10891 _376_/a_36_160# vdd -0.006711f
C10892 _147_ net23 0.011375f
C10893 _105_ ctlp[4] 0.002221f
C10894 FILLER_0_5_117/a_36_472# _360_/a_36_160# 0.003913f
C10895 _348_/a_49_472# vss 0.002301f
C10896 _417_/a_796_472# _006_ 0.014427f
C10897 FILLER_0_7_104/a_1468_375# _131_ 0.029718f
C10898 FILLER_0_7_146/a_124_375# _062_ 0.028312f
C10899 _301_/a_36_472# vss 0.003975f
C10900 _438_/a_448_472# _437_/a_36_151# 0.00198f
C10901 mask\[5\] _434_/a_2665_112# 0.003849f
C10902 net36 vss 1.788802f
C10903 _068_ _163_ 0.04926f
C10904 _072_ net21 0.062333f
C10905 _335_/a_49_472# _043_ 0.00367f
C10906 FILLER_0_18_37/a_1380_472# vdd 0.004422f
C10907 _317_/a_36_113# _123_ 0.037893f
C10908 _014_ calibrate 0.403103f
C10909 _053_ net23 0.031487f
C10910 net20 _411_/a_36_151# 0.011179f
C10911 _086_ _321_/a_2590_472# 0.001522f
C10912 output32/a_224_472# _418_/a_448_472# 0.008149f
C10913 _093_ FILLER_0_16_89/a_484_472# 0.001526f
C10914 _429_/a_2248_156# vdd -0.006752f
C10915 _429_/a_1204_472# vss 0.002428f
C10916 _367_/a_244_472# _154_ 0.001775f
C10917 FILLER_0_17_56/a_124_375# vdd 0.008529f
C10918 net79 net19 0.03862f
C10919 FILLER_0_12_220/a_1380_472# FILLER_0_12_236/a_36_472# 0.013277f
C10920 FILLER_0_13_212/a_36_472# mask\[0\] 0.001366f
C10921 net16 _180_ 0.00101f
C10922 FILLER_0_16_107/a_484_472# vss 0.004223f
C10923 FILLER_0_19_195/a_124_375# net21 0.039225f
C10924 _316_/a_124_24# vdd 0.033047f
C10925 _415_/a_448_472# net81 0.004045f
C10926 net79 _416_/a_796_472# 0.01137f
C10927 _176_ _180_ 0.030701f
C10928 net18 _044_ 0.174456f
C10929 net62 _416_/a_1000_472# 0.002399f
C10930 _413_/a_2248_156# FILLER_0_3_212/a_124_375# 0.030666f
C10931 _093_ _150_ 0.406318f
C10932 net20 _429_/a_2248_156# 0.027661f
C10933 FILLER_0_24_130/a_124_375# _050_ 0.007643f
C10934 _093_ FILLER_0_17_72/a_3172_472# 0.012002f
C10935 _193_/a_36_160# vss 0.035228f
C10936 ctlp[2] net78 0.369805f
C10937 _056_ _117_ 0.065147f
C10938 _098_ _022_ 0.013131f
C10939 _017_ vdd 0.26981f
C10940 net26 _424_/a_1308_423# 0.001179f
C10941 _120_ _389_/a_36_148# 0.022887f
C10942 _038_ _389_/a_36_148# 0.003749f
C10943 FILLER_0_10_247/a_36_472# vss 0.002828f
C10944 output44/a_224_472# net44 0.051347f
C10945 result[7] _419_/a_448_472# 0.021809f
C10946 FILLER_0_15_235/a_36_472# FILLER_0_15_228/a_36_472# 0.002765f
C10947 FILLER_0_9_105/a_572_375# FILLER_0_10_107/a_484_472# 0.001543f
C10948 _277_/a_36_160# net30 0.014059f
C10949 _090_ _113_ 0.263235f
C10950 FILLER_0_21_206/a_36_472# net33 0.001447f
C10951 net58 _425_/a_2248_156# 0.051603f
C10952 fanout51/a_36_113# FILLER_0_11_78/a_124_375# 0.005683f
C10953 _451_/a_36_151# net14 0.037503f
C10954 _285_/a_36_472# mask\[1\] 0.036335f
C10955 FILLER_0_5_72/a_1468_375# _164_ 0.040819f
C10956 FILLER_0_10_107/a_36_472# vdd 0.117291f
C10957 FILLER_0_10_107/a_572_375# vss 0.017711f
C10958 FILLER_0_15_228/a_36_472# vss 0.006585f
C10959 FILLER_0_11_282/a_36_472# _416_/a_448_472# 0.011962f
C10960 _452_/a_36_151# vss 0.02741f
C10961 _452_/a_448_472# vdd 0.019824f
C10962 trim_mask\[0\] FILLER_0_10_94/a_484_472# 0.015575f
C10963 net55 FILLER_0_11_78/a_484_472# 0.038269f
C10964 net20 _260_/a_244_472# 0.001593f
C10965 ctlp[5] mask\[7\] 0.131468f
C10966 _320_/a_1568_472# net79 0.001157f
C10967 _256_/a_36_68# _072_ 0.027152f
C10968 FILLER_0_21_142/a_36_472# net54 0.02217f
C10969 en vss 0.466499f
C10970 _068_ _117_ 0.011659f
C10971 FILLER_0_18_177/a_1828_472# net21 0.001887f
C10972 FILLER_0_12_124/a_36_472# vdd 0.040515f
C10973 FILLER_0_12_124/a_124_375# vss 0.012672f
C10974 fanout63/a_36_160# vdd 0.020165f
C10975 _187_ _095_ 0.00765f
C10976 _141_ _140_ 0.131685f
C10977 _425_/a_2248_156# calibrate 0.022237f
C10978 FILLER_0_9_142/a_36_472# vss 0.004305f
C10979 _216_/a_67_603# mask\[9\] 0.003086f
C10980 FILLER_0_5_128/a_484_472# _152_ 0.002283f
C10981 _248_/a_36_68# vdd 0.038887f
C10982 _012_ FILLER_0_21_60/a_124_375# 0.016032f
C10983 _118_ _121_ 0.02882f
C10984 _067_ cal_count\[0\] 0.201595f
C10985 FILLER_0_14_123/a_36_472# _043_ 0.001782f
C10986 FILLER_0_12_136/a_1380_472# net23 0.011488f
C10987 _174_ _181_ 0.079407f
C10988 cal_itt\[2\] FILLER_0_3_221/a_1380_472# 0.015024f
C10989 mask\[7\] _433_/a_36_151# 0.001832f
C10990 net57 _385_/a_36_68# 0.03315f
C10991 _024_ _435_/a_1000_472# 0.002902f
C10992 _417_/a_2665_112# vdd 0.03015f
C10993 FILLER_0_9_72/a_1020_375# vss 0.005622f
C10994 FILLER_0_9_72/a_1468_375# vdd 0.026475f
C10995 net64 _100_ 0.001674f
C10996 _114_ FILLER_0_12_136/a_124_375# 0.006974f
C10997 net20 fanout63/a_36_160# 0.084165f
C10998 net75 FILLER_0_6_239/a_124_375# 0.013962f
C10999 _111_ mask\[9\] 0.127919f
C11000 mask\[5\] FILLER_0_20_193/a_572_375# 0.036451f
C11001 net73 FILLER_0_19_111/a_484_472# 0.007404f
C11002 _093_ FILLER_0_18_139/a_1468_375# 0.004939f
C11003 net36 _195_/a_67_603# 0.034361f
C11004 _128_ vss 0.859962f
C11005 input1/a_36_113# vss 0.05331f
C11006 _421_/a_2665_112# _419_/a_2248_156# 0.001545f
C11007 _428_/a_36_151# _451_/a_36_151# 0.003608f
C11008 _152_ _163_ 0.05157f
C11009 FILLER_0_5_72/a_484_472# net47 0.00169f
C11010 _453_/a_1000_472# vss 0.001738f
C11011 _144_ _345_/a_36_160# 0.00465f
C11012 _311_/a_1212_473# vdd 0.001387f
C11013 output36/a_224_472# _045_ 0.041236f
C11014 FILLER_0_22_128/a_2724_472# _146_ 0.002471f
C11015 cal_count\[2\] FILLER_0_15_2/a_36_472# 0.037661f
C11016 _015_ _426_/a_1000_472# 0.033582f
C11017 _053_ _372_/a_2590_472# 0.001932f
C11018 _017_ _135_ 0.094281f
C11019 net52 FILLER_0_2_101/a_36_472# 0.00749f
C11020 net75 net19 1.345314f
C11021 FILLER_0_16_89/a_484_472# _136_ 0.032722f
C11022 _432_/a_36_151# vdd 0.173104f
C11023 trim_mask\[4\] _160_ 0.244284f
C11024 FILLER_0_18_2/a_124_375# vdd 0.008721f
C11025 FILLER_0_15_150/a_36_472# net23 0.010444f
C11026 FILLER_0_18_177/a_3172_472# net22 0.037136f
C11027 ctln[7] output15/a_224_472# 0.00838f
C11028 net47 _160_ 0.2966f
C11029 FILLER_0_18_2/a_1828_472# net55 0.011802f
C11030 _136_ FILLER_0_16_154/a_124_375# 0.00252f
C11031 _098_ _437_/a_2248_156# 0.008669f
C11032 output34/a_224_472# _199_/a_36_160# 0.003531f
C11033 net58 FILLER_0_8_263/a_36_472# 0.059769f
C11034 FILLER_0_11_142/a_36_472# FILLER_0_11_135/a_124_375# 0.012267f
C11035 _150_ _136_ 0.039815f
C11036 net54 FILLER_0_22_128/a_1380_472# 0.008765f
C11037 mask\[8\] _213_/a_255_603# 0.002776f
C11038 net35 _213_/a_67_603# 0.012955f
C11039 mask\[5\] FILLER_0_18_177/a_1468_375# 0.002726f
C11040 _140_ _148_ 0.011699f
C11041 FILLER_0_17_72/a_3172_472# _136_ 0.002925f
C11042 FILLER_0_16_89/a_124_375# _040_ 0.006315f
C11043 _431_/a_2248_156# _136_ 0.030673f
C11044 _270_/a_36_472# _087_ 0.02676f
C11045 vss _433_/a_1308_423# 0.002695f
C11046 _343_/a_257_69# _093_ 0.001043f
C11047 mask\[0\] _429_/a_796_472# 0.007281f
C11048 _448_/a_2248_156# net59 0.005684f
C11049 _005_ _192_/a_67_603# 0.013886f
C11050 _005_ vdd 0.506158f
C11051 _101_ mask\[1\] 0.033941f
C11052 net27 _323_/a_36_113# 0.010949f
C11053 FILLER_0_3_172/a_1020_375# net22 0.013048f
C11054 _150_ _438_/a_1000_472# 0.003452f
C11055 FILLER_0_18_53/a_124_375# vdd 0.022f
C11056 _114_ net14 0.127764f
C11057 _094_ _418_/a_448_472# 0.042782f
C11058 FILLER_0_18_107/a_932_472# FILLER_0_17_104/a_1380_472# 0.026657f
C11059 _412_/a_36_151# net76 0.001169f
C11060 _052_ _424_/a_1204_472# 0.002681f
C11061 FILLER_0_16_57/a_1020_375# _131_ 0.012481f
C11062 _004_ net19 0.112289f
C11063 FILLER_0_18_107/a_1916_375# _433_/a_36_151# 0.002709f
C11064 ctlp[4] result[8] 0.151286f
C11065 _180_ _041_ 0.00244f
C11066 FILLER_0_8_263/a_36_472# calibrate 0.006968f
C11067 FILLER_0_16_107/a_572_375# FILLER_0_16_115/a_36_472# 0.086635f
C11068 net72 FILLER_0_17_64/a_36_472# 0.001145f
C11069 _136_ _043_ 0.040107f
C11070 net76 FILLER_0_6_177/a_484_472# 0.016333f
C11071 result[5] net19 0.003542f
C11072 _430_/a_1000_472# _069_ 0.00929f
C11073 FILLER_0_4_107/a_36_472# _157_ 0.005289f
C11074 _445_/a_36_151# net40 0.007227f
C11075 FILLER_0_21_28/a_36_472# net40 0.032105f
C11076 net70 FILLER_0_13_100/a_124_375# 0.017886f
C11077 _321_/a_1602_69# _120_ 0.00262f
C11078 net41 _185_ 0.029318f
C11079 FILLER_0_18_2/a_1828_472# net17 0.008573f
C11080 _436_/a_448_472# FILLER_0_22_128/a_124_375# 0.006782f
C11081 net15 _216_/a_255_603# 0.002146f
C11082 net38 net55 0.10956f
C11083 net62 _043_ 0.00426f
C11084 FILLER_0_8_263/a_124_375# net64 0.004793f
C11085 output27/a_224_472# vss 0.027374f
C11086 _053_ FILLER_0_5_54/a_124_375# 0.001571f
C11087 FILLER_0_13_142/a_124_375# _043_ 0.009328f
C11088 FILLER_0_20_177/a_572_375# vdd -0.001627f
C11089 FILLER_0_20_177/a_124_375# vss 0.002674f
C11090 net81 _425_/a_1308_423# 0.004202f
C11091 net64 FILLER_0_14_235/a_124_375# 0.046554f
C11092 _070_ _067_ 0.001869f
C11093 _325_/a_224_472# _129_ 0.003137f
C11094 ctlp[3] _422_/a_448_472# 0.001441f
C11095 _093_ FILLER_0_18_209/a_484_472# 0.014737f
C11096 net16 _447_/a_36_151# 0.133348f
C11097 FILLER_0_16_89/a_1380_472# net36 0.001657f
C11098 _308_/a_848_380# _058_ 0.031449f
C11099 fanout53/a_36_160# net23 0.007461f
C11100 net74 _160_ 0.165289f
C11101 _396_/a_224_472# _177_ 0.001254f
C11102 _053_ net57 0.037224f
C11103 _114_ _428_/a_36_151# 0.008132f
C11104 FILLER_0_20_15/a_572_375# vdd 0.003301f
C11105 net65 FILLER_0_1_266/a_36_472# 0.003529f
C11106 _095_ _451_/a_2449_156# 0.001843f
C11107 _144_ _098_ 1.252524f
C11108 _321_/a_170_472# _118_ 0.034852f
C11109 _141_ FILLER_0_21_150/a_36_472# 0.002773f
C11110 _027_ net36 0.185347f
C11111 _065_ _238_/a_67_603# 0.005075f
C11112 cal_count\[2\] _452_/a_1353_112# 0.002558f
C11113 FILLER_0_17_104/a_124_375# _451_/a_448_472# 0.001718f
C11114 FILLER_0_17_104/a_572_375# _451_/a_36_151# 0.001619f
C11115 FILLER_0_5_212/a_124_375# _081_ 0.01149f
C11116 _441_/a_448_472# vdd 0.007984f
C11117 _441_/a_36_151# vss 0.015116f
C11118 _063_ _165_ 0.021839f
C11119 net64 _060_ 0.05104f
C11120 net55 _424_/a_36_151# 0.007344f
C11121 net38 net17 1.634286f
C11122 net48 _056_ 0.001581f
C11123 _065_ fanout68/a_36_113# 0.005586f
C11124 _058_ FILLER_0_9_105/a_572_375# 0.003832f
C11125 _077_ _134_ 0.043815f
C11126 _132_ net54 0.016007f
C11127 FILLER_0_4_197/a_484_472# _413_/a_36_151# 0.001512f
C11128 net52 _442_/a_2665_112# 0.031179f
C11129 FILLER_0_18_177/a_3172_472# vdd 0.002358f
C11130 _053_ _439_/a_2248_156# 0.002486f
C11131 net55 _067_ 0.053438f
C11132 _033_ FILLER_0_6_47/a_124_375# 0.002521f
C11133 _176_ FILLER_0_10_94/a_124_375# 0.009888f
C11134 _005_ _416_/a_1204_472# 0.014873f
C11135 _256_/a_2960_68# _056_ 0.001168f
C11136 net53 FILLER_0_16_154/a_124_375# 0.003458f
C11137 FILLER_0_9_60/a_484_472# vss 0.005321f
C11138 ctlp[3] _108_ 0.009437f
C11139 FILLER_0_15_142/a_484_472# _431_/a_2248_156# 0.016128f
C11140 _091_ _339_/a_36_160# 0.031941f
C11141 mask\[3\] net56 0.002632f
C11142 net25 _098_ 0.001267f
C11143 _098_ net23 0.036637f
C11144 ctlp[1] _421_/a_796_472# 0.001754f
C11145 _130_ FILLER_0_12_136/a_124_375# 0.010514f
C11146 vss _295_/a_36_472# 0.009751f
C11147 _114_ FILLER_0_11_109/a_36_472# 0.023029f
C11148 FILLER_0_17_142/a_124_375# _137_ 0.006974f
C11149 _429_/a_2665_112# _043_ 0.007641f
C11150 _431_/a_2248_156# net53 0.003335f
C11151 net41 _407_/a_36_472# 0.003257f
C11152 _155_ FILLER_0_6_90/a_572_375# 0.001562f
C11153 net41 cal_count\[0\] 0.001014f
C11154 FILLER_0_17_218/a_484_472# vss 0.035317f
C11155 _285_/a_36_472# _099_ 0.040922f
C11156 FILLER_0_3_172/a_1020_375# vdd 0.009809f
C11157 _131_ _372_/a_170_472# 0.002967f
C11158 _094_ mask\[1\] 0.49634f
C11159 _159_ _160_ 0.021804f
C11160 net76 net4 0.024291f
C11161 net63 FILLER_0_20_177/a_1468_375# 0.018435f
C11162 result[6] _420_/a_448_472# 0.017262f
C11163 _443_/a_2665_112# net22 0.00621f
C11164 _095_ net36 0.127549f
C11165 result[8] result[9] 0.242998f
C11166 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1468_375# 0.086635f
C11167 net16 _444_/a_36_151# 0.010514f
C11168 _091_ _273_/a_36_68# 0.00155f
C11169 FILLER_0_12_220/a_932_472# _223_/a_36_160# 0.001323f
C11170 _104_ output19/a_224_472# 0.064818f
C11171 fanout72/a_36_113# _449_/a_36_151# 0.032681f
C11172 fanout80/a_36_113# vdd 0.033884f
C11173 net50 _165_ 0.056964f
C11174 output28/a_224_472# net79 0.04262f
C11175 _423_/a_36_151# FILLER_0_23_44/a_36_472# 0.001723f
C11176 net48 _068_ 0.054333f
C11177 net78 mask\[7\] 0.001437f
C11178 net66 net17 0.023639f
C11179 net82 FILLER_0_2_171/a_124_375# 0.003818f
C11180 _098_ FILLER_0_15_212/a_484_472# 0.00912f
C11181 net53 _043_ 0.053033f
C11182 _050_ mask\[7\] 0.128172f
C11183 _428_/a_2560_156# net74 0.002759f
C11184 _430_/a_36_151# FILLER_0_18_209/a_36_472# 0.002841f
C11185 FILLER_0_21_28/a_3172_472# FILLER_0_21_60/a_36_472# 0.013276f
C11186 vss _416_/a_36_151# 0.044403f
C11187 _134_ _120_ 0.047627f
C11188 _067_ net17 0.17227f
C11189 _422_/a_448_472# _108_ 0.03293f
C11190 _154_ _160_ 0.395185f
C11191 FILLER_0_8_138/a_36_472# _059_ 0.02252f
C11192 mask\[8\] _149_ 0.0498f
C11193 fanout82/a_36_113# net37 0.046126f
C11194 _086_ FILLER_0_11_142/a_484_472# 0.008338f
C11195 cal_count\[3\] vdd 1.020669f
C11196 ctln[0] net40 0.001334f
C11197 FILLER_0_16_73/a_572_375# _040_ 0.014453f
C11198 result[2] FILLER_0_15_282/a_572_375# 0.0011f
C11199 _058_ _125_ 0.016525f
C11200 _422_/a_448_472# net19 0.003382f
C11201 output31/a_224_472# _417_/a_2248_156# 0.024448f
C11202 output46/a_224_472# FILLER_0_20_15/a_1020_375# 0.001274f
C11203 net23 _387_/a_36_113# 0.031688f
C11204 _059_ vdd 0.161836f
C11205 FILLER_0_19_47/a_36_472# _012_ 0.001667f
C11206 _028_ FILLER_0_6_47/a_3172_472# 0.015585f
C11207 _086_ FILLER_0_7_104/a_1468_375# 0.065371f
C11208 net80 _024_ 0.064854f
C11209 _098_ _434_/a_796_472# 0.001383f
C11210 _414_/a_2560_156# vss 0.001078f
C11211 mask\[4\] net21 0.049513f
C11212 net74 FILLER_0_13_80/a_124_375# 0.012889f
C11213 FILLER_0_14_91/a_124_375# _136_ 0.013064f
C11214 _210_/a_255_603# mask\[7\] 0.001329f
C11215 _118_ _122_ 0.046796f
C11216 _117_ _113_ 0.09166f
C11217 trim_mask\[2\] trim_mask\[1\] 0.002186f
C11218 _091_ _432_/a_2560_156# 0.001542f
C11219 trim_val\[4\] _037_ 0.258184f
C11220 mask\[4\] FILLER_0_19_171/a_932_472# 0.004669f
C11221 net52 FILLER_0_3_78/a_124_375# 0.017889f
C11222 _073_ net59 0.028673f
C11223 result[5] _419_/a_448_472# 0.00232f
C11224 FILLER_0_7_72/a_3260_375# vdd 0.008342f
C11225 _140_ _207_/a_67_603# 0.014923f
C11226 net34 _024_ 0.009705f
C11227 _118_ _227_/a_36_160# 0.017547f
C11228 FILLER_0_9_223/a_36_472# vss 0.019592f
C11229 _070_ net23 0.047632f
C11230 net50 net40 0.005105f
C11231 mask\[5\] output19/a_224_472# 0.092961f
C11232 FILLER_0_10_78/a_1468_375# _114_ 0.01836f
C11233 ctlp[7] _211_/a_36_160# 0.003488f
C11234 _095_ _452_/a_36_151# 0.002974f
C11235 net38 _446_/a_1308_423# 0.010331f
C11236 trim[0] _446_/a_36_151# 0.044586f
C11237 net49 FILLER_0_3_78/a_124_375# 0.001597f
C11238 _030_ FILLER_0_3_78/a_572_375# 0.007667f
C11239 _320_/a_672_472# vdd 0.008437f
C11240 _053_ FILLER_0_6_47/a_2276_472# 0.004472f
C11241 trim_mask\[2\] _157_ 0.002951f
C11242 _069_ _248_/a_36_68# 0.058746f
C11243 net50 FILLER_0_6_79/a_124_375# 0.004402f
C11244 _213_/a_67_603# vdd 0.014901f
C11245 net82 FILLER_0_3_172/a_2724_472# 0.007912f
C11246 FILLER_0_15_150/a_124_375# fanout53/a_36_160# 0.004079f
C11247 FILLER_0_21_206/a_36_472# net22 0.012952f
C11248 net34 FILLER_0_22_128/a_2812_375# 0.005158f
C11249 _093_ FILLER_0_18_107/a_3172_472# 0.008787f
C11250 _405_/a_255_603# vdd 0.001044f
C11251 _405_/a_67_603# vss 0.008564f
C11252 FILLER_0_4_123/a_36_472# fanout69/a_36_113# 0.007864f
C11253 vss FILLER_0_14_235/a_484_472# 0.003246f
C11254 FILLER_0_4_197/a_124_375# _088_ 0.024641f
C11255 _398_/a_36_113# cal_count\[2\] 0.004895f
C11256 _178_ _405_/a_67_603# 0.02427f
C11257 net27 FILLER_0_9_282/a_36_472# 0.002962f
C11258 _101_ _099_ 0.198807f
C11259 _070_ FILLER_0_11_109/a_124_375# 0.002358f
C11260 _122_ _123_ 0.242965f
C11261 _443_/a_2248_156# vss 0.008696f
C11262 _443_/a_2665_112# vdd 0.011824f
C11263 FILLER_0_22_86/a_484_472# _437_/a_448_472# 0.008036f
C11264 _123_ FILLER_0_7_233/a_124_375# 0.007717f
C11265 _073_ _122_ 0.002157f
C11266 FILLER_0_19_28/a_124_375# vdd 0.028695f
C11267 cal_count\[3\] _135_ 0.039115f
C11268 output14/a_224_472# net14 0.018674f
C11269 _446_/a_1308_423# net66 0.005976f
C11270 _429_/a_36_151# FILLER_0_13_206/a_36_472# 0.059367f
C11271 cal_count\[3\] _373_/a_244_68# 0.002341f
C11272 _155_ FILLER_0_7_104/a_36_472# 0.005042f
C11273 _449_/a_2665_112# FILLER_0_13_80/a_124_375# 0.010688f
C11274 _404_/a_36_472# _182_ 0.036415f
C11275 net75 output28/a_224_472# 0.00151f
C11276 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001597f
C11277 trim_mask\[1\] FILLER_0_4_91/a_124_375# 0.006803f
C11278 _423_/a_1000_472# vdd 0.001833f
C11279 _115_ net52 0.022268f
C11280 FILLER_0_22_177/a_36_472# _023_ 0.007019f
C11281 FILLER_0_16_89/a_1020_375# vdd 0.007416f
C11282 FILLER_0_3_204/a_36_472# vss 0.003572f
C11283 net57 _428_/a_2665_112# 0.027291f
C11284 net57 fanout53/a_36_160# 0.009946f
C11285 net62 result[2] 0.311075f
C11286 net41 net55 0.033821f
C11287 net74 _133_ 0.696379f
C11288 net47 FILLER_0_5_164/a_36_472# 0.046908f
C11289 trimb[3] output45/a_224_472# 0.076387f
C11290 _077_ FILLER_0_6_231/a_124_375# 0.009235f
C11291 FILLER_0_4_99/a_124_375# _365_/a_36_68# 0.001918f
C11292 net16 _054_ 0.044357f
C11293 output42/a_224_472# _039_ 0.001254f
C11294 FILLER_0_15_72/a_36_472# cal_count\[1\] 0.006408f
C11295 FILLER_0_14_91/a_124_375# net53 0.065572f
C11296 FILLER_0_20_193/a_572_375# _434_/a_2665_112# 0.002362f
C11297 _105_ net78 0.004705f
C11298 _440_/a_36_151# FILLER_0_6_47/a_1380_472# 0.001512f
C11299 net81 net59 0.074175f
C11300 FILLER_0_17_72/a_1828_472# vdd 0.001969f
C11301 FILLER_0_17_72/a_1380_472# vss 0.003698f
C11302 FILLER_0_20_169/a_124_375# _434_/a_36_151# 0.026916f
C11303 net82 _066_ 0.029681f
C11304 FILLER_0_8_127/a_36_472# _129_ 0.060819f
C11305 FILLER_0_5_136/a_36_472# vss 0.007658f
C11306 FILLER_0_12_20/a_36_472# _039_ 0.007881f
C11307 _004_ output28/a_224_472# 0.024204f
C11308 _035_ _380_/a_224_472# 0.001921f
C11309 _053_ _414_/a_1308_423# 0.029387f
C11310 mask\[5\] mask\[6\] 0.140269f
C11311 ctln[5] _448_/a_448_472# 0.010887f
C11312 FILLER_0_3_78/a_36_472# _164_ 0.022063f
C11313 _427_/a_2248_156# vss 0.018484f
C11314 _427_/a_2665_112# vdd 0.033395f
C11315 FILLER_0_19_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001597f
C11316 net19 _420_/a_36_151# 0.016882f
C11317 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_572_375# 0.086635f
C11318 _372_/a_170_472# _076_ 0.049892f
C11319 _372_/a_2034_472# _133_ 0.001257f
C11320 _436_/a_36_151# FILLER_0_22_107/a_484_472# 0.001723f
C11321 net16 vss 0.679042f
C11322 net27 fanout62/a_36_160# 0.005558f
C11323 net16 _178_ 0.30147f
C11324 _398_/a_36_113# _043_ 0.005985f
C11325 net76 FILLER_0_3_172/a_1468_375# 0.039469f
C11326 _176_ vss 0.761803f
C11327 _000_ _260_/a_36_68# 0.004354f
C11328 _114_ _439_/a_2665_112# 0.011015f
C11329 net57 _098_ 0.062604f
C11330 FILLER_0_5_212/a_36_472# net59 0.058827f
C11331 net34 output19/a_224_472# 0.122464f
C11332 net82 net23 0.18994f
C11333 FILLER_0_21_206/a_36_472# vdd 0.00971f
C11334 FILLER_0_21_206/a_124_375# vss 0.05074f
C11335 net41 net17 0.911377f
C11336 mask\[3\] FILLER_0_18_177/a_484_472# 0.005654f
C11337 net4 FILLER_0_12_236/a_124_375# 0.001558f
C11338 net41 trim_val\[1\] 0.001912f
C11339 output37/a_224_472# en 0.003788f
C11340 _077_ FILLER_0_8_239/a_36_472# 0.001289f
C11341 FILLER_0_6_90/a_124_375# _163_ 0.013948f
C11342 _094_ _099_ 0.193065f
C11343 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3260_375# 0.086635f
C11344 _414_/a_2248_156# _056_ 0.001452f
C11345 _292_/a_36_160# vss 0.009517f
C11346 FILLER_0_18_107/a_3260_375# _145_ 0.00346f
C11347 FILLER_0_4_49/a_124_375# net47 0.006524f
C11348 mask\[7\] _435_/a_36_151# 0.037736f
C11349 net72 _052_ 0.138281f
C11350 _000_ net4 0.036895f
C11351 fanout69/a_36_113# net69 0.040451f
C11352 _077_ FILLER_0_9_28/a_2276_472# 0.003256f
C11353 net22 FILLER_0_18_209/a_124_375# 0.012909f
C11354 net25 FILLER_0_22_86/a_124_375# 0.004298f
C11355 _053_ FILLER_0_6_177/a_572_375# 0.01663f
C11356 net81 FILLER_0_10_256/a_36_472# 0.089055f
C11357 _128_ FILLER_0_12_236/a_36_472# 0.001043f
C11358 _373_/a_1458_68# _113_ 0.001257f
C11359 mask\[5\] FILLER_0_19_171/a_1020_375# 0.007169f
C11360 _124_ vss 0.110847f
C11361 _443_/a_2665_112# FILLER_0_2_165/a_124_375# 0.006271f
C11362 _133_ _154_ 0.0133f
C11363 net81 net64 0.455159f
C11364 FILLER_0_5_109/a_484_472# _160_ 0.001598f
C11365 FILLER_0_18_139/a_124_375# vdd 0.023256f
C11366 mask\[0\] FILLER_0_14_235/a_572_375# 0.002003f
C11367 _274_/a_36_68# net79 0.009814f
C11368 net28 _005_ 0.080653f
C11369 _141_ _137_ 0.40175f
C11370 FILLER_0_9_72/a_572_375# _439_/a_36_151# 0.059049f
C11371 FILLER_0_5_72/a_1468_375# _440_/a_2248_156# 0.030666f
C11372 FILLER_0_5_72/a_1020_375# _440_/a_2665_112# 0.010688f
C11373 FILLER_0_15_282/a_124_375# output30/a_224_472# 0.029138f
C11374 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_572_375# 0.026339f
C11375 FILLER_0_3_172/a_572_375# FILLER_0_2_177/a_36_472# 0.001723f
C11376 net19 _419_/a_448_472# 0.037199f
C11377 FILLER_0_0_130/a_124_375# vdd 0.012493f
C11378 FILLER_0_5_212/a_36_472# _122_ 0.002272f
C11379 FILLER_0_12_28/a_36_472# _039_ 0.007926f
C11380 _405_/a_67_603# _184_ 0.010046f
C11381 _039_ net40 0.036781f
C11382 _036_ _441_/a_36_151# 0.005754f
C11383 FILLER_0_4_144/a_124_375# _370_/a_848_380# 0.005599f
C11384 result[7] _009_ 0.697145f
C11385 fanout71/a_36_113# vss 0.007654f
C11386 _257_/a_36_472# vss 0.023401f
C11387 _074_ _305_/a_36_159# 0.012602f
C11388 _431_/a_36_151# FILLER_0_18_107/a_3172_472# 0.00271f
C11389 _064_ output39/a_224_472# 0.107406f
C11390 _308_/a_848_380# _134_ 0.001299f
C11391 _016_ _428_/a_2248_156# 0.048889f
C11392 FILLER_0_12_136/a_572_375# FILLER_0_13_142/a_36_472# 0.001684f
C11393 _140_ _348_/a_257_69# 0.001089f
C11394 FILLER_0_1_204/a_124_375# net21 0.008041f
C11395 net18 FILLER_0_9_282/a_36_472# 0.041571f
C11396 net75 _426_/a_796_472# 0.003146f
C11397 net71 _437_/a_796_472# 0.006933f
C11398 _106_ net64 0.001587f
C11399 net57 _070_ 0.202843f
C11400 _435_/a_796_472# vdd 0.003478f
C11401 net38 _444_/a_1308_423# 0.007915f
C11402 net80 mask\[6\] 0.080689f
C11403 _187_ cal_count\[0\] 0.645851f
C11404 _016_ _114_ 0.041462f
C11405 FILLER_0_17_72/a_124_375# FILLER_0_15_72/a_36_472# 0.001512f
C11406 FILLER_0_20_87/a_36_472# _438_/a_448_472# 0.004782f
C11407 _103_ _418_/a_1204_472# 0.00582f
C11408 net69 _371_/a_36_113# 0.016091f
C11409 _013_ _183_ 0.00176f
C11410 net2 net59 0.334636f
C11411 _141_ _049_ 0.0035f
C11412 _089_ _414_/a_796_472# 0.001426f
C11413 _068_ net37 0.006392f
C11414 _449_/a_2560_156# net55 0.004835f
C11415 FILLER_0_18_76/a_572_375# vdd -0.009037f
C11416 FILLER_0_18_76/a_124_375# vss 0.006877f
C11417 _443_/a_36_151# trim_mask\[4\] 0.002625f
C11418 mask\[4\] _105_ 0.025209f
C11419 _087_ _074_ 0.004231f
C11420 _069_ cal_count\[3\] 0.012382f
C11421 _134_ FILLER_0_9_105/a_572_375# 0.02163f
C11422 _155_ net47 0.009532f
C11423 _083_ FILLER_0_3_221/a_1380_472# 0.00181f
C11424 net34 mask\[6\] 0.231853f
C11425 result[9] _421_/a_1000_472# 0.012144f
C11426 output8/a_224_472# net75 0.044765f
C11427 _099_ FILLER_0_14_235/a_572_375# 0.013281f
C11428 _069_ _059_ 0.002034f
C11429 FILLER_0_21_125/a_124_375# vdd -0.010326f
C11430 net41 _446_/a_1308_423# 0.056251f
C11431 _320_/a_36_472# _055_ 0.001393f
C11432 output22/a_224_472# ctlp[4] 0.008275f
C11433 net78 _419_/a_2248_156# 0.001614f
C11434 output37/a_224_472# output27/a_224_472# 0.012653f
C11435 fanout70/a_36_113# vdd 0.015969f
C11436 FILLER_0_15_142/a_36_472# vdd 0.106034f
C11437 FILLER_0_6_90/a_36_472# FILLER_0_4_91/a_124_375# 0.001188f
C11438 _448_/a_2248_156# trim_val\[4\] 0.001534f
C11439 net38 _452_/a_2449_156# 0.058386f
C11440 net57 net55 0.001926f
C11441 _371_/a_36_113# _152_ 0.001083f
C11442 output23/a_224_472# _049_ 0.001034f
C11443 _131_ _451_/a_3129_107# 0.001608f
C11444 _432_/a_2665_112# mask\[3\] 0.011428f
C11445 _128_ _426_/a_2248_156# 0.019019f
C11446 net75 FILLER_0_6_231/a_572_375# 0.002577f
C11447 FILLER_0_21_28/a_2812_375# vdd -0.014642f
C11448 FILLER_0_18_209/a_124_375# vdd 0.023676f
C11449 _040_ net14 0.069672f
C11450 fanout58/a_36_160# input4/a_36_68# 0.059453f
C11451 _320_/a_1120_472# _043_ 0.002242f
C11452 _041_ vss 0.012963f
C11453 _126_ _320_/a_36_472# 0.026216f
C11454 net16 _184_ 0.028159f
C11455 FILLER_0_21_28/a_36_472# FILLER_0_20_15/a_1468_375# 0.001723f
C11456 _402_/a_1948_68# _182_ 0.016049f
C11457 net36 FILLER_0_20_87/a_124_375# 0.005853f
C11458 ctln[3] net8 0.003753f
C11459 net49 _167_ 0.031111f
C11460 FILLER_0_2_93/a_124_375# _030_ 0.001641f
C11461 _412_/a_448_472# net18 0.049704f
C11462 net36 _451_/a_448_472# 0.042223f
C11463 _176_ _401_/a_36_68# 0.004263f
C11464 _354_/a_49_472# _433_/a_36_151# 0.001715f
C11465 fanout63/a_36_160# _282_/a_36_160# 0.23939f
C11466 trim_val\[1\] FILLER_0_5_54/a_124_375# 0.001814f
C11467 FILLER_0_7_72/a_2364_375# _053_ 0.015932f
C11468 _125_ _134_ 0.00437f
C11469 _093_ FILLER_0_17_104/a_932_472# 0.014431f
C11470 FILLER_0_5_212/a_36_472# FILLER_0_5_206/a_124_375# 0.016748f
C11471 FILLER_0_4_107/a_484_472# net47 0.001975f
C11472 _267_/a_36_472# vss 0.001495f
C11473 fanout62/a_36_160# net18 0.008106f
C11474 valid net59 0.577796f
C11475 FILLER_0_12_136/a_1468_375# state\[2\] 0.035275f
C11476 FILLER_0_18_209/a_484_472# _047_ 0.002188f
C11477 _091_ FILLER_0_18_177/a_1020_375# 0.002226f
C11478 trimb[4] net55 0.01379f
C11479 _139_ FILLER_0_15_180/a_484_472# 0.004763f
C11480 _095_ _405_/a_67_603# 0.012596f
C11481 output38/a_224_472# output39/a_224_472# 0.002978f
C11482 output28/a_224_472# net19 0.101711f
C11483 mask\[7\] _350_/a_257_69# 0.001135f
C11484 FILLER_0_15_150/a_36_472# net36 0.012318f
C11485 net74 _443_/a_36_151# 0.003682f
C11486 mask\[5\] FILLER_0_20_177/a_36_472# 0.017871f
C11487 _052_ FILLER_0_17_38/a_484_472# 0.001368f
C11488 FILLER_0_9_28/a_1020_375# net16 0.012909f
C11489 net15 _174_ 0.090215f
C11490 _449_/a_36_151# cal_count\[3\] 0.018365f
C11491 trim_mask\[2\] net66 0.036211f
C11492 _427_/a_2248_156# _071_ 0.001131f
C11493 FILLER_0_13_212/a_1380_472# FILLER_0_13_228/a_36_472# 0.013277f
C11494 net82 FILLER_0_3_142/a_36_472# 0.0172f
C11495 FILLER_0_3_172/a_2724_472# net21 0.009426f
C11496 net14 FILLER_0_10_94/a_572_375# 0.047331f
C11497 net52 net22 0.017993f
C11498 _305_/a_36_159# _081_ 0.039192f
C11499 _176_ _071_ 0.002542f
C11500 FILLER_0_17_72/a_1380_472# _027_ 0.00378f
C11501 FILLER_0_17_72/a_2276_472# _150_ 0.003968f
C11502 net52 FILLER_0_9_72/a_1380_472# 0.003507f
C11503 FILLER_0_13_142/a_932_472# net23 0.020589f
C11504 net70 _451_/a_1353_112# 0.00194f
C11505 FILLER_0_21_133/a_36_472# vdd 0.092168f
C11506 result[6] _421_/a_36_151# 0.032036f
C11507 _057_ _060_ 0.033334f
C11508 fanout72/a_36_113# _394_/a_56_524# 0.002775f
C11509 FILLER_0_21_28/a_484_472# FILLER_0_20_31/a_124_375# 0.001723f
C11510 result[7] FILLER_0_23_290/a_36_472# 0.013403f
C11511 _425_/a_1000_472# net37 0.002879f
C11512 _077_ FILLER_0_8_156/a_484_472# 0.006446f
C11513 fanout66/a_36_113# _440_/a_36_151# 0.017895f
C11514 net57 net82 0.91473f
C11515 _413_/a_2665_112# net82 0.004306f
C11516 net72 net40 0.001815f
C11517 _414_/a_1288_156# cal_itt\[3\] 0.001354f
C11518 _340_/a_36_160# _098_ 0.019601f
C11519 FILLER_0_18_2/a_3172_472# vdd 0.011201f
C11520 FILLER_0_13_80/a_36_472# _451_/a_3129_107# 0.001115f
C11521 net57 fanout57/a_36_113# 0.004316f
C11522 _132_ net74 0.031741f
C11523 trimb[4] net17 0.004628f
C11524 net41 _408_/a_1336_472# 0.063099f
C11525 trim_mask\[4\] net59 0.012971f
C11526 _085_ _055_ 0.240451f
C11527 _277_/a_36_160# _103_ 0.032112f
C11528 _432_/a_2665_112# FILLER_0_17_200/a_36_472# 0.007491f
C11529 output29/a_224_472# vss 0.013148f
C11530 _087_ _081_ 0.002169f
C11531 ctln[5] net12 0.41364f
C11532 net82 FILLER_0_3_221/a_932_472# 0.004092f
C11533 _426_/a_36_151# vss 0.003014f
C11534 _426_/a_448_472# vdd 0.042167f
C11535 _098_ _438_/a_1308_423# 0.004124f
C11536 FILLER_0_8_247/a_484_472# calibrate 0.009318f
C11537 FILLER_0_12_220/a_484_472# _090_ 0.006993f
C11538 FILLER_0_12_220/a_1468_375# _060_ 0.001429f
C11539 FILLER_0_7_72/a_1468_375# net52 0.003576f
C11540 _337_/a_49_472# mask\[2\] 0.00188f
C11541 _065_ _447_/a_1000_472# 0.03162f
C11542 output13/a_224_472# net59 0.007733f
C11543 _086_ _087_ 0.015938f
C11544 _021_ mask\[3\] 0.036781f
C11545 trim_mask\[2\] FILLER_0_3_54/a_124_375# 0.015198f
C11546 valid net64 0.022969f
C11547 _016_ _130_ 0.114514f
C11548 _088_ net82 0.160444f
C11549 _233_/a_36_160# vdd 0.064615f
C11550 _427_/a_36_151# net74 0.04306f
C11551 FILLER_0_2_93/a_572_375# net14 0.044606f
C11552 _175_ FILLER_0_15_72/a_36_472# 0.006746f
C11553 net72 FILLER_0_17_38/a_572_375# 0.010272f
C11554 result[9] net18 0.019413f
C11555 net73 _433_/a_36_151# 0.004541f
C11556 fanout53/a_36_160# net36 0.028652f
C11557 _190_/a_36_160# _043_ 0.06415f
C11558 FILLER_0_17_64/a_36_472# vdd 0.094397f
C11559 FILLER_0_17_64/a_124_375# vss 0.022351f
C11560 FILLER_0_17_142/a_572_375# vss 0.049716f
C11561 FILLER_0_17_142/a_36_472# vdd 0.108843f
C11562 _155_ _154_ 0.18488f
C11563 FILLER_0_6_47/a_572_375# vdd 0.003158f
C11564 _028_ _058_ 0.041158f
C11565 _057_ _116_ 0.028033f
C11566 _093_ FILLER_0_18_177/a_2364_375# 0.001989f
C11567 trim[0] vss 0.132654f
C11568 _072_ FILLER_0_10_214/a_124_375# 0.033245f
C11569 _427_/a_2248_156# _095_ 0.022479f
C11570 _321_/a_170_472# net74 0.020269f
C11571 _126_ _085_ 0.02154f
C11572 FILLER_0_2_93/a_124_375# trim_mask\[3\] 0.003033f
C11573 FILLER_0_4_177/a_572_375# net22 0.006125f
C11574 mask\[9\] FILLER_0_19_111/a_124_375# 0.031474f
C11575 net16 _095_ 0.042842f
C11576 FILLER_0_16_255/a_36_472# _417_/a_2665_112# 0.003221f
C11577 FILLER_0_24_290/a_124_375# FILLER_0_24_274/a_1468_375# 0.012001f
C11578 output15/a_224_472# _383_/a_36_472# 0.001154f
C11579 net42 net6 0.166896f
C11580 _176_ _095_ 0.064978f
C11581 FILLER_0_3_142/a_124_375# _443_/a_36_151# 0.059049f
C11582 _258_/a_36_160# net59 0.003167f
C11583 calibrate net23 0.032259f
C11584 result[5] _290_/a_224_472# 0.001638f
C11585 clk rstn 0.541051f
C11586 fanout54/a_36_160# net23 0.05522f
C11587 _339_/a_36_160# vdd 0.01226f
C11588 _162_ _061_ 0.001665f
C11589 net16 _036_ 0.637538f
C11590 _122_ net47 0.030693f
C11591 _045_ _006_ 0.00216f
C11592 _050_ _436_/a_448_472# 0.064832f
C11593 FILLER_0_16_37/a_36_472# net47 0.008304f
C11594 net20 _256_/a_244_497# 0.005033f
C11595 _098_ _348_/a_49_472# 0.011096f
C11596 _430_/a_448_472# net81 0.003775f
C11597 _301_/a_36_472# _098_ 0.010091f
C11598 net52 vdd 1.32956f
C11599 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_572_375# 0.086635f
C11600 _114_ _017_ 0.071595f
C11601 net36 _098_ 3.387566f
C11602 FILLER_0_8_24/a_36_472# net47 0.097212f
C11603 _076_ _313_/a_67_603# 0.024219f
C11604 _127_ _129_ 0.716384f
C11605 FILLER_0_17_104/a_36_472# _438_/a_2248_156# 0.001731f
C11606 _139_ _138_ 0.00256f
C11607 _057_ _118_ 0.055726f
C11608 FILLER_0_18_107/a_1828_472# vdd 0.004446f
C11609 cal_itt\[0\] _082_ 0.018597f
C11610 _434_/a_2665_112# mask\[6\] 0.026286f
C11611 trim_mask\[4\] _169_ 0.042442f
C11612 _273_/a_36_68# vdd 0.041825f
C11613 net35 _434_/a_2248_156# 0.026885f
C11614 _010_ FILLER_0_23_274/a_36_472# 0.008718f
C11615 net82 cal_itt\[0\] 0.063072f
C11616 _102_ vdd 0.211559f
C11617 _285_/a_36_472# _196_/a_36_160# 0.004619f
C11618 FILLER_0_7_104/a_1380_472# vss 0.003236f
C11619 _424_/a_796_472# vdd 0.001951f
C11620 FILLER_0_17_104/a_572_375# _040_ 0.001228f
C11621 _413_/a_2248_156# ctln[4] 0.001253f
C11622 net41 FILLER_0_16_37/a_124_375# 0.008195f
C11623 _030_ vss 0.117034f
C11624 net49 vdd 0.872948f
C11625 net47 _169_ 0.528536f
C11626 _089_ cal_itt\[3\] 0.049851f
C11627 net41 _444_/a_1308_423# 0.015841f
C11628 _320_/a_36_472# state\[1\] 0.013058f
C11629 output29/a_224_472# _416_/a_2248_156# 0.024448f
C11630 net81 mask\[2\] 0.002083f
C11631 net50 _168_ 0.306226f
C11632 _122_ FILLER_0_5_172/a_124_375# 0.001352f
C11633 _027_ FILLER_0_18_76/a_124_375# 0.001285f
C11634 net41 FILLER_0_8_24/a_572_375# 0.003909f
C11635 _173_ _408_/a_728_93# 0.022838f
C11636 mask\[4\] FILLER_0_18_139/a_1380_472# 0.003851f
C11637 FILLER_0_19_55/a_124_375# _052_ 0.053626f
C11638 net50 _441_/a_796_472# 0.010626f
C11639 FILLER_0_4_107/a_484_472# _154_ 0.040595f
C11640 _129_ FILLER_0_11_135/a_36_472# 0.078373f
C11641 _114_ FILLER_0_10_107/a_36_472# 0.00263f
C11642 FILLER_0_19_47/a_124_375# FILLER_0_18_37/a_1380_472# 0.001684f
C11643 _429_/a_2248_156# FILLER_0_13_228/a_36_472# 0.035805f
C11644 FILLER_0_9_223/a_484_472# _128_ 0.005152f
C11645 net20 _102_ 0.081029f
C11646 net61 vss 0.254538f
C11647 _258_/a_36_160# _122_ 0.00102f
C11648 net27 _425_/a_2248_156# 0.027078f
C11649 net18 _417_/a_1000_472# 0.056791f
C11650 FILLER_0_16_57/a_124_375# net15 0.001594f
C11651 output22/a_224_472# ctlp[5] 0.024131f
C11652 _417_/a_1204_472# net30 0.001496f
C11653 _417_/a_796_472# result[3] 0.001206f
C11654 _258_/a_36_160# FILLER_0_7_233/a_124_375# 0.001633f
C11655 _062_ _055_ 0.29425f
C11656 FILLER_0_9_28/a_1468_375# _054_ 0.005381f
C11657 _072_ _162_ 0.090175f
C11658 FILLER_0_12_136/a_572_375# vss 0.006091f
C11659 FILLER_0_12_136/a_1020_375# vdd 0.017472f
C11660 _441_/a_2248_156# _030_ 0.003495f
C11661 _149_ _026_ 0.243704f
C11662 _207_/a_67_603# _049_ 0.003205f
C11663 FILLER_0_21_28/a_2276_472# _423_/a_448_472# 0.008036f
C11664 _259_/a_271_68# net4 0.003663f
C11665 FILLER_0_8_239/a_124_375# vdd 0.035205f
C11666 _415_/a_2560_156# result[1] 0.002282f
C11667 result[7] FILLER_0_24_274/a_932_472# 0.006454f
C11668 _114_ FILLER_0_12_124/a_36_472# 0.003953f
C11669 output32/a_224_472# net18 0.022521f
C11670 _428_/a_36_151# FILLER_0_14_107/a_484_472# 0.059367f
C11671 _065_ output15/a_224_472# 0.037721f
C11672 net69 FILLER_0_2_111/a_1020_375# 0.018655f
C11673 _031_ FILLER_0_2_111/a_124_375# 0.05482f
C11674 FILLER_0_6_239/a_124_375# FILLER_0_6_231/a_572_375# 0.012001f
C11675 net61 _422_/a_1000_472# 0.001947f
C11676 FILLER_0_18_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001684f
C11677 _432_/a_2560_156# vdd 0.003219f
C11678 _106_ mask\[2\] 0.039965f
C11679 trimb[3] net38 0.002836f
C11680 net38 output6/a_224_472# 0.060017f
C11681 _414_/a_2560_156# _053_ 0.008732f
C11682 _098_ FILLER_0_15_228/a_36_472# 0.022074f
C11683 _267_/a_36_472# _071_ 0.001682f
C11684 net67 _190_/a_36_160# 0.023989f
C11685 FILLER_0_23_282/a_36_472# FILLER_0_23_274/a_36_472# 0.002296f
C11686 FILLER_0_9_223/a_124_375# vdd 0.006153f
C11687 _144_ mask\[7\] 0.111088f
C11688 _091_ _430_/a_36_151# 0.02228f
C11689 net20 FILLER_0_8_239/a_124_375# 0.004302f
C11690 net35 _025_ 0.02169f
C11691 _110_ _437_/a_36_151# 0.00125f
C11692 _093_ _304_/a_224_472# 0.002907f
C11693 _096_ _090_ 0.026104f
C11694 FILLER_0_19_142/a_36_472# FILLER_0_19_134/a_36_472# 0.002296f
C11695 net16 _402_/a_1296_93# 0.053493f
C11696 ctln[6] net22 0.014307f
C11697 FILLER_0_4_177/a_124_375# vss 0.002462f
C11698 FILLER_0_4_177/a_572_375# vdd 0.001622f
C11699 _255_/a_224_552# _062_ 0.009032f
C11700 net7 ctln[0] 0.001209f
C11701 _008_ _418_/a_36_151# 0.016984f
C11702 net15 FILLER_0_15_59/a_124_375# 0.007439f
C11703 net36 FILLER_0_15_180/a_124_375# 0.004275f
C11704 _406_/a_36_159# _278_/a_36_160# 0.001331f
C11705 _411_/a_1000_472# net75 0.03227f
C11706 FILLER_0_14_91/a_36_472# _176_ 0.076419f
C11707 _359_/a_36_488# vss 0.002427f
C11708 FILLER_0_21_133/a_124_375# FILLER_0_21_142/a_124_375# 0.003228f
C11709 FILLER_0_22_177/a_1468_375# _435_/a_36_151# 0.059049f
C11710 net51 _450_/a_3129_107# 0.030082f
C11711 mask\[4\] output18/a_224_472# 0.017718f
C11712 _035_ _446_/a_36_151# 0.012914f
C11713 output11/a_224_472# ctln[1] 0.004299f
C11714 FILLER_0_13_228/a_124_375# net4 0.002641f
C11715 _406_/a_36_159# vss 0.002509f
C11716 _086_ FILLER_0_5_117/a_36_472# 0.042352f
C11717 net57 FILLER_0_13_142/a_932_472# 0.01158f
C11718 net75 _265_/a_244_68# 0.046186f
C11719 _178_ _406_/a_36_159# 0.007052f
C11720 mask\[7\] net23 0.225177f
C11721 _091_ net79 0.052824f
C11722 FILLER_0_15_72/a_572_375# vdd 0.003801f
C11723 FILLER_0_15_72/a_124_375# vss 0.048711f
C11724 _101_ _196_/a_36_160# 0.009836f
C11725 FILLER_0_20_193/a_572_375# mask\[6\] 0.001262f
C11726 net43 FILLER_0_20_15/a_572_375# 0.003924f
C11727 _067_ output6/a_224_472# 0.001611f
C11728 net81 FILLER_0_15_212/a_572_375# 0.006974f
C11729 trim_mask\[3\] vss 0.156544f
C11730 net52 FILLER_0_2_165/a_124_375# 0.002214f
C11731 net27 FILLER_0_8_263/a_36_472# 0.003956f
C11732 FILLER_0_8_247/a_1380_472# vss 0.001338f
C11733 FILLER_0_18_2/a_3260_375# net41 0.042057f
C11734 net47 FILLER_0_4_91/a_572_375# 0.008167f
C11735 input2/a_36_113# rstn 0.002202f
C11736 _095_ _041_ 0.002104f
C11737 FILLER_0_16_73/a_484_472# net15 0.001946f
C11738 _085_ state\[1\] 0.182697f
C11739 _093_ FILLER_0_18_100/a_36_472# 0.077197f
C11740 net27 FILLER_0_14_235/a_572_375# 0.006429f
C11741 _441_/a_2665_112# net14 0.00104f
C11742 net55 net36 0.273956f
C11743 _083_ _260_/a_244_472# 0.00134f
C11744 net55 FILLER_0_18_37/a_932_472# 0.00769f
C11745 _020_ _137_ 0.228674f
C11746 ctlp[3] _009_ 0.018168f
C11747 net80 FILLER_0_17_161/a_36_472# 0.003342f
C11748 net15 trim_val\[3\] 0.068273f
C11749 FILLER_0_12_136/a_932_472# cal_count\[3\] 0.007247f
C11750 _067_ _171_ 0.007069f
C11751 net72 FILLER_0_17_56/a_36_472# 0.008058f
C11752 ctlp[7] output25/a_224_472# 0.002088f
C11753 _144_ FILLER_0_18_107/a_1916_375# 0.003148f
C11754 FILLER_0_17_226/a_124_375# mask\[3\] 0.010642f
C11755 _070_ FILLER_0_10_107/a_572_375# 0.003959f
C11756 net78 _421_/a_1000_472# 0.022212f
C11757 _229_/a_224_472# net22 0.007346f
C11758 net38 net3 0.103189f
C11759 _412_/a_448_472# net65 0.043862f
C11760 ctlp[8] vss 0.107975f
C11761 _441_/a_2665_112# _164_ 0.021931f
C11762 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3260_375# 0.001597f
C11763 _412_/a_2665_112# net1 0.063655f
C11764 FILLER_0_3_221/a_484_472# net59 0.001655f
C11765 _093_ FILLER_0_17_72/a_1020_375# 0.001994f
C11766 mask\[5\] output35/a_224_472# 0.003461f
C11767 output12/a_224_472# net76 0.00803f
C11768 _428_/a_1308_423# vdd 0.004352f
C11769 _098_ _433_/a_1308_423# 0.010653f
C11770 net22 _202_/a_36_160# 0.052766f
C11771 net10 net75 0.073869f
C11772 net38 _450_/a_1293_527# 0.001307f
C11773 _077_ _392_/a_36_68# 0.055912f
C11774 _011_ _422_/a_1204_472# 0.002176f
C11775 net4 _078_ 0.487587f
C11776 _437_/a_36_151# net14 0.014361f
C11777 net13 vss 0.071697f
C11778 _127_ FILLER_0_11_135/a_124_375# 0.040456f
C11779 _182_ FILLER_0_18_37/a_1380_472# 0.004074f
C11780 _079_ net59 0.102335f
C11781 net1 _265_/a_916_472# 0.002088f
C11782 ctlp[9] FILLER_0_23_44/a_932_472# 0.001195f
C11783 FILLER_0_21_142/a_484_472# FILLER_0_22_128/a_1916_375# 0.001543f
C11784 FILLER_0_11_142/a_124_375# net23 0.002992f
C11785 FILLER_0_13_80/a_36_472# FILLER_0_13_72/a_484_472# 0.013277f
C11786 _432_/a_796_472# net80 0.007731f
C11787 _074_ _061_ 0.007152f
C11788 _422_/a_448_472# _009_ 0.018984f
C11789 FILLER_0_16_57/a_1380_472# vdd 0.005673f
C11790 FILLER_0_16_57/a_932_472# vss 0.003388f
C11791 _077_ FILLER_0_10_78/a_1380_472# 0.001548f
C11792 _091_ _429_/a_2560_156# 0.001502f
C11793 ctln[6] vdd 0.116327f
C11794 net57 calibrate 0.037299f
C11795 _112_ _316_/a_1152_472# 0.001449f
C11796 net20 _256_/a_1164_497# 0.001462f
C11797 cal_count\[3\] FILLER_0_11_124/a_124_375# 0.002147f
C11798 _127_ _068_ 0.052712f
C11799 _128_ _070_ 1.279188f
C11800 _131_ _331_/a_244_472# 0.002331f
C11801 net15 _449_/a_1000_472# 0.056791f
C11802 FILLER_0_20_177/a_124_375# _098_ 0.018701f
C11803 _061_ _076_ 0.024289f
C11804 FILLER_0_15_212/a_1380_472# vss 0.007595f
C11805 _246_/a_36_68# vss 0.024639f
C11806 FILLER_0_15_212/a_484_472# mask\[1\] 0.007258f
C11807 FILLER_0_10_214/a_36_472# _060_ 0.001378f
C11808 net55 _452_/a_36_151# 0.042427f
C11809 net81 FILLER_0_15_205/a_124_375# 0.015134f
C11810 _431_/a_448_472# net70 0.002293f
C11811 _119_ FILLER_0_7_104/a_1380_472# 0.002603f
C11812 _076_ _311_/a_66_473# 0.003077f
C11813 FILLER_0_19_125/a_124_375# _433_/a_36_151# 0.001597f
C11814 _413_/a_2665_112# net21 0.002828f
C11815 _281_/a_672_472# vdd 0.001069f
C11816 _187_ _408_/a_1336_472# 0.002191f
C11817 result[7] FILLER_0_23_282/a_572_375# 0.015853f
C11818 _094_ net18 0.468109f
C11819 _093_ FILLER_0_19_142/a_124_375# 0.00346f
C11820 FILLER_0_7_162/a_124_375# net47 0.030995f
C11821 _425_/a_36_151# _316_/a_124_24# 0.036238f
C11822 FILLER_0_4_197/a_1020_375# FILLER_0_5_206/a_36_472# 0.001723f
C11823 net54 _436_/a_1308_423# 0.002665f
C11824 _245_/a_234_472# net47 0.00188f
C11825 net57 _333_/a_36_160# 0.008292f
C11826 _392_/a_36_68# _120_ 0.001738f
C11827 mask\[9\] _354_/a_49_472# 0.032687f
C11828 trim_mask\[1\] FILLER_0_6_47/a_36_472# 0.004319f
C11829 _414_/a_36_151# _087_ 0.010359f
C11830 _073_ FILLER_0_3_221/a_1020_375# 0.002563f
C11831 _434_/a_2248_156# vdd 0.019386f
C11832 FILLER_0_7_72/a_1380_472# net52 0.003507f
C11833 FILLER_0_5_88/a_36_472# _164_ 0.011718f
C11834 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_124_375# 0.005439f
C11835 _094_ _196_/a_36_160# 0.001668f
C11836 FILLER_0_1_98/a_124_375# trim_val\[3\] 0.001628f
C11837 _079_ _122_ 0.003853f
C11838 cal_itt\[1\] net59 0.227495f
C11839 _091_ FILLER_0_19_171/a_572_375# 0.013568f
C11840 FILLER_0_1_212/a_36_472# FILLER_0_1_204/a_124_375# 0.009654f
C11841 _009_ _108_ 1.645945f
C11842 _072_ _074_ 2.017168f
C11843 _421_/a_36_151# _419_/a_36_151# 0.561555f
C11844 _057_ _228_/a_36_68# 0.002062f
C11845 _043_ FILLER_0_12_196/a_124_375# 0.003935f
C11846 output27/a_224_472# fanout64/a_36_160# 0.027335f
C11847 FILLER_0_10_78/a_1380_472# _120_ 0.003228f
C11848 FILLER_0_15_290/a_124_375# vss 0.032056f
C11849 FILLER_0_15_290/a_36_472# vdd 0.092839f
C11850 net19 _009_ 0.055383f
C11851 _088_ net21 0.053843f
C11852 vdd FILLER_0_8_156/a_36_472# 0.002891f
C11853 vss FILLER_0_8_156/a_572_375# 0.007969f
C11854 state\[1\] _062_ 0.001179f
C11855 cal_count\[3\] FILLER_0_12_50/a_36_472# 0.063276f
C11856 net35 FILLER_0_22_128/a_2364_375# 0.012732f
C11857 net17 _452_/a_36_151# 0.041497f
C11858 _087_ _163_ 0.004829f
C11859 FILLER_0_9_28/a_1916_375# _054_ 0.005889f
C11860 _072_ _076_ 0.068172f
C11861 FILLER_0_18_100/a_36_472# _136_ 0.003419f
C11862 _216_/a_67_603# net36 0.028132f
C11863 FILLER_0_13_100/a_124_375# net14 0.041373f
C11864 net58 cal_itt\[0\] 0.229955f
C11865 net68 FILLER_0_6_47/a_1020_375# 0.029857f
C11866 _254_/a_448_472# _072_ 0.002611f
C11867 _074_ _014_ 0.001557f
C11868 _077_ _120_ 0.205715f
C11869 _064_ _445_/a_2665_112# 0.004701f
C11870 _185_ _405_/a_67_603# 0.060789f
C11871 FILLER_0_4_107/a_1380_472# FILLER_0_2_111/a_1020_375# 0.001512f
C11872 _052_ vdd 0.264744f
C11873 FILLER_0_5_128/a_124_375# _163_ 0.009765f
C11874 _114_ cal_count\[3\] 0.081644f
C11875 vdd _202_/a_36_160# 0.06338f
C11876 net61 _419_/a_1000_472# 0.017712f
C11877 net60 _419_/a_1308_423# 0.029697f
C11878 FILLER_0_4_177/a_36_472# net76 0.003007f
C11879 _111_ net36 0.102444f
C11880 _412_/a_2248_156# cal_itt\[1\] 0.005868f
C11881 FILLER_0_17_104/a_1468_375# vdd 0.022331f
C11882 output9/a_224_472# net19 0.070689f
C11883 _013_ FILLER_0_18_37/a_1468_375# 0.017213f
C11884 _431_/a_2665_112# FILLER_0_16_154/a_124_375# 0.006271f
C11885 FILLER_0_5_212/a_124_375# FILLER_0_4_213/a_36_472# 0.001723f
C11886 _175_ cal_count\[1\] 0.203153f
C11887 net62 FILLER_0_14_263/a_124_375# 0.037111f
C11888 _161_ _060_ 0.042838f
C11889 FILLER_0_16_89/a_572_375# _451_/a_448_472# 0.001597f
C11890 _025_ vdd 0.259346f
C11891 net54 _354_/a_257_69# 0.001135f
C11892 ctlp[1] FILLER_0_21_286/a_36_472# 0.014043f
C11893 _053_ _257_/a_36_472# 0.00507f
C11894 _188_ _039_ 0.002071f
C11895 _112_ net1 0.001653f
C11896 net34 output35/a_224_472# 0.0731f
C11897 _322_/a_124_24# _125_ 0.01165f
C11898 net78 net18 1.351707f
C11899 _440_/a_796_472# _029_ 0.009261f
C11900 _269_/a_36_472# vdd 0.03432f
C11901 _174_ net74 0.00916f
C11902 _119_ _359_/a_36_488# 0.003263f
C11903 net28 _426_/a_448_472# 0.00154f
C11904 _142_ net73 0.090025f
C11905 net40 _167_ 0.020177f
C11906 net16 FILLER_0_8_37/a_572_375# 0.004285f
C11907 net63 _434_/a_2560_156# 0.014333f
C11908 _015_ vss 0.090048f
C11909 net73 mask\[9\] 0.383862f
C11910 FILLER_0_15_116/a_572_375# net36 0.007321f
C11911 FILLER_0_2_111/a_124_375# _157_ 0.028285f
C11912 net39 _445_/a_2248_156# 0.003571f
C11913 FILLER_0_5_72/a_932_472# trim_mask\[1\] 0.014619f
C11914 mask\[2\] FILLER_0_15_212/a_36_472# 0.001181f
C11915 FILLER_0_12_136/a_124_375# _126_ 0.013041f
C11916 _428_/a_36_151# FILLER_0_13_100/a_124_375# 0.023595f
C11917 _038_ _120_ 0.00117f
C11918 _036_ _030_ 0.430683f
C11919 _247_/a_36_160# net22 0.048614f
C11920 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1468_375# 0.086742f
C11921 _235_/a_67_603# net40 0.001273f
C11922 FILLER_0_4_99/a_124_375# net14 0.003714f
C11923 _086_ _061_ 0.152228f
C11924 FILLER_0_20_193/a_124_375# vdd 0.009092f
C11925 _242_/a_36_160# _066_ 0.044262f
C11926 _176_ _451_/a_448_472# 0.007191f
C11927 FILLER_0_17_72/a_484_472# _131_ 0.002672f
C11928 FILLER_0_4_177/a_36_472# FILLER_0_2_177/a_124_375# 0.001512f
C11929 _081_ _001_ 0.012101f
C11930 trim[0] output41/a_224_472# 0.018464f
C11931 net16 _166_ 0.146913f
C11932 _079_ FILLER_0_5_206/a_124_375# 0.009128f
C11933 _086_ _311_/a_66_473# 0.007295f
C11934 _420_/a_36_151# _009_ 0.018171f
C11935 mask\[7\] _436_/a_2248_156# 0.003615f
C11936 output12/a_224_472# ctln[4] 0.041517f
C11937 _413_/a_36_151# FILLER_0_3_172/a_1468_375# 0.001252f
C11938 FILLER_0_15_116/a_36_472# net70 0.051129f
C11939 _116_ _161_ 0.008003f
C11940 FILLER_0_23_274/a_36_472# vss 0.002346f
C11941 fanout61/a_36_113# vdd 0.108255f
C11942 net26 _423_/a_1204_472# 0.001069f
C11943 net31 _102_ 0.060034f
C11944 net64 FILLER_0_9_282/a_484_472# 0.005717f
C11945 FILLER_0_5_212/a_124_375# net37 0.005414f
C11946 _432_/a_36_151# _137_ 0.051293f
C11947 FILLER_0_16_107/a_124_375# net36 0.001706f
C11948 _032_ trim_mask\[4\] 0.010578f
C11949 FILLER_0_5_54/a_1020_375# vss 0.003196f
C11950 FILLER_0_5_54/a_1468_375# vdd 0.014683f
C11951 net23 _242_/a_36_160# 0.007466f
C11952 FILLER_0_17_72/a_1916_375# net36 0.015395f
C11953 output42/a_224_472# vdd 0.04917f
C11954 FILLER_0_7_104/a_572_375# _154_ 0.020664f
C11955 _442_/a_1204_472# vdd 0.001128f
C11956 net16 _185_ 0.086347f
C11957 FILLER_0_21_125/a_124_375# _140_ 0.031374f
C11958 net34 _435_/a_2248_156# 0.01519f
C11959 FILLER_0_9_28/a_2276_472# net68 0.023299f
C11960 trim_val\[4\] trim_mask\[4\] 0.152123f
C11961 trim_val\[4\] net47 0.003977f
C11962 _126_ net14 0.238336f
C11963 FILLER_0_18_177/a_1020_375# vdd 0.040478f
C11964 FILLER_0_16_241/a_124_375# vdd 0.035603f
C11965 _449_/a_796_472# _067_ 0.004874f
C11966 net79 FILLER_0_11_282/a_36_472# 0.004358f
C11967 FILLER_0_12_20/a_36_472# vdd 0.068477f
C11968 FILLER_0_12_20/a_572_375# vss 0.054934f
C11969 _086_ _072_ 0.220767f
C11970 _450_/a_36_151# _039_ 0.018559f
C11971 _161_ _118_ 0.023939f
C11972 output13/a_224_472# trim_val\[4\] 0.001014f
C11973 _095_ _406_/a_36_159# 0.131137f
C11974 _132_ net70 0.534228f
C11975 _095_ FILLER_0_15_72/a_124_375# 0.001474f
C11976 FILLER_0_18_2/a_484_472# trimb[1] 0.009245f
C11977 _431_/a_1308_423# vss 0.003472f
C11978 net23 FILLER_0_16_154/a_36_472# 0.035678f
C11979 net20 FILLER_0_16_241/a_124_375# 0.002327f
C11980 net17 FILLER_0_20_15/a_124_375# 0.005919f
C11981 _370_/a_124_24# vdd 0.018613f
C11982 _410_/a_244_472# _042_ 0.003902f
C11983 _129_ _118_ 0.213736f
C11984 _352_/a_49_472# FILLER_0_22_128/a_36_472# 0.063744f
C11985 mask\[7\] FILLER_0_22_128/a_1020_375# 0.035799f
C11986 net72 FILLER_0_20_31/a_36_472# 0.002751f
C11987 _165_ vdd 0.168803f
C11988 FILLER_0_7_146/a_124_375# _059_ 0.029514f
C11989 net63 FILLER_0_20_193/a_36_472# 0.048818f
C11990 net70 _427_/a_36_151# 0.029237f
C11991 _439_/a_2560_156# vss 0.001309f
C11992 fanout53/a_36_160# _427_/a_2248_156# 0.027388f
C11993 FILLER_0_5_117/a_36_472# _163_ 0.007418f
C11994 _350_/a_49_472# _208_/a_36_160# 0.078981f
C11995 _444_/a_2665_112# FILLER_0_8_37/a_484_472# 0.001167f
C11996 _428_/a_796_472# _043_ 0.007935f
C11997 FILLER_0_21_28/a_2276_472# _424_/a_36_151# 0.001723f
C11998 net29 result[2] 0.001786f
C11999 FILLER_0_9_223/a_36_472# _070_ 0.006158f
C12000 _247_/a_36_160# vdd 0.060423f
C12001 _126_ _428_/a_36_151# 0.032026f
C12002 _130_ cal_count\[3\] 0.037708f
C12003 net74 _032_ 0.208799f
C12004 mask\[3\] FILLER_0_16_154/a_932_472# 0.002604f
C12005 _002_ FILLER_0_3_172/a_2276_472# 0.030358f
C12006 mask\[4\] net56 0.006006f
C12007 _341_/a_49_472# _141_ 0.006222f
C12008 _428_/a_448_472# _095_ 0.008804f
C12009 _443_/a_1000_472# _170_ 0.012879f
C12010 _061_ _090_ 0.00832f
C12011 _056_ _060_ 0.085489f
C12012 net15 _440_/a_448_472# 0.036624f
C12013 _077_ FILLER_0_9_72/a_932_472# 0.006408f
C12014 _119_ FILLER_0_8_156/a_572_375# 0.01739f
C12015 state\[2\] FILLER_0_13_142/a_1020_375# 0.007311f
C12016 net16 _407_/a_36_472# 0.027354f
C12017 net53 FILLER_0_13_142/a_36_472# 0.059367f
C12018 _414_/a_1308_423# net21 0.06986f
C12019 comp FILLER_0_12_2/a_36_472# 0.003875f
C12020 net16 cal_count\[0\] 0.152321f
C12021 FILLER_0_19_55/a_124_375# FILLER_0_17_56/a_36_472# 0.001338f
C12022 FILLER_0_21_133/a_36_472# _140_ 0.008378f
C12023 _142_ net56 0.028797f
C12024 result[6] _010_ 0.056004f
C12025 FILLER_0_24_274/a_36_472# vdd 0.107635f
C12026 FILLER_0_24_274/a_1468_375# vss 0.060201f
C12027 _062_ _160_ 0.001024f
C12028 FILLER_0_15_142/a_124_375# net23 0.002212f
C12029 _448_/a_2665_112# _170_ 0.002715f
C12030 _448_/a_1204_472# _037_ 0.008883f
C12031 net63 FILLER_0_18_177/a_1916_375# 0.040551f
C12032 FILLER_0_12_28/a_36_472# vdd 0.095598f
C12033 FILLER_0_12_28/a_124_375# vss 0.013117f
C12034 _430_/a_36_151# net22 0.005321f
C12035 ctln[2] rstn 0.017812f
C12036 _326_/a_36_160# _062_ 0.007797f
C12037 vdd net40 1.984115f
C12038 _437_/a_2665_112# _436_/a_36_151# 0.001466f
C12039 FILLER_0_22_128/a_1916_375# vss 0.018094f
C12040 FILLER_0_22_128/a_2364_375# vdd 0.015888f
C12041 output22/a_224_472# _435_/a_36_151# 0.12978f
C12042 fanout66/a_36_113# _029_ 0.001684f
C12043 _077_ _453_/a_2560_156# 0.001286f
C12044 net71 FILLER_0_22_107/a_572_375# 0.006403f
C12045 _284_/a_224_472# _094_ 0.001731f
C12046 _091_ net63 0.767908f
C12047 FILLER_0_3_78/a_124_375# _168_ 0.009374f
C12048 _315_/a_36_68# vss 0.02467f
C12049 net20 FILLER_0_24_274/a_36_472# 0.009746f
C12050 _126_ FILLER_0_11_109/a_36_472# 0.00136f
C12051 FILLER_0_16_73/a_36_472# _176_ 0.013449f
C12052 FILLER_0_6_79/a_124_375# vdd 0.015119f
C12053 _084_ vss 0.082779f
C12054 _098_ FILLER_0_21_206/a_124_375# 0.001882f
C12055 _093_ vss 2.002012f
C12056 _420_/a_36_151# FILLER_0_23_290/a_36_472# 0.001723f
C12057 FILLER_0_18_139/a_1380_472# net23 0.013087f
C12058 _053_ FILLER_0_6_47/a_124_375# 0.002541f
C12059 result[7] vdd 0.500292f
C12060 net82 FILLER_0_3_172/a_572_375# 0.010972f
C12061 _095_ _281_/a_234_472# 0.001467f
C12062 _035_ vss 0.105648f
C12063 FILLER_0_21_206/a_124_375# _205_/a_36_160# 0.03126f
C12064 FILLER_0_15_212/a_36_472# FILLER_0_15_205/a_124_375# 0.012267f
C12065 _136_ _018_ 0.002892f
C12066 _292_/a_36_160# _098_ 0.048643f
C12067 ctln[1] rstn 0.62944f
C12068 _093_ FILLER_0_18_107/a_1020_375# 0.006376f
C12069 FILLER_0_15_282/a_572_375# vss 0.058168f
C12070 FILLER_0_15_282/a_36_472# vdd 0.10628f
C12071 _120_ FILLER_0_9_72/a_932_472# 0.001709f
C12072 FILLER_0_17_38/a_572_375# vdd 0.01525f
C12073 _072_ _090_ 0.091468f
C12074 net79 net22 0.042486f
C12075 _032_ _159_ 0.053405f
C12076 net65 _425_/a_2248_156# 0.003451f
C12077 _173_ _450_/a_3129_107# 0.00264f
C12078 net81 fanout82/a_36_113# 0.061162f
C12079 _308_/a_848_380# _077_ 0.010515f
C12080 _198_/a_67_603# vdd 0.015843f
C12081 net48 _305_/a_36_159# 0.059079f
C12082 _116_ _056_ 0.30649f
C12083 _292_/a_36_160# _205_/a_36_160# 0.105676f
C12084 net20 result[7] 0.134149f
C12085 net73 _022_ 0.003246f
C12086 FILLER_0_17_72/a_3172_472# FILLER_0_17_104/a_36_472# 0.013277f
C12087 _276_/a_36_160# FILLER_0_18_209/a_484_472# 0.003913f
C12088 net36 net21 0.034415f
C12089 _086_ _331_/a_244_472# 0.001991f
C12090 _155_ _365_/a_36_68# 0.053708f
C12091 _115_ FILLER_0_9_105/a_124_375# 0.002316f
C12092 FILLER_0_6_47/a_3172_472# vss 0.014726f
C12093 net20 _198_/a_67_603# 0.013603f
C12094 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_572_375# 0.007947f
C12095 FILLER_0_4_197/a_1468_375# net59 0.050218f
C12096 net52 FILLER_0_6_47/a_2364_375# 0.002577f
C12097 _141_ _346_/a_257_69# 0.002092f
C12098 _070_ FILLER_0_5_136/a_36_472# 0.029293f
C12099 net57 FILLER_0_13_100/a_36_472# 0.077963f
C12100 FILLER_0_0_266/a_36_472# rstn 0.006108f
C12101 FILLER_0_3_142/a_124_375# _032_ 0.001153f
C12102 fanout71/a_36_113# _098_ 0.012725f
C12103 net32 _421_/a_2665_112# 0.019532f
C12104 _339_/a_36_160# _140_ 0.025058f
C12105 _020_ _334_/a_36_160# 0.028435f
C12106 FILLER_0_12_2/a_124_375# clkc 0.003601f
C12107 net33 _108_ 0.001901f
C12108 net39 _034_ 0.004367f
C12109 _032_ _442_/a_448_472# 0.001977f
C12110 _443_/a_448_472# _031_ 0.001143f
C12111 _443_/a_796_472# net69 0.020234f
C12112 net58 en 0.029072f
C12113 _056_ _118_ 0.028015f
C12114 net63 net33 0.048496f
C12115 net19 net33 0.254336f
C12116 net54 FILLER_0_22_107/a_124_375# 0.003502f
C12117 _405_/a_67_603# net17 0.014714f
C12118 _433_/a_36_151# _145_ 0.004437f
C12119 _430_/a_448_472# _019_ 0.019666f
C12120 _116_ _068_ 0.011673f
C12121 FILLER_0_10_247/a_124_375# net64 0.001597f
C12122 _176_ _070_ 0.467961f
C12123 _415_/a_36_151# vss 0.003124f
C12124 FILLER_0_4_99/a_124_375# _153_ 0.030839f
C12125 _236_/a_36_160# output39/a_224_472# 0.042231f
C12126 vss FILLER_0_5_148/a_484_472# 0.009015f
C12127 net32 ctlp[4] 0.001413f
C12128 _430_/a_36_151# vdd 0.112575f
C12129 _098_ FILLER_0_18_76/a_124_375# 0.001831f
C12130 FILLER_0_17_200/a_484_472# FILLER_0_18_177/a_3172_472# 0.026657f
C12131 net73 FILLER_0_18_107/a_484_472# 0.0052f
C12132 net29 FILLER_0_16_255/a_124_375# 0.085055f
C12133 FILLER_0_2_101/a_124_375# _156_ 0.022015f
C12134 net55 FILLER_0_17_72/a_1380_472# 0.021108f
C12135 _112_ net76 0.011948f
C12136 FILLER_0_12_20/a_484_472# _450_/a_448_472# 0.04564f
C12137 _422_/a_36_151# _010_ 0.006787f
C12138 _019_ mask\[2\] 0.155325f
C12139 FILLER_0_2_111/a_1380_472# vss 0.001679f
C12140 _260_/a_36_68# _080_ 0.001888f
C12141 FILLER_0_9_142/a_124_375# _122_ 0.004711f
C12142 net15 _394_/a_1936_472# 0.001592f
C12143 net41 _402_/a_56_567# 0.021641f
C12144 _445_/a_2248_156# net47 0.028909f
C12145 _440_/a_2665_112# vss 0.008703f
C12146 _029_ _365_/a_692_472# 0.001426f
C12147 _068_ _118_ 1.374452f
C12148 _070_ _124_ 0.114614f
C12149 trim_val\[2\] _381_/a_36_472# 0.005253f
C12150 _077_ _125_ 0.017422f
C12151 net16 net55 0.035875f
C12152 _219_/a_36_160# vss 0.00157f
C12153 net60 _421_/a_36_151# 0.224039f
C12154 _136_ vss 0.947188f
C12155 cal_count\[2\] cal_count\[1\] 0.067712f
C12156 FILLER_0_21_28/a_2724_472# _012_ 0.020109f
C12157 net55 _176_ 0.300149f
C12158 _128_ calibrate 0.039365f
C12159 FILLER_0_7_72/a_3172_472# net50 0.001428f
C12160 net4 _080_ 0.076128f
C12161 _017_ FILLER_0_14_107/a_484_472# 0.004583f
C12162 _144_ _354_/a_49_472# 0.03742f
C12163 net70 FILLER_0_14_107/a_1380_472# 0.003355f
C12164 net79 vdd 1.283563f
C12165 _114_ _267_/a_224_472# 0.001264f
C12166 net79 _192_/a_67_603# 0.017688f
C12167 state\[0\] _055_ 0.042917f
C12168 net81 _429_/a_448_472# 0.018517f
C12169 net62 vss 1.17087f
C12170 output47/a_224_472# net47 0.023797f
C12171 _303_/a_36_472# vdd 0.015964f
C12172 FILLER_0_1_266/a_36_472# net8 0.0138f
C12173 _386_/a_848_380# net22 0.00429f
C12174 _438_/a_1000_472# vss 0.001536f
C12175 net66 _440_/a_36_151# 0.041433f
C12176 FILLER_0_13_142/a_572_375# vdd 0.017472f
C12177 ctlp[1] _419_/a_2665_112# 0.009197f
C12178 FILLER_0_13_142/a_124_375# vss 0.009543f
C12179 ctln[1] _411_/a_1308_423# 0.037098f
C12180 _053_ _359_/a_36_488# 0.015831f
C12181 _257_/a_36_472# _070_ 0.002295f
C12182 _161_ _228_/a_36_68# 0.055774f
C12183 _374_/a_36_68# _062_ 0.004248f
C12184 _128_ net21 0.03068f
C12185 _077_ _251_/a_906_472# 0.001076f
C12186 FILLER_0_15_142/a_124_375# fanout73/a_36_113# 0.00146f
C12187 net20 net79 0.046876f
C12188 fanout82/a_36_113# net2 0.008681f
C12189 _199_/a_36_160# _046_ 0.017122f
C12190 _414_/a_796_472# cal_itt\[3\] 0.019699f
C12191 FILLER_0_3_204/a_36_472# net82 0.008268f
C12192 FILLER_0_5_72/a_1468_375# net49 0.001276f
C12193 _390_/a_244_472# _067_ 0.004031f
C12194 FILLER_0_1_98/a_36_472# _238_/a_67_603# 0.02529f
C12195 _308_/a_124_24# trim_mask\[0\] 0.018998f
C12196 net44 FILLER_0_15_2/a_572_375# 0.041552f
C12197 FILLER_0_15_2/a_36_472# vss 0.002136f
C12198 _431_/a_36_151# vss 0.00849f
C12199 net16 net17 0.034209f
C12200 _412_/a_796_472# net81 0.038712f
C12201 _412_/a_36_151# vss 0.003515f
C12202 _125_ _120_ 0.006198f
C12203 net68 FILLER_0_5_54/a_36_472# 0.012107f
C12204 net16 trim_val\[1\] 0.164715f
C12205 net15 FILLER_0_7_59/a_484_472# 0.015199f
C12206 mask\[4\] FILLER_0_18_177/a_484_472# 0.016924f
C12207 net15 _453_/a_36_151# 0.009841f
C12208 FILLER_0_16_255/a_36_472# _102_ 0.004641f
C12209 _414_/a_36_151# _072_ 0.033026f
C12210 net58 output27/a_224_472# 0.121438f
C12211 FILLER_0_18_171/a_124_375# _432_/a_36_151# 0.001597f
C12212 _447_/a_2248_156# net69 0.001126f
C12213 en clk 0.067072f
C12214 _133_ _062_ 1.210949f
C12215 _072_ FILLER_0_7_233/a_36_472# 0.00241f
C12216 FILLER_0_18_2/a_2364_375# _452_/a_1353_112# 0.001068f
C12217 FILLER_0_18_2/a_3260_375# _452_/a_36_151# 0.001597f
C12218 FILLER_0_18_2/a_572_375# _452_/a_3129_107# 0.001073f
C12219 _417_/a_1204_472# _006_ 0.014354f
C12220 FILLER_0_7_104/a_484_472# _131_ 0.00432f
C12221 net32 result[9] 0.001371f
C12222 net36 mask\[1\] 0.28584f
C12223 output27/a_224_472# calibrate 0.010614f
C12224 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_572_375# 0.026339f
C12225 _086_ _321_/a_3662_472# 0.002598f
C12226 _429_/a_2665_112# vss 0.012165f
C12227 output11/a_224_472# net65 0.001529f
C12228 _440_/a_2665_112# FILLER_0_5_88/a_124_375# 0.02132f
C12229 _367_/a_36_68# _154_ 0.028801f
C12230 FILLER_0_17_56/a_572_375# vss 0.05884f
C12231 FILLER_0_17_56/a_36_472# vdd 0.040007f
C12232 _442_/a_36_151# _371_/a_36_113# 0.001089f
C12233 _072_ _163_ 0.016226f
C12234 _148_ _436_/a_36_151# 0.032004f
C12235 input1/a_36_113# clk 0.001121f
C12236 _014_ FILLER_0_7_233/a_36_472# 0.002089f
C12237 _069_ _247_/a_36_160# 0.046764f
C12238 _422_/a_36_151# _299_/a_36_472# 0.004432f
C12239 _144_ net73 0.003657f
C12240 cal_count\[1\] _043_ 0.002223f
C12241 _316_/a_692_472# vdd 0.001634f
C12242 net79 _416_/a_1204_472# 0.006493f
C12243 _256_/a_36_68# _128_ 0.001702f
C12244 net55 FILLER_0_18_76/a_124_375# 0.001706f
C12245 FILLER_0_15_142/a_484_472# vss 0.029611f
C12246 net62 _416_/a_2248_156# 0.043158f
C12247 _093_ _027_ 0.047164f
C12248 vdd FILLER_0_13_290/a_124_375# 0.031436f
C12249 _424_/a_36_151# FILLER_0_18_37/a_572_375# 0.002807f
C12250 net20 _429_/a_2560_156# 0.002069f
C12251 FILLER_0_3_172/a_124_375# net59 0.001045f
C12252 _061_ _117_ 0.046662f
C12253 net53 vss 0.426484f
C12254 net26 _424_/a_1000_472# 0.003207f
C12255 _453_/a_448_472# _042_ 0.053209f
C12256 _453_/a_36_151# net51 0.012537f
C12257 result[8] FILLER_0_24_274/a_572_375# 0.00726f
C12258 net62 _195_/a_67_603# 0.002422f
C12259 FILLER_0_3_54/a_36_472# _160_ 0.00702f
C12260 _058_ FILLER_0_10_94/a_124_375# 0.001597f
C12261 _311_/a_66_473# _117_ 0.001055f
C12262 FILLER_0_20_177/a_124_375# FILLER_0_19_171/a_932_472# 0.001543f
C12263 _070_ _267_/a_36_472# 0.002617f
C12264 _386_/a_124_24# vss 0.009702f
C12265 _386_/a_848_380# vdd 0.054849f
C12266 net75 vdd 1.265616f
C12267 _260_/a_36_68# vss 0.030324f
C12268 _113_ _060_ 0.01991f
C12269 FILLER_0_19_171/a_572_375# vdd 0.022516f
C12270 FILLER_0_20_87/a_36_472# net14 0.001471f
C12271 output14/a_224_472# FILLER_0_0_130/a_124_375# 0.00515f
C12272 _085_ _121_ 0.027373f
C12273 FILLER_0_22_86/a_36_472# net71 0.005766f
C12274 net15 FILLER_0_13_72/a_572_375# 0.003021f
C12275 net15 fanout51/a_36_113# 0.001562f
C12276 _423_/a_2248_156# FILLER_0_23_60/a_124_375# 0.001901f
C12277 net58 _425_/a_2560_156# 0.004835f
C12278 fanout51/a_36_113# FILLER_0_11_78/a_36_472# 0.193759f
C12279 _451_/a_1353_112# net14 0.041814f
C12280 fanout68/a_36_113# net66 0.042828f
C12281 FILLER_0_5_72/a_484_472# _164_ 0.003769f
C12282 FILLER_0_10_107/a_484_472# vss 0.00298f
C12283 _321_/a_358_69# _121_ 0.00135f
C12284 fanout60/a_36_160# net18 0.004124f
C12285 mask\[1\] FILLER_0_15_228/a_36_472# 0.02055f
C12286 net14 _160_ 0.034023f
C12287 _088_ FILLER_0_4_213/a_124_375# 0.016013f
C12288 FILLER_0_7_72/a_2276_472# net14 0.004375f
C12289 _452_/a_1040_527# vdd 0.004153f
C12290 net20 net75 0.092951f
C12291 _242_/a_36_160# FILLER_0_5_148/a_572_375# 0.00805f
C12292 net63 net35 0.126544f
C12293 _346_/a_49_472# vdd -0.002208f
C12294 net55 _041_ 0.972122f
C12295 _089_ vdd 0.087336f
C12296 net4 vss 0.774455f
C12297 FILLER_0_18_177/a_2724_472# net21 0.048803f
C12298 FILLER_0_19_125/a_124_375# _022_ 0.055527f
C12299 net58 _416_/a_36_151# 0.001558f
C12300 _075_ _414_/a_2560_156# 0.026328f
C12301 _164_ _160_ 1.863027f
C12302 _425_/a_2560_156# calibrate 0.010842f
C12303 _376_/a_36_160# FILLER_0_5_88/a_36_472# 0.001448f
C12304 _016_ _126_ 0.051451f
C12305 _004_ vdd 0.448886f
C12306 _004_ _192_/a_67_603# 0.020219f
C12307 net15 net69 0.034091f
C12308 _308_/a_692_472# _115_ 0.001485f
C12309 _412_/a_796_472# net2 0.00566f
C12310 _406_/a_36_159# _185_ 0.001573f
C12311 _012_ FILLER_0_21_60/a_36_472# 0.017483f
C12312 net32 output32/a_224_472# 0.014826f
C12313 _440_/a_448_472# net47 0.016997f
C12314 FILLER_0_14_107/a_124_375# vss 0.002674f
C12315 result[5] vdd 0.142481f
C12316 FILLER_0_14_107/a_572_375# vdd 0.021509f
C12317 _305_/a_36_159# net37 0.015682f
C12318 FILLER_0_9_72/a_36_472# vss 0.0392f
C12319 FILLER_0_9_72/a_484_472# vdd 0.005654f
C12320 _056_ _228_/a_36_68# 0.043669f
C12321 _114_ FILLER_0_12_136/a_1020_375# 0.006974f
C12322 result[6] vss 0.310169f
C12323 _420_/a_36_151# FILLER_0_23_282/a_572_375# 0.059049f
C12324 mask\[5\] FILLER_0_20_193/a_484_472# 0.02147f
C12325 _389_/a_36_148# FILLER_0_10_94/a_124_375# 0.004673f
C12326 output10/a_224_472# _411_/a_2665_112# 0.008469f
C12327 net27 _415_/a_796_472# 0.004502f
C12328 _093_ FILLER_0_18_139/a_484_472# 0.008683f
C12329 fanout61/a_36_113# net77 0.052643f
C12330 net18 rstn 0.015842f
C12331 _010_ _419_/a_36_151# 0.002099f
C12332 _116_ _113_ 0.179616f
C12333 _289_/a_36_472# vdd 0.006886f
C12334 _095_ FILLER_0_14_123/a_36_472# 0.014431f
C12335 ctln[1] _411_/a_2560_156# 0.001413f
C12336 FILLER_0_5_72/a_1380_472# net47 0.003924f
C12337 _002_ _079_ 0.051048f
C12338 FILLER_0_19_187/a_36_472# _434_/a_36_151# 0.002398f
C12339 result[5] net20 0.045364f
C12340 fanout51/a_36_113# net51 0.013081f
C12341 output12/a_224_472# _413_/a_36_151# 0.006251f
C12342 _453_/a_2248_156# vss 0.031525f
C12343 _453_/a_2665_112# vdd 0.005481f
C12344 _127_ FILLER_0_11_142/a_484_472# 0.001177f
C12345 fanout68/a_36_113# FILLER_0_3_54/a_124_375# 0.015816f
C12346 _311_/a_1920_473# vdd 0.007492f
C12347 _015_ _426_/a_2248_156# 0.021465f
C12348 net17 _041_ 0.002779f
C12349 _053_ _372_/a_3662_472# 0.002006f
C12350 input2/a_36_113# en 0.002108f
C12351 net75 net9 0.006945f
C12352 FILLER_0_19_47/a_36_472# _424_/a_448_472# 0.004782f
C12353 FILLER_0_16_89/a_1380_472# _136_ 0.009079f
C12354 FILLER_0_18_2/a_124_375# net44 0.051228f
C12355 net63 FILLER_0_19_171/a_1468_375# 0.006671f
C12356 _087_ net37 0.23484f
C12357 net31 result[7] 0.231528f
C12358 net47 _034_ 0.052602f
C12359 net79 _283_/a_36_472# 0.010249f
C12360 net54 FILLER_0_22_86/a_1468_375# 0.001597f
C12361 output31/a_224_472# net62 0.030092f
C12362 FILLER_0_18_2/a_2724_472# net55 0.007511f
C12363 _136_ FILLER_0_16_154/a_1020_375# 0.004387f
C12364 _098_ _437_/a_2560_156# 0.001174f
C12365 fanout49/a_36_160# _030_ 0.017759f
C12366 FILLER_0_9_28/a_3260_375# vdd 0.017581f
C12367 mask\[5\] FILLER_0_18_177/a_2364_375# 0.002726f
C12368 FILLER_0_16_89/a_1020_375# _040_ 0.004252f
C12369 output35/a_224_472# output19/a_224_472# 0.015892f
C12370 _118_ _113_ 0.005092f
C12371 mask\[0\] _429_/a_1204_472# 0.005396f
C12372 _448_/a_2560_156# net59 0.007516f
C12373 vss _433_/a_1000_472# 0.002059f
C12374 _430_/a_36_151# _069_ 0.026308f
C12375 fanout69/a_36_113# FILLER_0_2_111/a_1468_375# 0.015816f
C12376 _027_ _438_/a_1000_472# 0.010911f
C12377 input1/a_36_113# input2/a_36_113# 0.029417f
C12378 FILLER_0_3_172/a_1916_375# net22 0.00941f
C12379 _111_ FILLER_0_18_76/a_124_375# 0.002494f
C12380 _029_ trim_mask\[1\] 1.002118f
C12381 FILLER_0_18_53/a_572_375# vss 0.057185f
C12382 FILLER_0_18_53/a_36_472# vdd 0.089087f
C12383 _077_ net68 0.003823f
C12384 _094_ _418_/a_796_472# 0.005889f
C12385 FILLER_0_17_133/a_124_375# vdd 0.010519f
C12386 input5/a_36_113# vdd 0.026855f
C12387 fanout76/a_36_160# net4 0.002206f
C12388 net54 _211_/a_36_160# 0.001244f
C12389 output22/a_224_472# net23 0.008048f
C12390 _052_ _424_/a_2665_112# 0.003027f
C12391 FILLER_0_16_57/a_36_472# _131_ 0.00864f
C12392 _121_ _062_ 0.001616f
C12393 _162_ FILLER_0_5_172/a_36_472# 0.001501f
C12394 net63 net22 0.223664f
C12395 _035_ output41/a_224_472# 0.002168f
C12396 fanout55/a_36_160# FILLER_0_13_80/a_124_375# 0.00805f
C12397 net55 FILLER_0_17_64/a_124_375# 0.020021f
C12398 ctlp[3] vdd 0.251098f
C12399 _445_/a_1308_423# net40 0.046345f
C12400 FILLER_0_7_104/a_932_472# _133_ 0.019721f
C12401 _131_ FILLER_0_11_109/a_124_375# 0.001048f
C12402 _017_ FILLER_0_13_100/a_124_375# 0.001274f
C12403 result[9] _420_/a_2665_112# 0.037019f
C12404 FILLER_0_10_28/a_124_375# vdd 0.039012f
C12405 net16 _408_/a_1336_472# 0.022364f
C12406 FILLER_0_18_2/a_2724_472# net17 0.017841f
C12407 trim[4] output42/a_224_472# 0.017153f
C12408 FILLER_0_9_105/a_124_375# vdd 0.029831f
C12409 _398_/a_36_113# _278_/a_36_160# 0.001636f
C12410 FILLER_0_13_142/a_1020_375# _043_ 0.005672f
C12411 FILLER_0_20_177/a_1468_375# vdd 0.016422f
C12412 _106_ _201_/a_67_603# 0.00327f
C12413 _069_ net79 0.045808f
C12414 net64 FILLER_0_14_235/a_36_472# 0.067888f
C12415 state\[0\] _426_/a_2665_112# 0.017088f
C12416 mask\[4\] _145_ 0.340415f
C12417 _343_/a_49_472# vss 0.002581f
C12418 _136_ _095_ 0.043768f
C12419 net35 _423_/a_2248_156# 0.003899f
C12420 mask\[8\] _423_/a_2665_112# 0.004281f
C12421 FILLER_0_17_226/a_124_375# FILLER_0_17_218/a_572_375# 0.012001f
C12422 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_124_375# 0.001597f
C12423 output48/a_224_472# en 0.003074f
C12424 net16 _447_/a_1308_423# 0.001178f
C12425 ctln[9] _447_/a_36_151# 0.010503f
C12426 ctln[1] cal_itt\[0\] 0.003349f
C12427 net15 _013_ 0.152142f
C12428 _398_/a_36_113# _178_ 0.004282f
C12429 net36 FILLER_0_15_212/a_124_375# 0.004391f
C12430 net56 net23 0.930833f
C12431 net36 _099_ 0.325141f
C12432 net70 FILLER_0_16_115/a_124_375# 0.025173f
C12433 FILLER_0_10_78/a_932_472# vss 0.002987f
C12434 _021_ mask\[4\] 0.018108f
C12435 net68 _120_ 0.001304f
C12436 _431_/a_448_472# FILLER_0_17_142/a_124_375# 0.006782f
C12437 _429_/a_36_151# FILLER_0_15_212/a_484_472# 0.001723f
C12438 FILLER_0_20_15/a_1468_375# vdd 0.009742f
C12439 mask\[3\] FILLER_0_17_226/a_36_472# 0.011509f
C12440 net81 _138_ 0.006815f
C12441 FILLER_0_1_98/a_124_375# ctln[7] 0.004533f
C12442 FILLER_0_4_107/a_124_375# _156_ 0.00268f
C12443 _321_/a_2590_472# _118_ 0.002396f
C12444 _422_/a_36_151# vss 0.014056f
C12445 _422_/a_448_472# vdd 0.032865f
C12446 net73 fanout73/a_36_113# 0.02062f
C12447 _168_ vdd 0.083621f
C12448 _008_ net30 1.112351f
C12449 _441_/a_1308_423# vss 0.016854f
C12450 _129_ net74 0.476969f
C12451 _031_ _369_/a_692_472# 0.00359f
C12452 _067_ FILLER_0_13_72/a_124_375# 0.001782f
C12453 vss _047_ 0.070755f
C12454 net55 _424_/a_1308_423# 0.00168f
C12455 _077_ net67 0.073924f
C12456 _064_ _446_/a_2248_156# 0.04774f
C12457 net52 FILLER_0_5_54/a_1380_472# 0.00179f
C12458 _413_/a_796_472# net65 0.006888f
C12459 trim_val\[1\] FILLER_0_6_47/a_124_375# 0.002577f
C12460 FILLER_0_21_133/a_36_472# FILLER_0_22_128/a_484_472# 0.026657f
C12461 _058_ FILLER_0_9_105/a_484_472# 0.00148f
C12462 FILLER_0_16_241/a_124_375# _282_/a_36_160# 0.005398f
C12463 FILLER_0_14_81/a_124_375# cal_count\[1\] 0.070473f
C12464 en_co_clk _067_ 0.272082f
C12465 FILLER_0_3_204/a_36_472# net21 0.01535f
C12466 _176_ FILLER_0_10_94/a_36_472# 0.009089f
C12467 _005_ _416_/a_2665_112# 0.014205f
C12468 result[7] net77 0.005269f
C12469 FILLER_0_18_139/a_572_375# FILLER_0_19_142/a_124_375# 0.026339f
C12470 net32 _094_ 0.027571f
C12471 _441_/a_1204_472# _168_ 0.009437f
C12472 _058_ vss 0.19427f
C12473 _077_ FILLER_0_11_64/a_36_472# 0.076102f
C12474 FILLER_0_13_212/a_36_472# FILLER_0_13_206/a_124_375# 0.016748f
C12475 FILLER_0_5_117/a_124_375# vdd 0.035079f
C12476 _131_ FILLER_0_17_104/a_124_375# 0.006681f
C12477 output35/a_224_472# mask\[6\] 0.069819f
C12478 FILLER_0_6_239/a_124_375# vdd 0.031271f
C12479 ctlp[1] _421_/a_1204_472# 0.003759f
C12480 net48 _001_ 0.006122f
C12481 FILLER_0_17_142/a_36_472# _137_ 0.003953f
C12482 fanout77/a_36_113# vss 0.004099f
C12483 FILLER_0_20_31/a_36_472# vdd 0.097195f
C12484 FILLER_0_20_31/a_124_375# vss 0.049142f
C12485 _155_ FILLER_0_6_90/a_484_472# 0.005297f
C12486 _444_/a_2248_156# FILLER_0_6_37/a_124_375# 0.001101f
C12487 _104_ _010_ 0.252687f
C12488 _144_ FILLER_0_19_125/a_124_375# 0.012834f
C12489 _028_ FILLER_0_6_79/a_36_472# 0.016281f
C12490 FILLER_0_3_172/a_1916_375# vdd -0.010166f
C12491 _359_/a_36_488# _070_ 0.028563f
C12492 _003_ net76 0.080782f
C12493 FILLER_0_15_290/a_36_472# output30/a_224_472# 0.001711f
C12494 result[6] _420_/a_796_472# 0.002296f
C12495 net63 FILLER_0_20_177/a_484_472# 0.002172f
C12496 FILLER_0_18_171/a_36_472# net80 0.041571f
C12497 _108_ vdd 0.298249f
C12498 net20 FILLER_0_6_239/a_124_375# 0.004897f
C12499 FILLER_0_9_28/a_3260_375# fanout67/a_36_160# 0.001925f
C12500 net16 FILLER_0_16_37/a_124_375# 0.033245f
C12501 net16 _444_/a_1308_423# 0.002172f
C12502 _170_ _066_ 0.189122f
C12503 output11/a_224_472# FILLER_0_0_232/a_124_375# 0.00515f
C12504 FILLER_0_15_142/a_124_375# net36 0.006533f
C12505 FILLER_0_4_123/a_36_472# trim_mask\[4\] 0.003692f
C12506 net63 vdd 1.002883f
C12507 net19 vdd 2.167778f
C12508 net28 net79 0.116857f
C12509 trim[4] net40 0.017911f
C12510 net16 FILLER_0_8_24/a_572_375# 0.002225f
C12511 net19 _192_/a_67_603# 0.003106f
C12512 _423_/a_36_151# FILLER_0_23_44/a_932_472# 0.001723f
C12513 _232_/a_67_603# net47 0.014888f
C12514 _415_/a_2560_156# net64 0.066438f
C12515 state\[2\] _043_ 0.028842f
C12516 _287_/a_36_472# _094_ 0.029751f
C12517 _098_ FILLER_0_15_212/a_1380_472# 0.009972f
C12518 output11/a_224_472# net11 0.003448f
C12519 FILLER_0_4_123/a_36_472# net47 0.012399f
C12520 output14/a_224_472# net52 0.02346f
C12521 _072_ net48 0.037795f
C12522 vss _416_/a_1308_423# 0.001962f
C12523 _274_/a_36_68# _091_ 0.025773f
C12524 _422_/a_796_472# _108_ 0.007356f
C12525 net20 _108_ 0.125627f
C12526 trim_mask\[1\] _163_ 0.166315f
C12527 _153_ _160_ 0.304792f
C12528 mask\[8\] _026_ 0.001638f
C12529 FILLER_0_15_142/a_484_472# _095_ 0.001509f
C12530 _126_ _017_ 0.071134f
C12531 net54 net71 0.536043f
C12532 net65 FILLER_0_2_171/a_124_375# 0.023202f
C12533 _188_ vdd 0.022839f
C12534 _281_/a_234_472# _098_ 0.003724f
C12535 _075_ _257_/a_36_472# 0.005709f
C12536 ctln[0] trim[2] 0.011834f
C12537 _175_ _043_ 0.001037f
C12538 FILLER_0_21_206/a_124_375# net21 0.035287f
C12539 _008_ _417_/a_36_151# 0.001136f
C12540 net63 net20 0.045207f
C12541 net20 net19 0.384932f
C12542 net76 net1 0.059026f
C12543 FILLER_0_11_64/a_36_472# _120_ 0.011673f
C12544 FILLER_0_11_64/a_36_472# _038_ 0.001822f
C12545 net46 FILLER_0_20_15/a_1020_375# 0.0302f
C12546 trimb[3] FILLER_0_20_15/a_124_375# 0.001391f
C12547 net53 _095_ 0.431214f
C12548 net13 _387_/a_36_113# 0.00189f
C12549 net23 _170_ 0.107532f
C12550 _098_ _434_/a_1204_472# 0.006257f
C12551 net48 _014_ 0.276733f
C12552 FILLER_0_14_91/a_36_472# _136_ 0.008573f
C12553 _389_/a_36_148# vss 0.001935f
C12554 net79 FILLER_0_12_236/a_572_375# 0.010684f
C12555 net7 vdd 0.321735f
C12556 _430_/a_2248_156# net63 0.051057f
C12557 _434_/a_448_472# _023_ 0.03093f
C12558 FILLER_0_4_49/a_572_375# net66 0.074393f
C12559 net55 _406_/a_36_159# 0.001219f
C12560 net16 trim_mask\[2\] 0.002527f
C12561 net32 net78 0.055231f
C12562 net52 FILLER_0_3_78/a_36_472# 0.034084f
C12563 _140_ FILLER_0_22_128/a_2364_375# 0.003037f
C12564 output28/a_224_472# FILLER_0_11_282/a_36_472# 0.008834f
C12565 net52 FILLER_0_2_127/a_36_472# 0.001964f
C12566 _435_/a_2248_156# mask\[6\] 0.001778f
C12567 _076_ net23 0.105196f
C12568 _028_ _077_ 0.017713f
C12569 _105_ _295_/a_36_472# 0.031356f
C12570 ctlp[7] _050_ 0.153673f
C12571 _030_ FILLER_0_3_78/a_484_472# 0.007736f
C12572 net49 FILLER_0_3_78/a_36_472# 0.059367f
C12573 FILLER_0_17_161/a_124_375# vdd 0.014253f
C12574 _055_ _311_/a_1212_473# 0.004259f
C12575 _432_/a_36_151# FILLER_0_16_154/a_1468_375# 0.001107f
C12576 _068_ net47 0.001491f
C12577 FILLER_0_12_124/a_36_472# _126_ 0.056268f
C12578 _009_ FILLER_0_23_290/a_36_472# 0.002345f
C12579 _291_/a_36_160# vss 0.012222f
C12580 cal input4/a_36_68# 0.054357f
C12581 _053_ FILLER_0_6_47/a_3172_472# 0.001777f
C12582 net57 _131_ 0.030577f
C12583 FILLER_0_15_150/a_124_375# net56 0.011873f
C12584 _412_/a_1204_472# net1 0.019647f
C12585 FILLER_0_4_123/a_36_472# net74 0.001578f
C12586 net19 net9 0.342451f
C12587 _412_/a_36_151# output37/a_224_472# 0.006358f
C12588 _074_ FILLER_0_5_172/a_36_472# 0.016713f
C12589 result[7] _421_/a_448_472# 0.018021f
C12590 state\[0\] _223_/a_36_160# 0.070065f
C12591 FILLER_0_3_172/a_2724_472# net65 0.001777f
C12592 FILLER_0_7_72/a_2276_472# _439_/a_2665_112# 0.001167f
C12593 output12/a_224_472# _448_/a_36_151# 0.069748f
C12594 _070_ _246_/a_36_68# 0.056186f
C12595 net79 net77 0.431572f
C12596 _420_/a_36_151# vdd 0.137919f
C12597 FILLER_0_20_107/a_36_472# _438_/a_2665_112# 0.035266f
C12598 _406_/a_36_159# net17 0.053547f
C12599 _095_ FILLER_0_14_107/a_124_375# 0.01418f
C12600 net4 FILLER_0_12_220/a_124_375# 0.016485f
C12601 _443_/a_2560_156# vss 0.002467f
C12602 FILLER_0_19_47/a_124_375# _052_ 0.019401f
C12603 _057_ _311_/a_254_473# 0.002364f
C12604 _228_/a_36_68# _113_ 0.021898f
C12605 _122_ _062_ 0.190871f
C12606 FILLER_0_19_28/a_572_375# vss 0.002775f
C12607 FILLER_0_19_28/a_36_472# vdd 0.052986f
C12608 trimb[1] FILLER_0_20_2/a_572_375# 0.003431f
C12609 _446_/a_1000_472# net66 0.006158f
C12610 vdd _450_/a_36_151# 0.08588f
C12611 cal_count\[3\] _373_/a_632_68# 0.004529f
C12612 _413_/a_2248_156# vss 0.004157f
C12613 trim_mask\[1\] FILLER_0_4_91/a_36_472# 0.26171f
C12614 _423_/a_2248_156# vdd 0.013707f
C12615 FILLER_0_16_57/a_932_472# net55 0.00179f
C12616 _115_ net50 0.008628f
C12617 ctlp[3] output20/a_224_472# 0.023589f
C12618 FILLER_0_14_181/a_36_472# _138_ 0.002748f
C12619 _062_ _227_/a_36_160# 0.015411f
C12620 FILLER_0_16_89/a_1468_375# vss 0.048986f
C12621 FILLER_0_16_89/a_36_472# vdd 0.040085f
C12622 trim_mask\[4\] net69 0.185121f
C12623 net57 net56 0.054294f
C12624 _022_ _145_ 0.199016f
C12625 _189_/a_67_603# _043_ 0.005635f
C12626 net75 cal_itt\[2\] 0.143064f
C12627 _081_ _066_ 0.061358f
C12628 net60 FILLER_0_17_282/a_36_472# 0.009978f
C12629 _214_/a_36_160# FILLER_0_23_88/a_36_472# 0.006647f
C12630 _077_ FILLER_0_6_231/a_36_472# 0.075292f
C12631 FILLER_0_4_123/a_36_472# _159_ 0.004956f
C12632 FILLER_0_14_91/a_36_472# net53 0.005849f
C12633 FILLER_0_4_49/a_124_375# _164_ 0.017213f
C12634 _440_/a_36_151# FILLER_0_6_47/a_2276_472# 0.001512f
C12635 _053_ _219_/a_36_160# 0.005244f
C12636 _181_ _402_/a_2172_497# 0.001555f
C12637 FILLER_0_17_72/a_2724_472# vdd 0.007064f
C12638 FILLER_0_17_72/a_2276_472# vss -0.001288f
C12639 FILLER_0_22_86/a_572_375# net14 0.009573f
C12640 _419_/a_448_472# vdd 0.022174f
C12641 _419_/a_36_151# vss -0.00139f
C12642 net35 net24 0.01339f
C12643 _132_ FILLER_0_18_107/a_932_472# 0.001369f
C12644 _402_/a_56_567# _452_/a_36_151# 0.001915f
C12645 _004_ net28 0.082388f
C12646 net43 net40 0.018193f
C12647 _035_ _166_ 0.034749f
C12648 FILLER_0_4_107/a_932_472# _158_ 0.029116f
C12649 _119_ _058_ 0.692466f
C12650 ctln[5] _448_/a_796_472# 0.001484f
C12651 _081_ net23 0.081773f
C12652 FILLER_0_4_123/a_36_472# _154_ 0.001043f
C12653 FILLER_0_6_239/a_36_472# net76 0.011803f
C12654 output20/a_224_472# _422_/a_448_472# 0.009204f
C12655 _427_/a_2560_156# vss 0.003576f
C12656 trim_mask\[4\] _152_ 0.224909f
C12657 ctln[2] en 0.001355f
C12658 net19 _420_/a_1308_423# 0.010051f
C12659 FILLER_0_13_142/a_1468_375# _225_/a_36_160# 0.027706f
C12660 FILLER_0_5_172/a_36_472# FILLER_0_5_164/a_484_472# 0.013276f
C12661 _372_/a_2590_472# _076_ 0.002268f
C12662 ctln[9] vss 0.167242f
C12663 net74 FILLER_0_13_72/a_572_375# 0.012891f
C12664 net20 _419_/a_448_472# 0.025583f
C12665 _269_/a_36_472# _083_ 0.015096f
C12666 _152_ net47 0.242864f
C12667 output42/a_224_472# FILLER_0_8_2/a_124_375# 0.030009f
C12668 trim_val\[4\] FILLER_0_3_172/a_124_375# 0.002076f
C12669 FILLER_0_1_204/a_36_472# net59 0.067975f
C12670 _086_ net23 0.037804f
C12671 net60 _010_ 0.108311f
C12672 mask\[3\] FILLER_0_18_177/a_1380_472# 0.005654f
C12673 FILLER_0_9_28/a_36_472# output42/a_224_472# 0.010684f
C12674 _072_ FILLER_0_12_220/a_36_472# 0.01861f
C12675 FILLER_0_22_128/a_2364_375# FILLER_0_21_150/a_36_472# 0.001543f
C12676 net4 FILLER_0_12_236/a_36_472# 0.016315f
C12677 _272_/a_36_472# net37 0.002669f
C12678 ctln[6] output14/a_224_472# 0.007421f
C12679 FILLER_0_6_90/a_36_472# _163_ 0.016147f
C12680 _186_ vdd 0.074983f
C12681 net61 ctlp[2] 0.022612f
C12682 net66 _029_ 0.056971f
C12683 net58 _426_/a_36_151# 0.002612f
C12684 _369_/a_692_472# _157_ 0.0025f
C12685 FILLER_0_4_49/a_36_472# net47 0.002964f
C12686 mask\[7\] _435_/a_1308_423# 0.028235f
C12687 _394_/a_728_93# cal_count\[1\] 0.057049f
C12688 mask\[3\] FILLER_0_17_218/a_124_375# 0.016168f
C12689 net74 net69 0.143604f
C12690 _155_ net14 0.10433f
C12691 FILLER_0_8_263/a_124_375# FILLER_0_8_247/a_1468_375# 0.012001f
C12692 net22 FILLER_0_18_209/a_36_472# 0.018061f
C12693 _053_ FILLER_0_6_177/a_484_472# 0.015994f
C12694 FILLER_0_8_107/a_36_472# FILLER_0_7_104/a_484_472# 0.026657f
C12695 mask\[5\] FILLER_0_19_171/a_36_472# 0.002923f
C12696 output20/a_224_472# _108_ 0.022243f
C12697 _149_ vss 0.005314f
C12698 FILLER_0_2_171/a_36_472# net59 0.066486f
C12699 FILLER_0_3_2/a_124_375# _446_/a_36_151# 0.023595f
C12700 net23 FILLER_0_22_128/a_1828_472# 0.003857f
C12701 _213_/a_67_603# _051_ 0.015959f
C12702 _426_/a_36_151# calibrate 0.004525f
C12703 FILLER_0_18_139/a_1020_375# vdd 0.001285f
C12704 FILLER_0_18_139/a_572_375# vss 0.009977f
C12705 mask\[0\] FILLER_0_14_235/a_484_472# 0.004688f
C12706 _335_/a_49_472# _098_ 0.001047f
C12707 result[2] FILLER_0_13_290/a_36_472# 0.016496f
C12708 output36/a_224_472# FILLER_0_15_282/a_124_375# 0.002977f
C12709 result[1] _005_ 0.001478f
C12710 _411_/a_1308_423# net65 0.004122f
C12711 net57 _170_ 0.057355f
C12712 _408_/a_56_524# _067_ 0.003678f
C12713 FILLER_0_14_181/a_36_472# _113_ 0.004214f
C12714 FILLER_0_9_72/a_1468_375# _439_/a_36_151# 0.005577f
C12715 net78 _420_/a_2665_112# 0.039469f
C12716 ctln[1] input1/a_36_113# 0.004419f
C12717 FILLER_0_5_148/a_36_472# _160_ 0.001025f
C12718 FILLER_0_15_282/a_36_472# output30/a_224_472# 0.001711f
C12719 FILLER_0_15_282/a_124_375# net30 0.00123f
C12720 FILLER_0_3_172/a_1020_375# FILLER_0_2_177/a_484_472# 0.001723f
C12721 FILLER_0_12_28/a_124_375# cal_count\[0\] 0.001414f
C12722 FILLER_0_0_130/a_36_472# vss 0.00351f
C12723 FILLER_0_10_256/a_124_375# _426_/a_36_151# 0.001597f
C12724 cal_count\[3\] _055_ 0.039546f
C12725 FILLER_0_18_177/a_2812_375# _202_/a_36_160# 0.026361f
C12726 FILLER_0_4_144/a_36_472# _370_/a_848_380# 0.15783f
C12727 _412_/a_796_472# cal_itt\[1\] 0.004226f
C12728 net57 _074_ 0.026184f
C12729 FILLER_0_14_81/a_124_375# _175_ 0.005719f
C12730 _064_ net39 0.558387f
C12731 net74 _152_ 1.007413f
C12732 _430_/a_2665_112# vss 0.031646f
C12733 _016_ _428_/a_2560_156# 0.003934f
C12734 FILLER_0_12_136/a_1020_375# FILLER_0_13_142/a_484_472# 0.001684f
C12735 net67 _221_/a_36_160# 0.008581f
C12736 result[5] net77 0.142532f
C12737 FILLER_0_1_204/a_124_375# net11 0.01048f
C12738 net75 _426_/a_1204_472# 0.001592f
C12739 input3/a_36_113# cal_count\[2\] 0.00555f
C12740 FILLER_0_18_2/a_3260_375# _041_ 0.001024f
C12741 result[0] fanout65/a_36_113# 0.001816f
C12742 net57 _076_ 0.028356f
C12743 _435_/a_1204_472# vdd 0.013805f
C12744 _028_ _363_/a_36_68# 0.015609f
C12745 net38 _444_/a_1000_472# 0.027886f
C12746 _136_ _451_/a_448_472# 0.047841f
C12747 net63 _069_ 0.04528f
C12748 FILLER_0_17_72/a_572_375# FILLER_0_15_72/a_484_472# 0.001512f
C12749 FILLER_0_13_212/a_36_472# _429_/a_1308_423# 0.009119f
C12750 _013_ _012_ 0.003113f
C12751 net38 FILLER_0_8_24/a_484_472# 0.001223f
C12752 _189_/a_67_603# FILLER_0_12_236/a_124_375# 0.00221f
C12753 _103_ _418_/a_2665_112# 0.0066f
C12754 net69 _159_ 0.010086f
C12755 _063_ _167_ 0.002201f
C12756 _413_/a_1000_472# net59 0.018099f
C12757 _443_/a_448_472# net23 0.038188f
C12758 FILLER_0_5_128/a_572_375# _133_ 0.00134f
C12759 FILLER_0_8_2/a_124_375# net40 0.002839f
C12760 output28/a_224_472# vdd 0.044767f
C12761 FILLER_0_18_76/a_36_472# vss 0.007456f
C12762 net73 net36 0.073334f
C12763 ctln[5] net59 0.030363f
C12764 FILLER_0_15_150/a_36_472# _136_ 0.002967f
C12765 _093_ _098_ 0.556613f
C12766 _126_ cal_count\[3\] 0.418508f
C12767 FILLER_0_9_28/a_36_472# net40 0.020589f
C12768 _134_ FILLER_0_9_105/a_484_472# 0.011499f
C12769 _292_/a_36_160# _105_ 0.027405f
C12770 net27 FILLER_0_10_247/a_36_472# 0.016681f
C12771 _372_/a_2034_472# _152_ 0.00171f
C12772 ctln[5] FILLER_0_0_198/a_124_375# 0.002726f
C12773 net34 _299_/a_36_472# 0.003396f
C12774 _077_ FILLER_0_7_72/a_484_472# 0.001332f
C12775 FILLER_0_10_37/a_36_472# _453_/a_36_151# 0.003462f
C12776 _099_ FILLER_0_14_235/a_484_472# 0.00281f
C12777 FILLER_0_21_125/a_572_375# vss 0.054783f
C12778 FILLER_0_21_125/a_36_472# vdd 0.007233f
C12779 net41 _446_/a_1000_472# 0.01097f
C12780 FILLER_0_4_107/a_36_472# trim_mask\[3\] 0.00152f
C12781 _134_ vss 0.088213f
C12782 _008_ _046_ 0.067769f
C12783 _137_ FILLER_0_17_104/a_1468_375# 0.002679f
C12784 _176_ _171_ 0.049997f
C12785 _077_ FILLER_0_12_50/a_124_375# 0.008485f
C12786 net69 _154_ 0.05211f
C12787 FILLER_0_20_193/a_36_472# FILLER_0_18_177/a_1916_375# 0.0027f
C12788 net54 FILLER_0_18_107/a_3260_375# 0.001619f
C12789 _042_ net51 0.026776f
C12790 output34/a_224_472# _102_ 0.008577f
C12791 FILLER_0_6_90/a_484_472# FILLER_0_4_91/a_572_375# 0.00108f
C12792 FILLER_0_11_64/a_124_375# vdd 0.045435f
C12793 _053_ net4 0.013559f
C12794 net57 en_co_clk 0.195533f
C12795 _104_ vss 0.564464f
C12796 _132_ _428_/a_36_151# 0.013691f
C12797 _159_ _152_ 0.035925f
C12798 _121_ FILLER_0_8_156/a_124_375# 0.033427f
C12799 net80 FILLER_0_19_171/a_36_472# 0.040915f
C12800 _442_/a_448_472# net69 0.004308f
C12801 _445_/a_36_151# vdd 0.052935f
C12802 net75 FILLER_0_6_231/a_484_472# 0.003485f
C12803 FILLER_0_21_28/a_3260_375# vss 0.054959f
C12804 FILLER_0_21_28/a_36_472# vdd 0.090954f
C12805 _144_ _145_ 0.671767f
C12806 FILLER_0_18_209/a_572_375# vss 0.007545f
C12807 FILLER_0_18_209/a_36_472# vdd 0.089327f
C12808 _320_/a_1792_472# _043_ 0.002235f
C12809 net52 FILLER_0_2_93/a_572_375# 0.007787f
C12810 fanout58/a_36_160# en 0.00568f
C12811 FILLER_0_7_162/a_124_375# _062_ 0.010242f
C12812 net31 net19 0.023019f
C12813 _126_ _320_/a_672_472# 0.003662f
C12814 _356_/a_36_472# net14 0.001801f
C12815 _346_/a_49_472# _140_ 0.003436f
C12816 net16 _179_ 0.007397f
C12817 FILLER_0_4_107/a_1380_472# trim_mask\[4\] 0.011766f
C12818 _074_ cal_itt\[0\] 0.076802f
C12819 net63 _435_/a_2665_112# 0.039512f
C12820 net36 _451_/a_1040_527# 0.00974f
C12821 _427_/a_448_472# net23 0.014853f
C12822 FILLER_0_3_142/a_36_472# _081_ 0.001386f
C12823 net76 FILLER_0_5_198/a_124_375# 0.006974f
C12824 FILLER_0_12_50/a_124_375# _120_ 0.002753f
C12825 FILLER_0_4_107/a_1380_472# net47 0.008874f
C12826 net79 output30/a_224_472# 0.078502f
C12827 fanout53/a_36_160# _136_ 0.001471f
C12828 _070_ _315_/a_36_68# 0.031892f
C12829 _132_ FILLER_0_11_109/a_36_472# 0.005748f
C12830 net38 output39/a_224_472# 0.036027f
C12831 net28 net19 0.115252f
C12832 _115_ _322_/a_848_380# 0.011372f
C12833 FILLER_0_20_107/a_124_375# vss 0.002749f
C12834 FILLER_0_20_107/a_36_472# vdd 0.117841f
C12835 mask\[5\] FILLER_0_20_177/a_932_472# 0.016114f
C12836 FILLER_0_12_20/a_572_375# net17 0.041149f
C12837 net23 _145_ 0.035734f
C12838 trim_mask\[2\] _030_ 1.467465f
C12839 _412_/a_1204_472# net76 0.020975f
C12840 net76 FILLER_0_2_177/a_124_375# 0.00439f
C12841 _428_/a_2665_112# FILLER_0_13_142/a_124_375# 0.003325f
C12842 result[1] _416_/a_448_472# 0.008784f
C12843 _104_ _107_ 0.021508f
C12844 _009_ FILLER_0_23_282/a_572_375# 0.016879f
C12845 net24 vdd 0.223761f
C12846 net14 FILLER_0_10_94/a_484_472# 0.020589f
C12847 mask\[5\] vss 0.528441f
C12848 _131_ net36 0.068899f
C12849 net57 _081_ 0.023513f
C12850 FILLER_0_18_2/a_484_472# net38 0.003391f
C12851 net53 _451_/a_448_472# 0.026909f
C12852 net70 _451_/a_836_156# 0.006451f
C12853 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_124_375# 0.026339f
C12854 result[6] _421_/a_1308_423# 0.023269f
C12855 FILLER_0_15_142/a_484_472# FILLER_0_15_150/a_36_472# 0.013277f
C12856 _114_ FILLER_0_13_142/a_572_375# 0.00191f
C12857 _408_/a_244_524# net47 0.001066f
C12858 _425_/a_2248_156# net37 0.01491f
C12859 _086_ net57 0.126563f
C12860 FILLER_0_16_107/a_484_472# _131_ 0.008223f
C12861 _274_/a_1164_497# net64 0.002049f
C12862 FILLER_0_15_150/a_36_472# net53 0.016925f
C12863 net58 FILLER_0_8_247/a_1380_472# 0.0597f
C12864 FILLER_0_4_197/a_484_472# net21 0.046864f
C12865 _413_/a_2665_112# net65 0.033675f
C12866 _012_ net71 0.004946f
C12867 _136_ _098_ 0.049635f
C12868 _414_/a_796_472# vdd 0.001497f
C12869 result[0] FILLER_0_9_290/a_124_375# 0.030628f
C12870 net61 _418_/a_448_472# 0.001253f
C12871 net29 vss 0.259409f
C12872 output39/a_224_472# net66 0.009679f
C12873 _093_ net55 0.182194f
C12874 _314_/a_224_472# net23 0.001238f
C12875 FILLER_0_10_78/a_572_375# FILLER_0_11_78/a_572_375# 0.05841f
C12876 _426_/a_796_472# vdd 0.007178f
C12877 _098_ _438_/a_1000_472# 0.001492f
C12878 FILLER_0_8_247/a_1380_472# calibrate 0.008605f
C12879 FILLER_0_12_220/a_484_472# _060_ 0.003379f
C12880 FILLER_0_7_72/a_1468_375# net50 0.020186f
C12881 _065_ _447_/a_2248_156# 0.038629f
C12882 fanout49/a_36_160# _440_/a_2665_112# 0.00631f
C12883 FILLER_0_16_107/a_572_375# net70 0.002193f
C12884 _008_ result[4] 0.134001f
C12885 _063_ vdd 0.201806f
C12886 mask\[5\] _107_ 0.01249f
C12887 _132_ FILLER_0_17_104/a_572_375# 0.003857f
C12888 _427_/a_1308_423# net74 0.005627f
C12889 FILLER_0_2_93/a_484_472# net14 0.019214f
C12890 _077_ _078_ 0.069858f
C12891 net55 FILLER_0_17_38/a_124_375# 0.003236f
C12892 net72 FILLER_0_17_38/a_484_472# 0.00547f
C12893 _323_/a_36_113# _060_ 0.002584f
C12894 FILLER_0_13_228/a_36_472# net79 0.006824f
C12895 _141_ _143_ 0.192528f
C12896 net36 _196_/a_36_160# 0.024527f
C12897 _131_ FILLER_0_10_107/a_572_375# 0.007252f
C12898 net56 net36 0.772486f
C12899 _132_ _148_ 0.002873f
C12900 net27 output27/a_224_472# 0.046353f
C12901 FILLER_0_17_142/a_484_472# vss 0.030872f
C12902 net17 FILLER_0_12_28/a_124_375# 0.009108f
C12903 ctln[0] vdd 0.051631f
C12904 output12/a_224_472# vss 0.013728f
C12905 _155_ _153_ 0.033366f
C12906 _057_ _085_ 0.543871f
C12907 _225_/a_36_160# vdd 0.058272f
C12908 FILLER_0_14_107/a_572_375# _451_/a_36_151# 0.02627f
C12909 FILLER_0_6_47/a_1468_375# vdd -0.014642f
C12910 _093_ FILLER_0_18_177/a_3260_375# 0.002695f
C12911 cal_count\[3\] state\[1\] 0.236393f
C12912 _427_/a_2560_156# _095_ 0.009888f
C12913 FILLER_0_2_93/a_36_472# trim_mask\[3\] 0.003417f
C12914 output8/a_224_472# vdd 0.023187f
C12915 _068_ FILLER_0_5_148/a_124_375# 0.003986f
C12916 FILLER_0_21_142/a_36_472# FILLER_0_22_128/a_1468_375# 0.001543f
C12917 FILLER_0_4_177/a_484_472# net22 0.006506f
C12918 net18 _193_/a_36_160# 0.114176f
C12919 mask\[9\] FILLER_0_19_111/a_36_472# 0.285112f
C12920 net61 mask\[7\] 0.071542f
C12921 _066_ _163_ 0.006401f
C12922 FILLER_0_12_124/a_124_375# _131_ 0.07304f
C12923 FILLER_0_17_38/a_572_375# _182_ 0.035561f
C12924 vdd FILLER_0_12_196/a_36_472# 0.019648f
C12925 vss FILLER_0_12_196/a_124_375# 0.042104f
C12926 output8/a_224_472# net20 0.084627f
C12927 fanout53/a_36_160# net53 0.014917f
C12928 _428_/a_2665_112# net53 0.002379f
C12929 trim_val\[2\] _164_ 0.005847f
C12930 cal_count\[1\] _180_ 0.300952f
C12931 _050_ _436_/a_796_472# 0.007055f
C12932 FILLER_0_19_195/a_124_375# FILLER_0_19_187/a_572_375# 0.012001f
C12933 _035_ net17 0.021052f
C12934 _081_ cal_itt\[0\] 0.036569f
C12935 net80 vss 0.347557f
C12936 FILLER_0_1_266/a_572_375# rstn 0.00328f
C12937 _444_/a_1204_472# net47 0.007847f
C12938 _414_/a_1308_423# _074_ 0.005458f
C12939 vss FILLER_0_6_231/a_124_375# 0.00353f
C12940 vdd FILLER_0_6_231/a_572_375# 0.018694f
C12941 net50 vdd 0.661261f
C12942 FILLER_0_15_10/a_36_472# FILLER_0_15_2/a_484_472# 0.013277f
C12943 FILLER_0_9_223/a_484_472# net4 0.047334f
C12944 net38 _245_/a_672_472# 0.006341f
C12945 _141_ _146_ 0.020044f
C12946 _068_ _313_/a_255_603# 0.001149f
C12947 net67 _450_/a_448_472# 0.068692f
C12948 _136_ _070_ 0.010577f
C12949 _019_ _138_ 0.003734f
C12950 net57 _443_/a_448_472# 0.001956f
C12951 _053_ _058_ 0.075418f
C12952 FILLER_0_18_107/a_2724_472# vdd 0.004677f
C12953 net23 _163_ 0.034799f
C12954 _084_ _082_ 0.044645f
C12955 _382_/a_224_472# vdd 0.001663f
C12956 result[7] FILLER_0_24_290/a_36_472# 0.005185f
C12957 _429_/a_2665_112# _098_ 0.003225f
C12958 _136_ FILLER_0_15_180/a_124_375# 0.002442f
C12959 net82 _084_ 0.020793f
C12960 FILLER_0_7_195/a_124_375# cal_itt\[3\] 0.034632f
C12961 _394_/a_728_93# _175_ 0.010801f
C12962 _424_/a_1204_472# vdd 0.001573f
C12963 FILLER_0_15_150/a_124_375# _427_/a_448_472# 0.008952f
C12964 FILLER_0_1_192/a_124_375# vdd 0.017212f
C12965 net41 _444_/a_1000_472# 0.002179f
C12966 net20 FILLER_0_6_231/a_572_375# 0.01215f
C12967 net34 vss 0.481379f
C12968 en net18 0.32189f
C12969 net65 cal_itt\[0\] 0.07564f
C12970 _008_ net64 0.001427f
C12971 net50 _441_/a_1204_472# 0.006986f
C12972 net52 _441_/a_2665_112# 0.004975f
C12973 FILLER_0_4_107/a_484_472# _153_ 0.026082f
C12974 FILLER_0_4_107/a_1380_472# _154_ 0.005297f
C12975 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_572_375# 0.086635f
C12976 cal_itt\[3\] net22 0.134309f
C12977 net60 vss 0.382678f
C12978 net54 FILLER_0_19_111/a_484_472# 0.00105f
C12979 output36/a_224_472# _417_/a_2665_112# 0.008243f
C12980 net29 _195_/a_67_603# 0.048817f
C12981 FILLER_0_21_133/a_124_375# net54 0.013027f
C12982 net18 _417_/a_2248_156# 0.001601f
C12983 FILLER_0_16_57/a_1020_375# net15 0.048731f
C12984 FILLER_0_7_72/a_3172_472# vdd 0.003913f
C12985 _417_/a_2665_112# net30 0.015638f
C12986 net33 FILLER_0_22_128/a_3260_375# 0.001178f
C12987 FILLER_0_12_136/a_1468_375# vss 0.043987f
C12988 _064_ net47 0.110169f
C12989 _441_/a_2665_112# net49 0.062459f
C12990 _274_/a_36_68# net20 0.021022f
C12991 output35/a_224_472# _435_/a_2248_156# 0.019736f
C12992 FILLER_0_21_206/a_36_472# _204_/a_67_603# 0.003123f
C12993 FILLER_0_5_172/a_36_472# _163_ 0.006934f
C12994 FILLER_0_8_239/a_36_472# vss 0.003115f
C12995 FILLER_0_19_134/a_124_375# _145_ 0.023167f
C12996 input1/a_36_113# net18 0.004922f
C12997 _074_ FILLER_0_6_177/a_572_375# 0.012642f
C12998 _428_/a_448_472# FILLER_0_14_107/a_932_472# 0.007f
C12999 FILLER_0_5_72/a_572_375# vdd -0.00211f
C13000 FILLER_0_5_72/a_124_375# vss 0.041166f
C13001 net41 FILLER_0_21_28/a_124_375# 0.003254f
C13002 _065_ net15 0.065255f
C13003 net69 FILLER_0_2_111/a_36_472# 0.010759f
C13004 _031_ FILLER_0_2_111/a_1020_375# 0.016661f
C13005 net61 _422_/a_2248_156# 0.027973f
C13006 FILLER_0_18_177/a_1828_472# FILLER_0_19_187/a_572_375# 0.001684f
C13007 net14 FILLER_0_4_91/a_572_375# 0.047331f
C13008 _420_/a_36_151# net77 0.023469f
C13009 _098_ FILLER_0_19_171/a_124_375# 0.040575f
C13010 _431_/a_2665_112# vss 0.033886f
C13011 _122_ FILLER_0_8_156/a_124_375# 0.032617f
C13012 _441_/a_36_151# _440_/a_36_151# 0.003983f
C13013 net38 net6 0.071232f
C13014 output45/a_224_472# trimb[2] 0.045907f
C13015 _267_/a_672_472# _071_ 0.00255f
C13016 net67 _043_ 0.003726f
C13017 FILLER_0_9_28/a_2276_472# vss -0.001894f
C13018 net42 net47 0.237866f
C13019 _093_ _111_ 0.555171f
C13020 _446_/a_448_472# net40 0.05302f
C13021 _426_/a_36_151# FILLER_0_8_247/a_124_375# 0.059049f
C13022 _012_ FILLER_0_23_44/a_932_472# 0.001572f
C13023 net34 _107_ 0.017589f
C13024 _227_/a_36_160# FILLER_0_8_156/a_124_375# 0.005398f
C13025 FILLER_0_4_177/a_484_472# vdd 0.010663f
C13026 FILLER_0_4_177/a_36_472# vss 0.001806f
C13027 _375_/a_960_497# vdd 0.004471f
C13028 _057_ _062_ 0.062063f
C13029 _081_ FILLER_0_5_148/a_572_375# 0.01425f
C13030 _421_/a_448_472# net19 0.058446f
C13031 _008_ _418_/a_1308_423# 0.027229f
C13032 net15 FILLER_0_15_59/a_36_472# 0.00464f
C13033 net36 FILLER_0_15_180/a_36_472# 0.007275f
C13034 _008_ _006_ 0.02963f
C13035 _020_ _431_/a_448_472# 0.05255f
C13036 _114_ _311_/a_1920_473# 0.005579f
C13037 _445_/a_2665_112# trim_mask\[1\] 0.00183f
C13038 _384_/a_224_472# _160_ 0.00324f
C13039 net27 _415_/a_1308_423# 0.02437f
C13040 FILLER_0_22_177/a_484_472# _435_/a_36_151# 0.001723f
C13041 net51 _450_/a_2449_156# 0.008215f
C13042 _276_/a_36_160# vss 0.02914f
C13043 _035_ _446_/a_1308_423# 0.002639f
C13044 net68 net67 0.147318f
C13045 _008_ _103_ 0.092504f
C13046 _292_/a_36_160# output18/a_224_472# 0.009736f
C13047 _021_ net57 0.00736f
C13048 FILLER_0_13_65/a_124_375# _043_ 0.013045f
C13049 FILLER_0_15_72/a_484_472# vdd 0.002283f
C13050 FILLER_0_15_72/a_36_472# vss 0.038986f
C13051 mask\[4\] FILLER_0_19_155/a_124_375# 0.043876f
C13052 _015_ calibrate 0.105287f
C13053 _105_ net61 0.020753f
C13054 _427_/a_2665_112# state\[1\] 0.021573f
C13055 _419_/a_448_472# net77 0.007659f
C13056 _067_ net6 0.015232f
C13057 net81 FILLER_0_15_212/a_1468_375# 0.006906f
C13058 net47 FILLER_0_4_91/a_484_472# 0.007531f
C13059 _414_/a_1308_423# _081_ 0.003429f
C13060 FILLER_0_10_256/a_124_375# _015_ 0.001151f
C13061 FILLER_0_3_2/a_124_375# vss 0.007235f
C13062 FILLER_0_3_2/a_36_472# vdd 0.106665f
C13063 output27/a_224_472# net18 0.058296f
C13064 net27 FILLER_0_14_235/a_484_472# 0.010072f
C13065 net75 _083_ 0.055491f
C13066 net50 fanout67/a_36_160# 0.007195f
C13067 _096_ _116_ 0.020685f
C13068 FILLER_0_1_98/a_124_375# _065_ 0.001136f
C13069 ctln[8] trim_val\[3\] 0.007f
C13070 _067_ _172_ 0.010195f
C13071 net55 FILLER_0_17_56/a_572_375# 0.020564f
C13072 cal_itt\[3\] vdd 0.571239f
C13073 _070_ FILLER_0_10_107/a_484_472# 0.007421f
C13074 FILLER_0_23_88/a_124_375# net14 0.002894f
C13075 FILLER_0_16_107/a_124_375# _093_ 0.003941f
C13076 _431_/a_1000_472# _020_ 0.009685f
C13077 _093_ FILLER_0_17_72/a_1916_375# 0.017467f
C13078 output28/a_224_472# net28 0.048681f
C13079 FILLER_0_9_223/a_572_375# vss 0.00704f
C13080 _056_ _311_/a_254_473# 0.005937f
C13081 _428_/a_1000_472# vdd 0.005345f
C13082 _098_ _433_/a_1000_472# 0.0184f
C13083 FILLER_0_3_204/a_124_375# net59 0.007104f
C13084 ctlp[7] net25 0.003141f
C13085 _009_ vdd 0.693198f
C13086 FILLER_0_16_255/a_36_472# net19 0.001273f
C13087 net4 _070_ 0.169392f
C13088 _437_/a_1308_423# net14 0.085815f
C13089 _068_ FILLER_0_9_142/a_124_375# 0.008226f
C13090 _076_ FILLER_0_9_142/a_36_472# 0.038562f
C13091 trim_mask\[4\] _369_/a_36_68# 0.00407f
C13092 _394_/a_1336_472# vdd 0.003226f
C13093 _106_ mask\[3\] 0.249479f
C13094 FILLER_0_11_142/a_36_472# net23 0.002015f
C13095 _081_ FILLER_0_6_177/a_572_375# 0.007285f
C13096 _412_/a_36_151# _082_ 0.016538f
C13097 _059_ _160_ 0.037235f
C13098 _422_/a_796_472# _009_ 0.001178f
C13099 net20 _009_ 0.026064f
C13100 output42/a_224_472# FILLER_0_8_24/a_124_375# 0.001168f
C13101 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_572_375# 0.086635f
C13102 _412_/a_36_151# net82 0.064296f
C13103 vdd _039_ 0.219985f
C13104 FILLER_0_18_107/a_932_472# FILLER_0_16_115/a_124_375# 0.001512f
C13105 fanout68/a_36_113# _441_/a_36_151# 0.138322f
C13106 _274_/a_1612_497# state\[0\] 0.001071f
C13107 _112_ _316_/a_1084_68# 0.005773f
C13108 _189_/a_67_603# FILLER_0_13_228/a_124_375# 0.00744f
C13109 FILLER_0_21_142/a_572_375# net54 0.043619f
C13110 output9/a_224_472# vdd 0.102412f
C13111 _128_ _076_ 0.04562f
C13112 net15 _449_/a_2248_156# 0.001705f
C13113 _016_ _427_/a_36_151# 0.00483f
C13114 _086_ FILLER_0_6_177/a_572_375# 0.012909f
C13115 FILLER_0_9_28/a_1828_472# net16 0.001946f
C13116 FILLER_0_20_177/a_1020_375# _098_ 0.013949f
C13117 _091_ _432_/a_1308_423# 0.008903f
C13118 FILLER_0_15_212/a_1380_472# mask\[1\] 0.041503f
C13119 net55 _452_/a_1353_112# 0.030679f
C13120 FILLER_0_5_164/a_124_375# _386_/a_848_380# 0.014613f
C13121 _068_ _311_/a_254_473# 0.002606f
C13122 state\[0\] net64 0.01679f
C13123 net25 FILLER_0_23_88/a_36_472# 0.192699f
C13124 result[7] FILLER_0_23_282/a_484_472# 0.013947f
C13125 FILLER_0_17_200/a_484_472# _430_/a_36_151# 0.001723f
C13126 net76 FILLER_0_1_192/a_36_472# 0.003817f
C13127 _334_/a_36_160# FILLER_0_17_104/a_1468_375# 0.027706f
C13128 net54 _436_/a_1000_472# 0.002051f
C13129 _427_/a_36_151# FILLER_0_14_123/a_124_375# 0.023595f
C13130 net57 _163_ 0.759175f
C13131 _173_ _042_ 0.002294f
C13132 _424_/a_2665_112# _423_/a_2248_156# 0.001314f
C13133 trim_mask\[1\] FILLER_0_6_47/a_932_472# 0.007542f
C13134 FILLER_0_7_72/a_1380_472# net50 0.077411f
C13135 _434_/a_2560_156# vdd 0.002922f
C13136 _434_/a_2665_112# vss 0.00127f
C13137 _067_ _450_/a_2225_156# 0.002584f
C13138 cal_itt\[3\] _251_/a_1130_472# 0.001099f
C13139 FILLER_0_15_116/a_572_375# _136_ 0.001706f
C13140 _000_ ctln[4] 0.002823f
C13141 net82 _316_/a_848_380# 0.087022f
C13142 _091_ FILLER_0_19_171/a_1468_375# 0.002731f
C13143 fanout61/a_36_113# _418_/a_36_151# 0.001442f
C13144 _322_/a_848_380# vdd 0.067623f
C13145 _322_/a_124_24# vss 0.003731f
C13146 net18 _416_/a_36_151# 0.027435f
C13147 FILLER_0_4_99/a_36_472# _030_ 0.002699f
C13148 _273_/a_36_68# _055_ 0.081216f
C13149 _231_/a_652_68# _062_ 0.001555f
C13150 _098_ _047_ 0.062495f
C13151 net75 _425_/a_36_151# 0.02868f
C13152 FILLER_0_12_136/a_1468_375# _071_ 0.002023f
C13153 FILLER_0_2_101/a_124_375# vss 0.04897f
C13154 FILLER_0_2_101/a_36_472# vdd 0.099518f
C13155 FILLER_0_4_144/a_124_375# vss 0.017638f
C13156 FILLER_0_4_144/a_572_375# vdd -0.013698f
C13157 output31/a_224_472# net60 0.216716f
C13158 vss FILLER_0_8_156/a_484_472# 0.004078f
C13159 _412_/a_2665_112# vss 0.011887f
C13160 _188_ FILLER_0_12_50/a_36_472# 0.006464f
C13161 net35 FILLER_0_22_128/a_3260_375# 0.012732f
C13162 net17 _452_/a_1353_112# 0.038603f
C13163 _205_/a_36_160# _047_ 0.013528f
C13164 _207_/a_67_603# _146_ 0.026192f
C13165 net55 _453_/a_2248_156# 0.001546f
C13166 net35 net33 1.594925f
C13167 _250_/a_36_68# state\[2\] 0.038165f
C13168 output10/a_224_472# vss 0.014205f
C13169 net58 _084_ 0.141836f
C13170 net68 FILLER_0_6_47/a_1916_375# 0.00799f
C13171 _265_/a_244_68# vdd 0.022571f
C13172 net15 _439_/a_1000_472# 0.001798f
C13173 FILLER_0_18_100/a_124_375# _438_/a_2665_112# 0.010688f
C13174 _086_ FILLER_0_10_107/a_572_375# 0.001179f
C13175 _431_/a_36_151# FILLER_0_15_116/a_572_375# 0.001543f
C13176 FILLER_0_16_107/a_124_375# _136_ 0.00661f
C13177 _415_/a_1308_423# net18 0.010051f
C13178 net60 _419_/a_1000_472# 0.028992f
C13179 net61 _419_/a_2248_156# 0.022159f
C13180 _020_ _132_ 0.037636f
C13181 FILLER_0_17_104/a_484_472# vdd 0.020339f
C13182 FILLER_0_17_104/a_36_472# vss 0.002744f
C13183 _444_/a_448_472# net40 0.055844f
C13184 net54 FILLER_0_22_128/a_124_375# 0.032013f
C13185 _091_ net22 0.031921f
C13186 FILLER_0_17_72/a_1916_375# _136_ 0.009573f
C13187 FILLER_0_8_24/a_124_375# net40 0.002431f
C13188 _450_/a_1697_156# net6 0.00236f
C13189 _153_ FILLER_0_4_91/a_572_375# 0.001735f
C13190 _093_ fanout54/a_36_160# 0.003506f
C13191 net4 _082_ 0.004529f
C13192 mask\[4\] FILLER_0_19_187/a_572_375# 0.00553f
C13193 _230_/a_244_68# _056_ 0.001844f
C13194 net82 net4 1.982825f
C13195 FILLER_0_9_223/a_124_375# _055_ 0.014525f
C13196 _274_/a_36_68# _069_ 0.02257f
C13197 _300_/a_224_472# _011_ 0.007508f
C13198 net55 FILLER_0_18_53/a_572_375# 0.015895f
C13199 fanout50/a_36_160# trim_val\[3\] 0.017252f
C13200 result[7] output34/a_224_472# 0.057094f
C13201 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1468_375# 0.001597f
C13202 net16 FILLER_0_8_37/a_484_472# 0.004272f
C13203 result[8] net61 0.001106f
C13204 _267_/a_224_472# state\[1\] 0.001937f
C13205 _008_ mask\[2\] 0.003475f
C13206 net65 en 0.001469f
C13207 FILLER_0_23_290/a_124_375# vss 0.033011f
C13208 FILLER_0_23_290/a_36_472# vdd 0.089567f
C13209 FILLER_0_15_116/a_484_472# net36 0.009319f
C13210 net39 _445_/a_2560_156# 0.003401f
C13211 _093_ net21 0.032584f
C13212 FILLER_0_16_89/a_572_375# _131_ 0.012481f
C13213 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_124_375# 0.026339f
C13214 FILLER_0_12_136/a_1020_375# _126_ 0.012732f
C13215 FILLER_0_4_197/a_932_472# net59 0.003599f
C13216 net80 FILLER_0_22_177/a_572_375# 0.005202f
C13217 output34/a_224_472# _198_/a_67_603# 0.00179f
C13218 net10 vdd 0.227004f
C13219 _086_ _128_ 0.085571f
C13220 _141_ mask\[2\] 0.084094f
C13221 FILLER_0_10_78/a_484_472# cal_count\[3\] 0.001112f
C13222 _050_ FILLER_0_22_107/a_572_375# 0.001825f
C13223 FILLER_0_20_193/a_572_375# vss 0.005887f
C13224 FILLER_0_20_193/a_36_472# vdd 0.091886f
C13225 _293_/a_36_472# vss 0.014842f
C13226 net73 fanout71/a_36_113# 0.004833f
C13227 FILLER_0_17_72/a_1380_472# _131_ 0.006873f
C13228 FILLER_0_4_177/a_484_472# FILLER_0_2_177/a_572_375# 0.001512f
C13229 _420_/a_1308_423# _009_ 0.014359f
C13230 net10 net20 0.02842f
C13231 _369_/a_36_68# _154_ 0.042308f
C13232 net34 FILLER_0_22_177/a_572_375# 0.006974f
C13233 _413_/a_36_151# FILLER_0_3_172/a_2364_375# 0.059049f
C13234 _070_ _058_ 0.07307f
C13235 net72 vdd 1.425686f
C13236 FILLER_0_15_116/a_572_375# net53 0.012526f
C13237 _085_ _161_ 0.008926f
C13238 _438_/a_448_472# net71 0.044454f
C13239 _421_/a_2665_112# _109_ 0.002029f
C13240 output8/a_224_472# cal_itt\[2\] 0.05561f
C13241 FILLER_0_5_109/a_572_375# FILLER_0_4_107/a_932_472# 0.001684f
C13242 _118_ _313_/a_67_603# 0.001793f
C13243 _101_ _100_ 0.012073f
C13244 _035_ trim_mask\[2\] 0.004455f
C13245 FILLER_0_5_54/a_36_472# vss 0.001756f
C13246 FILLER_0_5_54/a_484_472# vdd 0.003166f
C13247 net33 net22 0.066751f
C13248 net16 _131_ 0.001308f
C13249 output42/a_224_472# net44 0.079084f
C13250 _144_ _434_/a_36_151# 0.004055f
C13251 _176_ _131_ 1.798819f
C13252 FILLER_0_7_104/a_1468_375# _154_ 0.003683f
C13253 _431_/a_2560_156# FILLER_0_17_142/a_124_375# 0.001178f
C13254 _442_/a_2665_112# vdd 0.056153f
C13255 FILLER_0_21_125/a_36_472# _140_ 0.101284f
C13256 FILLER_0_10_37/a_124_375# net51 0.006198f
C13257 net34 _435_/a_2560_156# 0.002967f
C13258 _030_ _367_/a_692_472# 0.002082f
C13259 _149_ FILLER_0_20_87/a_124_375# 0.004191f
C13260 _079_ FILLER_0_5_212/a_124_375# 0.005363f
C13261 net15 FILLER_0_6_47/a_1380_472# 0.00464f
C13262 FILLER_0_16_241/a_36_472# vss 0.004432f
C13263 FILLER_0_18_177/a_1916_375# vdd 0.021f
C13264 net47 _450_/a_2449_156# 0.004488f
C13265 _449_/a_1204_472# _067_ 0.014354f
C13266 _415_/a_36_151# FILLER_0_10_256/a_124_375# 0.035117f
C13267 _112_ vss 0.145781f
C13268 FILLER_0_12_20/a_484_472# vss 0.001783f
C13269 _308_/a_1084_68# _115_ 0.001451f
C13270 _414_/a_2560_156# _074_ 0.001344f
C13271 _450_/a_1353_112# _039_ 0.019843f
C13272 FILLER_0_17_133/a_124_375# _137_ 0.009198f
C13273 _132_ _017_ 0.155924f
C13274 FILLER_0_18_2/a_2812_375# net40 0.018463f
C13275 net66 trim[3] 0.00567f
C13276 _091_ vdd 1.011371f
C13277 net16 FILLER_0_18_37/a_572_375# 0.03477f
C13278 FILLER_0_15_282/a_124_375# _006_ 0.002249f
C13279 _398_/a_36_113# net17 0.002702f
C13280 FILLER_0_17_72/a_1916_375# net53 0.001657f
C13281 FILLER_0_16_57/a_36_472# _183_ 0.004107f
C13282 _068_ _261_/a_36_160# 0.008557f
C13283 _133_ _059_ 0.039848f
C13284 net41 _450_/a_2225_156# 0.024042f
C13285 _104_ _421_/a_1308_423# 0.001621f
C13286 net17 FILLER_0_20_15/a_1020_375# 0.039975f
C13287 _370_/a_848_380# vss 0.051599f
C13288 _410_/a_36_68# net51 0.014342f
C13289 _131_ _124_ 0.002448f
C13290 mask\[7\] FILLER_0_22_128/a_1916_375# 0.007718f
C13291 trim_val\[3\] net14 0.01035f
C13292 _163_ FILLER_0_5_148/a_572_375# 0.001706f
C13293 FILLER_0_17_72/a_1020_375# _175_ 0.028592f
C13294 FILLER_0_18_177/a_3260_375# _047_ 0.030543f
C13295 cal_count\[2\] FILLER_0_15_10/a_124_375# 0.017594f
C13296 _070_ _389_/a_36_148# 0.010534f
C13297 _091_ net20 0.0557f
C13298 FILLER_0_7_162/a_36_472# net57 0.015199f
C13299 output33/a_224_472# net19 0.12997f
C13300 _093_ FILLER_0_18_61/a_124_375# 0.031062f
C13301 output27/a_224_472# net65 0.019729f
C13302 net38 FILLER_0_12_2/a_572_375# 0.00609f
C13303 FILLER_0_14_50/a_36_472# cal_count\[3\] 0.005814f
C13304 _431_/a_3041_156# vss 0.001312f
C13305 FILLER_0_21_28/a_3172_472# _424_/a_36_151# 0.001723f
C13306 trim_val\[3\] _164_ 0.018411f
C13307 net61 output18/a_224_472# 0.059062f
C13308 _002_ _413_/a_1000_472# 0.006249f
C13309 net52 _439_/a_36_151# 0.01388f
C13310 _115_ FILLER_0_9_72/a_1380_472# 0.007262f
C13311 FILLER_0_9_223/a_36_472# _076_ 0.00146f
C13312 _091_ _430_/a_2248_156# 0.053571f
C13313 _335_/a_49_472# mask\[1\] 0.032497f
C13314 FILLER_0_16_57/a_484_472# FILLER_0_15_59/a_124_375# 0.001543f
C13315 _394_/a_728_93# _043_ 0.00355f
C13316 _119_ _322_/a_124_24# 0.020461f
C13317 _136_ net21 0.022198f
C13318 _024_ vss 0.132549f
C13319 net58 _412_/a_36_151# 0.010226f
C13320 FILLER_0_12_124/a_36_472# _132_ 0.00101f
C13321 _128_ _090_ 0.018296f
C13322 _136_ _333_/a_36_160# 0.00842f
C13323 cal_count\[1\] vss 0.307993f
C13324 _428_/a_796_472# _095_ 0.00117f
C13325 _002_ FILLER_0_3_172/a_3172_472# 0.002313f
C13326 _341_/a_665_69# _141_ 0.001064f
C13327 _178_ cal_count\[1\] 0.470244f
C13328 _443_/a_2248_156# _170_ 0.068179f
C13329 _061_ _060_ 0.066418f
C13330 state\[2\] FILLER_0_13_142/a_36_472# 0.022678f
C13331 net53 FILLER_0_13_142/a_932_472# 0.059367f
C13332 net15 _440_/a_796_472# 0.005848f
C13333 _119_ FILLER_0_8_156/a_484_472# 0.00979f
C13334 _015_ FILLER_0_8_247/a_124_375# 0.00706f
C13335 FILLER_0_3_78/a_124_375# vdd 0.002419f
C13336 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_572_375# 0.086635f
C13337 _448_/a_2665_112# _037_ 0.042225f
C13338 _367_/a_36_68# net14 0.055776f
C13339 net44 net40 0.003336f
C13340 _161_ _062_ 0.046903f
C13341 vdd trim[2] 0.166648f
C13342 FILLER_0_22_128/a_2812_375# vss 0.004347f
C13343 FILLER_0_22_128/a_3260_375# vdd 0.005207f
C13344 output22/a_224_472# _435_/a_1308_423# 0.005111f
C13345 net71 FILLER_0_22_107/a_484_472# 0.00689f
C13346 FILLER_0_8_107/a_124_375# FILLER_0_10_107/a_36_472# 0.0027f
C13347 _100_ _094_ 0.031066f
C13348 result[6] ctlp[2] 0.001324f
C13349 net33 vdd 0.42212f
C13350 net27 _426_/a_36_151# 0.008613f
C13351 output15/a_224_472# FILLER_0_0_96/a_124_375# 0.00515f
C13352 _413_/a_36_151# net76 0.084453f
C13353 FILLER_0_3_78/a_36_472# _168_ 0.063262f
C13354 FILLER_0_20_15/a_1380_472# net40 0.014911f
C13355 _431_/a_796_472# net73 0.002306f
C13356 _414_/a_36_151# FILLER_0_6_177/a_572_375# 0.073306f
C13357 trimb[0] vdd 0.10929f
C13358 FILLER_0_6_79/a_36_472# vss 0.008693f
C13359 _129_ _062_ 0.20212f
C13360 _079_ FILLER_0_3_172/a_1828_472# 0.001638f
C13361 _053_ FILLER_0_6_47/a_1020_375# 0.015621f
C13362 _425_/a_36_151# net19 0.009499f
C13363 net76 _078_ 0.029213f
C13364 _406_/a_36_159# _402_/a_56_567# 0.001025f
C13365 net82 FILLER_0_3_172/a_1468_375# 0.010439f
C13366 FILLER_0_21_206/a_124_375# _048_ 0.018458f
C13367 FILLER_0_13_228/a_124_375# _043_ 0.133079f
C13368 FILLER_0_5_109/a_572_375# _163_ 0.003096f
C13369 FILLER_0_15_282/a_484_472# vss 0.005507f
C13370 trim_val\[0\] _164_ 0.133785f
C13371 net80 _147_ 0.022618f
C13372 FILLER_0_17_38/a_484_472# vdd 0.009211f
C13373 _072_ _060_ 0.080908f
C13374 FILLER_0_3_172/a_572_375# net65 0.008318f
C13375 FILLER_0_3_2/a_124_375# output41/a_224_472# 0.030009f
C13376 net79 _418_/a_36_151# 0.059124f
C13377 _392_/a_36_68# vss 0.002019f
C13378 vdd FILLER_0_3_212/a_36_472# 0.110132f
C13379 vss FILLER_0_3_212/a_124_375# 0.009048f
C13380 FILLER_0_6_177/a_572_375# _163_ 0.001839f
C13381 _116_ _061_ 0.04837f
C13382 _292_/a_36_160# _048_ 0.008475f
C13383 net63 _137_ 0.006317f
C13384 FILLER_0_17_282/a_124_375# vdd 0.004586f
C13385 _152_ _261_/a_36_160# 0.001102f
C13386 _316_/a_848_380# calibrate 0.012121f
C13387 _316_/a_124_24# _122_ 0.040082f
C13388 _414_/a_2560_156# _081_ 0.008322f
C13389 _116_ _311_/a_66_473# 0.001527f
C13390 _149_ _098_ 0.398643f
C13391 _131_ _041_ 0.035642f
C13392 _115_ FILLER_0_9_105/a_36_472# 0.004013f
C13393 _306_/a_36_68# vdd 0.044152f
C13394 net62 FILLER_0_21_286/a_572_375# 0.003744f
C13395 net34 _147_ 0.144404f
C13396 _449_/a_36_151# _394_/a_1336_472# 0.001582f
C13397 FILLER_0_10_107/a_36_472# FILLER_0_10_94/a_484_472# 0.001963f
C13398 _412_/a_448_472# net81 0.047334f
C13399 net52 FILLER_0_6_47/a_3260_375# 0.040612f
C13400 FILLER_0_10_78/a_1380_472# vss 0.002096f
C13401 _115_ vdd 0.455713f
C13402 _028_ FILLER_0_5_72/a_1020_375# 0.00123f
C13403 FILLER_0_23_60/a_124_375# vdd 0.031398f
C13404 mask\[9\] FILLER_0_20_98/a_124_375# 0.003444f
C13405 net55 FILLER_0_19_28/a_572_375# 0.002115f
C13406 _077_ FILLER_0_9_105/a_484_472# 0.002951f
C13407 _440_/a_2665_112# FILLER_0_4_91/a_124_375# 0.006271f
C13408 FILLER_0_12_2/a_36_472# clkc 0.004826f
C13409 FILLER_0_18_100/a_124_375# vdd 0.044014f
C13410 _431_/a_1204_472# _137_ 0.005886f
C13411 _096_ FILLER_0_14_181/a_36_472# 0.028078f
C13412 _066_ net37 0.006164f
C13413 _379_/a_36_472# _166_ 0.038062f
C13414 _443_/a_1204_472# net69 0.002642f
C13415 net58 net4 0.858616f
C13416 _061_ _118_ 0.268815f
C13417 _077_ vss 1.071923f
C13418 _426_/a_2665_112# FILLER_0_8_239/a_124_375# 0.010736f
C13419 net54 FILLER_0_22_107/a_36_472# 0.043792f
C13420 _143_ _432_/a_36_151# 0.001486f
C13421 net72 _403_/a_224_472# 0.002276f
C13422 _433_/a_1308_423# _145_ 0.026613f
C13423 net74 _372_/a_170_472# 0.079123f
C13424 _176_ _076_ 0.046873f
C13425 _118_ _311_/a_66_473# 0.008528f
C13426 _072_ _116_ 0.283323f
C13427 _328_/a_36_113# vss 0.044028f
C13428 _236_/a_36_160# net39 0.052649f
C13429 net35 net22 0.001381f
C13430 net23 FILLER_0_19_155/a_124_375# 0.001347f
C13431 FILLER_0_17_72/a_124_375# vss 0.048053f
C13432 FILLER_0_17_72/a_572_375# vdd 0.002455f
C13433 output19/a_224_472# vss 0.048948f
C13434 net41 trim[3] 0.005906f
C13435 cal_count\[3\] _121_ 0.011368f
C13436 FILLER_0_17_161/a_124_375# _137_ 0.016092f
C13437 net23 net37 0.01763f
C13438 _106_ _294_/a_224_472# 0.001038f
C13439 net73 FILLER_0_18_107/a_1380_472# 0.039646f
C13440 net4 calibrate 0.04302f
C13441 _412_/a_36_151# fanout81/a_36_160# 0.001725f
C13442 _430_/a_796_472# net21 0.015066f
C13443 FILLER_0_4_107/a_124_375# vss 0.00322f
C13444 FILLER_0_4_107/a_572_375# vdd 0.034678f
C13445 FILLER_0_9_270/a_124_375# vdd 0.013312f
C13446 net41 _402_/a_718_527# 0.019628f
C13447 _445_/a_2560_156# net47 0.014069f
C13448 net38 FILLER_0_20_2/a_572_375# 0.004413f
C13449 FILLER_0_21_125/a_572_375# _098_ 0.006462f
C13450 _053_ FILLER_0_9_28/a_2276_472# 0.002243f
C13451 ctlp[2] _422_/a_36_151# 0.068086f
C13452 _395_/a_36_488# vdd 0.066813f
C13453 fanout63/a_36_160# net64 0.016132f
C13454 net54 FILLER_0_20_98/a_36_472# 0.059367f
C13455 net57 FILLER_0_16_154/a_932_472# 0.003453f
C13456 cal_count\[2\] _180_ 0.153207f
C13457 FILLER_0_9_28/a_932_472# FILLER_0_10_37/a_36_472# 0.026657f
C13458 _120_ vss 0.42505f
C13459 _072_ _118_ 0.120452f
C13460 _038_ vss 0.373776f
C13461 net60 _421_/a_1308_423# 0.020693f
C13462 _136_ mask\[1\] 0.407932f
C13463 net48 cal_itt\[0\] 0.006171f
C13464 _257_/a_36_472# _074_ 0.011352f
C13465 _449_/a_2248_156# net74 0.004565f
C13466 en_co_clk _176_ 0.099475f
C13467 _401_/a_36_68# cal_count\[1\] 0.006747f
C13468 FILLER_0_4_197/a_572_375# net76 0.006026f
C13469 net41 _445_/a_2665_112# 0.056125f
C13470 _144_ _354_/a_665_69# 0.001518f
C13471 result[8] FILLER_0_23_274/a_36_472# 0.001908f
C13472 _009_ net77 0.001183f
C13473 FILLER_0_23_282/a_572_375# vdd -0.013698f
C13474 FILLER_0_23_282/a_124_375# vss 0.005048f
C13475 FILLER_0_17_200/a_484_472# net63 0.003767f
C13476 net81 _429_/a_796_472# 0.002847f
C13477 net62 mask\[1\] 0.227329f
C13478 net76 _263_/a_224_472# 0.00132f
C13479 _438_/a_2665_112# vdd 0.00587f
C13480 _438_/a_2248_156# vss 0.002607f
C13481 _030_ _440_/a_36_151# 0.001187f
C13482 fanout66/a_36_113# net15 0.024302f
C13483 FILLER_0_5_172/a_36_472# net37 0.013857f
C13484 FILLER_0_13_142/a_1468_375# vdd 0.028002f
C13485 ctlp[6] vdd 0.207209f
C13486 FILLER_0_13_142/a_1020_375# vss 0.005307f
C13487 _098_ FILLER_0_18_209/a_572_375# 0.001352f
C13488 _020_ FILLER_0_18_107/a_2364_375# 0.003755f
C13489 net52 FILLER_0_5_72/a_484_472# 0.050714f
C13490 net50 FILLER_0_5_72/a_1468_375# 0.001777f
C13491 _053_ _359_/a_1492_488# 0.001437f
C13492 _131_ FILLER_0_17_64/a_124_375# 0.005913f
C13493 _056_ _062_ 0.320621f
C13494 FILLER_0_5_128/a_124_375# net47 0.011156f
C13495 _413_/a_2248_156# net82 0.009308f
C13496 _115_ _135_ 0.004345f
C13497 output19/a_224_472# _107_ 0.005034f
C13498 _087_ FILLER_0_5_172/a_124_375# 0.003043f
C13499 net15 FILLER_0_9_72/a_124_375# 0.006492f
C13500 _390_/a_36_68# _067_ 0.029588f
C13501 net19 FILLER_0_14_263/a_36_472# 0.135429f
C13502 output29/a_224_472# net18 0.010345f
C13503 net44 FILLER_0_15_2/a_484_472# 0.047161f
C13504 net52 _160_ 0.133292f
C13505 _081_ FILLER_0_5_136/a_36_472# 0.0028f
C13506 _152_ FILLER_0_5_136/a_124_375# 0.039558f
C13507 mask\[4\] _201_/a_255_603# 0.002111f
C13508 FILLER_0_19_55/a_124_375# vdd 0.035786f
C13509 FILLER_0_3_204/a_36_472# net65 0.001777f
C13510 comp FILLER_0_15_2/a_124_375# 0.034135f
C13511 _412_/a_2665_112# output37/a_224_472# 0.002025f
C13512 net17 _190_/a_36_160# 0.04702f
C13513 _164_ FILLER_0_6_47/a_484_472# 0.012286f
C13514 net54 _433_/a_36_151# 0.00661f
C13515 _412_/a_448_472# net2 0.033994f
C13516 _050_ _210_/a_67_603# 0.006444f
C13517 net68 FILLER_0_5_54/a_932_472# 0.013043f
C13518 fanout72/a_36_113# _174_ 0.026207f
C13519 FILLER_0_20_107/a_124_375# _098_ 0.01186f
C13520 FILLER_0_11_282/a_36_472# vdd 0.106843f
C13521 FILLER_0_11_282/a_124_375# vss 0.005415f
C13522 mask\[4\] FILLER_0_18_177/a_1380_472# 0.016924f
C13523 net15 _453_/a_1308_423# 0.00293f
C13524 _132_ cal_count\[3\] 0.193553f
C13525 _091_ _069_ 0.741596f
C13526 net49 _160_ 1.243817f
C13527 _413_/a_2560_156# vss 0.001097f
C13528 _447_/a_2560_156# net69 0.001774f
C13529 FILLER_0_14_81/a_124_375# _394_/a_728_93# 0.004587f
C13530 FILLER_0_9_223/a_36_472# _090_ 0.001057f
C13531 mask\[5\] _098_ 1.316993f
C13532 FILLER_0_7_72/a_572_375# _028_ 0.003837f
C13533 _068_ _062_ 0.089152f
C13534 _070_ _134_ 0.087767f
C13535 _256_/a_36_68# net4 0.017783f
C13536 net64 _005_ 0.006192f
C13537 result[5] _418_/a_36_151# 0.009705f
C13538 mask\[6\] vss 0.348967f
C13539 _417_/a_2665_112# _006_ 0.023025f
C13540 FILLER_0_7_104/a_1380_472# _131_ 0.043557f
C13541 mask\[8\] vss 0.378558f
C13542 net35 vdd 1.0365f
C13543 mask\[5\] _205_/a_36_160# 0.003775f
C13544 _086_ _176_ 0.837546f
C13545 _273_/a_36_68# _223_/a_36_160# 0.002786f
C13546 _320_/a_36_472# _113_ 0.030365f
C13547 net56 FILLER_0_17_142/a_572_375# 0.014948f
C13548 fanout81/a_36_160# net4 0.002848f
C13549 _014_ _123_ 0.050082f
C13550 FILLER_0_9_28/a_1468_375# FILLER_0_8_37/a_484_472# 0.001723f
C13551 _429_/a_2665_112# mask\[1\] 0.001022f
C13552 _367_/a_36_68# _153_ 0.019803f
C13553 FILLER_0_17_56/a_484_472# vss 0.006298f
C13554 result[6] FILLER_0_21_286/a_572_375# 0.015047f
C13555 _093_ _099_ 0.001725f
C13556 _411_/a_2248_156# net75 0.032114f
C13557 _025_ _436_/a_36_151# 0.026707f
C13558 mask\[3\] _019_ 0.001403f
C13559 _449_/a_36_151# net72 0.039436f
C13560 fanout52/a_36_160# vss 0.010082f
C13561 FILLER_0_5_128/a_124_375# net74 0.013683f
C13562 _432_/a_1308_423# vdd 0.029938f
C13563 net79 _416_/a_2665_112# 0.035115f
C13564 _430_/a_1000_472# mask\[2\] 0.00785f
C13565 net55 FILLER_0_18_76/a_36_472# 0.003695f
C13566 _114_ _225_/a_36_160# 0.003628f
C13567 net62 _416_/a_2560_156# 0.010748f
C13568 _431_/a_2665_112# FILLER_0_15_150/a_36_472# 0.035266f
C13569 _424_/a_448_472# FILLER_0_18_37/a_1020_375# 0.001674f
C13570 vss FILLER_0_13_290/a_36_472# 0.009561f
C13571 cal_count\[3\] _408_/a_728_93# 0.040643f
C13572 _093_ FILLER_0_19_111/a_124_375# 0.00186f
C13573 _128_ _117_ 0.045015f
C13574 FILLER_0_2_111/a_124_375# trim_mask\[3\] 0.004993f
C13575 state\[2\] vss 0.185787f
C13576 _453_/a_796_472# _042_ 0.005463f
C13577 _453_/a_1308_423# net51 0.001804f
C13578 _136_ _171_ 0.008792f
C13579 _095_ cal_count\[1\] 0.853949f
C13580 result[8] FILLER_0_24_274/a_1468_375# 0.00726f
C13581 _091_ net31 0.001465f
C13582 _440_/a_448_472# _164_ 0.0036f
C13583 _058_ FILLER_0_10_94/a_36_472# 0.009346f
C13584 _086_ _124_ 0.063099f
C13585 FILLER_0_20_177/a_572_375# FILLER_0_19_171/a_1380_472# 0.001543f
C13586 _102_ net30 0.043037f
C13587 _448_/a_36_151# net76 0.03831f
C13588 result[7] _419_/a_1204_472# 0.018181f
C13589 FILLER_0_7_72/a_932_472# net52 0.008749f
C13590 _175_ vss 0.162988f
C13591 _010_ _420_/a_448_472# 0.027802f
C13592 vdd _167_ 0.012869f
C13593 output23/a_224_472# _208_/a_36_160# 0.014541f
C13594 FILLER_0_19_171/a_1468_375# vdd 0.064097f
C13595 FILLER_0_22_86/a_932_472# net71 0.005789f
C13596 net15 FILLER_0_13_72/a_484_472# 0.002925f
C13597 _451_/a_836_156# net14 0.00174f
C13598 net81 _001_ 0.012492f
C13599 FILLER_0_5_72/a_1380_472# _164_ 0.049427f
C13600 _119_ _077_ 2.584241f
C13601 FILLER_0_4_152/a_124_375# FILLER_0_4_144/a_572_375# 0.012001f
C13602 net61 net18 0.71051f
C13603 _088_ FILLER_0_4_213/a_36_472# 0.01735f
C13604 net55 FILLER_0_21_28/a_3260_375# 0.006399f
C13605 net72 FILLER_0_21_28/a_932_472# 0.015756f
C13606 _058_ calibrate 0.075294f
C13607 net21 _047_ 0.048701f
C13608 mask\[0\] _136_ 0.025838f
C13609 _235_/a_67_603# vdd 0.026582f
C13610 FILLER_0_7_195/a_124_375# vdd 0.007788f
C13611 _242_/a_36_160# FILLER_0_5_148/a_484_472# 0.003699f
C13612 _136_ FILLER_0_13_100/a_36_472# 0.005029f
C13613 _363_/a_36_68# vss 0.043707f
C13614 _003_ vss 0.095366f
C13615 trim_mask\[4\] FILLER_0_2_111/a_1468_375# 0.001226f
C13616 FILLER_0_5_128/a_124_375# _159_ 0.003644f
C13617 net62 mask\[0\] 0.552008f
C13618 _359_/a_36_488# _131_ 0.006398f
C13619 FILLER_0_10_37/a_124_375# _173_ 0.00262f
C13620 _431_/a_448_472# fanout70/a_36_113# 0.001157f
C13621 FILLER_0_5_117/a_36_472# net47 0.005919f
C13622 FILLER_0_7_72/a_1020_375# _028_ 0.003837f
C13623 net80 _098_ 1.289178f
C13624 _352_/a_49_472# mask\[7\] 0.001066f
C13625 _058_ net21 0.004383f
C13626 FILLER_0_16_107/a_124_375# FILLER_0_16_89/a_1468_375# 0.005439f
C13627 FILLER_0_17_200/a_572_375# _093_ 0.002355f
C13628 FILLER_0_18_100/a_36_472# FILLER_0_17_72/a_3172_472# 0.05841f
C13629 _033_ net67 0.148585f
C13630 net22 vdd 1.920713f
C13631 _440_/a_796_472# net47 0.002508f
C13632 FILLER_0_18_61/a_124_375# FILLER_0_18_53/a_572_375# 0.012001f
C13633 _412_/a_36_151# output48/a_224_472# 0.229574f
C13634 FILLER_0_14_107/a_1468_375# vdd 0.007687f
C13635 net57 net37 0.091923f
C13636 _152_ _062_ 0.097086f
C13637 FILLER_0_9_72/a_932_472# vss 0.007033f
C13638 FILLER_0_9_72/a_1380_472# vdd 0.007659f
C13639 output34/a_224_472# net19 0.001308f
C13640 _448_/a_36_151# FILLER_0_2_177/a_124_375# 0.001597f
C13641 _114_ FILLER_0_12_136/a_36_472# 0.003953f
C13642 _420_/a_36_151# FILLER_0_23_282/a_484_472# 0.001723f
C13643 _389_/a_36_148# FILLER_0_10_94/a_36_472# 0.001723f
C13644 FILLER_0_22_177/a_124_375# net33 0.013581f
C13645 _093_ FILLER_0_18_139/a_1380_472# 0.007013f
C13646 cal_itt\[3\] _375_/a_1612_497# 0.003901f
C13647 FILLER_0_16_107/a_572_375# net14 0.002308f
C13648 net15 FILLER_0_9_60/a_572_375# 0.047331f
C13649 net1 vss 0.161208f
C13650 FILLER_0_10_78/a_484_472# net52 0.004421f
C13651 _085_ _113_ 0.084246f
C13652 _119_ _120_ 0.036534f
C13653 _115_ _069_ 0.022355f
C13654 _410_/a_36_68# _173_ 0.009636f
C13655 net31 net33 0.002465f
C13656 _453_/a_2560_156# vss 0.00337f
C13657 _122_ _059_ 0.190023f
C13658 _015_ _426_/a_2560_156# 0.024461f
C13659 input5/a_36_113# net5 0.061819f
C13660 net2 input4/a_36_68# 0.031809f
C13661 FILLER_0_18_2/a_1020_375# net44 0.009108f
C13662 net33 _435_/a_2665_112# 0.005831f
C13663 ctln[7] ctln[8] 0.004643f
C13664 _221_/a_36_160# _054_ 0.02124f
C13665 net78 _109_ 0.001432f
C13666 _402_/a_1296_93# cal_count\[1\] 0.004472f
C13667 net75 _416_/a_2665_112# 0.001785f
C13668 _136_ FILLER_0_16_154/a_36_472# 0.00615f
C13669 _428_/a_448_472# _131_ 0.041178f
C13670 _443_/a_2665_112# net59 0.0434f
C13671 _059_ _227_/a_36_160# 0.099735f
C13672 net62 _099_ 0.062012f
C13673 FILLER_0_7_72/a_1468_375# vdd 0.001135f
C13674 _238_/a_67_603# trim_mask\[3\] 0.028437f
C13675 FILLER_0_16_89/a_36_472# _040_ 0.015634f
C13676 _072_ _228_/a_36_68# 0.005788f
C13677 vss _433_/a_2248_156# 0.034403f
C13678 vdd _433_/a_2665_112# 0.002569f
C13679 mask\[0\] _429_/a_2665_112# 0.016053f
C13680 _087_ _079_ 0.251042f
C13681 FILLER_0_21_125/a_484_472# FILLER_0_22_128/a_36_472# 0.026657f
C13682 net74 FILLER_0_2_111/a_1468_375# 0.003854f
C13683 net27 _015_ 0.103416f
C13684 _111_ FILLER_0_18_76/a_36_472# 0.006706f
C13685 FILLER_0_3_172/a_2812_375# net22 0.013048f
C13686 _308_/a_848_380# vss 0.043591f
C13687 FILLER_0_18_53/a_484_472# vss 0.003579f
C13688 _094_ _418_/a_1204_472# 0.009231f
C13689 _256_/a_36_68# _058_ 0.001402f
C13690 FILLER_0_17_133/a_36_472# vss 0.006791f
C13691 _189_/a_67_603# vss 0.004088f
C13692 net54 _050_ 0.040506f
C13693 _422_/a_36_151# mask\[7\] 0.043316f
C13694 FILLER_0_17_72/a_932_472# net71 0.001418f
C13695 _285_/a_36_472# _045_ 0.00269f
C13696 _052_ FILLER_0_21_60/a_124_375# 0.002308f
C13697 FILLER_0_16_57/a_932_472# _131_ 0.007885f
C13698 _086_ _267_/a_36_472# 0.070088f
C13699 _221_/a_36_160# vss 0.037067f
C13700 FILLER_0_9_60/a_572_375# net51 0.002279f
C13701 _078_ FILLER_0_6_231/a_36_472# 0.013046f
C13702 FILLER_0_21_133/a_36_472# FILLER_0_21_142/a_36_472# 0.001963f
C13703 _413_/a_36_151# FILLER_0_1_192/a_36_472# 0.046516f
C13704 _004_ _416_/a_2665_112# 0.002631f
C13705 net36 FILLER_0_16_115/a_36_472# 0.003805f
C13706 _379_/a_36_472# trim_val\[1\] 0.00909f
C13707 _321_/a_2034_472# _176_ 0.002722f
C13708 _069_ _395_/a_36_488# 0.042974f
C13709 _445_/a_1000_472# net40 0.015508f
C13710 _256_/a_3368_68# _076_ 0.001183f
C13711 net2 _001_ 0.081616f
C13712 _105_ result[6] 0.001477f
C13713 FILLER_0_10_28/a_36_472# vss 0.001102f
C13714 FILLER_0_15_235/a_124_375# vss 0.001993f
C13715 _432_/a_36_151# _097_ 0.003144f
C13716 FILLER_0_15_235/a_572_375# vdd -0.005887f
C13717 result[0] vss 0.291352f
C13718 fanout63/a_36_160# mask\[2\] 0.026642f
C13719 _053_ FILLER_0_5_54/a_36_472# 0.003309f
C13720 FILLER_0_9_105/a_36_472# vdd 0.009746f
C13721 FILLER_0_9_105/a_572_375# vss 0.020145f
C13722 FILLER_0_8_138/a_36_472# vdd 0.008749f
C13723 FILLER_0_13_142/a_36_472# _043_ 0.011974f
C13724 net81 _094_ 0.004737f
C13725 FILLER_0_20_177/a_36_472# vss 0.003944f
C13726 FILLER_0_20_177/a_484_472# vdd 0.010805f
C13727 net81 _425_/a_2248_156# 0.058229f
C13728 ctlp[3] output21/a_224_472# 0.021951f
C13729 FILLER_0_16_107/a_484_472# FILLER_0_16_115/a_36_472# 0.013276f
C13730 _126_ net79 0.085443f
C13731 FILLER_0_4_197/a_36_472# net76 0.003914f
C13732 FILLER_0_5_54/a_124_375# FILLER_0_6_47/a_932_472# 0.001597f
C13733 FILLER_0_16_57/a_124_375# FILLER_0_17_56/a_124_375# 0.026339f
C13734 _192_/a_67_603# vdd 0.027014f
C13735 FILLER_0_16_73/a_36_472# FILLER_0_15_72/a_36_472# 0.026657f
C13736 output16/a_224_472# _447_/a_2248_156# 0.001937f
C13737 net16 _447_/a_1000_472# 0.003207f
C13738 _013_ FILLER_0_21_28/a_1916_375# 0.006025f
C13739 FILLER_0_15_142/a_124_375# _136_ 0.001706f
C13740 net36 FILLER_0_15_212/a_1020_375# 0.004863f
C13741 _176_ _318_/a_224_472# 0.003019f
C13742 FILLER_0_2_165/a_124_375# net22 0.206491f
C13743 FILLER_0_18_107/a_572_375# vdd 0.00419f
C13744 FILLER_0_18_107/a_124_375# vss 0.003425f
C13745 _434_/a_36_151# _348_/a_49_472# 0.017459f
C13746 net20 vdd 2.14128f
C13747 _267_/a_224_472# _121_ 0.0029f
C13748 _422_/a_796_472# vdd 0.003546f
C13749 cal_count\[2\] _452_/a_3129_107# 0.008853f
C13750 _062_ _113_ 0.020368f
C13751 _106_ FILLER_0_17_218/a_572_375# 0.022684f
C13752 state\[2\] _071_ 0.04575f
C13753 net79 FILLER_0_12_220/a_572_375# 0.010889f
C13754 _441_/a_1000_472# vss 0.01858f
C13755 _242_/a_36_160# _386_/a_124_24# 0.031797f
C13756 _411_/a_1308_423# net8 0.0176f
C13757 _232_/a_67_603# _164_ 0.076123f
C13758 net55 _424_/a_1000_472# 0.001357f
C13759 _413_/a_2248_156# net21 0.009186f
C13760 mask\[3\] _092_ 0.040554f
C13761 _064_ _446_/a_2560_156# 0.029586f
C13762 _432_/a_36_151# mask\[2\] 0.031341f
C13763 FILLER_0_5_117/a_36_472# _154_ 0.005034f
C13764 net32 _295_/a_36_472# 0.002637f
C13765 _430_/a_2248_156# vdd 0.008989f
C13766 net76 _080_ 0.03728f
C13767 _447_/a_36_151# net68 0.040925f
C13768 _411_/a_2248_156# net19 0.001197f
C13769 _372_/a_358_69# _160_ 0.001562f
C13770 _415_/a_1204_472# _004_ 0.002391f
C13771 net53 FILLER_0_16_154/a_36_472# 0.006261f
C13772 _125_ vss 0.149512f
C13773 _024_ _147_ 0.006801f
C13774 FILLER_0_5_128/a_484_472# FILLER_0_5_136/a_36_472# 0.013276f
C13775 _091_ _140_ 0.006511f
C13776 _318_/a_224_472# _124_ 0.001288f
C13777 _131_ FILLER_0_17_104/a_1020_375# 0.006574f
C13778 FILLER_0_6_239/a_36_472# vss 0.003177f
C13779 ctlp[1] _421_/a_2665_112# 0.008695f
C13780 _130_ FILLER_0_12_136/a_36_472# 0.082451f
C13781 _430_/a_2248_156# net20 0.001893f
C13782 FILLER_0_17_200/a_124_375# mask\[3\] 0.01841f
C13783 net15 _423_/a_448_472# 0.004833f
C13784 FILLER_0_21_28/a_1468_375# _423_/a_36_151# 0.001543f
C13785 _226_/a_860_68# net21 0.00107f
C13786 _101_ _045_ 0.001111f
C13787 net41 _181_ 0.043679f
C13788 _449_/a_448_472# _038_ 0.064169f
C13789 FILLER_0_3_172/a_2812_375# vdd -0.012025f
C13790 FILLER_0_5_54/a_1020_375# _440_/a_36_151# 0.059049f
C13791 _359_/a_1044_488# _133_ 0.001894f
C13792 _359_/a_1492_488# _070_ 0.0043f
C13793 _359_/a_36_488# _076_ 0.005184f
C13794 FILLER_0_15_212/a_1468_375# FILLER_0_15_228/a_124_375# 0.012001f
C13795 net63 FILLER_0_20_177/a_1380_472# 0.011079f
C13796 result[6] _420_/a_1204_472# 0.002681f
C13797 _431_/a_1308_423# net73 0.039024f
C13798 FILLER_0_7_104/a_124_375# _058_ 0.006125f
C13799 FILLER_0_20_31/a_36_472# FILLER_0_20_15/a_1380_472# 0.013276f
C13800 _052_ FILLER_0_18_37/a_124_375# 0.03242f
C13801 _251_/a_906_472# vss 0.0016f
C13802 _104_ ctlp[2] 1.420577f
C13803 _163_ FILLER_0_5_136/a_36_472# 0.007779f
C13804 net81 FILLER_0_8_263/a_36_472# 0.007373f
C13805 _267_/a_36_472# _090_ 0.001109f
C13806 FILLER_0_21_286/a_124_375# _420_/a_36_151# 0.001597f
C13807 net9 vdd 0.190349f
C13808 result[1] net79 0.25261f
C13809 net36 FILLER_0_15_205/a_36_472# 0.005101f
C13810 _127_ net23 0.069001f
C13811 FILLER_0_15_142/a_36_472# _427_/a_36_151# 0.001723f
C13812 net81 FILLER_0_14_235/a_572_375# 0.029643f
C13813 net15 FILLER_0_17_72/a_484_472# 0.002925f
C13814 output21/a_224_472# _108_ 0.005356f
C13815 output17/a_224_472# vdd 0.026649f
C13816 vss _416_/a_1000_472# 0.001784f
C13817 _422_/a_1204_472# _108_ 0.015401f
C13818 output46/a_224_472# vss 0.00432f
C13819 mask\[4\] net54 0.009909f
C13820 _277_/a_36_160# _094_ 0.007538f
C13821 FILLER_0_5_109/a_36_472# vdd 0.042799f
C13822 _135_ vdd 0.018662f
C13823 FILLER_0_13_65/a_36_472# cal_count\[1\] 0.016393f
C13824 net57 _390_/a_36_68# 0.001112f
C13825 _105_ _422_/a_36_151# 0.030571f
C13826 net13 _170_ 0.001668f
C13827 state\[2\] _095_ 0.001426f
C13828 FILLER_0_11_142/a_572_375# cal_count\[3\] 0.014082f
C13829 _053_ FILLER_0_6_79/a_36_472# 0.001777f
C13830 _086_ FILLER_0_7_104/a_1380_472# 0.034829f
C13831 FILLER_0_22_177/a_572_375# mask\[6\] 0.002657f
C13832 net35 FILLER_0_22_177/a_124_375# 0.0073f
C13833 _098_ _434_/a_2665_112# 0.013854f
C13834 net15 trim_mask\[1\] 0.042093f
C13835 net15 output16/a_224_472# 0.013768f
C13836 FILLER_0_15_142/a_124_375# net53 0.033224f
C13837 FILLER_0_6_79/a_124_375# FILLER_0_6_47/a_3260_375# 0.012001f
C13838 _176_ FILLER_0_11_78/a_124_375# 0.004803f
C13839 net79 FILLER_0_12_236/a_484_472# 0.009305f
C13840 net54 mask\[9\] 0.094381f
C13841 _077_ FILLER_0_10_78/a_36_472# 0.002486f
C13842 _175_ _095_ 0.041931f
C13843 FILLER_0_18_2/a_2812_375# FILLER_0_19_28/a_36_472# 0.001684f
C13844 _434_/a_796_472# _023_ 0.002118f
C13845 FILLER_0_2_165/a_124_375# vdd 0.020315f
C13846 FILLER_0_4_49/a_124_375# net49 0.005427f
C13847 FILLER_0_4_49/a_484_472# net66 0.015555f
C13848 FILLER_0_5_198/a_572_375# net22 0.029657f
C13849 _140_ FILLER_0_22_128/a_3260_375# 0.003524f
C13850 _140_ net33 0.026401f
C13851 fanout67/a_36_160# vdd 0.018829f
C13852 _174_ cal_count\[3\] 0.053844f
C13853 net35 _435_/a_2665_112# 0.007912f
C13854 FILLER_0_4_185/a_124_375# _002_ 0.013895f
C13855 result[6] _419_/a_2248_156# 0.002634f
C13856 mask\[5\] ctlp[2] 0.104304f
C13857 trim_mask\[1\] FILLER_0_6_90/a_572_375# 0.001263f
C13858 FILLER_0_17_161/a_36_472# vss 0.003343f
C13859 output43/a_224_472# output46/a_224_472# 0.292611f
C13860 net69 net14 0.056927f
C13861 cal_count\[2\] _278_/a_36_160# 0.023061f
C13862 _018_ _043_ 0.0022f
C13863 FILLER_0_15_290/a_36_472# _417_/a_36_151# 0.027236f
C13864 cal en 0.482495f
C13865 net15 _447_/a_2665_112# 0.063341f
C13866 _323_/a_36_113# FILLER_0_10_247/a_124_375# 0.001846f
C13867 FILLER_0_14_107/a_36_472# _043_ 0.001661f
C13868 net79 state\[1\] 0.005861f
C13869 net73 _093_ 0.350073f
C13870 _370_/a_124_24# _160_ 0.001126f
C13871 net15 mask\[9\] 0.128816f
C13872 _165_ _160_ 0.008705f
C13873 _069_ net22 0.327999f
C13874 cal_count\[2\] vss 0.361185f
C13875 _178_ cal_count\[2\] 0.119443f
C13876 net69 _164_ 0.040362f
C13877 FILLER_0_11_101/a_572_375# FILLER_0_11_109/a_36_472# 0.086635f
C13878 net79 _007_ 0.096772f
C13879 _093_ FILLER_0_21_60/a_572_375# 0.011177f
C13880 FILLER_0_10_78/a_36_472# _120_ 0.004669f
C13881 _013_ _424_/a_448_472# 0.043803f
C13882 net72 FILLER_0_12_50/a_36_472# 0.002007f
C13883 _420_/a_1308_423# vdd 0.00284f
C13884 _420_/a_448_472# vss 0.007371f
C13885 _095_ FILLER_0_14_107/a_1020_375# 0.014156f
C13886 _094_ _045_ 0.102437f
C13887 net19 _416_/a_2665_112# 0.059453f
C13888 _086_ FILLER_0_4_177/a_124_375# 0.024433f
C13889 _053_ _077_ 0.123663f
C13890 net4 FILLER_0_12_220/a_1020_375# 0.020782f
C13891 input3/a_36_113# vss 0.043862f
C13892 cal input1/a_36_113# 0.025739f
C13893 FILLER_0_19_47/a_36_472# _052_ 0.015772f
C13894 _057_ _311_/a_1212_473# 0.004869f
C13895 _398_/a_36_113# net3 0.099638f
C13896 output46/a_224_472# net46 0.008691f
C13897 _444_/a_36_151# net67 0.055072f
C13898 _177_ _451_/a_3129_107# 0.043731f
C13899 net72 _394_/a_56_524# 0.066156f
C13900 FILLER_0_19_28/a_484_472# vss 0.001207f
C13901 net52 _443_/a_36_151# 0.020518f
C13902 valid _425_/a_2248_156# 0.00154f
C13903 result[9] ctlp[1] 0.074012f
C13904 net47 _365_/a_692_472# 0.002051f
C13905 trimb[1] FILLER_0_20_2/a_484_472# 0.003628f
C13906 ctln[7] net14 0.197449f
C13907 _446_/a_2248_156# net66 0.002766f
C13908 net76 vss 0.436111f
C13909 net44 _450_/a_36_151# 0.026203f
C13910 vss _450_/a_448_472# -0.001661f
C13911 FILLER_0_9_28/a_1916_375# _220_/a_67_603# 0.014522f
C13912 cal_count\[3\] _373_/a_1254_68# 0.001391f
C13913 FILLER_0_16_241/a_124_375# net30 0.028559f
C13914 net27 _415_/a_36_151# 0.019856f
C13915 _087_ FILLER_0_6_177/a_124_375# 0.001151f
C13916 _412_/a_448_472# cal_itt\[1\] 0.043203f
C13917 FILLER_0_19_28/a_36_472# FILLER_0_20_15/a_1380_472# 0.026657f
C13918 _322_/a_124_24# _070_ 0.033355f
C13919 _423_/a_2665_112# vss 0.016881f
C13920 _411_/a_2560_156# net8 0.013106f
C13921 FILLER_0_4_152/a_36_472# vdd 0.087397f
C13922 FILLER_0_8_138/a_124_375# _129_ 0.006506f
C13923 FILLER_0_16_89/a_932_472# vdd 0.002218f
C13924 FILLER_0_16_89/a_484_472# vss -0.001894f
C13925 _283_/a_36_472# vdd 0.092097f
C13926 trim_mask\[4\] _031_ 0.001262f
C13927 net40 _160_ 0.152292f
C13928 _076_ FILLER_0_8_156/a_572_375# 0.010751f
C13929 _074_ _265_/a_224_472# 0.001223f
C13930 FILLER_0_20_193/a_572_375# _098_ 0.078973f
C13931 FILLER_0_20_177/a_124_375# _434_/a_36_151# 0.059049f
C13932 _185_ cal_count\[1\] 0.001949f
C13933 FILLER_0_16_154/a_124_375# vss 0.004317f
C13934 FILLER_0_16_154/a_572_375# vdd 0.004706f
C13935 net31 net22 0.002533f
C13936 _448_/a_36_151# FILLER_0_1_192/a_36_472# 0.008172f
C13937 _253_/a_1100_68# _074_ 0.001563f
C13938 _150_ vss 0.016993f
C13939 _424_/a_36_151# _423_/a_36_151# 0.006746f
C13940 FILLER_0_20_193/a_572_375# _205_/a_36_160# 0.002828f
C13941 FILLER_0_4_49/a_36_472# _164_ 0.033727f
C13942 _440_/a_36_151# FILLER_0_6_47/a_3172_472# 0.001653f
C13943 output20/a_224_472# vdd 0.09529f
C13944 _105_ _291_/a_36_160# 0.002075f
C13945 FILLER_0_17_72/a_3172_472# vss 0.001338f
C13946 _083_ _265_/a_244_68# 0.004022f
C13947 _421_/a_36_151# _010_ 0.015107f
C13948 _389_/a_36_148# _171_ 0.023988f
C13949 net22 _435_/a_2665_112# 0.004214f
C13950 _431_/a_2248_156# vss 0.041929f
C13951 FILLER_0_5_198/a_572_375# vdd 0.005402f
C13952 FILLER_0_22_86/a_1468_375# net14 0.024975f
C13953 _106_ mask\[4\] 0.091207f
C13954 _132_ FILLER_0_18_107/a_1828_472# 0.045833f
C13955 _004_ result[1] 0.005653f
C13956 _432_/a_2248_156# mask\[3\] 0.002775f
C13957 _119_ _125_ 0.11554f
C13958 _043_ _278_/a_36_160# 0.004357f
C13959 ctln[5] _448_/a_1204_472# 0.005186f
C13960 FILLER_0_4_123/a_36_472# _153_ 0.001419f
C13961 output20/a_224_472# net20 0.024692f
C13962 ctln[2] net4 0.039098f
C13963 _093_ _131_ 0.254316f
C13964 FILLER_0_2_177/a_124_375# vss 0.00252f
C13965 FILLER_0_2_177/a_572_375# vdd 0.022268f
C13966 FILLER_0_5_109/a_484_472# FILLER_0_5_117/a_36_472# 0.013276f
C13967 net19 _420_/a_1000_472# 0.006558f
C13968 _372_/a_3126_472# _068_ 0.005304f
C13969 net74 FILLER_0_13_72/a_484_472# 0.007142f
C13970 trimb[0] net43 0.109028f
C13971 net27 net62 0.008623f
C13972 _043_ vss 1.362912f
C13973 _178_ _043_ 0.130207f
C13974 _211_/a_36_160# net14 0.005761f
C13975 _000_ _080_ 0.002867f
C13976 net68 _054_ 0.08092f
C13977 _292_/a_36_160# net32 0.011466f
C13978 _449_/a_1308_423# _453_/a_2665_112# 0.001066f
C13979 output35/a_224_472# vss 0.01667f
C13980 net34 ctlp[2] 0.953441f
C13981 mask\[3\] FILLER_0_18_177/a_2276_472# 0.01204f
C13982 _069_ vdd 0.985405f
C13983 result[9] FILLER_0_24_274/a_124_375# 0.008195f
C13984 _139_ net36 0.024268f
C13985 sample en 0.001572f
C13986 FILLER_0_13_212/a_124_375# net79 0.007396f
C13987 _016_ _129_ 0.002216f
C13988 net62 FILLER_0_13_212/a_572_375# 0.001597f
C13989 net76 fanout76/a_36_160# 0.004503f
C13990 _377_/a_36_472# _164_ 0.03259f
C13991 net73 _136_ 0.050578f
C13992 result[6] output18/a_224_472# 0.003068f
C13993 net4 FILLER_0_3_221/a_572_375# 0.030599f
C13994 mask\[7\] _435_/a_1000_472# 0.024725f
C13995 result[8] _422_/a_36_151# 0.001488f
C13996 ctln[1] net4 0.009703f
C13997 mask\[5\] net21 0.212814f
C13998 FILLER_0_9_28/a_2724_472# _453_/a_448_472# 0.008036f
C13999 _147_ mask\[6\] 0.103475f
C14000 _143_ _339_/a_36_160# 0.00507f
C14001 mask\[3\] FILLER_0_17_218/a_36_472# 0.015535f
C14002 _131_ FILLER_0_14_123/a_36_472# 0.029747f
C14003 _272_/a_36_472# _079_ 0.0237f
C14004 _091_ FILLER_0_13_228/a_36_472# 0.001826f
C14005 net68 vss 0.635359f
C14006 net25 FILLER_0_22_86/a_36_472# 0.001265f
C14007 cal_itt\[0\] net8 0.026229f
C14008 _110_ net71 0.004816f
C14009 mask\[5\] FILLER_0_19_171/a_932_472# 0.007596f
C14010 _026_ vss 0.005992f
C14011 _430_/a_2248_156# _069_ 0.042876f
C14012 net23 FILLER_0_22_128/a_2724_472# 0.054521f
C14013 net50 _447_/a_448_472# 0.001219f
C14014 output44/a_224_472# trimb[1] 0.046391f
C14015 _413_/a_448_472# vdd 0.016117f
C14016 _426_/a_1308_423# calibrate 0.001708f
C14017 FILLER_0_18_139/a_1468_375# vss 0.009191f
C14018 FILLER_0_18_139/a_36_472# vdd 0.089771f
C14019 FILLER_0_7_72/a_932_472# FILLER_0_6_79/a_124_375# 0.001723f
C14020 output36/a_224_472# FILLER_0_15_282/a_36_472# 0.008834f
C14021 _408_/a_718_524# _067_ 0.006516f
C14022 _093_ net56 0.040124f
C14023 FILLER_0_9_72/a_484_472# _439_/a_36_151# 0.001723f
C14024 FILLER_0_15_282/a_572_375# net18 0.00298f
C14025 net54 _022_ 0.004106f
C14026 FILLER_0_18_107/a_36_472# mask\[9\] 0.005458f
C14027 FILLER_0_22_177/a_124_375# vdd 0.001293f
C14028 FILLER_0_15_282/a_36_472# net30 0.001692f
C14029 FILLER_0_15_282/a_124_375# result[3] 0.004601f
C14030 cal_count\[2\] _184_ 0.033241f
C14031 trim_val\[3\] _441_/a_448_472# 0.00469f
C14032 _390_/a_244_472# _136_ 0.001777f
C14033 cal_count\[2\] _401_/a_36_68# 0.008136f
C14034 vss _156_ 0.089339f
C14035 _431_/a_36_151# net73 0.015086f
C14036 _426_/a_448_472# net64 0.054931f
C14037 _198_/a_67_603# net30 0.017304f
C14038 _064_ trim[1] 0.166575f
C14039 net31 vdd 0.542738f
C14040 _430_/a_2665_112# mask\[1\] 0.004574f
C14041 FILLER_0_12_136/a_1468_375# FILLER_0_13_142/a_932_472# 0.001684f
C14042 _104_ mask\[7\] 0.069172f
C14043 net67 _054_ 0.391592f
C14044 _439_/a_36_151# _453_/a_2665_112# 0.001738f
C14045 result[5] _007_ 0.0249f
C14046 _095_ _280_/a_224_472# 0.001416f
C14047 net35 _140_ 0.12583f
C14048 _308_/a_124_24# net14 0.005016f
C14049 net71 _437_/a_2665_112# 0.039687f
C14050 _081_ _265_/a_224_472# 0.008598f
C14051 _435_/a_2665_112# vdd 0.01769f
C14052 FILLER_0_17_72/a_3260_375# net14 0.040606f
C14053 _136_ _451_/a_1040_527# 0.00497f
C14054 _187_ _181_ 0.001158f
C14055 _449_/a_36_151# vdd 0.09324f
C14056 _210_/a_67_603# net23 0.005398f
C14057 net31 net20 0.238809f
C14058 _303_/a_36_472# FILLER_0_20_87/a_36_472# 0.005725f
C14059 _079_ _001_ 0.082209f
C14060 fanout65/a_36_113# vss 0.053899f
C14061 _443_/a_796_472# net23 0.002306f
C14062 _443_/a_448_472# net13 0.002263f
C14063 net28 vdd 0.489756f
C14064 net28 _192_/a_67_603# 0.119061f
C14065 _057_ cal_count\[3\] 0.416063f
C14066 _392_/a_36_68# cal_count\[0\] 0.038691f
C14067 _149_ _437_/a_448_472# 0.009274f
C14068 FILLER_0_8_127/a_124_375# vdd 0.019587f
C14069 net67 vss 0.435869f
C14070 _114_ _306_/a_36_68# 0.032258f
C14071 FILLER_0_9_28/a_1380_472# vdd 0.01306f
C14072 FILLER_0_11_124/a_36_472# _120_ 0.014712f
C14073 _131_ _136_ 1.42765f
C14074 ctln[4] vss 0.244634f
C14075 trim_val\[4\] _443_/a_2665_112# 0.018733f
C14076 cal_itt\[2\] vdd 0.267121f
C14077 _415_/a_36_151# net18 0.015992f
C14078 FILLER_0_21_125/a_484_472# vss 0.002399f
C14079 net41 _446_/a_2248_156# 0.016492f
C14080 net21 FILLER_0_12_196/a_124_375# 0.005374f
C14081 _176_ _172_ 0.043154f
C14082 _031_ _154_ 0.037238f
C14083 net69 _153_ 0.003678f
C14084 _114_ _115_ 0.148291f
C14085 FILLER_0_20_193/a_484_472# FILLER_0_18_177/a_2364_375# 0.0027f
C14086 sample output27/a_224_472# 0.006116f
C14087 _415_/a_2665_112# vdd 0.017004f
C14088 _053_ _363_/a_36_68# 0.021227f
C14089 net72 _182_ 0.044895f
C14090 ctln[3] _411_/a_36_151# 0.004014f
C14091 _053_ _003_ 0.021223f
C14092 net50 FILLER_0_8_24/a_124_375# 0.001597f
C14093 FILLER_0_11_64/a_36_472# vss 0.006069f
C14094 net80 net21 0.016911f
C14095 output13/a_224_472# _448_/a_2665_112# 0.027303f
C14096 FILLER_0_24_290/a_36_472# FILLER_0_23_290/a_36_472# 0.05841f
C14097 net73 net53 0.094507f
C14098 _132_ _428_/a_1308_423# 0.027389f
C14099 FILLER_0_12_236/a_572_375# vdd 0.024713f
C14100 FILLER_0_12_236/a_124_375# vss 0.001024f
C14101 net80 _333_/a_36_160# 0.001594f
C14102 net20 cal_itt\[2\] 0.715447f
C14103 mask\[5\] mask\[7\] 0.014384f
C14104 _376_/a_36_160# FILLER_0_5_72/a_1380_472# 0.035111f
C14105 net71 net14 0.147175f
C14106 FILLER_0_14_91/a_572_375# vdd -0.011429f
C14107 net63 FILLER_0_22_177/a_1020_375# 0.003419f
C14108 _442_/a_448_472# _031_ 0.019293f
C14109 _445_/a_1308_423# vdd 0.001478f
C14110 FILLER_0_21_28/a_932_472# vdd 0.04815f
C14111 FILLER_0_18_209/a_484_472# vss 0.005794f
C14112 net27 net4 0.025834f
C14113 net50 FILLER_0_2_93/a_572_375# 0.00275f
C14114 net52 FILLER_0_2_93/a_484_472# 0.009006f
C14115 _246_/a_36_68# _090_ 0.001712f
C14116 _077_ cal_count\[0\] 0.018501f
C14117 _423_/a_448_472# _012_ 0.038928f
C14118 _429_/a_36_151# _136_ 0.001188f
C14119 FILLER_0_13_65/a_124_375# vss 0.030194f
C14120 net41 _423_/a_36_151# 0.001134f
C14121 net34 net21 0.036237f
C14122 _104_ _422_/a_2248_156# 0.041703f
C14123 _000_ vss 0.205593f
C14124 _001_ cal_itt\[1\] 0.057933f
C14125 _152_ _153_ 0.002954f
C14126 _431_/a_36_151# _131_ 0.03645f
C14127 _074_ _084_ 0.110937f
C14128 FILLER_0_8_239/a_36_472# calibrate 0.008683f
C14129 net54 _437_/a_2248_156# 0.046559f
C14130 _013_ _217_/a_36_160# 0.001614f
C14131 FILLER_0_21_28/a_1020_375# _424_/a_36_151# 0.001252f
C14132 net76 FILLER_0_5_198/a_36_472# 0.003987f
C14133 FILLER_0_12_136/a_1380_472# state\[2\] 0.005779f
C14134 net62 net18 0.089041f
C14135 net15 net66 0.006618f
C14136 FILLER_0_14_50/a_124_375# cal_count\[1\] 0.023752f
C14137 net56 _136_ 0.462275f
C14138 _068_ _315_/a_716_497# 0.00217f
C14139 _076_ _315_/a_36_68# 0.001568f
C14140 _070_ _315_/a_1657_68# 0.001601f
C14141 net3 _190_/a_36_160# 0.013324f
C14142 _095_ cal_count\[2\] 0.270066f
C14143 output38/a_224_472# trim[1] 0.003114f
C14144 net38 net39 0.066083f
C14145 result[1] net19 0.084617f
C14146 net15 _067_ 0.042278f
C14147 trim_mask\[1\] net47 0.306848f
C14148 FILLER_0_12_20/a_484_472# net17 0.05005f
C14149 net77 vdd 0.526632f
C14150 _114_ _395_/a_36_488# 0.005314f
C14151 net62 _196_/a_36_160# 0.029171f
C14152 trim_val\[2\] net49 0.00301f
C14153 net76 FILLER_0_2_177/a_36_472# 0.003526f
C14154 output28/a_224_472# _416_/a_2665_112# 0.008243f
C14155 _009_ FILLER_0_23_282/a_484_472# 0.009744f
C14156 output14/a_224_472# _442_/a_2665_112# 0.009771f
C14157 net16 _450_/a_2225_156# 0.001015f
C14158 _150_ _027_ 0.006689f
C14159 FILLER_0_16_73/a_36_472# FILLER_0_17_72/a_124_375# 0.001723f
C14160 _112_ _425_/a_448_472# 0.002335f
C14161 net55 cal_count\[1\] 0.204733f
C14162 FILLER_0_18_2/a_1380_472# net38 0.029747f
C14163 FILLER_0_16_57/a_572_375# _176_ 0.006422f
C14164 net53 _451_/a_1040_527# 0.023651f
C14165 result[6] _421_/a_1000_472# 0.024206f
C14166 _120_ cal_count\[0\] 0.014209f
C14167 _131_ FILLER_0_17_56/a_572_375# 0.006224f
C14168 net16 _183_ 0.001103f
C14169 FILLER_0_15_116/a_36_472# FILLER_0_17_104/a_1468_375# 0.001512f
C14170 _114_ FILLER_0_13_142/a_1468_375# 0.001931f
C14171 _425_/a_2560_156# net37 0.002508f
C14172 _102_ _006_ 0.006115f
C14173 _176_ _183_ 0.024038f
C14174 FILLER_0_5_128/a_572_375# _152_ 0.00813f
C14175 _412_/a_36_151# net18 0.011383f
C14176 output33/a_224_472# net33 0.151281f
C14177 _028_ vss 0.410396f
C14178 _095_ _450_/a_448_472# 0.001393f
C14179 _104_ _105_ 0.931514f
C14180 _118_ net23 0.108864f
C14181 FILLER_0_4_177/a_124_375# _163_ 0.004052f
C14182 net35 FILLER_0_21_150/a_36_472# 0.004456f
C14183 _103_ _102_ 0.392644f
C14184 _431_/a_36_151# net56 0.001371f
C14185 FILLER_0_9_28/a_1020_375# net68 0.004803f
C14186 FILLER_0_16_107/a_36_472# net36 0.001245f
C14187 _091_ _137_ 0.486022f
C14188 FILLER_0_9_142/a_124_375# _313_/a_67_603# 0.029786f
C14189 net53 _131_ 0.059223f
C14190 FILLER_0_14_81/a_36_472# vdd 0.00958f
C14191 FILLER_0_14_81/a_124_375# vss 0.03341f
C14192 net60 _418_/a_448_472# 0.055895f
C14193 result[2] vss 0.327009f
C14194 net29 mask\[1\] 0.023266f
C14195 _413_/a_2248_156# FILLER_0_1_212/a_36_472# 0.035805f
C14196 FILLER_0_4_152/a_124_375# vdd -0.001403f
C14197 _426_/a_1204_472# vdd 0.003412f
C14198 net80 mask\[7\] 0.020051f
C14199 net46 FILLER_0_21_28/a_484_472# 0.001795f
C14200 net82 _370_/a_848_380# 0.014538f
C14201 _439_/a_2248_156# trim_mask\[0\] 0.005416f
C14202 _140_ _433_/a_2665_112# 0.001108f
C14203 _098_ _438_/a_2248_156# 0.002798f
C14204 FILLER_0_9_290/a_124_375# vss 0.033914f
C14205 FILLER_0_9_290/a_36_472# vdd 0.094552f
C14206 FILLER_0_12_220/a_1380_472# _060_ 0.01563f
C14207 net61 FILLER_0_21_286/a_484_472# 0.001829f
C14208 _144_ net54 0.095482f
C14209 _176_ FILLER_0_15_59/a_572_375# 0.007169f
C14210 _065_ _447_/a_2560_156# 0.012523f
C14211 _415_/a_448_472# net79 0.001602f
C14212 ctln[6] net59 0.001267f
C14213 _028_ FILLER_0_7_72/a_36_472# 0.020625f
C14214 mask\[9\] _012_ 0.008145f
C14215 trim[4] vdd 0.198218f
C14216 net79 _417_/a_36_151# 0.082646f
C14217 output27/a_224_472# FILLER_0_9_282/a_572_375# 0.029138f
C14218 _132_ FILLER_0_17_104/a_1468_375# 0.051996f
C14219 _427_/a_1000_472# net74 0.009646f
C14220 _077_ _070_ 0.29321f
C14221 net55 FILLER_0_17_38/a_36_472# 0.010728f
C14222 net62 _417_/a_448_472# 0.011318f
C14223 net34 mask\[7\] 0.901671f
C14224 FILLER_0_10_78/a_1468_375# _308_/a_124_24# 0.001565f
C14225 _411_/a_2665_112# vss 0.00238f
C14226 FILLER_0_6_47/a_2364_375# vdd 0.015888f
C14227 FILLER_0_6_47/a_1916_375# vss 0.005279f
C14228 _328_/a_36_113# _070_ 0.016264f
C14229 _321_/a_3662_472# net74 0.00253f
C14230 ctlp[1] net78 0.025929f
C14231 _068_ FILLER_0_5_148/a_36_472# 0.003015f
C14232 _104_ _298_/a_224_472# 0.001731f
C14233 FILLER_0_9_223/a_572_375# calibrate 0.002082f
C14234 _291_/a_36_160# output18/a_224_472# 0.001175f
C14235 _095_ _043_ 2.807456f
C14236 net60 mask\[7\] 0.001053f
C14237 mask\[5\] _105_ 0.706158f
C14238 FILLER_0_15_142/a_484_472# net56 0.003214f
C14239 output15/a_224_472# trim_mask\[3\] 0.024718f
C14240 cal_count\[2\] _402_/a_1296_93# 0.022009f
C14241 FILLER_0_17_38/a_484_472# _182_ 0.00527f
C14242 _320_/a_36_472# FILLER_0_13_206/a_36_472# 0.038251f
C14243 net54 net23 0.084191f
C14244 _428_/a_2665_112# state\[2\] 0.001746f
C14245 _140_ vdd 0.598538f
C14246 _282_/a_36_160# vdd 0.010099f
C14247 net56 net53 0.053535f
C14248 FILLER_0_6_90/a_124_375# net14 0.005361f
C14249 _050_ _436_/a_1204_472# 0.006724f
C14250 _081_ _084_ 0.016804f
C14251 result[4] FILLER_0_15_290/a_36_472# 0.001422f
C14252 net80 mask\[1\] 0.015535f
C14253 _161_ _311_/a_1212_473# 0.004138f
C14254 _098_ mask\[6\] 0.297837f
C14255 mask\[8\] _098_ 0.096999f
C14256 vdd FILLER_0_6_231/a_484_472# 0.004642f
C14257 vss FILLER_0_6_231/a_36_472# 0.0048f
C14258 _421_/a_36_151# vss 0.021759f
C14259 _421_/a_448_472# vdd 0.030898f
C14260 _086_ _315_/a_36_68# 0.003329f
C14261 _070_ _120_ 0.838223f
C14262 net67 _450_/a_1040_527# 0.032098f
C14263 _038_ _070_ 0.075667f
C14264 FILLER_0_18_107/a_3172_472# vss 0.006614f
C14265 net20 _282_/a_36_160# 0.016884f
C14266 _136_ FILLER_0_15_180/a_36_472# 0.006924f
C14267 _435_/a_36_151# _434_/a_1308_423# 0.001518f
C14268 _424_/a_2665_112# vdd 0.013636f
C14269 _424_/a_2248_156# vss 0.004855f
C14270 net26 FILLER_0_23_44/a_572_375# 0.003172f
C14271 FILLER_0_1_192/a_36_472# vss 0.004422f
C14272 net32 net61 0.056005f
C14273 net41 _444_/a_2248_156# 0.028267f
C14274 _320_/a_1568_472# state\[1\] 0.001531f
C14275 net4 net18 0.034592f
C14276 net20 FILLER_0_6_231/a_484_472# 0.017025f
C14277 result[2] _416_/a_2248_156# 0.001396f
C14278 net55 FILLER_0_17_72/a_124_375# 0.019544f
C14279 net20 _421_/a_448_472# 0.015767f
C14280 net15 net25 0.013745f
C14281 net65 _084_ 0.031674f
C14282 _096_ _320_/a_36_472# 0.052438f
C14283 _114_ _308_/a_1084_68# 0.00178f
C14284 net50 _441_/a_2665_112# 0.056602f
C14285 output37/a_224_472# net76 0.004028f
C14286 net68 _036_ 0.168017f
C14287 FILLER_0_23_290/a_36_472# FILLER_0_23_282/a_484_472# 0.013276f
C14288 _412_/a_2665_112# net58 0.006815f
C14289 _053_ _251_/a_906_472# 0.001696f
C14290 net82 FILLER_0_3_212/a_124_375# 0.015932f
C14291 net34 _422_/a_2248_156# 0.005617f
C14292 trim_mask\[1\] _154_ 0.004835f
C14293 result[6] net18 0.026875f
C14294 FILLER_0_8_37/a_124_375# vdd 0.029725f
C14295 _049_ FILLER_0_22_128/a_3260_375# 0.16381f
C14296 FILLER_0_12_136/a_484_472# vss 0.007054f
C14297 FILLER_0_12_136/a_932_472# vdd 0.005266f
C14298 net25 FILLER_0_23_44/a_1380_472# 0.0014f
C14299 output10/a_224_472# net58 0.025878f
C14300 _269_/a_36_472# net59 0.011985f
C14301 _340_/a_36_160# FILLER_0_20_169/a_36_472# 0.195478f
C14302 _412_/a_2560_156# net5 0.007446f
C14303 FILLER_0_21_28/a_1468_375# _012_ 0.00351f
C14304 _074_ FILLER_0_6_177/a_484_472# 0.002068f
C14305 FILLER_0_16_73/a_36_472# _175_ 0.006803f
C14306 FILLER_0_5_72/a_1468_375# vdd 0.001826f
C14307 FILLER_0_5_72/a_1020_375# vss 0.004157f
C14308 net21 _434_/a_2665_112# 0.004945f
C14309 net41 FILLER_0_21_28/a_1020_375# 0.010649f
C14310 _397_/a_36_472# net36 0.010045f
C14311 _065_ ctln[8] 0.193903f
C14312 net69 FILLER_0_2_111/a_932_472# 0.011453f
C14313 net14 FILLER_0_4_91/a_484_472# 0.020589f
C14314 _031_ FILLER_0_2_111/a_36_472# 0.034656f
C14315 net55 _120_ 0.001054f
C14316 FILLER_0_12_136/a_572_375# FILLER_0_11_142/a_36_472# 0.001543f
C14317 net55 _038_ 0.05656f
C14318 en_co_clk _136_ 0.034892f
C14319 _050_ FILLER_0_22_128/a_572_375# 0.002607f
C14320 net61 _422_/a_2560_156# 0.010748f
C14321 _289_/a_36_472# net30 0.009623f
C14322 FILLER_0_5_54/a_1020_375# _029_ 0.024737f
C14323 _315_/a_1229_68# _121_ 0.003401f
C14324 _122_ FILLER_0_8_156/a_36_472# 0.047846f
C14325 _183_ _041_ 0.001931f
C14326 _441_/a_36_151# _440_/a_1308_423# 0.001736f
C14327 net38 clkc 0.088241f
C14328 _451_/a_36_151# vdd 0.088651f
C14329 _154_ _157_ 0.447829f
C14330 _114_ FILLER_0_9_72/a_1380_472# 0.001043f
C14331 FILLER_0_9_28/a_484_472# net51 0.001023f
C14332 FILLER_0_21_286/a_124_375# _009_ 0.001024f
C14333 _446_/a_796_472# net40 0.001504f
C14334 FILLER_0_4_197/a_36_472# _413_/a_36_151# 0.001512f
C14335 _426_/a_36_151# FILLER_0_8_247/a_1020_375# 0.059049f
C14336 _144_ _350_/a_49_472# 0.033348f
C14337 _227_/a_36_160# FILLER_0_8_156/a_36_472# 0.006647f
C14338 FILLER_0_16_255/a_36_472# vdd 0.044615f
C14339 _081_ FILLER_0_5_148/a_484_472# 0.016132f
C14340 FILLER_0_9_28/a_572_375# net40 0.001406f
C14341 _421_/a_796_472# net19 0.009462f
C14342 _308_/a_124_24# _439_/a_2665_112# 0.002245f
C14343 net57 _116_ 0.069858f
C14344 _008_ _418_/a_1000_472# 0.01006f
C14345 FILLER_0_2_93/a_572_375# FILLER_0_2_101/a_36_472# 0.086635f
C14346 _114_ _311_/a_2700_473# 0.005178f
C14347 _253_/a_244_68# _073_ 0.002878f
C14348 FILLER_0_14_91/a_36_472# _043_ 0.001779f
C14349 FILLER_0_11_124/a_124_375# vdd 0.016626f
C14350 _186_ _402_/a_728_93# 0.002381f
C14351 _104_ result[8] 0.00201f
C14352 _168_ _160_ 0.03261f
C14353 _170_ _386_/a_124_24# 0.008511f
C14354 net16 _445_/a_2665_112# 0.061595f
C14355 net50 FILLER_0_5_88/a_36_472# 0.00867f
C14356 FILLER_0_22_177/a_1380_472# _435_/a_36_151# 0.001723f
C14357 _432_/a_2665_112# _093_ 0.02266f
C14358 _035_ _446_/a_1000_472# 0.00349f
C14359 result[7] _046_ 0.003397f
C14360 _408_/a_56_524# FILLER_0_12_20/a_572_375# 0.009967f
C14361 _105_ net34 0.784678f
C14362 _004_ _415_/a_448_472# 0.044374f
C14363 net43 vdd 0.210686f
C14364 mask\[4\] FILLER_0_19_155/a_36_472# 0.047448f
C14365 net41 net39 0.003649f
C14366 _372_/a_170_472# _062_ 0.014919f
C14367 net70 FILLER_0_11_101/a_484_472# 0.001474f
C14368 FILLER_0_14_91/a_124_375# _095_ 0.01418f
C14369 FILLER_0_12_124/a_124_375# _127_ 0.003767f
C14370 _350_/a_49_472# net23 0.002397f
C14371 net41 net51 0.031531f
C14372 _127_ FILLER_0_9_142/a_36_472# 0.004721f
C14373 _105_ net60 0.042726f
C14374 net43 FILLER_0_20_15/a_484_472# 0.001534f
C14375 fanout79/a_36_160# _094_ 0.008308f
C14376 _102_ mask\[2\] 0.036292f
C14377 _419_/a_796_472# net77 0.001053f
C14378 _198_/a_67_603# _046_ 0.007349f
C14379 net81 FILLER_0_15_212/a_484_472# 0.00169f
C14380 net57 _118_ 0.036179f
C14381 net2 rstn 0.002598f
C14382 FILLER_0_13_65/a_124_375# _095_ 0.002035f
C14383 FILLER_0_21_150/a_36_472# vdd 0.092128f
C14384 FILLER_0_21_150/a_124_375# vss 0.013882f
C14385 FILLER_0_5_117/a_124_375# _160_ 0.008534f
C14386 _162_ _058_ 0.015239f
C14387 mask\[0\] FILLER_0_12_196/a_124_375# 0.034009f
C14388 fanout50/a_36_160# _383_/a_36_472# 0.096296f
C14389 _096_ _085_ 0.0099f
C14390 _078_ _080_ 0.030094f
C14391 net26 vss 0.263774f
C14392 _101_ _285_/a_244_68# 0.001153f
C14393 net29 _099_ 0.358926f
C14394 ctln[7] FILLER_0_0_96/a_36_472# 0.01317f
C14395 FILLER_0_11_101/a_572_375# FILLER_0_10_107/a_36_472# 0.001684f
C14396 _127_ _128_ 0.257374f
C14397 net55 FILLER_0_17_56/a_484_472# 0.023554f
C14398 FILLER_0_4_177/a_36_472# FILLER_0_3_172/a_484_472# 0.026657f
C14399 vdd output30/a_224_472# 0.068123f
C14400 _074_ net4 0.088616f
C14401 FILLER_0_7_72/a_484_472# vss 0.003793f
C14402 _053_ net76 0.022571f
C14403 _131_ _058_ 0.031061f
C14404 FILLER_0_24_63/a_124_375# vdd 0.029514f
C14405 net54 FILLER_0_19_134/a_124_375# 0.002681f
C14406 FILLER_0_12_50/a_124_375# vss 0.004123f
C14407 FILLER_0_12_50/a_36_472# vdd 0.012805f
C14408 _093_ FILLER_0_17_72/a_2812_375# 0.019521f
C14409 net38 net47 0.352245f
C14410 output9/a_224_472# net5 0.005189f
C14411 output28/a_224_472# result[1] 0.054333f
C14412 mask\[5\] result[8] 0.003797f
C14413 _428_/a_2248_156# vdd 0.006977f
C14414 _098_ _433_/a_2248_156# 0.034774f
C14415 FILLER_0_20_193/a_572_375# net21 0.002103f
C14416 net75 _317_/a_36_113# 0.030797f
C14417 net38 _450_/a_1284_156# 0.001291f
C14418 FILLER_0_17_64/a_124_375# _183_ 0.001236f
C14419 net4 _076_ 1.140706f
C14420 _437_/a_1000_472# net14 0.028506f
C14421 en_co_clk net53 0.001712f
C14422 trim_mask\[4\] _158_ 0.022724f
C14423 _394_/a_56_524# vdd 0.010692f
C14424 _394_/a_728_93# vss 0.024106f
C14425 _114_ vdd 1.30767f
C14426 _161_ cal_count\[3\] 0.047389f
C14427 _415_/a_796_472# net81 0.002008f
C14428 _449_/a_448_472# FILLER_0_11_64/a_36_472# 0.001462f
C14429 output21/a_224_472# _009_ 0.004164f
C14430 net55 _175_ 0.142124f
C14431 net52 _032_ 0.009879f
C14432 _081_ FILLER_0_6_177/a_484_472# 0.010037f
C14433 _408_/a_728_93# net40 0.084147f
C14434 _422_/a_1204_472# _009_ 0.009783f
C14435 net44 _039_ 0.15647f
C14436 FILLER_0_17_226/a_36_472# FILLER_0_17_218/a_484_472# 0.013277f
C14437 _112_ calibrate 0.024557f
C14438 FILLER_0_7_72/a_572_375# vss 0.006884f
C14439 output37/a_224_472# fanout65/a_36_113# 0.013171f
C14440 FILLER_0_11_124/a_124_375# _135_ 0.004831f
C14441 _098_ FILLER_0_15_235/a_124_375# 0.012702f
C14442 output17/a_224_472# net43 0.006661f
C14443 _413_/a_2560_156# net82 0.00101f
C14444 _129_ cal_count\[3\] 0.005967f
C14445 net52 trim_val\[4\] 0.21532f
C14446 _412_/a_36_151# net65 0.015454f
C14447 _086_ FILLER_0_6_177/a_484_472# 0.017841f
C14448 fanout78/a_36_113# net79 0.029496f
C14449 FILLER_0_20_177/a_36_472# _098_ 0.015061f
C14450 net55 _452_/a_836_156# 0.010887f
C14451 _411_/a_2560_156# _073_ 0.002649f
C14452 FILLER_0_5_164/a_36_472# _386_/a_848_380# 0.001177f
C14453 _052_ FILLER_0_18_61/a_36_472# 0.001508f
C14454 _129_ _059_ 0.005414f
C14455 FILLER_0_14_81/a_124_375# _095_ 0.009791f
C14456 net66 net47 0.238874f
C14457 _068_ _311_/a_1212_473# 0.002835f
C14458 fanout77/a_36_113# net18 0.060158f
C14459 _111_ _303_/a_244_68# 0.001153f
C14460 _092_ FILLER_0_17_218/a_572_375# 0.006125f
C14461 _021_ _093_ 0.049589f
C14462 _065_ fanout50/a_36_160# 0.022932f
C14463 net54 _436_/a_2248_156# 0.043158f
C14464 _067_ net47 0.0609f
C14465 _149_ _354_/a_49_472# 0.017453f
C14466 _424_/a_36_151# _012_ 0.005964f
C14467 _104_ output18/a_224_472# 0.08426f
C14468 trim_mask\[1\] FILLER_0_6_47/a_1828_472# 0.007542f
C14469 _033_ _444_/a_36_151# 0.014843f
C14470 FILLER_0_18_177/a_36_472# FILLER_0_19_171/a_572_375# 0.001684f
C14471 _118_ _315_/a_244_497# 0.003007f
C14472 FILLER_0_21_125/a_36_472# _436_/a_36_151# 0.001695f
C14473 output36/a_224_472# net19 0.106928f
C14474 FILLER_0_8_2/a_124_375# vdd 0.016103f
C14475 _432_/a_2665_112# _136_ 0.002691f
C14476 FILLER_0_15_116/a_484_472# _136_ 0.002712f
C14477 net82 fanout52/a_36_160# 0.026154f
C14478 FILLER_0_9_28/a_36_472# vdd 0.086674f
C14479 net19 net30 0.311153f
C14480 FILLER_0_13_228/a_36_472# vdd 0.085375f
C14481 FILLER_0_13_228/a_124_375# vss 0.007465f
C14482 _091_ FILLER_0_19_171/a_484_472# 0.013944f
C14483 FILLER_0_19_47/a_124_375# vdd 0.025971f
C14484 _088_ _073_ 0.001254f
C14485 _432_/a_1308_423# _137_ 0.002078f
C14486 _286_/a_224_472# _005_ 0.001254f
C14487 net18 _416_/a_1308_423# 0.021956f
C14488 _091_ FILLER_0_18_171/a_124_375# 0.034351f
C14489 net75 _425_/a_1308_423# 0.034219f
C14490 _301_/a_36_472# FILLER_0_22_86/a_36_472# 0.010679f
C14491 mask\[8\] FILLER_0_22_86/a_124_375# 0.014263f
C14492 FILLER_0_13_65/a_36_472# _043_ 0.013651f
C14493 FILLER_0_15_10/a_36_472# vdd 0.086171f
C14494 FILLER_0_15_10/a_124_375# vss 0.002173f
C14495 _308_/a_848_380# _070_ 0.033275f
C14496 FILLER_0_4_144/a_36_472# vss 0.008308f
C14497 FILLER_0_4_144/a_484_472# vdd 0.004027f
C14498 _178_ FILLER_0_15_10/a_124_375# 0.002355f
C14499 _091_ fanout56/a_36_113# 0.001254f
C14500 net20 FILLER_0_13_228/a_36_472# 0.020589f
C14501 output19/a_224_472# ctlp[2] 0.04607f
C14502 net35 FILLER_0_22_128/a_484_472# 0.004578f
C14503 net17 _452_/a_836_156# 0.002817f
C14504 _053_ net68 0.239882f
C14505 _048_ _047_ 0.007849f
C14506 net35 _049_ 0.022439f
C14507 FILLER_0_10_78/a_124_375# cal_count\[3\] 0.012197f
C14508 FILLER_0_18_177/a_2812_375# net22 0.010501f
C14509 _185_ cal_count\[2\] 0.205002f
C14510 FILLER_0_4_197/a_124_375# net76 0.00811f
C14511 FILLER_0_18_2/a_1468_375# net55 0.007169f
C14512 _281_/a_672_472# _097_ 0.002131f
C14513 _114_ _135_ 0.018715f
C14514 _413_/a_36_151# vss 0.003285f
C14515 net60 _419_/a_2248_156# 0.047724f
C14516 net61 _419_/a_2560_156# 0.008214f
C14517 net54 FILLER_0_22_128/a_1020_375# 0.010068f
C14518 FILLER_0_17_104/a_1380_472# vdd 0.010877f
C14519 _444_/a_796_472# net40 0.005776f
C14520 _431_/a_2665_112# FILLER_0_16_154/a_36_472# 0.007491f
C14521 net4 _081_ 0.02226f
C14522 _070_ FILLER_0_9_105/a_572_375# 0.017191f
C14523 _013_ FILLER_0_18_37/a_1380_472# 0.01384f
C14524 mask\[5\] output18/a_224_472# 0.00133f
C14525 _432_/a_448_472# FILLER_0_19_171/a_572_375# 0.00184f
C14526 FILLER_0_17_72/a_2812_375# _136_ 0.017702f
C14527 FILLER_0_7_162/a_36_472# FILLER_0_8_156/a_572_375# 0.001543f
C14528 FILLER_0_16_89/a_484_472# _451_/a_448_472# 0.059367f
C14529 net10 _411_/a_2248_156# 0.002419f
C14530 _013_ FILLER_0_17_56/a_124_375# 0.001047f
C14531 net34 result[8] 0.076645f
C14532 FILLER_0_7_72/a_1020_375# vss 0.004851f
C14533 net74 _067_ 0.674895f
C14534 _083_ vdd 0.157549f
C14535 _078_ vss 0.367953f
C14536 mask\[4\] FILLER_0_19_187/a_484_472# 0.004669f
C14537 output31/a_224_472# FILLER_0_16_255/a_124_375# 0.001274f
C14538 FILLER_0_7_146/a_124_375# vdd 0.034288f
C14539 net52 trim_val\[3\] 0.082691f
C14540 _073_ cal_itt\[0\] 0.211566f
C14541 net24 _436_/a_36_151# 0.075327f
C14542 net55 FILLER_0_18_53/a_484_472# 0.012319f
C14543 _415_/a_448_472# net19 0.03569f
C14544 net65 net4 0.614946f
C14545 FILLER_0_2_111/a_36_472# _157_ 0.104961f
C14546 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_124_375# 0.026339f
C14547 _176_ _390_/a_36_68# 0.005007f
C14548 FILLER_0_16_89/a_1468_375# _131_ 0.016581f
C14549 net20 _083_ 0.230786f
C14550 FILLER_0_10_78/a_1380_472# FILLER_0_10_94/a_36_472# 0.013277f
C14551 _115_ FILLER_0_10_94/a_572_375# 0.00887f
C14552 FILLER_0_16_37/a_124_375# FILLER_0_17_38/a_36_472# 0.001723f
C14553 FILLER_0_12_136/a_932_472# _069_ 0.002161f
C14554 FILLER_0_12_136/a_36_472# _126_ 0.014981f
C14555 trim_val\[3\] net49 0.009336f
C14556 _065_ net14 0.005438f
C14557 _075_ _077_ 0.004518f
C14558 FILLER_0_20_193/a_36_472# FILLER_0_20_177/a_1380_472# 0.013276f
C14559 FILLER_0_18_2/a_1468_375# net17 0.004803f
C14560 trim_mask\[4\] _066_ 0.396509f
C14561 net1 _082_ 0.033169f
C14562 FILLER_0_8_107/a_36_472# _219_/a_36_160# 0.002767f
C14563 trim_val\[2\] net40 0.06019f
C14564 _415_/a_2665_112# FILLER_0_9_290/a_36_472# 0.007376f
C14565 _053_ net67 0.672744f
C14566 net82 net1 0.029512f
C14567 FILLER_0_20_193/a_484_472# vss 0.002439f
C14568 net47 _066_ 0.096823f
C14569 output33/a_224_472# vdd -0.031734f
C14570 _077_ FILLER_0_10_94/a_36_472# 0.001114f
C14571 FILLER_0_17_72/a_2276_472# _131_ 0.004125f
C14572 _065_ _164_ 0.006953f
C14573 _130_ vdd 0.046379f
C14574 trim[0] trim[3] 0.012429f
C14575 trim_val\[0\] FILLER_0_6_47/a_572_375# 0.03235f
C14576 _420_/a_1000_472# _009_ 0.019219f
C14577 _173_ _067_ 0.011854f
C14578 FILLER_0_11_101/a_124_375# _058_ 0.002209f
C14579 _056_ cal_count\[3\] 0.186969f
C14580 _158_ _154_ 0.008872f
C14581 _369_/a_36_68# _153_ 0.008048f
C14582 net34 FILLER_0_22_177/a_1468_375# 0.006974f
C14583 FILLER_0_15_116/a_484_472# net53 0.002804f
C14584 _413_/a_36_151# FILLER_0_3_172/a_3260_375# 0.059049f
C14585 _070_ _125_ 0.125523f
C14586 _076_ _058_ 0.912225f
C14587 net68 FILLER_0_8_37/a_572_375# 0.011704f
C14588 _438_/a_796_472# net71 0.00514f
C14589 cal_count\[3\] _453_/a_36_151# 0.023915f
C14590 trim_mask\[4\] net23 0.180803f
C14591 FILLER_0_18_177/a_2276_472# FILLER_0_19_195/a_124_375# 0.001684f
C14592 FILLER_0_15_72/a_124_375# FILLER_0_15_59/a_572_375# 0.003228f
C14593 _233_/a_36_160# _445_/a_2248_156# 0.00136f
C14594 FILLER_0_5_54/a_932_472# vss 0.003426f
C14595 FILLER_0_5_54/a_1380_472# vdd 0.008983f
C14596 net23 net47 0.090948f
C14597 _430_/a_2560_156# vss 0.002924f
C14598 _077_ calibrate 0.055446f
C14599 FILLER_0_17_72/a_36_472# net36 0.001121f
C14600 cal_count\[3\] FILLER_0_11_135/a_124_375# 0.004365f
C14601 result[4] net79 0.048452f
C14602 mask\[9\] _438_/a_448_472# 0.046823f
C14603 FILLER_0_5_164/a_124_375# vdd 0.00419f
C14604 output13/a_224_472# net23 0.00255f
C14605 _026_ FILLER_0_20_87/a_124_375# 0.031902f
C14606 _431_/a_2665_112# FILLER_0_18_139/a_1380_472# 0.001008f
C14607 _251_/a_906_472# _070_ 0.002124f
C14608 result[5] fanout78/a_36_113# 0.018989f
C14609 _033_ _054_ 0.003394f
C14610 net15 FILLER_0_6_47/a_2276_472# 0.049487f
C14611 _182_ vdd 0.161134f
C14612 FILLER_0_10_28/a_36_472# net17 0.012954f
C14613 net25 _012_ 0.001747f
C14614 cal_itt\[3\] _055_ 0.007428f
C14615 _141_ _346_/a_665_69# 0.002048f
C14616 FILLER_0_6_239/a_124_375# _317_/a_36_113# 0.002437f
C14617 FILLER_0_18_177/a_2812_375# vdd 0.003766f
C14618 _449_/a_2665_112# _067_ 0.03661f
C14619 mask\[7\] _024_ 0.122185f
C14620 output8/a_224_472# FILLER_0_3_221/a_124_375# 0.03228f
C14621 _077_ net21 0.032627f
C14622 _450_/a_836_156# _039_ 0.019042f
C14623 FILLER_0_11_101/a_572_375# cal_count\[3\] 0.002017f
C14624 net18 _419_/a_36_151# 0.021491f
C14625 net69 _384_/a_224_472# 0.002407f
C14626 net16 FILLER_0_18_37/a_1468_375# 0.002269f
C14627 FILLER_0_15_282/a_36_472# _006_ 0.003055f
C14628 net41 net47 0.19549f
C14629 net69 _441_/a_448_472# 0.028545f
C14630 _432_/a_2248_156# FILLER_0_18_177/a_1828_472# 0.035805f
C14631 result[7] _103_ 0.298427f
C14632 _432_/a_796_472# _098_ 0.038458f
C14633 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_572_375# 0.001597f
C14634 _068_ _059_ 0.255081f
C14635 state\[1\] _225_/a_36_160# 0.0535f
C14636 FILLER_0_18_171/a_36_472# vss 0.0032f
C14637 _425_/a_36_151# vdd 0.078723f
C14638 net81 cal_itt\[0\] 0.001048f
C14639 FILLER_0_5_172/a_36_472# net47 0.0015f
C14640 net17 FILLER_0_20_15/a_36_472# 0.004375f
C14641 _163_ FILLER_0_5_148/a_484_472# 0.002734f
C14642 _187_ net51 0.04894f
C14643 mask\[7\] FILLER_0_22_128/a_2812_375# 0.001476f
C14644 _033_ vss 0.019158f
C14645 net34 output18/a_224_472# 0.17524f
C14646 FILLER_0_17_226/a_124_375# _093_ 0.001604f
C14647 net4 _090_ 0.06324f
C14648 _255_/a_224_552# cal_itt\[3\] 0.003266f
C14649 FILLER_0_24_290/a_124_375# vss 0.034103f
C14650 FILLER_0_24_290/a_36_472# vdd 0.089567f
C14651 net53 _427_/a_448_472# 0.047356f
C14652 output14/a_224_472# vdd 0.054725f
C14653 calibrate _120_ 0.001106f
C14654 net31 FILLER_0_16_255/a_36_472# 0.003056f
C14655 _103_ _198_/a_67_603# 0.005362f
C14656 state\[1\] FILLER_0_12_196/a_36_472# 0.030132f
C14657 _105_ _293_/a_36_472# 0.004667f
C14658 _448_/a_448_472# net22 0.085004f
C14659 net38 FILLER_0_12_2/a_484_472# 0.002706f
C14660 FILLER_0_17_200/a_484_472# net22 0.020589f
C14661 _428_/a_2665_112# _043_ 0.021483f
C14662 mask\[4\] _092_ 0.072581f
C14663 fanout74/a_36_113# vss 0.048756f
C14664 net60 output18/a_224_472# 0.001518f
C14665 _008_ mask\[3\] 0.799138f
C14666 net50 _439_/a_36_151# 0.009774f
C14667 net52 _439_/a_1308_423# 0.033366f
C14668 _274_/a_36_68# FILLER_0_12_236/a_484_472# 0.001237f
C14669 _445_/a_2248_156# net49 0.029744f
C14670 _137_ vdd 0.945976f
C14671 fanout51/a_36_113# cal_count\[3\] 0.054567f
C14672 net74 net23 0.0064f
C14673 FILLER_0_4_185/a_36_472# net76 0.023698f
C14674 FILLER_0_16_57/a_932_472# FILLER_0_15_59/a_572_375# 0.001543f
C14675 _028_ _053_ 0.891578f
C14676 _250_/a_36_68# vss 0.005108f
C14677 _128_ _060_ 0.022833f
C14678 net79 net64 0.049663f
C14679 _013_ FILLER_0_18_53/a_124_375# 0.015996f
C14680 _180_ vss 0.106022f
C14681 mask\[3\] _141_ 0.361692f
C14682 _028_ FILLER_0_6_47/a_2812_375# 0.023189f
C14683 _178_ _180_ 0.004668f
C14684 output26/a_224_472# net26 0.047008f
C14685 _443_/a_2560_156# _170_ 0.00758f
C14686 _443_/a_2248_156# _037_ 0.005717f
C14687 net15 _440_/a_1204_472# 0.01349f
C14688 state\[2\] FILLER_0_13_142/a_932_472# 0.004118f
C14689 net16 _181_ 0.48682f
C14690 _114_ _069_ 0.029875f
C14691 _015_ FILLER_0_8_247/a_1020_375# 0.006994f
C14692 _043_ cal_count\[0\] 0.019077f
C14693 _421_/a_448_472# net77 0.003958f
C14694 FILLER_0_3_78/a_36_472# vdd 0.082597f
C14695 FILLER_0_3_78/a_572_375# vss 0.04008f
C14696 FILLER_0_2_127/a_36_472# vdd 0.08468f
C14697 FILLER_0_2_127/a_124_375# vss 0.008566f
C14698 _394_/a_728_93# _095_ 0.035417f
C14699 _132_ FILLER_0_14_107/a_572_375# 0.007439f
C14700 FILLER_0_4_152/a_36_472# FILLER_0_4_144/a_484_472# 0.013276f
C14701 FILLER_0_24_274/a_1380_472# vss 0.005744f
C14702 _308_/a_124_24# FILLER_0_9_72/a_1468_375# 0.007188f
C14703 _077_ _256_/a_36_68# 0.027906f
C14704 net63 FILLER_0_18_177/a_36_472# 0.015187f
C14705 FILLER_0_17_104/a_1468_375# FILLER_0_16_115/a_124_375# 0.026339f
C14706 en_co_clk _389_/a_36_148# 0.001249f
C14707 FILLER_0_22_128/a_484_472# vdd 0.002467f
C14708 _297_/a_36_472# _295_/a_36_472# 0.004259f
C14709 FILLER_0_22_128/a_36_472# vss 0.001309f
C14710 _449_/a_2248_156# fanout55/a_36_160# 0.027388f
C14711 _186_ _407_/a_244_68# 0.001153f
C14712 _049_ vdd 0.199608f
C14713 _086_ _058_ 0.054155f
C14714 net27 _426_/a_1308_423# 0.00384f
C14715 _098_ _043_ 0.032706f
C14716 _414_/a_36_151# FILLER_0_6_177/a_484_472# 0.006095f
C14717 net56 FILLER_0_18_139/a_572_375# 0.005919f
C14718 trimb[0] net44 0.00246f
C14719 output27/a_224_472# FILLER_0_8_263/a_124_375# 0.011584f
C14720 output35/a_224_472# _098_ 0.003653f
C14721 _441_/a_2248_156# FILLER_0_3_78/a_572_375# 0.001068f
C14722 _131_ _134_ 0.887647f
C14723 _088_ FILLER_0_3_172/a_2276_472# 0.024532f
C14724 _304_/a_224_472# vss 0.001746f
C14725 _053_ FILLER_0_6_47/a_1916_375# 0.008103f
C14726 _425_/a_1308_423# net19 0.058462f
C14727 output46/a_224_472# net17 0.082914f
C14728 output21/a_224_472# net33 0.001166f
C14729 FILLER_0_4_177/a_124_375# net37 0.00459f
C14730 FILLER_0_16_241/a_124_375# mask\[2\] 0.027201f
C14731 net75 net59 0.06935f
C14732 net82 FILLER_0_3_172/a_2364_375# 0.010439f
C14733 output35/a_224_472# _205_/a_36_160# 0.002043f
C14734 _411_/a_36_151# FILLER_0_0_232/a_36_472# 0.001723f
C14735 _093_ FILLER_0_18_107/a_2812_375# 0.00626f
C14736 _413_/a_2560_156# net21 0.002416f
C14737 net54 net36 0.005827f
C14738 _446_/a_448_472# vdd 0.006805f
C14739 _127_ _176_ 0.319517f
C14740 _128_ _116_ 0.069335f
C14741 net55 cal_count\[2\] 0.022989f
C14742 net79 _006_ 0.050445f
C14743 FILLER_0_6_177/a_484_472# _163_ 0.002256f
C14744 output48/a_224_472# _112_ 0.027383f
C14745 fanout80/a_36_113# _138_ 0.002489f
C14746 _322_/a_848_380# _126_ 0.002519f
C14747 _449_/a_36_151# FILLER_0_12_50/a_36_472# 0.003462f
C14748 net21 mask\[6\] 0.634881f
C14749 FILLER_0_17_282/a_36_472# vss 0.007765f
C14750 _152_ _059_ 0.038141f
C14751 output19/a_224_472# mask\[7\] 0.001181f
C14752 _316_/a_692_472# _122_ 0.002929f
C14753 _316_/a_1152_472# calibrate 0.001604f
C14754 FILLER_0_15_116/a_124_375# vdd 0.012886f
C14755 _026_ _098_ 0.197713f
C14756 _432_/a_448_472# net63 0.002757f
C14757 FILLER_0_9_142/a_36_472# _118_ 0.01533f
C14758 _076_ _226_/a_860_68# 0.001752f
C14759 _095_ FILLER_0_15_10/a_124_375# 0.023187f
C14760 net73 FILLER_0_17_142/a_484_472# 0.001122f
C14761 _412_/a_1000_472# vdd 0.002008f
C14762 _448_/a_448_472# vdd 0.02042f
C14763 FILLER_0_17_200/a_484_472# vdd 0.008335f
C14764 result[5] result[4] 0.090472f
C14765 FILLER_0_3_142/a_124_375# net23 0.25251f
C14766 FILLER_0_23_60/a_36_472# vss 0.006794f
C14767 net55 FILLER_0_19_28/a_484_472# 0.001426f
C14768 FILLER_0_3_142/a_36_472# trim_mask\[4\] 0.008297f
C14769 net15 net36 0.265646f
C14770 _440_/a_2665_112# FILLER_0_4_91/a_36_472# 0.007491f
C14771 net75 _122_ 0.052177f
C14772 _128_ _118_ 0.58787f
C14773 _127_ _124_ 0.035569f
C14774 _104_ net18 0.039321f
C14775 FILLER_0_18_100/a_36_472# vss 0.002412f
C14776 FILLER_0_7_59/a_124_375# net68 0.019553f
C14777 _379_/a_244_68# _160_ 0.001202f
C14778 FILLER_0_5_54/a_124_375# net47 0.012889f
C14779 _414_/a_2665_112# cal_itt\[3\] 0.02392f
C14780 _041_ FILLER_0_18_37/a_1468_375# 0.001032f
C14781 net55 _423_/a_2665_112# 0.002379f
C14782 net26 FILLER_0_21_28/a_1380_472# 0.035291f
C14783 net45 net40 0.029947f
C14784 _433_/a_1000_472# _145_ 0.004227f
C14785 FILLER_0_14_99/a_36_472# net14 0.036527f
C14786 cal_count\[2\] net17 0.074204f
C14787 net75 FILLER_0_10_256/a_36_472# 0.010024f
C14788 _376_/a_36_160# FILLER_0_6_90/a_124_375# 0.005705f
C14789 FILLER_0_14_263/a_124_375# vss 0.007923f
C14790 FILLER_0_14_263/a_36_472# vdd 0.02759f
C14791 _043_ FILLER_0_15_180/a_124_375# 0.003099f
C14792 _010_ vss 0.064717f
C14793 net57 trim_mask\[4\] 0.259381f
C14794 net75 net64 0.037337f
C14795 _072_ _085_ 0.408915f
C14796 _386_/a_848_380# _169_ 0.001355f
C14797 _386_/a_124_24# _163_ 0.001234f
C14798 _236_/a_36_160# trim[1] 0.003604f
C14799 net23 FILLER_0_19_155/a_36_472# 0.019429f
C14800 FILLER_0_17_72/a_1020_375# vss 0.005441f
C14801 FILLER_0_17_72/a_1468_375# vdd 0.003316f
C14802 net57 net47 0.279638f
C14803 _089_ _122_ 0.006163f
C14804 fanout49/a_36_160# _156_ 0.002871f
C14805 net73 FILLER_0_18_107/a_2276_472# 0.016723f
C14806 mask\[0\] _335_/a_665_69# 0.001711f
C14807 FILLER_0_4_107/a_1468_375# vdd 0.023541f
C14808 _273_/a_36_68# FILLER_0_10_214/a_36_472# 0.003036f
C14809 net58 net1 0.626432f
C14810 net4 FILLER_0_7_233/a_36_472# 0.036721f
C14811 FILLER_0_9_270/a_36_472# vdd 0.008742f
C14812 FILLER_0_9_270/a_572_375# vss 0.017196f
C14813 FILLER_0_5_109/a_124_375# _151_ 0.003377f
C14814 _032_ _370_/a_124_24# 0.007035f
C14815 FILLER_0_21_125/a_484_472# _098_ 0.002964f
C14816 net38 FILLER_0_20_2/a_484_472# 0.006727f
C14817 net17 _450_/a_448_472# 0.017832f
C14818 result[9] _418_/a_2665_112# 0.053489f
C14819 FILLER_0_16_241/a_36_472# _099_ 0.158391f
C14820 net52 FILLER_0_2_111/a_572_375# 0.00245f
C14821 output19/a_224_472# _422_/a_2248_156# 0.011418f
C14822 _063_ _160_ 0.091185f
C14823 mask\[4\] FILLER_0_19_195/a_36_472# 0.004669f
C14824 _004_ FILLER_0_10_256/a_36_472# 0.00402f
C14825 FILLER_0_21_142/a_484_472# vss 0.034607f
C14826 net52 _440_/a_448_472# 0.067294f
C14827 _004_ net64 0.001495f
C14828 net60 _421_/a_1000_472# 0.035511f
C14829 mask\[3\] FILLER_0_18_177/a_124_375# 0.002924f
C14830 net55 _043_ 0.053191f
C14831 fanout73/a_36_113# net74 0.04136f
C14832 input5/a_36_113# net59 0.257143f
C14833 net81 net36 0.030215f
C14834 _401_/a_36_68# _180_ 0.051459f
C14835 _179_ cal_count\[1\] 0.088667f
C14836 _091_ FILLER_0_16_154/a_1468_375# 0.003056f
C14837 net50 FILLER_0_8_37/a_36_472# 0.059367f
C14838 FILLER_0_23_282/a_36_472# vss 0.003317f
C14839 _141_ FILLER_0_19_155/a_572_375# 0.033271f
C14840 net81 _429_/a_1204_472# 0.005046f
C14841 FILLER_0_11_142/a_124_375# _120_ 0.036088f
C14842 net10 FILLER_0_1_212/a_124_375# 0.002314f
C14843 _198_/a_67_603# mask\[2\] 0.005143f
C14844 FILLER_0_3_142/a_36_472# net74 0.001098f
C14845 fanout64/a_36_160# fanout65/a_36_113# 0.001627f
C14846 mask\[7\] mask\[6\] 0.227476f
C14847 FILLER_0_13_142/a_36_472# vss 0.005768f
C14848 net49 _440_/a_448_472# 0.049861f
C14849 mask\[8\] mask\[7\] 0.021731f
C14850 net82 net76 0.061682f
C14851 _091_ _055_ 0.003332f
C14852 net52 FILLER_0_5_72/a_1380_472# 0.001523f
C14853 FILLER_0_7_59/a_124_375# net67 0.036499f
C14854 _061_ _062_ 0.344031f
C14855 FILLER_0_19_142/a_124_375# vss 0.032026f
C14856 FILLER_0_19_142/a_36_472# vdd 0.107105f
C14857 _431_/a_2665_112# net73 0.001495f
C14858 _040_ vdd 0.065702f
C14859 net74 _442_/a_1308_423# 0.001618f
C14860 FILLER_0_11_142/a_36_472# FILLER_0_13_142/a_124_375# 0.0027f
C14861 _062_ _311_/a_66_473# 0.027039f
C14862 _447_/a_448_472# vdd 0.014537f
C14863 _447_/a_36_151# vss 0.001541f
C14864 _250_/a_36_68# _071_ 0.199512f
C14865 cal_count\[3\] _113_ 0.093684f
C14866 _413_/a_2248_156# net65 0.036792f
C14867 FILLER_0_5_72/a_1380_472# net49 0.002057f
C14868 ctln[2] output10/a_224_472# 0.024524f
C14869 net57 net74 2.360287f
C14870 net50 _160_ 0.048787f
C14871 FILLER_0_7_72/a_2276_472# net50 0.030391f
C14872 FILLER_0_24_96/a_36_472# vss 0.003218f
C14873 net81 FILLER_0_10_247/a_36_472# 0.015109f
C14874 _137_ FILLER_0_16_154/a_572_375# 0.010132f
C14875 comp FILLER_0_15_2/a_36_472# 0.001941f
C14876 net17 _043_ 0.571818f
C14877 net54 _433_/a_1308_423# 0.004372f
C14878 fanout54/a_36_160# _433_/a_2248_156# 0.012122f
C14879 net29 _196_/a_36_160# 0.073294f
C14880 FILLER_0_5_72/a_124_375# _440_/a_36_151# 0.059049f
C14881 _105_ output19/a_224_472# 0.107668f
C14882 FILLER_0_12_28/a_36_472# _450_/a_3129_107# 0.009814f
C14883 mask\[4\] FILLER_0_18_177/a_2276_472# 0.016876f
C14884 _450_/a_3129_107# net40 0.034729f
C14885 _447_/a_2248_156# _441_/a_36_151# 0.035837f
C14886 net58 result[0] 0.443436f
C14887 net49 _034_ 0.031359f
C14888 result[7] _420_/a_2248_156# 0.034866f
C14889 _093_ FILLER_0_16_115/a_36_472# 0.001526f
C14890 FILLER_0_8_107/a_36_472# _058_ 0.015262f
C14891 net31 output33/a_224_472# 0.005087f
C14892 net22 net12 0.032084f
C14893 net81 FILLER_0_15_228/a_36_472# 0.003953f
C14894 cal_itt\[2\] _083_ 0.10423f
C14895 _053_ FILLER_0_7_72/a_484_472# 0.00887f
C14896 _239_/a_36_160# net40 0.010925f
C14897 vdd FILLER_0_10_94/a_572_375# 0.02784f
C14898 _444_/a_36_151# _054_ 0.011342f
C14899 output10/a_224_472# ctln[1] 0.083631f
C14900 output22/a_224_472# net80 0.00955f
C14901 net82 FILLER_0_2_177/a_124_375# 0.003837f
C14902 _072_ _062_ 0.025795f
C14903 _430_/a_36_151# mask\[2\] 0.016265f
C14904 mask\[5\] _048_ 0.062788f
C14905 _320_/a_1120_472# _090_ 0.001215f
C14906 _140_ FILLER_0_21_150/a_36_472# 0.015502f
C14907 FILLER_0_24_130/a_36_472# _050_ 0.008605f
C14908 net56 FILLER_0_17_142/a_484_472# 0.008895f
C14909 net81 en 0.071123f
C14910 result[0] calibrate 0.00287f
C14911 net68 net17 0.601273f
C14912 result[5] _103_ 0.425479f
C14913 output32/a_224_472# _418_/a_2665_112# 0.011048f
C14914 _363_/a_692_472# _028_ 0.001416f
C14915 result[6] FILLER_0_21_286/a_484_472# 0.011149f
C14916 _025_ _436_/a_1308_423# 0.006243f
C14917 _091_ FILLER_0_12_220/a_572_375# 0.003075f
C14918 net68 trim_val\[1\] 0.006974f
C14919 state\[0\] _323_/a_36_113# 0.016796f
C14920 output34/a_224_472# vdd 0.094191f
C14921 output44/a_224_472# net38 0.106923f
C14922 _091_ _432_/a_1204_472# 0.00563f
C14923 _444_/a_36_151# vss 0.003795f
C14924 _444_/a_448_472# vdd 0.03285f
C14925 FILLER_0_10_78/a_1020_375# net52 0.001158f
C14926 FILLER_0_3_172/a_1916_375# net59 0.001221f
C14927 _448_/a_2248_156# _443_/a_2248_156# 0.006556f
C14928 FILLER_0_7_72/a_572_375# _053_ 0.014569f
C14929 FILLER_0_8_24/a_124_375# vdd 0.01166f
C14930 output10/a_224_472# FILLER_0_0_266/a_36_472# 0.023414f
C14931 fanout59/a_36_160# vdd 0.02169f
C14932 _453_/a_1204_472# _042_ 0.002408f
C14933 _120_ _171_ 0.414533f
C14934 _136_ _172_ 0.024344f
C14935 _095_ _180_ 0.013383f
C14936 result[8] FILLER_0_24_274/a_484_472# 0.005458f
C14937 net20 output34/a_224_472# 0.023142f
C14938 output31/a_224_472# FILLER_0_17_282/a_36_472# 0.008834f
C14939 result[4] net19 0.015095f
C14940 net19 net59 0.0206f
C14941 FILLER_0_7_72/a_932_472# net50 0.074005f
C14942 result[7] _419_/a_2665_112# 0.002471f
C14943 FILLER_0_10_78/a_124_375# net52 0.008557f
C14944 _438_/a_36_151# net14 0.008367f
C14945 FILLER_0_2_93/a_572_375# vdd 0.022073f
C14946 _080_ vss 0.012982f
C14947 FILLER_0_19_171/a_484_472# vdd 0.009225f
C14948 FILLER_0_19_171/a_36_472# vss 0.001338f
C14949 ctln[7] FILLER_0_0_130/a_124_375# 0.002726f
C14950 trim[4] FILLER_0_8_2/a_124_375# 0.028454f
C14951 FILLER_0_18_171/a_124_375# vdd 0.021417f
C14952 mask\[8\] _437_/a_448_472# 0.008198f
C14953 net57 FILLER_0_3_142/a_124_375# 0.003738f
C14954 net23 FILLER_0_5_148/a_124_375# 0.01836f
C14955 net60 net18 0.949607f
C14956 _306_/a_36_68# _055_ 0.006686f
C14957 _452_/a_3129_107# vss 0.00145f
C14958 _452_/a_2225_156# vdd 0.005612f
C14959 fanout56/a_36_113# vdd 0.078814f
C14960 FILLER_0_6_239/a_124_375# _122_ 0.01772f
C14961 FILLER_0_7_195/a_36_472# vss 0.002568f
C14962 net47 FILLER_0_5_148/a_572_375# 0.062581f
C14963 net16 _446_/a_2248_156# 0.010032f
C14964 _105_ mask\[6\] 0.029716f
C14965 FILLER_0_22_86/a_124_375# _026_ 0.001024f
C14966 _253_/a_36_68# cal_itt\[0\] 0.001495f
C14967 _359_/a_1044_488# _129_ 0.001111f
C14968 net67 net17 0.04175f
C14969 FILLER_0_23_44/a_1020_375# vdd -0.014642f
C14970 net32 result[6] 0.048987f
C14971 net15 _441_/a_36_151# 0.01821f
C14972 net12 vdd 0.082923f
C14973 _165_ trim_val\[0\] 0.164683f
C14974 _018_ vss 0.022336f
C14975 _440_/a_1204_472# net47 0.006257f
C14976 _412_/a_36_151# net48 0.001091f
C14977 _418_/a_36_151# vdd 0.155643f
C14978 FILLER_0_14_107/a_484_472# vdd 0.030114f
C14979 FILLER_0_14_107/a_36_472# vss 0.003706f
C14980 _431_/a_2665_112# net56 0.048214f
C14981 _412_/a_2665_112# fanout58/a_36_160# 0.001221f
C14982 _136_ FILLER_0_16_115/a_36_472# 0.013477f
C14983 _448_/a_36_151# FILLER_0_2_177/a_36_472# 0.04556f
C14984 _114_ FILLER_0_12_136/a_932_472# 0.003953f
C14985 FILLER_0_3_172/a_2364_375# net21 0.004803f
C14986 FILLER_0_22_177/a_1020_375# net33 0.013731f
C14987 _433_/a_448_472# _022_ 0.074451f
C14988 _306_/a_36_68# _126_ 0.01893f
C14989 net36 _045_ 0.091033f
C14990 output21/a_224_472# net22 0.022576f
C14991 net15 FILLER_0_9_60/a_484_472# 0.020589f
C14992 _395_/a_1044_488# _071_ 0.001198f
C14993 _010_ _419_/a_1000_472# 0.001598f
C14994 FILLER_0_21_286/a_124_375# vdd 0.026138f
C14995 _445_/a_448_472# net17 0.038794f
C14996 net81 output27/a_224_472# 0.011872f
C14997 _086_ _134_ 0.020487f
C14998 net64 net19 0.029763f
C14999 _187_ _173_ 0.03421f
C15000 FILLER_0_17_200/a_484_472# _069_ 0.001396f
C15001 net63 net64 0.002181f
C15002 FILLER_0_7_72/a_1020_375# _053_ 0.014569f
C15003 _256_/a_2552_68# _072_ 0.001213f
C15004 net2 en 0.067828f
C15005 _053_ _078_ 0.137388f
C15006 net50 FILLER_0_7_59/a_572_375# 0.009554f
C15007 net33 _204_/a_67_603# 0.022193f
C15008 net63 FILLER_0_19_171/a_1380_472# 0.003014f
C15009 FILLER_0_18_2/a_2812_375# vdd 0.021655f
C15010 net54 FILLER_0_22_86/a_1380_472# 0.059367f
C15011 _136_ FILLER_0_16_154/a_932_472# 0.008185f
C15012 _334_/a_36_160# vdd 0.041716f
C15013 _088_ FILLER_0_3_221/a_484_472# 0.002245f
C15014 _395_/a_36_488# _055_ 0.002775f
C15015 net48 _316_/a_848_380# 0.026413f
C15016 FILLER_0_19_125/a_124_375# FILLER_0_18_107/a_2276_472# 0.001684f
C15017 _431_/a_36_151# FILLER_0_16_115/a_36_472# 0.004847f
C15018 net35 _051_ 0.019252f
C15019 mask\[5\] FILLER_0_18_177/a_484_472# 0.001063f
C15020 FILLER_0_14_81/a_124_375# net55 0.038949f
C15021 FILLER_0_16_89/a_932_472# _040_ 0.00702f
C15022 result[8] output19/a_224_472# 0.001465f
C15023 output35/a_224_472# ctlp[2] 0.001465f
C15024 output26/a_224_472# FILLER_0_23_60/a_36_472# 0.003292f
C15025 vss _433_/a_2560_156# 0.003477f
C15026 _079_ _088_ 0.012529f
C15027 net16 FILLER_0_6_37/a_36_472# 0.013074f
C15028 _074_ FILLER_0_6_231/a_124_375# 0.006087f
C15029 cal_count\[3\] FILLER_0_11_78/a_572_375# 0.010243f
C15030 _000_ net82 0.032846f
C15031 _005_ _044_ 0.50767f
C15032 ctlp[1] FILLER_0_24_274/a_572_375# 0.002408f
C15033 input1/a_36_113# net2 0.018839f
C15034 _091_ _432_/a_1000_472# 0.026097f
C15035 FILLER_0_3_172/a_36_472# net22 0.012287f
C15036 FILLER_0_5_109/a_572_375# net47 0.011047f
C15037 _094_ _418_/a_2665_112# 0.035668f
C15038 FILLER_0_12_136/a_572_375# _127_ 0.00116f
C15039 net5 vdd 0.516129f
C15040 _422_/a_1308_423# mask\[7\] 0.045368f
C15041 _411_/a_2248_156# vdd 0.006283f
C15042 fanout66/a_36_113# FILLER_0_3_54/a_36_472# 0.001645f
C15043 _086_ _267_/a_672_472# 0.004515f
C15044 _054_ vss 0.176655f
C15045 FILLER_0_9_60/a_484_472# net51 0.061362f
C15046 _003_ FILLER_0_5_181/a_124_375# 0.009929f
C15047 _076_ FILLER_0_6_231/a_124_375# 0.001382f
C15048 _070_ FILLER_0_6_231/a_36_472# 0.001096f
C15049 _058_ _117_ 0.003932f
C15050 _116_ _176_ 0.067051f
C15051 FILLER_0_5_128/a_36_472# _160_ 0.006214f
C15052 net19 _006_ 0.090449f
C15053 _321_/a_3126_472# _176_ 0.001932f
C15054 _069_ _395_/a_1492_488# 0.002565f
C15055 FILLER_0_16_37/a_124_375# cal_count\[2\] 0.008393f
C15056 _445_/a_2248_156# net40 0.004545f
C15057 net58 net76 0.700034f
C15058 net75 FILLER_0_8_247/a_572_375# 0.003962f
C15059 _446_/a_36_151# output41/a_224_472# 0.135198f
C15060 _412_/a_1308_423# net1 0.022273f
C15061 FILLER_0_15_235/a_484_472# vdd 0.006f
C15062 FILLER_0_15_235/a_36_472# vss 0.003138f
C15063 _408_/a_1336_472# _043_ 0.023648f
C15064 _408_/a_56_524# _190_/a_36_160# 0.004025f
C15065 _436_/a_2248_156# FILLER_0_22_128/a_572_375# 0.006739f
C15066 _436_/a_2665_112# FILLER_0_22_128/a_124_375# 0.004834f
C15067 FILLER_0_15_235/a_124_375# mask\[1\] 0.013103f
C15068 _093_ FILLER_0_19_155/a_124_375# 0.001864f
C15069 _053_ FILLER_0_5_54/a_932_472# 0.001578f
C15070 FILLER_0_9_105/a_484_472# vss 0.004412f
C15071 _178_ _278_/a_36_160# 0.269109f
C15072 FILLER_0_13_142/a_932_472# _043_ 0.011974f
C15073 FILLER_0_20_177/a_1380_472# vdd 0.009871f
C15074 FILLER_0_20_177/a_932_472# vss 0.001272f
C15075 net81 _425_/a_2560_156# 0.022037f
C15076 _103_ net19 0.047895f
C15077 output24/a_224_472# vss 0.004078f
C15078 FILLER_0_1_266/a_124_375# net19 0.007016f
C15079 FILLER_0_5_54/a_572_375# FILLER_0_6_47/a_1380_472# 0.001597f
C15080 ctlp[3] _422_/a_2665_112# 0.001024f
C15081 _012_ net36 0.053654f
C15082 net44 vdd 0.897202f
C15083 FILLER_0_16_57/a_572_375# FILLER_0_17_56/a_572_375# 0.026339f
C15084 FILLER_0_7_72/a_1916_375# _376_/a_36_160# 0.001925f
C15085 valid en 0.026142f
C15086 net48 net4 0.099614f
C15087 _178_ vss 0.150839f
C15088 _408_/a_728_93# _186_ 0.003815f
C15089 net36 FILLER_0_15_212/a_36_472# 0.005396f
C15090 output47/a_224_472# net40 0.002339f
C15091 net52 fanout51/a_36_113# 0.036773f
C15092 _095_ FILLER_0_13_142/a_36_472# 0.001782f
C15093 fanout66/a_36_113# _164_ 0.010496f
C15094 FILLER_0_17_56/a_572_375# _183_ 0.002605f
C15095 _429_/a_2248_156# FILLER_0_15_212/a_1468_375# 0.001068f
C15096 _176_ _118_ 0.392531f
C15097 _114_ _428_/a_2248_156# 0.004516f
C15098 FILLER_0_20_98/a_36_472# net14 0.024154f
C15099 FILLER_0_20_15/a_1380_472# vdd 0.007068f
C15100 cal_count\[3\] _042_ 0.001716f
C15101 _079_ cal_itt\[0\] 0.018495f
C15102 _008_ result[9] 0.048497f
C15103 output21/a_224_472# vdd 0.028725f
C15104 FILLER_0_18_107/a_1468_375# vdd 0.004726f
C15105 _098_ FILLER_0_21_150/a_124_375# 0.006526f
C15106 FILLER_0_4_107/a_36_472# _156_ 0.005297f
C15107 _289_/a_36_472# mask\[2\] 0.006392f
C15108 _321_/a_3126_472# _124_ 0.001072f
C15109 _076_ FILLER_0_8_239/a_36_472# 0.029514f
C15110 FILLER_0_12_50/a_124_375# cal_count\[0\] 0.002359f
C15111 _422_/a_1204_472# vdd 0.001062f
C15112 _106_ FILLER_0_17_218/a_484_472# 0.012952f
C15113 FILLER_0_18_139/a_572_375# _145_ 0.00346f
C15114 net79 FILLER_0_12_220/a_1468_375# 0.012754f
C15115 _441_/a_2665_112# vdd 0.012404f
C15116 _441_/a_2248_156# vss 0.005663f
C15117 net76 net21 0.041873f
C15118 FILLER_0_4_177/a_36_472# _074_ 0.002603f
C15119 _074_ _375_/a_692_497# 0.004556f
C15120 net55 _424_/a_2248_156# 0.057967f
C15121 output48/a_224_472# net1 0.006536f
C15122 FILLER_0_7_72/a_36_472# vss 0.033878f
C15123 trim_val\[4\] _386_/a_848_380# 0.007605f
C15124 FILLER_0_9_223/a_124_375# _068_ 0.010485f
C15125 _412_/a_1204_472# net58 0.018724f
C15126 FILLER_0_5_117/a_36_472# _153_ 0.028773f
C15127 _447_/a_1308_423# net68 0.006686f
C15128 _447_/a_36_151# _036_ 0.007244f
C15129 net52 net69 0.372114f
C15130 FILLER_0_18_139/a_484_472# FILLER_0_19_142/a_124_375# 0.001723f
C15131 net47 _452_/a_36_151# 0.021978f
C15132 _118_ _124_ 0.652002f
C15133 output43/a_224_472# vss -0.005182f
C15134 _131_ FILLER_0_17_104/a_36_472# 0.004125f
C15135 _091_ FILLER_0_13_212/a_124_375# 0.025558f
C15136 result[8] mask\[6\] 0.111221f
C15137 vss _107_ 0.186994f
C15138 net74 net36 0.012494f
C15139 net69 net49 0.051235f
C15140 _437_/a_36_151# vdd 0.115376f
C15141 FILLER_0_3_172/a_124_375# FILLER_0_2_171/a_124_375# 0.026339f
C15142 _449_/a_796_472# _038_ 0.018626f
C15143 cal_itt\[3\] _374_/a_36_68# 0.001569f
C15144 _306_/a_36_68# state\[1\] 0.028553f
C15145 _430_/a_1308_423# net63 0.01125f
C15146 FILLER_0_3_172/a_36_472# vdd 0.006145f
C15147 FILLER_0_3_172/a_3260_375# vss 0.054783f
C15148 FILLER_0_5_198/a_124_375# net21 0.029659f
C15149 output18/a_224_472# output19/a_224_472# 0.00124f
C15150 FILLER_0_15_290/a_36_472# result[3] 0.014709f
C15151 _412_/a_2665_112# net18 0.001321f
C15152 net16 _444_/a_2248_156# 0.065914f
C15153 _264_/a_224_472# _084_ 0.007508f
C15154 cal_itt\[1\] cal_itt\[0\] 0.055355f
C15155 _052_ FILLER_0_18_37/a_1020_375# 0.001287f
C15156 FILLER_0_21_286/a_36_472# _420_/a_36_151# 0.059367f
C15157 FILLER_0_10_28/a_36_472# output6/a_224_472# 0.010475f
C15158 _430_/a_1204_472# net63 0.013728f
C15159 net37 FILLER_0_5_148/a_484_472# 0.001212f
C15160 _077_ _439_/a_448_472# 0.052962f
C15161 net81 FILLER_0_14_235/a_484_472# 0.015266f
C15162 fanout76/a_36_160# vss 0.028897f
C15163 FILLER_0_18_76/a_572_375# net71 0.006025f
C15164 _144_ _433_/a_448_472# 0.075144f
C15165 ctln[7] net52 0.06558f
C15166 _043_ net21 0.033824f
C15167 _192_/a_67_603# _416_/a_2665_112# 0.012638f
C15168 vdd _416_/a_2665_112# 0.027256f
C15169 net46 vss 0.110452f
C15170 _422_/a_2665_112# _108_ 0.023365f
C15171 FILLER_0_7_195/a_124_375# _055_ 0.001597f
C15172 output35/a_224_472# net21 0.069263f
C15173 FILLER_0_5_88/a_36_472# vdd 0.090268f
C15174 FILLER_0_5_88/a_124_375# vss 0.015423f
C15175 FILLER_0_8_107/a_36_472# _134_ 0.005632f
C15176 FILLER_0_8_263/a_124_375# _426_/a_36_151# 0.001252f
C15177 _422_/a_2665_112# net19 0.006987f
C15178 mask\[3\] fanout63/a_36_160# 0.002585f
C15179 FILLER_0_10_214/a_36_472# _247_/a_36_160# 0.004828f
C15180 FILLER_0_11_142/a_484_472# cal_count\[3\] 0.014314f
C15181 FILLER_0_22_177/a_1468_375# mask\[6\] 0.002149f
C15182 net35 FILLER_0_22_177/a_1020_375# 0.008333f
C15183 _195_/a_67_603# vss 0.002638f
C15184 _130_ FILLER_0_11_124/a_124_375# 0.001943f
C15185 _189_/a_67_603# mask\[0\] 0.043158f
C15186 ctln[8] output16/a_224_472# 0.006971f
C15187 _013_ FILLER_0_17_64/a_36_472# 0.001991f
C15188 _008_ output32/a_224_472# 0.074809f
C15189 FILLER_0_15_72/a_124_375# FILLER_0_13_72/a_36_472# 0.001418f
C15190 net15 _176_ 0.038396f
C15191 FILLER_0_5_109/a_572_375# _154_ 0.014669f
C15192 _055_ net22 0.084669f
C15193 _176_ FILLER_0_11_78/a_36_472# 0.003603f
C15194 fanout81/a_36_160# net76 0.001905f
C15195 FILLER_0_18_2/a_3260_375# FILLER_0_19_28/a_484_472# 0.001684f
C15196 FILLER_0_2_165/a_36_472# vss 0.001099f
C15197 FILLER_0_4_49/a_36_472# net49 0.010951f
C15198 FILLER_0_9_223/a_572_375# _076_ 0.034523f
C15199 FILLER_0_5_198/a_484_472# net22 0.012457f
C15200 result[1] FILLER_0_11_282/a_36_472# 0.01775f
C15201 _140_ _049_ 0.003069f
C15202 FILLER_0_12_124/a_124_375# net74 0.049113f
C15203 _395_/a_36_488# state\[1\] 0.002702f
C15204 _116_ _267_/a_36_472# 0.029316f
C15205 _025_ FILLER_0_22_107/a_124_375# 0.001891f
C15206 fanout71/a_36_113# net54 0.001194f
C15207 trim_mask\[1\] FILLER_0_6_90/a_484_472# 0.014443f
C15208 FILLER_0_2_177/a_484_472# net22 0.001324f
C15209 output43/a_224_472# net46 0.0215f
C15210 net31 output34/a_224_472# 0.165772f
C15211 _031_ net14 0.00913f
C15212 _103_ _419_/a_448_472# 0.001207f
C15213 net72 FILLER_0_18_37/a_124_375# 0.05632f
C15214 cal net4 0.026084f
C15215 mask\[3\] _432_/a_36_151# 0.002148f
C15216 ctln[8] _447_/a_2665_112# 0.001271f
C15217 FILLER_0_14_107/a_932_472# _043_ 0.0017f
C15218 _051_ vdd 0.036931f
C15219 FILLER_0_13_100/a_124_375# vdd 0.039324f
C15220 FILLER_0_9_28/a_1020_375# _054_ 0.002273f
C15221 FILLER_0_8_138/a_124_375# _313_/a_67_603# 0.00744f
C15222 _077_ FILLER_0_7_72/a_2812_375# 0.002969f
C15223 _033_ _166_ 0.004448f
C15224 net26 net55 0.002901f
C15225 _136_ FILLER_0_14_99/a_124_375# 0.007209f
C15226 net34 FILLER_0_22_128/a_1828_472# 0.005158f
C15227 result[9] FILLER_0_23_274/a_124_375# 0.003102f
C15228 _184_ vss 0.068129f
C15229 _415_/a_1204_472# vdd 0.00108f
C15230 _178_ _184_ 0.436202f
C15231 state\[1\] FILLER_0_13_142/a_1468_375# 0.010245f
C15232 trim_mask\[2\] net68 0.099597f
C15233 result[7] _421_/a_1204_472# 0.014927f
C15234 _128_ net74 0.121254f
C15235 net63 _430_/a_448_472# 0.026599f
C15236 FILLER_0_11_101/a_484_472# FILLER_0_11_109/a_36_472# 0.013276f
C15237 _093_ FILLER_0_21_60/a_484_472# 0.001396f
C15238 mask\[5\] _145_ 0.012075f
C15239 _091_ _223_/a_36_160# 0.001976f
C15240 _130_ _428_/a_2248_156# 0.006602f
C15241 _013_ _424_/a_796_472# 0.032857f
C15242 _420_/a_796_472# vss 0.001659f
C15243 _095_ FILLER_0_14_107/a_36_472# 0.011439f
C15244 net16 net51 0.035455f
C15245 _086_ FILLER_0_4_177/a_36_472# 0.001464f
C15246 _086_ _375_/a_692_497# 0.002565f
C15247 FILLER_0_4_185/a_124_375# _087_ 0.120668f
C15248 fanout73/a_36_113# net70 0.00238f
C15249 _435_/a_2248_156# net21 0.012406f
C15250 _359_/a_1044_488# _152_ 0.001339f
C15251 net4 FILLER_0_12_220/a_36_472# 0.019348f
C15252 FILLER_0_10_28/a_124_375# _450_/a_3129_107# 0.010735f
C15253 _432_/a_2665_112# net80 0.041304f
C15254 FILLER_0_5_128/a_36_472# _133_ 0.001217f
C15255 output46/a_224_472# trimb[3] 0.050924f
C15256 _021_ mask\[5\] 0.001088f
C15257 FILLER_0_9_28/a_572_375# net50 0.002807f
C15258 _130_ _114_ 0.002404f
C15259 output47/a_224_472# FILLER_0_15_2/a_484_472# 0.038484f
C15260 _155_ net50 0.012085f
C15261 _444_/a_1308_423# net67 0.021684f
C15262 _177_ _451_/a_2449_156# 0.002085f
C15263 output23/a_224_472# ctlp[5] 0.005152f
C15264 net72 _394_/a_718_524# 0.001558f
C15265 net55 _394_/a_728_93# 0.0026f
C15266 net63 mask\[2\] 0.553545f
C15267 _136_ _139_ 0.394888f
C15268 net52 _443_/a_1308_423# 0.02003f
C15269 trim_mask\[2\] _156_ 0.018332f
C15270 _446_/a_2560_156# net66 0.002649f
C15271 _119_ vss 0.22921f
C15272 FILLER_0_17_72/a_36_472# FILLER_0_17_64/a_124_375# 0.009654f
C15273 _071_ vss 0.126519f
C15274 net35 _436_/a_36_151# 0.014669f
C15275 _305_/a_36_159# _316_/a_124_24# 0.003478f
C15276 FILLER_0_3_78/a_124_375# _160_ 0.003276f
C15277 _000_ net58 0.00389f
C15278 _322_/a_692_472# _070_ 0.002328f
C15279 net48 _251_/a_244_472# 0.001259f
C15280 net26 net17 0.132516f
C15281 _233_/a_36_160# FILLER_0_6_37/a_124_375# 0.001713f
C15282 FILLER_0_5_72/a_932_472# FILLER_0_6_79/a_36_472# 0.026657f
C15283 output35/a_224_472# mask\[7\] 0.004608f
C15284 ctln[4] net21 0.009947f
C15285 output31/a_224_472# vss -0.003316f
C15286 FILLER_0_16_89/a_1380_472# vss 0.005351f
C15287 net40 _034_ 0.04333f
C15288 _076_ FILLER_0_8_156/a_484_472# 0.008487f
C15289 net57 net70 0.012088f
C15290 _131_ cal_count\[1\] 0.001497f
C15291 _316_/a_848_380# net37 0.01216f
C15292 FILLER_0_20_193/a_484_472# _098_ 0.012457f
C15293 FILLER_0_9_28/a_1828_472# _120_ 0.00108f
C15294 FILLER_0_20_177/a_1020_375# _434_/a_36_151# 0.059049f
C15295 _275_/a_224_472# vss 0.001498f
C15296 FILLER_0_4_99/a_124_375# vdd 0.029154f
C15297 _185_ _180_ 0.001053f
C15298 net32 _419_/a_36_151# 0.006506f
C15299 FILLER_0_16_154/a_1020_375# vss 0.001453f
C15300 FILLER_0_16_154/a_1468_375# vdd 0.017574f
C15301 _068_ _229_/a_224_472# 0.002601f
C15302 _341_/a_49_472# vdd 0.026636f
C15303 _027_ vss 0.011873f
C15304 _055_ vdd 0.406945f
C15305 _424_/a_36_151# _423_/a_1308_423# 0.001722f
C15306 FILLER_0_20_193/a_484_472# _205_/a_36_160# 0.001684f
C15307 output22/a_224_472# _024_ 0.029795f
C15308 ctln[6] net69 0.003695f
C15309 net22 _204_/a_67_603# 0.006495f
C15310 _389_/a_36_148# _172_ 0.039684f
C15311 FILLER_0_22_86/a_484_472# net14 0.006746f
C15312 _065_ _441_/a_448_472# 0.001973f
C15313 _386_/a_124_24# net37 0.00431f
C15314 _132_ FILLER_0_18_107/a_2724_472# 0.002229f
C15315 _420_/a_2248_156# _108_ 0.021735f
C15316 _177_ net36 0.371814f
C15317 net20 _055_ 0.203142f
C15318 FILLER_0_2_177/a_484_472# vdd 0.008489f
C15319 _089_ _002_ 0.002349f
C15320 net19 _420_/a_2248_156# 0.058662f
C15321 FILLER_0_17_161/a_124_375# mask\[2\] 0.00227f
C15322 FILLER_0_13_142/a_1380_472# _225_/a_36_160# 0.004111f
C15323 net20 _419_/a_1204_472# 0.006482f
C15324 _142_ FILLER_0_17_142/a_124_375# 0.011387f
C15325 FILLER_0_15_116/a_124_375# _451_/a_36_151# 0.006111f
C15326 mask\[1\] _043_ 0.027561f
C15327 net76 FILLER_0_3_172/a_484_472# 0.002542f
C15328 _050_ net14 0.001835f
C15329 comp _190_/a_36_160# 0.001891f
C15330 _255_/a_224_552# vdd 0.082462f
C15331 _095_ _278_/a_36_160# 0.030448f
C15332 mask\[8\] _354_/a_49_472# 0.105272f
C15333 _126_ vdd 0.682779f
C15334 FILLER_0_24_96/a_124_375# output24/a_224_472# 0.00363f
C15335 _019_ net36 0.309649f
C15336 FILLER_0_13_206/a_124_375# net4 0.031251f
C15337 result[9] FILLER_0_24_274/a_1020_375# 0.001657f
C15338 net53 FILLER_0_14_99/a_124_375# 0.00494f
C15339 _412_/a_1308_423# net76 0.023786f
C15340 _414_/a_1000_472# _089_ 0.001754f
C15341 _008_ _094_ 0.234346f
C15342 FILLER_0_13_212/a_1020_375# net79 0.009597f
C15343 FILLER_0_24_96/a_124_375# vss 0.017357f
C15344 FILLER_0_17_226/a_36_472# _093_ 0.004282f
C15345 net62 FILLER_0_13_212/a_1468_375# 0.003327f
C15346 net4 net37 0.021795f
C15347 ctln[6] ctln[7] 0.00499f
C15348 _095_ vss 1.465527f
C15349 _178_ _095_ 0.839141f
C15350 FILLER_0_19_47/a_124_375# _182_ 0.001771f
C15351 FILLER_0_16_107/a_36_472# _093_ 0.001526f
C15352 net4 FILLER_0_3_221/a_1468_375# 0.006974f
C15353 _261_/a_36_160# net23 0.005015f
C15354 FILLER_0_18_171/a_36_472# _098_ 0.020038f
C15355 _326_/a_36_160# _115_ 0.051266f
C15356 mask\[7\] _435_/a_2248_156# 0.026974f
C15357 result[8] _422_/a_1308_423# 0.001356f
C15358 output8/a_224_472# net59 0.00398f
C15359 _414_/a_2665_112# net22 0.004067f
C15360 net58 FILLER_0_9_290/a_124_375# 0.001157f
C15361 net76 FILLER_0_5_181/a_124_375# 0.031324f
C15362 _021_ net80 0.254353f
C15363 net63 FILLER_0_15_212/a_572_375# 0.001597f
C15364 FILLER_0_1_212/a_124_375# vdd 0.020159f
C15365 output12/a_224_472# FILLER_0_0_198/a_36_472# 0.023414f
C15366 FILLER_0_15_142/a_572_375# vdd -0.013698f
C15367 _011_ net78 0.002956f
C15368 _036_ vss 0.161195f
C15369 cal_count\[1\] FILLER_0_13_80/a_36_472# 0.001559f
C15370 _084_ net8 0.001821f
C15371 net27 FILLER_0_11_282/a_124_375# 0.002857f
C15372 output26/a_224_472# vss 0.0137f
C15373 _077_ _162_ 0.013298f
C15374 FILLER_0_12_220/a_572_375# vdd -0.014642f
C15375 FILLER_0_12_220/a_124_375# vss 0.040895f
C15376 FILLER_0_4_197/a_1468_375# _088_ 0.012367f
C15377 fanout50/a_36_160# _447_/a_2665_112# 0.002885f
C15378 net58 _411_/a_2665_112# 0.018133f
C15379 _426_/a_1000_472# calibrate 0.002865f
C15380 FILLER_0_18_139/a_932_472# vdd 0.002904f
C15381 FILLER_0_18_139/a_484_472# vss 0.006719f
C15382 net20 FILLER_0_1_212/a_124_375# 0.084041f
C15383 FILLER_0_4_123/a_36_472# _370_/a_124_24# 0.003595f
C15384 result[9] FILLER_0_15_282/a_124_375# 0.001233f
C15385 _432_/a_1204_472# vdd 0.004019f
C15386 _408_/a_1936_472# _067_ 0.003007f
C15387 output25/a_224_472# _213_/a_67_603# 0.032497f
C15388 FILLER_0_21_125/a_484_472# mask\[7\] 0.003404f
C15389 FILLER_0_9_72/a_1380_472# _439_/a_36_151# 0.001723f
C15390 FILLER_0_15_282/a_484_472# net18 0.018113f
C15391 ctln[1] net1 0.003756f
C15392 trim_val\[3\] _168_ 0.271475f
C15393 FILLER_0_5_72/a_124_375# _029_ 0.010208f
C15394 FILLER_0_22_177/a_1020_375# vdd 0.001695f
C15395 FILLER_0_18_107/a_932_472# mask\[9\] 0.005296f
C15396 net19 _419_/a_2665_112# 0.00276f
C15397 output48/a_224_472# net76 0.069862f
C15398 _077_ _131_ 0.03465f
C15399 state\[1\] net22 0.007096f
C15400 _110_ mask\[9\] 0.00319f
C15401 _390_/a_244_472# _038_ 0.001278f
C15402 _390_/a_36_68# _136_ 0.032598f
C15403 net20 FILLER_0_12_220/a_572_375# 0.007386f
C15404 _447_/a_2248_156# _030_ 0.001588f
C15405 _104_ FILLER_0_17_226/a_124_375# 0.024833f
C15406 FILLER_0_4_144/a_124_375# _081_ 0.004558f
C15407 FILLER_0_18_139/a_124_375# FILLER_0_18_107/a_3260_375# 0.012552f
C15408 cal_count\[2\] _179_ 0.404284f
C15409 _081_ FILLER_0_8_156/a_484_472# 0.001772f
C15410 net7 _239_/a_36_160# 0.068281f
C15411 _426_/a_796_472# net64 0.006933f
C15412 FILLER_0_4_107/a_572_375# _160_ 0.008945f
C15413 FILLER_0_17_282/a_124_375# net30 0.001288f
C15414 FILLER_0_1_192/a_124_375# net59 0.014491f
C15415 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_124_375# 0.003732f
C15416 _418_/a_36_151# net77 0.019316f
C15417 FILLER_0_17_72/a_124_375# _131_ 0.006224f
C15418 net3 cal_count\[2\] 0.119728f
C15419 _081_ _265_/a_916_472# 0.002264f
C15420 _204_/a_67_603# vdd 0.039556f
C15421 _435_/a_1288_156# vdd 0.001119f
C15422 _367_/a_244_472# vdd 0.001113f
C15423 _105_ output35/a_224_472# 0.013092f
C15424 FILLER_0_10_78/a_572_375# _176_ 0.005927f
C15425 _449_/a_1308_423# vdd 0.002584f
C15426 _449_/a_448_472# vss 0.032274f
C15427 _008_ net78 0.032202f
C15428 _405_/a_67_603# net47 0.004116f
C15429 _153_ _365_/a_692_472# 0.002377f
C15430 FILLER_0_21_286/a_124_375# net77 0.00301f
C15431 _141_ FILLER_0_22_128/a_3172_472# 0.01947f
C15432 state\[0\] _072_ 0.030642f
C15433 output12/a_224_472# net11 0.009336f
C15434 _443_/a_1204_472# net23 0.026261f
C15435 result[1] vdd 0.221634f
C15436 net4 _264_/a_224_472# 0.001408f
C15437 en cal_itt\[1\] 0.028447f
C15438 input3/a_36_113# net3 0.015124f
C15439 _443_/a_2248_156# trim_mask\[4\] 0.002315f
C15440 _126_ _135_ 0.011447f
C15441 mask\[9\] _437_/a_2665_112# 0.014146f
C15442 _026_ _437_/a_448_472# 0.026072f
C15443 vss output41/a_224_472# -0.007739f
C15444 fanout49/a_36_160# FILLER_0_3_78/a_572_375# 0.00805f
C15445 net63 FILLER_0_15_205/a_124_375# 0.001597f
C15446 _451_/a_36_151# _040_ 0.018648f
C15447 trim_mask\[1\] net14 0.024935f
C15448 _413_/a_36_151# net82 0.00601f
C15449 net15 FILLER_0_17_64/a_124_375# 0.047331f
C15450 _122_ FILLER_0_6_231/a_572_375# 0.016091f
C15451 _131_ _120_ 0.191602f
C15452 net41 _446_/a_2560_156# 0.005695f
C15453 _104_ net32 0.342568f
C15454 FILLER_0_14_263/a_36_472# output30/a_224_472# 0.002002f
C15455 _031_ _153_ 0.009316f
C15456 _402_/a_728_93# vdd 0.050988f
C15457 _178_ _402_/a_1296_93# 0.062418f
C15458 FILLER_0_7_233/a_36_472# FILLER_0_6_231/a_124_375# 0.001684f
C15459 trim_mask\[1\] _164_ 0.195956f
C15460 net82 _078_ 0.00197f
C15461 net50 FILLER_0_8_24/a_36_472# 0.015187f
C15462 _363_/a_36_68# _151_ 0.020916f
C15463 _068_ _247_/a_36_160# 0.003213f
C15464 _132_ _428_/a_1000_472# 0.027767f
C15465 FILLER_0_12_236/a_36_472# vss 0.001526f
C15466 FILLER_0_12_236/a_484_472# vdd 0.00923f
C15467 output37/a_224_472# vss 0.026983f
C15468 FILLER_0_18_2/a_124_375# trimb[1] 0.01352f
C15469 FILLER_0_15_282/a_36_472# _417_/a_1308_423# 0.001295f
C15470 _414_/a_2665_112# vdd 0.006496f
C15471 FILLER_0_14_91/a_36_472# vss 0.001729f
C15472 FILLER_0_14_91/a_484_472# vdd 0.00605f
C15473 _157_ net14 0.026868f
C15474 _385_/a_36_68# vss 0.002408f
C15475 _442_/a_796_472# _031_ 0.013039f
C15476 _372_/a_170_472# _059_ 0.033956f
C15477 FILLER_0_16_73/a_124_375# _176_ 0.006386f
C15478 FILLER_0_21_28/a_1828_472# vdd 0.004227f
C15479 FILLER_0_21_28/a_1380_472# vss 0.001688f
C15480 FILLER_0_16_107/a_36_472# _136_ 0.011469f
C15481 mask\[0\] _043_ 0.929722f
C15482 net50 FILLER_0_2_93/a_484_472# 0.002377f
C15483 FILLER_0_3_221/a_124_375# vdd 0.008869f
C15484 _436_/a_36_151# vdd 0.078019f
C15485 output23/a_224_472# _050_ 0.014495f
C15486 _423_/a_796_472# _012_ 0.015809f
C15487 FILLER_0_17_282/a_124_375# _417_/a_36_151# 0.059049f
C15488 FILLER_0_1_192/a_36_472# net21 0.016033f
C15489 FILLER_0_13_100/a_36_472# _043_ 0.012726f
C15490 _093_ _397_/a_36_472# 0.001509f
C15491 _104_ _422_/a_2560_156# 0.003223f
C15492 net36 _438_/a_448_472# 0.034338f
C15493 mask\[9\] net14 0.090939f
C15494 _439_/a_36_151# vdd 0.095368f
C15495 _274_/a_36_68# net64 0.036017f
C15496 net81 _426_/a_36_151# 0.060652f
C15497 net36 _451_/a_2225_156# 0.044144f
C15498 net54 _437_/a_2560_156# 0.009745f
C15499 _013_ _052_ 0.284735f
C15500 net47 FILLER_0_5_136/a_36_472# 0.006139f
C15501 FILLER_0_21_28/a_1916_375# _424_/a_36_151# 0.059049f
C15502 net79 result[3] 0.138076f
C15503 state\[1\] vdd 0.544231f
C15504 FILLER_0_10_78/a_484_472# _115_ 0.005678f
C15505 net15 _030_ 0.355335f
C15506 mask\[5\] net32 0.304094f
C15507 FILLER_0_14_50/a_124_375# _180_ 0.022435f
C15508 _050_ _148_ 0.002456f
C15509 net1 fanout58/a_36_160# 0.060243f
C15510 _085_ net23 0.020463f
C15511 net3 _043_ 0.004313f
C15512 _091_ FILLER_0_18_177/a_36_472# 0.012695f
C15513 _095_ _184_ 0.265966f
C15514 net69 _370_/a_124_24# 0.001491f
C15515 _095_ _401_/a_36_68# 0.001398f
C15516 _341_/a_49_472# FILLER_0_16_154/a_572_375# 0.001643f
C15517 _007_ vdd 0.129966f
C15518 _321_/a_358_69# net23 0.001718f
C15519 _449_/a_2248_156# cal_count\[3\] 0.002041f
C15520 net16 net47 0.089651f
C15521 _002_ FILLER_0_3_172/a_1916_375# 0.047331f
C15522 _064_ net49 0.377675f
C15523 net28 _416_/a_2665_112# 0.008877f
C15524 ctln[3] net75 0.066513f
C15525 _432_/a_1000_472# vdd 0.010431f
C15526 _428_/a_2665_112# FILLER_0_13_142/a_36_472# 0.003706f
C15527 FILLER_0_0_266/a_124_375# vdd 0.006328f
C15528 fanout75/a_36_113# net1 0.011428f
C15529 FILLER_0_10_78/a_36_472# vss 0.008832f
C15530 FILLER_0_18_2/a_2276_472# net38 0.002313f
C15531 _112_ _081_ 0.037903f
C15532 FILLER_0_9_28/a_1468_375# _444_/a_2248_156# 0.001074f
C15533 FILLER_0_16_57/a_1468_375# _176_ 0.006445f
C15534 FILLER_0_4_49/a_572_375# FILLER_0_5_54/a_36_472# 0.001723f
C15535 FILLER_0_5_109/a_124_375# _163_ 0.002658f
C15536 result[6] _421_/a_2248_156# 0.031832f
C15537 cal_itt\[3\] net59 0.018616f
C15538 _131_ FILLER_0_17_56/a_484_472# 0.002672f
C15539 FILLER_0_3_142/a_36_472# _261_/a_36_160# 0.001542f
C15540 net67 output6/a_224_472# 0.070024f
C15541 _033_ net17 0.028529f
C15542 net18 FILLER_0_11_282/a_124_375# 0.042342f
C15543 FILLER_0_4_177/a_36_472# _163_ 0.002787f
C15544 _370_/a_124_24# _152_ 0.069015f
C15545 _370_/a_848_380# _081_ 0.035068f
C15546 FILLER_0_21_142/a_484_472# _098_ 0.001158f
C15547 _167_ _160_ 0.157458f
C15548 _053_ _054_ 0.015389f
C15549 net60 _418_/a_796_472# 0.008602f
C15550 trim[1] net66 0.007756f
C15551 net27 _189_/a_67_603# 0.008028f
C15552 net24 FILLER_0_23_88/a_124_375# 0.020193f
C15553 _069_ _055_ 0.741952f
C15554 _077_ _074_ 0.148596f
C15555 _091_ _432_/a_448_472# 0.050539f
C15556 _028_ FILLER_0_7_104/a_124_375# 0.008248f
C15557 _426_/a_2248_156# vss 0.002303f
C15558 _426_/a_2665_112# vdd 0.008893f
C15559 _070_ _310_/a_49_472# 0.00564f
C15560 _147_ vss 0.006333f
C15561 net74 FILLER_0_5_136/a_36_472# 0.003704f
C15562 _175_ _131_ 0.050098f
C15563 mask\[4\] _141_ 0.948091f
C15564 _444_/a_2665_112# _164_ 0.015644f
C15565 _176_ FILLER_0_15_59/a_484_472# 0.007596f
C15566 trim[4] net44 0.188184f
C15567 _132_ FILLER_0_17_104/a_484_472# 0.002737f
C15568 output27/a_224_472# FILLER_0_9_282/a_484_472# 0.001711f
C15569 output9/a_224_472# net59 0.051763f
C15570 net50 FILLER_0_4_91/a_572_375# 0.007234f
C15571 _077_ _076_ 1.895143f
C15572 net29 _287_/a_36_472# 0.002936f
C15573 _141_ _142_ 0.200324f
C15574 net70 net36 0.066607f
C15575 _053_ vss 0.85895f
C15576 net20 _426_/a_2665_112# 0.018602f
C15577 net27 result[0] 0.106157f
C15578 fanout74/a_36_113# net82 0.018392f
C15579 _274_/a_2552_68# vss 0.003123f
C15580 FILLER_0_4_185/a_124_375# _272_/a_36_472# 0.001781f
C15581 cal_itt\[3\] _122_ 0.03282f
C15582 _114_ FILLER_0_10_94/a_572_375# 0.008375f
C15583 FILLER_0_8_127/a_36_472# _058_ 0.003283f
C15584 _176_ net74 0.067915f
C15585 FILLER_0_6_47/a_2812_375# vss 0.035758f
C15586 FILLER_0_6_47/a_3260_375# vdd 0.003435f
C15587 FILLER_0_14_107/a_484_472# _451_/a_36_151# 0.001723f
C15588 net73 FILLER_0_17_133/a_36_472# 0.049294f
C15589 net79 _056_ 0.022406f
C15590 net15 FILLER_0_15_72/a_124_375# 0.006566f
C15591 net18 FILLER_0_13_290/a_36_472# 0.079901f
C15592 output35/a_224_472# result[8] 0.016867f
C15593 _332_/a_244_68# _135_ 0.001325f
C15594 _096_ cal_count\[3\] 0.016393f
C15595 FILLER_0_16_107/a_484_472# net70 0.002732f
C15596 cal_count\[2\] _402_/a_56_567# 0.07745f
C15597 _402_/a_1296_93# _401_/a_36_68# 0.001523f
C15598 net36 FILLER_0_15_228/a_124_375# 0.00167f
C15599 FILLER_0_13_65/a_36_472# vss 0.007545f
C15600 FILLER_0_4_99/a_36_472# _156_ 0.0255f
C15601 _053_ FILLER_0_7_72/a_36_472# 0.01287f
C15602 FILLER_0_13_212/a_124_375# vdd 0.010978f
C15603 _093_ FILLER_0_17_218/a_124_375# 0.003338f
C15604 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_572_375# 0.086635f
C15605 FILLER_0_6_90/a_36_472# net14 0.002705f
C15606 fanout67/a_36_160# _439_/a_36_151# 0.00246f
C15607 _050_ _436_/a_2665_112# 0.030939f
C15608 _062_ net23 0.061239f
C15609 FILLER_0_9_28/a_1468_375# net51 0.00111f
C15610 output38/a_224_472# net49 0.002434f
C15611 FILLER_0_7_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001723f
C15612 _377_/a_36_472# _165_ 0.025689f
C15613 FILLER_0_11_101/a_124_375# _120_ 0.008016f
C15614 net74 _124_ 0.180235f
C15615 net32 net34 0.330134f
C15616 _446_/a_36_151# net17 0.006518f
C15617 _076_ _120_ 0.736844f
C15618 _104_ _420_/a_2665_112# 0.053555f
C15619 net16 _173_ 0.029412f
C15620 net79 _286_/a_224_472# 0.001276f
C15621 ctln[2] net76 0.001008f
C15622 _025_ net71 0.030824f
C15623 FILLER_0_8_37/a_572_375# _054_ 0.137749f
C15624 _424_/a_2560_156# vss 0.001554f
C15625 vdd FILLER_0_21_60/a_124_375# 0.014029f
C15626 net32 net60 0.509175f
C15627 net73 FILLER_0_18_107/a_124_375# 0.003742f
C15628 net4 net8 0.00647f
C15629 _265_/a_244_68# net59 0.001147f
C15630 net55 FILLER_0_17_72/a_1020_375# 0.049648f
C15631 _422_/a_36_151# _421_/a_2248_156# 0.001189f
C15632 _096_ _320_/a_672_472# 0.0082f
C15633 output35/a_224_472# FILLER_0_22_177/a_1468_375# 0.018187f
C15634 _410_/a_36_68# cal_count\[3\] 0.001096f
C15635 _000_ _411_/a_1204_472# 0.002575f
C15636 mask\[9\] _148_ 0.01635f
C15637 result[9] _417_/a_2665_112# 0.060365f
C15638 output29/a_224_472# _045_ 0.002303f
C15639 FILLER_0_6_239/a_36_472# fanout75/a_36_113# 0.00191f
C15640 FILLER_0_16_57/a_932_472# net15 0.037807f
C15641 FILLER_0_1_98/a_36_472# net14 0.023583f
C15642 FILLER_0_8_37/a_572_375# vss 0.00282f
C15643 FILLER_0_8_37/a_36_472# vdd 0.135405f
C15644 _207_/a_67_603# FILLER_0_22_128/a_3172_472# 0.005759f
C15645 FILLER_0_12_136/a_1380_472# vss 0.031524f
C15646 _449_/a_2665_112# _176_ 0.048319f
C15647 FILLER_0_21_28/a_2364_375# _012_ 0.017669f
C15648 net65 FILLER_0_3_212/a_124_375# 0.003807f
C15649 net1 net18 0.047886f
C15650 FILLER_0_5_72/a_36_472# vss 0.031034f
C15651 FILLER_0_5_72/a_484_472# vdd 0.002735f
C15652 _031_ FILLER_0_2_111/a_932_472# 0.017509f
C15653 _270_/a_36_472# net76 0.009569f
C15654 FILLER_0_12_136/a_1020_375# FILLER_0_11_142/a_484_472# 0.001543f
C15655 en_co_clk _120_ 0.008507f
C15656 en_co_clk _038_ 0.014475f
C15657 _050_ FILLER_0_22_128/a_1468_375# 0.001661f
C15658 _098_ FILLER_0_19_171/a_36_472# 0.021559f
C15659 FILLER_0_5_54/a_572_375# trim_mask\[1\] 0.011664f
C15660 _075_ _078_ 0.001896f
C15661 FILLER_0_1_98/a_124_375# trim_mask\[3\] 0.058544f
C15662 FILLER_0_20_87/a_124_375# vss 0.00279f
C15663 FILLER_0_20_87/a_36_472# vdd 0.006784f
C15664 _127_ net53 0.00917f
C15665 fanout52/a_36_160# _170_ 0.024724f
C15666 _451_/a_1353_112# vdd 0.009693f
C15667 _153_ _157_ 0.050552f
C15668 FILLER_0_21_286/a_36_472# _009_ 0.003266f
C15669 _446_/a_1204_472# net40 0.026414f
C15670 FILLER_0_8_127/a_124_375# _126_ 0.001799f
C15671 _426_/a_36_151# FILLER_0_8_247/a_36_472# 0.001723f
C15672 _070_ FILLER_0_10_94/a_124_375# 0.008294f
C15673 _304_/a_224_472# _111_ 0.003461f
C15674 vss _166_ 0.011302f
C15675 FILLER_0_7_72/a_2276_472# vdd 0.004035f
C15676 vdd _160_ 0.606139f
C15677 FILLER_0_10_78/a_124_375# _453_/a_2665_112# 0.006271f
C15678 _086_ _077_ 0.058673f
C15679 _375_/a_36_68# vss 0.02182f
C15680 _326_/a_36_160# vdd 0.066545f
C15681 output10/a_224_472# FILLER_0_0_232/a_124_375# 0.00363f
C15682 FILLER_0_15_150/a_36_472# vss 0.00975f
C15683 FILLER_0_12_2/a_124_375# _450_/a_36_151# 0.001543f
C15684 net57 _085_ 0.211414f
C15685 _131_ FILLER_0_9_105/a_572_375# 0.031928f
C15686 _008_ _418_/a_2248_156# 0.047066f
C15687 FILLER_0_2_93/a_484_472# FILLER_0_2_101/a_36_472# 0.013277f
C15688 _185_ _278_/a_36_160# 0.001237f
C15689 net63 FILLER_0_19_187/a_124_375# 0.012282f
C15690 _165_ FILLER_0_6_37/a_124_375# 0.002884f
C15691 FILLER_0_11_124/a_36_472# vss 0.002545f
C15692 _267_/a_1792_472# _055_ 0.003058f
C15693 FILLER_0_19_55/a_36_472# net55 0.062683f
C15694 trimb[1] FILLER_0_19_28/a_124_375# 0.00285f
C15695 mask\[4\] FILLER_0_18_177/a_124_375# 0.016093f
C15696 _223_/a_36_160# vdd 0.018653f
C15697 _185_ vss 0.021437f
C15698 ctln[4] FILLER_0_1_212/a_36_472# 0.006408f
C15699 _413_/a_36_151# net21 0.012223f
C15700 fanout82/a_36_113# net19 0.021188f
C15701 _430_/a_36_151# _138_ 0.001123f
C15702 _178_ _185_ 0.979797f
C15703 FILLER_0_18_2/a_2724_472# net47 0.001551f
C15704 net66 FILLER_0_3_54/a_36_472# 0.008174f
C15705 _345_/a_36_160# vss 0.003697f
C15706 _372_/a_2590_472# _062_ 0.0012f
C15707 FILLER_0_14_91/a_36_472# _095_ 0.014431f
C15708 _350_/a_665_69# net23 0.001468f
C15709 _128_ FILLER_0_9_142/a_124_375# 0.004439f
C15710 FILLER_0_18_107/a_484_472# net14 0.002472f
C15711 mask\[5\] _434_/a_36_151# 0.00104f
C15712 net62 _100_ 0.006742f
C15713 net81 FILLER_0_15_212/a_1380_472# 0.003953f
C15714 _219_/a_36_160# trim_mask\[0\] 0.395762f
C15715 net20 _223_/a_36_160# 0.066119f
C15716 _091_ _143_ 0.007204f
C15717 FILLER_0_9_223/a_484_472# vss 0.006102f
C15718 ctln[3] net19 0.003077f
C15719 _372_/a_786_69# _163_ 0.001179f
C15720 FILLER_0_18_37/a_124_375# vdd 0.024546f
C15721 FILLER_0_0_130/a_124_375# _442_/a_36_151# 0.059049f
C15722 result[0] net18 0.085445f
C15723 _086_ _120_ 0.408014f
C15724 _447_/a_36_151# net17 0.001448f
C15725 _057_ _267_/a_1120_472# 0.001833f
C15726 _069_ state\[1\] 0.003884f
C15727 output36/a_224_472# vdd 0.145046f
C15728 _003_ _074_ 0.00476f
C15729 net79 _138_ 0.024731f
C15730 FILLER_0_4_177/a_484_472# FILLER_0_3_172/a_932_472# 0.026657f
C15731 vdd net30 0.636147f
C15732 fanout55/a_36_160# _067_ 0.126784f
C15733 _119_ _053_ 0.038651f
C15734 _131_ _125_ 0.013932f
C15735 _177_ _176_ 0.226424f
C15736 net66 _164_ 0.093385f
C15737 FILLER_0_5_72/a_1468_375# FILLER_0_5_88/a_36_472# 0.086635f
C15738 _059_ _313_/a_67_603# 0.061666f
C15739 FILLER_0_10_37/a_36_472# net16 0.012905f
C15740 _093_ FILLER_0_17_72/a_36_472# 0.001971f
C15741 _415_/a_36_151# FILLER_0_8_263/a_124_375# 0.001619f
C15742 FILLER_0_16_37/a_36_472# net72 0.005134f
C15743 _098_ _433_/a_2560_156# 0.004273f
C15744 fanout53/a_36_160# vss 0.006674f
C15745 _428_/a_2665_112# vss 0.005991f
C15746 FILLER_0_20_193/a_484_472# net21 0.00371f
C15747 output7/a_224_472# net41 0.003942f
C15748 _413_/a_1308_423# vdd 0.002686f
C15749 _437_/a_2248_156# net14 0.023718f
C15750 net20 net30 0.033149f
C15751 FILLER_0_24_63/a_36_472# vdd 0.055524f
C15752 _072_ _248_/a_36_68# 0.001683f
C15753 fanout75/a_36_113# net76 0.040306f
C15754 _074_ net1 0.128466f
C15755 _395_/a_36_488# _121_ 0.009689f
C15756 FILLER_0_21_142/a_36_472# net35 0.003079f
C15757 _415_/a_2665_112# result[1] 0.010555f
C15758 _408_/a_718_524# FILLER_0_12_28/a_124_375# 0.001192f
C15759 FILLER_0_13_80/a_124_375# vdd 0.018971f
C15760 _422_/a_2665_112# _009_ 0.061508f
C15761 _178_ _407_/a_36_472# 0.001699f
C15762 vss cal_count\[0\] 0.160743f
C15763 _432_/a_1308_423# FILLER_0_18_177/a_36_472# 0.009119f
C15764 _178_ cal_count\[0\] 0.011488f
C15765 _144_ _437_/a_2665_112# 0.001186f
C15766 _098_ FILLER_0_15_235/a_36_472# 0.093007f
C15767 FILLER_0_20_177/a_932_472# _098_ 0.008366f
C15768 FILLER_0_17_64/a_124_375# FILLER_0_15_59/a_484_472# 0.001188f
C15769 FILLER_0_9_28/a_1916_375# net51 0.001008f
C15770 net57 _062_ 0.067654f
C15771 net55 _452_/a_3129_107# 0.006395f
C15772 _413_/a_2560_156# net65 0.011101f
C15773 _092_ FILLER_0_17_218/a_484_472# 0.007838f
C15774 _444_/a_36_151# net17 0.001435f
C15775 _068_ _311_/a_1920_473# 0.001498f
C15776 net60 _420_/a_2665_112# 0.038894f
C15777 FILLER_0_18_177/a_2364_375# net21 0.018463f
C15778 _098_ vss 0.958032f
C15779 FILLER_0_17_200/a_124_375# FILLER_0_18_177/a_2724_472# 0.001597f
C15780 net15 FILLER_0_5_54/a_1020_375# 0.015944f
C15781 _065_ net52 0.017184f
C15782 _187_ _408_/a_1936_472# 0.017573f
C15783 FILLER_0_3_54/a_124_375# _164_ 0.008654f
C15784 _334_/a_36_160# FILLER_0_17_104/a_1380_472# 0.004111f
C15785 FILLER_0_16_73/a_36_472# vss 0.035175f
C15786 net54 _436_/a_2560_156# 0.010748f
C15787 FILLER_0_21_286/a_484_472# FILLER_0_23_290/a_124_375# 0.001404f
C15788 _091_ net64 0.079488f
C15789 trim_mask\[1\] FILLER_0_6_47/a_2724_472# 0.003645f
C15790 _424_/a_1308_423# _012_ 0.007041f
C15791 FILLER_0_7_72/a_1916_375# net52 0.001608f
C15792 FILLER_0_19_55/a_36_472# _216_/a_67_603# 0.00254f
C15793 net62 FILLER_0_14_235/a_124_375# 0.015659f
C15794 _033_ _444_/a_1308_423# 0.002877f
C15795 net44 FILLER_0_8_2/a_124_375# 0.083677f
C15796 FILLER_0_18_177/a_484_472# FILLER_0_19_171/a_1020_375# 0.001684f
C15797 FILLER_0_8_2/a_36_472# vss 0.004429f
C15798 _118_ _315_/a_36_68# 0.005792f
C15799 _415_/a_448_472# vdd 0.005273f
C15800 _205_/a_36_160# vss 0.003612f
C15801 cal_itt\[2\] FILLER_0_3_221/a_124_375# 0.006217f
C15802 ctln[1] ctln[4] 0.002283f
C15803 net80 _434_/a_36_151# 0.067037f
C15804 _417_/a_36_151# vdd 0.140703f
C15805 _057_ _225_/a_36_160# 0.026341f
C15806 _065_ net49 0.001576f
C15807 FILLER_0_10_78/a_484_472# vdd 0.004673f
C15808 net81 _015_ 0.002818f
C15809 FILLER_0_4_185/a_36_472# vss 0.002627f
C15810 _091_ FILLER_0_19_171/a_1380_472# 0.001044f
C15811 FILLER_0_19_47/a_572_375# vss 0.055293f
C15812 FILLER_0_19_47/a_36_472# vdd 0.072773f
C15813 FILLER_0_9_28/a_1828_472# net68 0.048468f
C15814 net18 _416_/a_1000_472# 0.046085f
C15815 mask\[3\] _102_ 0.142836f
C15816 _101_ _005_ 0.003946f
C15817 _421_/a_36_151# _419_/a_2248_156# 0.001203f
C15818 _431_/a_2248_156# net73 0.003228f
C15819 FILLER_0_4_197/a_572_375# net21 0.041173f
C15820 _374_/a_36_68# vdd 0.075685f
C15821 FILLER_0_12_136/a_1380_472# _071_ 0.004003f
C15822 net35 FILLER_0_22_86/a_572_375# 0.010986f
C15823 mask\[8\] FILLER_0_22_86/a_1020_375# 0.009431f
C15824 net75 _425_/a_1000_472# 0.038919f
C15825 net44 FILLER_0_15_10/a_36_472# 0.012286f
C15826 fanout49/a_36_160# vss 0.025717f
C15827 FILLER_0_7_59/a_124_375# vss 0.002006f
C15828 FILLER_0_7_59/a_572_375# vdd 0.005991f
C15829 FILLER_0_13_212/a_572_375# _043_ 0.01418f
C15830 FILLER_0_22_128/a_3260_375# _146_ 0.004692f
C15831 output42/a_224_472# net42 0.117956f
C15832 net35 FILLER_0_22_128/a_1380_472# 0.016004f
C15833 net79 _113_ 0.002432f
C15834 fanout64/a_36_160# vss 0.007097f
C15835 net33 _146_ 0.306187f
C15836 _069_ FILLER_0_13_212/a_124_375# 0.070185f
C15837 net59 FILLER_0_3_212/a_36_472# 0.058623f
C15838 _387_/a_36_113# vss 0.047621f
C15839 result[4] FILLER_0_17_282/a_124_375# 0.018106f
C15840 _131_ cal_count\[2\] 0.044147f
C15841 net68 FILLER_0_6_47/a_36_472# 0.001248f
C15842 FILLER_0_13_65/a_36_472# _095_ 0.003171f
C15843 ctln[1] _000_ 0.223573f
C15844 _185_ _184_ 0.047803f
C15845 net17 FILLER_0_23_44/a_572_375# 0.001332f
C15846 _291_/a_36_160# FILLER_0_17_226/a_36_472# 0.035111f
C15847 FILLER_0_18_2/a_2364_375# net55 0.005899f
C15848 _077_ FILLER_0_8_107/a_36_472# 0.007552f
C15849 fanout49/a_36_160# _441_/a_2248_156# 0.027388f
C15850 FILLER_0_4_49/a_124_375# _167_ 0.009437f
C15851 _003_ _081_ 0.041822f
C15852 _119_ _375_/a_36_68# 0.007338f
C15853 net60 _419_/a_2560_156# 0.006989f
C15854 net54 FILLER_0_22_128/a_1916_375# 0.001933f
C15855 _444_/a_1204_472# net40 0.017496f
C15856 FILLER_0_1_98/a_36_472# _153_ 0.001463f
C15857 _070_ FILLER_0_9_105/a_484_472# 0.020248f
C15858 _013_ FILLER_0_17_56/a_36_472# 0.002659f
C15859 _086_ _363_/a_36_68# 0.007567f
C15860 _440_/a_2248_156# trim_mask\[1\] 0.004408f
C15861 _133_ vdd 0.27652f
C15862 _070_ vss 1.363355f
C15863 _093_ net54 0.003211f
C15864 FILLER_0_17_72/a_1828_472# _438_/a_36_151# 0.001221f
C15865 _217_/a_36_160# _424_/a_36_151# 0.035111f
C15866 _406_/a_36_159# net47 0.034933f
C15867 FILLER_0_15_180/a_572_375# vdd 0.068901f
C15868 _429_/a_2665_112# FILLER_0_14_235/a_124_375# 0.006271f
C15869 FILLER_0_7_146/a_36_472# vss 0.029149f
C15870 net50 trim_val\[3\] 0.111824f
C15871 _073_ _084_ 0.048469f
C15872 FILLER_0_4_197/a_124_375# FILLER_0_5_198/a_36_472# 0.001723f
C15873 net1 _081_ 0.111227f
C15874 _321_/a_170_472# _395_/a_36_488# 0.007047f
C15875 FILLER_0_16_89/a_484_472# _131_ 0.01075f
C15876 _115_ FILLER_0_10_94/a_484_472# 0.015061f
C15877 FILLER_0_21_28/a_572_375# net40 0.001406f
C15878 FILLER_0_12_136/a_932_472# _126_ 0.014483f
C15879 _163_ FILLER_0_6_79/a_36_472# 0.001789f
C15880 net80 FILLER_0_22_177/a_484_472# 0.005297f
C15881 trim_mask\[2\] FILLER_0_3_78/a_572_375# 0.011713f
C15882 _321_/a_2034_472# _120_ 0.002489f
C15883 _300_/a_224_472# _009_ 0.001405f
C15884 FILLER_0_18_2/a_2364_375# net17 0.048345f
C15885 _317_/a_36_113# vdd 0.054289f
C15886 _063_ trim_val\[0\] 0.001978f
C15887 FILLER_0_14_50/a_36_472# vdd 0.081414f
C15888 FILLER_0_14_50/a_124_375# vss 0.002412f
C15889 _064_ net40 0.141744f
C15890 FILLER_0_6_239/a_36_472# _074_ 0.004715f
C15891 net77 _007_ 0.002591f
C15892 _093_ net15 0.145303f
C15893 _176_ _451_/a_2225_156# 0.030788f
C15894 net68 _440_/a_36_151# 0.080854f
C15895 FILLER_0_17_72/a_3172_472# _131_ 0.003717f
C15896 net67 FILLER_0_6_47/a_36_472# 0.004607f
C15897 _028_ _439_/a_448_472# 0.017606f
C15898 _086_ _311_/a_2180_473# 0.001744f
C15899 _420_/a_2248_156# _009_ 0.00681f
C15900 FILLER_0_16_89/a_124_375# net36 0.011956f
C15901 net1 net65 0.035488f
C15902 _061_ cal_count\[3\] 0.003415f
C15903 net20 _317_/a_36_113# 0.00189f
C15904 _115_ _122_ 0.004082f
C15905 net34 FILLER_0_22_177/a_484_472# 0.003953f
C15906 _020_ _142_ 0.010094f
C15907 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1468_375# 0.016748f
C15908 net76 net18 0.002264f
C15909 _076_ _125_ 0.009254f
C15910 net55 vss 0.947665f
C15911 net68 FILLER_0_8_37/a_484_472# 0.002696f
C15912 fanout49/a_36_160# FILLER_0_5_88/a_124_375# 0.001154f
C15913 _188_ _453_/a_36_151# 0.03354f
C15914 _407_/a_36_472# _184_ 0.004667f
C15915 _095_ _451_/a_448_472# 0.002474f
C15916 net42 net40 0.007686f
C15917 _005_ _094_ 0.162984f
C15918 _074_ _251_/a_906_472# 0.002887f
C15919 _144_ _141_ 0.095441f
C15920 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_572_375# 0.007947f
C15921 _063_ _445_/a_2248_156# 0.008121f
C15922 net17 _054_ 0.034759f
C15923 _115_ _227_/a_36_160# 0.00124f
C15924 ctlp[2] _299_/a_36_472# 0.012937f
C15925 _131_ _043_ 0.047425f
C15926 _053_ _385_/a_36_68# 0.018437f
C15927 FILLER_0_17_72/a_932_472# net36 0.00356f
C15928 FILLER_0_7_104/a_1380_472# _154_ 0.002799f
C15929 _359_/a_36_488# net74 0.037211f
C15930 _137_ _334_/a_36_160# 0.015722f
C15931 _442_/a_3041_156# vdd 0.001178f
C15932 mask\[9\] _438_/a_796_472# 0.004751f
C15933 FILLER_0_15_150/a_36_472# _095_ 0.001526f
C15934 net27 FILLER_0_12_236/a_124_375# 0.044776f
C15935 FILLER_0_5_164/a_572_375# vss 0.055055f
C15936 FILLER_0_5_164/a_36_472# vdd 0.004144f
C15937 net58 FILLER_0_9_270/a_572_375# 0.006256f
C15938 _126_ FILLER_0_11_124/a_124_375# 0.038971f
C15939 output13/a_224_472# net13 0.058196f
C15940 _030_ _154_ 0.004803f
C15941 output11/a_224_472# _411_/a_36_151# 0.095813f
C15942 _376_/a_36_160# trim_mask\[1\] 0.003111f
C15943 _091_ _430_/a_1308_423# 0.023198f
C15944 net50 trim_val\[0\] 0.390586f
C15945 net52 _442_/a_36_151# 0.029373f
C15946 ctln[1] _411_/a_2665_112# 0.004748f
C15947 FILLER_0_18_177/a_3260_375# vss 0.055219f
C15948 FILLER_0_18_177/a_36_472# vdd 0.110153f
C15949 _431_/a_448_472# vdd 0.001932f
C15950 output8/a_224_472# FILLER_0_3_221/a_1020_375# 0.03228f
C15951 net72 _174_ 0.199504f
C15952 _339_/a_36_160# FILLER_0_19_155/a_572_375# 0.003589f
C15953 net66 FILLER_0_5_54/a_572_375# 0.002203f
C15954 _450_/a_3129_107# _039_ 0.012762f
C15955 FILLER_0_11_101/a_484_472# cal_count\[3\] 0.00702f
C15956 net18 _419_/a_1308_423# 0.013637f
C15957 _095_ _185_ 0.034457f
C15958 net69 _168_ 0.035976f
C15959 _439_/a_36_151# FILLER_0_6_47/a_2364_375# 0.002807f
C15960 output27/a_224_472# _425_/a_2665_112# 0.021504f
C15961 net16 FILLER_0_18_37/a_484_472# 0.054878f
C15962 _091_ _430_/a_1204_472# 0.007301f
C15963 net17 vss 0.940703f
C15964 net69 _441_/a_796_472# 0.002057f
C15965 FILLER_0_21_142/a_36_472# vdd 0.111749f
C15966 FILLER_0_17_104/a_124_375# net14 0.010099f
C15967 _178_ net17 0.115251f
C15968 _141_ net23 0.782974f
C15969 _429_/a_36_151# _043_ 0.002771f
C15970 _072_ cal_count\[3\] 0.028346f
C15971 trim_val\[1\] vss 0.029927f
C15972 _431_/a_2248_156# net56 0.013627f
C15973 FILLER_0_16_73/a_484_472# FILLER_0_15_72/a_484_472# 0.026657f
C15974 _140_ _436_/a_36_151# 0.031519f
C15975 _425_/a_1308_423# vdd 0.021703f
C15976 FILLER_0_17_282/a_36_472# _418_/a_448_472# 0.011962f
C15977 net17 FILLER_0_20_15/a_932_472# 0.047256f
C15978 net37 FILLER_0_6_231/a_124_375# 0.001989f
C15979 mask\[7\] FILLER_0_22_128/a_36_472# 0.013408f
C15980 FILLER_0_17_282/a_124_375# _006_ 0.004694f
C15981 _114_ _055_ 0.071738f
C15982 _028_ FILLER_0_7_72/a_2812_375# 0.003873f
C15983 net4 _060_ 0.327437f
C15984 _057_ cal_itt\[3\] 0.014849f
C15985 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1468_375# 0.086635f
C15986 state\[2\] _427_/a_448_472# 0.00237f
C15987 net53 _427_/a_796_472# 0.001983f
C15988 net64 FILLER_0_9_270/a_124_375# 0.013532f
C15989 _067_ FILLER_0_12_20/a_124_375# 0.017026f
C15990 _082_ vss 0.053349f
C15991 result[0] net65 0.011634f
C15992 _144_ _148_ 0.038002f
C15993 FILLER_0_18_76/a_572_375# _438_/a_36_151# 0.059049f
C15994 net82 vss 0.550252f
C15995 _428_/a_448_472# net74 0.019814f
C15996 net61 ctlp[1] 2.770871f
C15997 net52 _439_/a_1000_472# 0.03537f
C15998 net50 _439_/a_1308_423# 0.008832f
C15999 _445_/a_2560_156# net49 0.001208f
C16000 net3 FILLER_0_15_10/a_124_375# 0.035504f
C16001 FILLER_0_4_49/a_124_375# vdd 0.008637f
C16002 _126_ _428_/a_2248_156# 0.001131f
C16003 _098_ FILLER_0_16_154/a_1020_375# 0.003386f
C16004 fanout57/a_36_113# vss 0.046378f
C16005 FILLER_0_12_136/a_124_375# net57 0.001727f
C16006 output23/a_224_472# net23 0.122379f
C16007 _432_/a_448_472# vdd 0.035246f
C16008 fanout54/a_36_160# FILLER_0_19_142/a_124_375# 0.005489f
C16009 output38/a_224_472# net40 0.072234f
C16010 _028_ _151_ 0.020076f
C16011 _106_ _093_ 0.045972f
C16012 _013_ FILLER_0_18_53/a_36_472# 0.013138f
C16013 _428_/a_2665_112# _095_ 0.001471f
C16014 fanout53/a_36_160# _095_ 0.007436f
C16015 _114_ _255_/a_224_552# 0.005131f
C16016 output43/a_224_472# net17 0.083607f
C16017 _043_ FILLER_0_13_80/a_36_472# 0.016194f
C16018 _136_ _337_/a_49_472# 0.058704f
C16019 _114_ _126_ 3.341247f
C16020 FILLER_0_5_54/a_124_375# FILLER_0_3_54/a_36_472# 0.001512f
C16021 _015_ FILLER_0_8_247/a_36_472# 0.005458f
C16022 _091_ _097_ 0.036863f
C16023 FILLER_0_3_78/a_484_472# vss 0.005811f
C16024 _176_ FILLER_0_10_107/a_124_375# 0.013408f
C16025 _132_ FILLER_0_14_107/a_1468_375# 0.019517f
C16026 FILLER_0_22_86/a_572_375# vdd 0.017472f
C16027 FILLER_0_22_86/a_124_375# vss 0.00285f
C16028 FILLER_0_11_78/a_124_375# _120_ 0.014367f
C16029 net63 FILLER_0_18_177/a_932_472# 0.063742f
C16030 net68 fanout68/a_36_113# 0.027807f
C16031 FILLER_0_22_128/a_1380_472# vdd 0.005746f
C16032 FILLER_0_22_128/a_932_472# vss 0.003452f
C16033 _058_ trim_mask\[0\] 0.076069f
C16034 net35 _146_ 0.096468f
C16035 _216_/a_67_603# vss 0.012211f
C16036 _095_ cal_count\[0\] 0.005211f
C16037 _074_ net76 0.026801f
C16038 net27 _426_/a_1000_472# 0.002971f
C16039 _086_ _125_ 0.490983f
C16040 mask\[5\] FILLER_0_19_187/a_572_375# 0.005529f
C16041 ctln[8] FILLER_0_0_96/a_124_375# 0.002726f
C16042 _116_ net4 0.00603f
C16043 _056_ _226_/a_1044_68# 0.002852f
C16044 net56 FILLER_0_18_139/a_1468_375# 0.065206f
C16045 _091_ _430_/a_448_472# 0.065306f
C16046 net80 _139_ 0.178583f
C16047 net27 FILLER_0_9_290/a_124_375# 0.002657f
C16048 _121_ vdd 0.106437f
C16049 fanout78/a_36_113# vdd 0.061637f
C16050 _415_/a_36_151# net81 0.046145f
C16051 _088_ FILLER_0_3_172/a_3172_472# 0.004381f
C16052 net31 net30 0.130396f
C16053 _425_/a_1000_472# net19 0.020388f
C16054 _111_ vss 0.233815f
C16055 net41 _217_/a_36_160# 0.004517f
C16056 _053_ FILLER_0_6_47/a_2812_375# 0.003818f
C16057 net46 net17 0.791341f
C16058 _445_/a_36_151# _034_ 0.005488f
C16059 FILLER_0_4_177/a_36_472# net37 0.004017f
C16060 _119_ _070_ 1.949038f
C16061 net64 FILLER_0_11_282/a_36_472# 0.003938f
C16062 net76 _076_ 0.003124f
C16063 _185_ _402_/a_1296_93# 0.001714f
C16064 _070_ _071_ 0.001757f
C16065 FILLER_0_14_50/a_124_375# _401_/a_36_68# 0.001129f
C16066 net82 FILLER_0_3_172/a_3260_375# 0.007693f
C16067 FILLER_0_5_54/a_124_375# _164_ 0.004076f
C16068 output35/a_224_472# _048_ 0.009509f
C16069 _095_ _098_ 0.057687f
C16070 _093_ FILLER_0_18_107/a_36_472# 0.008683f
C16071 net57 net14 0.05113f
C16072 trim_mask\[2\] _447_/a_36_151# 0.022881f
C16073 _093_ _302_/a_224_472# 0.011376f
C16074 _091_ mask\[2\] 2.252217f
C16075 FILLER_0_3_172/a_2364_375# net65 0.003745f
C16076 _128_ _085_ 0.004532f
C16077 net57 fanout55/a_36_160# 0.017476f
C16078 FILLER_0_4_177/a_572_375# _087_ 0.006527f
C16079 _046_ vdd 0.041841f
C16080 net48 _112_ 0.284235f
C16081 _277_/a_36_160# _093_ 0.018101f
C16082 net82 fanout76/a_36_160# 0.001033f
C16083 _155_ vdd 0.193832f
C16084 FILLER_0_9_28/a_572_375# vdd 0.023246f
C16085 _316_/a_848_380# _123_ 0.0018f
C16086 _443_/a_36_151# vdd 0.175472f
C16087 FILLER_0_15_116/a_36_472# vdd 0.013454f
C16088 _104_ FILLER_0_17_226/a_36_472# 0.013926f
C16089 FILLER_0_4_197/a_36_472# net21 0.011079f
C16090 net20 _046_ 0.194455f
C16091 net81 _136_ 0.021146f
C16092 _409_/a_245_68# cal_count\[3\] 0.001164f
C16093 _448_/a_796_472# vdd 0.002153f
C16094 _439_/a_2248_156# net14 0.001279f
C16095 _028_ FILLER_0_5_72/a_932_472# 0.003042f
C16096 net22 net59 0.195226f
C16097 net68 _220_/a_67_603# 0.030878f
C16098 _149_ FILLER_0_20_98/a_124_375# 0.020028f
C16099 net81 net62 0.245647f
C16100 FILLER_0_13_228/a_124_375# FILLER_0_12_220/a_1020_375# 0.05841f
C16101 FILLER_0_21_142/a_484_472# mask\[7\] 0.001603f
C16102 FILLER_0_16_57/a_124_375# net72 0.052543f
C16103 net15 FILLER_0_17_56/a_572_375# 0.007386f
C16104 FILLER_0_7_59/a_36_472# net68 0.050931f
C16105 FILLER_0_5_54/a_1020_375# net47 0.005159f
C16106 _414_/a_1000_472# cal_itt\[3\] 0.08528f
C16107 net26 FILLER_0_21_28/a_2276_472# 0.001561f
C16108 net57 _428_/a_36_151# 0.023215f
C16109 net32 output19/a_224_472# 0.101682f
C16110 _433_/a_2248_156# _145_ 0.009108f
C16111 net75 FILLER_0_0_232/a_36_472# 0.001514f
C16112 _184_ net17 0.007958f
C16113 _073_ _260_/a_36_68# 0.079772f
C16114 _376_/a_36_160# FILLER_0_6_90/a_36_472# 0.195478f
C16115 _043_ FILLER_0_15_180/a_36_472# 0.001219f
C16116 FILLER_0_24_130/a_124_375# output24/a_224_472# 0.00515f
C16117 FILLER_0_16_107/a_124_375# vss 0.002683f
C16118 _132_ vdd 0.960634f
C16119 ctln[6] _442_/a_36_151# 0.007031f
C16120 FILLER_0_24_130/a_124_375# vss 0.018125f
C16121 _003_ _414_/a_36_151# 0.021191f
C16122 FILLER_0_7_195/a_36_472# calibrate 0.010951f
C16123 FILLER_0_17_72/a_2364_375# vdd 0.002455f
C16124 FILLER_0_17_72/a_1916_375# vss 0.001345f
C16125 FILLER_0_12_20/a_572_375# net47 0.00139f
C16126 net55 _027_ 0.002104f
C16127 ctlp[2] vss 0.131085f
C16128 net73 FILLER_0_18_107/a_3172_472# 0.00533f
C16129 _412_/a_36_151# net81 0.014094f
C16130 FILLER_0_4_107/a_36_472# vss 0.002634f
C16131 FILLER_0_2_111/a_932_472# _158_ 0.00264f
C16132 FILLER_0_4_107/a_484_472# vdd 0.03151f
C16133 _000_ _411_/a_448_472# 0.073053f
C16134 FILLER_0_5_72/a_36_472# FILLER_0_6_47/a_2812_375# 0.001597f
C16135 _073_ net4 0.076114f
C16136 _427_/a_36_151# vdd 0.107344f
C16137 FILLER_0_7_195/a_36_472# net21 0.005469f
C16138 net72 FILLER_0_15_59/a_124_375# 0.022905f
C16139 _122_ net22 0.024638f
C16140 _043_ FILLER_0_13_72/a_124_375# 0.013517f
C16141 _424_/a_2248_156# FILLER_0_21_60/a_572_375# 0.030666f
C16142 _424_/a_2665_112# FILLER_0_21_60/a_124_375# 0.010688f
C16143 FILLER_0_12_220/a_124_375# _070_ 0.007554f
C16144 _363_/a_36_68# _163_ 0.005627f
C16145 trim_val\[2\] _167_ 0.011787f
C16146 trim_mask\[2\] FILLER_0_2_93/a_124_375# 0.046032f
C16147 net76 _081_ 0.706096f
C16148 mask\[3\] FILLER_0_16_241/a_124_375# 0.006824f
C16149 _091_ FILLER_0_15_212/a_572_375# 0.022582f
C16150 net60 _421_/a_2248_156# 0.036944f
C16151 mask\[3\] FILLER_0_18_177/a_1020_375# 0.002924f
C16152 _321_/a_170_472# vdd 0.060585f
C16153 en_co_clk _043_ 0.041355f
C16154 FILLER_0_14_50/a_124_375# _095_ 0.052375f
C16155 _179_ _180_ 0.018662f
C16156 _130_ _126_ 0.061836f
C16157 _155_ FILLER_0_5_109/a_36_472# 0.001872f
C16158 _144_ _207_/a_67_603# 0.064623f
C16159 FILLER_0_8_107/a_124_375# vdd 0.049132f
C16160 _114_ state\[1\] 0.087216f
C16161 _018_ net21 0.077174f
C16162 net79 _044_ 0.013636f
C16163 FILLER_0_18_2/a_3172_472# FILLER_0_18_37/a_36_472# 0.002765f
C16164 net81 _429_/a_2665_112# 0.012675f
C16165 FILLER_0_11_142/a_36_472# _120_ 0.040786f
C16166 _408_/a_1336_472# vss 0.001022f
C16167 _408_/a_728_93# vdd 0.024163f
C16168 _141_ FILLER_0_19_155/a_484_472# 0.015625f
C16169 _086_ net76 0.049988f
C16170 FILLER_0_13_142/a_1380_472# vdd 0.001977f
C16171 FILLER_0_13_142/a_932_472# vss 0.005192f
C16172 net49 _440_/a_796_472# 0.003597f
C16173 _128_ _062_ 0.025708f
C16174 mask\[7\] _299_/a_36_472# 0.033949f
C16175 net50 FILLER_0_5_72/a_1380_472# 0.002431f
C16176 _363_/a_244_472# _028_ 0.002693f
C16177 FILLER_0_7_59/a_36_472# net67 0.021549f
C16178 net38 FILLER_0_15_2/a_572_375# 0.007477f
C16179 _235_/a_255_603# trim_mask\[2\] 0.001488f
C16180 _235_/a_67_603# trim_val\[2\] 0.00747f
C16181 net55 _095_ 0.055644f
C16182 _143_ vdd 0.074199f
C16183 FILLER_0_11_142/a_484_472# FILLER_0_13_142/a_572_375# 0.0027f
C16184 _431_/a_796_472# net70 0.001754f
C16185 net76 net65 0.14935f
C16186 _062_ _311_/a_692_473# 0.008632f
C16187 _447_/a_796_472# vdd 0.001959f
C16188 FILLER_0_5_117/a_124_375# FILLER_0_4_107/a_1380_472# 0.001684f
C16189 net57 FILLER_0_8_156/a_124_375# 0.001628f
C16190 net24 FILLER_0_22_107/a_124_375# 0.001023f
C16191 net15 FILLER_0_9_72/a_36_472# 0.006905f
C16192 _356_/a_36_472# vdd 0.016338f
C16193 result[4] vdd 0.205815f
C16194 result[2] net18 0.086474f
C16195 FILLER_0_11_64/a_124_375# _453_/a_36_151# 0.005577f
C16196 _256_/a_2124_68# _070_ 0.002444f
C16197 net23 FILLER_0_22_128/a_1468_375# 0.001866f
C16198 net54 _352_/a_49_472# 0.003941f
C16199 net59 vdd 2.180407f
C16200 _137_ FILLER_0_16_154/a_1468_375# 0.014214f
C16201 net23 _207_/a_67_603# 0.002734f
C16202 _341_/a_49_472# _137_ 0.059288f
C16203 _315_/a_716_497# net23 0.004725f
C16204 fanout72/a_36_113# _067_ 0.005796f
C16205 net54 _433_/a_1000_472# 0.0025f
C16206 FILLER_0_0_198/a_124_375# vdd 0.04491f
C16207 output37/a_224_472# fanout64/a_36_160# 0.017421f
C16208 _075_ vss 0.046342f
C16209 _132_ _135_ 0.345161f
C16210 mask\[4\] FILLER_0_18_177/a_3172_472# 0.014657f
C16211 _450_/a_2449_156# net40 0.010265f
C16212 net15 _453_/a_2248_156# 0.044493f
C16213 net32 mask\[6\] 0.003248f
C16214 net20 result[4] 0.001673f
C16215 FILLER_0_8_127/a_124_375# _133_ 0.001928f
C16216 FILLER_0_21_125/a_124_375# _433_/a_36_151# 0.059049f
C16217 result[7] _420_/a_2560_156# 0.001179f
C16218 net20 net59 0.045227f
C16219 _214_/a_36_160# _213_/a_67_603# 0.002505f
C16220 net41 output40/a_224_472# 0.018977f
C16221 _095_ net17 0.172789f
C16222 vdd FILLER_0_10_94/a_484_472# 0.008627f
C16223 _444_/a_1308_423# _054_ 0.005457f
C16224 net58 vss 0.589419f
C16225 _077_ net48 0.142015f
C16226 FILLER_0_20_107/a_124_375# FILLER_0_20_98/a_124_375# 0.003228f
C16227 output33/a_224_472# _204_/a_67_603# 0.00401f
C16228 _146_ vdd 0.031209f
C16229 FILLER_0_14_81/a_36_472# FILLER_0_13_80/a_124_375# 0.001597f
C16230 FILLER_0_18_2/a_1828_472# _452_/a_448_472# 0.005748f
C16231 net82 FILLER_0_2_177/a_36_472# 0.001777f
C16232 result[8] FILLER_0_24_290/a_124_375# 0.00562f
C16233 FILLER_0_4_197/a_1380_472# net22 0.012286f
C16234 fanout59/a_36_160# net5 0.05829f
C16235 _035_ net47 0.101683f
C16236 FILLER_0_8_24/a_572_375# _054_ 0.004858f
C16237 _261_/a_36_160# FILLER_0_5_136/a_36_472# 0.00304f
C16238 cal_count\[1\] FILLER_0_15_59/a_572_375# 0.008797f
C16239 _093_ _012_ 0.141641f
C16240 FILLER_0_7_72/a_2364_375# FILLER_0_6_90/a_484_472# 0.001684f
C16241 net81 net4 0.003327f
C16242 _412_/a_1204_472# net65 0.001629f
C16243 _412_/a_2248_156# vdd 0.005671f
C16244 FILLER_0_0_130/a_124_375# _031_ 0.001861f
C16245 state\[0\] FILLER_0_12_220/a_1380_472# 0.003733f
C16246 net65 FILLER_0_2_177/a_124_375# 0.018094f
C16247 _036_ net17 0.153479f
C16248 _058_ _118_ 0.001451f
C16249 _449_/a_1000_472# net72 0.001247f
C16250 _449_/a_448_472# net55 0.004439f
C16251 output26/a_224_472# net17 0.004277f
C16252 _025_ _436_/a_1000_472# 0.061189f
C16253 _000_ _074_ 0.003542f
C16254 _070_ _385_/a_36_68# 0.049178f
C16255 _422_/a_36_151# _109_ 0.036674f
C16256 FILLER_0_5_206/a_124_375# net22 0.019537f
C16257 calibrate vss 1.140031f
C16258 _122_ vdd 0.379907f
C16259 _110_ net36 0.002287f
C16260 _412_/a_36_151# net2 0.003823f
C16261 fanout54/a_36_160# vss 0.061573f
C16262 net64 FILLER_0_15_235/a_572_375# 0.007219f
C16263 FILLER_0_16_37/a_36_472# vdd 0.142203f
C16264 FILLER_0_16_37/a_124_375# vss 0.021237f
C16265 _178_ FILLER_0_16_37/a_124_375# 0.036901f
C16266 FILLER_0_7_233/a_124_375# vdd 0.03915f
C16267 _044_ FILLER_0_13_290/a_124_375# 0.001855f
C16268 FILLER_0_10_256/a_124_375# vss 0.006036f
C16269 FILLER_0_10_256/a_36_472# vdd 0.025204f
C16270 FILLER_0_2_111/a_36_472# trim_mask\[3\] 0.007915f
C16271 FILLER_0_8_127/a_36_472# _322_/a_124_24# 0.00171f
C16272 _421_/a_36_151# net18 0.00659f
C16273 FILLER_0_8_24/a_572_375# vss 0.012859f
C16274 FILLER_0_8_24/a_36_472# vdd 0.007423f
C16275 _274_/a_1612_497# net20 0.002057f
C16276 _227_/a_36_160# vdd 0.007828f
C16277 net64 vdd 1.155692f
C16278 net20 _122_ 0.046817f
C16279 _453_/a_2248_156# net51 0.05329f
C16280 _120_ _172_ 0.010275f
C16281 _038_ _172_ 0.050158f
C16282 net21 vss 1.123312f
C16283 net35 FILLER_0_23_88/a_124_375# 0.009071f
C16284 result[8] FILLER_0_24_274/a_1380_472# 0.005458f
C16285 fanout51/a_36_113# FILLER_0_11_64/a_124_375# 0.002335f
C16286 net62 _045_ 0.029263f
C16287 _333_/a_36_160# vss 0.030799f
C16288 _169_ vdd 0.055642f
C16289 net38 _452_/a_448_472# 0.016895f
C16290 FILLER_0_4_49/a_572_375# net68 0.023227f
C16291 net20 FILLER_0_7_233/a_124_375# 0.017217f
C16292 mask\[3\] _198_/a_67_603# 0.024102f
C16293 net70 FILLER_0_18_107/a_1380_472# 0.00116f
C16294 FILLER_0_2_93/a_484_472# vdd 0.005163f
C16295 _072_ _267_/a_224_472# 0.004269f
C16296 _438_/a_1308_423# net14 0.005201f
C16297 FILLER_0_0_96/a_124_375# net14 0.077876f
C16298 FILLER_0_19_171/a_1380_472# vdd 0.03086f
C16299 FILLER_0_19_171/a_932_472# vss 0.001256f
C16300 net20 net64 0.374636f
C16301 _432_/a_1204_472# _137_ 0.006554f
C16302 _063_ _232_/a_67_603# 0.005404f
C16303 FILLER_0_14_91/a_124_375# en_co_clk 0.006788f
C16304 _069_ _121_ 0.137961f
C16305 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_124_375# 0.004426f
C16306 net23 FILLER_0_5_148/a_36_472# 0.011079f
C16307 FILLER_0_15_72/a_572_375# _451_/a_3129_107# 0.007026f
C16308 FILLER_0_21_133/a_36_472# _433_/a_36_151# 0.001723f
C16309 net44 _452_/a_2225_156# 0.044858f
C16310 _402_/a_728_93# _182_ 0.00263f
C16311 trim_val\[2\] vdd 0.160419f
C16312 trim_mask\[2\] vss 0.182675f
C16313 net47 FILLER_0_5_148/a_484_472# 0.009741f
C16314 net58 fanout76/a_36_160# 0.055026f
C16315 net17 output41/a_224_472# 0.030456f
C16316 FILLER_0_22_86/a_1020_375# _026_ 0.001032f
C16317 _253_/a_36_68# _084_ 0.029805f
C16318 _430_/a_1308_423# net22 0.035518f
C16319 FILLER_0_2_165/a_124_375# net59 0.00999f
C16320 _230_/a_652_68# _062_ 0.001144f
C16321 FILLER_0_23_44/a_36_472# vdd 0.01833f
C16322 FILLER_0_23_44/a_1468_375# vss 0.055902f
C16323 _053_ FILLER_0_7_59/a_124_375# 0.015298f
C16324 net15 _441_/a_1308_423# 0.009697f
C16325 _173_ FILLER_0_12_28/a_124_375# 0.009218f
C16326 _408_/a_1336_472# _184_ 0.003286f
C16327 _430_/a_1204_472# net22 0.028536f
C16328 _440_/a_2665_112# net47 0.014066f
C16329 _018_ mask\[1\] 0.001206f
C16330 _412_/a_36_151# valid 0.009757f
C16331 _418_/a_448_472# vss 0.005772f
C16332 _418_/a_1308_423# vdd 0.002258f
C16333 net80 _023_ 0.261119f
C16334 _006_ vdd 0.632993f
C16335 FILLER_0_14_107/a_1380_472# vdd 0.002511f
C16336 _112_ net37 0.070289f
C16337 _057_ _306_/a_36_68# 0.019072f
C16338 FILLER_0_3_172/a_3260_375# net21 0.049606f
C16339 clk vss 0.210484f
C16340 output12/a_224_472# _037_ 0.00827f
C16341 _056_ FILLER_0_12_196/a_36_472# 0.039555f
C16342 FILLER_0_22_177/a_36_472# net33 0.013661f
C16343 _433_/a_796_472# _022_ 0.025882f
C16344 FILLER_0_4_197/a_1380_472# vdd 0.00581f
C16345 fanout66/a_36_113# net49 0.001044f
C16346 cal_itt\[3\] _161_ 0.20195f
C16347 fanout65/a_36_113# net65 0.019148f
C16348 _259_/a_455_68# _076_ 0.002372f
C16349 _043_ _090_ 0.001578f
C16350 FILLER_0_21_286/a_572_375# vss 0.031895f
C16351 FILLER_0_21_286/a_36_472# vdd 0.008714f
C16352 FILLER_0_16_255/a_36_472# net30 0.00209f
C16353 mask\[3\] _430_/a_36_151# 0.005848f
C16354 FILLER_0_15_116/a_572_375# _095_ 0.00152f
C16355 net52 FILLER_0_9_72/a_124_375# 0.029702f
C16356 _256_/a_36_68# vss 0.055568f
C16357 _103_ vdd 0.590261f
C16358 net36 net14 0.037175f
C16359 mask\[5\] FILLER_0_20_169/a_36_472# 0.016469f
C16360 FILLER_0_21_28/a_1380_472# net17 0.001709f
C16361 net20 _256_/a_716_497# 0.007413f
C16362 net20 _006_ 0.014721f
C16363 FILLER_0_1_266/a_124_375# vdd -0.002281f
C16364 _021_ _432_/a_796_472# 0.001666f
C16365 net34 _023_ 0.00872f
C16366 FILLER_0_16_89/a_124_375# _176_ 0.002781f
C16367 fanout81/a_36_160# vss 0.02458f
C16368 FILLER_0_5_206/a_124_375# vdd 0.038311f
C16369 _053_ _070_ 2.345795f
C16370 FILLER_0_15_150/a_36_472# fanout53/a_36_160# 0.002059f
C16371 ctln[4] net65 0.020799f
C16372 net2 net4 0.854661f
C16373 _274_/a_2552_68# _070_ 0.001238f
C16374 net50 FILLER_0_7_59/a_484_472# 0.011974f
C16375 FILLER_0_16_107/a_484_472# net14 0.001528f
C16376 _144_ _348_/a_257_69# 0.001978f
C16377 FILLER_0_18_2/a_3260_375# vss 0.026159f
C16378 FILLER_0_18_2/a_36_472# vdd 0.104532f
C16379 net20 _103_ 0.261438f
C16380 _053_ FILLER_0_7_146/a_36_472# 0.001014f
C16381 _141_ _340_/a_36_160# 0.00584f
C16382 FILLER_0_18_61/a_124_375# vss 0.021307f
C16383 FILLER_0_18_61/a_36_472# vdd 0.08828f
C16384 ctlp[3] _296_/a_224_472# 0.005335f
C16385 _428_/a_1204_472# _131_ 0.012968f
C16386 FILLER_0_18_2/a_2812_375# FILLER_0_20_15/a_1380_472# 0.001338f
C16387 mask\[7\] vss 0.85153f
C16388 FILLER_0_3_204/a_124_375# _088_ 0.00269f
C16389 _325_/a_224_472# _120_ 0.00233f
C16390 mask\[5\] FILLER_0_18_177/a_1380_472# 0.001063f
C16391 net26 FILLER_0_18_37/a_572_375# 0.00109f
C16392 output46/a_224_472# FILLER_0_21_28/a_124_375# 0.003337f
C16393 FILLER_0_4_213/a_36_472# FILLER_0_3_212/a_124_375# 0.001597f
C16394 vdd FILLER_0_4_91/a_572_375# 0.019853f
C16395 _074_ FILLER_0_6_231/a_36_472# 0.004325f
C16396 net31 _046_ 0.008368f
C16397 _098_ FILLER_0_20_87/a_124_375# 0.019333f
C16398 cal_count\[3\] FILLER_0_11_78/a_484_472# 0.011737f
C16399 ctlp[1] FILLER_0_24_274/a_1468_375# 0.01305f
C16400 FILLER_0_3_172/a_932_472# net22 0.012284f
C16401 _427_/a_448_472# _043_ 0.002896f
C16402 FILLER_0_5_128/a_124_375# _370_/a_124_24# 0.023285f
C16403 _422_/a_1000_472# mask\[7\] 0.039617f
C16404 _016_ fanout73/a_36_113# 0.001731f
C16405 FILLER_0_16_73/a_484_472# FILLER_0_17_72/a_572_375# 0.001723f
C16406 _000_ net65 0.093773f
C16407 _086_ _267_/a_1568_472# 0.002143f
C16408 FILLER_0_18_177/a_1468_375# _139_ 0.001359f
C16409 output36/a_224_472# output30/a_224_472# 0.003578f
C16410 _076_ FILLER_0_6_231/a_36_472# 0.005517f
C16411 _407_/a_36_472# _185_ 0.009281f
C16412 _085_ _176_ 0.024708f
C16413 _185_ cal_count\[0\] 0.008096f
C16414 output30/a_224_472# net30 0.043557f
C16415 _430_/a_448_472# net22 0.036303f
C16416 _096_ _335_/a_257_69# 0.001084f
C16417 FILLER_0_18_107/a_2812_375# FILLER_0_17_133/a_36_472# 0.001543f
C16418 ctln[3] _411_/a_1000_472# 0.00283f
C16419 net74 _136_ 0.042043f
C16420 net75 FILLER_0_8_247/a_1468_375# 0.047331f
C16421 net16 _408_/a_1936_472# 0.022235f
C16422 _321_/a_170_472# _069_ 0.025551f
C16423 _408_/a_56_524# _043_ 0.10151f
C16424 _430_/a_1308_423# vdd 0.00218f
C16425 net7 _064_ 0.001538f
C16426 FILLER_0_12_136/a_36_472# FILLER_0_11_135/a_124_375# 0.001597f
C16427 _436_/a_2665_112# FILLER_0_22_128/a_1020_375# 0.029834f
C16428 FILLER_0_15_235/a_36_472# mask\[1\] 0.009316f
C16429 _093_ FILLER_0_19_155/a_36_472# 0.001737f
C16430 result[8] FILLER_0_23_282/a_36_472# 0.001908f
C16431 net74 FILLER_0_13_142/a_124_375# 0.002722f
C16432 FILLER_0_5_198/a_572_375# net59 0.00183f
C16433 _432_/a_1000_472# _137_ 0.008914f
C16434 FILLER_0_1_266/a_36_472# net19 0.07227f
C16435 FILLER_0_5_54/a_36_472# FILLER_0_6_47/a_932_472# 0.026657f
C16436 FILLER_0_5_54/a_1020_375# FILLER_0_6_47/a_1828_472# 0.001597f
C16437 mask\[7\] _107_ 0.13732f
C16438 _345_/a_36_160# _098_ 0.002041f
C16439 FILLER_0_17_200/a_36_472# _430_/a_36_151# 0.001723f
C16440 _428_/a_448_472# net70 0.007116f
C16441 mask\[2\] net22 0.034216f
C16442 net68 _029_ 0.094915f
C16443 FILLER_0_16_57/a_36_472# FILLER_0_17_56/a_124_375# 0.001723f
C16444 _016_ net57 0.028276f
C16445 _369_/a_244_472# vdd 0.001255f
C16446 mask\[1\] vss 0.46268f
C16447 _414_/a_36_151# net76 0.037157f
C16448 _192_/a_255_603# mask\[1\] 0.001059f
C16449 net36 FILLER_0_15_212/a_932_472# 0.008239f
C16450 _408_/a_1336_472# _095_ 0.011305f
C16451 _028_ _086_ 0.011526f
C16452 _119_ calibrate 0.062309f
C16453 _095_ FILLER_0_13_142/a_932_472# 0.001782f
C16454 fanout81/a_36_160# fanout76/a_36_160# 0.01081f
C16455 FILLER_0_2_177/a_572_375# net59 0.005397f
C16456 FILLER_0_11_142/a_124_375# vss 0.008766f
C16457 FILLER_0_11_142/a_572_375# vdd 0.014107f
C16458 _188_ _042_ 0.015684f
C16459 FILLER_0_12_136/a_484_472# _076_ 0.001683f
C16460 net80 FILLER_0_20_169/a_36_472# 0.024142f
C16461 _141_ _348_/a_49_472# 0.037821f
C16462 _079_ _084_ 0.046584f
C16463 _322_/a_848_380# _129_ 0.048486f
C16464 FILLER_0_18_107/a_2364_375# vdd 0.017472f
C16465 FILLER_0_7_72/a_1020_375# FILLER_0_5_72/a_932_472# 0.001512f
C16466 _434_/a_36_151# mask\[6\] 0.048644f
C16467 net24 FILLER_0_22_86/a_1468_375# 0.008075f
C16468 trim_mask\[4\] _386_/a_124_24# 0.040347f
C16469 _422_/a_2248_156# vss 0.001755f
C16470 _422_/a_2665_112# vdd 0.008306f
C16471 FILLER_0_7_104/a_572_375# vdd 0.038253f
C16472 FILLER_0_18_139/a_1468_375# _145_ 0.002318f
C16473 FILLER_0_7_72/a_2364_375# net14 0.005919f
C16474 net79 FILLER_0_12_220/a_484_472# 0.005464f
C16475 _441_/a_2560_156# vss 0.001374f
C16476 net47 _386_/a_124_24# 0.024696f
C16477 _053_ trim_val\[1\] 0.00385f
C16478 _029_ _156_ 0.018258f
C16479 _074_ _375_/a_1388_497# 0.005488f
C16480 net55 _424_/a_2560_156# 0.003707f
C16481 net48 net1 0.006424f
C16482 FILLER_0_7_162/a_124_375# vdd 0.011809f
C16483 fanout78/a_36_113# net77 0.036366f
C16484 _174_ vdd 0.18623f
C16485 mask\[0\] _018_ 0.328328f
C16486 _447_/a_1000_472# net68 0.006223f
C16487 _447_/a_1308_423# _036_ 0.003079f
C16488 net50 net69 0.634381f
C16489 net52 _031_ 0.633473f
C16490 FILLER_0_23_88/a_124_375# vdd 0.03583f
C16491 _093_ _177_ 0.001194f
C16492 ctln[3] net10 0.873575f
C16493 _033_ FILLER_0_6_47/a_36_472# 0.001185f
C16494 trimb[1] net40 0.00126f
C16495 net24 _211_/a_36_160# 0.021941f
C16496 FILLER_0_12_124/a_124_375# _428_/a_36_151# 0.058722f
C16497 input2/a_36_113# vss 0.055539f
C16498 _122_ FILLER_0_5_198/a_572_375# 0.001352f
C16499 net47 _452_/a_1353_112# 0.003681f
C16500 _126_ FILLER_0_10_94/a_572_375# 0.027249f
C16501 _208_/a_36_160# FILLER_0_22_128/a_3260_375# 0.001948f
C16502 _417_/a_36_151# output30/a_224_472# 0.004902f
C16503 _131_ FILLER_0_17_104/a_932_472# 0.002988f
C16504 _062_ _226_/a_276_68# 0.001286f
C16505 _091_ FILLER_0_13_212/a_1020_375# 0.00799f
C16506 _441_/a_448_472# net66 0.023761f
C16507 FILLER_0_21_142/a_36_472# _140_ 0.009261f
C16508 _097_ vdd 0.191424f
C16509 _437_/a_448_472# vss 0.001524f
C16510 _437_/a_1308_423# vdd 0.005139f
C16511 _077_ net37 0.003374f
C16512 cal_itt\[3\] _056_ 0.023192f
C16513 _449_/a_1204_472# _038_ 0.005899f
C16514 FILLER_0_18_177/a_1020_375# FILLER_0_19_187/a_36_472# 0.001684f
C16515 FILLER_0_3_172/a_932_472# vdd 0.009887f
C16516 _062_ FILLER_0_5_136/a_36_472# 0.001404f
C16517 _413_/a_448_472# net59 0.059041f
C16518 FILLER_0_5_54/a_932_472# _440_/a_36_151# 0.001723f
C16519 _091_ FILLER_0_10_214/a_36_472# 0.001357f
C16520 FILLER_0_5_198/a_36_472# net21 0.014911f
C16521 FILLER_0_16_73/a_572_375# _176_ 0.006454f
C16522 net41 _452_/a_448_472# 0.052165f
C16523 FILLER_0_7_104/a_36_472# _058_ 0.006613f
C16524 net38 cal_count\[3\] 0.002225f
C16525 FILLER_0_14_107/a_1020_375# FILLER_0_16_115/a_36_472# 0.001512f
C16526 net16 _444_/a_2560_156# 0.010829f
C16527 cal_itt\[1\] _084_ 0.495918f
C16528 FILLER_0_10_28/a_36_472# net6 0.038613f
C16529 _069_ _122_ 0.002164f
C16530 _077_ _439_/a_796_472# 0.007471f
C16531 net19 _044_ 0.138869f
C16532 _105_ vss 0.485198f
C16533 output10/a_224_472# net8 0.010088f
C16534 trim_val\[4\] net22 0.144267f
C16535 _430_/a_448_472# vdd 0.002959f
C16536 _102_ _094_ 0.727442f
C16537 ctlp[0] vdd 0.08832f
C16538 FILLER_0_18_76/a_484_472# net71 0.004649f
C16539 net53 net74 0.164124f
C16540 _144_ _433_/a_796_472# 0.008448f
C16541 net45 vdd 0.087369f
C16542 trimb[3] vss 0.161605f
C16543 mask\[2\] FILLER_0_15_235/a_572_375# 0.003879f
C16544 FILLER_0_5_181/a_124_375# vss 0.011456f
C16545 FILLER_0_5_181/a_36_472# vdd 0.081434f
C16546 FILLER_0_4_197/a_932_472# _088_ 0.014643f
C16547 _360_/a_36_160# vss 0.028817f
C16548 vss output6/a_224_472# 0.004205f
C16549 FILLER_0_9_28/a_124_375# net17 0.009179f
C16550 net34 _297_/a_36_472# 0.005603f
C16551 _106_ _291_/a_36_160# 0.054237f
C16552 FILLER_0_22_177/a_484_472# mask\[6\] 0.006573f
C16553 FILLER_0_22_177/a_124_375# _146_ 0.001864f
C16554 net35 FILLER_0_22_177/a_36_472# 0.005721f
C16555 mask\[2\] vdd 0.433058f
C16556 _098_ _205_/a_36_160# 0.033853f
C16557 mask\[9\] FILLER_0_18_76/a_572_375# 0.006158f
C16558 _195_/a_67_603# mask\[1\] 0.016836f
C16559 net15 ctln[9] 0.01475f
C16560 net70 FILLER_0_17_104/a_1020_375# 0.001894f
C16561 FILLER_0_5_109/a_572_375# _153_ 0.03228f
C16562 net76 FILLER_0_5_206/a_36_472# 0.00169f
C16563 _171_ vss 0.004501f
C16564 FILLER_0_13_206/a_36_472# net79 0.00402f
C16565 net54 _149_ 0.212511f
C16566 net54 FILLER_0_18_139/a_572_375# 0.00217f
C16567 output48/a_224_472# vss 0.006655f
C16568 net20 mask\[2\] 0.050364f
C16569 cal_itt\[2\] net59 0.014956f
C16570 _077_ FILLER_0_8_127/a_36_472# 0.003023f
C16571 cal_count\[3\] _067_ 0.478427f
C16572 mask\[4\] FILLER_0_18_209/a_124_375# 0.020811f
C16573 mask\[3\] _289_/a_36_472# 0.02347f
C16574 output42/a_224_472# _236_/a_36_160# 0.001892f
C16575 FILLER_0_8_247/a_124_375# vss 0.002674f
C16576 FILLER_0_8_247/a_572_375# vdd -0.007963f
C16577 _105_ _107_ 0.020727f
C16578 _085_ _267_/a_36_472# 0.034055f
C16579 ctln[4] FILLER_0_0_198/a_36_472# 0.02582f
C16580 output43/a_224_472# trimb[3] 0.070044f
C16581 _430_/a_2248_156# mask\[2\] 0.009336f
C16582 mask\[0\] vss 0.694674f
C16583 trim_val\[1\] _166_ 0.06773f
C16584 _399_/a_224_472# net72 0.002538f
C16585 _015_ FILLER_0_10_247/a_124_375# 0.001261f
C16586 _300_/a_224_472# vdd 0.001344f
C16587 _057_ net22 0.163773f
C16588 FILLER_0_13_100/a_36_472# vss 0.003094f
C16589 FILLER_0_5_206/a_124_375# FILLER_0_5_198/a_572_375# 0.012001f
C16590 _096_ net79 0.015605f
C16591 net34 FILLER_0_22_128/a_2724_472# 0.004465f
C16592 _441_/a_36_151# _164_ 0.008955f
C16593 trim_mask\[2\] _036_ 0.466145f
C16594 comp cal_count\[2\] 0.015029f
C16595 _179_ vss 0.089947f
C16596 _163_ _156_ 0.001616f
C16597 net3 _278_/a_36_160# 0.014154f
C16598 _178_ _179_ 0.063494f
C16599 _046_ _282_/a_36_160# 0.005584f
C16600 FILLER_0_20_107/a_36_472# net71 0.004375f
C16601 _185_ net17 0.270086f
C16602 _095_ FILLER_0_14_107/a_932_472# 0.014431f
C16603 _420_/a_2248_156# vdd 0.00331f
C16604 _411_/a_1204_472# vss 0.001746f
C16605 output17/a_224_472# ctlp[0] 0.018696f
C16606 FILLER_0_15_205/a_124_375# net22 0.049201f
C16607 net4 FILLER_0_12_220/a_932_472# 0.050731f
C16608 net45 output17/a_224_472# 0.01994f
C16609 net3 vss 0.02666f
C16610 net24 net71 0.015101f
C16611 cal net1 0.336092f
C16612 _032_ vdd 0.174834f
C16613 vdd FILLER_0_16_115/a_124_375# 0.020393f
C16614 net58 output37/a_224_472# 0.099539f
C16615 FILLER_0_10_256/a_36_472# net28 0.00136f
C16616 _178_ net3 0.257606f
C16617 _098_ FILLER_0_15_180/a_124_375# 0.019007f
C16618 comp input3/a_36_113# 0.022213f
C16619 _104_ _109_ 0.029532f
C16620 _242_/a_36_160# vss 0.032884f
C16621 _444_/a_1000_472# net67 0.025169f
C16622 FILLER_0_21_125/a_572_375# net54 0.024701f
C16623 _136_ _019_ 0.049263f
C16624 _113_ FILLER_0_12_196/a_36_472# 0.002495f
C16625 net52 _443_/a_1000_472# 0.016322f
C16626 net20 _420_/a_2248_156# 0.003737f
C16627 _446_/a_2665_112# net49 0.006979f
C16628 trim_val\[4\] vdd 0.245329f
C16629 net44 _450_/a_836_156# 0.006278f
C16630 FILLER_0_16_57/a_124_375# vdd 0.008567f
C16631 net67 FILLER_0_8_24/a_484_472# 0.001065f
C16632 vdd _450_/a_3129_107# 0.039939f
C16633 _028_ FILLER_0_8_107/a_36_472# 0.002173f
C16634 net35 _436_/a_1308_423# 0.008773f
C16635 result[4] net77 0.003336f
C16636 _091_ _429_/a_448_472# 0.034713f
C16637 ctln[4] FILLER_0_0_232/a_124_375# 0.002726f
C16638 FILLER_0_3_78/a_36_472# _160_ 0.006564f
C16639 _330_/a_224_472# _134_ 0.007508f
C16640 _174_ _401_/a_244_472# 0.001957f
C16641 net34 _210_/a_67_603# 0.01049f
C16642 net48 _251_/a_906_472# 0.001362f
C16643 _322_/a_848_380# _068_ 0.009682f
C16644 _063_ FILLER_0_6_37/a_124_375# 0.012149f
C16645 net52 _448_/a_2665_112# 0.039348f
C16646 trimb[0] FILLER_0_20_2/a_124_375# 0.006864f
C16647 ctln[4] net11 0.194506f
C16648 FILLER_0_15_212/a_124_375# vss 0.005813f
C16649 FILLER_0_15_212/a_572_375# vdd -0.014642f
C16650 _239_/a_36_160# vdd 0.042369f
C16651 output37/a_224_472# calibrate 0.013149f
C16652 _099_ vss 0.255039f
C16653 net57 _017_ 0.045694f
C16654 _093_ _438_/a_448_472# 0.0106f
C16655 net15 FILLER_0_18_76/a_36_472# 0.001341f
C16656 _131_ _180_ 0.016104f
C16657 calibrate _385_/a_36_68# 0.001996f
C16658 _415_/a_2665_112# net64 0.074373f
C16659 FILLER_0_20_177/a_36_472# _434_/a_36_151# 0.001723f
C16660 FILLER_0_20_177/a_1468_375# _434_/a_448_472# 0.008952f
C16661 FILLER_0_4_99/a_36_472# vss 0.002273f
C16662 net32 _419_/a_1308_423# 0.00191f
C16663 FILLER_0_16_154/a_484_472# vdd 0.001006f
C16664 FILLER_0_16_154/a_36_472# vss 0.005098f
C16665 FILLER_0_4_197/a_36_472# _270_/a_36_472# 0.004546f
C16666 _132_ _140_ 0.019255f
C16667 net64 FILLER_0_12_236/a_572_375# 0.005704f
C16668 net31 _006_ 0.307613f
C16669 net27 FILLER_0_9_270/a_572_375# 0.043797f
C16670 trim_mask\[1\] FILLER_0_6_47/a_572_375# 0.007164f
C16671 FILLER_0_19_111/a_572_375# vdd -0.008314f
C16672 ctln[6] _031_ 0.004486f
C16673 net75 _305_/a_36_159# 0.049563f
C16674 FILLER_0_16_73/a_36_472# net55 0.002576f
C16675 _065_ _168_ 0.020406f
C16676 _236_/a_36_160# net40 0.035082f
C16677 _421_/a_1000_472# _010_ 0.01379f
C16678 FILLER_0_22_86/a_1380_472# net14 0.039176f
C16679 _308_/a_124_24# net50 0.02221f
C16680 _419_/a_2665_112# vdd 0.030085f
C16681 _074_ _078_ 0.003088f
C16682 net31 _103_ 0.227588f
C16683 _000_ FILLER_0_0_232/a_124_375# 0.001391f
C16684 FILLER_0_15_59/a_124_375# vdd 0.017243f
C16685 net32 output35/a_224_472# 0.072991f
C16686 _412_/a_36_151# cal_itt\[1\] 0.025078f
C16687 FILLER_0_19_47/a_572_375# net55 0.003447f
C16688 _116_ FILLER_0_12_196/a_124_375# 0.005332f
C16689 _430_/a_1308_423# _069_ 0.024499f
C16690 net19 _420_/a_2560_156# 0.010978f
C16691 _076_ _078_ 0.012626f
C16692 net50 FILLER_0_6_37/a_124_375# 0.003821f
C16693 net54 FILLER_0_20_107/a_124_375# 0.072539f
C16694 _142_ FILLER_0_17_142/a_36_472# 0.011216f
C16695 mask\[7\] FILLER_0_22_177/a_572_375# 0.001315f
C16696 FILLER_0_15_116/a_36_472# _451_/a_36_151# 0.096503f
C16697 FILLER_0_19_195/a_124_375# _202_/a_36_160# 0.005489f
C16698 net76 FILLER_0_3_172/a_1380_472# 0.015215f
C16699 comp _043_ 0.003867f
C16700 FILLER_0_7_146/a_124_375# _133_ 0.001577f
C16701 _057_ vdd 0.801978f
C16702 net52 trim_mask\[1\] 0.04149f
C16703 net72 _453_/a_36_151# 0.001607f
C16704 result[8] vss 0.235206f
C16705 _079_ _260_/a_36_68# 0.043596f
C16706 _430_/a_1204_472# _069_ 0.001629f
C16707 result[9] FILLER_0_24_274/a_36_472# 0.009425f
C16708 _002_ net22 0.038848f
C16709 _064_ _445_/a_36_151# 0.03209f
C16710 FILLER_0_13_212/a_36_472# net79 0.006158f
C16711 cal_count\[3\] net23 0.045417f
C16712 _003_ net37 0.046745f
C16713 FILLER_0_18_177/a_3260_375# _205_/a_36_160# 0.001313f
C16714 mask\[4\] _339_/a_36_160# 0.003234f
C16715 net62 FILLER_0_13_212/a_484_472# 0.059367f
C16716 FILLER_0_3_204/a_36_472# FILLER_0_3_172/a_3172_472# 0.013276f
C16717 _069_ FILLER_0_11_142/a_572_375# 0.020472f
C16718 _095_ mask\[1\] 0.001297f
C16719 net49 trim_mask\[1\] 0.003402f
C16720 output39/a_224_472# net67 0.008957f
C16721 result[6] ctlp[1] 0.677825f
C16722 FILLER_0_18_107/a_3172_472# _145_ 0.002415f
C16723 net4 FILLER_0_3_221/a_484_472# 0.043027f
C16724 _059_ net23 0.265909f
C16725 mask\[7\] _435_/a_2560_156# 0.011544f
C16726 FILLER_0_16_73/a_484_472# vdd 0.003462f
C16727 result[8] _422_/a_1000_472# 0.001104f
C16728 FILLER_0_15_142/a_124_375# vss 0.009207f
C16729 net69 FILLER_0_2_101/a_36_472# 0.00845f
C16730 _075_ _053_ 0.634359f
C16731 _143_ _140_ 0.00806f
C16732 FILLER_0_15_205/a_124_375# vdd 0.015886f
C16733 _414_/a_1000_472# net22 0.001649f
C16734 FILLER_0_1_212/a_36_472# vss 0.00858f
C16735 _450_/a_1040_527# output6/a_224_472# 0.005581f
C16736 _450_/a_448_472# net6 0.041113f
C16737 FILLER_0_17_200/a_572_375# vss 0.017327f
C16738 _089_ _087_ 0.002217f
C16739 FILLER_0_19_125/a_36_472# vdd 0.003414f
C16740 _092_ _093_ 0.287983f
C16741 net52 _157_ 0.005889f
C16742 state\[0\] _128_ 0.228492f
C16743 trim_val\[3\] vdd 0.211478f
C16744 FILLER_0_5_128/a_36_472# _152_ 0.013822f
C16745 _079_ net4 0.023763f
C16746 _181_ cal_count\[1\] 0.186904f
C16747 result[7] result[9] 1.21288f
C16748 FILLER_0_12_220/a_1020_375# vss 0.004698f
C16749 FILLER_0_12_220/a_1468_375# vdd 0.002801f
C16750 _115_ _129_ 0.021405f
C16751 net63 mask\[3\] 0.37365f
C16752 net41 cal_count\[3\] 0.028902f
C16753 _132_ _451_/a_36_151# 0.007777f
C16754 net1 net37 0.00519f
C16755 _426_/a_2248_156# calibrate 0.004597f
C16756 cal_count\[3\] FILLER_0_11_109/a_124_375# 0.004618f
C16757 FILLER_0_18_139/a_1380_472# vss 0.009272f
C16758 net74 _058_ 0.026905f
C16759 net63 _434_/a_448_472# 0.008139f
C16760 result[9] FILLER_0_15_282/a_36_472# 0.003213f
C16761 _432_/a_36_151# net57 0.00484f
C16762 _093_ net70 0.001888f
C16763 _028_ _163_ 0.199021f
C16764 FILLER_0_9_28/a_2364_375# vdd 0.004562f
C16765 trim_val\[4\] FILLER_0_2_165/a_124_375# 0.009193f
C16766 output39/a_224_472# _445_/a_448_472# 0.009352f
C16767 FILLER_0_9_72/a_1468_375# _439_/a_2248_156# 0.001901f
C16768 FILLER_0_5_72/a_1020_375# _029_ 0.010208f
C16769 FILLER_0_22_177/a_1468_375# vss 0.028064f
C16770 FILLER_0_22_177/a_36_472# vdd 0.111906f
C16771 FILLER_0_17_200/a_124_375# _093_ 0.00419f
C16772 net48 net76 0.069349f
C16773 result[8] _107_ 0.041984f
C16774 _099_ _195_/a_67_603# 0.065049f
C16775 _390_/a_36_68# _038_ 0.019355f
C16776 net20 FILLER_0_12_220/a_1468_375# 0.016974f
C16777 _114_ _121_ 0.002513f
C16778 FILLER_0_16_89/a_572_375# net14 0.00106f
C16779 FILLER_0_4_144/a_36_472# _081_ 0.003547f
C16780 FILLER_0_21_125/a_124_375# _022_ 0.007023f
C16781 net7 _065_ 0.0295f
C16782 mask\[2\] FILLER_0_16_154/a_572_375# 0.026605f
C16783 _053_ calibrate 0.081635f
C16784 _401_/a_36_68# _179_ 0.007074f
C16785 FILLER_0_4_107/a_1468_375# _160_ 0.028099f
C16786 _443_/a_2665_112# _066_ 0.001654f
C16787 FILLER_0_4_213/a_124_375# vss 0.006145f
C16788 FILLER_0_4_213/a_572_375# vdd 0.026692f
C16789 net25 _213_/a_67_603# 0.027452f
C16790 net18 FILLER_0_17_282/a_36_472# 0.036965f
C16791 _024_ _023_ 0.005966f
C16792 _430_/a_796_472# _019_ 0.006511f
C16793 _070_ FILLER_0_5_164/a_572_375# 0.001083f
C16794 _140_ _146_ 0.135012f
C16795 _418_/a_36_151# _007_ 0.007397f
C16796 FILLER_0_22_86/a_124_375# _098_ 0.011864f
C16797 FILLER_0_17_72/a_1020_375# _131_ 0.005847f
C16798 fanout62/a_36_160# net79 0.011515f
C16799 _061_ _247_/a_36_160# 0.009993f
C16800 _115_ FILLER_0_10_78/a_1020_375# 0.064761f
C16801 _136_ _451_/a_2225_156# 0.01289f
C16802 _367_/a_36_68# vdd 0.010246f
C16803 _053_ net21 0.036284f
C16804 _449_/a_796_472# vss 0.00143f
C16805 FILLER_0_21_286/a_36_472# net77 0.001557f
C16806 _430_/a_448_472# _069_ 0.047845f
C16807 _106_ _104_ 0.17237f
C16808 net70 FILLER_0_14_123/a_36_472# 0.009456f
C16809 _103_ net77 0.004691f
C16810 _091_ FILLER_0_15_180/a_484_472# 0.001757f
C16811 net4 cal_itt\[1\] 0.048147f
C16812 FILLER_0_9_142/a_124_375# _315_/a_36_68# 0.028077f
C16813 _149_ _437_/a_1204_472# 0.024276f
C16814 _026_ _437_/a_796_472# 0.008884f
C16815 _115_ FILLER_0_10_78/a_124_375# 0.001718f
C16816 _111_ _098_ 0.014998f
C16817 mask\[3\] FILLER_0_17_161/a_124_375# 0.032905f
C16818 cal_count\[2\] _183_ 0.034303f
C16819 fanout49/a_36_160# FILLER_0_3_78/a_484_472# 0.003699f
C16820 _078_ _081_ 0.445443f
C16821 _451_/a_1353_112# _040_ 0.005265f
C16822 trim_val\[0\] vdd 0.056059f
C16823 net34 _109_ 0.001298f
C16824 output36/a_224_472# FILLER_0_14_263/a_36_472# 0.001711f
C16825 _122_ FILLER_0_6_231/a_484_472# 0.017477f
C16826 _123_ FILLER_0_6_231/a_124_375# 0.001259f
C16827 _069_ mask\[2\] 0.032781f
C16828 ctln[2] vss 0.256543f
C16829 _077_ FILLER_0_9_28/a_3172_472# 0.011059f
C16830 _176_ net14 0.031922f
C16831 FILLER_0_14_263/a_36_472# net30 0.003972f
C16832 net64 _282_/a_36_160# 0.014431f
C16833 _002_ vdd 0.152662f
C16834 output38/a_224_472# _445_/a_36_151# 0.199812f
C16835 FILLER_0_7_233/a_124_375# FILLER_0_6_231/a_484_472# 0.001684f
C16836 _413_/a_36_151# net65 0.033028f
C16837 sample result[0] 0.081581f
C16838 _176_ fanout55/a_36_160# 0.070942f
C16839 output18/a_224_472# vss 0.086897f
C16840 _016_ FILLER_0_12_124/a_124_375# 0.007335f
C16841 _449_/a_36_151# _174_ 0.002252f
C16842 net60 _109_ 0.021502f
C16843 _196_/a_36_160# FILLER_0_14_263/a_124_375# 0.005732f
C16844 net16 _164_ 0.015161f
C16845 _430_/a_1000_472# net36 0.001836f
C16846 FILLER_0_17_200/a_36_472# net63 0.005648f
C16847 _425_/a_36_151# _317_/a_36_113# 0.002361f
C16848 net34 net54 0.003682f
C16849 _137_ FILLER_0_15_180/a_572_375# 0.028083f
C16850 FILLER_0_18_2/a_1020_375# trimb[1] 0.01376f
C16851 _414_/a_1000_472# vdd 0.002568f
C16852 _072_ _247_/a_36_160# 0.005008f
C16853 net63 FILLER_0_22_177/a_932_472# 0.060639f
C16854 net80 _337_/a_49_472# 0.015686f
C16855 net18 FILLER_0_9_270/a_572_375# 0.005977f
C16856 output24/a_224_472# _436_/a_448_472# 0.009204f
C16857 output32/a_224_472# result[7] 0.063135f
C16858 _091_ FILLER_0_20_169/a_124_375# 0.003958f
C16859 _020_ net36 0.001995f
C16860 _445_/a_2248_156# vdd 0.018573f
C16861 _372_/a_2590_472# _059_ 0.002974f
C16862 FILLER_0_21_28/a_2724_472# vdd 0.001342f
C16863 _436_/a_1308_423# vdd 0.005258f
C16864 net55 net17 0.056153f
C16865 FILLER_0_3_221/a_572_375# vss 0.003292f
C16866 _114_ _132_ 0.08562f
C16867 _423_/a_1204_472# _012_ 0.003181f
C16868 ctln[1] vss 0.27233f
C16869 net36 _438_/a_796_472# 0.016855f
C16870 net16 _404_/a_36_472# 0.001126f
C16871 _428_/a_2248_156# _427_/a_36_151# 0.035837f
C16872 _439_/a_448_472# vss 0.036535f
C16873 _439_/a_1308_423# vdd 0.002368f
C16874 net81 _426_/a_1308_423# 0.002332f
C16875 _126_ FILLER_0_13_100/a_124_375# 0.00134f
C16876 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_124_375# 0.012222f
C16877 FILLER_0_9_28/a_124_375# FILLER_0_8_24/a_572_375# 0.05841f
C16878 FILLER_0_8_239/a_36_472# _123_ 0.011767f
C16879 mask\[0\] _095_ 0.006711f
C16880 net20 FILLER_0_3_221/a_1020_375# 0.025371f
C16881 FILLER_0_21_28/a_2812_375# _424_/a_36_151# 0.059049f
C16882 _427_/a_2665_112# net23 0.032729f
C16883 output47/a_224_472# vdd 0.028666f
C16884 _095_ FILLER_0_13_100/a_36_472# 0.003036f
C16885 FILLER_0_4_144/a_484_472# _443_/a_36_151# 0.002841f
C16886 net70 _136_ 0.032219f
C16887 _050_ _025_ 0.033887f
C16888 _091_ FILLER_0_18_177/a_932_472# 0.002113f
C16889 fanout62/a_36_160# FILLER_0_13_290/a_124_375# 0.001138f
C16890 mask\[7\] _147_ 0.295801f
C16891 trim[0] trim[1] 0.001567f
C16892 FILLER_0_10_37/a_124_375# FILLER_0_10_28/a_124_375# 0.003228f
C16893 _002_ FILLER_0_3_172/a_2812_375# 0.006403f
C16894 _190_/a_36_160# net47 0.001489f
C16895 ctlp[1] fanout77/a_36_113# 0.012793f
C16896 net50 FILLER_0_6_90/a_124_375# 0.041764f
C16897 FILLER_0_12_2/a_124_375# vdd 0.0247f
C16898 FILLER_0_0_266/a_36_472# vss 0.003738f
C16899 ctln[7] _442_/a_2665_112# 0.01075f
C16900 FILLER_0_7_72/a_36_472# _439_/a_448_472# 0.008036f
C16901 FILLER_0_10_214/a_36_472# net22 0.001634f
C16902 _112_ _425_/a_1204_472# 0.001132f
C16903 _375_/a_36_68# calibrate 0.048799f
C16904 FILLER_0_6_239/a_36_472# net37 0.004187f
C16905 net56 FILLER_0_19_142/a_124_375# 0.003154f
C16906 FILLER_0_16_57/a_484_472# _176_ 0.013507f
C16907 net3 _095_ 0.002383f
C16908 net53 _451_/a_2225_156# 0.011677f
C16909 result[6] _421_/a_2560_156# 0.006943f
C16910 FILLER_0_4_197/a_124_375# net21 0.018398f
C16911 net67 net6 0.345681f
C16912 FILLER_0_9_28/a_1828_472# _054_ 0.003145f
C16913 net15 FILLER_0_5_72/a_124_375# 0.006403f
C16914 _077_ _453_/a_448_472# 0.057515f
C16915 _176_ FILLER_0_11_109/a_36_472# 0.002951f
C16916 _208_/a_36_160# vdd 0.014709f
C16917 _431_/a_448_472# _137_ 0.008493f
C16918 net62 FILLER_0_15_228/a_124_375# 0.001408f
C16919 _415_/a_448_472# FILLER_0_9_270/a_36_472# 0.012285f
C16920 FILLER_0_21_150/a_36_472# _146_ 0.00236f
C16921 net55 _216_/a_67_603# 0.071821f
C16922 net80 net81 0.006516f
C16923 _370_/a_692_472# _152_ 0.005908f
C16924 _370_/a_1152_472# _081_ 0.001901f
C16925 _431_/a_36_151# net70 0.031018f
C16926 net57 cal_count\[3\] 0.02848f
C16927 _359_/a_36_488# _062_ 0.005596f
C16928 net69 FILLER_0_3_78/a_124_375# 0.004201f
C16929 _087_ FILLER_0_3_172/a_1916_375# 0.001223f
C16930 _115_ _068_ 0.889978f
C16931 fanout61/a_36_113# net78 0.009579f
C16932 _126_ _055_ 0.01647f
C16933 _028_ FILLER_0_7_104/a_1020_375# 0.004954f
C16934 _111_ net55 0.002855f
C16935 _013_ net72 0.006579f
C16936 FILLER_0_1_98/a_36_472# net52 0.005688f
C16937 FILLER_0_9_28/a_1828_472# vss 0.001663f
C16938 fanout67/a_36_160# trim_val\[0\] 0.003096f
C16939 _432_/a_2248_156# _093_ 0.012955f
C16940 FILLER_0_7_195/a_124_375# _161_ 0.005368f
C16941 _132_ FILLER_0_17_104/a_1380_472# 0.02114f
C16942 result[0] FILLER_0_9_282/a_572_375# 0.042859f
C16943 net50 FILLER_0_4_91/a_484_472# 0.008749f
C16944 net82 _082_ 0.286003f
C16945 _127_ _120_ 0.198577f
C16946 _144_ FILLER_0_21_125/a_124_375# 0.009117f
C16947 net62 _417_/a_1204_472# 0.001941f
C16948 _114_ FILLER_0_10_94/a_484_472# 0.011954f
C16949 _151_ vss 0.050544f
C16950 FILLER_0_8_127/a_36_472# _125_ 0.003088f
C16951 _415_/a_1204_472# result[1] 0.004051f
C16952 output48/a_224_472# output37/a_224_472# 0.005147f
C16953 FILLER_0_9_223/a_36_472# state\[0\] 0.002846f
C16954 output34/a_224_472# net30 0.002189f
C16955 FILLER_0_6_47/a_36_472# vss 0.002433f
C16956 FILLER_0_6_47/a_484_472# vdd 0.005065f
C16957 FILLER_0_9_282/a_124_375# vdd 0.01273f
C16958 _086_ _250_/a_36_68# 0.001132f
C16959 net15 FILLER_0_15_72/a_36_472# 0.007185f
C16960 net82 fanout57/a_36_113# 0.017696f
C16961 net34 _350_/a_49_472# 0.008001f
C16962 fanout58/a_36_160# vss 0.039959f
C16963 net27 vss 0.534444f
C16964 _057_ _069_ 0.053765f
C16965 mask\[8\] FILLER_0_22_107/a_572_375# 0.030641f
C16966 net35 FILLER_0_22_107/a_124_375# 0.010439f
C16967 _432_/a_448_472# _137_ 0.008956f
C16968 net16 _217_/a_36_160# 0.00629f
C16969 FILLER_0_16_255/a_36_472# _006_ 0.006621f
C16970 _431_/a_1000_472# _137_ 0.010168f
C16971 _053_ FILLER_0_7_104/a_124_375# 0.012564f
C16972 FILLER_0_11_135/a_36_472# _120_ 0.012562f
C16973 _106_ net34 0.013009f
C16974 cal_count\[2\] _402_/a_718_527# 0.004645f
C16975 mask\[0\] FILLER_0_12_236/a_36_472# 0.002801f
C16976 net32 _421_/a_36_151# 0.008275f
C16977 _402_/a_1296_93# _179_ 0.001692f
C16978 net70 net53 1.170795f
C16979 _322_/a_124_24# _118_ 0.04952f
C16980 FILLER_0_13_212/a_1020_375# vdd -0.014642f
C16981 FILLER_0_13_212/a_572_375# vss 0.007991f
C16982 _093_ FILLER_0_17_218/a_36_472# 0.006994f
C16983 _429_/a_2665_112# FILLER_0_15_228/a_124_375# 0.001077f
C16984 FILLER_0_19_55/a_36_472# FILLER_0_19_47/a_484_472# 0.013276f
C16985 _069_ FILLER_0_15_205/a_124_375# 0.002728f
C16986 net38 net49 0.117427f
C16987 FILLER_0_7_72/a_1468_375# FILLER_0_5_72/a_1380_472# 0.00108f
C16988 FILLER_0_10_78/a_1468_375# _176_ 0.013408f
C16989 mask\[4\] _202_/a_36_160# 0.007912f
C16990 _395_/a_244_68# _070_ 0.001481f
C16991 net52 _158_ 0.001338f
C16992 FILLER_0_11_101/a_36_472# _120_ 0.007656f
C16993 _421_/a_1204_472# vdd 0.002198f
C16994 FILLER_0_10_214/a_36_472# vdd 0.026621f
C16995 FILLER_0_10_214/a_124_375# vss 0.013034f
C16996 FILLER_0_15_142/a_124_375# _095_ 0.003935f
C16997 _446_/a_1308_423# net17 0.033125f
C16998 net73 vss 0.342554f
C16999 fanout63/a_36_160# net36 0.004435f
C17000 net79 _101_ 0.014383f
C17001 net31 _419_/a_2665_112# 0.004446f
C17002 net20 FILLER_0_13_212/a_1020_375# 0.003962f
C17003 _023_ mask\[6\] 0.077441f
C17004 ctlp[3] ctlp[4] 0.027598f
C17005 FILLER_0_8_37/a_484_472# _054_ 0.022621f
C17006 FILLER_0_19_187/a_124_375# vdd 0.030349f
C17007 _404_/a_36_472# _041_ 0.003068f
C17008 vss FILLER_0_21_60/a_572_375# 0.021222f
C17009 vdd FILLER_0_21_60/a_36_472# 0.08419f
C17010 net26 FILLER_0_23_44/a_484_472# 0.003796f
C17011 net73 FILLER_0_18_107/a_1020_375# 0.04487f
C17012 net20 _421_/a_1204_472# 0.019627f
C17013 _052_ mask\[9\] 0.007224f
C17014 _096_ _320_/a_1568_472# 0.001632f
C17015 _429_/a_448_472# net22 0.054866f
C17016 _429_/a_36_151# _018_ 0.118135f
C17017 FILLER_0_2_111/a_572_375# vdd 0.012666f
C17018 _315_/a_244_497# _059_ 0.00101f
C17019 fanout82/a_36_113# vdd 0.083174f
C17020 _410_/a_36_68# _188_ 0.007731f
C17021 _187_ cal_count\[3\] 0.031898f
C17022 result[5] result[9] 0.064058f
C17023 output44/a_224_472# _452_/a_1353_112# 0.001321f
C17024 _130_ _427_/a_36_151# 0.001056f
C17025 _440_/a_448_472# vdd 0.007263f
C17026 _440_/a_36_151# vss 0.016458f
C17027 output45/a_224_472# net40 0.001284f
C17028 _091_ _113_ 0.006236f
C17029 net76 net37 0.549565f
C17030 net29 _045_ 0.344478f
C17031 net58 fanout64/a_36_160# 0.002438f
C17032 _098_ net21 0.133694f
C17033 FILLER_0_8_37/a_484_472# vss 0.001267f
C17034 _077_ FILLER_0_9_60/a_124_375# 0.051389f
C17035 ctln[3] vdd 0.167569f
C17036 net66 net49 0.657679f
C17037 _083_ net59 0.408831f
C17038 _093_ _199_/a_36_160# 0.05226f
C17039 output25/a_224_472# net24 0.002325f
C17040 FILLER_0_21_28/a_3260_375# _012_ 0.016427f
C17041 _130_ _321_/a_170_472# 0.001018f
C17042 net1 net8 0.00497f
C17043 net70 FILLER_0_14_107/a_124_375# 0.029975f
C17044 FILLER_0_5_72/a_1380_472# vdd 0.001438f
C17045 FILLER_0_5_72/a_932_472# vss 0.003084f
C17046 _205_/a_36_160# net21 0.020847f
C17047 _098_ FILLER_0_19_171/a_932_472# 0.003573f
C17048 FILLER_0_20_2/a_124_375# vdd 0.010886f
C17049 FILLER_0_5_54/a_932_472# _029_ 0.014976f
C17050 FILLER_0_5_54/a_1468_375# trim_mask\[1\] 0.010901f
C17051 _075_ _070_ 0.009314f
C17052 ctlp[1] _419_/a_36_151# 0.015335f
C17053 _106_ _276_/a_36_160# 0.009097f
C17054 _086_ _310_/a_49_472# 0.013039f
C17055 fanout63/a_36_160# FILLER_0_15_228/a_36_472# 0.014197f
C17056 fanout64/a_36_160# calibrate 0.001117f
C17057 _451_/a_836_156# vdd 0.003786f
C17058 _232_/a_67_603# _167_ 0.014152f
C17059 _062_ FILLER_0_8_156/a_572_375# 0.002944f
C17060 _446_/a_2665_112# net40 0.027712f
C17061 _077_ trim_mask\[0\] 0.090587f
C17062 _070_ FILLER_0_10_94/a_36_472# 0.001866f
C17063 _448_/a_36_151# net65 0.001983f
C17064 _426_/a_36_151# FILLER_0_8_247/a_932_472# 0.001723f
C17065 net57 _427_/a_2665_112# 0.016685f
C17066 FILLER_0_5_198/a_124_375# net37 0.009149f
C17067 result[7] net78 0.019651f
C17068 vdd _034_ 0.424437f
C17069 _272_/a_36_472# _089_ 0.003862f
C17070 net42 _039_ 0.001096f
C17071 _443_/a_36_151# FILLER_0_2_127/a_36_472# 0.006095f
C17072 _162_ vss 0.08357f
C17073 _161_ vdd 0.262564f
C17074 FILLER_0_5_128/a_572_375# FILLER_0_5_136/a_36_472# 0.086635f
C17075 _421_/a_2665_112# net19 0.01849f
C17076 _131_ FILLER_0_9_105/a_484_472# 0.004364f
C17077 FILLER_0_8_138/a_36_472# _129_ 0.055537f
C17078 _008_ _418_/a_2560_156# 0.006651f
C17079 FILLER_0_13_206/a_124_375# _043_ 0.014212f
C17080 _379_/a_36_472# net47 0.016584f
C17081 net63 FILLER_0_19_187/a_36_472# 0.006753f
C17082 _282_/a_36_160# mask\[2\] 0.023533f
C17083 _095_ _402_/a_56_567# 0.010012f
C17084 _164_ FILLER_0_6_47/a_124_375# 0.069738f
C17085 _132_ _137_ 0.023462f
C17086 FILLER_0_18_2/a_572_375# output44/a_224_472# 0.001296f
C17087 state\[1\] _055_ 0.067603f
C17088 _129_ vdd 0.314544f
C17089 trimb[1] FILLER_0_19_28/a_36_472# 0.01233f
C17090 _131_ vss 0.549133f
C17091 mask\[4\] FILLER_0_18_177/a_1020_375# 0.015941f
C17092 _397_/a_36_472# _175_ 0.004667f
C17093 _070_ calibrate 0.675125f
C17094 _042_ _039_ 0.003075f
C17095 _165_ trim_mask\[1\] 0.002231f
C17096 ctlp[4] _108_ 0.002002f
C17097 net75 _001_ 0.056236f
C17098 output38/a_224_472# FILLER_0_3_2/a_36_472# 0.035046f
C17099 net16 _378_/a_224_472# 0.001007f
C17100 output9/a_224_472# FILLER_0_1_266/a_36_472# 0.001007f
C17101 FILLER_0_7_146/a_36_472# calibrate 0.060587f
C17102 _005_ _193_/a_36_160# 0.009892f
C17103 trim_mask\[2\] fanout49/a_36_160# 0.12844f
C17104 _372_/a_3662_472# _062_ 0.0012f
C17105 net79 _094_ 0.301878f
C17106 _418_/a_36_151# _417_/a_36_151# 0.005373f
C17107 FILLER_0_16_107/a_572_375# vdd 0.019922f
C17108 _070_ net21 0.03068f
C17109 _009_ _296_/a_224_472# 0.001278f
C17110 FILLER_0_20_87/a_36_472# _437_/a_36_151# 0.001723f
C17111 _052_ FILLER_0_21_28/a_1468_375# 0.001757f
C17112 _086_ _395_/a_1044_488# 0.001091f
C17113 FILLER_0_18_2/a_3172_472# net41 0.00982f
C17114 _021_ FILLER_0_18_171/a_36_472# 0.103755f
C17115 FILLER_0_18_37/a_1020_375# vdd 0.020683f
C17116 _413_/a_448_472# _002_ 0.044695f
C17117 _412_/a_448_472# net19 0.001526f
C17118 _056_ net22 0.075673f
C17119 _399_/a_224_472# vdd 0.001593f
C17120 _447_/a_1308_423# net17 0.002531f
C17121 _030_ net14 0.079892f
C17122 result[5] output32/a_224_472# 0.047325f
C17123 _093_ FILLER_0_16_89/a_124_375# 0.004086f
C17124 _429_/a_36_151# vss 0.026298f
C17125 _429_/a_448_472# vdd 0.008822f
C17126 _057_ _267_/a_1792_472# 0.003005f
C17127 _076_ _080_ 0.005433f
C17128 _126_ state\[1\] 1.191746f
C17129 FILLER_0_7_195/a_36_472# _074_ 0.008706f
C17130 FILLER_0_10_78/a_1020_375# vdd 0.002901f
C17131 net10 FILLER_0_0_232/a_36_472# 0.016287f
C17132 _238_/a_67_603# vss 0.008203f
C17133 net18 vss 1.110302f
C17134 _144_ FILLER_0_18_107/a_1828_472# 0.001169f
C17135 _413_/a_1204_472# net82 0.00291f
C17136 vdd result[3] 0.181788f
C17137 output46/a_224_472# FILLER_0_20_2/a_572_375# 0.03228f
C17138 _030_ _164_ 0.036025f
C17139 net52 _066_ 0.022601f
C17140 net20 _429_/a_448_472# 0.002244f
C17141 FILLER_0_4_197/a_484_472# FILLER_0_3_172/a_3172_472# 0.026657f
C17142 _093_ FILLER_0_17_72/a_932_472# 0.004367f
C17143 fanout68/a_36_113# vss 0.006152f
C17144 _411_/a_448_472# vss 0.009447f
C17145 net41 _233_/a_36_160# 0.053625f
C17146 net56 vss 0.367812f
C17147 FILLER_0_10_78/a_124_375# vdd -0.011193f
C17148 net75 _014_ 0.204357f
C17149 _143_ _137_ 0.009932f
C17150 _426_/a_2665_112# _055_ 0.00142f
C17151 _306_/a_36_68# _113_ 0.010109f
C17152 _437_/a_2560_156# net14 0.00349f
C17153 _004_ _101_ 0.001514f
C17154 FILLER_0_15_142/a_36_472# fanout73/a_36_113# 0.009544f
C17155 fanout70/a_36_113# fanout73/a_36_113# 0.001578f
C17156 trim_mask\[1\] FILLER_0_6_79/a_124_375# 0.0042f
C17157 _310_/a_49_472# _090_ 0.059827f
C17158 net52 net23 0.093434f
C17159 _068_ net22 0.088209f
C17160 _395_/a_1492_488# _121_ 0.002537f
C17161 vdd FILLER_0_22_107/a_124_375# 0.029828f
C17162 FILLER_0_13_80/a_36_472# vss 0.009445f
C17163 _141_ FILLER_0_17_142/a_572_375# 0.029028f
C17164 net58 _425_/a_448_472# 0.002474f
C17165 _132_ FILLER_0_15_116/a_124_375# 0.047331f
C17166 FILLER_0_8_247/a_36_472# FILLER_0_8_239/a_36_472# 0.002296f
C17167 sample fanout65/a_36_113# 0.050978f
C17168 _297_/a_36_472# mask\[6\] 0.02557f
C17169 net72 FILLER_0_21_28/a_572_375# 0.005742f
C17170 ctlp[0] net43 0.003786f
C17171 net45 net43 0.131763f
C17172 net78 net79 0.009641f
C17173 _256_/a_36_68# _070_ 0.019259f
C17174 _115_ _308_/a_124_24# 0.039354f
C17175 _054_ _220_/a_67_603# 0.004333f
C17176 net58 _082_ 0.004276f
C17177 net55 _452_/a_2449_156# 0.015878f
C17178 net58 net82 0.022761f
C17179 fanout80/a_36_113# net36 0.007625f
C17180 _444_/a_1308_423# net17 0.028709f
C17181 _068_ _311_/a_2700_473# 0.001846f
C17182 FILLER_0_18_177/a_3260_375# net21 0.005704f
C17183 _394_/a_56_524# _174_ 0.015122f
C17184 _098_ mask\[1\] 1.476748f
C17185 _065_ net50 0.123581f
C17186 _425_/a_36_151# _122_ 0.063131f
C17187 _425_/a_448_472# calibrate 0.105581f
C17188 result[9] _108_ 0.015443f
C17189 FILLER_0_8_24/a_572_375# net17 0.007101f
C17190 FILLER_0_3_204/a_36_472# FILLER_0_4_197/a_932_472# 0.026657f
C17191 _424_/a_1000_472# _012_ 0.00675f
C17192 _104_ ctlp[1] 0.076863f
C17193 net62 FILLER_0_14_235/a_36_472# 0.00534f
C17194 FILLER_0_7_72/a_1916_375# net50 0.059471f
C17195 _033_ _444_/a_1000_472# 0.00692f
C17196 _165_ _444_/a_2665_112# 0.044447f
C17197 result[9] net19 0.540761f
C17198 FILLER_0_18_177/a_932_472# FILLER_0_19_171/a_1468_375# 0.001684f
C17199 FILLER_0_12_136/a_1020_375# net23 0.005919f
C17200 _048_ vss 0.056146f
C17201 cal_itt\[2\] FILLER_0_3_221/a_1020_375# 0.010951f
C17202 FILLER_0_18_171/a_124_375# FILLER_0_18_177/a_36_472# 0.016748f
C17203 net80 _434_/a_1308_423# 0.006837f
C17204 _417_/a_448_472# vss 0.005289f
C17205 _417_/a_1308_423# vdd 0.002263f
C17206 net41 net49 0.392356f
C17207 _232_/a_67_603# vdd 0.007565f
C17208 FILLER_0_4_123/a_36_472# vdd 0.091386f
C17209 fanout76/a_36_160# net18 0.003319f
C17210 FILLER_0_4_123/a_124_375# vss 0.009712f
C17211 FILLER_0_19_47/a_484_472# vss 0.001338f
C17212 net82 calibrate 0.002345f
C17213 _220_/a_67_603# vss 0.001485f
C17214 _114_ _097_ 0.004412f
C17215 net18 _416_/a_2248_156# 0.002106f
C17216 FILLER_0_19_55/a_124_375# _013_ 0.009611f
C17217 trim_mask\[3\] net14 0.142743f
C17218 _421_/a_448_472# _419_/a_2665_112# 0.002393f
C17219 _056_ vdd 0.423512f
C17220 net35 FILLER_0_22_86/a_1468_375# 0.010438f
C17221 mask\[8\] FILLER_0_22_86/a_36_472# 0.012471f
C17222 _008_ net61 0.004059f
C17223 FILLER_0_5_72/a_124_375# net47 0.006974f
C17224 FILLER_0_7_59/a_36_472# vss 0.004006f
C17225 FILLER_0_7_59/a_484_472# vdd 0.00824f
C17226 _081_ _080_ 0.003905f
C17227 _453_/a_36_151# vdd 0.164654f
C17228 FILLER_0_13_212/a_1468_375# _043_ 0.01418f
C17229 FILLER_0_5_109/a_124_375# net47 0.010784f
C17230 FILLER_0_15_116/a_36_472# _040_ 0.002896f
C17231 net35 FILLER_0_22_128/a_2276_472# 0.014483f
C17232 net82 net21 0.037271f
C17233 net22 _201_/a_67_603# 0.004491f
C17234 trim_mask\[2\] net17 0.084388f
C17235 _049_ _146_ 0.042698f
C17236 _164_ trim_mask\[3\] 0.016366f
C17237 FILLER_0_19_125/a_124_375# vss 0.001974f
C17238 FILLER_0_16_89/a_124_375# _136_ 0.011795f
C17239 FILLER_0_12_2/a_572_375# net67 0.007509f
C17240 _170_ vss 0.280383f
C17241 net68 FILLER_0_6_47/a_932_472# 0.014935f
C17242 FILLER_0_11_135/a_124_375# vdd 0.042201f
C17243 _000_ FILLER_0_3_221/a_1468_375# 0.054354f
C17244 net35 _211_/a_36_160# 0.009886f
C17245 FILLER_0_18_2/a_3260_375# net55 0.004262f
C17246 FILLER_0_10_214/a_36_472# _069_ 0.085701f
C17247 _098_ _437_/a_448_472# 0.050691f
C17248 FILLER_0_4_49/a_36_472# _167_ 0.063278f
C17249 _074_ vss 0.404343f
C17250 _119_ _162_ 0.036701f
C17251 FILLER_0_11_101/a_572_375# FILLER_0_9_105/a_36_472# 0.0027f
C17252 net55 FILLER_0_18_61/a_124_375# 0.040701f
C17253 _004_ _094_ 0.213913f
C17254 _412_/a_1000_472# net59 0.00147f
C17255 net73 _095_ 0.003688f
C17256 _448_/a_448_472# net59 0.050956f
C17257 _286_/a_224_472# vdd 0.00154f
C17258 net3 _185_ 0.004236f
C17259 FILLER_0_11_101/a_572_375# vdd 0.023482f
C17260 _127_ _125_ 0.053419f
C17261 _092_ _291_/a_36_160# 0.03297f
C17262 _068_ vdd 0.793549f
C17263 _076_ vss 1.132839f
C17264 _106_ _293_/a_36_472# 0.04279f
C17265 result[5] _094_ 0.065897f
C17266 net15 cal_count\[1\] 0.089855f
C17267 _105_ _098_ 0.055065f
C17268 FILLER_0_17_72/a_2724_472# _438_/a_36_151# 0.002529f
C17269 _052_ _424_/a_36_151# 0.010844f
C17270 _119_ _131_ 0.073868f
C17271 _429_/a_2665_112# FILLER_0_14_235/a_36_472# 0.007491f
C17272 FILLER_0_15_180/a_36_472# vss 0.00138f
C17273 FILLER_0_15_180/a_484_472# vdd 0.037927f
C17274 _132_ _040_ 0.023821f
C17275 mask\[1\] FILLER_0_15_180/a_124_375# 0.004011f
C17276 FILLER_0_4_99/a_124_375# _160_ 0.005563f
C17277 _105_ _205_/a_36_160# 0.001167f
C17278 _289_/a_36_472# _094_ 0.00922f
C17279 _116_ _120_ 0.005759f
C17280 FILLER_0_21_133/a_36_472# _436_/a_2248_156# 0.001148f
C17281 FILLER_0_16_89/a_1380_472# _131_ 0.004201f
C17282 net73 FILLER_0_18_139/a_484_472# 0.00131f
C17283 trim_mask\[2\] FILLER_0_3_78/a_484_472# 0.008122f
C17284 output39/a_224_472# _033_ 0.045759f
C17285 output34/a_224_472# _046_ 0.006059f
C17286 output32/a_224_472# net19 0.08441f
C17287 FILLER_0_20_177/a_36_472# FILLER_0_20_169/a_36_472# 0.002296f
C17288 vdd FILLER_0_13_72/a_572_375# -0.001166f
C17289 vss FILLER_0_13_72/a_124_375# 0.043492f
C17290 fanout51/a_36_113# vdd 0.013496f
C17291 net75 FILLER_0_8_263/a_36_472# 0.020293f
C17292 _274_/a_36_68# FILLER_0_12_220/a_484_472# 0.001048f
C17293 _028_ _439_/a_796_472# 0.013039f
C17294 _055_ _223_/a_36_160# 0.012271f
C17295 FILLER_0_19_142/a_124_375# _145_ 0.009109f
C17296 output42/a_224_472# net38 0.066219f
C17297 _420_/a_2560_156# _009_ 0.001487f
C17298 sample FILLER_0_9_290/a_124_375# 0.00195f
C17299 FILLER_0_20_169/a_124_375# vdd 0.03036f
C17300 net34 FILLER_0_22_177/a_1380_472# 0.003953f
C17301 _259_/a_455_68# net37 0.0023f
C17302 en_co_clk vss 0.014954f
C17303 fanout81/a_36_160# net82 0.027351f
C17304 _056_ _373_/a_244_68# 0.00229f
C17305 cal_count\[3\] _453_/a_1000_472# 0.001123f
C17306 net19 _001_ 0.018424f
C17307 _181_ cal_count\[2\] 0.375819f
C17308 _069_ _161_ 0.017831f
C17309 _095_ _451_/a_1040_527# 0.002316f
C17310 _118_ _120_ 0.339442f
C17311 FILLER_0_15_72/a_36_472# FILLER_0_15_59/a_484_472# 0.001963f
C17312 output31/a_224_472# net18 0.009938f
C17313 _189_/a_67_603# _100_ 0.002818f
C17314 FILLER_0_17_72/a_1828_472# net36 0.028046f
C17315 _343_/a_665_69# mask\[3\] 0.001405f
C17316 _303_/a_36_472# mask\[9\] 0.013976f
C17317 net52 FILLER_0_3_142/a_36_472# 0.001122f
C17318 net69 vdd 1.102677f
C17319 vdd _201_/a_67_603# 0.031337f
C17320 mask\[9\] _438_/a_1204_472# 0.03521f
C17321 net58 FILLER_0_9_270/a_484_472# 0.061043f
C17322 net27 FILLER_0_12_236/a_36_472# 0.005414f
C17323 _030_ _153_ 0.026157f
C17324 FILLER_0_5_164/a_484_472# vss 0.003257f
C17325 ctln[6] net23 0.003826f
C17326 _077_ _073_ 0.009611f
C17327 _308_/a_848_380# trim_mask\[0\] 0.035693f
C17328 result[5] net78 0.020038f
C17329 fanout78/a_36_113# _418_/a_36_151# 0.030244f
C17330 FILLER_0_16_89/a_124_375# net53 0.001032f
C17331 _077_ _330_/a_224_472# 0.001921f
C17332 net52 _442_/a_1308_423# 0.017208f
C17333 FILLER_0_18_177/a_932_472# vdd 0.029926f
C17334 FILLER_0_18_177/a_484_472# vss -0.001894f
C17335 _005_ _416_/a_36_151# 0.018752f
C17336 output8/a_224_472# FILLER_0_3_221/a_36_472# 0.001699f
C17337 _131_ _095_ 0.043211f
C17338 _427_/a_2665_112# net36 0.009904f
C17339 result[9] _419_/a_448_472# 0.015767f
C17340 net56 FILLER_0_16_154/a_1020_375# 0.002321f
C17341 _339_/a_36_160# FILLER_0_19_155/a_484_472# 0.00304f
C17342 _450_/a_2449_156# _039_ 0.013285f
C17343 _115_ FILLER_0_11_78/a_572_375# 0.034089f
C17344 net18 _419_/a_1000_472# 0.008295f
C17345 FILLER_0_19_28/a_124_375# _452_/a_36_151# 0.002709f
C17346 _360_/a_36_160# _070_ 0.012463f
C17347 net57 net52 0.016136f
C17348 net16 FILLER_0_18_37/a_1380_472# 0.002932f
C17349 net69 _441_/a_1204_472# 0.014374f
C17350 FILLER_0_17_104/a_1020_375# net14 0.002226f
C17351 net63 FILLER_0_19_195/a_124_375# 0.017284f
C17352 _216_/a_67_603# FILLER_0_18_61/a_124_375# 0.014522f
C17353 _425_/a_1000_472# vdd 0.019072f
C17354 _096_ _225_/a_36_160# 0.004807f
C17355 _077_ net15 0.238832f
C17356 _069_ _429_/a_448_472# 0.035108f
C17357 net37 FILLER_0_6_231/a_36_472# 0.002982f
C17358 _152_ vdd 0.354509f
C17359 _081_ vss 0.733408f
C17360 net35 net71 0.042275f
C17361 mask\[7\] FILLER_0_22_128/a_932_472# 0.017448f
C17362 _256_/a_1612_497# _055_ 0.001438f
C17363 _070_ _171_ 0.084342f
C17364 net34 ctlp[1] 0.127025f
C17365 FILLER_0_5_109/a_124_375# _154_ 0.058658f
C17366 net64 FILLER_0_9_270/a_36_472# 0.014971f
C17367 net53 _427_/a_1204_472# 0.004293f
C17368 ctln[7] vdd 0.359832f
C17369 _067_ FILLER_0_12_20/a_36_472# 0.015608f
C17370 _448_/a_1204_472# net22 0.002283f
C17371 _086_ vss 0.615299f
C17372 net15 FILLER_0_17_72/a_124_375# 0.006492f
C17373 _098_ FILLER_0_15_212/a_124_375# 0.008125f
C17374 FILLER_0_18_76/a_484_472# _438_/a_36_151# 0.001723f
C17375 net60 ctlp[1] 0.073021f
C17376 _099_ _098_ 0.018316f
C17377 net50 _439_/a_1000_472# 0.005154f
C17378 net52 _439_/a_2248_156# 0.00258f
C17379 _138_ vdd 0.090752f
C17380 net23 FILLER_0_8_156/a_36_472# 0.004939f
C17381 FILLER_0_4_49/a_36_472# vdd 0.090733f
C17382 FILLER_0_4_144/a_124_375# trim_mask\[4\] 0.014395f
C17383 FILLER_0_4_49/a_572_375# vss 0.008729f
C17384 net54 _438_/a_2248_156# 0.014423f
C17385 output11/a_224_472# net75 0.015211f
C17386 net65 vss 0.471168f
C17387 trim[0] output40/a_224_472# 0.005306f
C17388 FILLER_0_4_144/a_124_375# net47 0.012023f
C17389 net38 net40 1.103743f
C17390 output31/a_224_472# _417_/a_448_472# 0.008149f
C17391 _098_ FILLER_0_19_111/a_124_375# 0.001331f
C17392 net56 _095_ 0.004847f
C17393 _114_ _057_ 0.30288f
C17394 ctlp[9] net26 0.02213f
C17395 _136_ _337_/a_665_69# 0.001794f
C17396 _413_/a_1204_472# net21 0.011236f
C17397 _093_ FILLER_0_17_142/a_124_375# 0.009328f
C17398 _015_ FILLER_0_8_247/a_932_472# 0.005458f
C17399 _176_ FILLER_0_10_107/a_36_472# 0.009019f
C17400 _117_ _310_/a_49_472# 0.018229f
C17401 _053_ FILLER_0_7_72/a_2812_375# 0.016329f
C17402 FILLER_0_9_28/a_3172_472# net68 0.007929f
C17403 _132_ FILLER_0_14_107/a_484_472# 0.005391f
C17404 FILLER_0_22_86/a_1468_375# vdd 0.035441f
C17405 net15 _120_ 0.028275f
C17406 _308_/a_124_24# FILLER_0_9_72/a_1380_472# 0.003595f
C17407 net15 _038_ 0.078028f
C17408 net76 _037_ 0.010891f
C17409 FILLER_0_11_78/a_36_472# _120_ 0.014169f
C17410 _038_ FILLER_0_11_78/a_36_472# 0.001782f
C17411 net63 FILLER_0_18_177/a_1828_472# 0.047684f
C17412 _036_ fanout68/a_36_113# 0.007847f
C17413 FILLER_0_17_104/a_1380_472# FILLER_0_16_115/a_124_375# 0.001723f
C17414 mask\[4\] FILLER_0_19_171/a_572_375# 0.006277f
C17415 FILLER_0_5_212/a_124_375# FILLER_0_3_212/a_36_472# 0.001512f
C17416 _077_ net51 0.76967f
C17417 _095_ FILLER_0_13_80/a_36_472# 0.004187f
C17418 FILLER_0_22_128/a_2276_472# vdd 0.00565f
C17419 FILLER_0_22_128/a_1828_472# vss 0.009137f
C17420 FILLER_0_9_290/a_124_375# FILLER_0_9_282/a_572_375# 0.012001f
C17421 _075_ calibrate 0.022901f
C17422 FILLER_0_8_127/a_124_375# _129_ 0.056784f
C17423 _119_ _074_ 0.153267f
C17424 net27 _426_/a_2248_156# 0.002303f
C17425 mask\[5\] FILLER_0_19_187/a_484_472# 0.007596f
C17426 net56 FILLER_0_18_139/a_484_472# 0.004375f
C17427 fanout59/a_36_160# net59 0.021522f
C17428 net80 _019_ 0.265857f
C17429 _430_/a_2665_112# _092_ 0.004778f
C17430 _143_ FILLER_0_18_171/a_124_375# 0.005331f
C17431 _053_ _151_ 0.538643f
C17432 _211_/a_36_160# vdd 0.030216f
C17433 FILLER_0_15_235/a_124_375# FILLER_0_14_235/a_124_375# 0.05841f
C17434 output32/a_224_472# _419_/a_448_472# 0.010723f
C17435 _094_ net19 0.06304f
C17436 net63 FILLER_0_17_218/a_572_375# 0.006355f
C17437 _425_/a_2248_156# net19 0.010557f
C17438 _013_ vdd 0.372605f
C17439 net41 _052_ 0.001927f
C17440 _445_/a_1308_423# _034_ 0.002494f
C17441 trimb[3] net17 0.005798f
C17442 mask\[4\] _346_/a_49_472# 0.079347f
C17443 net58 calibrate 0.205792f
C17444 _137_ _097_ 0.001654f
C17445 _119_ _076_ 0.083673f
C17446 net66 net40 0.124825f
C17447 net17 output6/a_224_472# 0.047757f
C17448 _185_ _402_/a_56_567# 0.107713f
C17449 net82 FILLER_0_3_172/a_484_472# 0.008052f
C17450 _075_ net21 0.012335f
C17451 net36 FILLER_0_18_76/a_572_375# 0.005153f
C17452 FILLER_0_14_50/a_124_375# _179_ 0.021823f
C17453 net54 mask\[8\] 0.162104f
C17454 _067_ FILLER_0_12_28/a_36_472# 0.0127f
C17455 _093_ FILLER_0_18_107/a_932_472# 0.008683f
C17456 _067_ net40 0.040115f
C17457 _093_ _110_ 0.08348f
C17458 _132_ _334_/a_36_160# 0.026495f
C17459 FILLER_0_3_172/a_3260_375# net65 0.002696f
C17460 _322_/a_124_24# net74 0.05722f
C17461 FILLER_0_4_177/a_484_472# _087_ 0.005486f
C17462 _255_/a_224_552# _374_/a_36_68# 0.00191f
C17463 ctlp[2] mask\[7\] 0.036719f
C17464 _432_/a_2665_112# vss 0.002577f
C17465 _069_ _056_ 0.035189f
C17466 fanout70/a_36_113# net36 0.007807f
C17467 FILLER_0_15_142/a_36_472# net36 0.015456f
C17468 FILLER_0_15_116/a_484_472# vss 0.003923f
C17469 _443_/a_1308_423# vdd 0.00203f
C17470 _443_/a_448_472# vss 0.030448f
C17471 _020_ _431_/a_796_472# 0.012284f
C17472 _412_/a_2248_156# fanout59/a_36_160# 0.007753f
C17473 _120_ net51 1.716752f
C17474 fanout76/a_36_160# net65 0.018025f
C17475 output48/a_224_472# _425_/a_448_472# 0.001155f
C17476 FILLER_0_9_28/a_2812_375# vdd 0.016637f
C17477 _448_/a_1204_472# vdd 0.002228f
C17478 net52 FILLER_0_6_47/a_2276_472# 0.003298f
C17479 calibrate net21 0.036773f
C17480 net15 mask\[8\] 0.02403f
C17481 result[4] _418_/a_36_151# 0.005556f
C17482 net12 net59 0.001028f
C17483 _090_ vss 0.267577f
C17484 _137_ mask\[2\] 0.440828f
C17485 _113_ vdd 0.774039f
C17486 _131_ _332_/a_36_472# 0.006825f
C17487 _425_/a_36_151# FILLER_0_8_247/a_572_375# 0.001597f
C17488 _392_/a_244_472# _067_ 0.001893f
C17489 FILLER_0_16_57/a_1020_375# net72 0.002937f
C17490 output48/a_224_472# _082_ 0.002393f
C17491 output37/a_224_472# net18 0.046654f
C17492 net15 FILLER_0_17_56/a_484_472# 0.001758f
C17493 _041_ FILLER_0_18_37/a_1380_472# 0.003776f
C17494 FILLER_0_5_54/a_36_472# net47 0.00679f
C17495 net68 _453_/a_448_472# 0.01245f
C17496 fanout59/a_36_160# net64 0.006298f
C17497 net57 _428_/a_1308_423# 0.018725f
C17498 FILLER_0_3_54/a_124_375# net40 0.005766f
C17499 output48/a_224_472# net82 0.048965f
C17500 _092_ FILLER_0_18_209/a_572_375# 0.00609f
C17501 net78 _108_ 0.056528f
C17502 _433_/a_2560_156# _145_ 0.007651f
C17503 FILLER_0_17_56/a_124_375# _041_ 0.001489f
C17504 net74 _372_/a_786_69# 0.00149f
C17505 _016_ FILLER_0_12_136/a_572_375# 0.00332f
C17506 net78 net19 0.507249f
C17507 FILLER_0_7_195/a_36_472# _414_/a_36_151# 0.001723f
C17508 _308_/a_124_24# vdd 0.011014f
C17509 _069_ _068_ 0.003779f
C17510 _053_ FILLER_0_8_37/a_484_472# 0.002095f
C17511 _000_ net8 0.021422f
C17512 FILLER_0_17_72/a_3260_375# vdd 0.007427f
C17513 _134_ FILLER_0_10_107/a_124_375# 0.009573f
C17514 FILLER_0_12_20/a_484_472# net47 0.020293f
C17515 _136_ FILLER_0_17_142/a_124_375# 0.001315f
C17516 cal_itt\[3\] _087_ 0.002881f
C17517 FILLER_0_8_263/a_36_472# net19 0.047387f
C17518 net3 net17 0.045911f
C17519 _132_ FILLER_0_18_107/a_1468_375# 0.089207f
C17520 FILLER_0_4_107/a_1380_472# vdd 0.007022f
C17521 vdd FILLER_0_6_37/a_124_375# 0.041381f
C17522 FILLER_0_5_72/a_484_472# FILLER_0_6_47/a_3260_375# 0.001597f
C17523 net15 _175_ 0.052586f
C17524 _415_/a_448_472# result[1] 0.005209f
C17525 _142_ FILLER_0_17_133/a_124_375# 0.022066f
C17526 _427_/a_448_472# vss 0.040679f
C17527 _427_/a_1308_423# vdd 0.002814f
C17528 trim_mask\[4\] _370_/a_848_380# 0.027744f
C17529 net72 FILLER_0_15_59/a_36_472# 0.049812f
C17530 net52 FILLER_0_2_111/a_484_472# 0.061249f
C17531 _029_ vss 0.11129f
C17532 _043_ FILLER_0_13_72/a_36_472# 0.017766f
C17533 ctlp[2] _422_/a_2248_156# 0.001328f
C17534 cal_count\[3\] _405_/a_67_603# 0.011131f
C17535 _370_/a_848_380# net47 0.004223f
C17536 _093_ net14 0.11038f
C17537 FILLER_0_2_101/a_124_375# _154_ 0.003932f
C17538 net58 fanout81/a_36_160# 0.013959f
C17539 trim_mask\[2\] FILLER_0_2_93/a_36_472# 0.281054f
C17540 _415_/a_2248_156# vdd 0.009114f
C17541 _053_ _162_ 0.00209f
C17542 _091_ FILLER_0_15_212/a_1468_375# 0.002531f
C17543 net52 _440_/a_1204_472# 0.003916f
C17544 _449_/a_36_151# _453_/a_36_151# 0.007757f
C17545 net60 _421_/a_2560_156# 0.001951f
C17546 vss _145_ 0.399701f
C17547 mask\[3\] FILLER_0_18_177/a_1916_375# 0.003052f
C17548 net5 net59 0.923076f
C17549 _291_/a_36_160# _199_/a_36_160# 0.005575f
C17550 _256_/a_36_68# calibrate 0.02084f
C17551 FILLER_0_8_107/a_36_472# vss 0.006371f
C17552 output34/a_224_472# _103_ 0.027876f
C17553 _091_ FILLER_0_16_154/a_1380_472# 0.00133f
C17554 _452_/a_448_472# _041_ 0.007f
C17555 _114_ _307_/a_672_472# 0.0018f
C17556 _091_ mask\[3\] 0.044304f
C17557 _119_ _086_ 0.419383f
C17558 _178_ _408_/a_56_524# 0.014421f
C17559 net71 vdd 0.775031f
C17560 net49 _440_/a_1204_472# 0.006692f
C17561 output39/a_224_472# _444_/a_36_151# 0.062717f
C17562 _086_ _071_ 0.041029f
C17563 _021_ vss 0.142648f
C17564 _053_ _131_ 0.086215f
C17565 net38 FILLER_0_15_2/a_484_472# 0.003391f
C17566 _235_/a_67_603# _064_ 0.003796f
C17567 en_co_clk _095_ 0.003753f
C17568 _350_/a_49_472# mask\[6\] 0.033488f
C17569 _035_ _164_ 0.056332f
C17570 FILLER_0_9_28/a_484_472# net40 0.020293f
C17571 _447_/a_1204_472# vdd 0.001085f
C17572 net57 FILLER_0_8_156/a_36_472# 0.001544f
C17573 _077_ FILLER_0_10_78/a_572_375# 0.001886f
C17574 _324_/a_224_472# _129_ 0.009728f
C17575 FILLER_0_24_96/a_36_472# ctlp[7] 0.001551f
C17576 net23 FILLER_0_22_128/a_2364_375# 0.018463f
C17577 FILLER_0_17_64/a_36_472# net36 0.00195f
C17578 _137_ FILLER_0_16_154/a_484_472# 0.00631f
C17579 _183_ _180_ 0.002621f
C17580 _412_/a_2248_156# net5 0.048919f
C17581 _314_/a_224_472# vss 0.001399f
C17582 _447_/a_2665_112# _168_ 0.001107f
C17583 FILLER_0_5_72/a_36_472# _440_/a_36_151# 0.001723f
C17584 _164_ FILLER_0_6_47/a_3172_472# 0.001058f
C17585 FILLER_0_10_78/a_484_472# _439_/a_36_151# 0.00271f
C17586 net54 _433_/a_2248_156# 0.04755f
C17587 FILLER_0_0_198/a_36_472# vss 0.00344f
C17588 _105_ ctlp[2] 0.223601f
C17589 fanout60/a_36_160# net79 0.069956f
C17590 net15 _453_/a_2560_156# 0.049334f
C17591 mask\[7\] net21 0.050718f
C17592 FILLER_0_21_125/a_36_472# _433_/a_36_151# 0.001723f
C17593 _363_/a_244_472# _053_ 0.001236f
C17594 FILLER_0_14_81/a_36_472# _394_/a_1936_472# 0.010394f
C17595 net74 _370_/a_848_380# 0.004546f
C17596 _365_/a_244_472# _156_ 0.003847f
C17597 _016_ _428_/a_448_472# 0.00347f
C17598 net41 net40 2.687418f
C17599 _444_/a_1000_472# _054_ 0.002998f
C17600 _411_/a_2665_112# net8 0.036782f
C17601 result[5] _418_/a_2248_156# 0.001309f
C17602 FILLER_0_20_107/a_36_472# FILLER_0_20_98/a_36_472# 0.001963f
C17603 FILLER_0_18_2/a_3172_472# _452_/a_36_151# 0.059367f
C17604 FILLER_0_18_2/a_2724_472# _452_/a_448_472# 0.008967f
C17605 _345_/a_36_160# net73 0.032139f
C17606 output47/a_224_472# FILLER_0_15_10/a_36_472# 0.038484f
C17607 net64 net5 0.098088f
C17608 FILLER_0_8_24/a_484_472# _054_ 0.009315f
C17609 _449_/a_36_151# FILLER_0_13_72/a_572_375# 0.035849f
C17610 _059_ FILLER_0_5_136/a_36_472# 0.001755f
C17611 _410_/a_36_68# _039_ 0.016062f
C17612 cal_count\[1\] FILLER_0_15_59/a_484_472# 0.006408f
C17613 _008_ _093_ 0.252609f
C17614 net65 FILLER_0_2_177/a_36_472# 0.016652f
C17615 _125_ _118_ 0.239695f
C17616 _354_/a_49_472# _098_ 0.009677f
C17617 _029_ FILLER_0_5_88/a_124_375# 0.006771f
C17618 net16 cal_count\[3\] 0.082821f
C17619 _103_ _418_/a_36_151# 0.032388f
C17620 FILLER_0_10_78/a_572_375# _120_ 0.006134f
C17621 _176_ cal_count\[3\] 0.067683f
C17622 _025_ _436_/a_2248_156# 0.001054f
C17623 _076_ _385_/a_36_68# 0.006512f
C17624 _414_/a_36_151# vss 0.002101f
C17625 _091_ FILLER_0_12_220/a_484_472# 0.001453f
C17626 ctlp[1] FILLER_0_23_290/a_124_375# 0.053745f
C17627 mask\[4\] net63 0.043339f
C17628 _078_ net37 0.459092f
C17629 net31 _201_/a_67_603# 0.015773f
C17630 FILLER_0_5_128/a_484_472# vss 0.004051f
C17631 net33 _434_/a_448_472# 0.003049f
C17632 net64 FILLER_0_15_235/a_484_472# 0.005893f
C17633 _141_ _093_ 0.396041f
C17634 _102_ net36 0.003446f
C17635 trim_mask\[2\] FILLER_0_4_91/a_124_375# 0.003591f
C17636 _444_/a_1204_472# vdd 0.001086f
C17637 _091_ _323_/a_36_113# 0.001651f
C17638 FILLER_0_7_233/a_36_472# vss 0.005354f
C17639 net7 output16/a_224_472# 0.001321f
C17640 FILLER_0_0_232/a_36_472# vdd 0.050082f
C17641 FILLER_0_0_232/a_124_375# vss 0.019863f
C17642 FILLER_0_16_73/a_124_375# FILLER_0_17_72/a_124_375# 0.026339f
C17643 FILLER_0_21_142/a_124_375# _433_/a_2560_156# 0.001178f
C17644 _088_ _269_/a_36_472# 0.004438f
C17645 net78 _419_/a_448_472# 0.0122f
C17646 net81 net1 0.03613f
C17647 net54 FILLER_0_18_107/a_124_375# 0.001636f
C17648 _219_/a_36_160# net14 0.048037f
C17649 _136_ net14 0.417108f
C17650 net11 vss 0.057193f
C17651 _453_/a_2560_156# net51 0.013556f
C17652 mask\[1\] net21 0.023956f
C17653 _440_/a_2665_112# _164_ 0.067034f
C17654 _375_/a_36_68# _162_ 0.011065f
C17655 _375_/a_1612_497# _161_ 0.003325f
C17656 _163_ vss 0.638066f
C17657 net38 _452_/a_1040_527# 0.002024f
C17658 FILLER_0_4_49/a_484_472# net68 0.027016f
C17659 FILLER_0_20_2/a_124_375# net43 0.001563f
C17660 _010_ _420_/a_2665_112# 0.029378f
C17661 _438_/a_1000_472# net14 0.003275f
C17662 _412_/a_2665_112# cal_itt\[1\] 0.015571f
C17663 FILLER_0_21_28/a_572_375# vdd 0.013051f
C17664 _451_/a_1697_156# net14 0.001298f
C17665 output15/a_224_472# vss 0.067969f
C17666 FILLER_0_14_91/a_36_472# en_co_clk 0.007733f
C17667 FILLER_0_11_78/a_572_375# vdd -0.006646f
C17668 FILLER_0_11_78/a_124_375# vss 0.006233f
C17669 FILLER_0_13_65/a_124_375# FILLER_0_13_72/a_36_472# 0.012267f
C17670 FILLER_0_15_72/a_484_472# _451_/a_3129_107# 0.005866f
C17671 fanout74/a_36_113# _371_/a_36_113# 0.01088f
C17672 _412_/a_1308_423# net58 0.037719f
C17673 FILLER_0_0_96/a_36_472# trim_mask\[3\] 0.005343f
C17674 net82 FILLER_0_4_213/a_124_375# 0.00123f
C17675 _064_ vdd 0.874293f
C17676 FILLER_0_6_239/a_36_472# _123_ 0.004433f
C17677 _053_ _220_/a_67_603# 0.065611f
C17678 net67 FILLER_0_9_60/a_124_375# 0.003083f
C17679 FILLER_0_22_86/a_36_472# _026_ 0.001503f
C17680 FILLER_0_22_86/a_932_472# _149_ 0.001205f
C17681 _253_/a_1732_68# cal_itt\[1\] 0.001829f
C17682 _131_ FILLER_0_11_124/a_36_472# 0.015445f
C17683 net63 _435_/a_36_151# 0.017194f
C17684 ctlp[4] _009_ 0.004522f
C17685 _058_ _062_ 1.676625f
C17686 FILLER_0_21_142/a_124_375# vss 0.009345f
C17687 _093_ FILLER_0_17_104/a_572_375# 0.01418f
C17688 output39/a_224_472# _054_ 0.002121f
C17689 net39 _221_/a_36_160# 0.059979f
C17690 FILLER_0_4_107/a_124_375# net47 0.004586f
C17691 _053_ FILLER_0_7_59/a_36_472# 0.073877f
C17692 mask\[5\] FILLER_0_19_195/a_36_472# 0.007596f
C17693 net15 _441_/a_1000_472# 0.025912f
C17694 FILLER_0_6_90/a_124_375# vdd 0.020992f
C17695 _371_/a_36_113# FILLER_0_2_127/a_124_375# 0.002437f
C17696 net42 vdd 0.178782f
C17697 output29/a_224_472# _005_ 0.021351f
C17698 net73 _098_ 0.004745f
C17699 _418_/a_796_472# vss 0.00145f
C17700 _256_/a_244_497# _128_ 0.002372f
C17701 FILLER_0_13_212/a_1468_375# FILLER_0_13_228/a_124_375# 0.012001f
C17702 FILLER_0_10_28/a_36_472# net51 0.00703f
C17703 _172_ FILLER_0_10_94/a_124_375# 0.003341f
C17704 _171_ FILLER_0_10_94/a_36_472# 0.001514f
C17705 FILLER_0_22_177/a_932_472# net33 0.014021f
C17706 _433_/a_1204_472# _022_ 0.005308f
C17707 _426_/a_2248_156# _076_ 0.015189f
C17708 FILLER_0_18_2/a_1020_375# net38 0.047331f
C17709 _053_ _074_ 0.503728f
C17710 net52 FILLER_0_9_72/a_1020_375# 0.00799f
C17711 FILLER_0_21_286/a_484_472# vss 0.008522f
C17712 FILLER_0_15_116/a_484_472# _095_ 0.001069f
C17713 net81 FILLER_0_15_235/a_124_375# 0.008139f
C17714 FILLER_0_13_142/a_572_375# net23 0.009573f
C17715 FILLER_0_4_99/a_36_472# FILLER_0_4_107/a_36_472# 0.002296f
C17716 net58 output48/a_224_472# 0.065357f
C17717 _057_ _310_/a_741_69# 0.001002f
C17718 FILLER_0_19_187/a_484_472# _434_/a_2665_112# 0.001868f
C17719 FILLER_0_1_266/a_36_472# vdd 0.008551f
C17720 FILLER_0_1_266/a_572_375# vss 0.001919f
C17721 ctln[2] net82 0.005498f
C17722 _069_ _113_ 0.027402f
C17723 _079_ _112_ 0.004464f
C17724 _042_ vdd 0.261947f
C17725 _117_ vss 0.048946f
C17726 _081_ _385_/a_36_68# 0.006303f
C17727 _331_/a_448_472# _134_ 0.001126f
C17728 _092_ _276_/a_36_160# 0.06772f
C17729 fanout56/a_36_113# _097_ 0.062226f
C17730 output9/a_224_472# _412_/a_448_472# 0.001025f
C17731 FILLER_0_5_206/a_36_472# vss 0.003493f
C17732 _053_ _076_ 0.108358f
C17733 _077_ net74 0.025882f
C17734 FILLER_0_15_150/a_36_472# net56 0.011741f
C17735 _273_/a_36_68# _128_ 0.005719f
C17736 FILLER_0_18_2/a_36_472# net44 0.011079f
C17737 FILLER_0_18_2/a_932_472# vdd 0.002342f
C17738 FILLER_0_18_2/a_484_472# vss 0.001228f
C17739 FILLER_0_17_226/a_124_375# vss 0.025007f
C17740 _114_ _161_ 0.024297f
C17741 _328_/a_36_113# net74 0.002214f
C17742 _428_/a_2665_112# _131_ 0.006081f
C17743 result[5] fanout60/a_36_160# 0.001585f
C17744 output48/a_224_472# calibrate 0.003223f
C17745 _093_ FILLER_0_19_134/a_36_472# 0.002415f
C17746 _132_ _126_ 0.247838f
C17747 _176_ FILLER_0_17_72/a_1828_472# 0.001028f
C17748 _431_/a_2560_156# _137_ 0.002967f
C17749 net53 net14 0.04525f
C17750 output37/a_224_472# net65 0.096416f
C17751 net82 FILLER_0_3_221/a_572_375# 0.005424f
C17752 mask\[5\] FILLER_0_18_177/a_2276_472# 0.001063f
C17753 net46 FILLER_0_21_28/a_124_375# 0.011995f
C17754 ctln[1] net82 0.001141f
C17755 vdd FILLER_0_4_91/a_484_472# 0.007304f
C17756 result[8] ctlp[2] 0.068359f
C17757 output25/a_224_472# net35 0.016177f
C17758 input2/a_36_113# clk 0.021981f
C17759 FILLER_0_8_247/a_124_375# calibrate 0.008393f
C17760 FILLER_0_12_220/a_124_375# _090_ 0.001521f
C17761 ctlp[1] FILLER_0_24_274/a_484_472# 0.001875f
C17762 net1 net2 0.624657f
C17763 FILLER_0_13_212/a_572_375# _070_ 0.003986f
C17764 FILLER_0_3_172/a_1828_472# net22 0.009883f
C17765 FILLER_0_5_212/a_124_375# vdd 0.024541f
C17766 FILLER_0_8_37/a_572_375# _220_/a_67_603# 0.00744f
C17767 FILLER_0_12_136/a_484_472# _127_ 0.005549f
C17768 _143_ FILLER_0_16_154/a_1468_375# 0.002033f
C17769 _422_/a_2248_156# mask\[7\] 0.015008f
C17770 _071_ _314_/a_224_472# 0.001359f
C17771 output36/a_224_472# net30 0.083671f
C17772 _116_ _043_ 0.002037f
C17773 _104_ _199_/a_36_160# 0.095519f
C17774 FILLER_0_10_214/a_124_375# _070_ 0.017713f
C17775 output30/a_224_472# result[3] 0.019025f
C17776 output38/a_224_472# vdd -0.006652f
C17777 net74 _120_ 0.027885f
C17778 net74 _038_ 0.055774f
C17779 _427_/a_448_472# _095_ 0.063616f
C17780 result[9] _009_ 0.19745f
C17781 net75 FILLER_0_8_247/a_484_472# 0.003007f
C17782 net32 vss 0.824307f
C17783 FILLER_0_16_37/a_124_375# _179_ 0.005434f
C17784 mask\[0\] net21 0.050431f
C17785 _446_/a_36_151# trim[3] 0.00699f
C17786 net16 _408_/a_2215_68# 0.002096f
C17787 FILLER_0_9_223/a_124_375# _128_ 0.004252f
C17788 _321_/a_170_472# _126_ 0.018831f
C17789 _408_/a_718_524# _043_ 0.003719f
C17790 FILLER_0_16_73/a_124_375# _175_ 0.005727f
C17791 _066_ _386_/a_848_380# 0.00416f
C17792 output24/a_224_472# ctlp[7] 0.060657f
C17793 fanout52/a_36_160# trim_mask\[4\] 0.014356f
C17794 FILLER_0_16_73/a_36_472# _131_ 0.008223f
C17795 FILLER_0_5_198/a_484_472# net59 0.059394f
C17796 FILLER_0_15_142/a_572_375# _427_/a_36_151# 0.059049f
C17797 ctlp[7] vss 0.036681f
C17798 FILLER_0_1_266/a_36_472# net9 0.041635f
C17799 FILLER_0_5_54/a_484_472# FILLER_0_6_47/a_1380_472# 0.026657f
C17800 FILLER_0_5_54/a_1468_375# FILLER_0_6_47/a_2276_472# 0.001597f
C17801 _428_/a_448_472# _017_ 0.056f
C17802 _428_/a_36_151# net53 0.001124f
C17803 fanout53/a_36_160# net56 0.196684f
C17804 _369_/a_36_68# vdd 0.042534f
C17805 FILLER_0_16_57/a_484_472# FILLER_0_17_56/a_572_375# 0.001723f
C17806 _044_ vdd 0.406979f
C17807 _274_/a_36_68# _072_ 0.001647f
C17808 _192_/a_67_603# _044_ 0.002571f
C17809 comp vss 0.148428f
C17810 _408_/a_56_524# _095_ 0.01643f
C17811 FILLER_0_20_169/a_124_375# _140_ 0.01799f
C17812 _177_ cal_count\[1\] 0.03631f
C17813 net76 _123_ 0.003431f
C17814 _144_ _346_/a_49_472# 0.036821f
C17815 FILLER_0_2_177/a_484_472# net59 0.007829f
C17816 FILLER_0_11_142/a_484_472# vdd 0.006641f
C17817 FILLER_0_11_142/a_36_472# vss 0.008744f
C17818 FILLER_0_12_136/a_1380_472# _076_ 0.001809f
C17819 _322_/a_1152_472# _129_ 0.002978f
C17820 FILLER_0_18_107/a_2812_375# vss 0.002392f
C17821 FILLER_0_18_107/a_3260_375# vdd 0.004983f
C17822 _073_ net76 0.040554f
C17823 _434_/a_1308_423# mask\[6\] 0.022677f
C17824 state\[1\] _121_ 0.006184f
C17825 FILLER_0_7_104/a_1468_375# vdd 0.026224f
C17826 FILLER_0_16_73/a_484_472# _040_ 0.004877f
C17827 _105_ mask\[7\] 0.486236f
C17828 _432_/a_2248_156# net80 0.059406f
C17829 _173_ _120_ 0.004205f
C17830 FILLER_0_18_139/a_484_472# _145_ 0.002415f
C17831 FILLER_0_3_221/a_36_472# FILLER_0_3_212/a_36_472# 0.001963f
C17832 net79 FILLER_0_12_220/a_1380_472# 0.010583f
C17833 net47 _386_/a_692_472# 0.003299f
C17834 output29/a_224_472# _416_/a_448_472# 0.008149f
C17835 _074_ _375_/a_36_68# 0.003157f
C17836 FILLER_0_7_162/a_36_472# vss 0.006392f
C17837 valid net1 0.00347f
C17838 _119_ _163_ 0.009297f
C17839 trim_val\[4\] _386_/a_1084_68# 0.002659f
C17840 net55 FILLER_0_21_60/a_572_375# 0.041903f
C17841 _053_ _081_ 0.698311f
C17842 fanout78/a_36_113# _007_ 0.003126f
C17843 trim_val\[1\] FILLER_0_6_47/a_36_472# 0.00351f
C17844 FILLER_0_16_57/a_1468_375# _175_ 0.001654f
C17845 net52 _441_/a_36_151# 0.013755f
C17846 net32 _107_ 0.003155f
C17847 FILLER_0_4_107/a_124_375# _154_ 0.00183f
C17848 _447_/a_1000_472# _036_ 0.002902f
C17849 net54 _150_ 0.001162f
C17850 FILLER_0_23_88/a_36_472# vss 0.003481f
C17851 _133_ _160_ 0.043549f
C17852 FILLER_0_19_125/a_124_375# _345_/a_36_160# 0.005398f
C17853 net24 _050_ 0.049889f
C17854 _122_ FILLER_0_5_198/a_484_472# 0.002999f
C17855 _346_/a_49_472# net23 0.022558f
C17856 _030_ _384_/a_224_472# 0.003019f
C17857 _086_ _053_ 0.091538f
C17858 _417_/a_1308_423# output30/a_224_472# 0.001434f
C17859 _417_/a_36_151# net30 0.010021f
C17860 net47 _452_/a_836_156# 0.002075f
C17861 input5/a_36_113# rstn 0.019149f
C17862 output34/a_224_472# _419_/a_2665_112# 0.010731f
C17863 FILLER_0_5_117/a_124_375# _158_ 0.001068f
C17864 _062_ _226_/a_860_68# 0.001842f
C17865 _091_ FILLER_0_13_212/a_36_472# 0.007355f
C17866 _072_ _375_/a_960_497# 0.001322f
C17867 _441_/a_448_472# _030_ 0.038429f
C17868 _441_/a_36_151# net49 0.010951f
C17869 _208_/a_36_160# _049_ 0.04568f
C17870 net75 _411_/a_1308_423# 0.028281f
C17871 FILLER_0_7_72/a_124_375# _028_ 0.017052f
C17872 net64 _055_ 0.00384f
C17873 net15 _423_/a_2665_112# 0.061217f
C17874 _437_/a_1000_472# vdd 0.001777f
C17875 result[7] FILLER_0_24_274/a_572_375# 0.006125f
C17876 _428_/a_36_151# FILLER_0_14_107/a_124_375# 0.001597f
C17877 cal_itt\[3\] _061_ 0.001311f
C17878 _449_/a_2665_112# _038_ 0.024406f
C17879 FILLER_0_18_177/a_1468_375# FILLER_0_19_187/a_484_472# 0.001684f
C17880 FILLER_0_3_172/a_1828_472# vdd 0.0083f
C17881 _131_ _070_ 0.161861f
C17882 _096_ _306_/a_36_68# 0.016266f
C17883 FILLER_0_7_104/a_932_472# _058_ 0.002096f
C17884 FILLER_0_5_109/a_124_375# _365_/a_36_68# 0.004633f
C17885 _052_ net36 0.005689f
C17886 _065_ _235_/a_67_603# 0.004135f
C17887 FILLER_0_19_171/a_36_472# _434_/a_36_151# 0.00271f
C17888 _052_ FILLER_0_18_37/a_932_472# 0.002749f
C17889 fanout75/a_36_113# _082_ 0.016843f
C17890 output9/a_224_472# input4/a_36_68# 0.009732f
C17891 FILLER_0_12_50/a_36_472# _453_/a_36_151# 0.001748f
C17892 _144_ _352_/a_257_69# 0.001662f
C17893 _077_ _439_/a_1204_472# 0.016471f
C17894 _132_ _436_/a_36_151# 0.00162f
C17895 _144_ _433_/a_1204_472# 0.009472f
C17896 state\[2\] net74 0.024462f
C17897 mask\[2\] FILLER_0_15_235/a_484_472# 0.004683f
C17898 FILLER_0_9_223/a_484_472# _076_ 0.001736f
C17899 _114_ _056_ 0.034246f
C17900 vss net6 0.096009f
C17901 result[8] net21 0.166555f
C17902 fanout82/a_36_113# _425_/a_36_151# 0.030783f
C17903 FILLER_0_23_88/a_124_375# _437_/a_36_151# 0.002709f
C17904 FILLER_0_22_177/a_1380_472# mask\[6\] 0.006573f
C17905 net35 FILLER_0_22_177/a_932_472# 0.00643f
C17906 _098_ _048_ 0.092201f
C17907 mask\[9\] FILLER_0_18_76/a_484_472# 0.002672f
C17908 _130_ _129_ 0.021732f
C17909 ctlp[1] FILLER_0_23_282/a_124_375# 0.00324f
C17910 ctln[8] ctln[9] 0.003265f
C17911 net15 _043_ 0.042278f
C17912 mask\[3\] net22 0.036607f
C17913 _431_/a_1308_423# _020_ 0.001997f
C17914 FILLER_0_14_181/a_124_375# vdd 0.040138f
C17915 net57 FILLER_0_13_142/a_572_375# 0.011369f
C17916 _172_ vss 0.054608f
C17917 net55 _131_ 0.314732f
C17918 net81 net76 0.236554f
C17919 net54 _026_ 0.006401f
C17920 cal_itt\[3\] _072_ 2.019868f
C17921 _205_/a_36_160# _048_ 0.040317f
C17922 net48 vss 0.161385f
C17923 _140_ FILLER_0_22_128/a_2276_472# 0.002954f
C17924 FILLER_0_17_200/a_572_375# net21 0.011557f
C17925 _188_ _067_ 0.001554f
C17926 _383_/a_36_472# vdd -0.002154f
C17927 mask\[4\] FILLER_0_18_209/a_36_472# 0.018888f
C17928 _219_/a_36_160# _439_/a_2665_112# 0.002537f
C17929 FILLER_0_8_247/a_1468_375# vdd 0.011086f
C17930 _114_ FILLER_0_11_101/a_572_375# 0.051108f
C17931 _085_ _267_/a_672_472# 0.006682f
C17932 _116_ _267_/a_1568_472# 0.001147f
C17933 _114_ _068_ 1.097353f
C17934 _421_/a_2665_112# net33 0.007127f
C17935 _415_/a_796_472# _004_ 0.005395f
C17936 net55 FILLER_0_18_37/a_572_375# 0.007169f
C17937 net72 FILLER_0_18_37/a_36_472# 0.043427f
C17938 _092_ _293_/a_36_472# 0.004828f
C17939 FILLER_0_12_136/a_572_375# cal_count\[3\] 0.005006f
C17940 mask\[0\] mask\[1\] 0.01742f
C17941 net76 FILLER_0_5_212/a_36_472# 0.00377f
C17942 net15 net68 0.205016f
C17943 FILLER_0_9_28/a_932_472# vdd 0.04397f
C17944 FILLER_0_9_223/a_36_472# _273_/a_36_68# 0.015795f
C17945 net34 _199_/a_36_160# 0.026709f
C17946 _414_/a_2665_112# net59 0.010265f
C17947 net47 _221_/a_36_160# 0.012197f
C17948 output25/a_224_472# vdd 0.03413f
C17949 _441_/a_1308_423# _164_ 0.001807f
C17950 FILLER_0_7_72/a_2724_472# _219_/a_36_160# 0.001448f
C17951 state\[1\] FILLER_0_13_142/a_1380_472# 0.006475f
C17952 ctln[2] net58 0.025352f
C17953 _290_/a_224_472# _094_ 0.003006f
C17954 FILLER_0_3_221/a_124_375# net59 0.008996f
C17955 _058_ net14 0.40635f
C17956 FILLER_0_4_99/a_124_375# FILLER_0_4_91/a_572_375# 0.012001f
C17957 FILLER_0_10_28/a_36_472# net47 0.002783f
C17958 _013_ _424_/a_2665_112# 0.001222f
C17959 net38 _450_/a_36_151# 0.035458f
C17960 _420_/a_2560_156# vdd 0.001652f
C17961 _011_ _422_/a_36_151# 0.015698f
C17962 _420_/a_2665_112# vss 0.001749f
C17963 _412_/a_1204_472# net81 0.003435f
C17964 _086_ _375_/a_36_68# 0.038443f
C17965 ctlp[4] net33 0.001734f
C17966 FILLER_0_16_241/a_124_375# net36 0.004069f
C17967 _018_ FILLER_0_15_205/a_36_472# 0.00273f
C17968 _276_/a_36_160# FILLER_0_17_218/a_36_472# 0.035111f
C17969 output26/a_224_472# FILLER_0_23_44/a_484_472# 0.0323f
C17970 vss FILLER_0_16_115/a_36_472# 0.003243f
C17971 _399_/a_224_472# _182_ 0.002729f
C17972 _098_ FILLER_0_15_180/a_36_472# 0.101593f
C17973 cal_count\[1\] _451_/a_2225_156# 0.006336f
C17974 _444_/a_2248_156# net67 0.028782f
C17975 FILLER_0_4_197/a_1020_375# net22 0.040565f
C17976 result[1] net64 0.048458f
C17977 FILLER_0_21_125/a_484_472# net54 0.022347f
C17978 net52 _443_/a_2248_156# 0.045316f
C17979 _086_ FILLER_0_11_124/a_36_472# 0.010729f
C17980 FILLER_0_2_93/a_572_375# _367_/a_36_68# 0.001069f
C17981 net41 FILLER_0_10_28/a_124_375# 0.003909f
C17982 mask\[9\] FILLER_0_20_107/a_36_472# 0.006047f
C17983 FILLER_0_16_57/a_572_375# vss 0.00372f
C17984 FILLER_0_16_57/a_1020_375# vdd 0.004428f
C17985 ctln[1] net58 0.014147f
C17986 vdd _450_/a_2449_156# 0.003646f
C17987 FILLER_0_16_37/a_36_472# _402_/a_728_93# 0.0108f
C17988 _387_/a_36_113# _170_ 0.017801f
C17989 net35 _436_/a_1000_472# 0.009213f
C17990 FILLER_0_4_123/a_124_375# _070_ 0.001677f
C17991 net55 FILLER_0_13_80/a_36_472# 0.016536f
C17992 _020_ _093_ 0.015474f
C17993 _062_ _134_ 0.024038f
C17994 _322_/a_1152_472# _068_ 0.001502f
C17995 _265_/a_244_68# _001_ 0.008874f
C17996 result[8] mask\[7\] 0.110637f
C17997 trimb[0] FILLER_0_20_2/a_36_472# 0.005458f
C17998 _183_ vss 0.009822f
C17999 _065_ vdd 0.646511f
C18000 _374_/a_244_472# _076_ 0.001567f
C18001 FILLER_0_15_212/a_1020_375# vss 0.035883f
C18002 FILLER_0_15_212/a_1468_375# vdd 0.010445f
C18003 FILLER_0_15_212/a_124_375# mask\[1\] 0.007876f
C18004 _414_/a_2665_112# _122_ 0.007441f
C18005 net68 net51 0.008885f
C18006 _099_ mask\[1\] 0.19135f
C18007 _063_ trim_mask\[1\] 0.127216f
C18008 _093_ _438_/a_796_472# 0.001924f
C18009 _316_/a_1084_68# net37 0.001574f
C18010 net16 _233_/a_36_160# 0.01152f
C18011 _141_ _343_/a_49_472# 0.04106f
C18012 FILLER_0_7_72/a_1916_375# vdd 0.015888f
C18013 _363_/a_36_68# _154_ 0.149319f
C18014 FILLER_0_20_177/a_932_472# _434_/a_36_151# 0.001723f
C18015 output7/a_224_472# ctln[9] 0.001987f
C18016 FILLER_0_16_154/a_932_472# vss 0.001652f
C18017 FILLER_0_16_154/a_1380_472# vdd 0.001901f
C18018 mask\[3\] vdd 0.340612f
C18019 net57 _386_/a_848_380# 0.041622f
C18020 net15 net67 0.109181f
C18021 net64 FILLER_0_12_236/a_484_472# 0.010321f
C18022 fanout68/a_36_113# net17 0.001252f
C18023 _119_ FILLER_0_7_162/a_36_472# 0.005739f
C18024 net27 FILLER_0_9_270/a_484_472# 0.023461f
C18025 trim_mask\[1\] FILLER_0_6_47/a_1468_375# 0.007169f
C18026 FILLER_0_19_111/a_484_472# vdd 0.009246f
C18027 net20 FILLER_0_15_212/a_1468_375# 0.006824f
C18028 net62 FILLER_0_15_282/a_124_375# 0.012711f
C18029 _434_/a_36_151# vss 0.006401f
C18030 _434_/a_448_472# vdd 0.020387f
C18031 _148_ _352_/a_49_472# 0.003082f
C18032 output8/a_224_472# output11/a_224_472# 0.003437f
C18033 FILLER_0_21_133/a_124_375# vdd 0.010519f
C18034 _411_/a_2560_156# net75 0.007047f
C18035 _000_ _073_ 0.222349f
C18036 _074_ _070_ 0.102481f
C18037 _053_ FILLER_0_8_107/a_36_472# 0.013669f
C18038 _163_ _385_/a_36_68# 0.012699f
C18039 mask\[3\] net20 0.047107f
C18040 FILLER_0_15_59/a_572_375# vss 0.018573f
C18041 FILLER_0_15_59/a_36_472# vdd 0.031071f
C18042 net76 net2 0.039533f
C18043 net15 FILLER_0_11_64/a_36_472# 0.020589f
C18044 _080_ net37 0.005467f
C18045 FILLER_0_19_47/a_484_472# net55 0.061087f
C18046 FILLER_0_11_101/a_124_375# _070_ 0.052406f
C18047 _260_/a_36_68# FILLER_0_3_221/a_1380_472# 0.001652f
C18048 _270_/a_36_472# net21 0.001606f
C18049 _070_ _076_ 0.198272f
C18050 mask\[7\] FILLER_0_22_177/a_1468_375# 0.001315f
C18051 fanout69/a_36_113# vss 0.002239f
C18052 net35 FILLER_0_22_128/a_124_375# 0.010439f
C18053 _430_/a_2248_156# mask\[3\] 0.004211f
C18054 trim_val\[4\] FILLER_0_3_172/a_36_472# 0.006208f
C18055 net76 FILLER_0_3_172/a_2276_472# 0.002531f
C18056 _162_ _312_/a_234_472# 0.003812f
C18057 FILLER_0_7_146/a_36_472# _076_ 0.001843f
C18058 FILLER_0_7_146/a_124_375# _068_ 0.033245f
C18059 net50 trim_mask\[1\] 0.502622f
C18060 state\[0\] net4 0.13193f
C18061 FILLER_0_13_65/a_124_375# net15 0.048002f
C18062 FILLER_0_22_128/a_2724_472# FILLER_0_21_150/a_124_375# 0.001543f
C18063 FILLER_0_24_96/a_124_375# ctlp[7] 0.004486f
C18064 result[9] FILLER_0_24_274/a_932_472# 0.001826f
C18065 _064_ _445_/a_1308_423# 0.01485f
C18066 net52 _176_ 0.004215f
C18067 net41 FILLER_0_20_31/a_36_472# 0.030033f
C18068 cal vss 0.424638f
C18069 FILLER_0_13_212/a_932_472# net79 0.006824f
C18070 _130_ FILLER_0_11_135/a_124_375# 0.001198f
C18071 net62 FILLER_0_13_212/a_1380_472# 0.059367f
C18072 ctln[2] clk 0.004558f
C18073 _140_ net71 0.005182f
C18074 _069_ FILLER_0_11_142/a_484_472# 0.005789f
C18075 net39 net67 0.049482f
C18076 net4 FILLER_0_3_221/a_1380_472# 0.003953f
C18077 FILLER_0_13_206/a_36_472# net22 0.053292f
C18078 net16 net49 0.055931f
C18079 _431_/a_36_151# FILLER_0_14_123/a_124_375# 0.002807f
C18080 net67 net51 0.010753f
C18081 FILLER_0_15_205/a_36_472# vss 0.003239f
C18082 FILLER_0_15_116/a_572_375# _131_ 0.051323f
C18083 net63 FILLER_0_15_212/a_484_472# 0.059367f
C18084 _450_/a_448_472# clkc 0.003011f
C18085 _450_/a_1040_527# net6 0.019715f
C18086 output47/a_224_472# _452_/a_2225_156# 0.012077f
C18087 _003_ _079_ 0.035497f
C18088 _089_ _088_ 0.009863f
C18089 _084_ _316_/a_124_24# 0.001501f
C18090 _372_/a_170_472# vdd 0.031606f
C18091 _181_ _180_ 0.216908f
C18092 ctln[2] fanout81/a_36_160# 0.003798f
C18093 FILLER_0_4_197/a_1020_375# vdd 0.002455f
C18094 ctlp[9] vss 0.013018f
C18095 FILLER_0_12_220/a_484_472# vdd 0.002383f
C18096 FILLER_0_12_220/a_36_472# vss 0.023702f
C18097 FILLER_0_11_64/a_36_472# net51 0.009015f
C18098 _142_ FILLER_0_18_107/a_2724_472# 0.001549f
C18099 net50 _447_/a_2665_112# 0.015374f
C18100 _363_/a_692_472# _086_ 0.001353f
C18101 _058_ FILLER_0_8_156/a_124_375# 0.006325f
C18102 ctln[1] clk 0.551557f
C18103 _087_ net22 0.028009f
C18104 net74 _125_ 0.071757f
C18105 _186_ _067_ 0.001907f
C18106 FILLER_0_17_200/a_36_472# vdd 0.001039f
C18107 _074_ FILLER_0_5_164/a_572_375# 0.001307f
C18108 _323_/a_36_113# vdd 0.009958f
C18109 net78 _009_ 0.02395f
C18110 net58 fanout58/a_36_160# 0.013794f
C18111 net39 _445_/a_448_472# 0.014537f
C18112 net27 net58 0.190417f
C18113 FILLER_0_5_72/a_36_472# _029_ 0.007282f
C18114 FILLER_0_5_72/a_572_375# trim_mask\[1\] 0.010714f
C18115 FILLER_0_22_177/a_484_472# vss -0.001894f
C18116 FILLER_0_22_177/a_932_472# vdd 0.029547f
C18117 valid net76 0.285892f
C18118 net20 FILLER_0_12_220/a_484_472# 0.001758f
C18119 _053_ _414_/a_36_151# 0.035994f
C18120 _020_ _136_ 0.022753f
C18121 FILLER_0_16_89/a_1468_375# net14 0.022582f
C18122 FILLER_0_21_125/a_36_472# _022_ 0.002295f
C18123 FILLER_0_18_139/a_36_472# FILLER_0_18_107/a_3260_375# 0.086905f
C18124 net7 net41 0.243942f
C18125 net75 cal_itt\[0\] 0.032053f
C18126 _426_/a_2665_112# net64 0.01548f
C18127 _046_ net30 0.006105f
C18128 mask\[2\] FILLER_0_16_154/a_1468_375# 0.014254f
C18129 _079_ net1 0.099822f
C18130 _063_ _444_/a_2665_112# 0.001996f
C18131 _028_ net15 0.223301f
C18132 _452_/a_36_151# net40 0.012138f
C18133 FILLER_0_4_107/a_484_472# _160_ 0.008194f
C18134 FILLER_0_4_213/a_484_472# vdd 0.007084f
C18135 FILLER_0_4_213/a_36_472# vss 0.003969f
C18136 _070_ FILLER_0_5_164/a_484_472# 0.003424f
C18137 _341_/a_49_472# mask\[2\] 0.026222f
C18138 FILLER_0_16_107/a_124_375# _131_ 0.016011f
C18139 _016_ net53 0.180698f
C18140 _086_ _374_/a_244_472# 0.001496f
C18141 net20 _323_/a_36_113# 0.002161f
C18142 FILLER_0_14_99/a_124_375# FILLER_0_14_107/a_36_472# 0.009654f
C18143 FILLER_0_21_142/a_572_375# _433_/a_2665_112# 0.001092f
C18144 _128_ _247_/a_36_160# 0.00163f
C18145 _091_ _274_/a_2960_68# 0.001338f
C18146 FILLER_0_18_2/a_3172_472# _041_ 0.001503f
C18147 FILLER_0_17_72/a_1916_375# _131_ 0.006589f
C18148 net27 calibrate 0.017426f
C18149 _415_/a_796_472# net19 0.001468f
C18150 _411_/a_2665_112# _073_ 0.009313f
C18151 net55 FILLER_0_13_72/a_124_375# 0.00281f
C18152 net80 _435_/a_448_472# 0.005274f
C18153 _105_ result[8] 0.011678f
C18154 _449_/a_2248_156# vdd -0.001225f
C18155 _449_/a_1204_472# vss 0.006048f
C18156 cal_count\[2\] net47 0.274891f
C18157 net26 _423_/a_36_151# 0.067024f
C18158 net53 FILLER_0_14_123/a_124_375# 0.003138f
C18159 _103_ _007_ 0.002514f
C18160 _053_ _163_ 0.763235f
C18161 net27 FILLER_0_10_256/a_124_375# 0.006216f
C18162 net82 _170_ 0.080348f
C18163 net28 _044_ 0.481924f
C18164 _091_ _072_ 0.162027f
C18165 mask\[0\] _099_ 0.00418f
C18166 _028_ FILLER_0_6_90/a_572_375# 0.015802f
C18167 fanout64/a_36_160# net65 0.214347f
C18168 _149_ _437_/a_2665_112# 0.020763f
C18169 _026_ _437_/a_1204_472# 0.022954f
C18170 FILLER_0_1_266/a_124_375# FILLER_0_0_266/a_124_375# 0.05841f
C18171 vss trim[3] 0.235724f
C18172 _074_ _082_ 0.069835f
C18173 _070_ _081_ 0.00804f
C18174 _451_/a_836_156# _040_ 0.016371f
C18175 _074_ net82 0.123449f
C18176 _414_/a_2248_156# vss 0.00384f
C18177 _430_/a_36_151# net36 0.003701f
C18178 _020_ _431_/a_36_151# 0.023081f
C18179 _442_/a_36_151# vdd 0.102701f
C18180 FILLER_0_14_181/a_36_472# _043_ 0.008613f
C18181 net34 _435_/a_448_472# 0.013341f
C18182 net27 _415_/a_1000_472# 0.017938f
C18183 net38 _445_/a_36_151# 0.112205f
C18184 net50 _444_/a_2665_112# 0.023342f
C18185 net15 FILLER_0_6_47/a_1916_375# 0.029774f
C18186 net25 _423_/a_2248_156# 0.005535f
C18187 _176_ FILLER_0_15_72/a_572_375# 0.005529f
C18188 _073_ FILLER_0_6_231/a_36_472# 0.001898f
C18189 _086_ _070_ 0.123033f
C18190 _114_ _113_ 0.201729f
C18191 net47 _450_/a_448_472# 0.012172f
C18192 _345_/a_36_160# _145_ 0.001141f
C18193 _305_/a_36_159# vdd 0.017293f
C18194 FILLER_0_21_142/a_572_375# vdd 0.002442f
C18195 fanout62/a_36_160# FILLER_0_11_282/a_36_472# 0.005262f
C18196 _028_ net51 0.002321f
C18197 FILLER_0_19_47/a_124_375# _013_ 0.023766f
C18198 net1 cal_itt\[1\] 0.229522f
C18199 _408_/a_56_524# _185_ 0.002484f
C18200 FILLER_0_13_206/a_36_472# vdd 0.011681f
C18201 FILLER_0_19_155/a_572_375# vdd 0.01384f
C18202 FILLER_0_19_155/a_124_375# vss 0.00336f
C18203 FILLER_0_13_206/a_124_375# vss 0.051723f
C18204 sample vss 0.276162f
C18205 _328_/a_36_113# net70 0.00292f
C18206 _137_ FILLER_0_15_180/a_484_472# 0.046411f
C18207 FILLER_0_18_2/a_1916_375# trimb[1] 0.001855f
C18208 FILLER_0_7_104/a_932_472# _134_ 0.004249f
C18209 net37 vss 0.666835f
C18210 trim[4] net42 0.016428f
C18211 net18 FILLER_0_9_270/a_484_472# 0.004375f
C18212 _445_/a_2560_156# vdd 0.002586f
C18213 _445_/a_2665_112# vss 0.004455f
C18214 FILLER_0_21_28/a_3172_472# vss 0.001574f
C18215 _436_/a_1000_472# vdd 0.006522f
C18216 FILLER_0_3_221/a_36_472# vdd 0.018263f
C18217 FILLER_0_3_221/a_1468_375# vss 0.004085f
C18218 _114_ _308_/a_124_24# 0.052818f
C18219 _423_/a_2665_112# _012_ 0.014394f
C18220 _432_/a_36_151# _093_ 0.018324f
C18221 FILLER_0_10_78/a_1468_375# _389_/a_36_148# 0.001699f
C18222 _303_/a_36_472# net36 0.006675f
C18223 net76 FILLER_0_5_172/a_124_375# 0.001526f
C18224 net36 _438_/a_1204_472# 0.012234f
C18225 FILLER_0_16_107/a_572_375# _040_ 0.001244f
C18226 _439_/a_796_472# vss 0.003859f
C18227 _149_ net14 0.102004f
C18228 FILLER_0_19_171/a_1468_375# FILLER_0_19_187/a_36_472# 0.086743f
C18229 net62 _429_/a_2248_156# 0.012262f
C18230 _087_ vdd 0.281159f
C18231 _105_ _204_/a_255_603# 0.002146f
C18232 _258_/a_36_160# net76 0.015203f
C18233 output47/a_224_472# net44 0.077292f
C18234 FILLER_0_10_78/a_932_472# _439_/a_2665_112# 0.001182f
C18235 net15 _424_/a_2248_156# 0.00415f
C18236 _445_/a_36_151# net66 0.058093f
C18237 FILLER_0_5_109/a_484_472# _363_/a_36_68# 0.001709f
C18238 _096_ vdd 0.557569f
C18239 net79 _193_/a_36_160# 0.010228f
C18240 FILLER_0_13_212/a_36_472# net22 0.002402f
C18241 FILLER_0_5_128/a_124_375# vdd 0.008803f
C18242 FILLER_0_10_37/a_36_472# FILLER_0_10_28/a_36_472# 0.001963f
C18243 FILLER_0_14_99/a_36_472# vdd 0.095251f
C18244 FILLER_0_14_99/a_124_375# vss 0.017196f
C18245 _008_ _419_/a_36_151# 0.014476f
C18246 mask\[3\] FILLER_0_16_154/a_572_375# 0.027873f
C18247 _043_ net47 0.043824f
C18248 net44 FILLER_0_12_2/a_124_375# 0.01836f
C18249 net50 FILLER_0_6_90/a_36_472# 0.049285f
C18250 FILLER_0_12_2/a_36_472# vdd 0.104425f
C18251 FILLER_0_12_2/a_572_375# vss 0.017629f
C18252 _122_ _160_ 0.004488f
C18253 _077_ FILLER_0_9_72/a_572_375# 0.008103f
C18254 _074_ _312_/a_234_472# 0.005755f
C18255 _162_ calibrate 0.228839f
C18256 FILLER_0_16_57/a_1380_472# _176_ 0.01346f
C18257 FILLER_0_10_37/a_124_375# vdd 0.048346f
C18258 ctln[1] input2/a_36_113# 0.05197f
C18259 result[4] net30 0.298966f
C18260 _091_ FILLER_0_17_218/a_572_375# 0.001927f
C18261 _448_/a_36_151# _037_ 0.012725f
C18262 _120_ FILLER_0_10_107/a_124_375# 0.001834f
C18263 net67 clkc 0.102244f
C18264 _105_ output18/a_224_472# 0.105478f
C18265 FILLER_0_8_127/a_36_472# vss 0.004344f
C18266 _077_ _453_/a_796_472# 0.003409f
C18267 FILLER_0_22_128/a_124_375# vdd 0.013058f
C18268 trimb[1] vdd 0.225206f
C18269 _217_/a_36_160# FILLER_0_19_28/a_572_375# 0.058908f
C18270 _058_ _439_/a_2665_112# 0.001029f
C18271 _139_ vss 0.052996f
C18272 _413_/a_1308_423# net59 0.018948f
C18273 valid fanout65/a_36_113# 0.001646f
C18274 trimb[1] FILLER_0_20_15/a_484_472# 0.001292f
C18275 FILLER_0_4_123/a_36_472# FILLER_0_4_107/a_1468_375# 0.086635f
C18276 ctlp[4] net22 0.257841f
C18277 net68 net47 0.063835f
C18278 _098_ _145_ 0.007514f
C18279 net41 _186_ 0.054661f
C18280 net69 FILLER_0_3_78/a_36_472# 0.002068f
C18281 FILLER_0_9_142/a_124_375# _120_ 0.04442f
C18282 FILLER_0_8_138/a_124_375# _058_ 0.009863f
C18283 net60 _418_/a_2665_112# 0.042307f
C18284 net69 FILLER_0_2_127/a_36_472# 0.019383f
C18285 _072_ _306_/a_36_68# 0.042843f
C18286 _057_ _055_ 0.290639f
C18287 mask\[3\] _069_ 0.025564f
C18288 state\[1\] _097_ 0.004171f
C18289 _134_ net14 0.001303f
C18290 net58 net18 0.091503f
C18291 _410_/a_36_68# vdd 0.039824f
C18292 _081_ _082_ 0.008298f
C18293 _028_ FILLER_0_7_104/a_36_472# 0.006408f
C18294 net64 _223_/a_36_160# 0.007842f
C18295 _070_ _090_ 0.369847f
C18296 trimb[2] vss 0.102375f
C18297 FILLER_0_0_130/a_124_375# net13 0.009149f
C18298 output14/a_224_472# ctln[7] 0.076006f
C18299 _397_/a_36_472# FILLER_0_17_72/a_1020_375# 0.001781f
C18300 net62 _248_/a_36_68# 0.002178f
C18301 _021_ _098_ 0.014179f
C18302 trim_val\[2\] _160_ 0.051804f
C18303 net54 FILLER_0_21_150/a_124_375# 0.007123f
C18304 result[0] FILLER_0_9_282/a_484_472# 0.018647f
C18305 _144_ FILLER_0_21_125/a_36_472# 0.008287f
C18306 net62 _417_/a_2665_112# 0.006083f
C18307 net47 _156_ 0.040298f
C18308 calibrate net18 0.014127f
C18309 net74 _043_ 0.65119f
C18310 _137_ _138_ 0.045916f
C18311 FILLER_0_6_47/a_1380_472# vdd 0.002735f
C18312 FILLER_0_9_282/a_36_472# vdd 0.106034f
C18313 FILLER_0_9_282/a_572_375# vss 0.058599f
C18314 _093_ FILLER_0_18_177/a_3172_472# 0.003708f
C18315 _013_ _182_ 0.001681f
C18316 _429_/a_36_151# net21 0.054289f
C18317 net82 net65 0.630327f
C18318 _255_/a_224_552# _057_ 0.024333f
C18319 _057_ _126_ 0.022413f
C18320 mask\[8\] FILLER_0_22_107/a_484_472# 0.024416f
C18321 net35 FILLER_0_22_107/a_36_472# 0.007196f
C18322 _432_/a_36_151# _136_ 0.004543f
C18323 net56 fanout54/a_36_160# 0.044466f
C18324 net16 _052_ 0.022236f
C18325 _193_/a_36_160# FILLER_0_13_290/a_124_375# 0.005732f
C18326 _053_ FILLER_0_7_104/a_1020_375# 0.002671f
C18327 result[4] _417_/a_36_151# 0.010571f
C18328 fanout57/a_36_113# net65 0.035361f
C18329 net32 _421_/a_1308_423# 0.005394f
C18330 _104_ _011_ 0.021454f
C18331 _053_ FILLER_0_7_162/a_36_472# 0.004888f
C18332 _322_/a_692_472# _118_ 0.002849f
C18333 _415_/a_1000_472# net18 0.006558f
C18334 FILLER_0_13_212/a_1468_375# vss 0.062822f
C18335 FILLER_0_13_212/a_36_472# vdd 0.105926f
C18336 output43/a_224_472# trimb[2] 0.005445f
C18337 _238_/a_67_603# FILLER_0_2_93/a_36_472# 0.002778f
C18338 ctlp[1] _420_/a_448_472# 0.038053f
C18339 net67 net47 0.126281f
C18340 cal_count\[3\] FILLER_0_12_28/a_124_375# 0.013328f
C18341 _421_/a_2665_112# vdd 0.029293f
C18342 FILLER_0_20_177/a_1380_472# FILLER_0_19_187/a_124_375# 0.001543f
C18343 _446_/a_1000_472# net17 0.031119f
C18344 net19 cal_itt\[0\] 0.111163f
C18345 _072_ _395_/a_36_488# 0.024944f
C18346 ctln[3] _411_/a_2248_156# 0.001208f
C18347 net75 FILLER_0_10_247/a_36_472# 0.001184f
C18348 net62 _005_ 0.097739f
C18349 _238_/a_67_603# trim_mask\[2\] 0.003021f
C18350 FILLER_0_8_107/a_36_472# _070_ 0.001287f
C18351 FILLER_0_8_107/a_124_375# _133_ 0.048874f
C18352 FILLER_0_19_187/a_36_472# vdd 0.09884f
C18353 FILLER_0_19_187/a_572_375# vss 0.055266f
C18354 vss FILLER_0_21_60/a_484_472# 0.004134f
C18355 ctln[5] output12/a_224_472# 0.069673f
C18356 net73 FILLER_0_18_107/a_1916_375# 0.014643f
C18357 _094_ FILLER_0_17_282/a_124_375# 0.001151f
C18358 FILLER_0_5_117/a_36_472# vdd 0.092171f
C18359 output35/a_224_472# FILLER_0_22_177/a_1380_472# 0.002486f
C18360 FILLER_0_2_111/a_1468_375# vdd 0.011806f
C18361 ctln[1] _411_/a_1204_472# 0.031348f
C18362 _429_/a_796_472# net22 0.020124f
C18363 net10 output11/a_224_472# 0.095679f
C18364 _431_/a_2665_112# FILLER_0_17_142/a_124_375# 0.004834f
C18365 trim_mask\[2\] fanout68/a_36_113# 0.003509f
C18366 FILLER_0_4_91/a_572_375# _160_ 0.007391f
C18367 net15 _394_/a_728_93# 0.085551f
C18368 net50 net66 0.016385f
C18369 net52 _030_ 0.035783f
C18370 _187_ _188_ 0.001453f
C18371 FILLER_0_11_109/a_36_472# _134_ 0.007739f
C18372 _445_/a_448_472# net47 0.005429f
C18373 ctlp[4] vdd 0.278868f
C18374 _440_/a_1308_423# vss 0.028595f
C18375 FILLER_0_8_138/a_36_472# _313_/a_67_603# 0.005759f
C18376 _149_ _148_ 0.001124f
C18377 output36/a_224_472# _006_ 0.022685f
C18378 FILLER_0_16_107/a_484_472# FILLER_0_14_107/a_572_375# 0.001404f
C18379 net66 _382_/a_224_472# 0.001902f
C18380 _379_/a_36_472# _164_ 0.026812f
C18381 net18 _418_/a_448_472# 0.026048f
C18382 _104_ _008_ 0.135471f
C18383 output26/a_224_472# ctlp[9] 0.034572f
C18384 _075_ _074_ 0.058521f
C18385 _006_ net30 0.284414f
C18386 _077_ _319_/a_672_472# 0.001602f
C18387 _077_ FILLER_0_9_60/a_36_472# 0.038809f
C18388 _030_ net49 0.046089f
C18389 clk net18 0.003519f
C18390 _313_/a_67_603# vdd -0.002183f
C18391 _390_/a_36_68# vss 0.002334f
C18392 net82 _443_/a_448_472# 0.007335f
C18393 _412_/a_448_472# vdd 0.011f
C18394 trimb[0] output45/a_224_472# 0.003753f
C18395 _431_/a_448_472# _132_ 0.003024f
C18396 _004_ FILLER_0_10_247/a_36_472# 0.001551f
C18397 _415_/a_448_472# net64 0.02484f
C18398 net70 FILLER_0_14_107/a_1020_375# 0.011157f
C18399 net44 FILLER_0_20_2/a_124_375# 0.001564f
C18400 _079_ net76 2.404004f
C18401 FILLER_0_20_2/a_572_375# vss 0.001471f
C18402 FILLER_0_20_2/a_36_472# vdd 0.102471f
C18403 output22/a_224_472# mask\[7\] 0.05527f
C18404 _103_ net30 0.013544f
C18405 _430_/a_36_151# FILLER_0_18_177/a_2724_472# 0.001512f
C18406 net58 _074_ 0.004651f
C18407 FILLER_0_5_54/a_484_472# trim_mask\[1\] 0.013584f
C18408 fanout62/a_36_160# vdd 0.059299f
C18409 _438_/a_36_151# vdd 0.111691f
C18410 ctlp[1] _419_/a_1308_423# 0.00678f
C18411 net25 net24 0.031854f
C18412 _405_/a_67_603# net40 0.015326f
C18413 _451_/a_3129_107# vdd 0.008569f
C18414 _137_ _113_ 0.030279f
C18415 _062_ FILLER_0_8_156/a_484_472# 0.006123f
C18416 FILLER_0_5_198/a_36_472# net37 0.0114f
C18417 _369_/a_244_472# _160_ 0.00146f
C18418 _294_/a_224_472# net20 0.008053f
C18419 _053_ net48 0.003159f
C18420 _074_ calibrate 0.046632f
C18421 FILLER_0_21_142/a_124_375# _098_ 0.006558f
C18422 _370_/a_848_380# FILLER_0_5_136/a_124_375# 0.014613f
C18423 net4 _248_/a_36_68# 0.054512f
C18424 net50 FILLER_0_3_54/a_124_375# 0.00189f
C18425 _442_/a_2665_112# _157_ 0.001587f
C18426 _079_ FILLER_0_5_198/a_124_375# 0.013896f
C18427 _095_ _402_/a_718_527# 0.002109f
C18428 _033_ FILLER_0_6_37/a_36_472# 0.017695f
C18429 _236_/a_36_160# vdd 0.023428f
C18430 _164_ FILLER_0_6_47/a_1020_375# 0.004285f
C18431 FILLER_0_18_2/a_1468_375# output44/a_224_472# 0.032639f
C18432 mask\[4\] FILLER_0_18_177/a_1916_375# 0.013466f
C18433 _076_ calibrate 1.005804f
C18434 _069_ FILLER_0_13_206/a_36_472# 0.005793f
C18435 _119_ FILLER_0_8_127/a_36_472# 0.053962f
C18436 _074_ net21 0.186175f
C18437 _447_/a_448_472# net69 0.001694f
C18438 net16 _165_ 0.021744f
C18439 _070_ FILLER_0_7_233/a_36_472# 0.07194f
C18440 _073_ _078_ 0.098575f
C18441 FILLER_0_13_65/a_124_375# net74 0.020091f
C18442 _154_ _156_ 0.019471f
C18443 _091_ mask\[4\] 0.071954f
C18444 _408_/a_56_524# net17 0.048018f
C18445 _177_ _150_ 0.002507f
C18446 mask\[5\] _141_ 0.241158f
C18447 net76 cal_itt\[1\] 0.027781f
C18448 _418_/a_1308_423# _417_/a_36_151# 0.001518f
C18449 net27 mask\[0\] 0.067038f
C18450 FILLER_0_17_226/a_36_472# vss 0.007552f
C18451 _417_/a_36_151# _006_ 0.015561f
C18452 _076_ net21 0.031683f
C18453 FILLER_0_7_104/a_124_375# _131_ 0.001291f
C18454 FILLER_0_9_28/a_36_472# net42 0.038355f
C18455 _052_ FILLER_0_21_28/a_2364_375# 0.002388f
C18456 fanout80/a_36_113# _136_ 0.006151f
C18457 _070_ _163_ 1.884485f
C18458 FILLER_0_18_37/a_1468_375# vss 0.054381f
C18459 FILLER_0_18_37/a_36_472# vdd 0.136723f
C18460 _061_ net22 0.123662f
C18461 _093_ FILLER_0_16_89/a_1020_375# 0.004133f
C18462 _333_/a_36_160# FILLER_0_15_180/a_36_472# 0.016014f
C18463 _429_/a_1308_423# vss 0.008906f
C18464 _429_/a_36_151# mask\[1\] 0.001021f
C18465 net52 trim_mask\[3\] 0.666362f
C18466 _057_ state\[1\] 0.284428f
C18467 _000_ _253_/a_36_68# 0.005121f
C18468 _317_/a_36_113# FILLER_0_7_233/a_124_375# 0.03227f
C18469 result[9] vdd 0.597071f
C18470 _331_/a_448_472# _120_ 0.001496f
C18471 _307_/a_672_472# _126_ 0.00121f
C18472 cal_count\[3\] _136_ 0.00703f
C18473 net8 vss 0.171128f
C18474 net79 _416_/a_36_151# 0.062626f
C18475 ctlp[5] net22 0.001542f
C18476 output46/a_224_472# FILLER_0_20_2/a_484_472# 0.001699f
C18477 _044_ output30/a_224_472# 0.00717f
C18478 net62 _416_/a_448_472# 0.009111f
C18479 net49 trim_mask\[3\] 0.03723f
C18480 FILLER_0_5_72/a_1380_472# FILLER_0_5_88/a_36_472# 0.013277f
C18481 FILLER_0_5_117/a_124_375# FILLER_0_5_109/a_572_375# 0.012001f
C18482 FILLER_0_9_28/a_3172_472# vss 0.001977f
C18483 _093_ FILLER_0_17_72/a_1828_472# 0.053526f
C18484 _413_/a_1204_472# net65 0.017514f
C18485 _196_/a_36_160# mask\[1\] 0.003254f
C18486 FILLER_0_3_2/a_36_472# net66 0.011419f
C18487 net41 _063_ 0.105528f
C18488 FILLER_0_14_99/a_124_375# _095_ 0.012128f
C18489 net20 result[9] 1.593573f
C18490 FILLER_0_7_195/a_124_375# _072_ 0.012244f
C18491 net38 _039_ 0.059899f
C18492 net16 net40 0.039189f
C18493 _147_ _434_/a_36_151# 0.001817f
C18494 _075_ _081_ 0.001195f
C18495 output41/a_224_472# trim[3] 0.042209f
C18496 FILLER_0_15_235/a_124_375# FILLER_0_15_228/a_124_375# 0.002868f
C18497 _412_/a_1204_472# cal_itt\[1\] 0.001547f
C18498 _122_ FILLER_0_5_164/a_36_472# 0.002232f
C18499 _310_/a_49_472# _060_ 0.001122f
C18500 net52 net13 0.018118f
C18501 vdd FILLER_0_22_107/a_36_472# 0.114332f
C18502 vss FILLER_0_22_107/a_572_375# 0.001944f
C18503 output8/a_224_472# _411_/a_1308_423# 0.005111f
C18504 output44/a_224_472# FILLER_0_20_15/a_36_472# 0.0323f
C18505 _141_ FILLER_0_17_142/a_484_472# 0.004527f
C18506 _423_/a_36_151# FILLER_0_23_60/a_36_472# 0.001723f
C18507 _104_ FILLER_0_23_274/a_124_375# 0.002159f
C18508 _181_ vss 0.003673f
C18509 _285_/a_36_472# vdd 0.073338f
C18510 _072_ net22 0.147672f
C18511 _132_ FILLER_0_15_116/a_36_472# 0.020589f
C18512 _178_ _181_ 0.188669f
C18513 _321_/a_170_472# _121_ 0.007364f
C18514 net60 _011_ 0.003094f
C18515 FILLER_0_10_37/a_36_472# net68 0.005405f
C18516 fanout49/a_36_160# FILLER_0_4_91/a_36_472# 0.001461f
C18517 net72 FILLER_0_21_28/a_1468_375# 0.001823f
C18518 net55 FILLER_0_11_78/a_124_375# 0.001597f
C18519 _256_/a_36_68# _076_ 0.079206f
C18520 net16 FILLER_0_17_38/a_572_375# 0.018281f
C18521 _272_/a_36_472# vdd 0.058326f
C18522 FILLER_0_5_164/a_572_375# _163_ 0.046852f
C18523 FILLER_0_5_164/a_36_472# _169_ 0.00284f
C18524 input4/a_36_68# vdd 0.09828f
C18525 _068_ _311_/a_3740_473# 0.001409f
C18526 _070_ _117_ 0.080445f
C18527 fanout66/a_36_113# vdd 0.049012f
C18528 _444_/a_1000_472# net17 0.02064f
C18529 net63 net36 0.010544f
C18530 net36 net19 0.031858f
C18531 FILLER_0_2_93/a_572_375# net69 0.015032f
C18532 ctlp[6] _050_ 0.100418f
C18533 net15 FILLER_0_5_54/a_932_472# 0.008904f
C18534 net41 net50 0.002438f
C18535 _425_/a_796_472# calibrate 0.025807f
C18536 _187_ _186_ 0.032149f
C18537 mask\[3\] _282_/a_36_160# 0.005823f
C18538 FILLER_0_8_24/a_484_472# net17 0.010321f
C18539 net58 net65 1.468105f
C18540 _140_ _434_/a_448_472# 0.00128f
C18541 _141_ net80 0.077957f
C18542 _424_/a_2248_156# _012_ 0.009377f
C18543 _023_ vss 0.114191f
C18544 _033_ _444_/a_2248_156# 0.011578f
C18545 _273_/a_36_68# _246_/a_36_68# 0.001168f
C18546 FILLER_0_21_133/a_124_375# _140_ 0.018383f
C18547 cal_itt\[2\] FILLER_0_3_221/a_36_472# 0.003825f
C18548 _067_ _039_ 0.221585f
C18549 net80 _434_/a_1000_472# 0.01421f
C18550 ctln[2] ctln[1] 0.047127f
C18551 _024_ _435_/a_448_472# 0.039244f
C18552 _417_/a_796_472# vss 0.001608f
C18553 FILLER_0_9_72/a_124_375# vdd -0.003896f
C18554 result[4] fanout78/a_36_113# 0.001531f
C18555 FILLER_0_20_98/a_124_375# vss 0.013019f
C18556 FILLER_0_20_98/a_36_472# vdd 0.095266f
C18557 _086_ calibrate 0.041755f
C18558 FILLER_0_10_214/a_36_472# _055_ 0.027657f
C18559 output37/a_224_472# sample 0.015298f
C18560 net73 FILLER_0_19_111/a_124_375# 0.005778f
C18561 _081_ net21 0.030964f
C18562 _093_ FILLER_0_18_139/a_124_375# 0.008393f
C18563 output37/a_224_472# net37 0.011407f
C18564 _127_ vss 0.343764f
C18565 FILLER_0_10_78/a_932_472# FILLER_0_9_72/a_1468_375# 0.001543f
C18566 output32/a_224_472# vdd 0.082664f
C18567 _061_ vdd 0.295557f
C18568 net35 FILLER_0_22_86/a_484_472# 0.008347f
C18569 mask\[8\] FILLER_0_22_86/a_932_472# 0.012284f
C18570 _008_ net60 0.314106f
C18571 FILLER_0_5_72/a_1020_375# net47 0.006974f
C18572 _385_/a_36_68# net37 0.047762f
C18573 FILLER_0_21_28/a_124_375# net17 0.005751f
C18574 net65 calibrate 0.012434f
C18575 FILLER_0_13_290/a_124_375# _416_/a_36_151# 0.026277f
C18576 FILLER_0_5_212/a_36_472# _078_ 0.002235f
C18577 FILLER_0_13_212/a_484_472# _043_ 0.011439f
C18578 _453_/a_1308_423# vdd 0.002896f
C18579 _453_/a_448_472# vss 0.00396f
C18580 _311_/a_66_473# vdd 0.106886f
C18581 net35 FILLER_0_22_128/a_3172_472# 0.014415f
C18582 net17 _452_/a_1697_156# 0.001184f
C18583 _015_ _426_/a_448_472# 0.035938f
C18584 net57 _267_/a_1120_472# 0.002885f
C18585 mask\[2\] net30 0.089173f
C18586 FILLER_0_16_89/a_1020_375# _136_ 0.019549f
C18587 _069_ FILLER_0_13_212/a_36_472# 0.047013f
C18588 ctln[1] FILLER_0_3_221/a_572_375# 0.001554f
C18589 ctlp[5] vdd 0.293399f
C18590 net82 _163_ 0.00269f
C18591 FILLER_0_12_2/a_484_472# net67 0.006435f
C18592 _397_/a_36_472# vss 0.003673f
C18593 _037_ vss 0.051886f
C18594 net68 FILLER_0_6_47/a_1828_472# 0.009096f
C18595 output32/a_224_472# net20 0.050019f
C18596 _028_ _154_ 0.174927f
C18597 FILLER_0_11_135/a_36_472# vss 0.006739f
C18598 output46/a_224_472# output44/a_224_472# 0.005749f
C18599 net65 net21 0.04444f
C18600 _001_ vdd 0.122898f
C18601 _131_ _179_ 0.034602f
C18602 net47 _380_/a_224_472# 0.001405f
C18603 ctln[2] FILLER_0_0_266/a_36_472# 0.049163f
C18604 net35 _050_ 0.28822f
C18605 _098_ _437_/a_796_472# 0.0049f
C18606 net63 FILLER_0_15_228/a_36_472# 0.001669f
C18607 net54 FILLER_0_22_128/a_36_472# 0.020739f
C18608 mask\[5\] FILLER_0_18_177/a_124_375# 0.002726f
C18609 _000_ _079_ 0.032884f
C18610 FILLER_0_9_223/a_124_375# _246_/a_36_68# 0.005308f
C18611 FILLER_0_14_91/a_572_375# FILLER_0_14_99/a_36_472# 0.086635f
C18612 FILLER_0_17_72/a_1828_472# _136_ 0.004161f
C18613 FILLER_0_16_89/a_36_472# _451_/a_2449_156# 0.001571f
C18614 vdd _433_/a_36_151# 0.086874f
C18615 mask\[0\] _429_/a_36_151# 0.026729f
C18616 _448_/a_796_472# net59 0.004855f
C18617 output23/a_224_472# net34 0.021474f
C18618 _093_ FILLER_0_18_76/a_572_375# 0.025143f
C18619 _122_ _121_ 0.034975f
C18620 _101_ vdd 0.02756f
C18621 FILLER_0_11_101/a_484_472# vdd 0.009482f
C18622 FILLER_0_11_101/a_36_472# vss 0.001641f
C18623 FILLER_0_14_91/a_124_375# _177_ 0.00134f
C18624 FILLER_0_18_100/a_124_375# mask\[9\] 0.005751f
C18625 _052_ _424_/a_1308_423# 0.008633f
C18626 mask\[1\] FILLER_0_15_180/a_36_472# 0.001145f
C18627 _072_ vdd 0.715894f
C18628 net35 _214_/a_36_160# 0.0116f
C18629 ctln[1] FILLER_0_0_266/a_36_472# 0.011046f
C18630 FILLER_0_4_185/a_36_472# FILLER_0_3_172/a_1380_472# 0.026657f
C18631 output39/a_224_472# net17 0.041253f
C18632 FILLER_0_1_98/a_36_472# _442_/a_2665_112# 0.002597f
C18633 _105_ _048_ 0.02699f
C18634 FILLER_0_4_107/a_572_375# _157_ 0.001032f
C18635 net76 FILLER_0_6_177/a_124_375# 0.00227f
C18636 _085_ _120_ 0.032964f
C18637 _161_ _055_ 0.078364f
C18638 FILLER_0_24_63/a_124_375# output25/a_224_472# 0.007304f
C18639 FILLER_0_19_195/a_124_375# vdd 0.03587f
C18640 net39 _033_ 0.607942f
C18641 _014_ vdd 0.035382f
C18642 _041_ net40 0.082688f
C18643 _053_ _414_/a_2248_156# 0.013478f
C18644 _360_/a_36_160# FILLER_0_4_123/a_124_375# 0.013555f
C18645 vss FILLER_0_13_72/a_36_472# 0.034188f
C18646 _093_ FILLER_0_18_209/a_124_375# 0.00333f
C18647 net68 _440_/a_1000_472# 0.002604f
C18648 _176_ _451_/a_3081_151# 0.001255f
C18649 net31 _421_/a_2665_112# 0.005428f
C18650 net67 FILLER_0_6_47/a_1828_472# 0.001175f
C18651 net15 _304_/a_224_472# 0.001451f
C18652 FILLER_0_16_89/a_36_472# net36 0.010907f
C18653 FILLER_0_20_169/a_36_472# vss 0.005112f
C18654 _074_ FILLER_0_3_172/a_484_472# 0.001763f
C18655 net20 _014_ 0.008597f
C18656 FILLER_0_16_107/a_36_472# FILLER_0_16_89/a_1380_472# 0.003468f
C18657 _413_/a_36_151# FILLER_0_3_172/a_2276_472# 0.001723f
C18658 _000_ cal_itt\[1\] 0.012692f
C18659 _432_/a_2665_112# net21 0.005773f
C18660 _429_/a_36_151# FILLER_0_15_212/a_124_375# 0.059049f
C18661 _415_/a_1308_423# _004_ 0.002098f
C18662 net26 _012_ 0.066032f
C18663 _255_/a_224_552# _161_ 0.025424f
C18664 _181_ _184_ 0.022711f
C18665 _181_ _401_/a_36_68# 0.010647f
C18666 net57 _225_/a_36_160# 0.022745f
C18667 output8/a_224_472# _413_/a_2665_112# 0.010726f
C18668 _053_ net37 0.080949f
C18669 FILLER_0_17_38/a_572_375# _041_ 0.021754f
C18670 FILLER_0_14_50/a_36_472# _174_ 0.015387f
C18671 FILLER_0_2_101/a_124_375# net14 0.0239f
C18672 _031_ vdd 0.327674f
C18673 _090_ net21 0.038093f
C18674 mask\[9\] _438_/a_2665_112# 0.040085f
C18675 net72 _424_/a_36_151# 0.09381f
C18676 _064_ _446_/a_448_472# 0.01156f
C18677 _235_/a_67_603# _446_/a_2665_112# 0.017036f
C18678 ctln[6] net13 0.065837f
C18679 _015_ FILLER_0_8_239/a_124_375# 0.007342f
C18680 _126_ _129_ 0.039006f
C18681 output20/a_224_472# result[9] 0.001884f
C18682 _077_ _062_ 0.037598f
C18683 net52 _442_/a_1000_472# 0.016308f
C18684 _072_ _251_/a_1130_472# 0.004007f
C18685 FILLER_0_18_177/a_1828_472# vdd 0.004845f
C18686 FILLER_0_18_177/a_1380_472# vss -0.001894f
C18687 _165_ FILLER_0_6_47/a_124_375# 0.014312f
C18688 net72 _067_ 0.055817f
C18689 _005_ _416_/a_1308_423# 0.020096f
C18690 FILLER_0_21_142/a_572_375# _140_ 0.018708f
C18691 output8/a_224_472# FILLER_0_3_221/a_932_472# 0.001699f
C18692 FILLER_0_14_81/a_124_375# _177_ 0.002725f
C18693 _441_/a_36_151# _168_ 0.033578f
C18694 fanout53/a_36_160# FILLER_0_16_154/a_932_472# 0.001426f
C18695 net66 FILLER_0_5_54/a_484_472# 0.001863f
C18696 FILLER_0_9_60/a_124_375# vss 0.003217f
C18697 FILLER_0_9_60/a_572_375# vdd 0.031403f
C18698 _140_ FILLER_0_19_155/a_572_375# 0.040109f
C18699 _115_ FILLER_0_11_78/a_484_472# 0.003641f
C18700 net18 _419_/a_2248_156# 0.014287f
C18701 _439_/a_1308_423# FILLER_0_6_47/a_3260_375# 0.001224f
C18702 FILLER_0_18_2/a_2724_472# net40 0.011079f
C18703 ctlp[1] _421_/a_36_151# 0.010453f
C18704 net15 FILLER_0_23_60/a_36_472# 0.004561f
C18705 net61 fanout61/a_36_113# 0.023179f
C18706 net69 _441_/a_2665_112# 0.014995f
C18707 FILLER_0_17_104/a_36_472# net14 0.012286f
C18708 comp net17 0.02802f
C18709 net41 _039_ 0.030362f
C18710 _094_ vdd 0.717159f
C18711 FILLER_0_17_218/a_572_375# vdd 0.019414f
C18712 FILLER_0_17_218/a_124_375# vss 0.012673f
C18713 _100_ vss 0.020176f
C18714 _425_/a_2248_156# vdd 0.010067f
C18715 _069_ _429_/a_796_472# 0.003099f
C18716 mask\[7\] FILLER_0_22_128/a_1828_472# 0.004503f
C18717 FILLER_0_11_101/a_124_375# _171_ 0.00105f
C18718 _297_/a_36_472# vss 0.003601f
C18719 FILLER_0_17_72/a_932_472# _175_ 0.003281f
C18720 _070_ _172_ 0.237178f
C18721 FILLER_0_0_198/a_124_375# net59 0.004565f
C18722 FILLER_0_5_109/a_124_375# _153_ 0.040726f
C18723 _170_ _241_/a_224_472# 0.001199f
C18724 FILLER_0_21_142/a_484_472# net54 0.038728f
C18725 FILLER_0_23_60/a_36_472# FILLER_0_23_44/a_1380_472# 0.013276f
C18726 net53 _427_/a_2665_112# 0.042564f
C18727 FILLER_0_4_197/a_1468_375# net76 0.007667f
C18728 trim_mask\[0\] vss 0.014228f
C18729 _103_ _046_ 0.010317f
C18730 fanout54/a_36_160# _145_ 0.009257f
C18731 net48 _070_ 0.264809f
C18732 _423_/a_36_151# FILLER_0_23_44/a_572_375# 0.059049f
C18733 _448_/a_2665_112# net22 0.010428f
C18734 net20 _094_ 0.677838f
C18735 net70 _043_ 0.045182f
C18736 _098_ FILLER_0_15_212/a_1020_375# 0.00918f
C18737 _428_/a_1204_472# net74 0.009712f
C18738 net50 _439_/a_2248_156# 0.007461f
C18739 FILLER_0_4_144/a_572_375# net23 0.019114f
C18740 _245_/a_672_472# net17 0.00121f
C18741 _367_/a_36_68# _160_ 0.013113f
C18742 FILLER_0_4_144/a_36_472# trim_mask\[4\] 0.017557f
C18743 FILLER_0_4_49/a_484_472# vss 0.002751f
C18744 _086_ FILLER_0_11_142/a_124_375# 0.009046f
C18745 _098_ FILLER_0_16_154/a_932_472# 0.001701f
C18746 FILLER_0_15_142/a_36_472# _136_ 0.003745f
C18747 fanout70/a_36_113# _136_ 0.002788f
C18748 trim[0] net40 0.005988f
C18749 FILLER_0_4_144/a_36_472# net47 0.008498f
C18750 _319_/a_672_472# _125_ 0.002725f
C18751 net54 FILLER_0_19_142/a_124_375# 0.056556f
C18752 _086_ FILLER_0_7_104/a_124_375# 0.001629f
C18753 _098_ FILLER_0_19_111/a_36_472# 0.003915f
C18754 _098_ _434_/a_36_151# 0.019342f
C18755 _412_/a_2248_156# net59 0.008792f
C18756 FILLER_0_19_47/a_572_375# _183_ 0.001186f
C18757 _415_/a_2665_112# fanout62/a_36_160# 0.016426f
C18758 _093_ FILLER_0_17_142/a_36_472# 0.011974f
C18759 _242_/a_36_160# _170_ 0.001933f
C18760 _117_ _310_/a_1133_69# 0.002654f
C18761 FILLER_0_22_86/a_36_472# vss 0.002319f
C18762 _132_ FILLER_0_14_107/a_1380_472# 0.049391f
C18763 _122_ net59 0.041453f
C18764 _189_/a_67_603# FILLER_0_14_235/a_36_472# 0.002778f
C18765 _274_/a_244_497# net64 0.004085f
C18766 net63 FILLER_0_18_177/a_2724_472# 0.001857f
C18767 en_co_clk _171_ 0.003472f
C18768 _140_ FILLER_0_22_128/a_124_375# 0.011452f
C18769 _155_ FILLER_0_4_91/a_572_375# 0.004038f
C18770 output45/a_224_472# vdd -0.026726f
C18771 FILLER_0_22_128/a_2724_472# vss 0.005195f
C18772 FILLER_0_22_128/a_3172_472# vdd 0.003395f
C18773 _108_ _295_/a_36_472# 0.014558f
C18774 _095_ _181_ 0.008117f
C18775 _299_/a_36_472# _109_ 0.030751f
C18776 net35 _435_/a_36_151# 0.038368f
C18777 FILLER_0_7_72/a_124_375# vss 0.044754f
C18778 net27 _426_/a_2560_156# 0.004199f
C18779 _056_ _055_ 0.155993f
C18780 net56 FILLER_0_18_139/a_1380_472# 0.048069f
C18781 net64 net59 0.005832f
C18782 net68 _381_/a_36_472# 0.003421f
C18783 output38/a_224_472# _446_/a_448_472# 0.007649f
C18784 net78 vdd 0.265913f
C18785 _050_ vdd 0.484554f
C18786 _431_/a_36_151# fanout70/a_36_113# 0.016241f
C18787 FILLER_0_15_235/a_572_375# FILLER_0_14_235/a_572_375# 0.05841f
C18788 _442_/a_2248_156# net14 0.025334f
C18789 net63 FILLER_0_17_218/a_484_472# 0.002672f
C18790 _445_/a_1000_472# _034_ 0.007034f
C18791 _445_/a_2665_112# _166_ 0.002292f
C18792 _053_ FILLER_0_6_47/a_932_472# 0.011457f
C18793 net15 _447_/a_36_151# 0.001598f
C18794 FILLER_0_11_142/a_572_375# _121_ 0.003107f
C18795 _030_ net40 0.002509f
C18796 net17 net6 0.063494f
C18797 _185_ _402_/a_718_527# 0.001973f
C18798 net36 FILLER_0_18_76/a_484_472# 0.005765f
C18799 net82 FILLER_0_3_172/a_1380_472# 0.007879f
C18800 FILLER_0_5_54/a_36_472# _164_ 0.003923f
C18801 FILLER_0_8_263/a_36_472# vdd 0.092694f
C18802 FILLER_0_8_263/a_124_375# vss 0.007944f
C18803 result[8] _048_ 0.006006f
C18804 _058_ _059_ 0.990213f
C18805 net34 FILLER_0_22_128/a_1468_375# 0.003214f
C18806 _093_ FILLER_0_18_107/a_1828_472# 0.001872f
C18807 vdd FILLER_0_14_235/a_572_375# 0.006167f
C18808 vss FILLER_0_14_235/a_124_375# 0.002686f
C18809 en_co_clk FILLER_0_13_100/a_36_472# 0.001752f
C18810 FILLER_0_22_86/a_124_375# FILLER_0_23_88/a_36_472# 0.001684f
C18811 net20 net78 1.100401f
C18812 _101_ _283_/a_36_472# 0.002471f
C18813 net34 _207_/a_67_603# 0.008585f
C18814 FILLER_0_3_172/a_484_472# net65 0.003678f
C18815 _322_/a_692_472# net74 0.003192f
C18816 _093_ _102_ 0.008937f
C18817 _098_ FILLER_0_15_205/a_36_472# 0.010528f
C18818 ctln[3] FILLER_0_0_266/a_124_375# 0.002726f
C18819 _446_/a_2665_112# vdd 0.044081f
C18820 mask\[4\] net22 0.075713f
C18821 _210_/a_67_603# vss 0.038142f
C18822 _255_/a_224_552# _056_ 0.033615f
C18823 _412_/a_1308_423# net65 0.024499f
C18824 _214_/a_36_160# vdd 0.010812f
C18825 _069_ _061_ 0.024151f
C18826 _086_ FILLER_0_5_181/a_124_375# 0.006872f
C18827 _161_ state\[1\] 0.002512f
C18828 _443_/a_796_472# vss 0.001654f
C18829 FILLER_0_7_72/a_3260_375# _058_ 0.00258f
C18830 _035_ net49 0.018245f
C18831 _112_ FILLER_0_8_247/a_932_472# 0.001185f
C18832 calibrate FILLER_0_7_233/a_36_472# 0.013262f
C18833 _068_ _055_ 0.443477f
C18834 FILLER_0_21_142/a_572_375# FILLER_0_21_150/a_36_472# 0.086635f
C18835 ctln[2] net18 0.106494f
C18836 _258_/a_36_160# _078_ 0.006096f
C18837 _414_/a_36_151# net21 0.007791f
C18838 net48 _425_/a_448_472# 0.013011f
C18839 _448_/a_2248_156# vss 0.003807f
C18840 _448_/a_2665_112# vdd 0.005876f
C18841 output48/a_224_472# _081_ 0.007705f
C18842 net52 FILLER_0_6_47/a_3172_472# 0.047876f
C18843 _122_ _227_/a_36_160# 0.005128f
C18844 result[7] net61 0.021122f
C18845 _060_ vss 0.318005f
C18846 _126_ FILLER_0_11_135/a_124_375# 0.008245f
C18847 output18/a_224_472# net18 0.01698f
C18848 result[4] _006_ 0.271278f
C18849 _155_ FILLER_0_7_104/a_572_375# 0.002336f
C18850 cal_itt\[3\] net57 0.001586f
C18851 FILLER_0_16_73/a_572_375# _175_ 0.138524f
C18852 _122_ _169_ 0.014463f
C18853 calibrate _163_ 0.026892f
C18854 _017_ _134_ 0.017998f
C18855 _423_/a_36_151# vss 0.012999f
C18856 _423_/a_448_472# vdd 0.01351f
C18857 FILLER_0_16_57/a_572_375# net55 0.004559f
C18858 FILLER_0_16_57/a_36_472# net72 0.040135f
C18859 FILLER_0_14_181/a_124_375# _137_ 0.006021f
C18860 net48 _082_ 0.003853f
C18861 _415_/a_1308_423# net19 0.001498f
C18862 _432_/a_2560_156# _093_ 0.007613f
C18863 FILLER_0_5_54/a_932_472# net47 0.006386f
C18864 FILLER_0_4_197/a_1380_472# net59 0.022002f
C18865 _430_/a_2665_112# fanout63/a_36_160# 0.010365f
C18866 net68 _453_/a_796_472# 0.001516f
C18867 FILLER_0_15_142/a_36_472# net53 0.080484f
C18868 fanout70/a_36_113# net53 0.031633f
C18869 _413_/a_1308_423# _002_ 0.002178f
C18870 cal_count\[3\] _389_/a_36_148# 0.024777f
C18871 net57 _428_/a_1000_472# 0.024803f
C18872 net16 FILLER_0_18_53/a_36_472# 0.001532f
C18873 _092_ FILLER_0_18_209/a_484_472# 0.006303f
C18874 FILLER_0_9_223/a_572_375# state\[0\] 0.079258f
C18875 net55 _183_ 0.024948f
C18876 net21 net11 0.10869f
C18877 output45/a_224_472# output17/a_224_472# 0.071473f
C18878 net32 ctlp[2] 0.097138f
C18879 FILLER_0_17_56/a_36_472# _041_ 0.004881f
C18880 _176_ FILLER_0_18_53/a_36_472# 0.001868f
C18881 net41 net72 0.319547f
C18882 _073_ _080_ 0.455535f
C18883 _118_ _311_/a_3220_473# 0.001133f
C18884 fanout60/a_36_160# FILLER_0_17_282/a_124_375# 0.005489f
C18885 _044_ FILLER_0_14_263/a_36_472# 0.002013f
C18886 _255_/a_224_552# _068_ 0.002412f
C18887 ctln[1] net18 0.004646f
C18888 FILLER_0_24_130/a_124_375# ctlp[7] 0.002726f
C18889 FILLER_0_18_100/a_36_472# FILLER_0_18_107/a_36_472# 0.002764f
C18890 output48/a_224_472# net65 0.015306f
C18891 _126_ _068_ 0.01065f
C18892 fanout62/a_36_160# FILLER_0_9_290/a_36_472# 0.001961f
C18893 FILLER_0_14_81/a_36_472# _451_/a_3129_107# 0.001557f
C18894 fanout55/a_36_160# cal_count\[1\] 0.007256f
C18895 mask\[4\] _433_/a_2665_112# 0.005353f
C18896 FILLER_0_5_206/a_124_375# net59 0.008027f
C18897 FILLER_0_17_72/a_36_472# vss 0.036865f
C18898 _134_ FILLER_0_10_107/a_36_472# 0.006746f
C18899 _072_ _069_ 0.265737f
C18900 _181_ _402_/a_1296_93# 0.040412f
C18901 net22 _435_/a_36_151# 0.001559f
C18902 ctln[1] _411_/a_448_472# 0.039538f
C18903 net16 FILLER_0_10_28/a_124_375# 0.002225f
C18904 _132_ FILLER_0_18_107/a_2364_375# 0.006403f
C18905 _075_ FILLER_0_5_206/a_36_472# 0.001503f
C18906 trimb[1] net43 0.004299f
C18907 vss FILLER_0_6_37/a_36_472# 0.006755f
C18908 _427_/a_796_472# vss 0.001131f
C18909 trim_mask\[4\] _370_/a_1152_472# 0.001449f
C18910 net17 _450_/a_2225_156# 0.033342f
C18911 net52 FILLER_0_2_111/a_1380_472# 0.050754f
C18912 trim_mask\[1\] vdd 0.241393f
C18913 output11/a_224_472# vdd 0.01016f
C18914 output16/a_224_472# vdd 0.006151f
C18915 _436_/a_36_151# FILLER_0_22_107/a_124_375# 0.026916f
C18916 _081_ _242_/a_36_160# 0.025059f
C18917 _033_ net47 0.056436f
C18918 net76 FILLER_0_3_172/a_124_375# 0.001186f
C18919 _444_/a_448_472# net42 0.002526f
C18920 _116_ vss 0.235141f
C18921 FILLER_0_12_220/a_36_472# _070_ 0.087648f
C18922 FILLER_0_7_146/a_124_375# _372_/a_170_472# 0.001188f
C18923 _091_ FILLER_0_15_212/a_484_472# 0.049391f
C18924 net52 _440_/a_2665_112# 0.005084f
C18925 mask\[4\] FILLER_0_20_177/a_484_472# 0.001215f
C18926 _321_/a_3662_472# vdd 0.001229f
C18927 _144_ FILLER_0_22_128/a_3260_375# 0.006444f
C18928 FILLER_0_8_24/a_124_375# net42 0.032303f
C18929 fanout74/a_36_113# trim_mask\[4\] 0.026261f
C18930 _144_ net33 0.042826f
C18931 _104_ fanout63/a_36_160# 0.007014f
C18932 trim[4] _236_/a_36_160# 0.004514f
C18933 _095_ FILLER_0_13_72/a_36_472# 0.00819f
C18934 output11/a_224_472# net20 0.036556f
C18935 FILLER_0_4_144/a_36_472# FILLER_0_3_142/a_124_375# 0.001543f
C18936 FILLER_0_6_79/a_36_472# _164_ 0.008685f
C18937 _452_/a_1040_527# _041_ 0.002066f
C18938 _094_ _283_/a_36_472# 0.004373f
C18939 mask\[4\] vdd 0.794539f
C18940 _046_ mask\[2\] 0.003147f
C18941 _114_ _096_ 0.066848f
C18942 net49 _440_/a_2665_112# 0.025303f
C18943 net39 _444_/a_36_151# 0.14155f
C18944 _157_ vdd 0.419501f
C18945 _020_ FILLER_0_18_107/a_2276_472# 0.004069f
C18946 _350_/a_665_69# mask\[6\] 0.001069f
C18947 _142_ vdd 0.090938f
C18948 _447_/a_2248_156# vss 0.003961f
C18949 _447_/a_2665_112# vdd 0.022038f
C18950 FILLER_0_18_107/a_1468_375# net71 0.001292f
C18951 FILLER_0_4_144/a_572_375# net57 0.001254f
C18952 _373_/a_1060_68# _090_ 0.002234f
C18953 FILLER_0_16_57/a_484_472# cal_count\[1\] 0.001664f
C18954 _118_ vss 0.217218f
C18955 _117_ net21 0.016722f
C18956 mask\[9\] vdd 0.940144f
C18957 net23 FILLER_0_22_128/a_3260_375# 0.012171f
C18958 _137_ FILLER_0_16_154/a_1380_472# 0.005667f
C18959 mask\[3\] _137_ 0.231419f
C18960 net54 _433_/a_2560_156# 0.014333f
C18961 FILLER_0_18_107/a_572_375# mask\[9\] 0.005368f
C18962 FILLER_0_17_64/a_36_472# FILLER_0_17_56/a_572_375# 0.086635f
C18963 sample fanout64/a_36_160# 0.007266f
C18964 net61 net79 0.159f
C18965 _431_/a_36_151# FILLER_0_18_107/a_1828_472# 0.001221f
C18966 _077_ net14 0.03359f
C18967 FILLER_0_2_111/a_572_375# _160_ 0.001049f
C18968 _365_/a_36_68# _156_ 0.027744f
C18969 _432_/a_2560_156# _136_ 0.001178f
C18970 net73 _131_ 0.022043f
C18971 FILLER_0_17_218/a_572_375# _069_ 0.001464f
C18972 FILLER_0_7_59/a_484_472# _439_/a_36_151# 0.001061f
C18973 _444_/a_2248_156# _054_ 0.002637f
C18974 net75 _426_/a_36_151# 0.070626f
C18975 _440_/a_448_472# _160_ 0.004748f
C18976 _127_ _332_/a_36_472# 0.00288f
C18977 _056_ state\[1\] 0.219625f
C18978 _109_ vss 0.023215f
C18979 net71 _437_/a_36_151# 0.055761f
C18980 FILLER_0_18_2/a_2724_472# _452_/a_1040_527# 0.001138f
C18981 FILLER_0_18_2/a_932_472# _452_/a_2225_156# 0.001256f
C18982 _328_/a_36_113# net14 0.002272f
C18983 _435_/a_36_151# vdd 0.059103f
C18984 net27 net18 0.092379f
C18985 _449_/a_36_151# FILLER_0_13_72/a_484_472# 0.001723f
C18986 output9/a_224_472# cal_itt\[0\] 0.008307f
C18987 fanout74/a_36_113# net74 0.007425f
C18988 _187_ _039_ 0.228074f
C18989 _139_ _098_ 0.026578f
C18990 _103_ _418_/a_1308_423# 0.004778f
C18991 _414_/a_2665_112# _068_ 0.002324f
C18992 _103_ _006_ 0.00205f
C18993 _070_ net37 0.036662f
C18994 _126_ _138_ 0.003253f
C18995 output24/a_224_472# net54 0.177947f
C18996 FILLER_0_15_116/a_36_472# FILLER_0_16_115/a_124_375# 0.001597f
C18997 _443_/a_36_151# _032_ 0.0737f
C18998 _422_/a_1000_472# _109_ 0.003473f
C18999 _110_ mask\[8\] 0.05045f
C19000 _413_/a_36_151# _079_ 0.0017f
C19001 _123_ vss 0.016878f
C19002 net81 _018_ 0.081888f
C19003 FILLER_0_7_146/a_36_472# net37 0.00208f
C19004 net54 vss 0.715177f
C19005 trim_mask\[2\] FILLER_0_4_91/a_36_472# 0.003327f
C19006 _444_/a_2248_156# vss 0.001329f
C19007 _444_/a_2665_112# vdd 0.029351f
C19008 result[9] _421_/a_448_472# 0.015264f
C19009 output20/a_224_472# net78 0.001495f
C19010 _073_ vss 0.216342f
C19011 _115_ net23 0.018953f
C19012 _204_/a_67_603# _201_/a_67_603# 0.001129f
C19013 net7 net16 0.033509f
C19014 trim_val\[4\] _443_/a_36_151# 0.009986f
C19015 net25 FILLER_0_23_60/a_124_375# 0.004431f
C19016 net69 _367_/a_244_472# 0.001708f
C19017 _442_/a_2248_156# _153_ 0.0011f
C19018 net74 FILLER_0_2_127/a_124_375# 0.001389f
C19019 _079_ _078_ 0.03338f
C19020 net78 _419_/a_796_472# 0.00376f
C19021 _120_ net14 0.024442f
C19022 _160_ _034_ 0.00905f
C19023 net29 _417_/a_2665_112# 0.002977f
C19024 _147_ _023_ 0.004036f
C19025 net65 FILLER_0_1_212/a_36_472# 0.004414f
C19026 _328_/a_36_113# _428_/a_36_151# 0.030244f
C19027 _438_/a_2248_156# net14 0.045909f
C19028 _339_/a_36_160# FILLER_0_19_171/a_124_375# 0.006021f
C19029 _337_/a_257_69# vdd 0.002972f
C19030 FILLER_0_7_162/a_36_472# calibrate 0.014431f
C19031 net31 _094_ 0.203395f
C19032 _034_ 0 0.304805f
C19033 _160_ 0 1.542665f
C19034 _166_ 0 0.299751f
C19035 trim[3] 0 1.777626f
C19036 output41/a_224_472# 0 2.38465f
C19037 clkc 0 0.763769f
C19038 net6 0 1.112469f
C19039 output6/a_224_472# 0 2.38465f
C19040 FILLER_0_12_196/a_36_472# 0 0.417394f
C19041 FILLER_0_12_196/a_124_375# 0 0.246306f
C19042 result[3] 0 0.50376f
C19043 net30 0 1.81422f
C19044 output30/a_224_472# 0 2.38465f
C19045 _047_ 0 0.374694f
C19046 _201_/a_67_603# 0 0.345683f
C19047 _416_/a_2560_156# 0 0.016968f
C19048 _416_/a_2665_112# 0 0.62251f
C19049 _416_/a_2248_156# 0 0.371662f
C19050 _416_/a_1204_472# 0 0.012971f
C19051 _416_/a_1000_472# 0 0.291735f
C19052 _416_/a_796_472# 0 0.023206f
C19053 _416_/a_1308_423# 0 0.279043f
C19054 _416_/a_448_472# 0 0.684413f
C19055 _416_/a_36_151# 0 1.43589f
C19056 FILLER_0_13_290/a_36_472# 0 0.417394f
C19057 FILLER_0_13_290/a_124_375# 0 0.246306f
C19058 _278_/a_36_160# 0 0.696445f
C19059 _145_ 0 0.546455f
C19060 FILLER_0_13_72/a_484_472# 0 0.345058f
C19061 FILLER_0_13_72/a_36_472# 0 0.404746f
C19062 FILLER_0_13_72/a_572_375# 0 0.232991f
C19063 FILLER_0_13_72/a_124_375# 0 0.185089f
C19064 FILLER_0_14_235/a_484_472# 0 0.345058f
C19065 FILLER_0_14_235/a_36_472# 0 0.404746f
C19066 FILLER_0_14_235/a_572_375# 0 0.232991f
C19067 FILLER_0_14_235/a_124_375# 0 0.185089f
C19068 _156_ 0 0.593796f
C19069 _107_ 0 0.391583f
C19070 _295_/a_36_472# 0 0.031137f
C19071 _022_ 0 0.387773f
C19072 _433_/a_2560_156# 0 0.016968f
C19073 _433_/a_2665_112# 0 0.62251f
C19074 _433_/a_2248_156# 0 0.371662f
C19075 _433_/a_1204_472# 0 0.012971f
C19076 _433_/a_1000_472# 0 0.291735f
C19077 _433_/a_796_472# 0 0.023206f
C19078 _433_/a_1308_423# 0 0.279043f
C19079 _433_/a_448_472# 0 0.684413f
C19080 _433_/a_36_151# 0 1.43589f
C19081 FILLER_0_5_148/a_484_472# 0 0.345058f
C19082 FILLER_0_5_148/a_36_472# 0 0.404746f
C19083 FILLER_0_5_148/a_572_375# 0 0.232991f
C19084 FILLER_0_5_148/a_124_375# 0 0.185089f
C19085 _167_ 0 0.285904f
C19086 _381_/a_36_472# 0 0.031137f
C19087 trim[2] 0 0.79181f
C19088 net40 0 1.845219f
C19089 output40/a_224_472# 0 2.38465f
C19090 cal_count\[0\] 0 0.893784f
C19091 _039_ 0 0.412301f
C19092 _450_/a_2449_156# 0 0.049992f
C19093 _450_/a_2225_156# 0 0.434082f
C19094 _450_/a_3129_107# 0 0.58406f
C19095 _450_/a_836_156# 0 0.019766f
C19096 _450_/a_1040_527# 0 0.302082f
C19097 _450_/a_1353_112# 0 0.286513f
C19098 _450_/a_448_472# 0 1.21246f
C19099 _450_/a_36_151# 0 1.31409f
C19100 rstn 0 1.86494f
C19101 FILLER_0_8_156/a_484_472# 0 0.345058f
C19102 FILLER_0_8_156/a_36_472# 0 0.404746f
C19103 FILLER_0_8_156/a_572_375# 0 0.232991f
C19104 FILLER_0_8_156/a_124_375# 0 0.185089f
C19105 FILLER_0_6_37/a_36_472# 0 0.417394f
C19106 FILLER_0_6_37/a_124_375# 0 0.246306f
C19107 FILLER_0_21_60/a_484_472# 0 0.345058f
C19108 FILLER_0_21_60/a_36_472# 0 0.404746f
C19109 FILLER_0_21_60/a_572_375# 0 0.232991f
C19110 FILLER_0_21_60/a_124_375# 0 0.185089f
C19111 FILLER_0_22_107/a_484_472# 0 0.345058f
C19112 FILLER_0_22_107/a_36_472# 0 0.404746f
C19113 FILLER_0_22_107/a_572_375# 0 0.232991f
C19114 FILLER_0_22_107/a_124_375# 0 0.185089f
C19115 FILLER_0_16_115/a_36_472# 0 0.417394f
C19116 FILLER_0_16_115/a_124_375# 0 0.246306f
C19117 FILLER_0_19_134/a_36_472# 0 0.417394f
C19118 FILLER_0_19_134/a_124_375# 0 0.246306f
C19119 FILLER_0_3_212/a_36_472# 0 0.417394f
C19120 FILLER_0_3_212/a_124_375# 0 0.246306f
C19121 FILLER_0_10_94/a_484_472# 0 0.345058f
C19122 FILLER_0_10_94/a_36_472# 0 0.404746f
C19123 FILLER_0_10_94/a_572_375# 0 0.232991f
C19124 FILLER_0_10_94/a_124_375# 0 0.185089f
C19125 FILLER_0_4_91/a_484_472# 0 0.345058f
C19126 FILLER_0_4_91/a_36_472# 0 0.404746f
C19127 FILLER_0_4_91/a_572_375# 0 0.232991f
C19128 FILLER_0_4_91/a_124_375# 0 0.185089f
C19129 net14 0 1.508711f
C19130 _202_/a_36_160# 0 0.696445f
C19131 FILLER_0_6_231/a_484_472# 0 0.345058f
C19132 FILLER_0_6_231/a_36_472# 0 0.404746f
C19133 FILLER_0_6_231/a_572_375# 0 0.232991f
C19134 FILLER_0_6_231/a_124_375# 0 0.185089f
C19135 vss 0 65.60368f
C19136 vdd 0 1.086009p
C19137 _006_ 0 0.41456f
C19138 _417_/a_2560_156# 0 0.016968f
C19139 _417_/a_2665_112# 0 0.62251f
C19140 _417_/a_2248_156# 0 0.371662f
C19141 _417_/a_1204_472# 0 0.012971f
C19142 _417_/a_1000_472# 0 0.291735f
C19143 _417_/a_796_472# 0 0.023206f
C19144 _417_/a_1308_423# 0 0.279043f
C19145 _417_/a_448_472# 0 0.684413f
C19146 _417_/a_36_151# 0 1.43589f
C19147 _146_ 0 0.35443f
C19148 mask\[6\] 0 1.246962f
C19149 _348_/a_49_472# 0 0.054843f
C19150 _365_/a_36_68# 0 0.150048f
C19151 _023_ 0 0.345812f
C19152 _434_/a_2560_156# 0 0.016968f
C19153 _434_/a_2665_112# 0 0.62251f
C19154 _434_/a_2248_156# 0 0.371662f
C19155 _434_/a_1204_472# 0 0.012971f
C19156 _434_/a_1000_472# 0 0.291735f
C19157 _434_/a_796_472# 0 0.023206f
C19158 _434_/a_1308_423# 0 0.279043f
C19159 _434_/a_448_472# 0 0.684413f
C19160 _434_/a_36_151# 0 1.43589f
C19161 FILLER_0_5_136/a_36_472# 0 0.417394f
C19162 FILLER_0_5_136/a_124_375# 0 0.246306f
C19163 FILLER_0_18_209/a_484_472# 0 0.345058f
C19164 FILLER_0_18_209/a_36_472# 0 0.404746f
C19165 FILLER_0_18_209/a_572_375# 0 0.232991f
C19166 FILLER_0_18_209/a_124_375# 0 0.185089f
C19167 FILLER_0_12_28/a_36_472# 0 0.417394f
C19168 FILLER_0_12_28/a_124_375# 0 0.246306f
C19169 _040_ 0 0.355703f
C19170 _451_/a_2449_156# 0 0.049992f
C19171 _451_/a_2225_156# 0 0.434082f
C19172 _451_/a_3129_107# 0 0.58406f
C19173 _451_/a_836_156# 0 0.019766f
C19174 _451_/a_1040_527# 0 0.302082f
C19175 _451_/a_1353_112# 0 0.286513f
C19176 _451_/a_448_472# 0 1.21246f
C19177 _451_/a_36_151# 0 1.31409f
C19178 FILLER_0_6_47/a_3172_472# 0 0.345058f
C19179 FILLER_0_6_47/a_2724_472# 0 0.33241f
C19180 FILLER_0_6_47/a_2276_472# 0 0.33241f
C19181 FILLER_0_6_47/a_1828_472# 0 0.33241f
C19182 FILLER_0_6_47/a_1380_472# 0 0.33241f
C19183 FILLER_0_6_47/a_932_472# 0 0.33241f
C19184 FILLER_0_6_47/a_484_472# 0 0.33241f
C19185 FILLER_0_6_47/a_36_472# 0 0.404746f
C19186 FILLER_0_6_47/a_3260_375# 0 0.233093f
C19187 FILLER_0_6_47/a_2812_375# 0 0.17167f
C19188 FILLER_0_6_47/a_2364_375# 0 0.17167f
C19189 FILLER_0_6_47/a_1916_375# 0 0.17167f
C19190 FILLER_0_6_47/a_1468_375# 0 0.17167f
C19191 FILLER_0_6_47/a_1020_375# 0 0.17167f
C19192 FILLER_0_6_47/a_572_375# 0 0.17167f
C19193 FILLER_0_6_47/a_124_375# 0 0.185915f
C19194 FILLER_0_21_150/a_36_472# 0 0.417394f
C19195 FILLER_0_21_150/a_124_375# 0 0.246306f
C19196 FILLER_0_15_180/a_484_472# 0 0.345058f
C19197 FILLER_0_15_180/a_36_472# 0 0.404746f
C19198 FILLER_0_15_180/a_572_375# 0 0.232991f
C19199 FILLER_0_15_180/a_124_375# 0 0.185089f
C19200 FILLER_0_22_128/a_3172_472# 0 0.345058f
C19201 FILLER_0_22_128/a_2724_472# 0 0.33241f
C19202 FILLER_0_22_128/a_2276_472# 0 0.33241f
C19203 FILLER_0_22_128/a_1828_472# 0 0.33241f
C19204 FILLER_0_22_128/a_1380_472# 0 0.33241f
C19205 FILLER_0_22_128/a_932_472# 0 0.33241f
C19206 FILLER_0_22_128/a_484_472# 0 0.33241f
C19207 FILLER_0_22_128/a_36_472# 0 0.404746f
C19208 FILLER_0_22_128/a_3260_375# 0 0.233093f
C19209 FILLER_0_22_128/a_2812_375# 0 0.17167f
C19210 FILLER_0_22_128/a_2364_375# 0 0.17167f
C19211 FILLER_0_22_128/a_1916_375# 0 0.17167f
C19212 FILLER_0_22_128/a_1468_375# 0 0.17167f
C19213 FILLER_0_22_128/a_1020_375# 0 0.17167f
C19214 FILLER_0_22_128/a_572_375# 0 0.17167f
C19215 FILLER_0_22_128/a_124_375# 0 0.185915f
C19216 FILLER_0_19_111/a_484_472# 0 0.345058f
C19217 FILLER_0_19_111/a_36_472# 0 0.404746f
C19218 FILLER_0_19_111/a_572_375# 0 0.232991f
C19219 FILLER_0_19_111/a_124_375# 0 0.185089f
C19220 FILLER_0_19_155/a_484_472# 0 0.345058f
C19221 FILLER_0_19_155/a_36_472# 0 0.404746f
C19222 FILLER_0_19_155/a_572_375# 0 0.232991f
C19223 FILLER_0_19_155/a_124_375# 0 0.185089f
C19224 net11 0 1.328455f
C19225 net21 0 1.922829f
C19226 _007_ 0 0.309495f
C19227 net77 0 1.39077f
C19228 _418_/a_2560_156# 0 0.016968f
C19229 _418_/a_2665_112# 0 0.62251f
C19230 _418_/a_2248_156# 0 0.371662f
C19231 _418_/a_1204_472# 0 0.012971f
C19232 _418_/a_1000_472# 0 0.291735f
C19233 _418_/a_796_472# 0 0.023206f
C19234 _418_/a_1308_423# 0 0.279043f
C19235 _418_/a_448_472# 0 0.684413f
C19236 _418_/a_36_151# 0 1.43589f
C19237 _220_/a_67_603# 0 0.345683f
C19238 FILLER_0_9_282/a_484_472# 0 0.345058f
C19239 FILLER_0_9_282/a_36_472# 0 0.404746f
C19240 FILLER_0_9_282/a_572_375# 0 0.232991f
C19241 FILLER_0_9_282/a_124_375# 0 0.185089f
C19242 FILLER_0_18_37/a_1380_472# 0 0.345058f
C19243 FILLER_0_18_37/a_932_472# 0 0.33241f
C19244 FILLER_0_18_37/a_484_472# 0 0.33241f
C19245 FILLER_0_18_37/a_36_472# 0 0.404746f
C19246 FILLER_0_18_37/a_1468_375# 0 0.233029f
C19247 FILLER_0_18_37/a_1020_375# 0 0.171606f
C19248 FILLER_0_18_37/a_572_375# 0 0.171606f
C19249 FILLER_0_18_37/a_124_375# 0 0.185399f
C19250 FILLER_0_2_127/a_36_472# 0 0.417394f
C19251 FILLER_0_2_127/a_124_375# 0 0.246306f
C19252 _157_ 0 0.531763f
C19253 _435_/a_2560_156# 0 0.016968f
C19254 _435_/a_2665_112# 0 0.62251f
C19255 _435_/a_2248_156# 0 0.371662f
C19256 _435_/a_1204_472# 0 0.012971f
C19257 _435_/a_1000_472# 0 0.291735f
C19258 _435_/a_796_472# 0 0.023206f
C19259 _435_/a_1308_423# 0 0.279043f
C19260 _435_/a_448_472# 0 0.684413f
C19261 _435_/a_36_151# 0 1.43589f
C19262 _108_ 0 0.411979f
C19263 _297_/a_36_472# 0 0.031137f
C19264 trim_mask\[3\] 0 1.081535f
C19265 _164_ 0 1.3268f
C19266 _383_/a_36_472# 0 0.031137f
C19267 _041_ 0 0.299289f
C19268 _452_/a_2449_156# 0 0.049992f
C19269 _452_/a_2225_156# 0 0.434082f
C19270 _452_/a_3129_107# 0 0.58406f
C19271 _452_/a_836_156# 0 0.019766f
C19272 _452_/a_1040_527# 0 0.302082f
C19273 _452_/a_1353_112# 0 0.286513f
C19274 _452_/a_448_472# 0 1.21246f
C19275 _452_/a_36_151# 0 1.31409f
C19276 FILLER_0_6_79/a_36_472# 0 0.417394f
C19277 FILLER_0_6_79/a_124_375# 0 0.246306f
C19278 net59 0 5.044369f
C19279 FILLER_0_15_59/a_484_472# 0 0.345058f
C19280 FILLER_0_15_59/a_36_472# 0 0.404746f
C19281 FILLER_0_15_59/a_572_375# 0 0.232991f
C19282 FILLER_0_15_59/a_124_375# 0 0.185089f
C19283 FILLER_0_3_221/a_1380_472# 0 0.345058f
C19284 FILLER_0_3_221/a_932_472# 0 0.33241f
C19285 FILLER_0_3_221/a_484_472# 0 0.33241f
C19286 FILLER_0_3_221/a_36_472# 0 0.404746f
C19287 FILLER_0_3_221/a_1468_375# 0 0.233029f
C19288 FILLER_0_3_221/a_1020_375# 0 0.171606f
C19289 FILLER_0_3_221/a_572_375# 0 0.171606f
C19290 FILLER_0_3_221/a_124_375# 0 0.185399f
C19291 FILLER_0_19_187/a_484_472# 0 0.345058f
C19292 FILLER_0_19_187/a_36_472# 0 0.404746f
C19293 FILLER_0_19_187/a_572_375# 0 0.232991f
C19294 FILLER_0_19_187/a_124_375# 0 0.185089f
C19295 FILLER_0_20_15/a_1380_472# 0 0.345058f
C19296 FILLER_0_20_15/a_932_472# 0 0.33241f
C19297 FILLER_0_20_15/a_484_472# 0 0.33241f
C19298 FILLER_0_20_15/a_36_472# 0 0.404746f
C19299 FILLER_0_20_15/a_1468_375# 0 0.233029f
C19300 FILLER_0_20_15/a_1020_375# 0 0.171606f
C19301 FILLER_0_20_15/a_572_375# 0 0.171606f
C19302 FILLER_0_20_15/a_124_375# 0 0.185399f
C19303 _204_/a_67_603# 0 0.345683f
C19304 _419_/a_2560_156# 0 0.016968f
C19305 _419_/a_2665_112# 0 0.62251f
C19306 _419_/a_2248_156# 0 0.371662f
C19307 _419_/a_1204_472# 0 0.012971f
C19308 _419_/a_1000_472# 0 0.291735f
C19309 _419_/a_796_472# 0 0.023206f
C19310 _419_/a_1308_423# 0 0.279043f
C19311 _419_/a_448_472# 0 0.684413f
C19312 _419_/a_36_151# 0 1.43589f
C19313 _054_ 0 0.522819f
C19314 _221_/a_36_160# 0 0.386641f
C19315 FILLER_0_9_270/a_484_472# 0 0.345058f
C19316 FILLER_0_9_270/a_36_472# 0 0.404746f
C19317 FILLER_0_9_270/a_572_375# 0 0.232991f
C19318 FILLER_0_9_270/a_124_375# 0 0.185089f
C19319 FILLER_0_1_192/a_36_472# 0 0.417394f
C19320 FILLER_0_1_192/a_124_375# 0 0.246306f
C19321 FILLER_0_13_80/a_36_472# 0 0.417394f
C19322 FILLER_0_13_80/a_124_375# 0 0.246306f
C19323 _153_ 0 1.165862f
C19324 _154_ 0 1.167112f
C19325 _367_/a_36_68# 0 0.150048f
C19326 _436_/a_2560_156# 0 0.016968f
C19327 _436_/a_2665_112# 0 0.62251f
C19328 _436_/a_2248_156# 0 0.371662f
C19329 _436_/a_1204_472# 0 0.012971f
C19330 _436_/a_1000_472# 0 0.291735f
C19331 _436_/a_796_472# 0 0.023206f
C19332 _436_/a_1308_423# 0 0.279043f
C19333 _436_/a_448_472# 0 0.684413f
C19334 _436_/a_36_151# 0 1.43589f
C19335 FILLER_0_10_107/a_484_472# 0 0.345058f
C19336 FILLER_0_10_107/a_36_472# 0 0.404746f
C19337 FILLER_0_10_107/a_572_375# 0 0.232991f
C19338 FILLER_0_10_107/a_124_375# 0 0.185089f
C19339 _168_ 0 0.336537f
C19340 net51 0 2.105066f
C19341 _042_ 0 0.323587f
C19342 _453_/a_2560_156# 0 0.016968f
C19343 _453_/a_2665_112# 0 0.62251f
C19344 _453_/a_2248_156# 0 0.371662f
C19345 _453_/a_1204_472# 0 0.012971f
C19346 _453_/a_1000_472# 0 0.291735f
C19347 _453_/a_796_472# 0 0.023206f
C19348 _453_/a_1308_423# 0 0.279043f
C19349 _453_/a_448_472# 0 0.684413f
C19350 _453_/a_36_151# 0 1.43589f
C19351 FILLER_0_19_142/a_36_472# 0 0.417394f
C19352 FILLER_0_19_142/a_124_375# 0 0.246306f
C19353 _048_ 0 0.358805f
C19354 _205_/a_36_160# 0 0.696445f
C19355 net43 0 1.236377f
C19356 FILLER_0_3_78/a_484_472# 0 0.345058f
C19357 FILLER_0_3_78/a_36_472# 0 0.404746f
C19358 FILLER_0_3_78/a_572_375# 0 0.232991f
C19359 FILLER_0_3_78/a_124_375# 0 0.185089f
C19360 _437_/a_2560_156# 0 0.016968f
C19361 _437_/a_2665_112# 0 0.62251f
C19362 _437_/a_2248_156# 0 0.371662f
C19363 _437_/a_1204_472# 0 0.012971f
C19364 _437_/a_1000_472# 0 0.291735f
C19365 _437_/a_796_472# 0 0.023206f
C19366 _437_/a_1308_423# 0 0.279043f
C19367 _437_/a_448_472# 0 0.684413f
C19368 _437_/a_36_151# 0 1.43589f
C19369 _109_ 0 0.319326f
C19370 _299_/a_36_472# 0 0.031137f
C19371 net37 0 1.529713f
C19372 _385_/a_36_68# 0 0.112263f
C19373 FILLER_0_0_266/a_36_472# 0 0.417394f
C19374 FILLER_0_0_266/a_124_375# 0 0.246306f
C19375 net12 0 1.263595f
C19376 net22 0 2.108509f
C19377 FILLER_0_9_290/a_36_472# 0 0.417394f
C19378 FILLER_0_9_290/a_124_375# 0 0.246306f
C19379 _223_/a_36_160# 0 0.696445f
C19380 FILLER_0_14_263/a_36_472# 0 0.417394f
C19381 FILLER_0_14_263/a_124_375# 0 0.246306f
C19382 _158_ 0 0.309522f
C19383 _369_/a_36_68# 0 0.150048f
C19384 net71 0 1.420869f
C19385 _438_/a_2560_156# 0 0.016968f
C19386 _438_/a_2665_112# 0 0.62251f
C19387 _438_/a_2248_156# 0 0.371662f
C19388 _438_/a_1204_472# 0 0.012971f
C19389 _438_/a_1000_472# 0 0.291735f
C19390 _438_/a_796_472# 0 0.023206f
C19391 _438_/a_1308_423# 0 0.279043f
C19392 _438_/a_448_472# 0 0.684413f
C19393 _438_/a_36_151# 0 1.43589f
C19394 FILLER_0_23_274/a_36_472# 0 0.417394f
C19395 FILLER_0_23_274/a_124_375# 0 0.246306f
C19396 FILLER_0_17_282/a_36_472# 0 0.417394f
C19397 FILLER_0_17_282/a_124_375# 0 0.246306f
C19398 FILLER_0_5_198/a_484_472# 0 0.345058f
C19399 FILLER_0_5_198/a_36_472# 0 0.404746f
C19400 FILLER_0_5_198/a_572_375# 0 0.232991f
C19401 FILLER_0_5_198/a_124_375# 0 0.185089f
C19402 _163_ 0 1.03762f
C19403 _169_ 0 0.245383f
C19404 _386_/a_848_380# 0 0.40208f
C19405 _386_/a_124_24# 0 0.591898f
C19406 FILLER_0_20_2/a_484_472# 0 0.345058f
C19407 FILLER_0_20_2/a_36_472# 0 0.404746f
C19408 FILLER_0_20_2/a_572_375# 0 0.232991f
C19409 FILLER_0_20_2/a_124_375# 0 0.185089f
C19410 FILLER_0_16_154/a_1380_472# 0 0.345058f
C19411 FILLER_0_16_154/a_932_472# 0 0.33241f
C19412 FILLER_0_16_154/a_484_472# 0 0.33241f
C19413 FILLER_0_16_154/a_36_472# 0 0.404746f
C19414 FILLER_0_16_154/a_1468_375# 0 0.233029f
C19415 FILLER_0_16_154/a_1020_375# 0 0.171606f
C19416 FILLER_0_16_154/a_572_375# 0 0.171606f
C19417 FILLER_0_16_154/a_124_375# 0 0.185399f
C19418 FILLER_0_0_232/a_36_472# 0 0.417394f
C19419 FILLER_0_0_232/a_124_375# 0 0.246306f
C19420 FILLER_0_19_195/a_36_472# 0 0.417394f
C19421 FILLER_0_19_195/a_124_375# 0 0.246306f
C19422 _049_ 0 0.329957f
C19423 net33 0 1.934915f
C19424 _207_/a_67_603# 0 0.345683f
C19425 FILLER_0_3_54/a_36_472# 0 0.417394f
C19426 FILLER_0_3_54/a_124_375# 0 0.246306f
C19427 FILLER_0_2_101/a_36_472# 0 0.417394f
C19428 FILLER_0_2_101/a_124_375# 0 0.246306f
C19429 trim_mask\[0\] 0 0.605753f
C19430 _439_/a_2560_156# 0 0.016968f
C19431 _439_/a_2665_112# 0 0.62251f
C19432 _439_/a_2248_156# 0 0.371662f
C19433 _439_/a_1204_472# 0 0.012971f
C19434 _439_/a_1000_472# 0 0.291735f
C19435 _439_/a_796_472# 0 0.023206f
C19436 _439_/a_1308_423# 0 0.279043f
C19437 _439_/a_448_472# 0 0.684413f
C19438 _439_/a_36_151# 0 1.43589f
C19439 _066_ 0 0.333041f
C19440 FILLER_0_23_44/a_1380_472# 0 0.345058f
C19441 FILLER_0_23_44/a_932_472# 0 0.33241f
C19442 FILLER_0_23_44/a_484_472# 0 0.33241f
C19443 FILLER_0_23_44/a_36_472# 0 0.404746f
C19444 FILLER_0_23_44/a_1468_375# 0 0.233029f
C19445 FILLER_0_23_44/a_1020_375# 0 0.171606f
C19446 FILLER_0_23_44/a_572_375# 0 0.171606f
C19447 FILLER_0_23_44/a_124_375# 0 0.185399f
C19448 FILLER_0_23_88/a_36_472# 0 0.417394f
C19449 FILLER_0_23_88/a_124_375# 0 0.246306f
C19450 FILLER_0_5_164/a_484_472# 0 0.345058f
C19451 FILLER_0_5_164/a_36_472# 0 0.404746f
C19452 FILLER_0_5_164/a_572_375# 0 0.232991f
C19453 FILLER_0_5_164/a_124_375# 0 0.185089f
C19454 _060_ 0 2.485177f
C19455 _113_ 0 2.833205f
C19456 _090_ 0 2.629271f
C19457 _310_/a_49_472# 0 0.098072f
C19458 _037_ 0 0.467089f
C19459 _170_ 0 0.413995f
C19460 _387_/a_36_113# 0 0.418095f
C19461 _208_/a_36_160# 0 0.696445f
C19462 FILLER_0_18_76/a_484_472# 0 0.345058f
C19463 FILLER_0_18_76/a_36_472# 0 0.404746f
C19464 FILLER_0_18_76/a_572_375# 0 0.232991f
C19465 FILLER_0_18_76/a_124_375# 0 0.185089f
C19466 _225_/a_36_160# 0 0.386641f
C19467 FILLER_0_2_177/a_484_472# 0 0.345058f
C19468 FILLER_0_2_177/a_36_472# 0 0.404746f
C19469 FILLER_0_2_177/a_572_375# 0 0.232991f
C19470 FILLER_0_2_177/a_124_375# 0 0.185089f
C19471 FILLER_0_2_111/a_1380_472# 0 0.345058f
C19472 FILLER_0_2_111/a_932_472# 0 0.33241f
C19473 FILLER_0_2_111/a_484_472# 0 0.33241f
C19474 FILLER_0_2_111/a_36_472# 0 0.404746f
C19475 FILLER_0_2_111/a_1468_375# 0 0.233029f
C19476 FILLER_0_2_111/a_1020_375# 0 0.171606f
C19477 FILLER_0_2_111/a_572_375# 0 0.171606f
C19478 FILLER_0_2_111/a_124_375# 0 0.185399f
C19479 FILLER_0_15_228/a_36_472# 0 0.417394f
C19480 FILLER_0_15_228/a_124_375# 0 0.246306f
C19481 net47 0 2.314376f
C19482 _242_/a_36_160# 0 0.696445f
C19483 _117_ 0 1.266251f
C19484 _311_/a_66_473# 0 0.11665f
C19485 _043_ 0 0.487279f
C19486 _190_/a_36_160# 0 0.696445f
C19487 FILLER_0_9_105/a_484_472# 0 0.345058f
C19488 FILLER_0_9_105/a_36_472# 0 0.404746f
C19489 FILLER_0_9_105/a_572_375# 0 0.232991f
C19490 FILLER_0_9_105/a_124_375# 0 0.185089f
C19491 FILLER_0_13_100/a_36_472# 0 0.417394f
C19492 FILLER_0_13_100/a_124_375# 0 0.246306f
C19493 FILLER_0_22_177/a_1380_472# 0 0.345058f
C19494 FILLER_0_22_177/a_932_472# 0 0.33241f
C19495 FILLER_0_22_177/a_484_472# 0 0.33241f
C19496 FILLER_0_22_177/a_36_472# 0 0.404746f
C19497 FILLER_0_22_177/a_1468_375# 0 0.233029f
C19498 FILLER_0_22_177/a_1020_375# 0 0.171606f
C19499 FILLER_0_22_177/a_572_375# 0 0.171606f
C19500 FILLER_0_22_177/a_124_375# 0 0.185399f
C19501 FILLER_0_15_2/a_484_472# 0 0.345058f
C19502 FILLER_0_15_2/a_36_472# 0 0.404746f
C19503 FILLER_0_15_2/a_572_375# 0 0.232991f
C19504 FILLER_0_15_2/a_124_375# 0 0.185089f
C19505 FILLER_0_15_10/a_36_472# 0 0.417394f
C19506 FILLER_0_15_10/a_124_375# 0 0.246306f
C19507 FILLER_0_19_171/a_1380_472# 0 0.345058f
C19508 FILLER_0_19_171/a_932_472# 0 0.33241f
C19509 FILLER_0_19_171/a_484_472# 0 0.33241f
C19510 FILLER_0_19_171/a_36_472# 0 0.404746f
C19511 FILLER_0_19_171/a_1468_375# 0 0.233029f
C19512 FILLER_0_19_171/a_1020_375# 0 0.171606f
C19513 FILLER_0_19_171/a_572_375# 0 0.171606f
C19514 FILLER_0_19_171/a_124_375# 0 0.185399f
C19515 net13 0 1.176306f
C19516 net23 0 2.091399f
C19517 FILLER_0_20_87/a_36_472# 0 0.417394f
C19518 FILLER_0_20_87/a_124_375# 0 0.246306f
C19519 FILLER_0_20_98/a_36_472# 0 0.417394f
C19520 FILLER_0_20_98/a_124_375# 0 0.246306f
C19521 _055_ 0 1.782885f
C19522 FILLER_0_18_53/a_484_472# 0 0.345058f
C19523 FILLER_0_18_53/a_36_472# 0 0.404746f
C19524 FILLER_0_18_53/a_572_375# 0 0.232991f
C19525 FILLER_0_18_53/a_124_375# 0 0.185089f
C19526 FILLER_0_2_165/a_36_472# 0 0.417394f
C19527 FILLER_0_2_165/a_124_375# 0 0.246306f
C19528 FILLER_0_15_205/a_36_472# 0 0.417394f
C19529 FILLER_0_15_205/a_124_375# 0 0.246306f
C19530 FILLER_0_23_282/a_484_472# 0 0.345058f
C19531 FILLER_0_23_282/a_36_472# 0 0.404746f
C19532 FILLER_0_23_282/a_572_375# 0 0.232991f
C19533 FILLER_0_23_282/a_124_375# 0 0.185089f
C19534 net42 0 1.067446f
C19535 net17 0 2.210219f
C19536 _172_ 0 0.265782f
C19537 _171_ 0 0.300355f
C19538 _389_/a_36_148# 0 0.388358f
C19539 _080_ 0 0.328202f
C19540 _260_/a_36_68# 0 0.112263f
C19541 FILLER_0_0_96/a_36_472# 0 0.417394f
C19542 FILLER_0_0_96/a_124_375# 0 0.246306f
C19543 FILLER_0_9_72/a_1380_472# 0 0.345058f
C19544 FILLER_0_9_72/a_932_472# 0 0.33241f
C19545 FILLER_0_9_72/a_484_472# 0 0.33241f
C19546 FILLER_0_9_72/a_36_472# 0 0.404746f
C19547 FILLER_0_9_72/a_1468_375# 0 0.233029f
C19548 FILLER_0_9_72/a_1020_375# 0 0.171606f
C19549 FILLER_0_9_72/a_572_375# 0 0.171606f
C19550 FILLER_0_9_72/a_124_375# 0 0.185399f
C19551 FILLER_0_20_31/a_36_472# 0 0.417394f
C19552 FILLER_0_20_31/a_124_375# 0 0.246306f
C19553 _227_/a_36_160# 0 0.386641f
C19554 _120_ 0 1.533088f
C19555 _313_/a_67_603# 0 0.345683f
C19556 FILLER_0_5_172/a_36_472# 0 0.417394f
C19557 FILLER_0_5_172/a_124_375# 0 0.246306f
C19558 FILLER_0_12_20/a_484_472# 0 0.345058f
C19559 FILLER_0_12_20/a_36_472# 0 0.404746f
C19560 FILLER_0_12_20/a_572_375# 0 0.232991f
C19561 FILLER_0_12_20/a_124_375# 0 0.185089f
C19562 _134_ 0 0.365972f
C19563 _062_ 0 1.717773f
C19564 _059_ 0 1.686761f
C19565 _261_/a_36_160# 0 0.386641f
C19566 _044_ 0 0.388801f
C19567 mask\[1\] 0 1.295078f
C19568 _192_/a_67_603# 0 0.345683f
C19569 FILLER_0_13_142/a_1380_472# 0 0.345058f
C19570 FILLER_0_13_142/a_932_472# 0 0.33241f
C19571 FILLER_0_13_142/a_484_472# 0 0.33241f
C19572 FILLER_0_13_142/a_36_472# 0 0.404746f
C19573 FILLER_0_13_142/a_1468_375# 0 0.233029f
C19574 FILLER_0_13_142/a_1020_375# 0 0.171606f
C19575 FILLER_0_13_142/a_572_375# 0 0.171606f
C19576 FILLER_0_13_142/a_124_375# 0 0.185399f
C19577 FILLER_0_9_60/a_484_472# 0 0.345058f
C19578 FILLER_0_9_60/a_36_472# 0 0.404746f
C19579 FILLER_0_9_60/a_572_375# 0 0.232991f
C19580 FILLER_0_9_60/a_124_375# 0 0.185089f
C19581 FILLER_0_7_233/a_36_472# 0 0.417394f
C19582 FILLER_0_7_233/a_124_375# 0 0.246306f
C19583 _228_/a_36_68# 0 0.69549f
C19584 FILLER_0_21_206/a_36_472# 0 0.417394f
C19585 FILLER_0_21_206/a_124_375# 0 0.246306f
C19586 _067_ 0 0.851951f
C19587 _135_ 0 0.339478f
C19588 _193_/a_36_160# 0 0.696445f
C19589 _180_ 0 0.390598f
C19590 cal_count\[1\] 0 1.568289f
C19591 FILLER_0_4_213/a_484_472# 0 0.345058f
C19592 FILLER_0_4_213/a_36_472# 0 0.404746f
C19593 FILLER_0_4_213/a_572_375# 0 0.232991f
C19594 FILLER_0_4_213/a_124_375# 0 0.185089f
C19595 FILLER_0_11_282/a_36_472# 0 0.417394f
C19596 FILLER_0_11_282/a_124_375# 0 0.246306f
C19597 FILLER_0_18_61/a_36_472# 0 0.417394f
C19598 FILLER_0_18_61/a_124_375# 0 0.246306f
C19599 FILLER_0_15_235/a_484_472# 0 0.345058f
C19600 FILLER_0_15_235/a_36_472# 0 0.404746f
C19601 FILLER_0_15_235/a_572_375# 0 0.232991f
C19602 FILLER_0_15_235/a_124_375# 0 0.185089f
C19603 FILLER_0_23_290/a_36_472# 0 0.417394f
C19604 FILLER_0_23_290/a_124_375# 0 0.246306f
C19605 _121_ 0 0.532847f
C19606 _315_/a_36_68# 0 0.052951f
C19607 _246_/a_36_68# 0 0.69549f
C19608 FILLER_0_5_181/a_36_472# 0 0.417394f
C19609 FILLER_0_5_181/a_124_375# 0 0.246306f
C19610 _082_ 0 0.619901f
C19611 net8 0 1.163723f
C19612 net18 0 2.032159f
C19613 _332_/a_36_472# 0 0.031137f
C19614 _179_ 0 0.336984f
C19615 _401_/a_36_68# 0 0.112263f
C19616 FILLER_0_14_107/a_1380_472# 0 0.345058f
C19617 FILLER_0_14_107/a_932_472# 0 0.33241f
C19618 FILLER_0_14_107/a_484_472# 0 0.33241f
C19619 FILLER_0_14_107/a_36_472# 0 0.404746f
C19620 FILLER_0_14_107/a_1468_375# 0 0.233029f
C19621 FILLER_0_14_107/a_1020_375# 0 0.171606f
C19622 FILLER_0_14_107/a_572_375# 0 0.171606f
C19623 FILLER_0_14_107/a_124_375# 0 0.185399f
C19624 _097_ 0 0.592554f
C19625 FILLER_0_1_204/a_36_472# 0 0.417394f
C19626 FILLER_0_1_204/a_124_375# 0 0.246306f
C19627 FILLER_0_15_72/a_484_472# 0 0.345058f
C19628 FILLER_0_15_72/a_36_472# 0 0.404746f
C19629 FILLER_0_15_72/a_572_375# 0 0.232991f
C19630 FILLER_0_15_72/a_124_375# 0 0.185089f
C19631 FILLER_0_17_104/a_1380_472# 0 0.345058f
C19632 FILLER_0_17_104/a_932_472# 0 0.33241f
C19633 FILLER_0_17_104/a_484_472# 0 0.33241f
C19634 FILLER_0_17_104/a_36_472# 0 0.404746f
C19635 FILLER_0_17_104/a_1468_375# 0 0.233029f
C19636 FILLER_0_17_104/a_1020_375# 0 0.171606f
C19637 FILLER_0_17_104/a_572_375# 0 0.171606f
C19638 FILLER_0_17_104/a_124_375# 0 0.185399f
C19639 FILLER_0_8_37/a_484_472# 0 0.345058f
C19640 FILLER_0_8_37/a_36_472# 0 0.404746f
C19641 FILLER_0_8_37/a_572_375# 0 0.232991f
C19642 FILLER_0_8_37/a_124_375# 0 0.185089f
C19643 FILLER_0_15_212/a_1380_472# 0 0.345058f
C19644 FILLER_0_15_212/a_932_472# 0 0.33241f
C19645 FILLER_0_15_212/a_484_472# 0 0.33241f
C19646 FILLER_0_15_212/a_36_472# 0 0.404746f
C19647 FILLER_0_15_212/a_1468_375# 0 0.233029f
C19648 FILLER_0_15_212/a_1020_375# 0 0.171606f
C19649 FILLER_0_15_212/a_572_375# 0 0.171606f
C19650 FILLER_0_15_212/a_124_375# 0 0.185399f
C19651 FILLER_0_23_60/a_36_472# 0 0.417394f
C19652 FILLER_0_23_60/a_124_375# 0 0.246306f
C19653 _123_ 0 0.344874f
C19654 _122_ 0 0.600118f
C19655 calibrate 0 1.343796f
C19656 _316_/a_848_380# 0 0.40208f
C19657 _316_/a_124_24# 0 0.591898f
C19658 _247_/a_36_160# 0 0.696445f
C19659 FILLER_0_12_50/a_36_472# 0 0.417394f
C19660 FILLER_0_12_50/a_124_375# 0 0.246306f
C19661 _084_ 0 0.296163f
C19662 cal_itt\[0\] 0 1.831055f
C19663 cal_itt\[1\] 0 1.705665f
C19664 FILLER_0_11_109/a_36_472# 0 0.417394f
C19665 FILLER_0_11_109/a_124_375# 0 0.246306f
C19666 _182_ 0 0.34197f
C19667 _402_/a_1948_68# 0 0.022025f
C19668 _402_/a_718_527# 0 0.001795f
C19669 _402_/a_56_567# 0 0.424713f
C19670 _402_/a_728_93# 0 0.65929f
C19671 _402_/a_1296_93# 0 0.317801f
C19672 _045_ 0 0.349338f
C19673 mask\[2\] 0 1.335688f
C19674 _195_/a_67_603# 0 0.345683f
C19675 _333_/a_36_160# 0 0.386641f
C19676 _098_ 0 1.816151f
C19677 _147_ 0 0.322539f
C19678 _350_/a_49_472# 0 0.054843f
C19679 FILLER_0_12_236/a_484_472# 0 0.345058f
C19680 FILLER_0_12_236/a_36_472# 0 0.404746f
C19681 FILLER_0_12_236/a_572_375# 0 0.232991f
C19682 FILLER_0_12_236/a_124_375# 0 0.185089f
C19683 FILLER_0_2_171/a_36_472# 0 0.417394f
C19684 FILLER_0_2_171/a_124_375# 0 0.246306f
C19685 _014_ 0 0.363432f
C19686 _317_/a_36_113# 0 0.418095f
C19687 _248_/a_36_68# 0 0.69549f
C19688 FILLER_0_17_38/a_484_472# 0 0.345058f
C19689 FILLER_0_17_38/a_36_472# 0 0.404746f
C19690 FILLER_0_17_38/a_572_375# 0 0.232991f
C19691 FILLER_0_17_38/a_124_375# 0 0.185089f
C19692 _001_ 0 0.285216f
C19693 _265_/a_244_68# 0 0.138666f
C19694 _196_/a_36_160# 0 0.696445f
C19695 FILLER_0_6_90/a_484_472# 0 0.345058f
C19696 FILLER_0_6_90/a_36_472# 0 0.404746f
C19697 FILLER_0_6_90/a_572_375# 0 0.232991f
C19698 FILLER_0_6_90/a_124_375# 0 0.185089f
C19699 _183_ 0 0.356629f
C19700 _334_/a_36_160# 0 0.386641f
C19701 _282_/a_36_160# 0 0.386641f
C19702 _024_ 0 0.451815f
C19703 _009_ 0 0.397943f
C19704 _420_/a_2560_156# 0 0.016968f
C19705 _420_/a_2665_112# 0 0.62251f
C19706 _420_/a_2248_156# 0 0.371662f
C19707 _420_/a_1204_472# 0 0.012971f
C19708 _420_/a_1000_472# 0 0.291735f
C19709 _420_/a_796_472# 0 0.023206f
C19710 _420_/a_1308_423# 0 0.279043f
C19711 _420_/a_448_472# 0 0.684413f
C19712 _420_/a_36_151# 0 1.43589f
C19713 clk 0 1.162312f
C19714 FILLER_0_8_2/a_36_472# 0 0.417394f
C19715 FILLER_0_8_2/a_124_375# 0 0.246306f
C19716 FILLER_0_8_24/a_484_472# 0 0.345058f
C19717 FILLER_0_8_24/a_36_472# 0 0.404746f
C19718 FILLER_0_8_24/a_572_375# 0 0.232991f
C19719 FILLER_0_8_24/a_124_375# 0 0.185089f
C19720 _124_ 0 0.294081f
C19721 _118_ 0 1.378735f
C19722 _071_ 0 1.600488f
C19723 net9 0 1.13171f
C19724 net19 0 1.889339f
C19725 _138_ 0 0.33132f
C19726 _137_ 0 1.178616f
C19727 _335_/a_49_472# 0 0.054843f
C19728 _404_/a_36_472# 0 0.031137f
C19729 FILLER_0_20_107/a_36_472# 0 0.417394f
C19730 FILLER_0_20_107/a_124_375# 0 0.246306f
C19731 FILLER_0_9_142/a_36_472# 0 0.417394f
C19732 FILLER_0_9_142/a_124_375# 0 0.246306f
C19733 _099_ 0 1.152785f
C19734 _283_/a_36_472# 0 0.031137f
C19735 mask\[7\] 0 1.477838f
C19736 _352_/a_49_472# 0 0.054843f
C19737 _010_ 0 0.377779f
C19738 _421_/a_2560_156# 0 0.016968f
C19739 _421_/a_2665_112# 0 0.62251f
C19740 _421_/a_2248_156# 0 0.371662f
C19741 _421_/a_1204_472# 0 0.012971f
C19742 _421_/a_1000_472# 0 0.291735f
C19743 _421_/a_796_472# 0 0.023206f
C19744 _421_/a_1308_423# 0 0.279043f
C19745 _421_/a_448_472# 0 0.684413f
C19746 _421_/a_36_151# 0 1.43589f
C19747 FILLER_0_1_212/a_36_472# 0 0.417394f
C19748 FILLER_0_1_212/a_124_375# 0 0.246306f
C19749 FILLER_0_8_239/a_36_472# 0 0.417394f
C19750 FILLER_0_8_239/a_124_375# 0 0.246306f
C19751 _125_ 0 1.526603f
C19752 _058_ 0 1.483584f
C19753 FILLER_0_6_177/a_484_472# 0 0.345058f
C19754 FILLER_0_6_177/a_36_472# 0 0.404746f
C19755 FILLER_0_6_177/a_572_375# 0 0.232991f
C19756 FILLER_0_6_177/a_124_375# 0 0.185089f
C19757 state\[1\] 0 2.652405f
C19758 _267_/a_36_472# 0 0.137725f
C19759 _184_ 0 0.350066f
C19760 cal_count\[2\] 0 1.971854f
C19761 _405_/a_67_603# 0 0.345683f
C19762 _018_ 0 0.358633f
C19763 _046_ 0 0.361963f
C19764 _198_/a_67_603# 0 0.345683f
C19765 _094_ 0 1.263877f
C19766 _100_ 0 0.333135f
C19767 net36 0 2.262756f
C19768 FILLER_0_17_133/a_36_472# 0 0.417394f
C19769 FILLER_0_17_133/a_124_375# 0 0.246306f
C19770 _025_ 0 0.350324f
C19771 _148_ 0 0.325709f
C19772 _422_/a_2560_156# 0 0.016968f
C19773 _422_/a_2665_112# 0 0.62251f
C19774 _422_/a_2248_156# 0 0.371662f
C19775 _422_/a_1204_472# 0 0.012971f
C19776 _422_/a_1000_472# 0 0.291735f
C19777 _422_/a_796_472# 0 0.023206f
C19778 _422_/a_1308_423# 0 0.279043f
C19779 _422_/a_448_472# 0 0.684413f
C19780 _422_/a_36_151# 0 1.43589f
C19781 FILLER_0_1_266/a_484_472# 0 0.345058f
C19782 FILLER_0_1_266/a_36_472# 0 0.404746f
C19783 FILLER_0_1_266/a_572_375# 0 0.232991f
C19784 FILLER_0_1_266/a_124_375# 0 0.185089f
C19785 _152_ 0 0.918583f
C19786 _081_ 0 1.140656f
C19787 _370_/a_848_380# 0 0.40208f
C19788 _370_/a_124_24# 0 0.591898f
C19789 FILLER_0_24_274/a_1380_472# 0 0.345058f
C19790 FILLER_0_24_274/a_932_472# 0 0.33241f
C19791 FILLER_0_24_274/a_484_472# 0 0.33241f
C19792 FILLER_0_24_274/a_36_472# 0 0.404746f
C19793 FILLER_0_24_274/a_1468_375# 0 0.233029f
C19794 FILLER_0_24_274/a_1020_375# 0 0.171606f
C19795 FILLER_0_24_274/a_572_375# 0 0.171606f
C19796 FILLER_0_24_274/a_124_375# 0 0.185399f
C19797 _185_ 0 0.386917f
C19798 _406_/a_36_159# 0 0.374116f
C19799 _337_/a_49_472# 0 0.054843f
C19800 _199_/a_36_160# 0 0.696445f
C19801 _285_/a_36_472# 0 0.031137f
C19802 _354_/a_49_472# 0 0.054843f
C19803 _012_ 0 0.75195f
C19804 _423_/a_2560_156# 0 0.016968f
C19805 _423_/a_2665_112# 0 0.62251f
C19806 _423_/a_2248_156# 0 0.371662f
C19807 _423_/a_1204_472# 0 0.012971f
C19808 _423_/a_1000_472# 0 0.291735f
C19809 _423_/a_796_472# 0 0.023206f
C19810 _423_/a_1308_423# 0 0.279043f
C19811 _423_/a_448_472# 0 0.684413f
C19812 _423_/a_36_151# 0 1.43589f
C19813 FILLER_0_5_88/a_36_472# 0 0.417394f
C19814 FILLER_0_5_88/a_124_375# 0 0.246306f
C19815 trim_mask\[1\] 0 1.020743f
C19816 _029_ 0 0.308904f
C19817 _440_/a_2560_156# 0 0.016968f
C19818 _440_/a_2665_112# 0 0.62251f
C19819 _440_/a_2248_156# 0 0.371662f
C19820 _440_/a_1204_472# 0 0.012971f
C19821 _440_/a_1000_472# 0 0.291735f
C19822 _440_/a_796_472# 0 0.023206f
C19823 _440_/a_1308_423# 0 0.279043f
C19824 _440_/a_448_472# 0 0.684413f
C19825 _440_/a_36_151# 0 1.43589f
C19826 _159_ 0 0.351814f
C19827 _371_/a_36_113# 0 0.418095f
C19828 FILLER_0_17_56/a_484_472# 0 0.345058f
C19829 FILLER_0_17_56/a_36_472# 0 0.404746f
C19830 FILLER_0_17_56/a_572_375# 0 0.232991f
C19831 FILLER_0_17_56/a_124_375# 0 0.185089f
C19832 _083_ 0 0.527882f
C19833 _078_ 0 0.904554f
C19834 _269_/a_36_472# 0 0.031137f
C19835 _181_ 0 0.829168f
C19836 _407_/a_36_472# 0 0.031137f
C19837 _019_ 0 0.32907f
C19838 _139_ 0 0.346404f
C19839 FILLER_0_14_123/a_36_472# 0 0.417394f
C19840 FILLER_0_14_123/a_124_375# 0 0.246306f
C19841 _005_ 0 0.340993f
C19842 _101_ 0 0.280497f
C19843 _424_/a_2560_156# 0 0.016968f
C19844 _424_/a_2665_112# 0 0.62251f
C19845 _424_/a_2248_156# 0 0.371662f
C19846 _424_/a_1204_472# 0 0.012971f
C19847 _424_/a_1000_472# 0 0.291735f
C19848 _424_/a_796_472# 0 0.023206f
C19849 _424_/a_1308_423# 0 0.279043f
C19850 _424_/a_448_472# 0 0.684413f
C19851 _424_/a_36_151# 0 1.43589f
C19852 _026_ 0 0.320379f
C19853 _149_ 0 0.305496f
C19854 FILLER_0_5_54/a_1380_472# 0 0.345058f
C19855 FILLER_0_5_54/a_932_472# 0 0.33241f
C19856 FILLER_0_5_54/a_484_472# 0 0.33241f
C19857 FILLER_0_5_54/a_36_472# 0 0.404746f
C19858 FILLER_0_5_54/a_1468_375# 0 0.233029f
C19859 FILLER_0_5_54/a_1020_375# 0 0.171606f
C19860 FILLER_0_5_54/a_572_375# 0 0.171606f
C19861 FILLER_0_5_54/a_124_375# 0 0.185399f
C19862 FILLER_0_17_142/a_484_472# 0 0.345058f
C19863 FILLER_0_17_142/a_36_472# 0 0.404746f
C19864 FILLER_0_17_142/a_572_375# 0 0.232991f
C19865 FILLER_0_17_142/a_124_375# 0 0.185089f
C19866 _068_ 0 3.162692f
C19867 _076_ 0 3.812442f
C19868 _133_ 0 1.430901f
C19869 _070_ 0 3.115722f
C19870 _372_/a_170_472# 0 0.077257f
C19871 net49 0 5.140563f
C19872 _030_ 0 0.307083f
C19873 net66 0 1.472669f
C19874 _441_/a_2560_156# 0 0.016968f
C19875 _441_/a_2665_112# 0 0.62251f
C19876 _441_/a_2248_156# 0 0.371662f
C19877 _441_/a_1204_472# 0 0.012971f
C19878 _441_/a_1000_472# 0 0.291735f
C19879 _441_/a_796_472# 0 0.023206f
C19880 _441_/a_1308_423# 0 0.279043f
C19881 _441_/a_448_472# 0 0.684413f
C19882 _441_/a_36_151# 0 1.43589f
C19883 FILLER_0_5_206/a_36_472# 0 0.417394f
C19884 FILLER_0_5_206/a_124_375# 0 0.246306f
C19885 fanout49/a_36_160# 0 0.696445f
C19886 FILLER_0_8_247/a_1380_472# 0 0.345058f
C19887 FILLER_0_8_247/a_932_472# 0 0.33241f
C19888 FILLER_0_8_247/a_484_472# 0 0.33241f
C19889 FILLER_0_8_247/a_36_472# 0 0.404746f
C19890 FILLER_0_8_247/a_1468_375# 0 0.233029f
C19891 FILLER_0_8_247/a_1020_375# 0 0.171606f
C19892 FILLER_0_8_247/a_572_375# 0 0.171606f
C19893 FILLER_0_8_247/a_124_375# 0 0.185399f
C19894 FILLER_0_12_220/a_1380_472# 0 0.345058f
C19895 FILLER_0_12_220/a_932_472# 0 0.33241f
C19896 FILLER_0_12_220/a_484_472# 0 0.33241f
C19897 FILLER_0_12_220/a_36_472# 0 0.404746f
C19898 FILLER_0_12_220/a_1468_375# 0 0.233029f
C19899 FILLER_0_12_220/a_1020_375# 0 0.171606f
C19900 FILLER_0_12_220/a_572_375# 0 0.171606f
C19901 FILLER_0_12_220/a_124_375# 0 0.185399f
C19902 FILLER_0_21_286/a_484_472# 0 0.345058f
C19903 FILLER_0_21_286/a_36_472# 0 0.404746f
C19904 FILLER_0_21_286/a_572_375# 0 0.232991f
C19905 FILLER_0_21_286/a_124_375# 0 0.185089f
C19906 _140_ 0 1.276518f
C19907 _339_/a_36_160# 0 0.386641f
C19908 _095_ 0 2.689027f
C19909 _186_ 0 0.580923f
C19910 _408_/a_1936_472# 0 0.009918f
C19911 _408_/a_718_524# 0 0.005143f
C19912 _408_/a_56_524# 0 0.41096f
C19913 _408_/a_728_93# 0 0.654825f
C19914 _408_/a_1336_472# 0 0.316639f
C19915 FILLER_0_20_169/a_36_472# 0 0.417394f
C19916 FILLER_0_20_169/a_124_375# 0 0.246306f
C19917 _210_/a_67_603# 0 0.345683f
C19918 _425_/a_2560_156# 0 0.016968f
C19919 _425_/a_2665_112# 0 0.62251f
C19920 _425_/a_2248_156# 0 0.371662f
C19921 _425_/a_1204_472# 0 0.012971f
C19922 _425_/a_1000_472# 0 0.291735f
C19923 _425_/a_796_472# 0 0.023206f
C19924 _425_/a_1308_423# 0 0.279043f
C19925 _425_/a_448_472# 0 0.684413f
C19926 _425_/a_36_151# 0 1.43589f
C19927 net5 0 0.610761f
C19928 input5/a_36_113# 0 0.418095f
C19929 FILLER_0_11_78/a_484_472# 0 0.345058f
C19930 FILLER_0_11_78/a_36_472# 0 0.404746f
C19931 FILLER_0_11_78/a_572_375# 0 0.232991f
C19932 FILLER_0_11_78/a_124_375# 0 0.185089f
C19933 _102_ 0 0.335308f
C19934 _287_/a_36_472# 0 0.031137f
C19935 mask\[9\] 0 1.383606f
C19936 _356_/a_36_472# 0 0.031137f
C19937 _031_ 0 0.417351f
C19938 net69 0 1.020293f
C19939 _442_/a_2560_156# 0 0.016968f
C19940 _442_/a_2665_112# 0 0.62251f
C19941 _442_/a_2248_156# 0 0.371662f
C19942 _442_/a_1204_472# 0 0.012971f
C19943 _442_/a_1000_472# 0 0.291735f
C19944 _442_/a_796_472# 0 0.023206f
C19945 _442_/a_1308_423# 0 0.279043f
C19946 _442_/a_448_472# 0 0.684413f
C19947 _442_/a_36_151# 0 1.43589f
C19948 net64 0 2.598514f
C19949 fanout59/a_36_160# 0 0.696445f
C19950 FILLER_0_14_99/a_36_472# 0 0.417394f
C19951 FILLER_0_14_99/a_124_375# 0 0.246306f
C19952 _038_ 0 0.362839f
C19953 _136_ 0 1.345638f
C19954 _390_/a_36_68# 0 0.150048f
C19955 FILLER_0_15_282/a_484_472# 0 0.345058f
C19956 FILLER_0_15_282/a_36_472# 0 0.404746f
C19957 FILLER_0_15_282/a_572_375# 0 0.232991f
C19958 FILLER_0_15_282/a_124_375# 0 0.185089f
C19959 FILLER_0_11_124/a_36_472# 0 0.417394f
C19960 FILLER_0_11_124/a_124_375# 0 0.246306f
C19961 FILLER_0_11_135/a_36_472# 0 0.417394f
C19962 FILLER_0_11_135/a_124_375# 0 0.246306f
C19963 _188_ 0 0.349407f
C19964 cal_count\[3\] 0 1.862896f
C19965 _050_ 0 0.622354f
C19966 _211_/a_36_160# 0 0.386641f
C19967 net4 0 2.711508f
C19968 en 0 0.833743f
C19969 input4/a_36_68# 0 0.69549f
C19970 _426_/a_2560_156# 0 0.016968f
C19971 _426_/a_2665_112# 0 0.62251f
C19972 _426_/a_2248_156# 0 0.371662f
C19973 _426_/a_1204_472# 0 0.012971f
C19974 _426_/a_1000_472# 0 0.291735f
C19975 _426_/a_796_472# 0 0.023206f
C19976 _426_/a_1308_423# 0 0.279043f
C19977 _426_/a_448_472# 0 0.684413f
C19978 _426_/a_36_151# 0 1.43589f
C19979 _027_ 0 0.302949f
C19980 _150_ 0 0.320497f
C19981 FILLER_0_18_107/a_3172_472# 0 0.345058f
C19982 FILLER_0_18_107/a_2724_472# 0 0.33241f
C19983 FILLER_0_18_107/a_2276_472# 0 0.33241f
C19984 FILLER_0_18_107/a_1828_472# 0 0.33241f
C19985 FILLER_0_18_107/a_1380_472# 0 0.33241f
C19986 FILLER_0_18_107/a_932_472# 0 0.33241f
C19987 FILLER_0_18_107/a_484_472# 0 0.33241f
C19988 FILLER_0_18_107/a_36_472# 0 0.404746f
C19989 FILLER_0_18_107/a_3260_375# 0 0.233093f
C19990 FILLER_0_18_107/a_2812_375# 0 0.17167f
C19991 FILLER_0_18_107/a_2364_375# 0 0.17167f
C19992 FILLER_0_18_107/a_1916_375# 0 0.17167f
C19993 FILLER_0_18_107/a_1468_375# 0 0.17167f
C19994 FILLER_0_18_107/a_1020_375# 0 0.17167f
C19995 FILLER_0_18_107/a_572_375# 0 0.17167f
C19996 FILLER_0_18_107/a_124_375# 0 0.185915f
C19997 trim_mask\[4\] 0 0.987791f
C19998 _032_ 0 0.34876f
C19999 _443_/a_2560_156# 0 0.016968f
C20000 _443_/a_2665_112# 0 0.62251f
C20001 _443_/a_2248_156# 0 0.371662f
C20002 _443_/a_1204_472# 0 0.012971f
C20003 _443_/a_1000_472# 0 0.291735f
C20004 _443_/a_796_472# 0 0.023206f
C20005 _443_/a_1308_423# 0 0.279043f
C20006 _443_/a_448_472# 0 0.684413f
C20007 _443_/a_36_151# 0 1.43589f
C20008 _061_ 0 0.84986f
C20009 _056_ 0 2.393362f
C20010 _374_/a_36_68# 0 0.112263f
C20011 fanout58/a_36_160# 0 0.696445f
C20012 net74 0 1.237373f
C20013 fanout69/a_36_113# 0 0.418095f
C20014 _173_ 0 0.339446f
C20015 FILLER_0_3_142/a_36_472# 0 0.417394f
C20016 FILLER_0_3_142/a_124_375# 0 0.246306f
C20017 FILLER_0_17_64/a_36_472# 0 0.417394f
C20018 FILLER_0_17_64/a_124_375# 0 0.246306f
C20019 FILLER_0_11_101/a_484_472# 0 0.345058f
C20020 FILLER_0_11_101/a_36_472# 0 0.404746f
C20021 FILLER_0_11_101/a_572_375# 0 0.232991f
C20022 FILLER_0_11_101/a_124_375# 0 0.185089f
C20023 FILLER_0_22_86/a_1380_472# 0 0.345058f
C20024 FILLER_0_22_86/a_932_472# 0 0.33241f
C20025 FILLER_0_22_86/a_484_472# 0 0.33241f
C20026 FILLER_0_22_86/a_36_472# 0 0.404746f
C20027 FILLER_0_22_86/a_1468_375# 0 0.233029f
C20028 FILLER_0_22_86/a_1020_375# 0 0.171606f
C20029 FILLER_0_22_86/a_572_375# 0 0.171606f
C20030 FILLER_0_22_86/a_124_375# 0 0.185399f
C20031 net24 0 1.61895f
C20032 net3 0 0.740676f
C20033 input3/a_36_113# 0 0.418095f
C20034 _103_ 0 0.350464f
C20035 _289_/a_36_472# 0 0.031137f
C20036 _151_ 0 0.300777f
C20037 _427_/a_2560_156# 0 0.016968f
C20038 _427_/a_2665_112# 0 0.91969f
C20039 _427_/a_2248_156# 0 0.30886f
C20040 _427_/a_1204_472# 0 0.012971f
C20041 _427_/a_1000_472# 0 0.291735f
C20042 _427_/a_796_472# 0 0.023206f
C20043 _427_/a_1308_423# 0 0.279043f
C20044 _427_/a_448_472# 0 0.684413f
C20045 _427_/a_36_151# 0 1.43587f
C20046 FILLER_0_17_161/a_36_472# 0 0.417394f
C20047 FILLER_0_17_161/a_124_375# 0 0.246306f
C20048 FILLER_0_18_139/a_1380_472# 0 0.345058f
C20049 FILLER_0_18_139/a_932_472# 0 0.33241f
C20050 FILLER_0_18_139/a_484_472# 0 0.33241f
C20051 FILLER_0_18_139/a_36_472# 0 0.404746f
C20052 FILLER_0_18_139/a_1468_375# 0 0.233029f
C20053 FILLER_0_18_139/a_1020_375# 0 0.171606f
C20054 FILLER_0_18_139/a_572_375# 0 0.171606f
C20055 FILLER_0_18_139/a_124_375# 0 0.185399f
C20056 _161_ 0 0.592909f
C20057 _162_ 0 0.597238f
C20058 _375_/a_36_68# 0 0.048026f
C20059 trim_val\[0\] 0 0.742779f
C20060 net67 0 1.662327f
C20061 _444_/a_2560_156# 0 0.016968f
C20062 _444_/a_2665_112# 0 0.62251f
C20063 _444_/a_2248_156# 0 0.371662f
C20064 _444_/a_1204_472# 0 0.012971f
C20065 _444_/a_1000_472# 0 0.291735f
C20066 _444_/a_796_472# 0 0.023206f
C20067 _444_/a_1308_423# 0 0.279043f
C20068 _444_/a_448_472# 0 0.684413f
C20069 _444_/a_36_151# 0 1.43589f
C20070 net65 0 0.804072f
C20071 fanout57/a_36_113# 0 0.418095f
C20072 fanout68/a_36_113# 0 0.418095f
C20073 FILLER_0_12_2/a_484_472# 0 0.345058f
C20074 FILLER_0_12_2/a_36_472# 0 0.404746f
C20075 FILLER_0_12_2/a_572_375# 0 0.232991f
C20076 FILLER_0_12_2/a_124_375# 0 0.185089f
C20077 net79 0 1.584979f
C20078 fanout79/a_36_160# 0 0.386641f
C20079 _392_/a_36_68# 0 0.112263f
C20080 FILLER_0_13_228/a_36_472# 0 0.417394f
C20081 FILLER_0_13_228/a_124_375# 0 0.246306f
C20082 FILLER_0_13_206/a_36_472# 0 0.417394f
C20083 FILLER_0_13_206/a_124_375# 0 0.246306f
C20084 FILLER_0_20_177/a_1380_472# 0 0.345058f
C20085 FILLER_0_20_177/a_932_472# 0 0.33241f
C20086 FILLER_0_20_177/a_484_472# 0 0.33241f
C20087 FILLER_0_20_177/a_36_472# 0 0.404746f
C20088 FILLER_0_20_177/a_1468_375# 0 0.233029f
C20089 FILLER_0_20_177/a_1020_375# 0 0.171606f
C20090 FILLER_0_20_177/a_572_375# 0 0.171606f
C20091 FILLER_0_20_177/a_124_375# 0 0.185399f
C20092 _051_ 0 0.349381f
C20093 _213_/a_67_603# 0 0.345683f
C20094 net2 0 0.461658f
C20095 input2/a_36_113# 0 0.418095f
C20096 _129_ 0 0.926508f
C20097 _131_ 0 1.734297f
C20098 _359_/a_36_488# 0 0.101145f
C20099 FILLER_0_11_64/a_36_472# 0 0.417394f
C20100 FILLER_0_11_64/a_124_375# 0 0.246306f
C20101 state\[2\] 0 0.607433f
C20102 net53 0 4.483899f
C20103 _017_ 0 0.334329f
C20104 net70 0 1.238296f
C20105 _428_/a_2560_156# 0 0.016968f
C20106 _428_/a_2665_112# 0 0.62251f
C20107 _428_/a_2248_156# 0 0.371662f
C20108 _428_/a_1204_472# 0 0.012971f
C20109 _428_/a_1000_472# 0 0.291735f
C20110 _428_/a_796_472# 0 0.023206f
C20111 _428_/a_1308_423# 0 0.279043f
C20112 _428_/a_448_472# 0 0.684413f
C20113 _428_/a_36_151# 0 1.43589f
C20114 FILLER_0_5_72/a_1380_472# 0 0.345058f
C20115 FILLER_0_5_72/a_932_472# 0 0.33241f
C20116 FILLER_0_5_72/a_484_472# 0 0.33241f
C20117 FILLER_0_5_72/a_36_472# 0 0.404746f
C20118 FILLER_0_5_72/a_1468_375# 0 0.233029f
C20119 FILLER_0_5_72/a_1020_375# 0 0.171606f
C20120 FILLER_0_5_72/a_572_375# 0 0.171606f
C20121 FILLER_0_5_72/a_124_375# 0 0.185399f
C20122 _376_/a_36_160# 0 0.386641f
C20123 trim_val\[1\] 0 0.683578f
C20124 _445_/a_2560_156# 0 0.016968f
C20125 _445_/a_2665_112# 0 0.62251f
C20126 _445_/a_2248_156# 0 0.371662f
C20127 _445_/a_1204_472# 0 0.012971f
C20128 _445_/a_1000_472# 0 0.291735f
C20129 _445_/a_796_472# 0 0.023206f
C20130 _445_/a_1308_423# 0 0.279043f
C20131 _445_/a_448_472# 0 0.684413f
C20132 _445_/a_36_151# 0 1.43589f
C20133 fanout67/a_36_160# 0 0.386641f
C20134 fanout56/a_36_113# 0 0.418095f
C20135 net78 0 0.686263f
C20136 fanout78/a_36_113# 0 0.418095f
C20137 _174_ 0 0.979741f
C20138 FILLER_0_0_198/a_36_472# 0 0.417394f
C20139 FILLER_0_0_198/a_124_375# 0 0.246306f
C20140 FILLER_0_15_290/a_36_472# 0 0.417394f
C20141 FILLER_0_15_290/a_124_375# 0 0.246306f
C20142 FILLER_0_24_290/a_36_472# 0 0.417394f
C20143 FILLER_0_24_290/a_124_375# 0 0.246306f
C20144 FILLER_0_4_107/a_1380_472# 0 0.345058f
C20145 FILLER_0_4_107/a_932_472# 0 0.33241f
C20146 FILLER_0_4_107/a_484_472# 0 0.33241f
C20147 FILLER_0_4_107/a_36_472# 0 0.404746f
C20148 FILLER_0_4_107/a_1468_375# 0 0.233029f
C20149 FILLER_0_4_107/a_1020_375# 0 0.171606f
C20150 FILLER_0_4_107/a_572_375# 0 0.171606f
C20151 FILLER_0_4_107/a_124_375# 0 0.185399f
C20152 FILLER_0_7_104/a_1380_472# 0 0.345058f
C20153 FILLER_0_7_104/a_932_472# 0 0.33241f
C20154 FILLER_0_7_104/a_484_472# 0 0.33241f
C20155 FILLER_0_7_104/a_36_472# 0 0.404746f
C20156 FILLER_0_7_104/a_1468_375# 0 0.233029f
C20157 FILLER_0_7_104/a_1020_375# 0 0.171606f
C20158 FILLER_0_7_104/a_572_375# 0 0.171606f
C20159 FILLER_0_7_104/a_124_375# 0 0.185399f
C20160 _214_/a_36_160# 0 0.386641f
C20161 net1 0 0.364811f
C20162 input1/a_36_113# 0 0.418095f
C20163 _429_/a_2560_156# 0 0.016968f
C20164 _429_/a_2665_112# 0 0.62251f
C20165 _429_/a_2248_156# 0 0.371662f
C20166 _429_/a_1204_472# 0 0.012971f
C20167 _429_/a_1000_472# 0 0.291735f
C20168 _429_/a_796_472# 0 0.023206f
C20169 _429_/a_1308_423# 0 0.279043f
C20170 _429_/a_448_472# 0 0.684413f
C20171 _429_/a_36_151# 0 1.43589f
C20172 _011_ 0 0.278979f
C20173 _377_/a_36_472# 0 0.031137f
C20174 fanout66/a_36_113# 0 0.418095f
C20175 _035_ 0 0.327801f
C20176 _446_/a_2560_156# 0 0.016968f
C20177 _446_/a_2665_112# 0 0.62251f
C20178 _446_/a_2248_156# 0 0.371662f
C20179 _446_/a_1204_472# 0 0.012971f
C20180 _446_/a_1000_472# 0 0.291735f
C20181 _446_/a_796_472# 0 0.023206f
C20182 _446_/a_1308_423# 0 0.279043f
C20183 _446_/a_448_472# 0 0.684413f
C20184 _446_/a_36_151# 0 1.43589f
C20185 fanout77/a_36_113# 0 0.418095f
C20186 FILLER_0_5_212/a_36_472# 0 0.417394f
C20187 FILLER_0_5_212/a_124_375# 0 0.246306f
C20188 fanout55/a_36_160# 0 0.696445f
C20189 _175_ 0 0.344159f
C20190 _394_/a_1936_472# 0 0.009918f
C20191 _394_/a_718_524# 0 0.005143f
C20192 _394_/a_56_524# 0 0.41096f
C20193 _394_/a_728_93# 0 0.654825f
C20194 _394_/a_1336_472# 0 0.316639f
C20195 FILLER_0_3_172/a_3172_472# 0 0.345058f
C20196 FILLER_0_3_172/a_2724_472# 0 0.33241f
C20197 FILLER_0_3_172/a_2276_472# 0 0.33241f
C20198 FILLER_0_3_172/a_1828_472# 0 0.33241f
C20199 FILLER_0_3_172/a_1380_472# 0 0.33241f
C20200 FILLER_0_3_172/a_932_472# 0 0.33241f
C20201 FILLER_0_3_172/a_484_472# 0 0.33241f
C20202 FILLER_0_3_172/a_36_472# 0 0.404746f
C20203 FILLER_0_3_172/a_3260_375# 0 0.233093f
C20204 FILLER_0_3_172/a_2812_375# 0 0.17167f
C20205 FILLER_0_3_172/a_2364_375# 0 0.17167f
C20206 FILLER_0_3_172/a_1916_375# 0 0.17167f
C20207 FILLER_0_3_172/a_1468_375# 0 0.17167f
C20208 FILLER_0_3_172/a_1020_375# 0 0.17167f
C20209 FILLER_0_3_172/a_572_375# 0 0.17167f
C20210 FILLER_0_3_172/a_124_375# 0 0.185915f
C20211 FILLER_0_17_72/a_3172_472# 0 0.345058f
C20212 FILLER_0_17_72/a_2724_472# 0 0.33241f
C20213 FILLER_0_17_72/a_2276_472# 0 0.33241f
C20214 FILLER_0_17_72/a_1828_472# 0 0.33241f
C20215 FILLER_0_17_72/a_1380_472# 0 0.33241f
C20216 FILLER_0_17_72/a_932_472# 0 0.33241f
C20217 FILLER_0_17_72/a_484_472# 0 0.33241f
C20218 FILLER_0_17_72/a_36_472# 0 0.404746f
C20219 FILLER_0_17_72/a_3260_375# 0 0.233093f
C20220 FILLER_0_17_72/a_2812_375# 0 0.17167f
C20221 FILLER_0_17_72/a_2364_375# 0 0.17167f
C20222 FILLER_0_17_72/a_1916_375# 0 0.17167f
C20223 FILLER_0_17_72/a_1468_375# 0 0.17167f
C20224 FILLER_0_17_72/a_1020_375# 0 0.17167f
C20225 FILLER_0_17_72/a_572_375# 0 0.17167f
C20226 FILLER_0_17_72/a_124_375# 0 0.185915f
C20227 FILLER_0_2_93/a_484_472# 0 0.345058f
C20228 FILLER_0_2_93/a_36_472# 0 0.404746f
C20229 FILLER_0_2_93/a_572_375# 0 0.232991f
C20230 FILLER_0_2_93/a_124_375# 0 0.185089f
C20231 FILLER_0_11_142/a_484_472# 0 0.345058f
C20232 FILLER_0_11_142/a_36_472# 0 0.404746f
C20233 FILLER_0_11_142/a_572_375# 0 0.232991f
C20234 FILLER_0_11_142/a_124_375# 0 0.185089f
C20235 net25 0 1.803174f
C20236 _232_/a_67_603# 0 0.345683f
C20237 net35 0 1.844415f
C20238 mask\[8\] 0 1.276111f
C20239 _301_/a_36_472# 0 0.031137f
C20240 _033_ 0 0.323682f
C20241 _165_ 0 0.331995f
C20242 FILLER_0_3_2/a_36_472# 0 0.417394f
C20243 FILLER_0_3_2/a_124_375# 0 0.246306f
C20244 trim_val\[3\] 0 0.719615f
C20245 _036_ 0 0.369206f
C20246 net68 0 1.735004f
C20247 _447_/a_2560_156# 0 0.016968f
C20248 _447_/a_2665_112# 0 0.62251f
C20249 _447_/a_2248_156# 0 0.371662f
C20250 _447_/a_1204_472# 0 0.012971f
C20251 _447_/a_1000_472# 0 0.291735f
C20252 _447_/a_796_472# 0 0.023206f
C20253 _447_/a_1308_423# 0 0.279043f
C20254 _447_/a_448_472# 0 0.684413f
C20255 _447_/a_36_151# 0 1.43589f
C20256 FILLER_0_19_28/a_484_472# 0 0.345058f
C20257 FILLER_0_19_28/a_36_472# 0 0.404746f
C20258 FILLER_0_19_28/a_572_375# 0 0.232991f
C20259 FILLER_0_19_28/a_124_375# 0 0.185089f
C20260 fanout65/a_36_113# 0 0.418095f
C20261 fanout76/a_36_160# 0 0.386641f
C20262 net54 0 5.456963f
C20263 fanout54/a_36_160# 0 0.696445f
C20264 FILLER_0_4_49/a_484_472# 0 0.345058f
C20265 FILLER_0_4_49/a_36_472# 0 0.404746f
C20266 FILLER_0_4_49/a_572_375# 0 0.232991f
C20267 FILLER_0_4_49/a_124_375# 0 0.185089f
C20268 _176_ 0 0.804011f
C20269 _085_ 0 2.280803f
C20270 _116_ 0 1.959915f
C20271 _395_/a_36_488# 0 0.101145f
C20272 FILLER_0_14_50/a_36_472# 0 0.417394f
C20273 FILLER_0_14_50/a_124_375# 0 0.246306f
C20274 FILLER_0_8_263/a_36_472# 0 0.417394f
C20275 FILLER_0_8_263/a_124_375# 0 0.246306f
C20276 FILLER_0_0_130/a_36_472# 0 0.417394f
C20277 FILLER_0_0_130/a_124_375# 0 0.246306f
C20278 FILLER_0_16_255/a_36_472# 0 0.417394f
C20279 FILLER_0_16_255/a_124_375# 0 0.246306f
C20280 FILLER_0_7_59/a_484_472# 0 0.345058f
C20281 FILLER_0_7_59/a_36_472# 0 0.404746f
C20282 FILLER_0_7_59/a_572_375# 0 0.232991f
C20283 FILLER_0_7_59/a_124_375# 0 0.185089f
C20284 ctlp[2] 0 0.17528f
C20285 output19/a_224_472# 0 2.38465f
C20286 FILLER_0_7_146/a_36_472# 0 0.417394f
C20287 FILLER_0_7_146/a_124_375# 0 0.246306f
C20288 _216_/a_67_603# 0 0.345683f
C20289 FILLER_0_15_116/a_484_472# 0 0.345058f
C20290 FILLER_0_15_116/a_36_472# 0 0.404746f
C20291 FILLER_0_15_116/a_572_375# 0 0.232991f
C20292 FILLER_0_15_116/a_124_375# 0 0.185089f
C20293 _063_ 0 0.370155f
C20294 _233_/a_36_160# 0 0.386641f
C20295 FILLER_0_21_28/a_3172_472# 0 0.345058f
C20296 FILLER_0_21_28/a_2724_472# 0 0.33241f
C20297 FILLER_0_21_28/a_2276_472# 0 0.33241f
C20298 FILLER_0_21_28/a_1828_472# 0 0.33241f
C20299 FILLER_0_21_28/a_1380_472# 0 0.33241f
C20300 FILLER_0_21_28/a_932_472# 0 0.33241f
C20301 FILLER_0_21_28/a_484_472# 0 0.33241f
C20302 FILLER_0_21_28/a_36_472# 0 0.404746f
C20303 FILLER_0_21_28/a_3260_375# 0 0.233093f
C20304 FILLER_0_21_28/a_2812_375# 0 0.17167f
C20305 FILLER_0_21_28/a_2364_375# 0 0.17167f
C20306 FILLER_0_21_28/a_1916_375# 0 0.17167f
C20307 FILLER_0_21_28/a_1468_375# 0 0.17167f
C20308 FILLER_0_21_28/a_1020_375# 0 0.17167f
C20309 FILLER_0_21_28/a_572_375# 0 0.17167f
C20310 FILLER_0_21_28/a_124_375# 0 0.185915f
C20311 _110_ 0 0.323912f
C20312 _379_/a_36_472# 0 0.031137f
C20313 trim_val\[4\] 0 0.662409f
C20314 net76 0 1.454269f
C20315 _448_/a_2560_156# 0 0.016968f
C20316 _448_/a_2665_112# 0 0.62251f
C20317 _448_/a_2248_156# 0 0.371662f
C20318 _448_/a_1204_472# 0 0.012971f
C20319 _448_/a_1000_472# 0 0.291735f
C20320 _448_/a_796_472# 0 0.023206f
C20321 _448_/a_1308_423# 0 0.279043f
C20322 _448_/a_448_472# 0 0.684413f
C20323 _448_/a_36_151# 0 1.43589f
C20324 fanout64/a_36_160# 0 0.386641f
C20325 fanout75/a_36_113# 0 0.418095f
C20326 _250_/a_36_68# 0 0.69549f
C20327 net56 0 0.843396f
C20328 fanout53/a_36_160# 0 0.696445f
C20329 _177_ 0 0.358286f
C20330 result[2] 0 0.230851f
C20331 net29 0 1.802718f
C20332 output29/a_224_472# 0 2.38465f
C20333 ctlp[1] 0 0.17418f
C20334 output18/a_224_472# 0 2.38465f
C20335 FILLER_0_14_181/a_36_472# 0 0.417394f
C20336 FILLER_0_14_181/a_124_375# 0 0.246306f
C20337 _052_ 0 0.569133f
C20338 _217_/a_36_160# 0 0.386641f
C20339 net44 0 1.407054f
C20340 _303_/a_36_472# 0 0.031137f
C20341 en_co_clk 0 0.346872f
C20342 net55 0 5.119958f
C20343 net72 0 1.366255f
C20344 _449_/a_2560_156# 0 0.016968f
C20345 _449_/a_2665_112# 0 0.62251f
C20346 _449_/a_2248_156# 0 0.371662f
C20347 _449_/a_1204_472# 0 0.012971f
C20348 _449_/a_1000_472# 0 0.291735f
C20349 _449_/a_796_472# 0 0.023206f
C20350 _449_/a_1308_423# 0 0.279043f
C20351 _449_/a_448_472# 0 0.684413f
C20352 _449_/a_36_151# 0 1.43589f
C20353 fanout52/a_36_160# 0 0.696445f
C20354 net82 0 0.706042f
C20355 fanout74/a_36_113# 0 0.418095f
C20356 FILLER_0_10_28/a_36_472# 0 0.417394f
C20357 FILLER_0_10_28/a_124_375# 0 0.246306f
C20358 mask\[0\] 0 2.242948f
C20359 _320_/a_36_472# 0 0.137725f
C20360 fanout63/a_36_160# 0 0.696445f
C20361 FILLER_0_14_81/a_36_472# 0 0.417394f
C20362 FILLER_0_14_81/a_124_375# 0 0.246306f
C20363 _397_/a_36_472# 0 0.031137f
C20364 FILLER_0_13_212/a_1380_472# 0 0.345058f
C20365 FILLER_0_13_212/a_932_472# 0 0.33241f
C20366 FILLER_0_13_212/a_484_472# 0 0.33241f
C20367 FILLER_0_13_212/a_36_472# 0 0.404746f
C20368 FILLER_0_13_212/a_1468_375# 0 0.233029f
C20369 FILLER_0_13_212/a_1020_375# 0 0.171606f
C20370 FILLER_0_13_212/a_572_375# 0 0.171606f
C20371 FILLER_0_13_212/a_124_375# 0 0.185399f
C20372 trim[1] 0 0.793787f
C20373 net39 0 1.445128f
C20374 output39/a_224_472# 0 2.38465f
C20375 result[1] 0 0.229507f
C20376 net28 0 1.759728f
C20377 output28/a_224_472# 0 2.38465f
C20378 ctlp[0] 0 1.002286f
C20379 output17/a_224_472# 0 2.38465f
C20380 FILLER_0_16_37/a_36_472# 0 0.417394f
C20381 FILLER_0_16_37/a_124_375# 0 0.246306f
C20382 net26 0 1.671545f
C20383 _064_ 0 0.581481f
C20384 trim_val\[2\] 0 0.65354f
C20385 trim_mask\[2\] 0 0.92551f
C20386 _235_/a_67_603# 0 0.345683f
C20387 _013_ 0 0.48783f
C20388 _111_ 0 0.369652f
C20389 FILLER_0_18_177/a_3172_472# 0 0.345058f
C20390 FILLER_0_18_177/a_2724_472# 0 0.33241f
C20391 FILLER_0_18_177/a_2276_472# 0 0.33241f
C20392 FILLER_0_18_177/a_1828_472# 0 0.33241f
C20393 FILLER_0_18_177/a_1380_472# 0 0.33241f
C20394 FILLER_0_18_177/a_932_472# 0 0.33241f
C20395 FILLER_0_18_177/a_484_472# 0 0.33241f
C20396 FILLER_0_18_177/a_36_472# 0 0.404746f
C20397 FILLER_0_18_177/a_3260_375# 0 0.233093f
C20398 FILLER_0_18_177/a_2812_375# 0 0.17167f
C20399 FILLER_0_18_177/a_2364_375# 0 0.17167f
C20400 FILLER_0_18_177/a_1916_375# 0 0.17167f
C20401 FILLER_0_18_177/a_1468_375# 0 0.17167f
C20402 FILLER_0_18_177/a_1020_375# 0 0.17167f
C20403 FILLER_0_18_177/a_572_375# 0 0.17167f
C20404 FILLER_0_18_177/a_124_375# 0 0.185915f
C20405 FILLER_0_18_100/a_36_472# 0 0.417394f
C20406 FILLER_0_18_100/a_124_375# 0 0.246306f
C20407 _073_ 0 0.953711f
C20408 _126_ 0 2.036767f
C20409 _069_ 0 2.034557f
C20410 _321_/a_170_472# 0 0.077257f
C20411 fanout51/a_36_113# 0 0.418095f
C20412 net62 0 4.932099f
C20413 fanout62/a_36_160# 0 0.696445f
C20414 fanout73/a_36_113# 0 0.418095f
C20415 FILLER_0_19_47/a_484_472# 0 0.345058f
C20416 FILLER_0_19_47/a_36_472# 0 0.404746f
C20417 FILLER_0_19_47/a_572_375# 0 0.232991f
C20418 FILLER_0_19_47/a_124_375# 0 0.185089f
C20419 FILLER_0_14_91/a_484_472# 0 0.345058f
C20420 FILLER_0_14_91/a_36_472# 0 0.404746f
C20421 FILLER_0_14_91/a_572_375# 0 0.232991f
C20422 FILLER_0_14_91/a_124_375# 0 0.185089f
C20423 FILLER_0_10_214/a_36_472# 0 0.417394f
C20424 FILLER_0_10_214/a_124_375# 0 0.246306f
C20425 FILLER_0_10_247/a_36_472# 0 0.417394f
C20426 FILLER_0_10_247/a_124_375# 0 0.246306f
C20427 _178_ 0 1.252435f
C20428 _398_/a_36_113# 0 0.418095f
C20429 FILLER_0_16_241/a_36_472# 0 0.417394f
C20430 FILLER_0_16_241/a_124_375# 0 0.246306f
C20431 trim[0] 0 0.796081f
C20432 net38 0 1.529392f
C20433 output38/a_224_472# 0 2.38465f
C20434 ctln[9] 0 0.904836f
C20435 net16 0 1.295744f
C20436 output16/a_224_472# 0 2.38465f
C20437 result[0] 0 0.56622f
C20438 output27/a_224_472# 0 2.38465f
C20439 _219_/a_36_160# 0 0.386641f
C20440 FILLER_0_20_193/a_484_472# 0 0.345058f
C20441 FILLER_0_20_193/a_36_472# 0 0.404746f
C20442 FILLER_0_20_193/a_572_375# 0 0.232991f
C20443 FILLER_0_20_193/a_124_375# 0 0.185089f
C20444 _236_/a_36_160# 0 0.696445f
C20445 _112_ 0 0.308886f
C20446 _305_/a_36_159# 0 0.374116f
C20447 _074_ 0 1.813232f
C20448 _253_/a_36_68# 0 0.061249f
C20449 net50 0 4.486121f
C20450 net52 0 3.536016f
C20451 fanout50/a_36_160# 0 0.696445f
C20452 FILLER_0_10_37/a_36_472# 0 0.417394f
C20453 FILLER_0_10_37/a_124_375# 0 0.246306f
C20454 fanout72/a_36_113# 0 0.418095f
C20455 fanout61/a_36_113# 0 0.418095f
C20456 _128_ 0 0.447252f
C20457 _127_ 0 1.291729f
C20458 _322_/a_848_380# 0 0.40208f
C20459 _322_/a_124_24# 0 0.591898f
C20460 _088_ 0 0.457961f
C20461 _079_ 0 1.114894f
C20462 _087_ 0 0.601674f
C20463 _270_/a_36_472# 0 0.031137f
C20464 FILLER_0_4_123/a_36_472# 0 0.417394f
C20465 FILLER_0_4_123/a_124_375# 0 0.246306f
C20466 FILLER_0_17_218/a_484_472# 0 0.345058f
C20467 FILLER_0_17_218/a_36_472# 0 0.404746f
C20468 FILLER_0_17_218/a_572_375# 0 0.232991f
C20469 FILLER_0_17_218/a_124_375# 0 0.185089f
C20470 sample 0 0.508149f
C20471 output37/a_224_472# 0 2.38465f
C20472 valid 0 0.272072f
C20473 net48 0 1.219262f
C20474 output48/a_224_472# 0 2.38465f
C20475 ctln[8] 0 1.547984f
C20476 net15 0 1.440851f
C20477 output15/a_224_472# 0 2.38465f
C20478 ctlp[9] 0 0.73349f
C20479 output26/a_224_472# 0 2.38465f
C20480 FILLER_0_16_57/a_1380_472# 0 0.345058f
C20481 FILLER_0_16_57/a_932_472# 0 0.33241f
C20482 FILLER_0_16_57/a_484_472# 0 0.33241f
C20483 FILLER_0_16_57/a_36_472# 0 0.404746f
C20484 FILLER_0_16_57/a_1468_375# 0 0.233029f
C20485 FILLER_0_16_57/a_1020_375# 0 0.171606f
C20486 FILLER_0_16_57/a_572_375# 0 0.171606f
C20487 FILLER_0_16_57/a_124_375# 0 0.185399f
C20488 _306_/a_36_68# 0 0.69549f
C20489 _072_ 0 2.604301f
C20490 fanout82/a_36_113# 0 0.418095f
C20491 _015_ 0 0.406653f
C20492 _323_/a_36_113# 0 0.418095f
C20493 net60 0 5.024503f
C20494 net61 0 1.666523f
C20495 fanout60/a_36_160# 0 0.696445f
C20496 fanout71/a_36_113# 0 0.418095f
C20497 FILLER_0_6_239/a_36_472# 0 0.417394f
C20498 FILLER_0_6_239/a_124_375# 0 0.246306f
C20499 FILLER_0_4_99/a_36_472# 0 0.417394f
C20500 FILLER_0_4_99/a_124_375# 0 0.246306f
C20501 net57 0 1.383718f
C20502 FILLER_0_10_256/a_36_472# 0 0.417394f
C20503 FILLER_0_10_256/a_124_375# 0 0.246306f
C20504 cal_itt\[3\] 0 1.854962f
C20505 _340_/a_36_160# 0 0.386641f
C20506 FILLER_0_4_177/a_484_472# 0 0.345058f
C20507 FILLER_0_4_177/a_36_472# 0 0.404746f
C20508 FILLER_0_4_177/a_572_375# 0 0.232991f
C20509 FILLER_0_4_177/a_124_375# 0 0.185089f
C20510 FILLER_0_4_144/a_484_472# 0 0.345058f
C20511 FILLER_0_4_144/a_36_472# 0 0.404746f
C20512 FILLER_0_4_144/a_572_375# 0 0.232991f
C20513 FILLER_0_4_144/a_124_375# 0 0.185089f
C20514 ctln[7] 0 1.265946f
C20515 output14/a_224_472# 0 2.38465f
C20516 result[9] 0 0.8197f
C20517 output36/a_224_472# 0 2.38465f
C20518 trimb[4] 0 0.752332f
C20519 output47/a_224_472# 0 2.38465f
C20520 ctlp[8] 0 1.136333f
C20521 output25/a_224_472# 0 2.38465f
C20522 FILLER_0_12_136/a_1380_472# 0 0.345058f
C20523 FILLER_0_12_136/a_932_472# 0 0.33241f
C20524 FILLER_0_12_136/a_484_472# 0 0.33241f
C20525 FILLER_0_12_136/a_36_472# 0 0.404746f
C20526 FILLER_0_12_136/a_1468_375# 0 0.233029f
C20527 FILLER_0_12_136/a_1020_375# 0 0.171606f
C20528 FILLER_0_12_136/a_572_375# 0 0.171606f
C20529 FILLER_0_12_136/a_124_375# 0 0.185399f
C20530 FILLER_0_16_89/a_1380_472# 0 0.345058f
C20531 FILLER_0_16_89/a_932_472# 0 0.33241f
C20532 FILLER_0_16_89/a_484_472# 0 0.33241f
C20533 FILLER_0_16_89/a_36_472# 0 0.404746f
C20534 FILLER_0_16_89/a_1468_375# 0 0.233029f
C20535 FILLER_0_16_89/a_1020_375# 0 0.171606f
C20536 FILLER_0_16_89/a_572_375# 0 0.171606f
C20537 FILLER_0_16_89/a_124_375# 0 0.185399f
C20538 FILLER_0_21_125/a_484_472# 0 0.345058f
C20539 FILLER_0_21_125/a_36_472# 0 0.404746f
C20540 FILLER_0_21_125/a_572_375# 0 0.232991f
C20541 FILLER_0_21_125/a_124_375# 0 0.185089f
C20542 _238_/a_67_603# 0 0.345683f
C20543 _096_ 0 2.205532f
C20544 _093_ 0 1.893313f
C20545 FILLER_0_19_55/a_36_472# 0 0.417394f
C20546 FILLER_0_19_55/a_124_375# 0 0.246306f
C20547 net81 0 1.738987f
C20548 fanout81/a_36_160# 0 0.386641f
C20549 _057_ 0 1.600886f
C20550 _255_/a_224_552# 0 1.31114f
C20551 net73 0 1.058857f
C20552 fanout70/a_36_113# 0 0.418095f
C20553 _003_ 0 0.3064f
C20554 _089_ 0 0.36777f
C20555 _272_/a_36_472# 0 0.031137f
C20556 _187_ 0 0.311229f
C20557 _410_/a_36_68# 0 0.112263f
C20558 _141_ 0 1.249289f
C20559 mask\[3\] 0 1.26722f
C20560 _341_/a_49_472# 0 0.054843f
C20561 cal 0 0.793393f
C20562 FILLER_0_7_195/a_36_472# 0 0.417394f
C20563 FILLER_0_7_195/a_124_375# 0 0.246306f
C20564 FILLER_0_7_162/a_36_472# 0 0.417394f
C20565 FILLER_0_7_162/a_124_375# 0 0.246306f
C20566 ctln[6] 0 1.451644f
C20567 output13/a_224_472# 0 2.38465f
C20568 FILLER_0_18_2/a_3172_472# 0 0.345058f
C20569 FILLER_0_18_2/a_2724_472# 0 0.33241f
C20570 FILLER_0_18_2/a_2276_472# 0 0.33241f
C20571 FILLER_0_18_2/a_1828_472# 0 0.33241f
C20572 FILLER_0_18_2/a_1380_472# 0 0.33241f
C20573 FILLER_0_18_2/a_932_472# 0 0.33241f
C20574 FILLER_0_18_2/a_484_472# 0 0.33241f
C20575 FILLER_0_18_2/a_36_472# 0 0.404746f
C20576 FILLER_0_18_2/a_3260_375# 0 0.233093f
C20577 FILLER_0_18_2/a_2812_375# 0 0.17167f
C20578 FILLER_0_18_2/a_2364_375# 0 0.17167f
C20579 FILLER_0_18_2/a_1916_375# 0 0.17167f
C20580 FILLER_0_18_2/a_1468_375# 0 0.17167f
C20581 FILLER_0_18_2/a_1020_375# 0 0.17167f
C20582 FILLER_0_18_2/a_572_375# 0 0.17167f
C20583 FILLER_0_18_2/a_124_375# 0 0.185915f
C20584 trimb[3] 0 0.34698f
C20585 net46 0 1.13395f
C20586 output46/a_224_472# 0 2.38465f
C20587 result[8] 0 0.68837f
C20588 output35/a_224_472# 0 2.38465f
C20589 ctlp[7] 0 0.83567f
C20590 output24/a_224_472# 0 2.38465f
C20591 FILLER_0_8_107/a_36_472# 0 0.417394f
C20592 FILLER_0_8_107/a_124_375# 0 0.246306f
C20593 FILLER_0_12_124/a_36_472# 0 0.417394f
C20594 FILLER_0_12_124/a_124_375# 0 0.246306f
C20595 net41 0 1.746759f
C20596 _065_ 0 0.523724f
C20597 _239_/a_36_160# 0 0.696445f
C20598 FILLER_0_1_98/a_36_472# 0 0.417394f
C20599 FILLER_0_1_98/a_124_375# 0 0.246306f
C20600 _115_ 0 1.281516f
C20601 _114_ 0 2.293579f
C20602 _308_/a_848_380# 0 0.40208f
C20603 _308_/a_124_24# 0 0.591898f
C20604 _256_/a_36_68# 0 0.063181f
C20605 FILLER_0_10_78/a_1380_472# 0 0.345058f
C20606 FILLER_0_10_78/a_932_472# 0 0.33241f
C20607 FILLER_0_10_78/a_484_472# 0 0.33241f
C20608 FILLER_0_10_78/a_36_472# 0 0.404746f
C20609 FILLER_0_10_78/a_1468_375# 0 0.233029f
C20610 FILLER_0_10_78/a_1020_375# 0 0.171606f
C20611 FILLER_0_10_78/a_572_375# 0 0.171606f
C20612 FILLER_0_10_78/a_124_375# 0 0.185399f
C20613 _130_ 0 0.304085f
C20614 net80 0 1.375599f
C20615 fanout80/a_36_113# 0 0.418095f
C20616 net58 0 5.308423f
C20617 _000_ 0 0.382358f
C20618 net75 0 1.474299f
C20619 _411_/a_2560_156# 0 0.016968f
C20620 _411_/a_2665_112# 0 0.62251f
C20621 _411_/a_2248_156# 0 0.371662f
C20622 _411_/a_1204_472# 0 0.012971f
C20623 _411_/a_1000_472# 0 0.291735f
C20624 _411_/a_796_472# 0 0.023206f
C20625 _411_/a_1308_423# 0 0.279043f
C20626 _411_/a_448_472# 0 0.684413f
C20627 _411_/a_36_151# 0 1.43589f
C20628 state\[0\] 0 0.680109f
C20629 _273_/a_36_68# 0 0.69549f
C20630 _142_ 0 0.324372f
C20631 FILLER_0_9_223/a_484_472# 0 0.345058f
C20632 FILLER_0_9_223/a_36_472# 0 0.404746f
C20633 FILLER_0_9_223/a_572_375# 0 0.232991f
C20634 FILLER_0_9_223/a_124_375# 0 0.185089f
C20635 FILLER_0_4_197/a_1380_472# 0 0.345058f
C20636 FILLER_0_4_197/a_932_472# 0 0.33241f
C20637 FILLER_0_4_197/a_484_472# 0 0.33241f
C20638 FILLER_0_4_197/a_36_472# 0 0.404746f
C20639 FILLER_0_4_197/a_1468_375# 0 0.233029f
C20640 FILLER_0_4_197/a_1020_375# 0 0.171606f
C20641 FILLER_0_4_197/a_572_375# 0 0.171606f
C20642 FILLER_0_4_197/a_124_375# 0 0.185399f
C20643 FILLER_0_17_226/a_36_472# 0 0.417394f
C20644 FILLER_0_17_226/a_124_375# 0 0.246306f
C20645 FILLER_0_5_109/a_484_472# 0 0.345058f
C20646 FILLER_0_5_109/a_36_472# 0 0.404746f
C20647 FILLER_0_5_109/a_572_375# 0 0.232991f
C20648 FILLER_0_5_109/a_124_375# 0 0.185089f
C20649 ctln[5] 0 1.585113f
C20650 output12/a_224_472# 0 2.38465f
C20651 result[7] 0 0.24756f
C20652 net34 0 1.724665f
C20653 output34/a_224_472# 0 2.38465f
C20654 trimb[2] 0 0.839614f
C20655 net45 0 1.12041f
C20656 output45/a_224_472# 0 2.38465f
C20657 ctlp[6] 0 1.243017f
C20658 output23/a_224_472# 0 2.38465f
C20659 FILLER_0_15_142/a_484_472# 0 0.345058f
C20660 FILLER_0_15_142/a_36_472# 0 0.404746f
C20661 FILLER_0_15_142/a_572_375# 0 0.232991f
C20662 FILLER_0_15_142/a_124_375# 0 0.185089f
C20663 _077_ 0 1.645892f
C20664 _075_ 0 0.374516f
C20665 _257_/a_36_472# 0 0.031137f
C20666 _326_/a_36_160# 0 0.696445f
C20667 _412_/a_2560_156# 0 0.016968f
C20668 _412_/a_2665_112# 0 0.62251f
C20669 _412_/a_2248_156# 0 0.371662f
C20670 _412_/a_1204_472# 0 0.012971f
C20671 _412_/a_1000_472# 0 0.291735f
C20672 _412_/a_796_472# 0 0.023206f
C20673 _412_/a_1308_423# 0 0.279043f
C20674 _412_/a_448_472# 0 0.684413f
C20675 _412_/a_36_151# 0 1.43589f
C20676 _091_ 0 1.841339f
C20677 _274_/a_36_68# 0 0.063181f
C20678 _143_ 0 0.329289f
C20679 mask\[4\] 0 1.300438f
C20680 _343_/a_49_472# 0 0.054843f
C20681 FILLER_0_13_65/a_36_472# 0 0.417394f
C20682 FILLER_0_13_65/a_124_375# 0 0.246306f
C20683 _360_/a_36_160# 0 0.386641f
C20684 FILLER_0_4_185/a_36_472# 0 0.417394f
C20685 FILLER_0_4_185/a_124_375# 0 0.246306f
C20686 FILLER_0_4_152/a_36_472# 0 0.417394f
C20687 FILLER_0_4_152/a_124_375# 0 0.246306f
C20688 _291_/a_36_160# 0 0.386641f
C20689 ctln[2] 0 1.833091f
C20690 output9/a_224_472# 0 2.38465f
C20691 ctln[4] 0 1.461847f
C20692 output11/a_224_472# 0 2.38465f
C20693 trimb[1] 0 0.378532f
C20694 output44/a_224_472# 0 2.38465f
C20695 result[6] 0 0.19512f
C20696 output33/a_224_472# 0 2.38465f
C20697 ctlp[5] 0 1.282822f
C20698 output22/a_224_472# 0 2.38465f
C20699 FILLER_0_8_127/a_36_472# 0 0.417394f
C20700 FILLER_0_8_127/a_124_375# 0 0.246306f
C20701 FILLER_0_8_138/a_36_472# 0 0.417394f
C20702 FILLER_0_8_138/a_124_375# 0 0.246306f
C20703 FILLER_0_21_133/a_36_472# 0 0.417394f
C20704 FILLER_0_21_133/a_124_375# 0 0.246306f
C20705 FILLER_0_24_130/a_36_472# 0 0.417394f
C20706 FILLER_0_24_130/a_124_375# 0 0.246306f
C20707 FILLER_0_18_171/a_36_472# 0 0.417394f
C20708 FILLER_0_18_171/a_124_375# 0 0.246306f
C20709 _258_/a_36_160# 0 0.386641f
C20710 _016_ 0 0.314121f
C20711 _327_/a_36_472# 0 0.031137f
C20712 _189_/a_67_603# 0 0.345683f
C20713 FILLER_0_24_63/a_36_472# 0 0.417394f
C20714 FILLER_0_24_63/a_124_375# 0 0.246306f
C20715 FILLER_0_24_96/a_36_472# 0 0.417394f
C20716 FILLER_0_24_96/a_124_375# 0 0.246306f
C20717 cal_itt\[2\] 0 1.473514f
C20718 _002_ 0 0.289553f
C20719 _413_/a_2560_156# 0 0.016968f
C20720 _413_/a_2665_112# 0 0.62251f
C20721 _413_/a_2248_156# 0 0.371662f
C20722 _413_/a_1204_472# 0 0.012971f
C20723 _413_/a_1000_472# 0 0.291735f
C20724 _413_/a_796_472# 0 0.023206f
C20725 _413_/a_1308_423# 0 0.279043f
C20726 _413_/a_448_472# 0 0.684413f
C20727 _413_/a_36_151# 0 1.43589f
C20728 _092_ 0 0.680239f
C20729 FILLER_0_7_72/a_3172_472# 0 0.345058f
C20730 FILLER_0_7_72/a_2724_472# 0 0.33241f
C20731 FILLER_0_7_72/a_2276_472# 0 0.33241f
C20732 FILLER_0_7_72/a_1828_472# 0 0.33241f
C20733 FILLER_0_7_72/a_1380_472# 0 0.33241f
C20734 FILLER_0_7_72/a_932_472# 0 0.33241f
C20735 FILLER_0_7_72/a_484_472# 0 0.33241f
C20736 FILLER_0_7_72/a_36_472# 0 0.404746f
C20737 FILLER_0_7_72/a_3260_375# 0 0.233093f
C20738 FILLER_0_7_72/a_2812_375# 0 0.17167f
C20739 FILLER_0_7_72/a_2364_375# 0 0.17167f
C20740 FILLER_0_7_72/a_1916_375# 0 0.17167f
C20741 FILLER_0_7_72/a_1468_375# 0 0.17167f
C20742 FILLER_0_7_72/a_1020_375# 0 0.17167f
C20743 FILLER_0_7_72/a_572_375# 0 0.17167f
C20744 FILLER_0_7_72/a_124_375# 0 0.185915f
C20745 _086_ 0 2.45259f
C20746 _119_ 0 1.237181f
C20747 net63 0 5.362473f
C20748 _430_/a_2560_156# 0 0.016968f
C20749 _430_/a_2665_112# 0 0.62251f
C20750 _430_/a_2248_156# 0 0.371662f
C20751 _430_/a_1204_472# 0 0.012971f
C20752 _430_/a_1000_472# 0 0.291735f
C20753 _430_/a_796_472# 0 0.023206f
C20754 _430_/a_1308_423# 0 0.279043f
C20755 _430_/a_448_472# 0 0.684413f
C20756 _430_/a_36_151# 0 1.43589f
C20757 _292_/a_36_160# 0 0.386641f
C20758 comp 0 1.022965f
C20759 ctln[1] 0 1.11973f
C20760 output8/a_224_472# 0 2.38465f
C20761 ctln[3] 0 0.835391f
C20762 output10/a_224_472# 0 2.38465f
C20763 result[5] 0 0.206867f
C20764 net32 0 1.78884f
C20765 output32/a_224_472# 0 2.38465f
C20766 trimb[0] 0 0.847787f
C20767 output43/a_224_472# 0 2.38465f
C20768 ctlp[4] 0 0.37565f
C20769 output21/a_224_472# 0 2.38465f
C20770 _053_ 0 1.705161f
C20771 FILLER_0_16_107/a_484_472# 0 0.345058f
C20772 FILLER_0_16_107/a_36_472# 0 0.404746f
C20773 FILLER_0_16_107/a_572_375# 0 0.232991f
C20774 FILLER_0_16_107/a_124_375# 0 0.185089f
C20775 FILLER_0_3_204/a_36_472# 0 0.417394f
C20776 FILLER_0_3_204/a_124_375# 0 0.246306f
C20777 FILLER_0_9_28/a_3172_472# 0 0.345058f
C20778 FILLER_0_9_28/a_2724_472# 0 0.33241f
C20779 FILLER_0_9_28/a_2276_472# 0 0.33241f
C20780 FILLER_0_9_28/a_1828_472# 0 0.33241f
C20781 FILLER_0_9_28/a_1380_472# 0 0.33241f
C20782 FILLER_0_9_28/a_932_472# 0 0.33241f
C20783 FILLER_0_9_28/a_484_472# 0 0.33241f
C20784 FILLER_0_9_28/a_36_472# 0 0.404746f
C20785 FILLER_0_9_28/a_3260_375# 0 0.233093f
C20786 FILLER_0_9_28/a_2812_375# 0 0.17167f
C20787 FILLER_0_9_28/a_2364_375# 0 0.17167f
C20788 FILLER_0_9_28/a_1916_375# 0 0.17167f
C20789 FILLER_0_9_28/a_1468_375# 0 0.17167f
C20790 FILLER_0_9_28/a_1020_375# 0 0.17167f
C20791 FILLER_0_9_28/a_572_375# 0 0.17167f
C20792 FILLER_0_9_28/a_124_375# 0 0.185915f
C20793 _132_ 0 1.491425f
C20794 _328_/a_36_113# 0 0.418095f
C20795 _414_/a_2560_156# 0 0.016968f
C20796 _414_/a_2665_112# 0 0.62251f
C20797 _414_/a_2248_156# 0 0.371662f
C20798 _414_/a_1204_472# 0 0.012971f
C20799 _414_/a_1000_472# 0 0.291735f
C20800 _414_/a_796_472# 0 0.023206f
C20801 _414_/a_1308_423# 0 0.279043f
C20802 _414_/a_448_472# 0 0.684413f
C20803 _414_/a_36_151# 0 1.43589f
C20804 _276_/a_36_160# 0 0.386641f
C20805 _144_ 0 1.173846f
C20806 _345_/a_36_160# 0 0.386641f
C20807 _155_ 0 0.638535f
C20808 _020_ 0 0.316793f
C20809 _431_/a_2560_156# 0 0.016968f
C20810 _431_/a_2665_112# 0 0.62251f
C20811 _431_/a_2248_156# 0 0.371662f
C20812 _431_/a_1204_472# 0 0.012971f
C20813 _431_/a_1000_472# 0 0.291735f
C20814 _431_/a_796_472# 0 0.023206f
C20815 _431_/a_1308_423# 0 0.279043f
C20816 _431_/a_448_472# 0 0.684413f
C20817 _431_/a_36_151# 0 1.43589f
C20818 _105_ 0 1.21281f
C20819 _293_/a_36_472# 0 0.031137f
C20820 FILLER_0_5_128/a_484_472# 0 0.345058f
C20821 FILLER_0_5_128/a_36_472# 0 0.404746f
C20822 FILLER_0_5_128/a_572_375# 0 0.232991f
C20823 FILLER_0_5_128/a_124_375# 0 0.185089f
C20824 FILLER_0_5_117/a_36_472# 0 0.417394f
C20825 FILLER_0_5_117/a_124_375# 0 0.246306f
C20826 ctln[0] 0 1.423102f
C20827 net7 0 1.174913f
C20828 output7/a_224_472# 0 2.38465f
C20829 trim[4] 0 0.763069f
C20830 output42/a_224_472# 0 2.38465f
C20831 result[4] 0 0.038878f
C20832 net31 0 1.912935f
C20833 output31/a_224_472# 0 2.38465f
C20834 ctlp[3] 0 1.14968f
C20835 output20/a_224_472# 0 2.38465f
C20836 FILLER_0_16_73/a_484_472# 0 0.345058f
C20837 FILLER_0_16_73/a_36_472# 0 0.404746f
C20838 FILLER_0_16_73/a_572_375# 0 0.232991f
C20839 FILLER_0_16_73/a_124_375# 0 0.185089f
C20840 FILLER_0_21_142/a_484_472# 0 0.345058f
C20841 FILLER_0_21_142/a_36_472# 0 0.404746f
C20842 FILLER_0_21_142/a_572_375# 0 0.232991f
C20843 FILLER_0_21_142/a_124_375# 0 0.185089f
C20844 FILLER_0_15_150/a_36_472# 0 0.417394f
C20845 FILLER_0_15_150/a_124_375# 0 0.246306f
C20846 FILLER_0_19_125/a_36_472# 0 0.417394f
C20847 FILLER_0_19_125/a_124_375# 0 0.246306f
C20848 net10 0 1.480101f
C20849 net20 0 2.034189f
C20850 _277_/a_36_160# 0 0.386641f
C20851 net27 0 2.023744f
C20852 _004_ 0 0.390107f
C20853 _415_/a_2560_156# 0 0.016968f
C20854 _415_/a_2665_112# 0 0.62251f
C20855 _415_/a_2248_156# 0 0.371662f
C20856 _415_/a_1204_472# 0 0.012971f
C20857 _415_/a_1000_472# 0 0.291735f
C20858 _415_/a_796_472# 0 0.023206f
C20859 _415_/a_1308_423# 0 0.279043f
C20860 _415_/a_448_472# 0 0.684413f
C20861 _415_/a_36_151# 0 1.43589f
C20862 mask\[5\] 0 1.334568f
C20863 _346_/a_49_472# 0 0.054843f
C20864 _028_ 0 0.386029f
C20865 _363_/a_36_68# 0 0.150048f
C20866 _021_ 0 0.316776f
C20867 _432_/a_2560_156# 0 0.016968f
C20868 _432_/a_2665_112# 0 0.62251f
C20869 _432_/a_2248_156# 0 0.371662f
C20870 _432_/a_1204_472# 0 0.012971f
C20871 _432_/a_1000_472# 0 0.291735f
C20872 _432_/a_796_472# 0 0.023206f
C20873 _432_/a_1308_423# 0 0.279043f
C20874 _432_/a_448_472# 0 0.684413f
C20875 _432_/a_36_151# 0 1.43589f
C20876 _008_ 0 0.423631f
C20877 _104_ 0 1.435764f
C20878 _106_ 0 0.378703f
C20879 FILLER_0_17_200/a_484_472# 0 0.345058f
C20880 FILLER_0_17_200/a_36_472# 0 0.404746f
C20881 FILLER_0_17_200/a_572_375# 0 0.232991f
C20882 FILLER_0_17_200/a_124_375# 0 0.185089f
.ends

.subckt saradc vss vdd vinp vinn result[0] result[1] result[2] result[3] result[4]
+ result[5] result[6] result[7] result[8] result[9] valid cal en clk rstn
Xlatch_0 latch_0/Q latch_0/Qn latch_0/R latch_0/S latch_0/tutyuu1 latch_0/tutyuu2
+ vdd vdd latch
Xbuffer_0 sarlogic_0/clkc buffer_0/buf_out buffer_0/inv2_0/inv_in vdd buffer
Xdacp_0 vinp vdd dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9 dacp_0/ctl10 dacp_0/sample dacp_0/ctl2
+ dacp_0/ctl1 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/ndum dacp_0/ctl4 dacp_0/ctl6
+ dacp_0/bootstrapped_sw_p_0/enb dacp_0/dac_out dacp_0/ctl3 dacp_0/bootstrapped_sw_p_0/vg
+ dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n9 dacp_0/ctl5 dacp_0/carray_p_0/n7 vdd dacp_0/bootstrapped_sw_p_0/vbsh
+ vdd dacp_0/bootstrapped_sw_p_0/vbsl dacp
Xdacn_0 vinn dacn_0/ctl1 dacn_0/ctl2 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5 dacn_0/ctl6
+ dacn_0/ctl7 dacn_0/ctl8 dacn_0/ctl9 dacn_0/ctl10 dacn_0/bootstrapped_sw_n_0/vg dacn_0/bootstrapped_sw_n_0/enb
+ dacn_0/carray_n_0/n9 dacp_0/sample dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n0 vdd
+ dacn_0/carray_n_0/n8 dacn_0/bootstrapped_sw_n_0/vbsh dacn_0/dac_out vdd vdd dacn_0/bootstrapped_sw_n_0/vbsl
+ dacn_0/carray_n_0/ndum dacn
Xcomparator_0 sarlogic_0/trim[1] sarlogic_0/trim[0] sarlogic_0/trim[4] sarlogic_0/trimb[4]
+ sarlogic_0/trimb[1] sarlogic_0/trimb[0] sarlogic_0/trimb[2] sarlogic_0/trimb[3]
+ dacp_0/dac_out dacn_0/dac_out comparator_0/in comparator_0/ip comparator_0/diff
+ comparator_0/trim_right_0/n3 comparator_0/trim_left_0/n4 comparator_0/trim_left_0/n2
+ comparator_0/trim_left_0/n3 buffer_0/buf_out sarlogic_0/trim[3] latch_0/S sarlogic_0/trim[2]
+ vdd latch_0/R comparator_0/trim_right_0/n4 comparator_0/trim_right_0/n2 vdd comparator
Xmim_cap_boss_0 vss vdd vdd mim_cap_boss
Xsarlogic_0 dacn_0/ctl10 dacn_0/ctl1 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5 dacn_0/ctl6
+ dacn_0/ctl8 dacp_0/ctl10 dacp_0/ctl1 dacp_0/ctl2 dacp_0/ctl3 dacp_0/ctl4 dacp_0/ctl5
+ dacp_0/ctl6 dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9 clk sarlogic_0/clkc latch_0/Q en
+ result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7]
+ result[8] result[9] rstn dacp_0/sample sarlogic_0/trim[0] sarlogic_0/trim[1] sarlogic_0/trim[2]
+ sarlogic_0/trim[3] sarlogic_0/trim[4] sarlogic_0/trimb[0] sarlogic_0/trimb[1] sarlogic_0/trimb[2]
+ sarlogic_0/trimb[3] sarlogic_0/trimb[4] valid sarlogic_0/net10 sarlogic_0/output13/a_224_472#
+ sarlogic_0/output23/a_224_472# sarlogic_0/net59 sarlogic_0/net16 sarlogic_0/net27
+ sarlogic_0/output25/a_224_472# sarlogic_0/cal_itt\[1\] sarlogic_0/fanout65/a_36_113#
+ dacn_0/ctl2 dacn_0/ctl7 sarlogic_0/net15 dacn_0/ctl9 sarlogic_0/output10/a_224_472#
+ sarlogic_0/net26 sarlogic_0/net24 sarlogic_0/output11/a_224_472# sarlogic_0/output21/a_224_472#
+ sarlogic_0/net14 sarlogic_0/output12/a_224_472# sarlogic_0/output22/a_224_472# cal
+ sarlogic_0/net62 sarlogic_0/net20 vdd vdd sarlogic
Xmim_cap_boss_1 vss vdd vdd mim_cap_boss
C0 dacp_0/dac_out vdd 1.335938f
C1 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n9 87.10268f
C2 comparator_0/trim_left_0/n4 comparator_0/trim_left_0/n2 0.128631f
C3 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n1 0.134826f
C4 dacp_0/ctl6 dacp_0/ctl5 3.114209f
C5 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n6 14.716789f
C6 dacp_0/ctl6 vdd 1.604297f
C7 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n2 0.213096f
C8 vdd rstn 3.591095f
C9 sarlogic_0/trimb[2] vdd 0.775533f
C10 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n4 2.84323f
C11 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n5 3.36878f
C12 dacp_0/ctl8 dacp_0/ctl7 2.592389f
C13 dacn_0/dac_out dacn_0/carray_n_0/n0 1.702719f
C14 dacn_0/carray_n_0/n6 dacn_0/dac_out 0.105055p
C15 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n6 0.614078f
C16 en vdd 3.37982f
C17 dacn_0/bootstrapped_sw_n_0/vbsh dacp_0/bootstrapped_sw_p_0/vbsh 0.302212f
C18 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n0 0.097254f
C19 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n8 11.2161f
C20 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n1 0.134705f
C21 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n0 0.06073f
C22 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n6 34.326103f
C23 dacp_0/bootstrapped_sw_p_0/vbsl dacn_0/bootstrapped_sw_n_0/vbsl 0.256194f
C24 comparator_0/in vdd 3.523928f
C25 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/ndum 0.06073f
C26 dacp_0/bootstrapped_sw_p_0/vbsh vdd 0.507196f
C27 dacn_0/ctl8 dacn_0/ctl9 2.33149f
C28 dacn_0/carray_n_0/n1 dacn_0/carray_n_0/n5 0.134705f
C29 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n4 3.740573f
C30 result[8] result[9] 3.472163f
C31 valid cal 3.472163f
C32 dacp_0/carray_p_0/n1 dacp_0/carray_p_0/ndum 8.161697f
C33 vss clk 8.402781f
C34 result[0] result[1] 3.472163f
C35 vinn vss 13.325f
C36 sarlogic_0/output10/a_224_472# vdd 0.006335f
C37 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n6 0.025424f
C38 comparator_0/trim_left_0/n4 vdd 0.117372f
C39 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n5 7.399346f
C40 dacp_0/sample clk 0.171212f
C41 result[4] vss 8.402781f
C42 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n3 0.336612f
C43 dacn_0/carray_n_0/n3 dacn_0/carray_n_0/n0 0.051666f
C44 comparator_0/ip vdd 3.523929f
C45 latch_0/Q vdd 0.493384f
C46 vinp vdd 4.8626f
C47 result[4] dacp_0/sample 0.160929f
C48 valid vss 8.4233f
C49 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n2 0.207999f
C50 dacp_0/dac_out dacp_0/bootstrapped_sw_p_0/vbsl -0.018699f
C51 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n5 5.60732f
C52 dacn_0/ctl9 vdd 1.645072f
C53 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n4 3.740573f
C54 dacp_0/carray_p_0/n7 vdd 0.040786f
C55 sarlogic_0/trimb[3] vdd 1.519255f
C56 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n5 28.589401f
C57 comparator_0/trim_right_0/n4 comparator_0/trim_right_0/n2 0.128631f
C58 dacp_0/sample valid 0.161748f
C59 latch_0/R latch_0/Q 0.001492f
C60 dacp_0/carray_p_0/n2 dacp_0/carray_p_0/ndum 0.041162f
C61 sarlogic_0/output11/a_224_472# vdd 0.006847f
C62 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/ndum 0.097254f
C63 cal vss 8.402781f
C64 dacp_0/ctl8 vdd 1.685297f
C65 vss m5_121784_n195240# 0.79769p
C66 sarlogic_0/output13/a_224_472# vdd 0.006752f
C67 dacn_0/carray_n_0/n2 dacn_0/dac_out 6.640605f
C68 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/ndum 0.025424f
C69 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n8 0.770114f
C70 latch_0/Qn vdd 0.148748f
C71 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n2 0.485242f
C72 dacp_0/bootstrapped_sw_p_0/vbsh dacn_0/bootstrapped_sw_n_0/vbsl 0.015167f
C73 sarlogic_0/trim[2] sarlogic_0/trim[0] 3.076354f
C74 dacn_0/ctl2 vdd 2.454649f
C75 dacp_0/sample cal 0.161292f
C76 dacp_0/dac_out dacp_0/carray_p_0/n0 1.702719f
C77 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n0 0.025424f
C78 dacn_0/ctl1 vdd 2.70229f
C79 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n0 0.051666f
C80 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n2 0.041162f
C81 dacn_0/carray_n_0/n4 dacn_0/dac_out 26.32268f
C82 dacp_0/ctl5 dacp_0/ctl4 3.375109f
C83 sarlogic_0/net10 vdd 0.001258f
C84 dacn_0/ctl10 dacn_0/ctl9 2.076967f
C85 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n8 2.84323f
C86 sarlogic_0/trim[1] vdd 0.763954f
C87 dacp_0/ctl4 vdd 1.829149f
C88 sarlogic_0/output23/a_224_472# vdd 0.005853f
C89 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n7 1.70387f
C90 dacp_0/ctl3 dacp_0/ctl2 3.896919f
C91 sarlogic_0/trim[0] vdd 0.764556f
C92 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n3 22.8406f
C93 dacn_0/ctl2 dacn_0/ctl3 3.89692f
C94 comparator_0/trim_left_0/n3 vdd 0.230601f
C95 dacp_0/sample sarlogic_0/cal_itt\[1\] 0.004307f
C96 dacp_0/dac_out dacp_0/carray_p_0/n3 13.201303f
C97 sarlogic_0/net16 vdd 0.001182f
C98 vinp dacp_0/bootstrapped_sw_p_0/vbsl 0.007238f
C99 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n5 7.399346f
C100 dacp_0/carray_p_0/n8 vdd 0.075671f
C101 dacn_0/dac_out dacn_0/carray_n_0/n5 52.565514f
C102 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n5 5.60732f
C103 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n5 3.36878f
C104 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/ndum 0.025424f
C105 dacp_0/dac_out dacp_0/bootstrapped_sw_p_0/vbsh -0.004073f
C106 sarlogic_0/trim[4] vdd 1.198372f
C107 clk vdd 3.532875f
C108 result[4] result[5] 3.472163f
C109 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n5 27.491999f
C110 sarlogic_0/net20 vdd 0.004671f
C111 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/ndum 0.127951f
C112 vinn vdd 4.8626f
C113 comparator_0/trim_right_0/n2 vdd 0.0311f
C114 dacp_0/ctl9 vdd 1.724922f
C115 sarlogic_0/trimb[4] vdd 1.196384f
C116 comparator_0/ip comparator_0/trim_right_0/n3 6.42492f
C117 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n3 25.8929f
C118 comparator_0/ip comparator_0/trim_right_0/n0 1.60623f
C119 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/ndum 0.025424f
C120 dacn_0/bootstrapped_sw_n_0/enb vdd 0.019924f
C121 comparator_0/trim_right_0/n4 comparator_0/trim_right_0/n1 0.032158f
C122 result[4] vdd 3.379693f
C123 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n5 0.025424f
C124 vss m5_n161680_n110000# 0.79769p
C125 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n2 0.207877f
C126 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n0 0.099202f
C127 result[2] vss 8.402781f
C128 latch_0/S latch_0/Qn 0.014677f
C129 buffer_0/buf_out vdd 0.967639f
C130 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n0 0.06073f
C131 valid vdd 3.414013f
C132 dacn_0/carray_n_0/n3 dacn_0/carray_n_0/n5 0.346757f
C133 sarlogic_0/trim[2] sarlogic_0/trim[3] 2.938384f
C134 dacp_0/ctl3 vdd 2.055974f
C135 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/n1 8.469266f
C136 result[2] dacp_0/sample 0.160984f
C137 sarlogic_0/trimb[3] dacp_0/ctl10 0.087957f
C138 comparator_0/trim_left_0/n4 comparator_0/in 12.849839f
C139 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n1 0.342393f
C140 dacp_0/sample dacp_0/carray_p_0/ndum 0.002948f
C141 sarlogic_0/trimb[0] vdd 0.764556f
C142 cal vdd 3.379693f
C143 sarlogic_0/trimb[1] sarlogic_0/trimb[4] 2.912714f
C144 m5_121784_n195240# vdd 0.107014p
C145 buffer_0/buf_out latch_0/R 0.078509f
C146 dacp_0/dac_out dacp_0/carray_p_0/n7 0.210031p
C147 sarlogic_0/output22/a_224_472# vdd 0.006461f
C148 dacp_0/carray_p_0/n9 vdd 0.09396f
C149 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n0 0.040502f
C150 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n6 0.614078f
C151 dacp_0/dac_out dacp_0/carray_p_0/n1 3.365905f
C152 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n3 0.891504f
C153 sarlogic_0/output21/a_224_472# vdd 0.00611f
C154 sarlogic_0/trim[3] vdd 1.519256f
C155 sarlogic_0/trimb[2] sarlogic_0/trimb[3] 2.930414f
C156 result[5] vss 8.402781f
C157 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n1 0.137399f
C158 vinn dacn_0/bootstrapped_sw_n_0/vbsl 0.007238f
C159 sarlogic_0/clkc buffer_0/inv2_0/inv_in 0.002377f
C160 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/ndum 0.025424f
C161 dacn_0/carray_n_0/n5 dacn_0/carray_n_0/n0 0.025424f
C162 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n5 28.589401f
C163 dacp_0/sample result[5] 0.160929f
C164 sarlogic_0/trimb[1] sarlogic_0/trimb[0] 2.974034f
C165 dacp_0/carray_p_0/n0 dacp_0/carray_p_0/n2 0.099202f
C166 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n0 0.097254f
C167 dacp_0/sample vdd 18.621128f
C168 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n0 0.025424f
C169 result[4] result[3] 3.472163f
C170 sarlogic_0/fanout65/a_36_113# dacp_0/sample 0.001365f
C171 dacn_0/ctl4 dacn_0/ctl5 3.37511f
C172 result[7] vss 8.402781f
C173 dacn_0/ctl5 vdd 1.681347f
C174 dacn_0/bootstrapped_sw_n_0/vg vdd 0.015751f
C175 sarlogic_0/net15 vdd 0.00664f
C176 latch_0/tutyuu1 vdd 0.022865f
C177 dacp_0/dac_out dacp_0/carray_p_0/n2 6.640605f
C178 sarlogic_0/clkc vdd 0.309923f
C179 dacn_0/ctl10 sarlogic_0/trim[3] 0.097876f
C180 vdd sarlogic_0/net14 0.005269f
C181 dacp_0/carray_p_0/n8 dacp_0/dac_out 0.420151p
C182 dacp_0/sample result[7] 0.161003f
C183 comparator_0/trim_right_0/n4 vdd 0.117372f
C184 dacp_0/dac_out dacp_0/carray_p_0/n6 0.105055p
C185 dacp_0/ctl9 dacp_0/ctl10 2.076966f
C186 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n2 22.8406f
C187 dacp_0/ctl1 dacp_0/ctl2 4.157828f
C188 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n3 1.46111f
C189 dacp_0/ctl7 vdd 1.581332f
C190 comparator_0/trim_left_0/n3 comparator_0/in 6.42492f
C191 dacp_0/sample sarlogic_0/net62 0.160765f
C192 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n3 0.336612f
C193 dacn_0/carray_n_0/n9 vdd 0.09396f
C194 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n2 0.213096f
C195 sarlogic_0/net26 vdd 0.001136f
C196 m5_n161680_n110000# vdd 0.107014p
C197 dacp_0/ctl2 vdd 2.536638f
C198 clk rstn 3.472163f
C199 dacn_0/dac_out dacn_0/carray_n_0/n1 3.365905f
C200 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n1 0.278221f
C201 result[2] vdd 3.379693f
C202 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n1 0.205173f
C203 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n1 0.205173f
C204 en clk 3.472163f
C205 comparator_0/in comparator_0/trim_left_0/n0 1.60623f
C206 dacn_0/ctl8 dacn_0/ctl7 2.59239f
C207 result[0] vss 8.4233f
C208 dacn_0/ctl8 vdd 1.526202f
C209 comparator_0/trim_left_0/n3 comparator_0/trim_left_0/n4 0.241184f
C210 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n5 0.207999f
C211 dacp_0/sample dacn_0/carray_n_0/ndum 0.002948f
C212 comparator_0/trim_left_0/n2 vdd 0.0311f
C213 result[9] vss 8.4233f
C214 dacn_0/carray_n_0/n9 dacn_0/dac_out 0.846152p
C215 dacp_0/sample sarlogic_0/net59 0.022016f
C216 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n0 0.184985f
C217 buffer_0/inv2_0/inv_in vdd 0.165047f
C218 dacp_0/sample result[0] 0.161748f
C219 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n8 87.10268f
C220 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n7 29.516087f
C221 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n1 8.161697f
C222 sarlogic_0/trim[2] vdd 0.776953f
C223 result[8] vss 8.402781f
C224 sarlogic_0/net24 vdd 0.004775f
C225 vss result[3] 8.402781f
C226 comparator_0/trim_left_0/n4 comparator_0/trim_left_0/n0 0.032158f
C227 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n0 0.040502f
C228 dacp_0/sample result[9] 0.161326f
C229 dacn_0/carray_n_0/n3 dacn_0/carray_n_0/n1 0.137399f
C230 buffer_0/buf_out comparator_0/in 0.052543f
C231 comparator_0/trim_left_0/n1 comparator_0/in 1.60623f
C232 dacn_0/ctl2 dacn_0/ctl1 4.157831f
C233 dacp_0/sample result[8] 0.161003f
C234 dacp_0/carray_p_0/n9 dacp_0/dac_out 0.846152p
C235 dacp_0/sample result[3] 0.160929f
C236 sarlogic_0/trimb[0] sarlogic_0/trimb[2] 3.076354f
C237 result[5] vdd 3.379693f
C238 dacn_0/carray_n_0/n4 dacn_0/carray_n_0/n5 27.491999f
C239 dacp_0/ctl1 vdd 2.707573f
C240 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/ndum 0.127951f
C241 result[1] vss 8.402781f
C242 result[6] vss 8.402781f
C243 dacn_0/ctl5 dacn_0/ctl6 3.114201f
C244 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n3 1.911224f
C245 comparator_0/ip comparator_0/trim_right_0/n2 3.21246f
C246 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n2 0.485242f
C247 dacn_0/bootstrapped_sw_n_0/vbsh vdd 0.507197f
C248 dacp_0/carray_p_0/n4 dacp_0/dac_out 26.32268f
C249 cal en 3.472141f
C250 latch_0/S latch_0/tutyuu1 0.005953f
C251 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n7 50.178104f
C252 dacp_0/ctl5 vdd 1.681347f
C253 dacn_0/ctl7 vdd 1.585582f
C254 dacn_0/ctl4 vdd 1.827967f
C255 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n3 1.911224f
C256 comparator_0/trim_right_0/n1 comparator_0/trim_right_0/n0 0.032158f
C257 dacp_0/carray_p_0/n7 dacp_0/carray_p_0/n6 34.326103f
C258 dacp_0/sample result[1] 0.160984f
C259 result[6] dacp_0/sample 0.161003f
C260 comparator_0/trim_left_0/n1 comparator_0/trim_left_0/n4 0.032158f
C261 dacp_0/carray_p_0/n1 dacp_0/carray_p_0/n2 16.597801f
C262 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n3 25.8929f
C263 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n1 0.278221f
C264 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n1 0.134562f
C265 result[7] vdd 3.37982f
C266 sarlogic_0/output12/a_224_472# vdd 0.006182f
C267 latch_0/R vdd 1.621428f
C268 vss rstn 8.4233f
C269 dacn_0/bootstrapped_sw_n_0/vbsh dacn_0/dac_out -0.004073f
C270 dacp_0/ctl9 dacp_0/ctl8 2.331489f
C271 comparator_0/trim_right_0/n4 comparator_0/trim_right_0/n3 0.241184f
C272 result[2] result[3] 3.472163f
C273 dacn_0/carray_n_0/n6 dacn_0/carray_n_0/n1 0.134562f
C274 dacn_0/carray_n_0/n1 dacn_0/carray_n_0/n0 8.469266f
C275 dacn_0/dac_out vdd 1.335938f
C276 comparator_0/trim_right_0/n4 comparator_0/trim_right_0/n0 0.032158f
C277 dacn_0/ctl4 dacn_0/ctl3 3.636021f
C278 vss en 8.402781f
C279 dacn_0/ctl3 vdd 2.054162f
C280 dacn_0/carray_n_0/n8 vdd 0.075671f
C281 sarlogic_0/trim[0] sarlogic_0/trim[1] 2.966054f
C282 dacn_0/carray_n_0/n7 vdd 0.040786f
C283 dacp_0/sample rstn 0.161326f
C284 dacp_0/carray_p_0/n5 dacp_0/carray_p_0/n0 0.025424f
C285 sarlogic_0/trimb[1] vdd 0.765374f
C286 dacp_0/sample en 0.18575f
C287 result[2] result[1] 3.472163f
C288 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n0 0.184985f
C289 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n6 14.716789f
C290 dacn_0/ctl10 vdd 1.583664f
C291 sarlogic_0/trim[4] sarlogic_0/trim[1] 2.904734f
C292 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n2 0.770114f
C293 dacp_0/dac_out dacp_0/carray_p_0/n5 52.565514f
C294 dacn_0/dac_out dacn_0/carray_n_0/n8 0.420151p
C295 dacn_0/carray_n_0/n7 dacn_0/dac_out 0.210031p
C296 dacp_0/ctl7 dacp_0/ctl6 2.853299f
C297 dacp_0/carray_p_0/n6 dacp_0/carray_p_0/n2 0.207877f
C298 result[0] vdd 3.414013f
C299 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n8 50.178104f
C300 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n7 29.516087f
C301 dacp_0/carray_p_0/n8 dacp_0/carray_p_0/n6 11.2161f
C302 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/n5 0.346757f
C303 dacp_0/dac_out dacp_0/carray_p_0/ndum 1.640173f
C304 dacn_0/bootstrapped_sw_n_0/vbsh dacp_0/bootstrapped_sw_p_0/vbsl 0.015167f
C305 dacn_0/bootstrapped_sw_n_0/vbsl vdd 1.612052f
C306 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n1 0.342393f
C307 vinp vss 13.325f
C308 result[9] vdd 3.595587f
C309 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n7 1.70387f
C310 dacp_0/bootstrapped_sw_p_0/vbsl vdd 1.612052f
C311 comparator_0/trim_right_0/n1 comparator_0/ip 1.60623f
C312 dacp_0/carray_p_0/n3 dacp_0/carray_p_0/ndum 0.025424f
C313 latch_0/tutyuu2 vdd 0.087409f
C314 result[8] vdd 3.838088f
C315 dacn_0/carray_n_0/ndum dacn_0/dac_out 1.640173f
C316 vdd result[3] 3.379693f
C317 latch_0/S vdd 1.883988f
C318 dacp_0/carray_p_0/n4 dacp_0/carray_p_0/n1 0.134826f
C319 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n8 0.097254f
C320 dacn_0/ctl7 dacn_0/ctl6 2.853301f
C321 dacn_0/ctl6 vdd 1.606092f
C322 result[6] result[5] 3.472163f
C323 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/ndum 0.06073f
C324 dacp_0/ctl4 dacp_0/ctl3 3.636019f
C325 dacn_0/dac_out dacn_0/carray_n_0/n3 13.201303f
C326 dacn_0/carray_n_0/n8 dacn_0/carray_n_0/n3 1.46111f
C327 result[7] result[8] 3.472163f
C328 dacn_0/carray_n_0/n7 dacn_0/carray_n_0/n3 0.891504f
C329 dacn_0/dac_out dacn_0/bootstrapped_sw_n_0/vbsl -0.018699f
C330 dacn_0/carray_n_0/n2 dacn_0/carray_n_0/n1 16.597801f
C331 latch_0/R latch_0/tutyuu2 0.005568f
C332 comparator_0/trim_right_0/n3 vdd 0.2306f
C333 result[1] vdd 3.379693f
C334 result[6] vdd 3.379693f
C335 latch_0/S latch_0/R 0.183801f
C336 comparator_0/trim_right_0/n4 comparator_0/ip 12.849839f
C337 comparator_0/trim_left_0/n1 comparator_0/trim_left_0/n0 0.032158f
C338 comparator_0/in comparator_0/trim_left_0/n2 3.21246f
C339 dacp_0/bootstrapped_sw_p_0/enb vdd 0.019924f
C340 sarlogic_0/output25/a_224_472# vdd 0.005027f
C341 dacp_0/ctl10 vdd 1.583664f
C342 result[6] result[7] 3.472163f
C343 dacp_0/sample sarlogic_0/net27 0.004307f
C344 dacp_0/bootstrapped_sw_p_0/vg vdd 0.015751f
C345 dacn_0/carray_n_0/ndum dacn_0/carray_n_0/n3 0.025424f
C346 dacn_0/carray_n_0/n9 dacn_0/carray_n_0/n2 0.996568f
C347 dacp_0/carray_p_0/n9 dacp_0/carray_p_0/n2 0.996568f
C348 m5_121784_n195240# 0 0.191258p $ **FLOATING
C349 m5_n161680_n110000# 0 0.191258p $ **FLOATING
C350 sarlogic_0/_034_ 0 0.304805f
C351 sarlogic_0/_160_ 0 1.542665f
C352 sarlogic_0/_166_ 0 0.299751f
C353 sarlogic_0/output41/a_224_472# 0 2.38465f
C354 sarlogic_0/net6 0 1.112469f
C355 sarlogic_0/output6/a_224_472# 0 2.38465f
C356 sarlogic_0/FILLER_0_12_196/a_36_472# 0 0.417394f
C357 sarlogic_0/FILLER_0_12_196/a_124_375# 0 0.246306f
C358 result[3] 0 16.841412f
C359 sarlogic_0/net30 0 1.81422f
C360 sarlogic_0/output30/a_224_472# 0 2.38465f
C361 sarlogic_0/_047_ 0 0.374694f
C362 sarlogic_0/_201_/a_67_603# 0 0.345683f
C363 sarlogic_0/_416_/a_2560_156# 0 0.016968f
C364 sarlogic_0/_416_/a_2665_112# 0 0.62251f
C365 sarlogic_0/_416_/a_2248_156# 0 0.371662f
C366 sarlogic_0/_416_/a_1204_472# 0 0.012971f
C367 sarlogic_0/_416_/a_1000_472# 0 0.291735f
C368 sarlogic_0/_416_/a_796_472# 0 0.023206f
C369 sarlogic_0/_416_/a_1308_423# 0 0.279043f
C370 sarlogic_0/_416_/a_448_472# 0 0.684413f
C371 sarlogic_0/_416_/a_36_151# 0 1.43589f
C372 sarlogic_0/FILLER_0_13_290/a_36_472# 0 0.417394f
C373 sarlogic_0/FILLER_0_13_290/a_124_375# 0 0.246306f
C374 sarlogic_0/_278_/a_36_160# 0 0.696445f
C375 sarlogic_0/_145_ 0 0.546455f
C376 sarlogic_0/FILLER_0_13_72/a_484_472# 0 0.345058f
C377 sarlogic_0/FILLER_0_13_72/a_36_472# 0 0.404746f
C378 sarlogic_0/FILLER_0_13_72/a_572_375# 0 0.232991f
C379 sarlogic_0/FILLER_0_13_72/a_124_375# 0 0.185089f
C380 sarlogic_0/FILLER_0_14_235/a_484_472# 0 0.345058f
C381 sarlogic_0/FILLER_0_14_235/a_36_472# 0 0.404746f
C382 sarlogic_0/FILLER_0_14_235/a_572_375# 0 0.232991f
C383 sarlogic_0/FILLER_0_14_235/a_124_375# 0 0.185089f
C384 sarlogic_0/_156_ 0 0.593796f
C385 sarlogic_0/_107_ 0 0.391583f
C386 sarlogic_0/_295_/a_36_472# 0 0.031137f
C387 sarlogic_0/_022_ 0 0.387773f
C388 sarlogic_0/_433_/a_2560_156# 0 0.016968f
C389 sarlogic_0/_433_/a_2665_112# 0 0.62251f
C390 sarlogic_0/_433_/a_2248_156# 0 0.371662f
C391 sarlogic_0/_433_/a_1204_472# 0 0.012971f
C392 sarlogic_0/_433_/a_1000_472# 0 0.291735f
C393 sarlogic_0/_433_/a_796_472# 0 0.023206f
C394 sarlogic_0/_433_/a_1308_423# 0 0.279043f
C395 sarlogic_0/_433_/a_448_472# 0 0.684413f
C396 sarlogic_0/_433_/a_36_151# 0 1.43589f
C397 sarlogic_0/FILLER_0_5_148/a_484_472# 0 0.345058f
C398 sarlogic_0/FILLER_0_5_148/a_36_472# 0 0.404746f
C399 sarlogic_0/FILLER_0_5_148/a_572_375# 0 0.232991f
C400 sarlogic_0/FILLER_0_5_148/a_124_375# 0 0.185089f
C401 sarlogic_0/_167_ 0 0.285904f
C402 sarlogic_0/_381_/a_36_472# 0 0.031137f
C403 sarlogic_0/net40 0 1.845219f
C404 sarlogic_0/output40/a_224_472# 0 2.38465f
C405 sarlogic_0/cal_count\[0\] 0 0.893784f
C406 sarlogic_0/_039_ 0 0.412301f
C407 sarlogic_0/_450_/a_2449_156# 0 0.049992f
C408 sarlogic_0/_450_/a_2225_156# 0 0.434082f
C409 sarlogic_0/_450_/a_3129_107# 0 0.58406f
C410 sarlogic_0/_450_/a_836_156# 0 0.019766f
C411 sarlogic_0/_450_/a_1040_527# 0 0.302082f
C412 sarlogic_0/_450_/a_1353_112# 0 0.286513f
C413 sarlogic_0/_450_/a_448_472# 0 1.21246f
C414 sarlogic_0/_450_/a_36_151# 0 1.31409f
C415 rstn 0 22.56473f
C416 sarlogic_0/FILLER_0_8_156/a_484_472# 0 0.345058f
C417 sarlogic_0/FILLER_0_8_156/a_36_472# 0 0.404746f
C418 sarlogic_0/FILLER_0_8_156/a_572_375# 0 0.232991f
C419 sarlogic_0/FILLER_0_8_156/a_124_375# 0 0.185089f
C420 sarlogic_0/FILLER_0_6_37/a_36_472# 0 0.417394f
C421 sarlogic_0/FILLER_0_6_37/a_124_375# 0 0.246306f
C422 sarlogic_0/FILLER_0_21_60/a_484_472# 0 0.345058f
C423 sarlogic_0/FILLER_0_21_60/a_36_472# 0 0.404746f
C424 sarlogic_0/FILLER_0_21_60/a_572_375# 0 0.232991f
C425 sarlogic_0/FILLER_0_21_60/a_124_375# 0 0.185089f
C426 sarlogic_0/FILLER_0_22_107/a_484_472# 0 0.345058f
C427 sarlogic_0/FILLER_0_22_107/a_36_472# 0 0.404746f
C428 sarlogic_0/FILLER_0_22_107/a_572_375# 0 0.232991f
C429 sarlogic_0/FILLER_0_22_107/a_124_375# 0 0.185089f
C430 sarlogic_0/FILLER_0_16_115/a_36_472# 0 0.417394f
C431 sarlogic_0/FILLER_0_16_115/a_124_375# 0 0.246306f
C432 sarlogic_0/FILLER_0_19_134/a_36_472# 0 0.417394f
C433 sarlogic_0/FILLER_0_19_134/a_124_375# 0 0.246306f
C434 sarlogic_0/FILLER_0_3_212/a_36_472# 0 0.417394f
C435 sarlogic_0/FILLER_0_3_212/a_124_375# 0 0.246306f
C436 sarlogic_0/FILLER_0_10_94/a_484_472# 0 0.345058f
C437 sarlogic_0/FILLER_0_10_94/a_36_472# 0 0.404746f
C438 sarlogic_0/FILLER_0_10_94/a_572_375# 0 0.232991f
C439 sarlogic_0/FILLER_0_10_94/a_124_375# 0 0.185089f
C440 sarlogic_0/FILLER_0_4_91/a_484_472# 0 0.345058f
C441 sarlogic_0/FILLER_0_4_91/a_36_472# 0 0.404746f
C442 sarlogic_0/FILLER_0_4_91/a_572_375# 0 0.232991f
C443 sarlogic_0/FILLER_0_4_91/a_124_375# 0 0.185089f
C444 sarlogic_0/net14 0 1.508711f
C445 sarlogic_0/_202_/a_36_160# 0 0.696445f
C446 sarlogic_0/FILLER_0_6_231/a_484_472# 0 0.345058f
C447 sarlogic_0/FILLER_0_6_231/a_36_472# 0 0.404746f
C448 sarlogic_0/FILLER_0_6_231/a_572_375# 0 0.232991f
C449 sarlogic_0/FILLER_0_6_231/a_124_375# 0 0.185089f
C450 vdd 0 16.260454p
C451 sarlogic_0/_006_ 0 0.41456f
C452 sarlogic_0/_417_/a_2560_156# 0 0.016968f
C453 sarlogic_0/_417_/a_2665_112# 0 0.62251f
C454 sarlogic_0/_417_/a_2248_156# 0 0.371662f
C455 sarlogic_0/_417_/a_1204_472# 0 0.012971f
C456 sarlogic_0/_417_/a_1000_472# 0 0.291735f
C457 sarlogic_0/_417_/a_796_472# 0 0.023206f
C458 sarlogic_0/_417_/a_1308_423# 0 0.279043f
C459 sarlogic_0/_417_/a_448_472# 0 0.684413f
C460 sarlogic_0/_417_/a_36_151# 0 1.43589f
C461 sarlogic_0/_146_ 0 0.35443f
C462 sarlogic_0/mask\[6\] 0 1.246962f
C463 sarlogic_0/_348_/a_49_472# 0 0.054843f
C464 sarlogic_0/_365_/a_36_68# 0 0.150048f
C465 sarlogic_0/_023_ 0 0.345812f
C466 sarlogic_0/_434_/a_2560_156# 0 0.016968f
C467 sarlogic_0/_434_/a_2665_112# 0 0.62251f
C468 sarlogic_0/_434_/a_2248_156# 0 0.371662f
C469 sarlogic_0/_434_/a_1204_472# 0 0.012971f
C470 sarlogic_0/_434_/a_1000_472# 0 0.291735f
C471 sarlogic_0/_434_/a_796_472# 0 0.023206f
C472 sarlogic_0/_434_/a_1308_423# 0 0.279043f
C473 sarlogic_0/_434_/a_448_472# 0 0.684413f
C474 sarlogic_0/_434_/a_36_151# 0 1.43589f
C475 sarlogic_0/FILLER_0_5_136/a_36_472# 0 0.417394f
C476 sarlogic_0/FILLER_0_5_136/a_124_375# 0 0.246306f
C477 sarlogic_0/FILLER_0_18_209/a_484_472# 0 0.345058f
C478 sarlogic_0/FILLER_0_18_209/a_36_472# 0 0.404746f
C479 sarlogic_0/FILLER_0_18_209/a_572_375# 0 0.232991f
C480 sarlogic_0/FILLER_0_18_209/a_124_375# 0 0.185089f
C481 sarlogic_0/FILLER_0_12_28/a_36_472# 0 0.417394f
C482 sarlogic_0/FILLER_0_12_28/a_124_375# 0 0.246306f
C483 sarlogic_0/_040_ 0 0.355703f
C484 sarlogic_0/_451_/a_2449_156# 0 0.049992f
C485 sarlogic_0/_451_/a_2225_156# 0 0.434082f
C486 sarlogic_0/_451_/a_3129_107# 0 0.58406f
C487 sarlogic_0/_451_/a_836_156# 0 0.019766f
C488 sarlogic_0/_451_/a_1040_527# 0 0.302082f
C489 sarlogic_0/_451_/a_1353_112# 0 0.286513f
C490 sarlogic_0/_451_/a_448_472# 0 1.21246f
C491 sarlogic_0/_451_/a_36_151# 0 1.31409f
C492 sarlogic_0/FILLER_0_6_47/a_3172_472# 0 0.345058f
C493 sarlogic_0/FILLER_0_6_47/a_2724_472# 0 0.33241f
C494 sarlogic_0/FILLER_0_6_47/a_2276_472# 0 0.33241f
C495 sarlogic_0/FILLER_0_6_47/a_1828_472# 0 0.33241f
C496 sarlogic_0/FILLER_0_6_47/a_1380_472# 0 0.33241f
C497 sarlogic_0/FILLER_0_6_47/a_932_472# 0 0.33241f
C498 sarlogic_0/FILLER_0_6_47/a_484_472# 0 0.33241f
C499 sarlogic_0/FILLER_0_6_47/a_36_472# 0 0.404746f
C500 sarlogic_0/FILLER_0_6_47/a_3260_375# 0 0.233093f
C501 sarlogic_0/FILLER_0_6_47/a_2812_375# 0 0.17167f
C502 sarlogic_0/FILLER_0_6_47/a_2364_375# 0 0.17167f
C503 sarlogic_0/FILLER_0_6_47/a_1916_375# 0 0.17167f
C504 sarlogic_0/FILLER_0_6_47/a_1468_375# 0 0.17167f
C505 sarlogic_0/FILLER_0_6_47/a_1020_375# 0 0.17167f
C506 sarlogic_0/FILLER_0_6_47/a_572_375# 0 0.17167f
C507 sarlogic_0/FILLER_0_6_47/a_124_375# 0 0.185915f
C508 sarlogic_0/FILLER_0_21_150/a_36_472# 0 0.417394f
C509 sarlogic_0/FILLER_0_21_150/a_124_375# 0 0.246306f
C510 sarlogic_0/FILLER_0_15_180/a_484_472# 0 0.345058f
C511 sarlogic_0/FILLER_0_15_180/a_36_472# 0 0.404746f
C512 sarlogic_0/FILLER_0_15_180/a_572_375# 0 0.232991f
C513 sarlogic_0/FILLER_0_15_180/a_124_375# 0 0.185089f
C514 sarlogic_0/FILLER_0_22_128/a_3172_472# 0 0.345058f
C515 sarlogic_0/FILLER_0_22_128/a_2724_472# 0 0.33241f
C516 sarlogic_0/FILLER_0_22_128/a_2276_472# 0 0.33241f
C517 sarlogic_0/FILLER_0_22_128/a_1828_472# 0 0.33241f
C518 sarlogic_0/FILLER_0_22_128/a_1380_472# 0 0.33241f
C519 sarlogic_0/FILLER_0_22_128/a_932_472# 0 0.33241f
C520 sarlogic_0/FILLER_0_22_128/a_484_472# 0 0.33241f
C521 sarlogic_0/FILLER_0_22_128/a_36_472# 0 0.404746f
C522 sarlogic_0/FILLER_0_22_128/a_3260_375# 0 0.233093f
C523 sarlogic_0/FILLER_0_22_128/a_2812_375# 0 0.17167f
C524 sarlogic_0/FILLER_0_22_128/a_2364_375# 0 0.17167f
C525 sarlogic_0/FILLER_0_22_128/a_1916_375# 0 0.17167f
C526 sarlogic_0/FILLER_0_22_128/a_1468_375# 0 0.17167f
C527 sarlogic_0/FILLER_0_22_128/a_1020_375# 0 0.17167f
C528 sarlogic_0/FILLER_0_22_128/a_572_375# 0 0.17167f
C529 sarlogic_0/FILLER_0_22_128/a_124_375# 0 0.185915f
C530 sarlogic_0/FILLER_0_19_111/a_484_472# 0 0.345058f
C531 sarlogic_0/FILLER_0_19_111/a_36_472# 0 0.404746f
C532 sarlogic_0/FILLER_0_19_111/a_572_375# 0 0.232991f
C533 sarlogic_0/FILLER_0_19_111/a_124_375# 0 0.185089f
C534 sarlogic_0/FILLER_0_19_155/a_484_472# 0 0.345058f
C535 sarlogic_0/FILLER_0_19_155/a_36_472# 0 0.404746f
C536 sarlogic_0/FILLER_0_19_155/a_572_375# 0 0.232991f
C537 sarlogic_0/FILLER_0_19_155/a_124_375# 0 0.185089f
C538 sarlogic_0/net11 0 1.328455f
C539 sarlogic_0/net21 0 1.922829f
C540 sarlogic_0/_007_ 0 0.309495f
C541 sarlogic_0/net77 0 1.39077f
C542 sarlogic_0/_418_/a_2560_156# 0 0.016968f
C543 sarlogic_0/_418_/a_2665_112# 0 0.62251f
C544 sarlogic_0/_418_/a_2248_156# 0 0.371662f
C545 sarlogic_0/_418_/a_1204_472# 0 0.012971f
C546 sarlogic_0/_418_/a_1000_472# 0 0.291735f
C547 sarlogic_0/_418_/a_796_472# 0 0.023206f
C548 sarlogic_0/_418_/a_1308_423# 0 0.279043f
C549 sarlogic_0/_418_/a_448_472# 0 0.684413f
C550 sarlogic_0/_418_/a_36_151# 0 1.43589f
C551 sarlogic_0/_220_/a_67_603# 0 0.345683f
C552 sarlogic_0/FILLER_0_9_282/a_484_472# 0 0.345058f
C553 sarlogic_0/FILLER_0_9_282/a_36_472# 0 0.404746f
C554 sarlogic_0/FILLER_0_9_282/a_572_375# 0 0.232991f
C555 sarlogic_0/FILLER_0_9_282/a_124_375# 0 0.185089f
C556 sarlogic_0/FILLER_0_18_37/a_1380_472# 0 0.345058f
C557 sarlogic_0/FILLER_0_18_37/a_932_472# 0 0.33241f
C558 sarlogic_0/FILLER_0_18_37/a_484_472# 0 0.33241f
C559 sarlogic_0/FILLER_0_18_37/a_36_472# 0 0.404746f
C560 sarlogic_0/FILLER_0_18_37/a_1468_375# 0 0.233029f
C561 sarlogic_0/FILLER_0_18_37/a_1020_375# 0 0.171606f
C562 sarlogic_0/FILLER_0_18_37/a_572_375# 0 0.171606f
C563 sarlogic_0/FILLER_0_18_37/a_124_375# 0 0.185399f
C564 sarlogic_0/FILLER_0_2_127/a_36_472# 0 0.417394f
C565 sarlogic_0/FILLER_0_2_127/a_124_375# 0 0.246306f
C566 sarlogic_0/_157_ 0 0.531763f
C567 sarlogic_0/_435_/a_2560_156# 0 0.016968f
C568 sarlogic_0/_435_/a_2665_112# 0 0.62251f
C569 sarlogic_0/_435_/a_2248_156# 0 0.371662f
C570 sarlogic_0/_435_/a_1204_472# 0 0.012971f
C571 sarlogic_0/_435_/a_1000_472# 0 0.291735f
C572 sarlogic_0/_435_/a_796_472# 0 0.023206f
C573 sarlogic_0/_435_/a_1308_423# 0 0.279043f
C574 sarlogic_0/_435_/a_448_472# 0 0.684413f
C575 sarlogic_0/_435_/a_36_151# 0 1.43589f
C576 sarlogic_0/_108_ 0 0.411979f
C577 sarlogic_0/_297_/a_36_472# 0 0.031137f
C578 sarlogic_0/trim_mask\[3\] 0 1.081535f
C579 sarlogic_0/_164_ 0 1.3268f
C580 sarlogic_0/_383_/a_36_472# 0 0.031137f
C581 sarlogic_0/_041_ 0 0.299289f
C582 sarlogic_0/_452_/a_2449_156# 0 0.049992f
C583 sarlogic_0/_452_/a_2225_156# 0 0.434082f
C584 sarlogic_0/_452_/a_3129_107# 0 0.58406f
C585 sarlogic_0/_452_/a_836_156# 0 0.019766f
C586 sarlogic_0/_452_/a_1040_527# 0 0.302082f
C587 sarlogic_0/_452_/a_1353_112# 0 0.286513f
C588 sarlogic_0/_452_/a_448_472# 0 1.21246f
C589 sarlogic_0/_452_/a_36_151# 0 1.31409f
C590 sarlogic_0/FILLER_0_6_79/a_36_472# 0 0.417394f
C591 sarlogic_0/FILLER_0_6_79/a_124_375# 0 0.246306f
C592 sarlogic_0/net59 0 5.044369f
C593 sarlogic_0/FILLER_0_15_59/a_484_472# 0 0.345058f
C594 sarlogic_0/FILLER_0_15_59/a_36_472# 0 0.404746f
C595 sarlogic_0/FILLER_0_15_59/a_572_375# 0 0.232991f
C596 sarlogic_0/FILLER_0_15_59/a_124_375# 0 0.185089f
C597 sarlogic_0/FILLER_0_3_221/a_1380_472# 0 0.345058f
C598 sarlogic_0/FILLER_0_3_221/a_932_472# 0 0.33241f
C599 sarlogic_0/FILLER_0_3_221/a_484_472# 0 0.33241f
C600 sarlogic_0/FILLER_0_3_221/a_36_472# 0 0.404746f
C601 sarlogic_0/FILLER_0_3_221/a_1468_375# 0 0.233029f
C602 sarlogic_0/FILLER_0_3_221/a_1020_375# 0 0.171606f
C603 sarlogic_0/FILLER_0_3_221/a_572_375# 0 0.171606f
C604 sarlogic_0/FILLER_0_3_221/a_124_375# 0 0.185399f
C605 sarlogic_0/FILLER_0_19_187/a_484_472# 0 0.345058f
C606 sarlogic_0/FILLER_0_19_187/a_36_472# 0 0.404746f
C607 sarlogic_0/FILLER_0_19_187/a_572_375# 0 0.232991f
C608 sarlogic_0/FILLER_0_19_187/a_124_375# 0 0.185089f
C609 sarlogic_0/FILLER_0_20_15/a_1380_472# 0 0.345058f
C610 sarlogic_0/FILLER_0_20_15/a_932_472# 0 0.33241f
C611 sarlogic_0/FILLER_0_20_15/a_484_472# 0 0.33241f
C612 sarlogic_0/FILLER_0_20_15/a_36_472# 0 0.404746f
C613 sarlogic_0/FILLER_0_20_15/a_1468_375# 0 0.233029f
C614 sarlogic_0/FILLER_0_20_15/a_1020_375# 0 0.171606f
C615 sarlogic_0/FILLER_0_20_15/a_572_375# 0 0.171606f
C616 sarlogic_0/FILLER_0_20_15/a_124_375# 0 0.185399f
C617 sarlogic_0/_204_/a_67_603# 0 0.345683f
C618 sarlogic_0/_419_/a_2560_156# 0 0.016968f
C619 sarlogic_0/_419_/a_2665_112# 0 0.62251f
C620 sarlogic_0/_419_/a_2248_156# 0 0.371662f
C621 sarlogic_0/_419_/a_1204_472# 0 0.012971f
C622 sarlogic_0/_419_/a_1000_472# 0 0.291735f
C623 sarlogic_0/_419_/a_796_472# 0 0.023206f
C624 sarlogic_0/_419_/a_1308_423# 0 0.279043f
C625 sarlogic_0/_419_/a_448_472# 0 0.684413f
C626 sarlogic_0/_419_/a_36_151# 0 1.43589f
C627 sarlogic_0/_054_ 0 0.522819f
C628 sarlogic_0/_221_/a_36_160# 0 0.386641f
C629 sarlogic_0/FILLER_0_9_270/a_484_472# 0 0.345058f
C630 sarlogic_0/FILLER_0_9_270/a_36_472# 0 0.404746f
C631 sarlogic_0/FILLER_0_9_270/a_572_375# 0 0.232991f
C632 sarlogic_0/FILLER_0_9_270/a_124_375# 0 0.185089f
C633 sarlogic_0/FILLER_0_1_192/a_36_472# 0 0.417394f
C634 sarlogic_0/FILLER_0_1_192/a_124_375# 0 0.246306f
C635 sarlogic_0/FILLER_0_13_80/a_36_472# 0 0.417394f
C636 sarlogic_0/FILLER_0_13_80/a_124_375# 0 0.246306f
C637 sarlogic_0/_153_ 0 1.165862f
C638 sarlogic_0/_154_ 0 1.167112f
C639 sarlogic_0/_367_/a_36_68# 0 0.150048f
C640 sarlogic_0/_436_/a_2560_156# 0 0.016968f
C641 sarlogic_0/_436_/a_2665_112# 0 0.62251f
C642 sarlogic_0/_436_/a_2248_156# 0 0.371662f
C643 sarlogic_0/_436_/a_1204_472# 0 0.012971f
C644 sarlogic_0/_436_/a_1000_472# 0 0.291735f
C645 sarlogic_0/_436_/a_796_472# 0 0.023206f
C646 sarlogic_0/_436_/a_1308_423# 0 0.279043f
C647 sarlogic_0/_436_/a_448_472# 0 0.684413f
C648 sarlogic_0/_436_/a_36_151# 0 1.43589f
C649 sarlogic_0/FILLER_0_10_107/a_484_472# 0 0.345058f
C650 sarlogic_0/FILLER_0_10_107/a_36_472# 0 0.404746f
C651 sarlogic_0/FILLER_0_10_107/a_572_375# 0 0.232991f
C652 sarlogic_0/FILLER_0_10_107/a_124_375# 0 0.185089f
C653 sarlogic_0/_168_ 0 0.336537f
C654 sarlogic_0/net51 0 2.105066f
C655 sarlogic_0/_042_ 0 0.323587f
C656 sarlogic_0/_453_/a_2560_156# 0 0.016968f
C657 sarlogic_0/_453_/a_2665_112# 0 0.62251f
C658 sarlogic_0/_453_/a_2248_156# 0 0.371662f
C659 sarlogic_0/_453_/a_1204_472# 0 0.012971f
C660 sarlogic_0/_453_/a_1000_472# 0 0.291735f
C661 sarlogic_0/_453_/a_796_472# 0 0.023206f
C662 sarlogic_0/_453_/a_1308_423# 0 0.279043f
C663 sarlogic_0/_453_/a_448_472# 0 0.684413f
C664 sarlogic_0/_453_/a_36_151# 0 1.43589f
C665 sarlogic_0/FILLER_0_19_142/a_36_472# 0 0.417394f
C666 sarlogic_0/FILLER_0_19_142/a_124_375# 0 0.246306f
C667 sarlogic_0/_048_ 0 0.358805f
C668 sarlogic_0/_205_/a_36_160# 0 0.696445f
C669 sarlogic_0/net43 0 1.236377f
C670 sarlogic_0/FILLER_0_3_78/a_484_472# 0 0.345058f
C671 sarlogic_0/FILLER_0_3_78/a_36_472# 0 0.404746f
C672 sarlogic_0/FILLER_0_3_78/a_572_375# 0 0.232991f
C673 sarlogic_0/FILLER_0_3_78/a_124_375# 0 0.185089f
C674 sarlogic_0/_437_/a_2560_156# 0 0.016968f
C675 sarlogic_0/_437_/a_2665_112# 0 0.62251f
C676 sarlogic_0/_437_/a_2248_156# 0 0.371662f
C677 sarlogic_0/_437_/a_1204_472# 0 0.012971f
C678 sarlogic_0/_437_/a_1000_472# 0 0.291735f
C679 sarlogic_0/_437_/a_796_472# 0 0.023206f
C680 sarlogic_0/_437_/a_1308_423# 0 0.279043f
C681 sarlogic_0/_437_/a_448_472# 0 0.684413f
C682 sarlogic_0/_437_/a_36_151# 0 1.43589f
C683 sarlogic_0/_109_ 0 0.319326f
C684 sarlogic_0/_299_/a_36_472# 0 0.031137f
C685 sarlogic_0/net37 0 1.529713f
C686 sarlogic_0/_385_/a_36_68# 0 0.112263f
C687 sarlogic_0/FILLER_0_0_266/a_36_472# 0 0.417394f
C688 sarlogic_0/FILLER_0_0_266/a_124_375# 0 0.246306f
C689 sarlogic_0/net12 0 1.263595f
C690 sarlogic_0/net22 0 2.108509f
C691 sarlogic_0/FILLER_0_9_290/a_36_472# 0 0.417394f
C692 sarlogic_0/FILLER_0_9_290/a_124_375# 0 0.246306f
C693 sarlogic_0/_223_/a_36_160# 0 0.696445f
C694 sarlogic_0/FILLER_0_14_263/a_36_472# 0 0.417394f
C695 sarlogic_0/FILLER_0_14_263/a_124_375# 0 0.246306f
C696 sarlogic_0/_158_ 0 0.309522f
C697 sarlogic_0/_369_/a_36_68# 0 0.150048f
C698 sarlogic_0/net71 0 1.420869f
C699 sarlogic_0/_438_/a_2560_156# 0 0.016968f
C700 sarlogic_0/_438_/a_2665_112# 0 0.62251f
C701 sarlogic_0/_438_/a_2248_156# 0 0.371662f
C702 sarlogic_0/_438_/a_1204_472# 0 0.012971f
C703 sarlogic_0/_438_/a_1000_472# 0 0.291735f
C704 sarlogic_0/_438_/a_796_472# 0 0.023206f
C705 sarlogic_0/_438_/a_1308_423# 0 0.279043f
C706 sarlogic_0/_438_/a_448_472# 0 0.684413f
C707 sarlogic_0/_438_/a_36_151# 0 1.43589f
C708 sarlogic_0/FILLER_0_23_274/a_36_472# 0 0.417394f
C709 sarlogic_0/FILLER_0_23_274/a_124_375# 0 0.246306f
C710 sarlogic_0/FILLER_0_17_282/a_36_472# 0 0.417394f
C711 sarlogic_0/FILLER_0_17_282/a_124_375# 0 0.246306f
C712 sarlogic_0/FILLER_0_5_198/a_484_472# 0 0.345058f
C713 sarlogic_0/FILLER_0_5_198/a_36_472# 0 0.404746f
C714 sarlogic_0/FILLER_0_5_198/a_572_375# 0 0.232991f
C715 sarlogic_0/FILLER_0_5_198/a_124_375# 0 0.185089f
C716 sarlogic_0/_163_ 0 1.03762f
C717 sarlogic_0/_169_ 0 0.245383f
C718 sarlogic_0/_386_/a_848_380# 0 0.40208f
C719 sarlogic_0/_386_/a_124_24# 0 0.591898f
C720 sarlogic_0/FILLER_0_20_2/a_484_472# 0 0.345058f
C721 sarlogic_0/FILLER_0_20_2/a_36_472# 0 0.404746f
C722 sarlogic_0/FILLER_0_20_2/a_572_375# 0 0.232991f
C723 sarlogic_0/FILLER_0_20_2/a_124_375# 0 0.185089f
C724 sarlogic_0/FILLER_0_16_154/a_1380_472# 0 0.345058f
C725 sarlogic_0/FILLER_0_16_154/a_932_472# 0 0.33241f
C726 sarlogic_0/FILLER_0_16_154/a_484_472# 0 0.33241f
C727 sarlogic_0/FILLER_0_16_154/a_36_472# 0 0.404746f
C728 sarlogic_0/FILLER_0_16_154/a_1468_375# 0 0.233029f
C729 sarlogic_0/FILLER_0_16_154/a_1020_375# 0 0.171606f
C730 sarlogic_0/FILLER_0_16_154/a_572_375# 0 0.171606f
C731 sarlogic_0/FILLER_0_16_154/a_124_375# 0 0.185399f
C732 sarlogic_0/FILLER_0_0_232/a_36_472# 0 0.417394f
C733 sarlogic_0/FILLER_0_0_232/a_124_375# 0 0.246306f
C734 sarlogic_0/FILLER_0_19_195/a_36_472# 0 0.417394f
C735 sarlogic_0/FILLER_0_19_195/a_124_375# 0 0.246306f
C736 sarlogic_0/_049_ 0 0.329957f
C737 sarlogic_0/net33 0 1.934915f
C738 sarlogic_0/_207_/a_67_603# 0 0.345683f
C739 sarlogic_0/FILLER_0_3_54/a_36_472# 0 0.417394f
C740 sarlogic_0/FILLER_0_3_54/a_124_375# 0 0.246306f
C741 sarlogic_0/FILLER_0_2_101/a_36_472# 0 0.417394f
C742 sarlogic_0/FILLER_0_2_101/a_124_375# 0 0.246306f
C743 sarlogic_0/trim_mask\[0\] 0 0.605753f
C744 sarlogic_0/_439_/a_2560_156# 0 0.016968f
C745 sarlogic_0/_439_/a_2665_112# 0 0.62251f
C746 sarlogic_0/_439_/a_2248_156# 0 0.371662f
C747 sarlogic_0/_439_/a_1204_472# 0 0.012971f
C748 sarlogic_0/_439_/a_1000_472# 0 0.291735f
C749 sarlogic_0/_439_/a_796_472# 0 0.023206f
C750 sarlogic_0/_439_/a_1308_423# 0 0.279043f
C751 sarlogic_0/_439_/a_448_472# 0 0.684413f
C752 sarlogic_0/_439_/a_36_151# 0 1.43589f
C753 sarlogic_0/_066_ 0 0.333041f
C754 sarlogic_0/FILLER_0_23_44/a_1380_472# 0 0.345058f
C755 sarlogic_0/FILLER_0_23_44/a_932_472# 0 0.33241f
C756 sarlogic_0/FILLER_0_23_44/a_484_472# 0 0.33241f
C757 sarlogic_0/FILLER_0_23_44/a_36_472# 0 0.404746f
C758 sarlogic_0/FILLER_0_23_44/a_1468_375# 0 0.233029f
C759 sarlogic_0/FILLER_0_23_44/a_1020_375# 0 0.171606f
C760 sarlogic_0/FILLER_0_23_44/a_572_375# 0 0.171606f
C761 sarlogic_0/FILLER_0_23_44/a_124_375# 0 0.185399f
C762 sarlogic_0/FILLER_0_23_88/a_36_472# 0 0.417394f
C763 sarlogic_0/FILLER_0_23_88/a_124_375# 0 0.246306f
C764 sarlogic_0/FILLER_0_5_164/a_484_472# 0 0.345058f
C765 sarlogic_0/FILLER_0_5_164/a_36_472# 0 0.404746f
C766 sarlogic_0/FILLER_0_5_164/a_572_375# 0 0.232991f
C767 sarlogic_0/FILLER_0_5_164/a_124_375# 0 0.185089f
C768 sarlogic_0/_060_ 0 2.485177f
C769 sarlogic_0/_113_ 0 2.833205f
C770 sarlogic_0/_090_ 0 2.629271f
C771 sarlogic_0/_310_/a_49_472# 0 0.098072f
C772 sarlogic_0/_037_ 0 0.467089f
C773 sarlogic_0/_170_ 0 0.413995f
C774 sarlogic_0/_387_/a_36_113# 0 0.418095f
C775 sarlogic_0/_208_/a_36_160# 0 0.696445f
C776 sarlogic_0/FILLER_0_18_76/a_484_472# 0 0.345058f
C777 sarlogic_0/FILLER_0_18_76/a_36_472# 0 0.404746f
C778 sarlogic_0/FILLER_0_18_76/a_572_375# 0 0.232991f
C779 sarlogic_0/FILLER_0_18_76/a_124_375# 0 0.185089f
C780 sarlogic_0/_225_/a_36_160# 0 0.386641f
C781 sarlogic_0/FILLER_0_2_177/a_484_472# 0 0.345058f
C782 sarlogic_0/FILLER_0_2_177/a_36_472# 0 0.404746f
C783 sarlogic_0/FILLER_0_2_177/a_572_375# 0 0.232991f
C784 sarlogic_0/FILLER_0_2_177/a_124_375# 0 0.185089f
C785 sarlogic_0/FILLER_0_2_111/a_1380_472# 0 0.345058f
C786 sarlogic_0/FILLER_0_2_111/a_932_472# 0 0.33241f
C787 sarlogic_0/FILLER_0_2_111/a_484_472# 0 0.33241f
C788 sarlogic_0/FILLER_0_2_111/a_36_472# 0 0.404746f
C789 sarlogic_0/FILLER_0_2_111/a_1468_375# 0 0.233029f
C790 sarlogic_0/FILLER_0_2_111/a_1020_375# 0 0.171606f
C791 sarlogic_0/FILLER_0_2_111/a_572_375# 0 0.171606f
C792 sarlogic_0/FILLER_0_2_111/a_124_375# 0 0.185399f
C793 sarlogic_0/FILLER_0_15_228/a_36_472# 0 0.417394f
C794 sarlogic_0/FILLER_0_15_228/a_124_375# 0 0.246306f
C795 sarlogic_0/net47 0 2.314376f
C796 sarlogic_0/_242_/a_36_160# 0 0.696445f
C797 sarlogic_0/_117_ 0 1.266251f
C798 sarlogic_0/_311_/a_66_473# 0 0.11665f
C799 sarlogic_0/_043_ 0 0.487279f
C800 sarlogic_0/_190_/a_36_160# 0 0.696445f
C801 sarlogic_0/FILLER_0_9_105/a_484_472# 0 0.345058f
C802 sarlogic_0/FILLER_0_9_105/a_36_472# 0 0.404746f
C803 sarlogic_0/FILLER_0_9_105/a_572_375# 0 0.232991f
C804 sarlogic_0/FILLER_0_9_105/a_124_375# 0 0.185089f
C805 sarlogic_0/FILLER_0_13_100/a_36_472# 0 0.417394f
C806 sarlogic_0/FILLER_0_13_100/a_124_375# 0 0.246306f
C807 sarlogic_0/FILLER_0_22_177/a_1380_472# 0 0.345058f
C808 sarlogic_0/FILLER_0_22_177/a_932_472# 0 0.33241f
C809 sarlogic_0/FILLER_0_22_177/a_484_472# 0 0.33241f
C810 sarlogic_0/FILLER_0_22_177/a_36_472# 0 0.404746f
C811 sarlogic_0/FILLER_0_22_177/a_1468_375# 0 0.233029f
C812 sarlogic_0/FILLER_0_22_177/a_1020_375# 0 0.171606f
C813 sarlogic_0/FILLER_0_22_177/a_572_375# 0 0.171606f
C814 sarlogic_0/FILLER_0_22_177/a_124_375# 0 0.185399f
C815 sarlogic_0/FILLER_0_15_2/a_484_472# 0 0.345058f
C816 sarlogic_0/FILLER_0_15_2/a_36_472# 0 0.404746f
C817 sarlogic_0/FILLER_0_15_2/a_572_375# 0 0.232991f
C818 sarlogic_0/FILLER_0_15_2/a_124_375# 0 0.185089f
C819 sarlogic_0/FILLER_0_15_10/a_36_472# 0 0.417394f
C820 sarlogic_0/FILLER_0_15_10/a_124_375# 0 0.246306f
C821 sarlogic_0/FILLER_0_19_171/a_1380_472# 0 0.345058f
C822 sarlogic_0/FILLER_0_19_171/a_932_472# 0 0.33241f
C823 sarlogic_0/FILLER_0_19_171/a_484_472# 0 0.33241f
C824 sarlogic_0/FILLER_0_19_171/a_36_472# 0 0.404746f
C825 sarlogic_0/FILLER_0_19_171/a_1468_375# 0 0.233029f
C826 sarlogic_0/FILLER_0_19_171/a_1020_375# 0 0.171606f
C827 sarlogic_0/FILLER_0_19_171/a_572_375# 0 0.171606f
C828 sarlogic_0/FILLER_0_19_171/a_124_375# 0 0.185399f
C829 sarlogic_0/net13 0 1.176306f
C830 sarlogic_0/net23 0 2.091399f
C831 sarlogic_0/FILLER_0_20_87/a_36_472# 0 0.417394f
C832 sarlogic_0/FILLER_0_20_87/a_124_375# 0 0.246306f
C833 sarlogic_0/FILLER_0_20_98/a_36_472# 0 0.417394f
C834 sarlogic_0/FILLER_0_20_98/a_124_375# 0 0.246306f
C835 sarlogic_0/_055_ 0 1.782885f
C836 sarlogic_0/FILLER_0_18_53/a_484_472# 0 0.345058f
C837 sarlogic_0/FILLER_0_18_53/a_36_472# 0 0.404746f
C838 sarlogic_0/FILLER_0_18_53/a_572_375# 0 0.232991f
C839 sarlogic_0/FILLER_0_18_53/a_124_375# 0 0.185089f
C840 sarlogic_0/FILLER_0_2_165/a_36_472# 0 0.417394f
C841 sarlogic_0/FILLER_0_2_165/a_124_375# 0 0.246306f
C842 sarlogic_0/FILLER_0_15_205/a_36_472# 0 0.417394f
C843 sarlogic_0/FILLER_0_15_205/a_124_375# 0 0.246306f
C844 sarlogic_0/FILLER_0_23_282/a_484_472# 0 0.345058f
C845 sarlogic_0/FILLER_0_23_282/a_36_472# 0 0.404746f
C846 sarlogic_0/FILLER_0_23_282/a_572_375# 0 0.232991f
C847 sarlogic_0/FILLER_0_23_282/a_124_375# 0 0.185089f
C848 sarlogic_0/net42 0 1.067446f
C849 sarlogic_0/net17 0 2.210219f
C850 sarlogic_0/_172_ 0 0.265782f
C851 sarlogic_0/_171_ 0 0.300355f
C852 sarlogic_0/_389_/a_36_148# 0 0.388358f
C853 sarlogic_0/_080_ 0 0.328202f
C854 sarlogic_0/_260_/a_36_68# 0 0.112263f
C855 sarlogic_0/FILLER_0_0_96/a_36_472# 0 0.417394f
C856 sarlogic_0/FILLER_0_0_96/a_124_375# 0 0.246306f
C857 sarlogic_0/FILLER_0_9_72/a_1380_472# 0 0.345058f
C858 sarlogic_0/FILLER_0_9_72/a_932_472# 0 0.33241f
C859 sarlogic_0/FILLER_0_9_72/a_484_472# 0 0.33241f
C860 sarlogic_0/FILLER_0_9_72/a_36_472# 0 0.404746f
C861 sarlogic_0/FILLER_0_9_72/a_1468_375# 0 0.233029f
C862 sarlogic_0/FILLER_0_9_72/a_1020_375# 0 0.171606f
C863 sarlogic_0/FILLER_0_9_72/a_572_375# 0 0.171606f
C864 sarlogic_0/FILLER_0_9_72/a_124_375# 0 0.185399f
C865 sarlogic_0/FILLER_0_20_31/a_36_472# 0 0.417394f
C866 sarlogic_0/FILLER_0_20_31/a_124_375# 0 0.246306f
C867 sarlogic_0/_227_/a_36_160# 0 0.386641f
C868 sarlogic_0/_120_ 0 1.533088f
C869 sarlogic_0/_313_/a_67_603# 0 0.345683f
C870 sarlogic_0/FILLER_0_5_172/a_36_472# 0 0.417394f
C871 sarlogic_0/FILLER_0_5_172/a_124_375# 0 0.246306f
C872 sarlogic_0/FILLER_0_12_20/a_484_472# 0 0.345058f
C873 sarlogic_0/FILLER_0_12_20/a_36_472# 0 0.404746f
C874 sarlogic_0/FILLER_0_12_20/a_572_375# 0 0.232991f
C875 sarlogic_0/FILLER_0_12_20/a_124_375# 0 0.185089f
C876 sarlogic_0/_134_ 0 0.365972f
C877 sarlogic_0/_062_ 0 1.717773f
C878 sarlogic_0/_059_ 0 1.686761f
C879 sarlogic_0/_261_/a_36_160# 0 0.386641f
C880 sarlogic_0/_044_ 0 0.388801f
C881 sarlogic_0/mask\[1\] 0 1.295078f
C882 sarlogic_0/_192_/a_67_603# 0 0.345683f
C883 sarlogic_0/FILLER_0_13_142/a_1380_472# 0 0.345058f
C884 sarlogic_0/FILLER_0_13_142/a_932_472# 0 0.33241f
C885 sarlogic_0/FILLER_0_13_142/a_484_472# 0 0.33241f
C886 sarlogic_0/FILLER_0_13_142/a_36_472# 0 0.404746f
C887 sarlogic_0/FILLER_0_13_142/a_1468_375# 0 0.233029f
C888 sarlogic_0/FILLER_0_13_142/a_1020_375# 0 0.171606f
C889 sarlogic_0/FILLER_0_13_142/a_572_375# 0 0.171606f
C890 sarlogic_0/FILLER_0_13_142/a_124_375# 0 0.185399f
C891 sarlogic_0/FILLER_0_9_60/a_484_472# 0 0.345058f
C892 sarlogic_0/FILLER_0_9_60/a_36_472# 0 0.404746f
C893 sarlogic_0/FILLER_0_9_60/a_572_375# 0 0.232991f
C894 sarlogic_0/FILLER_0_9_60/a_124_375# 0 0.185089f
C895 sarlogic_0/FILLER_0_7_233/a_36_472# 0 0.417394f
C896 sarlogic_0/FILLER_0_7_233/a_124_375# 0 0.246306f
C897 sarlogic_0/_228_/a_36_68# 0 0.69549f
C898 sarlogic_0/FILLER_0_21_206/a_36_472# 0 0.417394f
C899 sarlogic_0/FILLER_0_21_206/a_124_375# 0 0.246306f
C900 sarlogic_0/_067_ 0 0.851951f
C901 sarlogic_0/_135_ 0 0.339478f
C902 sarlogic_0/_193_/a_36_160# 0 0.696445f
C903 sarlogic_0/_180_ 0 0.390598f
C904 sarlogic_0/cal_count\[1\] 0 1.568289f
C905 sarlogic_0/FILLER_0_4_213/a_484_472# 0 0.345058f
C906 sarlogic_0/FILLER_0_4_213/a_36_472# 0 0.404746f
C907 sarlogic_0/FILLER_0_4_213/a_572_375# 0 0.232991f
C908 sarlogic_0/FILLER_0_4_213/a_124_375# 0 0.185089f
C909 sarlogic_0/FILLER_0_11_282/a_36_472# 0 0.417394f
C910 sarlogic_0/FILLER_0_11_282/a_124_375# 0 0.246306f
C911 sarlogic_0/FILLER_0_18_61/a_36_472# 0 0.417394f
C912 sarlogic_0/FILLER_0_18_61/a_124_375# 0 0.246306f
C913 sarlogic_0/FILLER_0_15_235/a_484_472# 0 0.345058f
C914 sarlogic_0/FILLER_0_15_235/a_36_472# 0 0.404746f
C915 sarlogic_0/FILLER_0_15_235/a_572_375# 0 0.232991f
C916 sarlogic_0/FILLER_0_15_235/a_124_375# 0 0.185089f
C917 sarlogic_0/FILLER_0_23_290/a_36_472# 0 0.417394f
C918 sarlogic_0/FILLER_0_23_290/a_124_375# 0 0.246306f
C919 sarlogic_0/_121_ 0 0.532847f
C920 sarlogic_0/_315_/a_36_68# 0 0.052951f
C921 sarlogic_0/_246_/a_36_68# 0 0.69549f
C922 sarlogic_0/FILLER_0_5_181/a_36_472# 0 0.417394f
C923 sarlogic_0/FILLER_0_5_181/a_124_375# 0 0.246306f
C924 sarlogic_0/_082_ 0 0.619901f
C925 sarlogic_0/net8 0 1.163723f
C926 sarlogic_0/net18 0 2.032159f
C927 sarlogic_0/_332_/a_36_472# 0 0.031137f
C928 sarlogic_0/_179_ 0 0.336984f
C929 sarlogic_0/_401_/a_36_68# 0 0.112263f
C930 sarlogic_0/FILLER_0_14_107/a_1380_472# 0 0.345058f
C931 sarlogic_0/FILLER_0_14_107/a_932_472# 0 0.33241f
C932 sarlogic_0/FILLER_0_14_107/a_484_472# 0 0.33241f
C933 sarlogic_0/FILLER_0_14_107/a_36_472# 0 0.404746f
C934 sarlogic_0/FILLER_0_14_107/a_1468_375# 0 0.233029f
C935 sarlogic_0/FILLER_0_14_107/a_1020_375# 0 0.171606f
C936 sarlogic_0/FILLER_0_14_107/a_572_375# 0 0.171606f
C937 sarlogic_0/FILLER_0_14_107/a_124_375# 0 0.185399f
C938 sarlogic_0/_097_ 0 0.592554f
C939 sarlogic_0/FILLER_0_1_204/a_36_472# 0 0.417394f
C940 sarlogic_0/FILLER_0_1_204/a_124_375# 0 0.246306f
C941 sarlogic_0/FILLER_0_15_72/a_484_472# 0 0.345058f
C942 sarlogic_0/FILLER_0_15_72/a_36_472# 0 0.404746f
C943 sarlogic_0/FILLER_0_15_72/a_572_375# 0 0.232991f
C944 sarlogic_0/FILLER_0_15_72/a_124_375# 0 0.185089f
C945 sarlogic_0/FILLER_0_17_104/a_1380_472# 0 0.345058f
C946 sarlogic_0/FILLER_0_17_104/a_932_472# 0 0.33241f
C947 sarlogic_0/FILLER_0_17_104/a_484_472# 0 0.33241f
C948 sarlogic_0/FILLER_0_17_104/a_36_472# 0 0.404746f
C949 sarlogic_0/FILLER_0_17_104/a_1468_375# 0 0.233029f
C950 sarlogic_0/FILLER_0_17_104/a_1020_375# 0 0.171606f
C951 sarlogic_0/FILLER_0_17_104/a_572_375# 0 0.171606f
C952 sarlogic_0/FILLER_0_17_104/a_124_375# 0 0.185399f
C953 sarlogic_0/FILLER_0_8_37/a_484_472# 0 0.345058f
C954 sarlogic_0/FILLER_0_8_37/a_36_472# 0 0.404746f
C955 sarlogic_0/FILLER_0_8_37/a_572_375# 0 0.232991f
C956 sarlogic_0/FILLER_0_8_37/a_124_375# 0 0.185089f
C957 sarlogic_0/FILLER_0_15_212/a_1380_472# 0 0.345058f
C958 sarlogic_0/FILLER_0_15_212/a_932_472# 0 0.33241f
C959 sarlogic_0/FILLER_0_15_212/a_484_472# 0 0.33241f
C960 sarlogic_0/FILLER_0_15_212/a_36_472# 0 0.404746f
C961 sarlogic_0/FILLER_0_15_212/a_1468_375# 0 0.233029f
C962 sarlogic_0/FILLER_0_15_212/a_1020_375# 0 0.171606f
C963 sarlogic_0/FILLER_0_15_212/a_572_375# 0 0.171606f
C964 sarlogic_0/FILLER_0_15_212/a_124_375# 0 0.185399f
C965 sarlogic_0/FILLER_0_23_60/a_36_472# 0 0.417394f
C966 sarlogic_0/FILLER_0_23_60/a_124_375# 0 0.246306f
C967 sarlogic_0/_123_ 0 0.344874f
C968 sarlogic_0/_122_ 0 0.600118f
C969 sarlogic_0/calibrate 0 1.343796f
C970 sarlogic_0/_316_/a_848_380# 0 0.40208f
C971 sarlogic_0/_316_/a_124_24# 0 0.591898f
C972 sarlogic_0/_247_/a_36_160# 0 0.696445f
C973 sarlogic_0/FILLER_0_12_50/a_36_472# 0 0.417394f
C974 sarlogic_0/FILLER_0_12_50/a_124_375# 0 0.246306f
C975 sarlogic_0/_084_ 0 0.296163f
C976 sarlogic_0/cal_itt\[0\] 0 1.831055f
C977 sarlogic_0/cal_itt\[1\] 0 1.705665f
C978 sarlogic_0/FILLER_0_11_109/a_36_472# 0 0.417394f
C979 sarlogic_0/FILLER_0_11_109/a_124_375# 0 0.246306f
C980 sarlogic_0/_182_ 0 0.34197f
C981 sarlogic_0/_402_/a_1948_68# 0 0.022025f
C982 sarlogic_0/_402_/a_718_527# 0 0.001795f
C983 sarlogic_0/_402_/a_56_567# 0 0.424713f
C984 sarlogic_0/_402_/a_728_93# 0 0.65929f
C985 sarlogic_0/_402_/a_1296_93# 0 0.317801f
C986 sarlogic_0/_045_ 0 0.349338f
C987 sarlogic_0/mask\[2\] 0 1.335688f
C988 sarlogic_0/_195_/a_67_603# 0 0.345683f
C989 sarlogic_0/_333_/a_36_160# 0 0.386641f
C990 sarlogic_0/_098_ 0 1.816151f
C991 sarlogic_0/_147_ 0 0.322539f
C992 sarlogic_0/_350_/a_49_472# 0 0.054843f
C993 sarlogic_0/FILLER_0_12_236/a_484_472# 0 0.345058f
C994 sarlogic_0/FILLER_0_12_236/a_36_472# 0 0.404746f
C995 sarlogic_0/FILLER_0_12_236/a_572_375# 0 0.232991f
C996 sarlogic_0/FILLER_0_12_236/a_124_375# 0 0.185089f
C997 sarlogic_0/FILLER_0_2_171/a_36_472# 0 0.417394f
C998 sarlogic_0/FILLER_0_2_171/a_124_375# 0 0.246306f
C999 sarlogic_0/_014_ 0 0.363432f
C1000 sarlogic_0/_317_/a_36_113# 0 0.418095f
C1001 sarlogic_0/_248_/a_36_68# 0 0.69549f
C1002 sarlogic_0/FILLER_0_17_38/a_484_472# 0 0.345058f
C1003 sarlogic_0/FILLER_0_17_38/a_36_472# 0 0.404746f
C1004 sarlogic_0/FILLER_0_17_38/a_572_375# 0 0.232991f
C1005 sarlogic_0/FILLER_0_17_38/a_124_375# 0 0.185089f
C1006 sarlogic_0/_001_ 0 0.285216f
C1007 sarlogic_0/_265_/a_244_68# 0 0.138666f
C1008 sarlogic_0/_196_/a_36_160# 0 0.696445f
C1009 sarlogic_0/FILLER_0_6_90/a_484_472# 0 0.345058f
C1010 sarlogic_0/FILLER_0_6_90/a_36_472# 0 0.404746f
C1011 sarlogic_0/FILLER_0_6_90/a_572_375# 0 0.232991f
C1012 sarlogic_0/FILLER_0_6_90/a_124_375# 0 0.185089f
C1013 sarlogic_0/_183_ 0 0.356629f
C1014 sarlogic_0/_334_/a_36_160# 0 0.386641f
C1015 sarlogic_0/_282_/a_36_160# 0 0.386641f
C1016 sarlogic_0/_024_ 0 0.451815f
C1017 sarlogic_0/_009_ 0 0.397943f
C1018 sarlogic_0/_420_/a_2560_156# 0 0.016968f
C1019 sarlogic_0/_420_/a_2665_112# 0 0.62251f
C1020 sarlogic_0/_420_/a_2248_156# 0 0.371662f
C1021 sarlogic_0/_420_/a_1204_472# 0 0.012971f
C1022 sarlogic_0/_420_/a_1000_472# 0 0.291735f
C1023 sarlogic_0/_420_/a_796_472# 0 0.023206f
C1024 sarlogic_0/_420_/a_1308_423# 0 0.279043f
C1025 sarlogic_0/_420_/a_448_472# 0 0.684413f
C1026 sarlogic_0/_420_/a_36_151# 0 1.43589f
C1027 clk 0 17.49988f
C1028 sarlogic_0/FILLER_0_8_2/a_36_472# 0 0.417394f
C1029 sarlogic_0/FILLER_0_8_2/a_124_375# 0 0.246306f
C1030 sarlogic_0/FILLER_0_8_24/a_484_472# 0 0.345058f
C1031 sarlogic_0/FILLER_0_8_24/a_36_472# 0 0.404746f
C1032 sarlogic_0/FILLER_0_8_24/a_572_375# 0 0.232991f
C1033 sarlogic_0/FILLER_0_8_24/a_124_375# 0 0.185089f
C1034 sarlogic_0/_124_ 0 0.294081f
C1035 sarlogic_0/_118_ 0 1.378735f
C1036 sarlogic_0/_071_ 0 1.600488f
C1037 sarlogic_0/net9 0 1.13171f
C1038 sarlogic_0/net19 0 1.889339f
C1039 sarlogic_0/_138_ 0 0.33132f
C1040 sarlogic_0/_137_ 0 1.178616f
C1041 sarlogic_0/_335_/a_49_472# 0 0.054843f
C1042 sarlogic_0/_404_/a_36_472# 0 0.031137f
C1043 sarlogic_0/FILLER_0_20_107/a_36_472# 0 0.417394f
C1044 sarlogic_0/FILLER_0_20_107/a_124_375# 0 0.246306f
C1045 sarlogic_0/FILLER_0_9_142/a_36_472# 0 0.417394f
C1046 sarlogic_0/FILLER_0_9_142/a_124_375# 0 0.246306f
C1047 sarlogic_0/_099_ 0 1.152785f
C1048 sarlogic_0/_283_/a_36_472# 0 0.031137f
C1049 sarlogic_0/mask\[7\] 0 1.477838f
C1050 sarlogic_0/_352_/a_49_472# 0 0.054843f
C1051 sarlogic_0/_010_ 0 0.377779f
C1052 sarlogic_0/_421_/a_2560_156# 0 0.016968f
C1053 sarlogic_0/_421_/a_2665_112# 0 0.62251f
C1054 sarlogic_0/_421_/a_2248_156# 0 0.371662f
C1055 sarlogic_0/_421_/a_1204_472# 0 0.012971f
C1056 sarlogic_0/_421_/a_1000_472# 0 0.291735f
C1057 sarlogic_0/_421_/a_796_472# 0 0.023206f
C1058 sarlogic_0/_421_/a_1308_423# 0 0.279043f
C1059 sarlogic_0/_421_/a_448_472# 0 0.684413f
C1060 sarlogic_0/_421_/a_36_151# 0 1.43589f
C1061 sarlogic_0/FILLER_0_1_212/a_36_472# 0 0.417394f
C1062 sarlogic_0/FILLER_0_1_212/a_124_375# 0 0.246306f
C1063 sarlogic_0/FILLER_0_8_239/a_36_472# 0 0.417394f
C1064 sarlogic_0/FILLER_0_8_239/a_124_375# 0 0.246306f
C1065 sarlogic_0/_125_ 0 1.526603f
C1066 sarlogic_0/_058_ 0 1.483584f
C1067 sarlogic_0/FILLER_0_6_177/a_484_472# 0 0.345058f
C1068 sarlogic_0/FILLER_0_6_177/a_36_472# 0 0.404746f
C1069 sarlogic_0/FILLER_0_6_177/a_572_375# 0 0.232991f
C1070 sarlogic_0/FILLER_0_6_177/a_124_375# 0 0.185089f
C1071 sarlogic_0/state\[1\] 0 2.652405f
C1072 sarlogic_0/_267_/a_36_472# 0 0.137725f
C1073 sarlogic_0/_184_ 0 0.350066f
C1074 sarlogic_0/cal_count\[2\] 0 1.971854f
C1075 sarlogic_0/_405_/a_67_603# 0 0.345683f
C1076 sarlogic_0/_018_ 0 0.358633f
C1077 sarlogic_0/_046_ 0 0.361963f
C1078 sarlogic_0/_198_/a_67_603# 0 0.345683f
C1079 sarlogic_0/_094_ 0 1.263877f
C1080 sarlogic_0/_100_ 0 0.333135f
C1081 sarlogic_0/net36 0 2.262756f
C1082 sarlogic_0/FILLER_0_17_133/a_36_472# 0 0.417394f
C1083 sarlogic_0/FILLER_0_17_133/a_124_375# 0 0.246306f
C1084 sarlogic_0/_025_ 0 0.350324f
C1085 sarlogic_0/_148_ 0 0.325709f
C1086 sarlogic_0/_422_/a_2560_156# 0 0.016968f
C1087 sarlogic_0/_422_/a_2665_112# 0 0.62251f
C1088 sarlogic_0/_422_/a_2248_156# 0 0.371662f
C1089 sarlogic_0/_422_/a_1204_472# 0 0.012971f
C1090 sarlogic_0/_422_/a_1000_472# 0 0.291735f
C1091 sarlogic_0/_422_/a_796_472# 0 0.023206f
C1092 sarlogic_0/_422_/a_1308_423# 0 0.279043f
C1093 sarlogic_0/_422_/a_448_472# 0 0.684413f
C1094 sarlogic_0/_422_/a_36_151# 0 1.43589f
C1095 sarlogic_0/FILLER_0_1_266/a_484_472# 0 0.345058f
C1096 sarlogic_0/FILLER_0_1_266/a_36_472# 0 0.404746f
C1097 sarlogic_0/FILLER_0_1_266/a_572_375# 0 0.232991f
C1098 sarlogic_0/FILLER_0_1_266/a_124_375# 0 0.185089f
C1099 sarlogic_0/_152_ 0 0.918583f
C1100 sarlogic_0/_081_ 0 1.140656f
C1101 sarlogic_0/_370_/a_848_380# 0 0.40208f
C1102 sarlogic_0/_370_/a_124_24# 0 0.591898f
C1103 sarlogic_0/FILLER_0_24_274/a_1380_472# 0 0.345058f
C1104 sarlogic_0/FILLER_0_24_274/a_932_472# 0 0.33241f
C1105 sarlogic_0/FILLER_0_24_274/a_484_472# 0 0.33241f
C1106 sarlogic_0/FILLER_0_24_274/a_36_472# 0 0.404746f
C1107 sarlogic_0/FILLER_0_24_274/a_1468_375# 0 0.233029f
C1108 sarlogic_0/FILLER_0_24_274/a_1020_375# 0 0.171606f
C1109 sarlogic_0/FILLER_0_24_274/a_572_375# 0 0.171606f
C1110 sarlogic_0/FILLER_0_24_274/a_124_375# 0 0.185399f
C1111 sarlogic_0/_185_ 0 0.386917f
C1112 sarlogic_0/_406_/a_36_159# 0 0.374116f
C1113 sarlogic_0/_337_/a_49_472# 0 0.054843f
C1114 sarlogic_0/_199_/a_36_160# 0 0.696445f
C1115 sarlogic_0/_285_/a_36_472# 0 0.031137f
C1116 sarlogic_0/_354_/a_49_472# 0 0.054843f
C1117 sarlogic_0/_012_ 0 0.75195f
C1118 sarlogic_0/_423_/a_2560_156# 0 0.016968f
C1119 sarlogic_0/_423_/a_2665_112# 0 0.62251f
C1120 sarlogic_0/_423_/a_2248_156# 0 0.371662f
C1121 sarlogic_0/_423_/a_1204_472# 0 0.012971f
C1122 sarlogic_0/_423_/a_1000_472# 0 0.291735f
C1123 sarlogic_0/_423_/a_796_472# 0 0.023206f
C1124 sarlogic_0/_423_/a_1308_423# 0 0.279043f
C1125 sarlogic_0/_423_/a_448_472# 0 0.684413f
C1126 sarlogic_0/_423_/a_36_151# 0 1.43589f
C1127 sarlogic_0/FILLER_0_5_88/a_36_472# 0 0.417394f
C1128 sarlogic_0/FILLER_0_5_88/a_124_375# 0 0.246306f
C1129 sarlogic_0/trim_mask\[1\] 0 1.020743f
C1130 sarlogic_0/_029_ 0 0.308904f
C1131 sarlogic_0/_440_/a_2560_156# 0 0.016968f
C1132 sarlogic_0/_440_/a_2665_112# 0 0.62251f
C1133 sarlogic_0/_440_/a_2248_156# 0 0.371662f
C1134 sarlogic_0/_440_/a_1204_472# 0 0.012971f
C1135 sarlogic_0/_440_/a_1000_472# 0 0.291735f
C1136 sarlogic_0/_440_/a_796_472# 0 0.023206f
C1137 sarlogic_0/_440_/a_1308_423# 0 0.279043f
C1138 sarlogic_0/_440_/a_448_472# 0 0.684413f
C1139 sarlogic_0/_440_/a_36_151# 0 1.43589f
C1140 sarlogic_0/_159_ 0 0.351814f
C1141 sarlogic_0/_371_/a_36_113# 0 0.418095f
C1142 sarlogic_0/FILLER_0_17_56/a_484_472# 0 0.345058f
C1143 sarlogic_0/FILLER_0_17_56/a_36_472# 0 0.404746f
C1144 sarlogic_0/FILLER_0_17_56/a_572_375# 0 0.232991f
C1145 sarlogic_0/FILLER_0_17_56/a_124_375# 0 0.185089f
C1146 sarlogic_0/_083_ 0 0.527882f
C1147 sarlogic_0/_078_ 0 0.904554f
C1148 sarlogic_0/_269_/a_36_472# 0 0.031137f
C1149 sarlogic_0/_181_ 0 0.829168f
C1150 sarlogic_0/_407_/a_36_472# 0 0.031137f
C1151 sarlogic_0/_019_ 0 0.32907f
C1152 sarlogic_0/_139_ 0 0.346404f
C1153 sarlogic_0/FILLER_0_14_123/a_36_472# 0 0.417394f
C1154 sarlogic_0/FILLER_0_14_123/a_124_375# 0 0.246306f
C1155 sarlogic_0/_005_ 0 0.340993f
C1156 sarlogic_0/_101_ 0 0.280497f
C1157 sarlogic_0/_424_/a_2560_156# 0 0.016968f
C1158 sarlogic_0/_424_/a_2665_112# 0 0.62251f
C1159 sarlogic_0/_424_/a_2248_156# 0 0.371662f
C1160 sarlogic_0/_424_/a_1204_472# 0 0.012971f
C1161 sarlogic_0/_424_/a_1000_472# 0 0.291735f
C1162 sarlogic_0/_424_/a_796_472# 0 0.023206f
C1163 sarlogic_0/_424_/a_1308_423# 0 0.279043f
C1164 sarlogic_0/_424_/a_448_472# 0 0.684413f
C1165 sarlogic_0/_424_/a_36_151# 0 1.43589f
C1166 sarlogic_0/_026_ 0 0.320379f
C1167 sarlogic_0/_149_ 0 0.305496f
C1168 sarlogic_0/FILLER_0_5_54/a_1380_472# 0 0.345058f
C1169 sarlogic_0/FILLER_0_5_54/a_932_472# 0 0.33241f
C1170 sarlogic_0/FILLER_0_5_54/a_484_472# 0 0.33241f
C1171 sarlogic_0/FILLER_0_5_54/a_36_472# 0 0.404746f
C1172 sarlogic_0/FILLER_0_5_54/a_1468_375# 0 0.233029f
C1173 sarlogic_0/FILLER_0_5_54/a_1020_375# 0 0.171606f
C1174 sarlogic_0/FILLER_0_5_54/a_572_375# 0 0.171606f
C1175 sarlogic_0/FILLER_0_5_54/a_124_375# 0 0.185399f
C1176 sarlogic_0/FILLER_0_17_142/a_484_472# 0 0.345058f
C1177 sarlogic_0/FILLER_0_17_142/a_36_472# 0 0.404746f
C1178 sarlogic_0/FILLER_0_17_142/a_572_375# 0 0.232991f
C1179 sarlogic_0/FILLER_0_17_142/a_124_375# 0 0.185089f
C1180 sarlogic_0/_068_ 0 3.162692f
C1181 sarlogic_0/_076_ 0 3.812442f
C1182 sarlogic_0/_133_ 0 1.430901f
C1183 sarlogic_0/_070_ 0 3.115722f
C1184 sarlogic_0/_372_/a_170_472# 0 0.077257f
C1185 sarlogic_0/net49 0 5.140563f
C1186 sarlogic_0/_030_ 0 0.307083f
C1187 sarlogic_0/net66 0 1.472669f
C1188 sarlogic_0/_441_/a_2560_156# 0 0.016968f
C1189 sarlogic_0/_441_/a_2665_112# 0 0.62251f
C1190 sarlogic_0/_441_/a_2248_156# 0 0.371662f
C1191 sarlogic_0/_441_/a_1204_472# 0 0.012971f
C1192 sarlogic_0/_441_/a_1000_472# 0 0.291735f
C1193 sarlogic_0/_441_/a_796_472# 0 0.023206f
C1194 sarlogic_0/_441_/a_1308_423# 0 0.279043f
C1195 sarlogic_0/_441_/a_448_472# 0 0.684413f
C1196 sarlogic_0/_441_/a_36_151# 0 1.43589f
C1197 sarlogic_0/FILLER_0_5_206/a_36_472# 0 0.417394f
C1198 sarlogic_0/FILLER_0_5_206/a_124_375# 0 0.246306f
C1199 sarlogic_0/fanout49/a_36_160# 0 0.696445f
C1200 sarlogic_0/FILLER_0_8_247/a_1380_472# 0 0.345058f
C1201 sarlogic_0/FILLER_0_8_247/a_932_472# 0 0.33241f
C1202 sarlogic_0/FILLER_0_8_247/a_484_472# 0 0.33241f
C1203 sarlogic_0/FILLER_0_8_247/a_36_472# 0 0.404746f
C1204 sarlogic_0/FILLER_0_8_247/a_1468_375# 0 0.233029f
C1205 sarlogic_0/FILLER_0_8_247/a_1020_375# 0 0.171606f
C1206 sarlogic_0/FILLER_0_8_247/a_572_375# 0 0.171606f
C1207 sarlogic_0/FILLER_0_8_247/a_124_375# 0 0.185399f
C1208 sarlogic_0/FILLER_0_12_220/a_1380_472# 0 0.345058f
C1209 sarlogic_0/FILLER_0_12_220/a_932_472# 0 0.33241f
C1210 sarlogic_0/FILLER_0_12_220/a_484_472# 0 0.33241f
C1211 sarlogic_0/FILLER_0_12_220/a_36_472# 0 0.404746f
C1212 sarlogic_0/FILLER_0_12_220/a_1468_375# 0 0.233029f
C1213 sarlogic_0/FILLER_0_12_220/a_1020_375# 0 0.171606f
C1214 sarlogic_0/FILLER_0_12_220/a_572_375# 0 0.171606f
C1215 sarlogic_0/FILLER_0_12_220/a_124_375# 0 0.185399f
C1216 sarlogic_0/FILLER_0_21_286/a_484_472# 0 0.345058f
C1217 sarlogic_0/FILLER_0_21_286/a_36_472# 0 0.404746f
C1218 sarlogic_0/FILLER_0_21_286/a_572_375# 0 0.232991f
C1219 sarlogic_0/FILLER_0_21_286/a_124_375# 0 0.185089f
C1220 sarlogic_0/_140_ 0 1.276518f
C1221 sarlogic_0/_339_/a_36_160# 0 0.386641f
C1222 sarlogic_0/_095_ 0 2.689027f
C1223 sarlogic_0/_186_ 0 0.580923f
C1224 sarlogic_0/_408_/a_1936_472# 0 0.009918f
C1225 sarlogic_0/_408_/a_718_524# 0 0.005143f
C1226 sarlogic_0/_408_/a_56_524# 0 0.41096f
C1227 sarlogic_0/_408_/a_728_93# 0 0.654825f
C1228 sarlogic_0/_408_/a_1336_472# 0 0.316639f
C1229 sarlogic_0/FILLER_0_20_169/a_36_472# 0 0.417394f
C1230 sarlogic_0/FILLER_0_20_169/a_124_375# 0 0.246306f
C1231 sarlogic_0/_210_/a_67_603# 0 0.345683f
C1232 sarlogic_0/_425_/a_2560_156# 0 0.016968f
C1233 sarlogic_0/_425_/a_2665_112# 0 0.62251f
C1234 sarlogic_0/_425_/a_2248_156# 0 0.371662f
C1235 sarlogic_0/_425_/a_1204_472# 0 0.012971f
C1236 sarlogic_0/_425_/a_1000_472# 0 0.291735f
C1237 sarlogic_0/_425_/a_796_472# 0 0.023206f
C1238 sarlogic_0/_425_/a_1308_423# 0 0.279043f
C1239 sarlogic_0/_425_/a_448_472# 0 0.684413f
C1240 sarlogic_0/_425_/a_36_151# 0 1.43589f
C1241 sarlogic_0/net5 0 0.610761f
C1242 sarlogic_0/input5/a_36_113# 0 0.418095f
C1243 sarlogic_0/FILLER_0_11_78/a_484_472# 0 0.345058f
C1244 sarlogic_0/FILLER_0_11_78/a_36_472# 0 0.404746f
C1245 sarlogic_0/FILLER_0_11_78/a_572_375# 0 0.232991f
C1246 sarlogic_0/FILLER_0_11_78/a_124_375# 0 0.185089f
C1247 sarlogic_0/_102_ 0 0.335308f
C1248 sarlogic_0/_287_/a_36_472# 0 0.031137f
C1249 sarlogic_0/mask\[9\] 0 1.383606f
C1250 sarlogic_0/_356_/a_36_472# 0 0.031137f
C1251 sarlogic_0/_031_ 0 0.417351f
C1252 sarlogic_0/net69 0 1.020293f
C1253 sarlogic_0/_442_/a_2560_156# 0 0.016968f
C1254 sarlogic_0/_442_/a_2665_112# 0 0.62251f
C1255 sarlogic_0/_442_/a_2248_156# 0 0.371662f
C1256 sarlogic_0/_442_/a_1204_472# 0 0.012971f
C1257 sarlogic_0/_442_/a_1000_472# 0 0.291735f
C1258 sarlogic_0/_442_/a_796_472# 0 0.023206f
C1259 sarlogic_0/_442_/a_1308_423# 0 0.279043f
C1260 sarlogic_0/_442_/a_448_472# 0 0.684413f
C1261 sarlogic_0/_442_/a_36_151# 0 1.43589f
C1262 sarlogic_0/net64 0 2.598514f
C1263 sarlogic_0/fanout59/a_36_160# 0 0.696445f
C1264 sarlogic_0/FILLER_0_14_99/a_36_472# 0 0.417394f
C1265 sarlogic_0/FILLER_0_14_99/a_124_375# 0 0.246306f
C1266 sarlogic_0/_038_ 0 0.362839f
C1267 sarlogic_0/_136_ 0 1.345638f
C1268 sarlogic_0/_390_/a_36_68# 0 0.150048f
C1269 sarlogic_0/FILLER_0_15_282/a_484_472# 0 0.345058f
C1270 sarlogic_0/FILLER_0_15_282/a_36_472# 0 0.404746f
C1271 sarlogic_0/FILLER_0_15_282/a_572_375# 0 0.232991f
C1272 sarlogic_0/FILLER_0_15_282/a_124_375# 0 0.185089f
C1273 sarlogic_0/FILLER_0_11_124/a_36_472# 0 0.417394f
C1274 sarlogic_0/FILLER_0_11_124/a_124_375# 0 0.246306f
C1275 sarlogic_0/FILLER_0_11_135/a_36_472# 0 0.417394f
C1276 sarlogic_0/FILLER_0_11_135/a_124_375# 0 0.246306f
C1277 sarlogic_0/_188_ 0 0.349407f
C1278 sarlogic_0/cal_count\[3\] 0 1.862896f
C1279 sarlogic_0/_050_ 0 0.622354f
C1280 sarlogic_0/_211_/a_36_160# 0 0.386641f
C1281 sarlogic_0/net4 0 2.711508f
C1282 en 0 17.135206f
C1283 sarlogic_0/input4/a_36_68# 0 0.69549f
C1284 sarlogic_0/_426_/a_2560_156# 0 0.016968f
C1285 sarlogic_0/_426_/a_2665_112# 0 0.62251f
C1286 sarlogic_0/_426_/a_2248_156# 0 0.371662f
C1287 sarlogic_0/_426_/a_1204_472# 0 0.012971f
C1288 sarlogic_0/_426_/a_1000_472# 0 0.291735f
C1289 sarlogic_0/_426_/a_796_472# 0 0.023206f
C1290 sarlogic_0/_426_/a_1308_423# 0 0.279043f
C1291 sarlogic_0/_426_/a_448_472# 0 0.684413f
C1292 sarlogic_0/_426_/a_36_151# 0 1.43589f
C1293 sarlogic_0/_027_ 0 0.302949f
C1294 sarlogic_0/_150_ 0 0.320497f
C1295 sarlogic_0/FILLER_0_18_107/a_3172_472# 0 0.345058f
C1296 sarlogic_0/FILLER_0_18_107/a_2724_472# 0 0.33241f
C1297 sarlogic_0/FILLER_0_18_107/a_2276_472# 0 0.33241f
C1298 sarlogic_0/FILLER_0_18_107/a_1828_472# 0 0.33241f
C1299 sarlogic_0/FILLER_0_18_107/a_1380_472# 0 0.33241f
C1300 sarlogic_0/FILLER_0_18_107/a_932_472# 0 0.33241f
C1301 sarlogic_0/FILLER_0_18_107/a_484_472# 0 0.33241f
C1302 sarlogic_0/FILLER_0_18_107/a_36_472# 0 0.404746f
C1303 sarlogic_0/FILLER_0_18_107/a_3260_375# 0 0.233093f
C1304 sarlogic_0/FILLER_0_18_107/a_2812_375# 0 0.17167f
C1305 sarlogic_0/FILLER_0_18_107/a_2364_375# 0 0.17167f
C1306 sarlogic_0/FILLER_0_18_107/a_1916_375# 0 0.17167f
C1307 sarlogic_0/FILLER_0_18_107/a_1468_375# 0 0.17167f
C1308 sarlogic_0/FILLER_0_18_107/a_1020_375# 0 0.17167f
C1309 sarlogic_0/FILLER_0_18_107/a_572_375# 0 0.17167f
C1310 sarlogic_0/FILLER_0_18_107/a_124_375# 0 0.185915f
C1311 sarlogic_0/trim_mask\[4\] 0 0.987791f
C1312 sarlogic_0/_032_ 0 0.34876f
C1313 sarlogic_0/_443_/a_2560_156# 0 0.016968f
C1314 sarlogic_0/_443_/a_2665_112# 0 0.62251f
C1315 sarlogic_0/_443_/a_2248_156# 0 0.371662f
C1316 sarlogic_0/_443_/a_1204_472# 0 0.012971f
C1317 sarlogic_0/_443_/a_1000_472# 0 0.291735f
C1318 sarlogic_0/_443_/a_796_472# 0 0.023206f
C1319 sarlogic_0/_443_/a_1308_423# 0 0.279043f
C1320 sarlogic_0/_443_/a_448_472# 0 0.684413f
C1321 sarlogic_0/_443_/a_36_151# 0 1.43589f
C1322 sarlogic_0/_061_ 0 0.84986f
C1323 sarlogic_0/_056_ 0 2.393362f
C1324 sarlogic_0/_374_/a_36_68# 0 0.112263f
C1325 sarlogic_0/fanout58/a_36_160# 0 0.696445f
C1326 sarlogic_0/net74 0 1.237373f
C1327 sarlogic_0/fanout69/a_36_113# 0 0.418095f
C1328 sarlogic_0/_173_ 0 0.339446f
C1329 sarlogic_0/FILLER_0_3_142/a_36_472# 0 0.417394f
C1330 sarlogic_0/FILLER_0_3_142/a_124_375# 0 0.246306f
C1331 sarlogic_0/FILLER_0_17_64/a_36_472# 0 0.417394f
C1332 sarlogic_0/FILLER_0_17_64/a_124_375# 0 0.246306f
C1333 sarlogic_0/FILLER_0_11_101/a_484_472# 0 0.345058f
C1334 sarlogic_0/FILLER_0_11_101/a_36_472# 0 0.404746f
C1335 sarlogic_0/FILLER_0_11_101/a_572_375# 0 0.232991f
C1336 sarlogic_0/FILLER_0_11_101/a_124_375# 0 0.185089f
C1337 sarlogic_0/FILLER_0_22_86/a_1380_472# 0 0.345058f
C1338 sarlogic_0/FILLER_0_22_86/a_932_472# 0 0.33241f
C1339 sarlogic_0/FILLER_0_22_86/a_484_472# 0 0.33241f
C1340 sarlogic_0/FILLER_0_22_86/a_36_472# 0 0.404746f
C1341 sarlogic_0/FILLER_0_22_86/a_1468_375# 0 0.233029f
C1342 sarlogic_0/FILLER_0_22_86/a_1020_375# 0 0.171606f
C1343 sarlogic_0/FILLER_0_22_86/a_572_375# 0 0.171606f
C1344 sarlogic_0/FILLER_0_22_86/a_124_375# 0 0.185399f
C1345 sarlogic_0/net24 0 1.61895f
C1346 sarlogic_0/net3 0 0.740676f
C1347 sarlogic_0/input3/a_36_113# 0 0.418095f
C1348 sarlogic_0/_103_ 0 0.350464f
C1349 sarlogic_0/_289_/a_36_472# 0 0.031137f
C1350 sarlogic_0/_151_ 0 0.300777f
C1351 sarlogic_0/_427_/a_2560_156# 0 0.016968f
C1352 sarlogic_0/_427_/a_2665_112# 0 0.91969f
C1353 sarlogic_0/_427_/a_2248_156# 0 0.30886f
C1354 sarlogic_0/_427_/a_1204_472# 0 0.012971f
C1355 sarlogic_0/_427_/a_1000_472# 0 0.291735f
C1356 sarlogic_0/_427_/a_796_472# 0 0.023206f
C1357 sarlogic_0/_427_/a_1308_423# 0 0.279043f
C1358 sarlogic_0/_427_/a_448_472# 0 0.684413f
C1359 sarlogic_0/_427_/a_36_151# 0 1.43587f
C1360 sarlogic_0/FILLER_0_17_161/a_36_472# 0 0.417394f
C1361 sarlogic_0/FILLER_0_17_161/a_124_375# 0 0.246306f
C1362 sarlogic_0/FILLER_0_18_139/a_1380_472# 0 0.345058f
C1363 sarlogic_0/FILLER_0_18_139/a_932_472# 0 0.33241f
C1364 sarlogic_0/FILLER_0_18_139/a_484_472# 0 0.33241f
C1365 sarlogic_0/FILLER_0_18_139/a_36_472# 0 0.404746f
C1366 sarlogic_0/FILLER_0_18_139/a_1468_375# 0 0.233029f
C1367 sarlogic_0/FILLER_0_18_139/a_1020_375# 0 0.171606f
C1368 sarlogic_0/FILLER_0_18_139/a_572_375# 0 0.171606f
C1369 sarlogic_0/FILLER_0_18_139/a_124_375# 0 0.185399f
C1370 sarlogic_0/_161_ 0 0.592909f
C1371 sarlogic_0/_162_ 0 0.597238f
C1372 sarlogic_0/_375_/a_36_68# 0 0.048026f
C1373 sarlogic_0/trim_val\[0\] 0 0.742779f
C1374 sarlogic_0/net67 0 1.662327f
C1375 sarlogic_0/_444_/a_2560_156# 0 0.016968f
C1376 sarlogic_0/_444_/a_2665_112# 0 0.62251f
C1377 sarlogic_0/_444_/a_2248_156# 0 0.371662f
C1378 sarlogic_0/_444_/a_1204_472# 0 0.012971f
C1379 sarlogic_0/_444_/a_1000_472# 0 0.291735f
C1380 sarlogic_0/_444_/a_796_472# 0 0.023206f
C1381 sarlogic_0/_444_/a_1308_423# 0 0.279043f
C1382 sarlogic_0/_444_/a_448_472# 0 0.684413f
C1383 sarlogic_0/_444_/a_36_151# 0 1.43589f
C1384 sarlogic_0/net65 0 0.804072f
C1385 sarlogic_0/fanout57/a_36_113# 0 0.418095f
C1386 sarlogic_0/fanout68/a_36_113# 0 0.418095f
C1387 sarlogic_0/FILLER_0_12_2/a_484_472# 0 0.345058f
C1388 sarlogic_0/FILLER_0_12_2/a_36_472# 0 0.404746f
C1389 sarlogic_0/FILLER_0_12_2/a_572_375# 0 0.232991f
C1390 sarlogic_0/FILLER_0_12_2/a_124_375# 0 0.185089f
C1391 sarlogic_0/net79 0 1.584979f
C1392 sarlogic_0/fanout79/a_36_160# 0 0.386641f
C1393 sarlogic_0/_392_/a_36_68# 0 0.112263f
C1394 sarlogic_0/FILLER_0_13_228/a_36_472# 0 0.417394f
C1395 sarlogic_0/FILLER_0_13_228/a_124_375# 0 0.246306f
C1396 sarlogic_0/FILLER_0_13_206/a_36_472# 0 0.417394f
C1397 sarlogic_0/FILLER_0_13_206/a_124_375# 0 0.246306f
C1398 sarlogic_0/FILLER_0_20_177/a_1380_472# 0 0.345058f
C1399 sarlogic_0/FILLER_0_20_177/a_932_472# 0 0.33241f
C1400 sarlogic_0/FILLER_0_20_177/a_484_472# 0 0.33241f
C1401 sarlogic_0/FILLER_0_20_177/a_36_472# 0 0.404746f
C1402 sarlogic_0/FILLER_0_20_177/a_1468_375# 0 0.233029f
C1403 sarlogic_0/FILLER_0_20_177/a_1020_375# 0 0.171606f
C1404 sarlogic_0/FILLER_0_20_177/a_572_375# 0 0.171606f
C1405 sarlogic_0/FILLER_0_20_177/a_124_375# 0 0.185399f
C1406 sarlogic_0/_051_ 0 0.349381f
C1407 sarlogic_0/_213_/a_67_603# 0 0.345683f
C1408 sarlogic_0/net2 0 0.461658f
C1409 sarlogic_0/input2/a_36_113# 0 0.418095f
C1410 sarlogic_0/_129_ 0 0.926508f
C1411 sarlogic_0/_131_ 0 1.734297f
C1412 sarlogic_0/_359_/a_36_488# 0 0.101145f
C1413 sarlogic_0/FILLER_0_11_64/a_36_472# 0 0.417394f
C1414 sarlogic_0/FILLER_0_11_64/a_124_375# 0 0.246306f
C1415 sarlogic_0/state\[2\] 0 0.607433f
C1416 sarlogic_0/net53 0 4.483899f
C1417 sarlogic_0/_017_ 0 0.334329f
C1418 sarlogic_0/net70 0 1.238296f
C1419 sarlogic_0/_428_/a_2560_156# 0 0.016968f
C1420 sarlogic_0/_428_/a_2665_112# 0 0.62251f
C1421 sarlogic_0/_428_/a_2248_156# 0 0.371662f
C1422 sarlogic_0/_428_/a_1204_472# 0 0.012971f
C1423 sarlogic_0/_428_/a_1000_472# 0 0.291735f
C1424 sarlogic_0/_428_/a_796_472# 0 0.023206f
C1425 sarlogic_0/_428_/a_1308_423# 0 0.279043f
C1426 sarlogic_0/_428_/a_448_472# 0 0.684413f
C1427 sarlogic_0/_428_/a_36_151# 0 1.43589f
C1428 sarlogic_0/FILLER_0_5_72/a_1380_472# 0 0.345058f
C1429 sarlogic_0/FILLER_0_5_72/a_932_472# 0 0.33241f
C1430 sarlogic_0/FILLER_0_5_72/a_484_472# 0 0.33241f
C1431 sarlogic_0/FILLER_0_5_72/a_36_472# 0 0.404746f
C1432 sarlogic_0/FILLER_0_5_72/a_1468_375# 0 0.233029f
C1433 sarlogic_0/FILLER_0_5_72/a_1020_375# 0 0.171606f
C1434 sarlogic_0/FILLER_0_5_72/a_572_375# 0 0.171606f
C1435 sarlogic_0/FILLER_0_5_72/a_124_375# 0 0.185399f
C1436 sarlogic_0/_376_/a_36_160# 0 0.386641f
C1437 sarlogic_0/trim_val\[1\] 0 0.683578f
C1438 sarlogic_0/_445_/a_2560_156# 0 0.016968f
C1439 sarlogic_0/_445_/a_2665_112# 0 0.62251f
C1440 sarlogic_0/_445_/a_2248_156# 0 0.371662f
C1441 sarlogic_0/_445_/a_1204_472# 0 0.012971f
C1442 sarlogic_0/_445_/a_1000_472# 0 0.291735f
C1443 sarlogic_0/_445_/a_796_472# 0 0.023206f
C1444 sarlogic_0/_445_/a_1308_423# 0 0.279043f
C1445 sarlogic_0/_445_/a_448_472# 0 0.684413f
C1446 sarlogic_0/_445_/a_36_151# 0 1.43589f
C1447 sarlogic_0/fanout67/a_36_160# 0 0.386641f
C1448 sarlogic_0/fanout56/a_36_113# 0 0.418095f
C1449 sarlogic_0/net78 0 0.686263f
C1450 sarlogic_0/fanout78/a_36_113# 0 0.418095f
C1451 sarlogic_0/_174_ 0 0.979741f
C1452 sarlogic_0/FILLER_0_0_198/a_36_472# 0 0.417394f
C1453 sarlogic_0/FILLER_0_0_198/a_124_375# 0 0.246306f
C1454 sarlogic_0/FILLER_0_15_290/a_36_472# 0 0.417394f
C1455 sarlogic_0/FILLER_0_15_290/a_124_375# 0 0.246306f
C1456 sarlogic_0/FILLER_0_24_290/a_36_472# 0 0.417394f
C1457 sarlogic_0/FILLER_0_24_290/a_124_375# 0 0.246306f
C1458 sarlogic_0/FILLER_0_4_107/a_1380_472# 0 0.345058f
C1459 sarlogic_0/FILLER_0_4_107/a_932_472# 0 0.33241f
C1460 sarlogic_0/FILLER_0_4_107/a_484_472# 0 0.33241f
C1461 sarlogic_0/FILLER_0_4_107/a_36_472# 0 0.404746f
C1462 sarlogic_0/FILLER_0_4_107/a_1468_375# 0 0.233029f
C1463 sarlogic_0/FILLER_0_4_107/a_1020_375# 0 0.171606f
C1464 sarlogic_0/FILLER_0_4_107/a_572_375# 0 0.171606f
C1465 sarlogic_0/FILLER_0_4_107/a_124_375# 0 0.185399f
C1466 sarlogic_0/FILLER_0_7_104/a_1380_472# 0 0.345058f
C1467 sarlogic_0/FILLER_0_7_104/a_932_472# 0 0.33241f
C1468 sarlogic_0/FILLER_0_7_104/a_484_472# 0 0.33241f
C1469 sarlogic_0/FILLER_0_7_104/a_36_472# 0 0.404746f
C1470 sarlogic_0/FILLER_0_7_104/a_1468_375# 0 0.233029f
C1471 sarlogic_0/FILLER_0_7_104/a_1020_375# 0 0.171606f
C1472 sarlogic_0/FILLER_0_7_104/a_572_375# 0 0.171606f
C1473 sarlogic_0/FILLER_0_7_104/a_124_375# 0 0.185399f
C1474 sarlogic_0/_214_/a_36_160# 0 0.386641f
C1475 sarlogic_0/net1 0 0.364811f
C1476 sarlogic_0/input1/a_36_113# 0 0.418095f
C1477 sarlogic_0/_429_/a_2560_156# 0 0.016968f
C1478 sarlogic_0/_429_/a_2665_112# 0 0.62251f
C1479 sarlogic_0/_429_/a_2248_156# 0 0.371662f
C1480 sarlogic_0/_429_/a_1204_472# 0 0.012971f
C1481 sarlogic_0/_429_/a_1000_472# 0 0.291735f
C1482 sarlogic_0/_429_/a_796_472# 0 0.023206f
C1483 sarlogic_0/_429_/a_1308_423# 0 0.279043f
C1484 sarlogic_0/_429_/a_448_472# 0 0.684413f
C1485 sarlogic_0/_429_/a_36_151# 0 1.43589f
C1486 sarlogic_0/_011_ 0 0.278979f
C1487 sarlogic_0/_377_/a_36_472# 0 0.031137f
C1488 sarlogic_0/fanout66/a_36_113# 0 0.418095f
C1489 sarlogic_0/_035_ 0 0.327801f
C1490 sarlogic_0/_446_/a_2560_156# 0 0.016968f
C1491 sarlogic_0/_446_/a_2665_112# 0 0.62251f
C1492 sarlogic_0/_446_/a_2248_156# 0 0.371662f
C1493 sarlogic_0/_446_/a_1204_472# 0 0.012971f
C1494 sarlogic_0/_446_/a_1000_472# 0 0.291735f
C1495 sarlogic_0/_446_/a_796_472# 0 0.023206f
C1496 sarlogic_0/_446_/a_1308_423# 0 0.279043f
C1497 sarlogic_0/_446_/a_448_472# 0 0.684413f
C1498 sarlogic_0/_446_/a_36_151# 0 1.43589f
C1499 sarlogic_0/fanout77/a_36_113# 0 0.418095f
C1500 sarlogic_0/FILLER_0_5_212/a_36_472# 0 0.417394f
C1501 sarlogic_0/FILLER_0_5_212/a_124_375# 0 0.246306f
C1502 sarlogic_0/fanout55/a_36_160# 0 0.696445f
C1503 sarlogic_0/_175_ 0 0.344159f
C1504 sarlogic_0/_394_/a_1936_472# 0 0.009918f
C1505 sarlogic_0/_394_/a_718_524# 0 0.005143f
C1506 sarlogic_0/_394_/a_56_524# 0 0.41096f
C1507 sarlogic_0/_394_/a_728_93# 0 0.654825f
C1508 sarlogic_0/_394_/a_1336_472# 0 0.316639f
C1509 sarlogic_0/FILLER_0_3_172/a_3172_472# 0 0.345058f
C1510 sarlogic_0/FILLER_0_3_172/a_2724_472# 0 0.33241f
C1511 sarlogic_0/FILLER_0_3_172/a_2276_472# 0 0.33241f
C1512 sarlogic_0/FILLER_0_3_172/a_1828_472# 0 0.33241f
C1513 sarlogic_0/FILLER_0_3_172/a_1380_472# 0 0.33241f
C1514 sarlogic_0/FILLER_0_3_172/a_932_472# 0 0.33241f
C1515 sarlogic_0/FILLER_0_3_172/a_484_472# 0 0.33241f
C1516 sarlogic_0/FILLER_0_3_172/a_36_472# 0 0.404746f
C1517 sarlogic_0/FILLER_0_3_172/a_3260_375# 0 0.233093f
C1518 sarlogic_0/FILLER_0_3_172/a_2812_375# 0 0.17167f
C1519 sarlogic_0/FILLER_0_3_172/a_2364_375# 0 0.17167f
C1520 sarlogic_0/FILLER_0_3_172/a_1916_375# 0 0.17167f
C1521 sarlogic_0/FILLER_0_3_172/a_1468_375# 0 0.17167f
C1522 sarlogic_0/FILLER_0_3_172/a_1020_375# 0 0.17167f
C1523 sarlogic_0/FILLER_0_3_172/a_572_375# 0 0.17167f
C1524 sarlogic_0/FILLER_0_3_172/a_124_375# 0 0.185915f
C1525 sarlogic_0/FILLER_0_17_72/a_3172_472# 0 0.345058f
C1526 sarlogic_0/FILLER_0_17_72/a_2724_472# 0 0.33241f
C1527 sarlogic_0/FILLER_0_17_72/a_2276_472# 0 0.33241f
C1528 sarlogic_0/FILLER_0_17_72/a_1828_472# 0 0.33241f
C1529 sarlogic_0/FILLER_0_17_72/a_1380_472# 0 0.33241f
C1530 sarlogic_0/FILLER_0_17_72/a_932_472# 0 0.33241f
C1531 sarlogic_0/FILLER_0_17_72/a_484_472# 0 0.33241f
C1532 sarlogic_0/FILLER_0_17_72/a_36_472# 0 0.404746f
C1533 sarlogic_0/FILLER_0_17_72/a_3260_375# 0 0.233093f
C1534 sarlogic_0/FILLER_0_17_72/a_2812_375# 0 0.17167f
C1535 sarlogic_0/FILLER_0_17_72/a_2364_375# 0 0.17167f
C1536 sarlogic_0/FILLER_0_17_72/a_1916_375# 0 0.17167f
C1537 sarlogic_0/FILLER_0_17_72/a_1468_375# 0 0.17167f
C1538 sarlogic_0/FILLER_0_17_72/a_1020_375# 0 0.17167f
C1539 sarlogic_0/FILLER_0_17_72/a_572_375# 0 0.17167f
C1540 sarlogic_0/FILLER_0_17_72/a_124_375# 0 0.185915f
C1541 sarlogic_0/FILLER_0_2_93/a_484_472# 0 0.345058f
C1542 sarlogic_0/FILLER_0_2_93/a_36_472# 0 0.404746f
C1543 sarlogic_0/FILLER_0_2_93/a_572_375# 0 0.232991f
C1544 sarlogic_0/FILLER_0_2_93/a_124_375# 0 0.185089f
C1545 sarlogic_0/FILLER_0_11_142/a_484_472# 0 0.345058f
C1546 sarlogic_0/FILLER_0_11_142/a_36_472# 0 0.404746f
C1547 sarlogic_0/FILLER_0_11_142/a_572_375# 0 0.232991f
C1548 sarlogic_0/FILLER_0_11_142/a_124_375# 0 0.185089f
C1549 sarlogic_0/net25 0 1.803174f
C1550 sarlogic_0/_232_/a_67_603# 0 0.345683f
C1551 sarlogic_0/net35 0 1.844415f
C1552 sarlogic_0/mask\[8\] 0 1.276111f
C1553 sarlogic_0/_301_/a_36_472# 0 0.031137f
C1554 sarlogic_0/_033_ 0 0.323682f
C1555 sarlogic_0/_165_ 0 0.331995f
C1556 sarlogic_0/FILLER_0_3_2/a_36_472# 0 0.417394f
C1557 sarlogic_0/FILLER_0_3_2/a_124_375# 0 0.246306f
C1558 sarlogic_0/trim_val\[3\] 0 0.719615f
C1559 sarlogic_0/_036_ 0 0.369206f
C1560 sarlogic_0/net68 0 1.735004f
C1561 sarlogic_0/_447_/a_2560_156# 0 0.016968f
C1562 sarlogic_0/_447_/a_2665_112# 0 0.62251f
C1563 sarlogic_0/_447_/a_2248_156# 0 0.371662f
C1564 sarlogic_0/_447_/a_1204_472# 0 0.012971f
C1565 sarlogic_0/_447_/a_1000_472# 0 0.291735f
C1566 sarlogic_0/_447_/a_796_472# 0 0.023206f
C1567 sarlogic_0/_447_/a_1308_423# 0 0.279043f
C1568 sarlogic_0/_447_/a_448_472# 0 0.684413f
C1569 sarlogic_0/_447_/a_36_151# 0 1.43589f
C1570 sarlogic_0/FILLER_0_19_28/a_484_472# 0 0.345058f
C1571 sarlogic_0/FILLER_0_19_28/a_36_472# 0 0.404746f
C1572 sarlogic_0/FILLER_0_19_28/a_572_375# 0 0.232991f
C1573 sarlogic_0/FILLER_0_19_28/a_124_375# 0 0.185089f
C1574 sarlogic_0/fanout65/a_36_113# 0 0.418095f
C1575 sarlogic_0/fanout76/a_36_160# 0 0.386641f
C1576 sarlogic_0/net54 0 5.456963f
C1577 sarlogic_0/fanout54/a_36_160# 0 0.696445f
C1578 sarlogic_0/FILLER_0_4_49/a_484_472# 0 0.345058f
C1579 sarlogic_0/FILLER_0_4_49/a_36_472# 0 0.404746f
C1580 sarlogic_0/FILLER_0_4_49/a_572_375# 0 0.232991f
C1581 sarlogic_0/FILLER_0_4_49/a_124_375# 0 0.185089f
C1582 sarlogic_0/_176_ 0 0.804011f
C1583 sarlogic_0/_085_ 0 2.280803f
C1584 sarlogic_0/_116_ 0 1.959915f
C1585 sarlogic_0/_395_/a_36_488# 0 0.101145f
C1586 sarlogic_0/FILLER_0_14_50/a_36_472# 0 0.417394f
C1587 sarlogic_0/FILLER_0_14_50/a_124_375# 0 0.246306f
C1588 sarlogic_0/FILLER_0_8_263/a_36_472# 0 0.417394f
C1589 sarlogic_0/FILLER_0_8_263/a_124_375# 0 0.246306f
C1590 sarlogic_0/FILLER_0_0_130/a_36_472# 0 0.417394f
C1591 sarlogic_0/FILLER_0_0_130/a_124_375# 0 0.246306f
C1592 sarlogic_0/FILLER_0_16_255/a_36_472# 0 0.417394f
C1593 sarlogic_0/FILLER_0_16_255/a_124_375# 0 0.246306f
C1594 sarlogic_0/FILLER_0_7_59/a_484_472# 0 0.345058f
C1595 sarlogic_0/FILLER_0_7_59/a_36_472# 0 0.404746f
C1596 sarlogic_0/FILLER_0_7_59/a_572_375# 0 0.232991f
C1597 sarlogic_0/FILLER_0_7_59/a_124_375# 0 0.185089f
C1598 sarlogic_0/output19/a_224_472# 0 2.38465f
C1599 sarlogic_0/FILLER_0_7_146/a_36_472# 0 0.417394f
C1600 sarlogic_0/FILLER_0_7_146/a_124_375# 0 0.246306f
C1601 sarlogic_0/_216_/a_67_603# 0 0.345683f
C1602 sarlogic_0/FILLER_0_15_116/a_484_472# 0 0.345058f
C1603 sarlogic_0/FILLER_0_15_116/a_36_472# 0 0.404746f
C1604 sarlogic_0/FILLER_0_15_116/a_572_375# 0 0.232991f
C1605 sarlogic_0/FILLER_0_15_116/a_124_375# 0 0.185089f
C1606 sarlogic_0/_063_ 0 0.370155f
C1607 sarlogic_0/_233_/a_36_160# 0 0.386641f
C1608 sarlogic_0/FILLER_0_21_28/a_3172_472# 0 0.345058f
C1609 sarlogic_0/FILLER_0_21_28/a_2724_472# 0 0.33241f
C1610 sarlogic_0/FILLER_0_21_28/a_2276_472# 0 0.33241f
C1611 sarlogic_0/FILLER_0_21_28/a_1828_472# 0 0.33241f
C1612 sarlogic_0/FILLER_0_21_28/a_1380_472# 0 0.33241f
C1613 sarlogic_0/FILLER_0_21_28/a_932_472# 0 0.33241f
C1614 sarlogic_0/FILLER_0_21_28/a_484_472# 0 0.33241f
C1615 sarlogic_0/FILLER_0_21_28/a_36_472# 0 0.404746f
C1616 sarlogic_0/FILLER_0_21_28/a_3260_375# 0 0.233093f
C1617 sarlogic_0/FILLER_0_21_28/a_2812_375# 0 0.17167f
C1618 sarlogic_0/FILLER_0_21_28/a_2364_375# 0 0.17167f
C1619 sarlogic_0/FILLER_0_21_28/a_1916_375# 0 0.17167f
C1620 sarlogic_0/FILLER_0_21_28/a_1468_375# 0 0.17167f
C1621 sarlogic_0/FILLER_0_21_28/a_1020_375# 0 0.17167f
C1622 sarlogic_0/FILLER_0_21_28/a_572_375# 0 0.17167f
C1623 sarlogic_0/FILLER_0_21_28/a_124_375# 0 0.185915f
C1624 sarlogic_0/_110_ 0 0.323912f
C1625 sarlogic_0/_379_/a_36_472# 0 0.031137f
C1626 sarlogic_0/trim_val\[4\] 0 0.662409f
C1627 sarlogic_0/net76 0 1.454269f
C1628 sarlogic_0/_448_/a_2560_156# 0 0.016968f
C1629 sarlogic_0/_448_/a_2665_112# 0 0.62251f
C1630 sarlogic_0/_448_/a_2248_156# 0 0.371662f
C1631 sarlogic_0/_448_/a_1204_472# 0 0.012971f
C1632 sarlogic_0/_448_/a_1000_472# 0 0.291735f
C1633 sarlogic_0/_448_/a_796_472# 0 0.023206f
C1634 sarlogic_0/_448_/a_1308_423# 0 0.279043f
C1635 sarlogic_0/_448_/a_448_472# 0 0.684413f
C1636 sarlogic_0/_448_/a_36_151# 0 1.43589f
C1637 sarlogic_0/fanout64/a_36_160# 0 0.386641f
C1638 sarlogic_0/fanout75/a_36_113# 0 0.418095f
C1639 sarlogic_0/_250_/a_36_68# 0 0.69549f
C1640 sarlogic_0/net56 0 0.843396f
C1641 sarlogic_0/fanout53/a_36_160# 0 0.696445f
C1642 sarlogic_0/_177_ 0 0.358286f
C1643 result[2] 0 16.5685f
C1644 sarlogic_0/net29 0 1.802718f
C1645 sarlogic_0/output29/a_224_472# 0 2.38465f
C1646 sarlogic_0/output18/a_224_472# 0 2.38465f
C1647 sarlogic_0/FILLER_0_14_181/a_36_472# 0 0.417394f
C1648 sarlogic_0/FILLER_0_14_181/a_124_375# 0 0.246306f
C1649 sarlogic_0/_052_ 0 0.569133f
C1650 sarlogic_0/_217_/a_36_160# 0 0.386641f
C1651 sarlogic_0/net44 0 1.407054f
C1652 sarlogic_0/_303_/a_36_472# 0 0.031137f
C1653 sarlogic_0/en_co_clk 0 0.346872f
C1654 sarlogic_0/net55 0 5.119958f
C1655 sarlogic_0/net72 0 1.366255f
C1656 sarlogic_0/_449_/a_2560_156# 0 0.016968f
C1657 sarlogic_0/_449_/a_2665_112# 0 0.62251f
C1658 sarlogic_0/_449_/a_2248_156# 0 0.371662f
C1659 sarlogic_0/_449_/a_1204_472# 0 0.012971f
C1660 sarlogic_0/_449_/a_1000_472# 0 0.291735f
C1661 sarlogic_0/_449_/a_796_472# 0 0.023206f
C1662 sarlogic_0/_449_/a_1308_423# 0 0.279043f
C1663 sarlogic_0/_449_/a_448_472# 0 0.684413f
C1664 sarlogic_0/_449_/a_36_151# 0 1.43589f
C1665 sarlogic_0/fanout52/a_36_160# 0 0.696445f
C1666 sarlogic_0/net82 0 0.706042f
C1667 sarlogic_0/fanout74/a_36_113# 0 0.418095f
C1668 sarlogic_0/FILLER_0_10_28/a_36_472# 0 0.417394f
C1669 sarlogic_0/FILLER_0_10_28/a_124_375# 0 0.246306f
C1670 sarlogic_0/mask\[0\] 0 2.242948f
C1671 sarlogic_0/_320_/a_36_472# 0 0.137725f
C1672 sarlogic_0/fanout63/a_36_160# 0 0.696445f
C1673 sarlogic_0/FILLER_0_14_81/a_36_472# 0 0.417394f
C1674 sarlogic_0/FILLER_0_14_81/a_124_375# 0 0.246306f
C1675 sarlogic_0/_397_/a_36_472# 0 0.031137f
C1676 sarlogic_0/FILLER_0_13_212/a_1380_472# 0 0.345058f
C1677 sarlogic_0/FILLER_0_13_212/a_932_472# 0 0.33241f
C1678 sarlogic_0/FILLER_0_13_212/a_484_472# 0 0.33241f
C1679 sarlogic_0/FILLER_0_13_212/a_36_472# 0 0.404746f
C1680 sarlogic_0/FILLER_0_13_212/a_1468_375# 0 0.233029f
C1681 sarlogic_0/FILLER_0_13_212/a_1020_375# 0 0.171606f
C1682 sarlogic_0/FILLER_0_13_212/a_572_375# 0 0.171606f
C1683 sarlogic_0/FILLER_0_13_212/a_124_375# 0 0.185399f
C1684 sarlogic_0/net39 0 1.445128f
C1685 sarlogic_0/output39/a_224_472# 0 2.38465f
C1686 result[1] 0 16.567158f
C1687 sarlogic_0/net28 0 1.759728f
C1688 sarlogic_0/output28/a_224_472# 0 2.38465f
C1689 sarlogic_0/output17/a_224_472# 0 2.38465f
C1690 sarlogic_0/FILLER_0_16_37/a_36_472# 0 0.417394f
C1691 sarlogic_0/FILLER_0_16_37/a_124_375# 0 0.246306f
C1692 sarlogic_0/net26 0 1.671545f
C1693 sarlogic_0/_064_ 0 0.581481f
C1694 sarlogic_0/trim_val\[2\] 0 0.65354f
C1695 sarlogic_0/trim_mask\[2\] 0 0.92551f
C1696 sarlogic_0/_235_/a_67_603# 0 0.345683f
C1697 sarlogic_0/_013_ 0 0.48783f
C1698 sarlogic_0/_111_ 0 0.369652f
C1699 sarlogic_0/FILLER_0_18_177/a_3172_472# 0 0.345058f
C1700 sarlogic_0/FILLER_0_18_177/a_2724_472# 0 0.33241f
C1701 sarlogic_0/FILLER_0_18_177/a_2276_472# 0 0.33241f
C1702 sarlogic_0/FILLER_0_18_177/a_1828_472# 0 0.33241f
C1703 sarlogic_0/FILLER_0_18_177/a_1380_472# 0 0.33241f
C1704 sarlogic_0/FILLER_0_18_177/a_932_472# 0 0.33241f
C1705 sarlogic_0/FILLER_0_18_177/a_484_472# 0 0.33241f
C1706 sarlogic_0/FILLER_0_18_177/a_36_472# 0 0.404746f
C1707 sarlogic_0/FILLER_0_18_177/a_3260_375# 0 0.233093f
C1708 sarlogic_0/FILLER_0_18_177/a_2812_375# 0 0.17167f
C1709 sarlogic_0/FILLER_0_18_177/a_2364_375# 0 0.17167f
C1710 sarlogic_0/FILLER_0_18_177/a_1916_375# 0 0.17167f
C1711 sarlogic_0/FILLER_0_18_177/a_1468_375# 0 0.17167f
C1712 sarlogic_0/FILLER_0_18_177/a_1020_375# 0 0.17167f
C1713 sarlogic_0/FILLER_0_18_177/a_572_375# 0 0.17167f
C1714 sarlogic_0/FILLER_0_18_177/a_124_375# 0 0.185915f
C1715 sarlogic_0/FILLER_0_18_100/a_36_472# 0 0.417394f
C1716 sarlogic_0/FILLER_0_18_100/a_124_375# 0 0.246306f
C1717 sarlogic_0/_073_ 0 0.953711f
C1718 sarlogic_0/_126_ 0 2.036767f
C1719 sarlogic_0/_069_ 0 2.034557f
C1720 sarlogic_0/_321_/a_170_472# 0 0.077257f
C1721 sarlogic_0/fanout51/a_36_113# 0 0.418095f
C1722 sarlogic_0/net62 0 4.932099f
C1723 sarlogic_0/fanout62/a_36_160# 0 0.696445f
C1724 sarlogic_0/fanout73/a_36_113# 0 0.418095f
C1725 sarlogic_0/FILLER_0_19_47/a_484_472# 0 0.345058f
C1726 sarlogic_0/FILLER_0_19_47/a_36_472# 0 0.404746f
C1727 sarlogic_0/FILLER_0_19_47/a_572_375# 0 0.232991f
C1728 sarlogic_0/FILLER_0_19_47/a_124_375# 0 0.185089f
C1729 sarlogic_0/FILLER_0_14_91/a_484_472# 0 0.345058f
C1730 sarlogic_0/FILLER_0_14_91/a_36_472# 0 0.404746f
C1731 sarlogic_0/FILLER_0_14_91/a_572_375# 0 0.232991f
C1732 sarlogic_0/FILLER_0_14_91/a_124_375# 0 0.185089f
C1733 sarlogic_0/FILLER_0_10_214/a_36_472# 0 0.417394f
C1734 sarlogic_0/FILLER_0_10_214/a_124_375# 0 0.246306f
C1735 sarlogic_0/FILLER_0_10_247/a_36_472# 0 0.417394f
C1736 sarlogic_0/FILLER_0_10_247/a_124_375# 0 0.246306f
C1737 sarlogic_0/_178_ 0 1.252435f
C1738 sarlogic_0/_398_/a_36_113# 0 0.418095f
C1739 sarlogic_0/FILLER_0_16_241/a_36_472# 0 0.417394f
C1740 sarlogic_0/FILLER_0_16_241/a_124_375# 0 0.246306f
C1741 sarlogic_0/net38 0 1.529392f
C1742 sarlogic_0/output38/a_224_472# 0 2.38465f
C1743 sarlogic_0/net16 0 1.295744f
C1744 sarlogic_0/output16/a_224_472# 0 2.38465f
C1745 result[0] 0 21.268515f
C1746 sarlogic_0/output27/a_224_472# 0 2.38465f
C1747 sarlogic_0/_219_/a_36_160# 0 0.386641f
C1748 sarlogic_0/FILLER_0_20_193/a_484_472# 0 0.345058f
C1749 sarlogic_0/FILLER_0_20_193/a_36_472# 0 0.404746f
C1750 sarlogic_0/FILLER_0_20_193/a_572_375# 0 0.232991f
C1751 sarlogic_0/FILLER_0_20_193/a_124_375# 0 0.185089f
C1752 sarlogic_0/_236_/a_36_160# 0 0.696445f
C1753 sarlogic_0/_112_ 0 0.308886f
C1754 sarlogic_0/_305_/a_36_159# 0 0.374116f
C1755 sarlogic_0/_074_ 0 1.813232f
C1756 sarlogic_0/_253_/a_36_68# 0 0.061249f
C1757 sarlogic_0/net50 0 4.486121f
C1758 sarlogic_0/net52 0 3.536016f
C1759 sarlogic_0/fanout50/a_36_160# 0 0.696445f
C1760 sarlogic_0/FILLER_0_10_37/a_36_472# 0 0.417394f
C1761 sarlogic_0/FILLER_0_10_37/a_124_375# 0 0.246306f
C1762 sarlogic_0/fanout72/a_36_113# 0 0.418095f
C1763 sarlogic_0/fanout61/a_36_113# 0 0.418095f
C1764 sarlogic_0/_128_ 0 0.447252f
C1765 sarlogic_0/_127_ 0 1.291729f
C1766 sarlogic_0/_322_/a_848_380# 0 0.40208f
C1767 sarlogic_0/_322_/a_124_24# 0 0.591898f
C1768 sarlogic_0/_088_ 0 0.457961f
C1769 sarlogic_0/_079_ 0 1.114894f
C1770 sarlogic_0/_087_ 0 0.601674f
C1771 sarlogic_0/_270_/a_36_472# 0 0.031137f
C1772 sarlogic_0/FILLER_0_4_123/a_36_472# 0 0.417394f
C1773 sarlogic_0/FILLER_0_4_123/a_124_375# 0 0.246306f
C1774 sarlogic_0/FILLER_0_17_218/a_484_472# 0 0.345058f
C1775 sarlogic_0/FILLER_0_17_218/a_36_472# 0 0.404746f
C1776 sarlogic_0/FILLER_0_17_218/a_572_375# 0 0.232991f
C1777 sarlogic_0/FILLER_0_17_218/a_124_375# 0 0.185089f
C1778 sarlogic_0/output37/a_224_472# 0 2.38465f
C1779 valid 0 20.974365f
C1780 sarlogic_0/net48 0 1.219262f
C1781 sarlogic_0/output48/a_224_472# 0 2.38465f
C1782 sarlogic_0/net15 0 1.440851f
C1783 sarlogic_0/output15/a_224_472# 0 2.38465f
C1784 sarlogic_0/output26/a_224_472# 0 2.38465f
C1785 sarlogic_0/FILLER_0_16_57/a_1380_472# 0 0.345058f
C1786 sarlogic_0/FILLER_0_16_57/a_932_472# 0 0.33241f
C1787 sarlogic_0/FILLER_0_16_57/a_484_472# 0 0.33241f
C1788 sarlogic_0/FILLER_0_16_57/a_36_472# 0 0.404746f
C1789 sarlogic_0/FILLER_0_16_57/a_1468_375# 0 0.233029f
C1790 sarlogic_0/FILLER_0_16_57/a_1020_375# 0 0.171606f
C1791 sarlogic_0/FILLER_0_16_57/a_572_375# 0 0.171606f
C1792 sarlogic_0/FILLER_0_16_57/a_124_375# 0 0.185399f
C1793 sarlogic_0/_306_/a_36_68# 0 0.69549f
C1794 sarlogic_0/_072_ 0 2.604301f
C1795 sarlogic_0/fanout82/a_36_113# 0 0.418095f
C1796 sarlogic_0/_015_ 0 0.406653f
C1797 sarlogic_0/_323_/a_36_113# 0 0.418095f
C1798 sarlogic_0/net60 0 5.024503f
C1799 sarlogic_0/net61 0 1.666523f
C1800 sarlogic_0/fanout60/a_36_160# 0 0.696445f
C1801 sarlogic_0/fanout71/a_36_113# 0 0.418095f
C1802 sarlogic_0/FILLER_0_6_239/a_36_472# 0 0.417394f
C1803 sarlogic_0/FILLER_0_6_239/a_124_375# 0 0.246306f
C1804 sarlogic_0/FILLER_0_4_99/a_36_472# 0 0.417394f
C1805 sarlogic_0/FILLER_0_4_99/a_124_375# 0 0.246306f
C1806 sarlogic_0/net57 0 1.383718f
C1807 sarlogic_0/FILLER_0_10_256/a_36_472# 0 0.417394f
C1808 sarlogic_0/FILLER_0_10_256/a_124_375# 0 0.246306f
C1809 sarlogic_0/cal_itt\[3\] 0 1.854962f
C1810 sarlogic_0/_340_/a_36_160# 0 0.386641f
C1811 sarlogic_0/FILLER_0_4_177/a_484_472# 0 0.345058f
C1812 sarlogic_0/FILLER_0_4_177/a_36_472# 0 0.404746f
C1813 sarlogic_0/FILLER_0_4_177/a_572_375# 0 0.232991f
C1814 sarlogic_0/FILLER_0_4_177/a_124_375# 0 0.185089f
C1815 sarlogic_0/FILLER_0_4_144/a_484_472# 0 0.345058f
C1816 sarlogic_0/FILLER_0_4_144/a_36_472# 0 0.404746f
C1817 sarlogic_0/FILLER_0_4_144/a_572_375# 0 0.232991f
C1818 sarlogic_0/FILLER_0_4_144/a_124_375# 0 0.185089f
C1819 sarlogic_0/output14/a_224_472# 0 2.38465f
C1820 result[9] 0 21.520042f
C1821 sarlogic_0/output36/a_224_472# 0 2.38465f
C1822 sarlogic_0/output47/a_224_472# 0 2.38465f
C1823 sarlogic_0/output25/a_224_472# 0 2.38465f
C1824 sarlogic_0/FILLER_0_12_136/a_1380_472# 0 0.345058f
C1825 sarlogic_0/FILLER_0_12_136/a_932_472# 0 0.33241f
C1826 sarlogic_0/FILLER_0_12_136/a_484_472# 0 0.33241f
C1827 sarlogic_0/FILLER_0_12_136/a_36_472# 0 0.404746f
C1828 sarlogic_0/FILLER_0_12_136/a_1468_375# 0 0.233029f
C1829 sarlogic_0/FILLER_0_12_136/a_1020_375# 0 0.171606f
C1830 sarlogic_0/FILLER_0_12_136/a_572_375# 0 0.171606f
C1831 sarlogic_0/FILLER_0_12_136/a_124_375# 0 0.185399f
C1832 sarlogic_0/FILLER_0_16_89/a_1380_472# 0 0.345058f
C1833 sarlogic_0/FILLER_0_16_89/a_932_472# 0 0.33241f
C1834 sarlogic_0/FILLER_0_16_89/a_484_472# 0 0.33241f
C1835 sarlogic_0/FILLER_0_16_89/a_36_472# 0 0.404746f
C1836 sarlogic_0/FILLER_0_16_89/a_1468_375# 0 0.233029f
C1837 sarlogic_0/FILLER_0_16_89/a_1020_375# 0 0.171606f
C1838 sarlogic_0/FILLER_0_16_89/a_572_375# 0 0.171606f
C1839 sarlogic_0/FILLER_0_16_89/a_124_375# 0 0.185399f
C1840 sarlogic_0/FILLER_0_21_125/a_484_472# 0 0.345058f
C1841 sarlogic_0/FILLER_0_21_125/a_36_472# 0 0.404746f
C1842 sarlogic_0/FILLER_0_21_125/a_572_375# 0 0.232991f
C1843 sarlogic_0/FILLER_0_21_125/a_124_375# 0 0.185089f
C1844 sarlogic_0/_238_/a_67_603# 0 0.345683f
C1845 sarlogic_0/_096_ 0 2.205532f
C1846 sarlogic_0/_093_ 0 1.893313f
C1847 sarlogic_0/FILLER_0_19_55/a_36_472# 0 0.417394f
C1848 sarlogic_0/FILLER_0_19_55/a_124_375# 0 0.246306f
C1849 sarlogic_0/net81 0 1.738987f
C1850 sarlogic_0/fanout81/a_36_160# 0 0.386641f
C1851 sarlogic_0/_057_ 0 1.600886f
C1852 sarlogic_0/_255_/a_224_552# 0 1.31114f
C1853 sarlogic_0/net73 0 1.058857f
C1854 sarlogic_0/fanout70/a_36_113# 0 0.418095f
C1855 sarlogic_0/_003_ 0 0.3064f
C1856 sarlogic_0/_089_ 0 0.36777f
C1857 sarlogic_0/_272_/a_36_472# 0 0.031137f
C1858 sarlogic_0/_187_ 0 0.311229f
C1859 sarlogic_0/_410_/a_36_68# 0 0.112263f
C1860 sarlogic_0/_141_ 0 1.249289f
C1861 sarlogic_0/mask\[3\] 0 1.26722f
C1862 sarlogic_0/_341_/a_49_472# 0 0.054843f
C1863 cal 0 17.131042f
C1864 sarlogic_0/FILLER_0_7_195/a_36_472# 0 0.417394f
C1865 sarlogic_0/FILLER_0_7_195/a_124_375# 0 0.246306f
C1866 sarlogic_0/FILLER_0_7_162/a_36_472# 0 0.417394f
C1867 sarlogic_0/FILLER_0_7_162/a_124_375# 0 0.246306f
C1868 sarlogic_0/output13/a_224_472# 0 2.38465f
C1869 sarlogic_0/FILLER_0_18_2/a_3172_472# 0 0.345058f
C1870 sarlogic_0/FILLER_0_18_2/a_2724_472# 0 0.33241f
C1871 sarlogic_0/FILLER_0_18_2/a_2276_472# 0 0.33241f
C1872 sarlogic_0/FILLER_0_18_2/a_1828_472# 0 0.33241f
C1873 sarlogic_0/FILLER_0_18_2/a_1380_472# 0 0.33241f
C1874 sarlogic_0/FILLER_0_18_2/a_932_472# 0 0.33241f
C1875 sarlogic_0/FILLER_0_18_2/a_484_472# 0 0.33241f
C1876 sarlogic_0/FILLER_0_18_2/a_36_472# 0 0.404746f
C1877 sarlogic_0/FILLER_0_18_2/a_3260_375# 0 0.233093f
C1878 sarlogic_0/FILLER_0_18_2/a_2812_375# 0 0.17167f
C1879 sarlogic_0/FILLER_0_18_2/a_2364_375# 0 0.17167f
C1880 sarlogic_0/FILLER_0_18_2/a_1916_375# 0 0.17167f
C1881 sarlogic_0/FILLER_0_18_2/a_1468_375# 0 0.17167f
C1882 sarlogic_0/FILLER_0_18_2/a_1020_375# 0 0.17167f
C1883 sarlogic_0/FILLER_0_18_2/a_572_375# 0 0.17167f
C1884 sarlogic_0/FILLER_0_18_2/a_124_375# 0 0.185915f
C1885 sarlogic_0/net46 0 1.13395f
C1886 sarlogic_0/output46/a_224_472# 0 2.38465f
C1887 result[8] 0 17.026022f
C1888 sarlogic_0/output35/a_224_472# 0 2.38465f
C1889 sarlogic_0/output24/a_224_472# 0 2.38465f
C1890 sarlogic_0/FILLER_0_8_107/a_36_472# 0 0.417394f
C1891 sarlogic_0/FILLER_0_8_107/a_124_375# 0 0.246306f
C1892 sarlogic_0/FILLER_0_12_124/a_36_472# 0 0.417394f
C1893 sarlogic_0/FILLER_0_12_124/a_124_375# 0 0.246306f
C1894 sarlogic_0/net41 0 1.746759f
C1895 sarlogic_0/_065_ 0 0.523724f
C1896 sarlogic_0/_239_/a_36_160# 0 0.696445f
C1897 sarlogic_0/FILLER_0_1_98/a_36_472# 0 0.417394f
C1898 sarlogic_0/FILLER_0_1_98/a_124_375# 0 0.246306f
C1899 sarlogic_0/_115_ 0 1.281516f
C1900 sarlogic_0/_114_ 0 2.293579f
C1901 sarlogic_0/_308_/a_848_380# 0 0.40208f
C1902 sarlogic_0/_308_/a_124_24# 0 0.591898f
C1903 sarlogic_0/_256_/a_36_68# 0 0.063181f
C1904 sarlogic_0/FILLER_0_10_78/a_1380_472# 0 0.345058f
C1905 sarlogic_0/FILLER_0_10_78/a_932_472# 0 0.33241f
C1906 sarlogic_0/FILLER_0_10_78/a_484_472# 0 0.33241f
C1907 sarlogic_0/FILLER_0_10_78/a_36_472# 0 0.404746f
C1908 sarlogic_0/FILLER_0_10_78/a_1468_375# 0 0.233029f
C1909 sarlogic_0/FILLER_0_10_78/a_1020_375# 0 0.171606f
C1910 sarlogic_0/FILLER_0_10_78/a_572_375# 0 0.171606f
C1911 sarlogic_0/FILLER_0_10_78/a_124_375# 0 0.185399f
C1912 sarlogic_0/_130_ 0 0.304085f
C1913 sarlogic_0/net80 0 1.375599f
C1914 sarlogic_0/fanout80/a_36_113# 0 0.418095f
C1915 sarlogic_0/net58 0 5.308423f
C1916 sarlogic_0/_000_ 0 0.382358f
C1917 sarlogic_0/net75 0 1.474299f
C1918 sarlogic_0/_411_/a_2560_156# 0 0.016968f
C1919 sarlogic_0/_411_/a_2665_112# 0 0.62251f
C1920 sarlogic_0/_411_/a_2248_156# 0 0.371662f
C1921 sarlogic_0/_411_/a_1204_472# 0 0.012971f
C1922 sarlogic_0/_411_/a_1000_472# 0 0.291735f
C1923 sarlogic_0/_411_/a_796_472# 0 0.023206f
C1924 sarlogic_0/_411_/a_1308_423# 0 0.279043f
C1925 sarlogic_0/_411_/a_448_472# 0 0.684413f
C1926 sarlogic_0/_411_/a_36_151# 0 1.43589f
C1927 sarlogic_0/state\[0\] 0 0.680109f
C1928 sarlogic_0/_273_/a_36_68# 0 0.69549f
C1929 sarlogic_0/_142_ 0 0.324372f
C1930 sarlogic_0/FILLER_0_9_223/a_484_472# 0 0.345058f
C1931 sarlogic_0/FILLER_0_9_223/a_36_472# 0 0.404746f
C1932 sarlogic_0/FILLER_0_9_223/a_572_375# 0 0.232991f
C1933 sarlogic_0/FILLER_0_9_223/a_124_375# 0 0.185089f
C1934 sarlogic_0/FILLER_0_4_197/a_1380_472# 0 0.345058f
C1935 sarlogic_0/FILLER_0_4_197/a_932_472# 0 0.33241f
C1936 sarlogic_0/FILLER_0_4_197/a_484_472# 0 0.33241f
C1937 sarlogic_0/FILLER_0_4_197/a_36_472# 0 0.404746f
C1938 sarlogic_0/FILLER_0_4_197/a_1468_375# 0 0.233029f
C1939 sarlogic_0/FILLER_0_4_197/a_1020_375# 0 0.171606f
C1940 sarlogic_0/FILLER_0_4_197/a_572_375# 0 0.171606f
C1941 sarlogic_0/FILLER_0_4_197/a_124_375# 0 0.185399f
C1942 sarlogic_0/FILLER_0_17_226/a_36_472# 0 0.417394f
C1943 sarlogic_0/FILLER_0_17_226/a_124_375# 0 0.246306f
C1944 sarlogic_0/FILLER_0_5_109/a_484_472# 0 0.345058f
C1945 sarlogic_0/FILLER_0_5_109/a_36_472# 0 0.404746f
C1946 sarlogic_0/FILLER_0_5_109/a_572_375# 0 0.232991f
C1947 sarlogic_0/FILLER_0_5_109/a_124_375# 0 0.185089f
C1948 sarlogic_0/output12/a_224_472# 0 2.38465f
C1949 result[7] 0 16.58521f
C1950 sarlogic_0/net34 0 1.724665f
C1951 sarlogic_0/output34/a_224_472# 0 2.38465f
C1952 sarlogic_0/net45 0 1.12041f
C1953 sarlogic_0/output45/a_224_472# 0 2.38465f
C1954 sarlogic_0/output23/a_224_472# 0 2.38465f
C1955 sarlogic_0/FILLER_0_15_142/a_484_472# 0 0.345058f
C1956 sarlogic_0/FILLER_0_15_142/a_36_472# 0 0.404746f
C1957 sarlogic_0/FILLER_0_15_142/a_572_375# 0 0.232991f
C1958 sarlogic_0/FILLER_0_15_142/a_124_375# 0 0.185089f
C1959 sarlogic_0/_077_ 0 1.645892f
C1960 sarlogic_0/_075_ 0 0.374516f
C1961 sarlogic_0/_257_/a_36_472# 0 0.031137f
C1962 sarlogic_0/_326_/a_36_160# 0 0.696445f
C1963 sarlogic_0/_412_/a_2560_156# 0 0.016968f
C1964 sarlogic_0/_412_/a_2665_112# 0 0.62251f
C1965 sarlogic_0/_412_/a_2248_156# 0 0.371662f
C1966 sarlogic_0/_412_/a_1204_472# 0 0.012971f
C1967 sarlogic_0/_412_/a_1000_472# 0 0.291735f
C1968 sarlogic_0/_412_/a_796_472# 0 0.023206f
C1969 sarlogic_0/_412_/a_1308_423# 0 0.279043f
C1970 sarlogic_0/_412_/a_448_472# 0 0.684413f
C1971 sarlogic_0/_412_/a_36_151# 0 1.43589f
C1972 sarlogic_0/_091_ 0 1.841339f
C1973 sarlogic_0/_274_/a_36_68# 0 0.063181f
C1974 sarlogic_0/_143_ 0 0.329289f
C1975 sarlogic_0/mask\[4\] 0 1.300438f
C1976 sarlogic_0/_343_/a_49_472# 0 0.054843f
C1977 sarlogic_0/FILLER_0_13_65/a_36_472# 0 0.417394f
C1978 sarlogic_0/FILLER_0_13_65/a_124_375# 0 0.246306f
C1979 sarlogic_0/_360_/a_36_160# 0 0.386641f
C1980 sarlogic_0/FILLER_0_4_185/a_36_472# 0 0.417394f
C1981 sarlogic_0/FILLER_0_4_185/a_124_375# 0 0.246306f
C1982 sarlogic_0/FILLER_0_4_152/a_36_472# 0 0.417394f
C1983 sarlogic_0/FILLER_0_4_152/a_124_375# 0 0.246306f
C1984 sarlogic_0/_291_/a_36_160# 0 0.386641f
C1985 sarlogic_0/output9/a_224_472# 0 2.38465f
C1986 sarlogic_0/output11/a_224_472# 0 2.38465f
C1987 sarlogic_0/output44/a_224_472# 0 2.38465f
C1988 result[6] 0 16.532772f
C1989 sarlogic_0/output33/a_224_472# 0 2.38465f
C1990 sarlogic_0/output22/a_224_472# 0 2.38465f
C1991 sarlogic_0/FILLER_0_8_127/a_36_472# 0 0.417394f
C1992 sarlogic_0/FILLER_0_8_127/a_124_375# 0 0.246306f
C1993 sarlogic_0/FILLER_0_8_138/a_36_472# 0 0.417394f
C1994 sarlogic_0/FILLER_0_8_138/a_124_375# 0 0.246306f
C1995 sarlogic_0/FILLER_0_21_133/a_36_472# 0 0.417394f
C1996 sarlogic_0/FILLER_0_21_133/a_124_375# 0 0.246306f
C1997 sarlogic_0/FILLER_0_24_130/a_36_472# 0 0.417394f
C1998 sarlogic_0/FILLER_0_24_130/a_124_375# 0 0.246306f
C1999 sarlogic_0/FILLER_0_18_171/a_36_472# 0 0.417394f
C2000 sarlogic_0/FILLER_0_18_171/a_124_375# 0 0.246306f
C2001 sarlogic_0/_258_/a_36_160# 0 0.386641f
C2002 sarlogic_0/_016_ 0 0.314121f
C2003 sarlogic_0/_327_/a_36_472# 0 0.031137f
C2004 sarlogic_0/_189_/a_67_603# 0 0.345683f
C2005 sarlogic_0/FILLER_0_24_63/a_36_472# 0 0.417394f
C2006 sarlogic_0/FILLER_0_24_63/a_124_375# 0 0.246306f
C2007 sarlogic_0/FILLER_0_24_96/a_36_472# 0 0.417394f
C2008 sarlogic_0/FILLER_0_24_96/a_124_375# 0 0.246306f
C2009 sarlogic_0/cal_itt\[2\] 0 1.473514f
C2010 sarlogic_0/_002_ 0 0.289553f
C2011 sarlogic_0/_413_/a_2560_156# 0 0.016968f
C2012 sarlogic_0/_413_/a_2665_112# 0 0.62251f
C2013 sarlogic_0/_413_/a_2248_156# 0 0.371662f
C2014 sarlogic_0/_413_/a_1204_472# 0 0.012971f
C2015 sarlogic_0/_413_/a_1000_472# 0 0.291735f
C2016 sarlogic_0/_413_/a_796_472# 0 0.023206f
C2017 sarlogic_0/_413_/a_1308_423# 0 0.279043f
C2018 sarlogic_0/_413_/a_448_472# 0 0.684413f
C2019 sarlogic_0/_413_/a_36_151# 0 1.43589f
C2020 sarlogic_0/_092_ 0 0.680239f
C2021 sarlogic_0/FILLER_0_7_72/a_3172_472# 0 0.345058f
C2022 sarlogic_0/FILLER_0_7_72/a_2724_472# 0 0.33241f
C2023 sarlogic_0/FILLER_0_7_72/a_2276_472# 0 0.33241f
C2024 sarlogic_0/FILLER_0_7_72/a_1828_472# 0 0.33241f
C2025 sarlogic_0/FILLER_0_7_72/a_1380_472# 0 0.33241f
C2026 sarlogic_0/FILLER_0_7_72/a_932_472# 0 0.33241f
C2027 sarlogic_0/FILLER_0_7_72/a_484_472# 0 0.33241f
C2028 sarlogic_0/FILLER_0_7_72/a_36_472# 0 0.404746f
C2029 sarlogic_0/FILLER_0_7_72/a_3260_375# 0 0.233093f
C2030 sarlogic_0/FILLER_0_7_72/a_2812_375# 0 0.17167f
C2031 sarlogic_0/FILLER_0_7_72/a_2364_375# 0 0.17167f
C2032 sarlogic_0/FILLER_0_7_72/a_1916_375# 0 0.17167f
C2033 sarlogic_0/FILLER_0_7_72/a_1468_375# 0 0.17167f
C2034 sarlogic_0/FILLER_0_7_72/a_1020_375# 0 0.17167f
C2035 sarlogic_0/FILLER_0_7_72/a_572_375# 0 0.17167f
C2036 sarlogic_0/FILLER_0_7_72/a_124_375# 0 0.185915f
C2037 sarlogic_0/_086_ 0 2.45259f
C2038 sarlogic_0/_119_ 0 1.237181f
C2039 sarlogic_0/net63 0 5.362473f
C2040 sarlogic_0/_430_/a_2560_156# 0 0.016968f
C2041 sarlogic_0/_430_/a_2665_112# 0 0.62251f
C2042 sarlogic_0/_430_/a_2248_156# 0 0.371662f
C2043 sarlogic_0/_430_/a_1204_472# 0 0.012971f
C2044 sarlogic_0/_430_/a_1000_472# 0 0.291735f
C2045 sarlogic_0/_430_/a_796_472# 0 0.023206f
C2046 sarlogic_0/_430_/a_1308_423# 0 0.279043f
C2047 sarlogic_0/_430_/a_448_472# 0 0.684413f
C2048 sarlogic_0/_430_/a_36_151# 0 1.43589f
C2049 sarlogic_0/_292_/a_36_160# 0 0.386641f
C2050 sarlogic_0/output8/a_224_472# 0 2.38465f
C2051 sarlogic_0/output10/a_224_472# 0 2.38465f
C2052 result[5] 0 16.544518f
C2053 sarlogic_0/net32 0 1.78884f
C2054 sarlogic_0/output32/a_224_472# 0 2.38465f
C2055 sarlogic_0/output43/a_224_472# 0 2.38465f
C2056 sarlogic_0/output21/a_224_472# 0 2.38465f
C2057 sarlogic_0/_053_ 0 1.705161f
C2058 sarlogic_0/FILLER_0_16_107/a_484_472# 0 0.345058f
C2059 sarlogic_0/FILLER_0_16_107/a_36_472# 0 0.404746f
C2060 sarlogic_0/FILLER_0_16_107/a_572_375# 0 0.232991f
C2061 sarlogic_0/FILLER_0_16_107/a_124_375# 0 0.185089f
C2062 sarlogic_0/FILLER_0_3_204/a_36_472# 0 0.417394f
C2063 sarlogic_0/FILLER_0_3_204/a_124_375# 0 0.246306f
C2064 sarlogic_0/FILLER_0_9_28/a_3172_472# 0 0.345058f
C2065 sarlogic_0/FILLER_0_9_28/a_2724_472# 0 0.33241f
C2066 sarlogic_0/FILLER_0_9_28/a_2276_472# 0 0.33241f
C2067 sarlogic_0/FILLER_0_9_28/a_1828_472# 0 0.33241f
C2068 sarlogic_0/FILLER_0_9_28/a_1380_472# 0 0.33241f
C2069 sarlogic_0/FILLER_0_9_28/a_932_472# 0 0.33241f
C2070 sarlogic_0/FILLER_0_9_28/a_484_472# 0 0.33241f
C2071 sarlogic_0/FILLER_0_9_28/a_36_472# 0 0.404746f
C2072 sarlogic_0/FILLER_0_9_28/a_3260_375# 0 0.233093f
C2073 sarlogic_0/FILLER_0_9_28/a_2812_375# 0 0.17167f
C2074 sarlogic_0/FILLER_0_9_28/a_2364_375# 0 0.17167f
C2075 sarlogic_0/FILLER_0_9_28/a_1916_375# 0 0.17167f
C2076 sarlogic_0/FILLER_0_9_28/a_1468_375# 0 0.17167f
C2077 sarlogic_0/FILLER_0_9_28/a_1020_375# 0 0.17167f
C2078 sarlogic_0/FILLER_0_9_28/a_572_375# 0 0.17167f
C2079 sarlogic_0/FILLER_0_9_28/a_124_375# 0 0.185915f
C2080 sarlogic_0/_132_ 0 1.491425f
C2081 sarlogic_0/_328_/a_36_113# 0 0.418095f
C2082 sarlogic_0/_414_/a_2560_156# 0 0.016968f
C2083 sarlogic_0/_414_/a_2665_112# 0 0.62251f
C2084 sarlogic_0/_414_/a_2248_156# 0 0.371662f
C2085 sarlogic_0/_414_/a_1204_472# 0 0.012971f
C2086 sarlogic_0/_414_/a_1000_472# 0 0.291735f
C2087 sarlogic_0/_414_/a_796_472# 0 0.023206f
C2088 sarlogic_0/_414_/a_1308_423# 0 0.279043f
C2089 sarlogic_0/_414_/a_448_472# 0 0.684413f
C2090 sarlogic_0/_414_/a_36_151# 0 1.43589f
C2091 sarlogic_0/_276_/a_36_160# 0 0.386641f
C2092 sarlogic_0/_144_ 0 1.173846f
C2093 sarlogic_0/_345_/a_36_160# 0 0.386641f
C2094 sarlogic_0/_155_ 0 0.638535f
C2095 sarlogic_0/_020_ 0 0.316793f
C2096 sarlogic_0/_431_/a_2560_156# 0 0.016968f
C2097 sarlogic_0/_431_/a_2665_112# 0 0.62251f
C2098 sarlogic_0/_431_/a_2248_156# 0 0.371662f
C2099 sarlogic_0/_431_/a_1204_472# 0 0.012971f
C2100 sarlogic_0/_431_/a_1000_472# 0 0.291735f
C2101 sarlogic_0/_431_/a_796_472# 0 0.023206f
C2102 sarlogic_0/_431_/a_1308_423# 0 0.279043f
C2103 sarlogic_0/_431_/a_448_472# 0 0.684413f
C2104 sarlogic_0/_431_/a_36_151# 0 1.43589f
C2105 sarlogic_0/_105_ 0 1.21281f
C2106 sarlogic_0/_293_/a_36_472# 0 0.031137f
C2107 sarlogic_0/FILLER_0_5_128/a_484_472# 0 0.345058f
C2108 sarlogic_0/FILLER_0_5_128/a_36_472# 0 0.404746f
C2109 sarlogic_0/FILLER_0_5_128/a_572_375# 0 0.232991f
C2110 sarlogic_0/FILLER_0_5_128/a_124_375# 0 0.185089f
C2111 sarlogic_0/FILLER_0_5_117/a_36_472# 0 0.417394f
C2112 sarlogic_0/FILLER_0_5_117/a_124_375# 0 0.246306f
C2113 sarlogic_0/net7 0 1.174913f
C2114 sarlogic_0/output7/a_224_472# 0 2.38465f
C2115 sarlogic_0/output42/a_224_472# 0 2.38465f
C2116 result[4] 0 16.37653f
C2117 sarlogic_0/net31 0 1.912935f
C2118 sarlogic_0/output31/a_224_472# 0 2.38465f
C2119 sarlogic_0/output20/a_224_472# 0 2.38465f
C2120 sarlogic_0/FILLER_0_16_73/a_484_472# 0 0.345058f
C2121 sarlogic_0/FILLER_0_16_73/a_36_472# 0 0.404746f
C2122 sarlogic_0/FILLER_0_16_73/a_572_375# 0 0.232991f
C2123 sarlogic_0/FILLER_0_16_73/a_124_375# 0 0.185089f
C2124 sarlogic_0/FILLER_0_21_142/a_484_472# 0 0.345058f
C2125 sarlogic_0/FILLER_0_21_142/a_36_472# 0 0.404746f
C2126 sarlogic_0/FILLER_0_21_142/a_572_375# 0 0.232991f
C2127 sarlogic_0/FILLER_0_21_142/a_124_375# 0 0.185089f
C2128 sarlogic_0/FILLER_0_15_150/a_36_472# 0 0.417394f
C2129 sarlogic_0/FILLER_0_15_150/a_124_375# 0 0.246306f
C2130 sarlogic_0/FILLER_0_19_125/a_36_472# 0 0.417394f
C2131 sarlogic_0/FILLER_0_19_125/a_124_375# 0 0.246306f
C2132 sarlogic_0/net10 0 1.480101f
C2133 sarlogic_0/net20 0 2.034189f
C2134 sarlogic_0/_277_/a_36_160# 0 0.386641f
C2135 sarlogic_0/net27 0 2.023744f
C2136 sarlogic_0/_004_ 0 0.390107f
C2137 sarlogic_0/_415_/a_2560_156# 0 0.016968f
C2138 sarlogic_0/_415_/a_2665_112# 0 0.62251f
C2139 sarlogic_0/_415_/a_2248_156# 0 0.371662f
C2140 sarlogic_0/_415_/a_1204_472# 0 0.012971f
C2141 sarlogic_0/_415_/a_1000_472# 0 0.291735f
C2142 sarlogic_0/_415_/a_796_472# 0 0.023206f
C2143 sarlogic_0/_415_/a_1308_423# 0 0.279043f
C2144 sarlogic_0/_415_/a_448_472# 0 0.684413f
C2145 sarlogic_0/_415_/a_36_151# 0 1.43589f
C2146 sarlogic_0/mask\[5\] 0 1.334568f
C2147 sarlogic_0/_346_/a_49_472# 0 0.054843f
C2148 sarlogic_0/_028_ 0 0.386029f
C2149 sarlogic_0/_363_/a_36_68# 0 0.150048f
C2150 sarlogic_0/_021_ 0 0.316776f
C2151 sarlogic_0/_432_/a_2560_156# 0 0.016968f
C2152 sarlogic_0/_432_/a_2665_112# 0 0.62251f
C2153 sarlogic_0/_432_/a_2248_156# 0 0.371662f
C2154 sarlogic_0/_432_/a_1204_472# 0 0.012971f
C2155 sarlogic_0/_432_/a_1000_472# 0 0.291735f
C2156 sarlogic_0/_432_/a_796_472# 0 0.023206f
C2157 sarlogic_0/_432_/a_1308_423# 0 0.279043f
C2158 sarlogic_0/_432_/a_448_472# 0 0.684413f
C2159 sarlogic_0/_432_/a_36_151# 0 1.43589f
C2160 sarlogic_0/_008_ 0 0.423631f
C2161 sarlogic_0/_104_ 0 1.435764f
C2162 sarlogic_0/_106_ 0 0.378703f
C2163 sarlogic_0/FILLER_0_17_200/a_484_472# 0 0.345058f
C2164 sarlogic_0/FILLER_0_17_200/a_36_472# 0 0.404746f
C2165 sarlogic_0/FILLER_0_17_200/a_572_375# 0 0.232991f
C2166 sarlogic_0/FILLER_0_17_200/a_124_375# 0 0.185089f
C2167 vss 0 10.515274p
C2168 comparator_0/trim_left_0/n0 0 0.627477f
C2169 comparator_0/trim_left_0/n1 0 0.643951f
C2170 comparator_0/trim_left_0/n4 0 4.635427f
C2171 comparator_0/in 0 -7.798843f
C2172 comparator_0/trim_left_0/n3 0 3.342805f
C2173 comparator_0/trim_left_0/n2 0 1.998525f
C2174 sarlogic_0/trim[3] 0 10.909932f
C2175 sarlogic_0/trim[2] 0 5.259631f
C2176 sarlogic_0/trim[1] 0 5.593644f
C2177 sarlogic_0/trim[0] 0 4.848347f
C2178 sarlogic_0/trim[4] 0 10.616135f
C2179 latch_0/S 0 6.241351f
C2180 latch_0/R 0 4.698747f
C2181 sarlogic_0/trimb[1] 0 5.208551f
C2182 sarlogic_0/trimb[4] 0 10.649281f
C2183 sarlogic_0/trimb[2] 0 5.266952f
C2184 sarlogic_0/trimb[0] 0 4.941973f
C2185 sarlogic_0/trimb[3] 0 9.450794f
C2186 comparator_0/trim_right_0/n0 0 0.627477f
C2187 comparator_0/trim_right_0/n1 0 0.643951f
C2188 comparator_0/trim_right_0/n4 0 4.635427f
C2189 comparator_0/ip 0 -7.798843f
C2190 comparator_0/trim_right_0/n3 0 3.342805f
C2191 comparator_0/trim_right_0/n2 0 1.998525f
C2192 comparator_0/diff 0 0.212313f
C2193 buffer_0/buf_out 0 8.064797f
C2194 dacn_0/carray_n_0/n9 0 14.963586f
C2195 dacn_0/dac_out 0 -0.683058p
C2196 dacn_0/carray_n_0/n8 0 40.580837f
C2197 dacn_0/carray_n_0/n7 0 56.915478f
C2198 dacn_0/carray_n_0/n6 0 53.64827f
C2199 dacn_0/carray_n_0/n0 0 17.632519f
C2200 dacn_0/carray_n_0/n1 0 17.795374f
C2201 dacn_0/carray_n_0/n2 0 30.783176f
C2202 dacn_0/carray_n_0/n3 0 34.265587f
C2203 dacn_0/carray_n_0/n4 0 39.983223f
C2204 dacn_0/carray_n_0/n5 0 48.00648f
C2205 vinn 0 27.34083f
C2206 dacn_0/bootstrapped_sw_n_0/vg 0 1.498165f
C2207 dacn_0/bootstrapped_sw_n_0/vbsh 0 14.27723f
C2208 dacn_0/bootstrapped_sw_n_0/vbsl 0 7.956583f
C2209 dacp_0/sample 0 92.15834f
C2210 dacn_0/bootstrapped_sw_n_0/vs 0 0.053987f
C2211 dacn_0/bootstrapped_sw_n_0/enb 0 1.502816f
C2212 dacn_0/ctl9 0 7.033419f
C2213 dacn_0/ctl8 0 7.441137f
C2214 dacn_0/ctl7 0 10.297702f
C2215 dacn_0/ctl6 0 11.395121f
C2216 dacn_0/ctl5 0 12.440359f
C2217 dacn_0/ctl4 0 13.228794f
C2218 dacn_0/ctl3 0 13.514038f
C2219 dacn_0/ctl1 0 20.84428f
C2220 dacn_0/ctl10 0 9.550506f
C2221 dacn_0/ctl2 0 15.423438f
C2222 dacn_0/carray_n_0/ndum 0 14.881693f
C2223 dacp_0/carray_p_0/n2 0 30.783176f
C2224 dacp_0/carray_p_0/n3 0 34.265587f
C2225 dacp_0/carray_p_0/n4 0 39.983223f
C2226 dacp_0/carray_p_0/n5 0 48.00648f
C2227 dacp_0/carray_p_0/n9 0 14.963586f
C2228 dacp_0/dac_out 0 -0.681098p
C2229 dacp_0/carray_p_0/n8 0 40.580837f
C2230 dacp_0/carray_p_0/n7 0 56.915478f
C2231 dacp_0/carray_p_0/n6 0 53.64827f
C2232 dacp_0/carray_p_0/n0 0 17.632519f
C2233 dacp_0/carray_p_0/n1 0 17.795374f
C2234 dacp_0/bootstrapped_sw_p_0/vs 0 0.053987f
C2235 dacp_0/bootstrapped_sw_p_0/enb 0 1.502816f
C2236 vinp 0 27.34083f
C2237 dacp_0/bootstrapped_sw_p_0/vg 0 1.498165f
C2238 dacp_0/bootstrapped_sw_p_0/vbsh 0 14.27723f
C2239 dacp_0/bootstrapped_sw_p_0/vbsl 0 7.956583f
C2240 dacp_0/ctl9 0 6.604383f
C2241 dacp_0/ctl8 0 7.029485f
C2242 dacp_0/ctl7 0 9.867429f
C2243 dacp_0/ctl6 0 11.186495f
C2244 dacp_0/ctl5 0 12.138051f
C2245 dacp_0/ctl4 0 12.142579f
C2246 dacp_0/ctl3 0 13.828307f
C2247 dacp_0/ctl1 0 19.89871f
C2248 dacp_0/ctl10 0 9.136993f
C2249 dacp_0/ctl2 0 13.765609f
C2250 dacp_0/carray_p_0/ndum 0 14.881693f
C2251 sarlogic_0/clkc 0 7.220488f
C2252 buffer_0/inv2_0/inv_in 0 0.832311f
C2253 latch_0/Qn 0 0.887927f
C2254 latch_0/Q 0 7.192533f
C2255 latch_0/tutyuu2 0 0.717123f
C2256 latch_0/tutyuu1 0 0.717027f
.ends

