* NGSPICE file created from mim_cap_30_30.ext - technology: gf180mcuD

.subckt cap_mim_2p0fF_RCWXT2
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
.ends


* Top level circuit mim_cap_30_30

Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2
.end

