* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

.subckt XM2_x4_latch G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_x4_latch G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt x4_latch inv_out inv_in vdd vss
XXM2_x4_latch_0 inv_in inv_out vdd vdd XM2_x4_latch
XXM1_x4_latch_0 inv_in inv_out vss vss XM1_x4_latch
.ends

.subckt XM2_x3_latch G D w_n319_n356# S
MX0 S G D w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_x3_latch G D a_n319_n324# S
MX0 S G D a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt x3_latch inv_out inv_in vdd vss
XXM2_x3_latch_0 inv_in inv_out vdd vdd XM2_x3_latch
XXM1_x3_latch_0 inv_in inv_out vss vss XM1_x3_latch
.ends

.subckt XM4_latch G D a_n319_n324# S a_n319_252#
MX0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_x2_latch G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_x2_latch G a_n320_n324# D a_n318_252# S
MX0 D G S a_n320_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt x2_latch inv_out inv_in XM1_x2_latch_0/a_n318_252# vdd vss
XXM2_x2_latch_0 inv_in inv_out vdd vdd XM2_x2_latch
XXM1_x2_latch_0 inv_in vss inv_out XM1_x2_latch_0/a_n318_252# vss XM1_x2_latch
.ends

.subckt XM3_latch G D a_n319_n324# S a_n319_252#
MX0 D G S a_n319_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_x1_latch G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_x1_latch G D a_n318_252# a_n318_n324# S
MX0 D G S a_n318_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt x1_latch inv_out inv_in XM1_x1_latch_0/a_n318_252# vdd vss
XXM2_x1_latch_0 inv_in inv_out vdd vdd XM2_x1_latch
XXM1_x1_latch_0 inv_in inv_out XM1_x1_latch_0/a_n318_252# vss vss XM1_x1_latch
.ends

.subckt latch Q Qn R S tutyuu1 tutyuu2 vdd vss
Xx4_latch_0 tutyuu1 S vdd vss x4_latch
Xx3_latch_0 tutyuu2 R vdd vss x3_latch
XXM4_latch_0 tutyuu2 Q vss vss vss XM4_latch
Xx2_latch_0 Qn Q vss vdd vss x2_latch
XXM3_latch_0 tutyuu1 Qn vss vss vss XM3_latch
Xx1_latch_0 Q Qn vss vdd vss x1_latch
.ends

.subckt XM1_inv2 VSUBS G D S
MX0 D G S VSUBS nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_inv2 VSUBS G D S
MX0 D G S VSUBS pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt inv2 inv_out inv_in vss
XXM1_inv2_0 vss inv_in inv_out vss XM1_inv2
XXM2_inv2_0 vss inv_in inv_out vss XM2_inv2
.ends

.subckt XM1_inv1 VSUBS G D S
MX0 D G S VSUBS nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_inv1 VSUBS G D S
MX0 D G S VSUBS pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt inv1 inv_out inv_in vss
XXM1_inv1_0 vss inv_in inv_out vss XM1_inv1
XXM2_inv1_0 vss inv_in inv_out vss XM2_inv1
.ends

.subckt buffer buf_in buf_out vss
Xinv2_0 buf_out inv2_0/inv_in vss inv2
Xinv1_0 inv2_0/inv_in buf_in vss inv1
.ends

.subckt inv_p VSS ZN I VDD VPW VNW
MX0 VDD I ZN VNW pfet_06v0 ad=1.21p pd=4.42u as=0.457p ps=1.97u w=1.22u l=0.5u M=2
MX1 ZN I VSS VPW nfet_06v0 ad=0.225p pd=1.37u as=0.508p ps=2.88u w=0.82u l=0.6u M=2
.ends

.subckt inv_renketu_p inv_p_3/I inv_p_9/ZN inv_p_6/ZN inv_p_6/I inv_p_8/I inv_p_0/ZN
+ inv_p_8/ZN inv_p_5/ZN inv_p_7/I inv_p_2/I inv_p_0/I inv_p_2/ZN inv_p_4/ZN inv_p_9/I
+ inv_p_10/I inv_p_7/ZN inv_p_5/I inv_p_1/ZN inv_p_3/ZN inv_p_4/I inv_p_10/ZN inv_p_1/I
+ vdd vss
Xinv_p_0 vss inv_p_0/ZN inv_p_0/I vdd vss vdd inv_p
Xinv_p_1 vss inv_p_1/ZN inv_p_1/I vdd vss vdd inv_p
Xinv_p_2 vss inv_p_2/ZN inv_p_2/I vdd vss vdd inv_p
Xinv_p_3 vss inv_p_3/ZN inv_p_3/I vdd vss vdd inv_p
Xinv_p_4 vss inv_p_4/ZN inv_p_4/I vdd vss vdd inv_p
Xinv_p_5 vss inv_p_5/ZN inv_p_5/I vdd vss vdd inv_p
Xinv_p_6 vss inv_p_6/ZN inv_p_6/I vdd vss vdd inv_p
Xinv_p_7 vss inv_p_7/ZN inv_p_7/I vdd vss vdd inv_p
Xinv_p_8 vss inv_p_8/ZN inv_p_8/I vdd vss vdd inv_p
Xinv_p_9 vss inv_p_9/ZN inv_p_9/I vdd vss vdd inv_p
Xinv_p_10 vss inv_p_10/ZN inv_p_10/I vdd vss vdd inv_p
.ends

.subckt XMs2_bs_p G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM3_bs_p G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM2_bs_inv_p G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_bs_inv_p G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt bs_inv_p inv_out vdd inv_in vss
XXM2_bs_inv_p_0 inv_in inv_out vdd vdd XM2_bs_inv_p
XXM1_bs_inv_p_0 inv_in inv_out vss vss XM1_bs_inv_p
.ends

.subckt XM4_bs_p G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt bs_cap_p I1_1_1_R0_BOT I1_1_1_R0_TOP
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.3u c_length=12.3u
.ends

.subckt XMs_bs_p G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM1_bs_p G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XMs1_bs_p G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_bs_p G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt bootstrapped_sw_p vdd en enb bs_in bs_out vg vs vbsh vbsl vss
XXMs2_bs_p_0 enb vss vss vss vs XMs2_bs_p
XXM3_bs_p_0 enb vg vbsh vbsh XM3_bs_p
Xbs_inv_p_0 enb vdd en vss bs_inv_p
XXM4_bs_p_0 vg vdd vbsh vbsh XM4_bs_p
Xbs_cap_p_0 vbsl vbsh bs_cap_p
Xbs_cap_p_1 vbsl vbsh bs_cap_p
Xbs_cap_p_2 vbsl vbsh bs_cap_p
Xbs_cap_p_3 vbsl vbsh bs_cap_p
Xbs_cap_p_4 vbsl vbsh bs_cap_p
XXMs_bs_p_0 vg bs_out vss bs_in XMs_bs_p
XXM1_bs_p_0 vg vbsl vss vss bs_in XM1_bs_p
XXMs1_bs_p_0 vdd vs vss vg XMs1_bs_p
XXM2_bs_p_0 enb vbsl vss vss vss XM2_bs_p
.ends

.subckt dacp dac_in dac_out dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10
+ sample vdd_uq0 vdd vss
Xinv_renketu_p_0 ctl1 carray_p_0/n8 carray_p_0/n5 ctl5 ctl7 carray_p_0/ndum carray_p_0/n7
+ carray_p_0/n4 ctl6 ctl10 dum carray_p_0/n0 carray_p_0/n3 ctl8 ctl9 carray_p_0/n6
+ ctl4 carray_p_0/n2 carray_p_0/n1 ctl3 carray_p_0/n9 ctl2 vdd vss inv_renketu_p
Xbootstrapped_sw_p_0 vdd_uq0 sample bootstrapped_sw_p_0/enb dac_in dac_out bootstrapped_sw_p_0/vg
+ bootstrapped_sw_p_0/vs bootstrapped_sw_p_0/vbsh bootstrapped_sw_p_0/vbsl vss bootstrapped_sw_p
.ends

.subckt inv_n VSS ZN I VDD VPW VNW
MX0 VDD I ZN VNW pfet_06v0 ad=1.21p pd=4.42u as=0.457p ps=1.97u w=1.22u l=0.5u M=2
MX1 ZN I VSS VPW nfet_06v0 ad=0.225p pd=1.37u as=0.508p ps=2.88u w=0.82u l=0.6u M=2
.ends

.subckt inv_renketu_n inv_n_3/I inv_n_9/ZN inv_n_6/ZN inv_n_6/I inv_n_8/I inv_n_0/ZN
+ inv_n_8/ZN inv_n_5/ZN inv_n_7/I inv_n_2/I inv_n_0/I inv_n_2/ZN inv_n_4/ZN inv_n_9/I
+ inv_n_10/I inv_n_7/ZN inv_n_5/I inv_n_1/ZN inv_n_3/ZN vdd inv_n_4/I inv_n_10/ZN
+ inv_n_1/I vss
Xinv_n_0 vss inv_n_0/ZN inv_n_0/I vdd vss vdd inv_n
Xinv_n_1 vss inv_n_1/ZN inv_n_1/I vdd vss vdd inv_n
Xinv_n_2 vss inv_n_2/ZN inv_n_2/I vdd vss vdd inv_n
Xinv_n_3 vss inv_n_3/ZN inv_n_3/I vdd vss vdd inv_n
Xinv_n_4 vss inv_n_4/ZN inv_n_4/I vdd vss vdd inv_n
Xinv_n_5 vss inv_n_5/ZN inv_n_5/I vdd vss vdd inv_n
Xinv_n_6 vss inv_n_6/ZN inv_n_6/I vdd vss vdd inv_n
Xinv_n_7 vss inv_n_7/ZN inv_n_7/I vdd vss vdd inv_n
Xinv_n_8 vss inv_n_8/ZN inv_n_8/I vdd vss vdd inv_n
Xinv_n_9 vss inv_n_9/ZN inv_n_9/I vdd vss vdd inv_n
Xinv_n_10 vss inv_n_10/ZN inv_n_10/I vdd vss vdd inv_n
.ends

.subckt XMs1_bs_n G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_bs_n G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XMs2_bs_n G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM3_bs_n G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_bs_inv_n G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_bs_inv_n G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt bs_inv_n inv_out vdd inv_in vss
XXM1_bs_inv_n_0 inv_in inv_out vss vss XM1_bs_inv_n
XXM2_bs_inv_n_0 inv_in inv_out vdd vdd XM2_bs_inv_n
.ends

.subckt XM4_bs_n G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt bs_cap_n I1_1_1_R0_BOT I1_1_1_R0_TOP
X0 I1_1_1_R0_TOP I1_1_1_R0_BOT cap_mim_2f0fF c_width=12.3u c_length=12.3u
.ends

.subckt XMs_bs_n G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM1_bs_n G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt bootstrapped_sw_n vdd en enb bs_in bs_out vg vs vbsh vbsl vss
XXMs1_bs_n_0 vdd vs vss vg XMs1_bs_n
XXM2_bs_n_0 enb vbsl vss vss vss XM2_bs_n
XXMs2_bs_n_0 enb vss vss vss vs XMs2_bs_n
XXM3_bs_n_0 enb vg vbsh vbsh XM3_bs_n
Xbs_inv_n_0 enb vdd en vss bs_inv_n
XXM4_bs_n_0 vg vdd vbsh vbsh XM4_bs_n
Xbs_cap_n_0 vbsl vbsh bs_cap_n
Xbs_cap_n_1 vbsl vbsh bs_cap_n
Xbs_cap_n_2 vbsl vbsh bs_cap_n
Xbs_cap_n_4 vbsl vbsh bs_cap_n
Xbs_cap_n_3 vbsl vbsh bs_cap_n
XXMs_bs_n_0 vg bs_out vss bs_in XMs_bs_n
XXM1_bs_n_0 vg vbsl vss vss bs_in XM1_bs_n
.ends

.subckt dacn dac_in dac_out dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10
+ sample vdd_uq0 vdd vss
Xinv_renketu_n_0 ctl1 carray_n_0/n8 carray_n_0/n5 ctl5 ctl7 carray_n_0/ndum carray_n_0/n7
+ carray_n_0/n4 ctl6 ctl10 dum carray_n_0/n0 carray_n_0/n3 ctl8 ctl9 carray_n_0/n6
+ ctl4 carray_n_0/n2 carray_n_0/n1 vdd ctl3 carray_n_0/n9 ctl2 vss inv_renketu_n
Xbootstrapped_sw_n_0 vdd_uq0 sample bootstrapped_sw_n_0/enb dac_in dac_out bootstrapped_sw_n_0/vg
+ bootstrapped_sw_n_0/vs bootstrapped_sw_n_0/vbsh bootstrapped_sw_n_0/vbsl vss bootstrapped_sw_n
.ends

.subckt XMdiff_cmp a_192_n100# a_n280_n100# a_n192_n183# a_n52_n100# a_n424_n324#
+ a_52_n183#
MX0 a_192_n100# a_52_n183# a_n52_n100# a_n424_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
MX1 a_n52_n100# a_n192_n183# a_n280_n100# a_n424_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM3_trims_right a_n2052_n100# a_n2668_n324# a_n1808_n100# a_n1948_n183# a_n1564_n100#
+ a_n2524_n100# a_n1704_n183# a_n2296_n100# a_n2192_n183# a_n2436_n183#
MX0 a_n2052_n100# a_n2192_n183# a_n2296_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX1 a_n1564_n100# a_n1704_n183# a_n1808_n100# a_n2668_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
MX2 a_n1808_n100# a_n1948_n183# a_n2052_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX3 a_n2296_n100# a_n2436_n183# a_n2524_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM0_trims_right G D a_n5334_252# a_n5334_n324# S
MX0 S G D a_n5334_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_trims_right a_n4456_n324# a_n3948_n183# a_n3808_n100# a_n4280_n100# a_n4052_n100#
+ a_n4192_n183# a_n4456_252#
MX0 a_n4052_n100# a_n4192_n183# a_n4280_n100# a_n4456_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
MX1 a_n3808_n100# a_n3948_n183# a_n4052_n100# a_n4456_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
.ends

.subckt XM4_trims_right a_436_n100# a_192_n100# a_n1188_n324# a_n296_n100# a_784_n183#
+ a_n192_n183# a_n436_n183# a_540_n183# a_n52_n100# a_924_n100# a_680_n100# a_n1012_n100#
+ a_n784_n100# a_n924_n183# a_n680_n183# a_n540_n100# a_296_n183# a_52_n183#
MX0 a_436_n100# a_296_n183# a_192_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX1 a_n784_n100# a_n924_n183# a_n1012_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
MX2 a_192_n100# a_52_n183# a_n52_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX3 a_680_n100# a_540_n183# a_436_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX4 a_924_n100# a_784_n183# a_680_n100# a_n1188_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
MX5 a_n52_n100# a_n192_n183# a_n296_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX6 a_n296_n100# a_n436_n183# a_n540_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX7 a_n540_n100# a_n680_n183# a_n784_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
.ends

.subckt XM1_trims_right G D a_n5302_n324# S a_n5302_252#
MX0 D G S a_n5302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt trim_switch_right d_0 d_4 d_1 d_2 d_3 n4 n2 n3 n1 n0 VSUBS
XXM3_trims_right_0 n3 VSUBS VSUBS d_3 n3 n3 d_3 VSUBS d_3 d_3 XM3_trims_right
XXM0_trims_right_0 d_0 n0 VSUBS VSUBS VSUBS XM0_trims_right
XXM2_trims_right_0 VSUBS d_2 n2 n2 VSUBS d_2 VSUBS XM2_trims_right
XXM4_trims_right_0 n4 VSUBS VSUBS VSUBS d_4 d_4 d_4 d_4 n4 n4 VSUBS n4 VSUBS d_4 d_4
+ n4 d_4 d_4 XM4_trims_right
XXM1_trims_right_0 d_1 n1 VSUBS VSUBS VSUBS XM1_trims_right
.ends

.subckt trim_right d_0 d_4 d_1 d_2 d_3 drain n1 n4 n0 n2 n3 vss
Xtrim_switch_right_0 d_0 d_4 d_1 d_2 d_3 n4 n2 n3 n1 n0 vss trim_switch_right
.ends

.subckt XMinp_cmp G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM4_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XMl4_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XMinn_cmp G D a_n302_n324# a_n302_252# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XMl3_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM3_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XMl2_cmp G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XM1_cmp G D w_n319_n356# S
MX0 D G S w_n319_n356# pfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.55u
.ends

.subckt XMl1_cmp G D a_n302_n324# S
MX0 D G S a_n302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM4_trims_left a_436_n100# a_192_n100# a_n1188_n324# a_n296_n100# a_784_n183#
+ a_n192_n183# a_n436_n183# a_540_n183# a_n52_n100# a_924_n100# a_680_n100# a_n1012_n100#
+ a_n784_n100# a_n924_n183# a_n680_n183# a_n540_n100# a_296_n183# a_52_n183#
MX0 a_436_n100# a_296_n183# a_192_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX1 a_n784_n100# a_n924_n183# a_n1012_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
MX2 a_192_n100# a_52_n183# a_n52_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX3 a_680_n100# a_540_n183# a_436_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX4 a_924_n100# a_784_n183# a_680_n100# a_n1188_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
MX5 a_n52_n100# a_n192_n183# a_n296_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX6 a_n296_n100# a_n436_n183# a_n540_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX7 a_n540_n100# a_n680_n183# a_n784_n100# a_n1188_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
.ends

.subckt XM0_trims_left G D a_n5334_252# a_n5334_n324# S
MX0 S G D a_n5334_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM1_trims_left G D a_n5302_n324# S a_n5302_252#
MX0 D G S a_n5302_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt XM2_trims_left a_n4456_n324# a_n3948_n183# a_n3808_n100# a_n4280_n100# a_n4052_n100#
+ a_n4192_n183# a_n4456_252#
MX0 a_n4052_n100# a_n4192_n183# a_n4280_n100# a_n4456_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
MX1 a_n3808_n100# a_n3948_n183# a_n4052_n100# a_n4456_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
.ends

.subckt XM3_trims_left a_n2052_n100# a_n2668_n324# a_n1808_n100# a_n1948_n183# a_n1564_n100#
+ a_n2524_n100# a_n1704_n183# a_n2296_n100# a_n2192_n183# a_n2436_n183#
MX0 a_n2052_n100# a_n2192_n183# a_n2296_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX1 a_n1564_n100# a_n1704_n183# a_n1808_n100# a_n2668_n324# nfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.7u
MX2 a_n1808_n100# a_n1948_n183# a_n2052_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.7u
MX3 a_n2296_n100# a_n2436_n183# a_n2524_n100# a_n2668_n324# nfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.7u
.ends

.subckt trim_switch_left d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 VSUBS
XXM4_trims_left_0 n4 VSUBS VSUBS VSUBS d_4 d_4 d_4 d_4 n4 n4 VSUBS n4 VSUBS d_4 d_4
+ n4 d_4 d_4 XM4_trims_left
XXM0_trims_left_0 d_0 n0 VSUBS VSUBS VSUBS XM0_trims_left
XXM1_trims_left_0 d_1 n1 VSUBS VSUBS VSUBS XM1_trims_left
XXM2_trims_left_0 VSUBS d_2 n2 n2 VSUBS d_2 VSUBS XM2_trims_left
XXM3_trims_left_0 n3 VSUBS VSUBS d_3 n3 n3 d_3 VSUBS d_3 d_3 XM3_trims_left
.ends

.subckt trim_left d_0 d_4 d_1 d_2 d_3 drain n1 n4 n0 n2 n3 vss
Xtrim_switch_left_0 d_0 d_4 d_1 d_2 d_3 n1 n4 n0 n2 n3 vss trim_switch_left
.ends

.subckt comparator trim1 trim0 trim2 trim3 trim4 trimb4 trimb1 trimb0 trimb2 trimb3
+ vp vn outp outn in ip clkc diff vdd vss
XXMdiff_cmp_0 vss vss clkc diff vss clkc XMdiff_cmp
Xtrim_right_0 trimb0 trimb4 trimb1 trimb2 trimb3 ip trim_right_0/n1 trim_right_0/n4
+ trim_right_0/n0 trim_right_0/n2 trim_right_0/n3 vss trim_right
XXMinp_cmp_0 vp ip vss vss diff XMinp_cmp
XXM4_cmp_0 clkc ip vdd vdd XM4_cmp
XXMl4_cmp_0 outn outp vdd vdd XMl4_cmp
XXMinn_cmp_0 vn in vss vss diff XMinn_cmp
XXMl3_cmp_0 outp outn vdd vdd XMl3_cmp
XXM3_cmp_0 clkc outp vdd vdd XM3_cmp
XXMl2_cmp_0 outn outp vss ip XMl2_cmp
XXM2_cmp_0 clkc outn vdd vdd XM2_cmp
XXM1_cmp_0 clkc in vdd vdd XM1_cmp
XXMl1_cmp_0 outp outn vss in XMl1_cmp
Xtrim_left_0 trim0 trim4 trim1 trim2 trim3 in trim_left_0/n1 trim_left_0/n4 trim_left_0/n0
+ trim_left_0/n2 trim_left_0/n3 vss trim_left
.ends

.subckt cap_mim_2p0fF_RCWXT2$1 m4_n3120_n3000# m4_n3240_n3120#
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30_flip cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ cap_mim_2p0fF_RCWXT2$1
.ends

.subckt cap_mim_2p0fF_RCWXT2 m4_n3120_n3000# m4_n3240_n3120#
X0 m4_n3120_n3000# m4_n3240_n3120# cap_mim_2f0fF c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30 cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3120_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3240_n3120#
+ cap_mim_2p0fF_RCWXT2
.ends

.subckt mim_cap1 vss vdd
Xmim_cap_30_30_flip_233 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_222 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_200 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_211 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_68 vss vdd mim_cap_30_30
Xmim_cap_30_30_57 vss vdd mim_cap_30_30
Xmim_cap_30_30_79 vss vdd mim_cap_30_30
Xmim_cap_30_30_13 vss vdd mim_cap_30_30
Xmim_cap_30_30_24 vss vdd mim_cap_30_30
Xmim_cap_30_30_46 vss vdd mim_cap_30_30
Xmim_cap_30_30_35 vss vdd mim_cap_30_30
Xmim_cap_30_30_213 vss vdd mim_cap_30_30
Xmim_cap_30_30_224 vss vdd mim_cap_30_30
Xmim_cap_30_30_202 vss vdd mim_cap_30_30
Xmim_cap_30_30_235 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_212 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_234 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_223 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_201 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_58 vss vdd mim_cap_30_30
Xmim_cap_30_30_69 vss vdd mim_cap_30_30
Xmim_cap_30_30_14 vss vdd mim_cap_30_30
Xmim_cap_30_30_25 vss vdd mim_cap_30_30
Xmim_cap_30_30_47 vss vdd mim_cap_30_30
Xmim_cap_30_30_36 vss vdd mim_cap_30_30
Xmim_cap_30_30_214 vss vdd mim_cap_30_30
Xmim_cap_30_30_225 vss vdd mim_cap_30_30
Xmim_cap_30_30_203 vss vdd mim_cap_30_30
Xmim_cap_30_30_236 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_224 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_213 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_235 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_202 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_59 vss vdd mim_cap_30_30
Xmim_cap_30_30_15 vss vdd mim_cap_30_30
Xmim_cap_30_30_48 vss vdd mim_cap_30_30
Xmim_cap_30_30_26 vss vdd mim_cap_30_30
Xmim_cap_30_30_37 vss vdd mim_cap_30_30
Xmim_cap_30_30_226 vss vdd mim_cap_30_30
Xmim_cap_30_30_204 vss vdd mim_cap_30_30
Xmim_cap_30_30_237 vss vdd mim_cap_30_30
Xmim_cap_30_30_215 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_225 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_214 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_236 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_203 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_16 vss vdd mim_cap_30_30
Xmim_cap_30_30_49 vss vdd mim_cap_30_30
Xmim_cap_30_30_38 vss vdd mim_cap_30_30
Xmim_cap_30_30_27 vss vdd mim_cap_30_30
Xmim_cap_30_30_227 vss vdd mim_cap_30_30
Xmim_cap_30_30_238 vss vdd mim_cap_30_30
Xmim_cap_30_30_205 vss vdd mim_cap_30_30
Xmim_cap_30_30_216 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_226 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_215 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_237 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_204 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_17 vss vdd mim_cap_30_30
Xmim_cap_30_30_28 vss vdd mim_cap_30_30
Xmim_cap_30_30_39 vss vdd mim_cap_30_30
Xmim_cap_30_30_228 vss vdd mim_cap_30_30
Xmim_cap_30_30_217 vss vdd mim_cap_30_30
Xmim_cap_30_30_239 vss vdd mim_cap_30_30
Xmim_cap_30_30_206 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_227 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_216 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_238 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_205 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_18 vss vdd mim_cap_30_30
Xmim_cap_30_30_29 vss vdd mim_cap_30_30
Xmim_cap_30_30_229 vss vdd mim_cap_30_30
Xmim_cap_30_30_218 vss vdd mim_cap_30_30
Xmim_cap_30_30_207 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_228 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_217 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_206 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_239 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_19 vss vdd mim_cap_30_30
Xmim_cap_30_30_219 vss vdd mim_cap_30_30
Xmim_cap_30_30_208 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_229 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_218 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_207 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_209 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_219 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_208 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_190 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_209 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_90 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_180 vss vdd mim_cap_30_30
Xmim_cap_30_30_191 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_80 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_91 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_190 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_170 vss vdd mim_cap_30_30
Xmim_cap_30_30_181 vss vdd mim_cap_30_30
Xmim_cap_30_30_192 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_81 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_70 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_92 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_0 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_191 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_180 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_0 vss vdd mim_cap_30_30
Xmim_cap_30_30_160 vss vdd mim_cap_30_30
Xmim_cap_30_30_193 vss vdd mim_cap_30_30
Xmim_cap_30_30_182 vss vdd mim_cap_30_30
Xmim_cap_30_30_171 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_60 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_82 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_71 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_93 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_1 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_170 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_192 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_181 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_1 vss vdd mim_cap_30_30
Xmim_cap_30_30_183 vss vdd mim_cap_30_30
Xmim_cap_30_30_172 vss vdd mim_cap_30_30
Xmim_cap_30_30_150 vss vdd mim_cap_30_30
Xmim_cap_30_30_194 vss vdd mim_cap_30_30
Xmim_cap_30_30_161 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_83 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_72 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_94 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_50 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_61 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_2 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_160 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_193 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_182 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_171 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_2 vss vdd mim_cap_30_30
Xmim_cap_30_30_173 vss vdd mim_cap_30_30
Xmim_cap_30_30_162 vss vdd mim_cap_30_30
Xmim_cap_30_30_184 vss vdd mim_cap_30_30
Xmim_cap_30_30_195 vss vdd mim_cap_30_30
Xmim_cap_30_30_140 vss vdd mim_cap_30_30
Xmim_cap_30_30_151 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_73 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_84 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_95 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_51 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_40 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_62 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_3 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_161 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_172 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_194 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_183 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_150 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_3 vss vdd mim_cap_30_30
Xmim_cap_30_30_174 vss vdd mim_cap_30_30
Xmim_cap_30_30_152 vss vdd mim_cap_30_30
Xmim_cap_30_30_141 vss vdd mim_cap_30_30
Xmim_cap_30_30_196 vss vdd mim_cap_30_30
Xmim_cap_30_30_130 vss vdd mim_cap_30_30
Xmim_cap_30_30_185 vss vdd mim_cap_30_30
Xmim_cap_30_30_163 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_30 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_74 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_85 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_52 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_96 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_41 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_63 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_4 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_151 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_162 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_140 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_173 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_184 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_195 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_4 vss vdd mim_cap_30_30
Xmim_cap_30_30_131 vss vdd mim_cap_30_30
Xmim_cap_30_30_120 vss vdd mim_cap_30_30
Xmim_cap_30_30_153 vss vdd mim_cap_30_30
Xmim_cap_30_30_186 vss vdd mim_cap_30_30
Xmim_cap_30_30_142 vss vdd mim_cap_30_30
Xmim_cap_30_30_197 vss vdd mim_cap_30_30
Xmim_cap_30_30_164 vss vdd mim_cap_30_30
Xmim_cap_30_30_175 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_31 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_75 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_20 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_64 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_86 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_42 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_53 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_97 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_5 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_152 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_163 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_141 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_174 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_130 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_196 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_185 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_5 vss vdd mim_cap_30_30
Xmim_cap_30_30_154 vss vdd mim_cap_30_30
Xmim_cap_30_30_176 vss vdd mim_cap_30_30
Xmim_cap_30_30_165 vss vdd mim_cap_30_30
Xmim_cap_30_30_110 vss vdd mim_cap_30_30
Xmim_cap_30_30_132 vss vdd mim_cap_30_30
Xmim_cap_30_30_121 vss vdd mim_cap_30_30
Xmim_cap_30_30_143 vss vdd mim_cap_30_30
Xmim_cap_30_30_198 vss vdd mim_cap_30_30
Xmim_cap_30_30_187 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_76 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_21 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_65 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_10 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_32 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_43 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_54 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_87 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_98 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_6 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_153 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_164 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_175 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_131 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_142 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_120 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_197 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_186 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_6 vss vdd mim_cap_30_30
Xmim_cap_30_30_155 vss vdd mim_cap_30_30
Xmim_cap_30_30_166 vss vdd mim_cap_30_30
Xmim_cap_30_30_111 vss vdd mim_cap_30_30
Xmim_cap_30_30_100 vss vdd mim_cap_30_30
Xmim_cap_30_30_133 vss vdd mim_cap_30_30
Xmim_cap_30_30_144 vss vdd mim_cap_30_30
Xmim_cap_30_30_122 vss vdd mim_cap_30_30
Xmim_cap_30_30_199 vss vdd mim_cap_30_30
Xmim_cap_30_30_188 vss vdd mim_cap_30_30
Xmim_cap_30_30_177 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_77 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_22 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_66 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_11 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_99 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_33 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_44 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_55 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_88 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_7 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_110 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_121 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_154 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_176 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_143 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_198 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_187 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_132 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_165 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_7 vss vdd mim_cap_30_30
Xmim_cap_30_30_156 vss vdd mim_cap_30_30
Xmim_cap_30_30_167 vss vdd mim_cap_30_30
Xmim_cap_30_30_178 vss vdd mim_cap_30_30
Xmim_cap_30_30_101 vss vdd mim_cap_30_30
Xmim_cap_30_30_112 vss vdd mim_cap_30_30
Xmim_cap_30_30_145 vss vdd mim_cap_30_30
Xmim_cap_30_30_123 vss vdd mim_cap_30_30
Xmim_cap_30_30_189 vss vdd mim_cap_30_30
Xmim_cap_30_30_134 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_23 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_67 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_78 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_12 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_34 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_56 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_45 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_89 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_8 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_100 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_111 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_177 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_188 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_133 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_122 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_199 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_144 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_155 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_166 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_8 vss vdd mim_cap_30_30
Xmim_cap_30_30_168 vss vdd mim_cap_30_30
Xmim_cap_30_30_157 vss vdd mim_cap_30_30
Xmim_cap_30_30_179 vss vdd mim_cap_30_30
Xmim_cap_30_30_102 vss vdd mim_cap_30_30
Xmim_cap_30_30_113 vss vdd mim_cap_30_30
Xmim_cap_30_30_135 vss vdd mim_cap_30_30
Xmim_cap_30_30_146 vss vdd mim_cap_30_30
Xmim_cap_30_30_124 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_68 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_79 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_24 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_13 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_35 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_57 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_46 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_9 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_156 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_145 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_101 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_112 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_123 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_178 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_134 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_189 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_167 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_9 vss vdd mim_cap_30_30
Xmim_cap_30_30_103 vss vdd mim_cap_30_30
Xmim_cap_30_30_114 vss vdd mim_cap_30_30
Xmim_cap_30_30_136 vss vdd mim_cap_30_30
Xmim_cap_30_30_147 vss vdd mim_cap_30_30
Xmim_cap_30_30_125 vss vdd mim_cap_30_30
Xmim_cap_30_30_169 vss vdd mim_cap_30_30
Xmim_cap_30_30_158 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_14 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_69 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_25 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_58 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_36 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_47 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_157 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_168 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_146 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_113 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_102 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_135 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_124 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_179 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_104 vss vdd mim_cap_30_30
Xmim_cap_30_30_115 vss vdd mim_cap_30_30
Xmim_cap_30_30_137 vss vdd mim_cap_30_30
Xmim_cap_30_30_148 vss vdd mim_cap_30_30
Xmim_cap_30_30_126 vss vdd mim_cap_30_30
Xmim_cap_30_30_159 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_15 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_26 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_59 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_37 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_48 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_158 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_147 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_169 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_114 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_103 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_136 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_125 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_105 vss vdd mim_cap_30_30
Xmim_cap_30_30_116 vss vdd mim_cap_30_30
Xmim_cap_30_30_149 vss vdd mim_cap_30_30
Xmim_cap_30_30_138 vss vdd mim_cap_30_30
Xmim_cap_30_30_127 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_16 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_27 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_38 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_49 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_115 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_104 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_137 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_126 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_148 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_159 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_117 vss vdd mim_cap_30_30
Xmim_cap_30_30_106 vss vdd mim_cap_30_30
Xmim_cap_30_30_139 vss vdd mim_cap_30_30
Xmim_cap_30_30_128 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_17 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_28 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_39 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_149 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_116 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_105 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_138 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_127 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_118 vss vdd mim_cap_30_30
Xmim_cap_30_30_107 vss vdd mim_cap_30_30
Xmim_cap_30_30_129 vss vdd mim_cap_30_30
Xmim_cap_30_30_90 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_29 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_18 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_117 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_106 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_139 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_128 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_119 vss vdd mim_cap_30_30
Xmim_cap_30_30_108 vss vdd mim_cap_30_30
Xmim_cap_30_30_80 vss vdd mim_cap_30_30
Xmim_cap_30_30_91 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_19 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_118 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_107 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_129 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_109 vss vdd mim_cap_30_30
Xmim_cap_30_30_70 vss vdd mim_cap_30_30
Xmim_cap_30_30_81 vss vdd mim_cap_30_30
Xmim_cap_30_30_92 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_119 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_108 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_82 vss vdd mim_cap_30_30
Xmim_cap_30_30_60 vss vdd mim_cap_30_30
Xmim_cap_30_30_71 vss vdd mim_cap_30_30
Xmim_cap_30_30_93 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_109 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_50 vss vdd mim_cap_30_30
Xmim_cap_30_30_83 vss vdd mim_cap_30_30
Xmim_cap_30_30_72 vss vdd mim_cap_30_30
Xmim_cap_30_30_61 vss vdd mim_cap_30_30
Xmim_cap_30_30_94 vss vdd mim_cap_30_30
Xmim_cap_30_30_73 vss vdd mim_cap_30_30
Xmim_cap_30_30_84 vss vdd mim_cap_30_30
Xmim_cap_30_30_62 vss vdd mim_cap_30_30
Xmim_cap_30_30_95 vss vdd mim_cap_30_30
Xmim_cap_30_30_51 vss vdd mim_cap_30_30
Xmim_cap_30_30_40 vss vdd mim_cap_30_30
Xmim_cap_30_30_74 vss vdd mim_cap_30_30
Xmim_cap_30_30_52 vss vdd mim_cap_30_30
Xmim_cap_30_30_85 vss vdd mim_cap_30_30
Xmim_cap_30_30_63 vss vdd mim_cap_30_30
Xmim_cap_30_30_96 vss vdd mim_cap_30_30
Xmim_cap_30_30_30 vss vdd mim_cap_30_30
Xmim_cap_30_30_41 vss vdd mim_cap_30_30
Xmim_cap_30_30_230 vss vdd mim_cap_30_30
Xmim_cap_30_30_75 vss vdd mim_cap_30_30
Xmim_cap_30_30_20 vss vdd mim_cap_30_30
Xmim_cap_30_30_64 vss vdd mim_cap_30_30
Xmim_cap_30_30_86 vss vdd mim_cap_30_30
Xmim_cap_30_30_53 vss vdd mim_cap_30_30
Xmim_cap_30_30_31 vss vdd mim_cap_30_30
Xmim_cap_30_30_42 vss vdd mim_cap_30_30
Xmim_cap_30_30_97 vss vdd mim_cap_30_30
Xmim_cap_30_30_220 vss vdd mim_cap_30_30
Xmim_cap_30_30_231 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_230 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_65 vss vdd mim_cap_30_30
Xmim_cap_30_30_76 vss vdd mim_cap_30_30
Xmim_cap_30_30_10 vss vdd mim_cap_30_30
Xmim_cap_30_30_54 vss vdd mim_cap_30_30
Xmim_cap_30_30_21 vss vdd mim_cap_30_30
Xmim_cap_30_30_87 vss vdd mim_cap_30_30
Xmim_cap_30_30_32 vss vdd mim_cap_30_30
Xmim_cap_30_30_43 vss vdd mim_cap_30_30
Xmim_cap_30_30_98 vss vdd mim_cap_30_30
Xmim_cap_30_30_221 vss vdd mim_cap_30_30
Xmim_cap_30_30_232 vss vdd mim_cap_30_30
Xmim_cap_30_30_210 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_231 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_220 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_66 vss vdd mim_cap_30_30
Xmim_cap_30_30_77 vss vdd mim_cap_30_30
Xmim_cap_30_30_11 vss vdd mim_cap_30_30
Xmim_cap_30_30_22 vss vdd mim_cap_30_30
Xmim_cap_30_30_88 vss vdd mim_cap_30_30
Xmim_cap_30_30_44 vss vdd mim_cap_30_30
Xmim_cap_30_30_99 vss vdd mim_cap_30_30
Xmim_cap_30_30_33 vss vdd mim_cap_30_30
Xmim_cap_30_30_55 vss vdd mim_cap_30_30
Xmim_cap_30_30_222 vss vdd mim_cap_30_30
Xmim_cap_30_30_233 vss vdd mim_cap_30_30
Xmim_cap_30_30_200 vss vdd mim_cap_30_30
Xmim_cap_30_30_211 vss vdd mim_cap_30_30
Xmim_cap_30_30_flip_232 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_221 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_flip_210 vss vdd mim_cap_30_30_flip
Xmim_cap_30_30_67 vss vdd mim_cap_30_30
Xmim_cap_30_30_12 vss vdd mim_cap_30_30
Xmim_cap_30_30_23 vss vdd mim_cap_30_30
Xmim_cap_30_30_56 vss vdd mim_cap_30_30
Xmim_cap_30_30_78 vss vdd mim_cap_30_30
Xmim_cap_30_30_89 vss vdd mim_cap_30_30
Xmim_cap_30_30_45 vss vdd mim_cap_30_30
Xmim_cap_30_30_34 vss vdd mim_cap_30_30
Xmim_cap_30_30_212 vss vdd mim_cap_30_30
Xmim_cap_30_30_234 vss vdd mim_cap_30_30
Xmim_cap_30_30_223 vss vdd mim_cap_30_30
Xmim_cap_30_30_201 vss vdd mim_cap_30_30
.ends

.subckt cap_mim_2p0fF_DMYL6H m4_n114303_n17580# m4_n114183_n17460#
X0 m4_n114183_n17460# m4_n114303_n17580# cap_mim_2f0fF c_width=100u c_length=100u
.ends

.subckt mim_cap_100_100 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_n114303_n17580# cap_mim_2p0fF_DMYL6H_0/m4_n114183_n17460#
+ cap_mim_2p0fF_DMYL6H
.ends

.subckt cap_mim_2p0fF_RCWXT2$2 m4_n3148_n3000# m4_n3268_n3120#
X0 m4_n3148_n3000# m4_n3268_n3120# cap_mim_2f0fF c_width=30u c_length=30u
.ends

.subckt mim_cap_30_30$1 cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120# cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000#
Xcap_mim_2p0fF_RCWXT2_0 cap_mim_2p0fF_RCWXT2_0/m4_n3148_n3000# cap_mim_2p0fF_RCWXT2_0/m4_n3268_n3120#
+ cap_mim_2p0fF_RCWXT2$2
.ends

.subckt cap_mim_2p0fF_DMYL6H$1 m4_93823_n2660# m4_93943_n2540#
X0 m4_93943_n2540# m4_93823_n2660# cap_mim_2f0fF c_width=100u c_length=100u
.ends

.subckt mim_cap_100_100$1 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
Xcap_mim_2p0fF_DMYL6H_0 cap_mim_2p0fF_DMYL6H_0/m4_93823_n2660# cap_mim_2p0fF_DMYL6H_0/m4_93943_n2540#
+ cap_mim_2p0fF_DMYL6H$1
.ends

.subckt mim_cap2 vss vdd
Xmim_cap_100_100_1 vss vdd mim_cap_100_100
Xmim_cap_100_100_0 vss vdd mim_cap_100_100
Xmim_cap_100_100_2 vss vdd mim_cap_100_100
Xmim_cap_100_100_3 vss vdd mim_cap_100_100
Xmim_cap_30_30$1_20 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_0 vss vdd mim_cap_30_30$1
Xmim_cap_100_100_4 vss vdd mim_cap_100_100
Xmim_cap_30_30$1_22 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_21 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_11 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_10 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_1 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_23 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_12 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_2 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_24 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_13 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_3 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_14 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_4 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_15 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_6 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_5 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_16 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_7 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_17 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_8 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_18 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_9 vss vdd mim_cap_30_30$1
Xmim_cap_30_30$1_19 vss vdd mim_cap_30_30$1
Xmim_cap_100_100$1_0 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_1 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_2 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_4 vss vdd mim_cap_100_100$1
Xmim_cap_100_100$1_3 vss vdd mim_cap_100_100$1
.ends

.subckt mim_cap_boss vdd vdd_uq0 vss
Xmim_cap1_0 vss vdd mim_cap1
Xmim_cap2_0 vss vdd_uq0 mim_cap2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VPW VNW
MX0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VPW VNW
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.205p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.205p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VPW VNW
MX0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
MX1 VSS RN a_1456_156# VPW nfet_06v0 ad=0.202p pd=1.48u as=43.2f ps=0.6u w=0.36u l=0.6u
MX2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.535p pd=3.31u as=0.535p ps=3.31u w=1.22u l=0.5u
MX3 a_796_472# D VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX4 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.122p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
MX5 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
MX6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.203p pd=1.3u as=0.203p ps=1.3u w=0.78u l=0.5u
MX7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.254p pd=1.51u as=0.242p ps=1.46u w=0.505u l=0.5u
MX8 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.201p pd=1.48u as=0.201p ps=1.48u w=0.36u l=0.6u
MX9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
MX10 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.2f pd=0.6u as=43.2f ps=0.6u w=0.36u l=0.6u
MX11 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.201p pd=1.48u as=0.202p ps=1.48u w=0.36u l=0.6u
MX12 Q a_2665_112# VSS VPW nfet_06v0 ad=0.359p pd=2.51u as=0.359p ps=2.51u w=0.815u l=0.6u
MX13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
MX14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.203p pd=1.3u as=0.203p ps=1.3u w=0.78u l=0.5u
MX15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.343p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
MX16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.295p ps=1.74u w=1u l=0.5u
MX17 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.201p ps=1.48u w=0.36u l=0.6u
MX18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
MX19 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
MX20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.203p ps=1.3u w=0.78u l=0.5u
MX21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.131p pd=1.02u as=0.254p ps=1.51u w=0.505u l=0.5u
MX22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
MX23 a_3041_156# RN VSS VPW nfet_06v0 ad=0.134p pd=1.1u as=0.122p ps=1.04u w=0.36u l=0.6u
MX24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.295p pd=1.74u as=0.131p ps=1.02u w=0.505u l=0.5u
MX25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.242p pd=1.46u as=0.222p ps=1.89u w=0.505u l=0.5u
MX26 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
MX27 a_796_472# D VDD VNW pfet_06v0 ad=0.203p pd=1.3u as=0.343p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
MX1 VSS A1 ZN VPW nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
MX2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.409p pd=1.89u as=0.537p ps=3.32u w=1.22u l=0.5u
MX3 ZN A2 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VPW VNW
MX0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
MX1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
MX2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.659p ps=3.52u w=1.22u l=0.5u
MX3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.378p ps=1.84u w=1.22u l=0.5u
MX4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
MX5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
MX6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
MX7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.13p ps=1.13u w=0.815u l=0.6u
MX1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
MX2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
MX3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
MX4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
MX5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.13p pd=1.13u as=0.359p ps=2.51u w=0.815u l=0.6u
MX6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.13p pd=1.13u as=0.212p ps=1.34u w=0.815u l=0.6u
MX7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.359p pd=2.51u as=0.13p ps=1.13u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VPW VNW
MX0 Z a_36_160# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.234p ps=1.56u w=0.82u l=0.6u
MX1 Z a_36_160# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.353p ps=1.96u w=1.22u l=0.5u
MX2 VDD I a_36_160# VNW pfet_06v0 ad=0.353p pd=1.96u as=0.249p ps=2.01u w=0.565u l=0.5u
MX3 VSS I a_36_160# VPW nfet_06v0 ad=0.234p pd=1.56u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VPW VNW
MX0 ZN I VSS VPW nfet_06v0 ad=0.211p pd=1.84u as=0.211p ps=1.84u w=0.48u l=0.6u
MX1 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VPW VNW
MX0 ZN I VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=0.6u
MX1 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VPW VNW
MX0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VPW VNW
MX0 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u M=4
MX1 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u M=8
MX2 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u M=4
MX3 VSS a_224_472# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u M=8
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VPW VNW
MX0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
MX1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.257p pd=1.56u as=0.131p ps=1.14u w=0.82u l=0.6u
MX2 VDD B a_36_472# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.45p ps=1.96u w=1.22u l=0.5u
MX3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
MX4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.45p pd=1.96u as=0.316p ps=1.74u w=1.22u l=0.5u
MX5 VSS B ZN VPW nfet_06v0 ad=0.224p pd=1.9u as=0.257p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VPW VNW
MX0 VDD I a_36_113# VNW pfet_06v0 ad=0.401p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
MX1 Z a_36_113# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.401p ps=1.92u w=1.22u l=0.5u
MX2 Z a_36_113# VSS VPW nfet_06v0 ad=0.218p pd=1.87u as=0.153p ps=1.19u w=0.495u l=0.6u
MX3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.19u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
MX1 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
MX2 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
MX3 ZN A1 VDD VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
MX4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
MX5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VPW VNW
MX0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u
MX1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
MX2 VDD A1 ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.294p ps=1.65u w=1.13u l=0.5u
MX3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VPW VNW
MX0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.5u
MX1 Z a_67_603# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.229p ps=1.58u w=0.82u l=0.6u
MX2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.387p pd=2.08u as=0.147p ps=1.09u w=0.565u l=0.5u
MX3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.229p pd=1.58u as=93.6f ps=0.88u w=0.36u l=0.6u
MX4 Z a_67_603# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.387p ps=2.08u w=1.22u l=0.5u
MX5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VPW VNW
MX0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.377p pd=1.81u as=0.46p ps=1.93u w=1.1u l=0.5u
MX1 VDD C ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u M=4
MX2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u M=4
MX3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
MX4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
MX5 a_2124_68# B a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
MX6 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.361p ps=2.52u w=0.82u l=0.6u M=4
MX7 VSS C a_2960_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
MX8 VDD B ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u M=4
MX9 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
MX10 a_36_68# B a_3368_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
MX11 a_244_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.482p ps=3.07u w=1.1u l=0.5u
MX12 VSS C a_2124_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX13 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
MX14 a_36_68# B a_2552_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
MX15 a_2552_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX16 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
MX17 a_3368_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX18 a_2960_68# B a_36_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX19 ZN A1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VPW VNW
MX0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.449p ps=2.92u w=1.02u l=0.5u
MX1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.18u as=0.158p ps=1.6u w=0.36u l=0.6u
MX2 VDD a_36_160# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u M=2
MX3 VSS a_36_160# Z VPW nfet_06v0 ad=0.213p pd=1.85u as=0.126p ps=1u w=0.485u l=0.6u M=2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VPW VNW
MX0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
MX4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
MX7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VPW VNW
MX0 Z a_36_68# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.494p ps=2.03u w=1.22u l=0.5u M=2
MX1 VSS I a_36_68# VPW nfet_06v0 ad=0.291p pd=1.53u as=0.361p ps=2.52u w=0.82u l=0.6u
MX2 Z a_36_68# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.291p ps=1.53u w=0.82u l=0.6u M=2
MX3 VDD I a_36_68# VNW pfet_06v0 ad=0.494p pd=2.03u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VPW VNW
MX0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.146p pd=1.46u as=0.317p ps=1.74u w=1.22u l=0.5u
MX1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
MX2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
MX3 Z a_124_24# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u M=2
MX4 a_848_380# S VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
MX5 VDD a_124_24# Z VNW pfet_06v0 ad=0.439p pd=1.94u as=0.348p ps=1.79u w=1.22u l=0.5u M=2
MX6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.146p ps=1.46u w=1.22u l=0.5u
MX7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.476p pd=2u as=0.439p ps=1.94u w=1.22u l=0.5u
MX8 a_848_380# S VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
MX9 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.197p ps=1.3u w=0.82u l=0.6u
MX10 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.197p pd=1.3u as=0.213p ps=1.34u w=0.82u l=0.6u
MX11 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.476p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VPW VNW
MX0 VSS B a_36_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
MX1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
MX2 VDD B ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.425p ps=1.94u w=1.13u l=0.5u
MX3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
MX4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.425p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
MX5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VPW VNW
MX0 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u M=4
MX1 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u M=2
MX2 VSS a_224_552# Z VPW nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u M=4
MX3 a_224_552# I VSS VPW nfet_06v0 ad=0.514p pd=2.91u as=0.266p ps=2.09u w=0.605u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VPW VNW
MX0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.409p pd=1.89u as=0.348p ps=1.79u w=1.22u l=0.5u
MX1 ZN A1 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u M=2
MX2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
MX3 a_234_472# A2 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
MX4 VDD A2 a_672_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
MX5 VSS A2 ZN VPW nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u M=2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
MX1 ZN A1 VSS VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
MX2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
MX3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.317p ps=1.74u w=1.22u l=0.5u
MX4 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
MX5 ZN A3 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 VDD A1 ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.522p ps=2.05u w=0.985u l=0.5u M=4
MX1 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.416p ps=1.9u w=0.82u l=0.6u M=3
MX2 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.305p ps=1.61u w=0.985u l=0.5u M=4
MX3 a_36_68# A2 a_672_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX4 a_1732_68# A2 a_1528_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.172p ps=1.24u w=0.82u l=0.6u
MX5 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.305p ps=1.61u w=0.985u l=0.5u M=4
MX6 a_244_68# A2 a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.361p ps=2.52u w=0.82u l=0.6u
MX7 a_1528_68# A3 VSS VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
MX8 a_1100_68# A2 a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
MX9 ZN A1 a_1732_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.172p ps=1.24u w=0.82u l=0.6u
MX10 VSS A3 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX11 VSS A3 a_1100_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX12 a_672_68# A3 VSS VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VPW VNW
MX0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.406p pd=2.05u as=0.156p ps=1.12u w=0.6u l=0.5u
MX1 Z a_36_159# VDD VNW pfet_06v0 ad=0.535p pd=3.31u as=0.406p ps=2.05u w=1.22u l=0.5u
MX2 Z a_36_159# VSS VPW nfet_06v0 ad=0.359p pd=2.51u as=0.234p ps=1.55u w=0.815u l=0.6u
MX3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.234p pd=1.55u as=58.4f ps=0.685u w=0.365u l=0.6u
MX4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.4f pd=0.685u as=0.161p ps=1.61u w=0.365u l=0.6u
MX5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VPW VNW
MX0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.598p pd=3.42u as=0.317p ps=1.74u w=1.22u l=0.5u
MX1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
MX2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
MX3 VSS C ZN VPW nfet_06v0 ad=0.254p pd=1.61u as=0.12p ps=0.98u w=0.46u l=0.6u M=4
MX4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u M=4
MX5 ZN B VSS VPW nfet_06v0 ad=0.12p pd=0.98u as=0.238p ps=1.51u w=0.46u l=0.6u M=4
MX6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
MX7 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.162p ps=1.19u w=0.77u l=0.6u
MX8 VDD C a_3126_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.317p ps=1.74u w=1.22u l=0.5u
MX9 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.238p pd=1.51u as=0.123p ps=1.09u w=0.77u l=0.6u
MX10 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
MX11 a_170_472# A2 ZN VNW pfet_06v0 ad=0.451p pd=1.96u as=0.317p ps=1.74u w=1.22u l=0.5u M=4
MX12 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.451p ps=1.96u w=1.22u l=0.5u
MX13 a_2590_472# C VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
MX14 a_358_69# A2 VSS VPW nfet_06v0 ad=0.162p pd=1.19u as=0.447p ps=2.7u w=0.77u l=0.6u
MX15 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
MX16 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.317p ps=1.74u w=1.22u l=0.5u
MX17 VDD C a_2034_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.378p ps=1.84u w=1.22u l=0.5u
MX18 a_786_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
MX19 a_3662_472# C VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u M=3
MX2 ZN A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u M=4
MX3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX5 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u M=4
MX6 VSS A3 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u M=4
MX7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX8 VDD A3 a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX9 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX10 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX11 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX12 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.348p ps=1.79u w=1.22u l=0.5u
MX1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
MX2 ZN A3 VSS VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u M=2
MX3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
MX4 ZN A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u M=2
MX5 ZN A2 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u M=2
MX6 a_906_472# A1 ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
MX7 ZN A1 a_468_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
MX8 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VPW VNW
MX0 VSS B ZN VPW nfet_06v0 ad=0.227p pd=1.91u as=0.134p ps=1.03u w=0.515u l=0.6u M=2
MX1 VSS C ZN VPW nfet_06v0 ad=0.134p pd=1.03u as=0.134p ps=1.03u w=0.515u l=0.6u M=2
MX2 a_244_68# A2 VSS VPW nfet_06v0 ad=93.6f pd=1.02u as=0.343p ps=2.44u w=0.78u l=0.6u
MX3 ZN A1 a_244_68# VPW nfet_06v0 ad=0.203p pd=1.3u as=93.6f ps=1.02u w=0.78u l=0.6u
MX4 VDD C a_1044_488# VNW pfet_06v0 ad=0.353p pd=1.76u as=0.353p ps=1.76u w=1.14u l=0.5u
MX5 ZN A1 a_36_488# VNW pfet_06v0 ad=0.296p pd=1.66u as=0.308p ps=1.68u w=1.14u l=0.5u M=2
MX6 ZN A2 a_36_488# VNW pfet_06v0 ad=0.296p pd=1.66u as=0.502p ps=3.16u w=1.14u l=0.5u M=2
MX7 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.353p pd=1.76u as=0.296p ps=1.66u w=1.14u l=0.5u
MX8 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.502p pd=3.16u as=0.353p ps=1.76u w=1.14u l=0.5u
MX9 a_636_68# A1 ZN VPW nfet_06v0 ad=93.6f pd=1.02u as=0.203p ps=1.3u w=0.78u l=0.6u
MX10 a_1492_488# C VDD VNW pfet_06v0 ad=0.353p pd=1.76u as=0.353p ps=1.76u w=1.14u l=0.5u
MX11 VSS A2 a_636_68# VPW nfet_06v0 ad=0.233p pd=1.48u as=93.6f ps=1.02u w=0.78u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VPW VNW
MX0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=93.6f ps=0.88u w=0.36u l=0.6u
MX1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.161p ps=1.13u w=0.565u l=0.5u
MX2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.249p ps=2.01u w=0.565u l=0.5u
MX3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.5u
MX4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161p pd=1.13u as=0.194p ps=1.41u w=0.565u l=0.5u
MX5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.5u
MX6 VSS A1 a_56_524# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
MX7 a_1336_472# a_728_93# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.41u as=93.6f ps=0.88u w=0.36u l=0.5u
MX9 a_56_524# A2 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX10 VSS A3 a_1336_472# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.6f ps=0.88u w=0.36u l=0.6u
MX11 a_2215_68# A3 Z VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX12 VSS a_728_93# a_2215_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
MX13 Z a_1336_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
MX14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
MX15 a_728_93# a_56_524# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
MX16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
MX17 VSS A2 a_952_93# VPW nfet_06v0 ad=0.158p pd=1.6u as=57.6f ps=0.68u w=0.36u l=0.6u
MX18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.353p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
MX19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.353p ps=1.96u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VPW VNW
MX0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
MX1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
MX2 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u M=2
MX3 VDD A1 ZN VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u M=2
MX4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VPW VNW
MX0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
MX1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.339p pd=1.71u as=0.46p ps=1.93u w=1.1u l=0.5u
MX2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u M=2
MX3 VSS B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u M=2
MX4 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u M=2
MX5 ZN B VDD VNW pfet_06v0 ad=0.281p pd=1.6u as=0.529p ps=3.14u w=1.08u l=0.5u M=2
MX6 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u M=2
MX7 a_692_497# A3 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.392p ps=1.81u w=1.1u l=0.5u
MX8 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.46p pd=1.93u as=0.339p ps=1.71u w=1.1u l=0.5u
MX9 ZN A1 a_960_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.339p ps=1.71u w=1.1u l=0.5u
MX10 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VPW VNW
MX0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
MX1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u M=2
MX2 VSS RN a_1456_156# VPW nfet_06v0 ad=0.202p pd=1.48u as=43.2f ps=0.6u w=0.36u l=0.6u
MX3 a_796_472# D VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX4 VSS a_2665_112# a_2560_156# VPW nfet_06v0 ad=0.122p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
MX5 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.203p pd=1.3u as=0.203p ps=1.3u w=0.78u l=0.5u
MX6 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.254p pd=1.51u as=0.242p ps=1.46u w=0.505u l=0.5u
MX7 a_2248_156# a_448_472# a_1308_423# VPW nfet_06v0 ad=0.201p pd=1.48u as=0.201p ps=1.48u w=0.36u l=0.6u
MX8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
MX9 a_1456_156# a_1308_423# a_1288_156# VPW nfet_06v0 ad=43.2f pd=0.6u as=43.2f ps=0.6u w=0.36u l=0.6u
MX10 a_1308_423# a_1000_472# VSS VPW nfet_06v0 ad=0.201p pd=1.48u as=0.202p ps=1.48u w=0.36u l=0.6u
MX11 Q a_2665_112# VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.359p ps=2.51u w=0.815u l=0.6u M=2
MX12 a_2665_112# a_2248_156# a_3041_156# VPW nfet_06v0 ad=0.359p pd=2.51u as=0.217p ps=1.51u w=0.815u l=0.6u
MX13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
MX14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.203p pd=1.3u as=0.203p ps=1.3u w=0.78u l=0.5u
MX15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.343p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
MX16 a_2560_156# a_36_151# a_2248_156# VPW nfet_06v0 ad=94.5f pd=0.885u as=0.201p ps=1.48u w=0.36u l=0.6u
MX17 a_1288_156# a_448_472# a_1000_472# VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
MX18 a_2665_112# RN VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.338p ps=1.96u w=1.22u l=0.5u
MX19 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.203p ps=1.3u w=0.78u l=0.5u
MX20 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.131p pd=1.02u as=0.254p ps=1.51u w=0.505u l=0.5u
MX21 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
MX22 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
MX23 a_3041_156# RN VSS VPW nfet_06v0 ad=0.217p pd=1.51u as=0.122p ps=1.04u w=0.36u l=0.6u
MX24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.338p pd=1.96u as=0.131p ps=1.02u w=0.505u l=0.5u
MX25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.242p pd=1.46u as=0.222p ps=1.89u w=0.505u l=0.5u
MX26 a_1000_472# a_36_151# a_796_472# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
MX27 a_796_472# D VDD VNW pfet_06v0 ad=0.203p pd=1.3u as=0.343p ps=2.44u w=0.78u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VPW VNW
MX0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.172p ps=1.24u w=0.82u l=0.6u
MX1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
MX2 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.372p ps=2.57u w=0.845u l=0.5u M=2
MX3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.152p pd=1.19u as=0.361p ps=2.52u w=0.82u l=0.6u
MX4 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u M=2
MX5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.152p ps=1.19u w=0.82u l=0.6u
MX6 VDD A2 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u M=2
MX7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX8 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u M=2
MX9 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.152p pd=1.19u as=0.213p ps=1.34u w=0.82u l=0.6u
MX10 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
MX11 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.152p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VPW VNW
MX0 ZN I VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u M=2
MX1 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u M=2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
MX1 a_244_68# A1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
MX2 a_244_68# A3 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
MX3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
MX4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
MX5 ZN B1 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
MX6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
MX7 VSS A2 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
MX8 a_244_68# B2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
MX9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=93.6f ps=0.88u w=0.36u l=0.6u
MX1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.103p pd=0.93u as=0.158p ps=1.6u w=0.36u l=0.5u
MX2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.146p pd=1.08u as=0.16p ps=1.13u w=0.56u l=0.5u
MX3 ZN A3 a_1948_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.213p ps=1.34u w=0.82u l=0.6u
MX4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.339p pd=1.71u as=0.352p ps=1.89u w=1.1u l=0.5u
MX5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.526p ps=2.05u w=1.1u l=0.5u
MX6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.16p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
MX7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.246p pd=2u as=0.146p ps=1.08u w=0.56u l=0.5u
MX8 VSS A1 a_56_567# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
MX9 VSS A3 a_1504_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.6f ps=0.68u w=0.36u l=0.6u
MX10 a_1948_68# a_728_93# ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.416p ps=1.9u w=0.82u l=0.6u
MX11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.526p pd=2.05u as=0.339p ps=1.71u w=1.1u l=0.5u
MX12 a_1504_93# a_728_93# a_1296_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=0.158p ps=1.6u w=0.36u l=0.6u
MX13 a_56_567# A2 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX14 a_1948_68# a_1296_93# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
MX15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.146p pd=1.08u as=0.246p ps=2u w=0.56u l=0.5u
MX16 a_728_93# a_56_567# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
MX17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352p pd=1.89u as=0.146p ps=1.08u w=0.56u l=0.5u
MX18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.103p ps=0.93u w=0.36u l=0.5u
MX19 VSS A2 a_952_93# VPW nfet_06v0 ad=0.158p pd=1.6u as=57.6f ps=0.68u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VPW VNW
MX0 a_1229_68# B a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.215p ps=1.35u w=0.82u l=0.6u
MX1 VDD B ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u M=2
MX2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u M=2
MX3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
MX4 a_36_68# B a_1657_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
MX5 ZN A2 a_36_68# VPW nfet_06v0 ad=0.312p pd=1.68u as=0.361p ps=2.52u w=0.82u l=0.6u M=2
MX6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.379p pd=1.82u as=0.46p ps=1.93u w=1.1u l=0.5u
MX7 a_244_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.482p ps=3.07u w=1.1u l=0.5u
MX8 a_1657_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX9 VDD C ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u M=2
MX10 VSS C a_1229_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
MX11 ZN A1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VPW VNW
MX0 Z a_36_148# VDD VNW pfet_06v0 ad=0.535p pd=3.31u as=0.427p ps=2.17u w=1.22u l=0.5u
MX1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.8f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
MX2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.242p ps=1.63u w=0.775u l=0.6u
MX3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.242p pd=1.63u as=79.8f ps=0.8u w=0.38u l=0.6u
MX4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.167p ps=1.64u w=0.38u l=0.6u
MX5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.139p pd=1.05u as=0.235p ps=1.95u w=0.535u l=0.5u
MX6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.139p pd=1.05u as=0.139p ps=1.05u w=0.535u l=0.5u
MX7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.427p pd=2.17u as=0.139p ps=1.05u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VPW VNW
MX0 ZN A1 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u M=2
MX1 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
MX2 a_860_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
MX3 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u M=2
MX4 VDD A3 ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u M=2
MX5 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
MX6 a_276_68# A3 VSS VPW nfet_06v0 ad=0.115p pd=1.1u as=0.361p ps=2.52u w=0.82u l=0.6u
MX7 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.115p ps=1.1u w=0.82u l=0.6u
MX8 ZN A1 a_452_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VPW VNW
MX0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX1 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u M=4
MX2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.456p pd=1.96u as=0.486p ps=2.02u w=1.22u l=0.5u
MX5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.486p ps=2.02u w=1.22u l=0.5u
MX6 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX7 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.456p ps=1.96u w=1.22u l=0.5u
MX8 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX9 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u M=4
MX10 VDD A4 a_254_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.346p ps=1.78u w=1.22u l=0.5u
MX11 VSS A4 ZN VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u M=4
MX12 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u M=4
MX13 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
MX14 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX15 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346p pd=1.78u as=0.535p ps=3.31u w=1.22u l=0.5u
MX16 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
MX17 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.377p ps=1.83u w=1.22u l=0.5u
MX18 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
MX19 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VPW VNW
MX0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=93f ps=1.01u w=0.775u l=0.6u
MX1 VDD B a_49_472# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.535p ps=3.31u w=1.22u l=0.5u M=2
MX2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.328p ps=1.75u w=1.22u l=0.5u M=2
MX3 a_741_69# A2 VSS VPW nfet_06v0 ad=93f pd=1.01u as=0.24p ps=1.48u w=0.775u l=0.6u
MX4 ZN B VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u M=2
MX5 a_49_472# A2 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u M=2
MX6 ZN A1 a_741_69# VPW nfet_06v0 ad=0.201p pd=1.29u as=93f ps=1.01u w=0.775u l=0.6u
MX7 a_1133_69# A1 ZN VPW nfet_06v0 ad=93f pd=1.01u as=0.201p ps=1.29u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VPW VNW
MX0 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.457p ps=1.97u w=1.22u l=0.5u M=2
MX1 ZN I VSS VPW nfet_06v0 ad=0.225p pd=1.37u as=0.361p ps=2.52u w=0.82u l=0.6u M=2
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VPW VNW
MX0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
MX1 a_1353_112# SETN a_1697_156# VPW nfet_06v0 ad=0.199p pd=1.46u as=86.4f ps=0.84u w=0.36u l=0.6u
MX2 a_836_156# D VDD VNW pfet_06v0 ad=0.131p pd=1.02u as=0.227p ps=1.91u w=0.505u l=0.5u
MX3 a_1040_527# a_36_151# a_836_156# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
MX4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.193p pd=1.27u as=0.131p ps=1.02u w=0.505u l=0.5u
MX5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.108p pd=0.935u as=0.278p ps=2.17u w=0.415u l=0.5u
MX6 VSS a_1353_112# a_1284_156# VPW nfet_06v0 ad=93.6f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
MX7 a_2225_156# a_448_472# a_1353_112# VPW nfet_06v0 ad=93.6f pd=0.88u as=0.199p ps=1.46u w=0.36u l=0.6u
MX8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
MX9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.183p pd=1.71u as=0.108p ps=0.935u w=0.415u l=0.5u
MX10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.328p pd=1.62u as=0.203p ps=1.3u w=0.78u l=0.5u
MX11 Q a_3129_107# VSS VPW nfet_06v0 ad=0.359p pd=2.51u as=0.359p ps=2.51u w=0.815u l=0.6u
MX12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
MX13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.203p pd=1.3u as=0.343p ps=2.44u w=0.78u l=0.5u
MX14 VSS a_3129_107# a_3081_151# VPW nfet_06v0 ad=0.15p pd=1.14u as=48.6f ps=0.645u w=0.405u l=0.6u
MX15 a_836_156# D VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
MX16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
MX17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.152p pd=1.11u as=0.397p ps=2.18u w=0.585u l=0.5u
MX18 a_3129_107# a_2225_156# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.15p ps=1.14u w=0.405u l=0.6u
MX19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.415p pd=2.65u as=0.152p ps=1.11u w=0.585u l=0.5u
MX20 a_1284_156# a_448_472# a_1040_527# VPW nfet_06v0 ad=62.1f pd=0.705u as=93.6f ps=0.88u w=0.36u l=0.6u
MX21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.397p pd=2.18u as=0.101p ps=0.905u w=0.505u l=0.5u
MX22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.656p pd=3.51u as=0.535p ps=3.31u w=1.22u l=0.5u
MX23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.343p pd=2.44u as=0.328p ps=1.62u w=0.78u l=0.5u
MX24 a_2449_156# a_36_151# a_2225_156# VPW nfet_06v0 ad=0.29p pd=2.33u as=93.6f ps=0.88u w=0.36u l=0.6u
MX25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.193p ps=1.27u w=0.505u l=0.5u
MX26 a_1697_156# a_1040_527# VSS VPW nfet_06v0 ad=86.4f pd=0.84u as=93.6f ps=0.88u w=0.36u l=0.6u
MX27 a_3081_151# SETN a_2449_156# VPW nfet_06v0 ad=48.6f pd=0.645u as=0.312p ps=2.38u w=0.405u l=0.6u
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctln[8]
+ ctln[9] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8]
+ ctlp[9] cal clk clkc comp en result[0] result[1] result[2] result[3] result[4] result[5]
+ result[6] result[7] result[8] result[9] rstn sample trim[0] trim[1] trim[2] trim[3]
+ trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] valid vdd vss
XFILLER_0_17_200 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_432_ _021_ mask\[3\] net63 vss net80 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_294_ vdd vss _008_ _104_ _106_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput7 ctln[0] net7 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
X_431_ _020_ mask\[2\] net53 vss net70 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_293_ net31 vdd vss _106_ mask\[4\] _105_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_362_ vdd vss trim_mask\[1\] _155_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_276_ vss _093_ _092_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_345_ vss _144_ _132_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_204 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _078_ vdd vss _080_ _073_ _076_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout79_I vss net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__358__I vss _053_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_430_ _019_ mask\[1\] net63 vss net80 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_292_ vss _105_ _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_361_ vdd vss _154_ _086_ _119_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_344_ vdd vss _143_ _021_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__191__I vss net17 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_96 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_327_ _131_ vdd vss _016_ _127_ _130_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_189_ vdd vss _043_ net27 mask\[0\] vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_258_ vss _079_ _078_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput33 result[6] net33 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput22 ctlp[5] net22 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__292__I vss _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_257_ _077_ vdd vss _078_ _053_ _075_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_326_ _131_ vss vdd _125_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_309_ vss _116_ net4 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__301__A2 vss _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 ctlp[6] net23 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_273_ vss _090_ state\[0\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
X_342_ vdd vss _142_ _020_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout80 vss net80 net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_325_ vdd vss _130_ _118_ _129_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_98 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ vss vdd gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_124 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 ctln[6] net13 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput24 ctlp[7] net24 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_272_ _089_ vdd vss _003_ _079_ _087_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_410_ vdd _188_ _187_ _042_ _120_ vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout81 vss net81 net82 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_255_ _076_ vss vdd _057_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output40_I vss net40 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_324_ vdd vss _129_ calibrate _062_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout70 vss net70 net73 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__304__A1 vss _093_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_55 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_307_ vdd vss _114_ _113_ _096_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput36 result[9] net36 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 ctlp[8] net25 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__200__I vss net20 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_99 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout60 net60 vss vdd net61 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout71 vss net71 net73 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_323_ vss _015_ _128_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_306_ vss _113_ _057_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
X_237_ vdd vss net40 net45 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_57 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ vss vdd gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_10_37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net50 vss vdd net52 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_305_ vdd vss _112_ net1 _081_ vss vdd gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ net40 vss vdd _064_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vss net22 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_214 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__209__I vss net23 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_91 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_output19_I vss net19 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_252_ vdd vss cal_itt\[0\] _073_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout62 net62 vss vdd net64 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vss net51 net52 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout73 vss net73 net74 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_100 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xfanout63 net63 vss vdd net64 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout52 net52 vss vdd net57 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout74 vss net74 net82 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_449_ _038_ en_co_clk net55 vss net72 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_181 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_217_ vss net26 _052_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput18 ctlp[1] net18 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_250_ vss _072_ _071_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout53 net53 vss vdd net56 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout75 vss net75 net76 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__216__A2 vss net36 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_302_ vdd vss _012_ _093_ _110_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_233_ vss net39 _063_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_146 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ vdd vss _052_ mask\[9\] net36 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput19 ctlp[2] net19 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_378_ vdd vss _033_ _160_ _165_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout66 vss net66 net68 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd vss _011_ _104_ _109_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vss _164_ _163_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd vss _062_ _060_ _061_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ _017_ state\[2\] net53 vss net70 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vss net2 clk vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output22_I vss net22 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_206 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__282__I vss _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout57 vss net57 net65 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout79 vss net79 net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout68 vss net68 net69 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] vss vdd gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_139 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__277__I vss _093_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_427_ _016_ state\[1\] net53 vdd vss net70 vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_17_161 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__385__A2 vss net47 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_358_ vdd vss _053_ _151_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_289_ net30 vdd vss _103_ mask\[3\] _099_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout58 net58 vss vdd net59 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout69 vss net69 net74 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_374_ vdd _061_ _056_ _162_ calibrate vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 vss net4 en vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
X_426_ _015_ state\[0\] net64 vss net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_211_ vss net24 _050_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput5 vss net5 rstn vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_78 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_210_ vdd vss _050_ mask\[7\] net34 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] vss vdd gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_206 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net49 vss vdd net50 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_17_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__303__A2 vss _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_54 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_286_ vdd vss _005_ _094_ _101_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_355_ vdd vss _149_ _026_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_14_123 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vss _032_ _159_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_285_ net28 vdd vss _101_ mask\[1\] _099_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_423_ _012_ net35 net55 vss net72 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_199_ net20 vss vdd _046_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] vss vdd gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ vss vdd gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_284_ vdd vss _004_ _094_ _100_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_422_ _011_ net34 net61 vss net78 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output36_I vss net36 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_353_ vdd vss _148_ _025_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_336_ vdd vss _138_ _018_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_198_ vdd vss _046_ mask\[3\] net30 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_266_ vdd vss _055_ _085_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_197_ vdd vss net19 net9 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vss cal_count\[3\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd vss _124_ _115_ _118_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_403_ vdd vss _183_ cal_count\[2\] _176_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vss net41 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_334_ vss _137_ _132_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_196_ net19 vss vdd _045_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ vss _070_ _069_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_38 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_317_ vss _014_ _123_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__409__A2 vss _077_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_171 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] vss vdd gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_109 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_50 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate vss vdd gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_212 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_60 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_104 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_280_ vdd vss _097_ _095_ _096_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_332_ _126_ vdd vss _017_ _127_ _135_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_401_ vdd _180_ _179_ _181_ _174_ vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_194_ vss net8 net18 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_246_ vss _068_ _055_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_290 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_213 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout76_I vss net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_193_ net18 vss vdd _044_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_400_ vdd vss _180_ cal_count\[1\] _178_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_262_ vdd vss cal_itt\[1\] _082_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_331_ _134_ vdd vss _135_ _086_ _132_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__303__B vss net36 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_245_ vdd vss net6 _067_ net67 vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_314_ vdd vss _121_ _085_ _069_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_206 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_261_ vss _081_ _059_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_192_ vdd vss _044_ mask\[1\] net28 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_330_ vdd vss _134_ _133_ _062_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ vdd vss _120_ _059_ _119_ vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__190__I vss _043_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_244_ vdd vss en_co_clk _067_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__257__A1 vss _053_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_96 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_260_ vdd _080_ _079_ _000_ _073_ vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_191_ vdd vss net17 net7 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_389_ _171_ vdd vss _172_ _115_ _120_ vss vdd gf180mcu_fd_sc_mcu7t5v0__and3_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd vss net47 net42 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_87 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_98 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_242_ net47 vss vdd _066_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_15_228 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_164 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_310_ _090_ vdd vss _117_ _060_ _113_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_88 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd vss _049_ mask\[6\] net33 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ vss vdd gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_240_ vdd vss net41 net46 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_274 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss vss vdd gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_368_ vdd vss trim_mask\[4\] _158_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_78 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_222_ vdd vss net38 net43 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_384_ vdd vss _036_ _160_ _168_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_10_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vss net38 _054_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ _008_ net31 net60 vss net77 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vss net59 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 vss vdd gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__408__A2 vss cal_count\[3\] vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_127 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_366_ vdd vss trim_mask\[3\] _157_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd vss _054_ trim_val\[0\] _053_ vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
X_418_ _007_ net30 net60 vss net77 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_349_ vdd vss _146_ _023_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output21_I vss net21 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_28 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd vss _035_ _160_ _167_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 vss vdd gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_18_209 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ vss vdd gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_279_ vdd vss _096_ _090_ state\[1\] vss vdd gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_6_231 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_91 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output14_I vss net14 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_212 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_94 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_134 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I vss rstn vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_156 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__243__I vss net47 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput40 trim[2] net40 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 vss vdd gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_5_148 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ vss vdd gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_416_ _005_ net28 net62 vss net79 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_13_290 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_347_ vdd vss _145_ _022_ vss vdd gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 vss vdd gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_201_ vdd vss _047_ mask\[4\] net31 vss vdd gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd vss vdd gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_196 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 result[3] net30 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ vss vdd gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput6 clkc net6 vdd vss vss vdd gf180mcu_fd_sc_mcu7t5v0__buf_8
.ends

.subckt saradc vinp vinn result[0] result[1] result[2] result[3] result[4] result[5]
+ result[6] result[7] result[8] result[9] valid cal en clk rstn vss
Xlatch_0 latch_0/Q latch_0/Qn latch_0/R latch_0/S latch_0/tutyuu1 latch_0/tutyuu2
+ vss vss latch
Xbuffer_0 sarlogic_0/clkc buffer_0/buf_out vss buffer
Xdacp_0 vinp dacp_0/dac_out vss dacp_0/ctl1 dacp_0/ctl2 dacp_0/ctl3 dacp_0/ctl4 dacp_0/ctl5
+ dacp_0/ctl6 dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9 dacp_0/ctl10 dacp_0/sample vss vss
+ vss dacp
Xdacn_0 vinn dacn_0/dac_out vss dacn_0/ctl1 dacn_0/ctl2 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5
+ dacn_0/ctl6 dacn_0/ctl7 dacn_0/ctl8 dacn_0/ctl9 dacn_0/ctl10 dacp_0/sample vss vss
+ vss dacn
Xcomparator_0 sarlogic_0/trim[1] sarlogic_0/trim[0] sarlogic_0/trim[2] sarlogic_0/trim[3]
+ sarlogic_0/trim[4] sarlogic_0/trimb[4] sarlogic_0/trimb[1] sarlogic_0/trimb[0] sarlogic_0/trimb[2]
+ sarlogic_0/trimb[3] dacp_0/dac_out dacn_0/dac_out latch_0/S latch_0/R comparator_0/in
+ comparator_0/ip buffer_0/buf_out comparator_0/diff vss vss comparator
Xmim_cap_boss_0 vss vss vss mim_cap_boss
Xsarlogic_0 dacn_0/ctl10 dacn_0/ctl1 dacn_0/ctl2 dacn_0/ctl3 dacn_0/ctl4 dacn_0/ctl5
+ dacn_0/ctl6 dacn_0/ctl7 dacn_0/ctl8 dacn_0/ctl9 dacp_0/ctl10 dacp_0/ctl1 dacp_0/ctl2
+ dacp_0/ctl3 dacp_0/ctl4 dacp_0/ctl5 dacp_0/ctl6 dacp_0/ctl7 dacp_0/ctl8 dacp_0/ctl9
+ cal clk sarlogic_0/clkc latch_0/Q en result[0] result[1] result[2] result[3] result[4]
+ result[5] result[6] result[7] result[8] result[9] rstn dacp_0/sample sarlogic_0/trim[0]
+ sarlogic_0/trim[1] sarlogic_0/trim[2] sarlogic_0/trim[3] sarlogic_0/trim[4] sarlogic_0/trimb[0]
+ sarlogic_0/trimb[1] sarlogic_0/trimb[2] sarlogic_0/trimb[3] sarlogic_0/trimb[4]
+ valid vss vss sarlogic
Xmim_cap_boss_1 vss vss vss mim_cap_boss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xsaradc io_in[30] io_in[32] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] io_out[10] io_out[11] io_out[12] io_out[2] io_in[3] io_in[2] io_in[1]
+ io_in[0] vss saradc
.ends

