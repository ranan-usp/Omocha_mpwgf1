magic
tech gf180mcuD
magscale 1 5
timestamp 1701229122
<< obsm1 >>
rect 672 1538 17384 11398
<< metal2 >>
rect 896 12600 952 13000
rect 2688 12600 2744 13000
rect 4480 12600 4536 13000
rect 6272 12600 6328 13000
rect 8064 12600 8120 13000
rect 9856 12600 9912 13000
rect 11648 12600 11704 13000
rect 13440 12600 13496 13000
rect 15232 12600 15288 13000
rect 17024 12600 17080 13000
rect 896 0 952 400
rect 2688 0 2744 400
rect 4480 0 4536 400
rect 6272 0 6328 400
rect 8064 0 8120 400
rect 9856 0 9912 400
rect 11648 0 11704 400
rect 13440 0 13496 400
rect 15232 0 15288 400
rect 17024 0 17080 400
<< obsm2 >>
rect 854 12570 866 12642
rect 982 12570 2658 12642
rect 2774 12570 4450 12642
rect 4566 12570 6242 12642
rect 6358 12570 8034 12642
rect 8150 12570 9826 12642
rect 9942 12570 11618 12642
rect 11734 12570 13410 12642
rect 13526 12570 15202 12642
rect 15318 12570 16994 12642
rect 17110 12570 17370 12642
rect 854 430 17370 12570
rect 854 350 866 430
rect 982 350 2658 430
rect 2774 350 4450 430
rect 4566 350 6242 430
rect 6358 350 8034 430
rect 8150 350 9826 430
rect 9942 350 11618 430
rect 11734 350 13410 430
rect 13526 350 15202 430
rect 15318 350 16994 430
rect 17110 350 17370 430
<< metal3 >>
rect 17600 12320 18000 12376
rect 0 11984 400 12040
rect 17600 11536 18000 11592
rect 0 10976 400 11032
rect 17600 10752 18000 10808
rect 0 9968 400 10024
rect 17600 9968 18000 10024
rect 17600 9184 18000 9240
rect 0 8960 400 9016
rect 17600 8400 18000 8456
rect 0 7952 400 8008
rect 17600 7616 18000 7672
rect 0 6944 400 7000
rect 17600 6832 18000 6888
rect 17600 6048 18000 6104
rect 0 5936 400 5992
rect 17600 5264 18000 5320
rect 0 4928 400 4984
rect 17600 4480 18000 4536
rect 0 3920 400 3976
rect 17600 3696 18000 3752
rect 0 2912 400 2968
rect 17600 2912 18000 2968
rect 17600 2128 18000 2184
rect 0 1904 400 1960
rect 17600 1344 18000 1400
rect 0 896 400 952
rect 17600 560 18000 616
<< obsm3 >>
rect 400 12290 17570 12362
rect 400 12070 17600 12290
rect 430 11954 17600 12070
rect 400 11622 17600 11954
rect 400 11506 17570 11622
rect 400 11062 17600 11506
rect 430 10946 17600 11062
rect 400 10838 17600 10946
rect 400 10722 17570 10838
rect 400 10054 17600 10722
rect 430 9938 17570 10054
rect 400 9270 17600 9938
rect 400 9154 17570 9270
rect 400 9046 17600 9154
rect 430 8930 17600 9046
rect 400 8486 17600 8930
rect 400 8370 17570 8486
rect 400 8038 17600 8370
rect 430 7922 17600 8038
rect 400 7702 17600 7922
rect 400 7586 17570 7702
rect 400 7030 17600 7586
rect 430 6918 17600 7030
rect 430 6914 17570 6918
rect 400 6802 17570 6914
rect 400 6134 17600 6802
rect 400 6022 17570 6134
rect 430 6018 17570 6022
rect 430 5906 17600 6018
rect 400 5350 17600 5906
rect 400 5234 17570 5350
rect 400 5014 17600 5234
rect 430 4898 17600 5014
rect 400 4566 17600 4898
rect 400 4450 17570 4566
rect 400 4006 17600 4450
rect 430 3890 17600 4006
rect 400 3782 17600 3890
rect 400 3666 17570 3782
rect 400 2998 17600 3666
rect 430 2882 17570 2998
rect 400 2214 17600 2882
rect 400 2098 17570 2214
rect 400 1990 17600 2098
rect 430 1874 17600 1990
rect 400 1430 17600 1874
rect 400 1314 17570 1430
rect 400 982 17600 1314
rect 430 866 17600 982
rect 400 646 17600 866
rect 400 574 17570 646
<< metal4 >>
rect 2671 1538 2831 11398
rect 4750 1538 4910 11398
rect 6829 1538 6989 11398
rect 8908 1538 9068 11398
rect 10987 1538 11147 11398
rect 13066 1538 13226 11398
rect 15145 1538 15305 11398
rect 17224 1538 17384 11398
<< obsm4 >>
rect 9646 4769 10066 6599
<< labels >>
rlabel metal3 s 17600 2912 18000 2968 6 cal
port 1 nsew signal input
rlabel metal3 s 17600 1344 18000 1400 6 clk
port 2 nsew signal input
rlabel metal3 s 0 5936 400 5992 6 clkc
port 3 nsew signal output
rlabel metal3 s 0 6944 400 7000 6 comp
port 4 nsew signal input
rlabel metal2 s 896 0 952 400 6 ctln[0]
port 5 nsew signal output
rlabel metal2 s 17024 0 17080 400 6 ctln[1]
port 6 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 ctln[2]
port 7 nsew signal output
rlabel metal2 s 13440 0 13496 400 6 ctln[3]
port 8 nsew signal output
rlabel metal2 s 11648 0 11704 400 6 ctln[4]
port 9 nsew signal output
rlabel metal2 s 9856 0 9912 400 6 ctln[5]
port 10 nsew signal output
rlabel metal2 s 8064 0 8120 400 6 ctln[6]
port 11 nsew signal output
rlabel metal2 s 6272 0 6328 400 6 ctln[7]
port 12 nsew signal output
rlabel metal2 s 4480 0 4536 400 6 ctln[8]
port 13 nsew signal output
rlabel metal2 s 2688 0 2744 400 6 ctln[9]
port 14 nsew signal output
rlabel metal2 s 896 12600 952 13000 6 ctlp[0]
port 15 nsew signal output
rlabel metal2 s 17024 12600 17080 13000 6 ctlp[1]
port 16 nsew signal output
rlabel metal2 s 15232 12600 15288 13000 6 ctlp[2]
port 17 nsew signal output
rlabel metal2 s 13440 12600 13496 13000 6 ctlp[3]
port 18 nsew signal output
rlabel metal2 s 11648 12600 11704 13000 6 ctlp[4]
port 19 nsew signal output
rlabel metal2 s 9856 12600 9912 13000 6 ctlp[5]
port 20 nsew signal output
rlabel metal2 s 8064 12600 8120 13000 6 ctlp[6]
port 21 nsew signal output
rlabel metal2 s 6272 12600 6328 13000 6 ctlp[7]
port 22 nsew signal output
rlabel metal2 s 4480 12600 4536 13000 6 ctlp[8]
port 23 nsew signal output
rlabel metal2 s 2688 12600 2744 13000 6 ctlp[9]
port 24 nsew signal output
rlabel metal3 s 17600 2128 18000 2184 6 en
port 25 nsew signal input
rlabel metal3 s 17600 5264 18000 5320 6 result[0]
port 26 nsew signal output
rlabel metal3 s 17600 6048 18000 6104 6 result[1]
port 27 nsew signal output
rlabel metal3 s 17600 6832 18000 6888 6 result[2]
port 28 nsew signal output
rlabel metal3 s 17600 7616 18000 7672 6 result[3]
port 29 nsew signal output
rlabel metal3 s 17600 8400 18000 8456 6 result[4]
port 30 nsew signal output
rlabel metal3 s 17600 9184 18000 9240 6 result[5]
port 31 nsew signal output
rlabel metal3 s 17600 9968 18000 10024 6 result[6]
port 32 nsew signal output
rlabel metal3 s 17600 10752 18000 10808 6 result[7]
port 33 nsew signal output
rlabel metal3 s 17600 11536 18000 11592 6 result[8]
port 34 nsew signal output
rlabel metal3 s 17600 12320 18000 12376 6 result[9]
port 35 nsew signal output
rlabel metal3 s 17600 560 18000 616 6 rstn
port 36 nsew signal input
rlabel metal3 s 17600 4480 18000 4536 6 sample
port 37 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 trim[0]
port 38 nsew signal output
rlabel metal3 s 0 3920 400 3976 6 trim[1]
port 39 nsew signal output
rlabel metal3 s 0 1904 400 1960 6 trim[2]
port 40 nsew signal output
rlabel metal3 s 0 896 400 952 6 trim[3]
port 41 nsew signal output
rlabel metal3 s 0 4928 400 4984 6 trim[4]
port 42 nsew signal output
rlabel metal3 s 0 9968 400 10024 6 trimb[0]
port 43 nsew signal output
rlabel metal3 s 0 8960 400 9016 6 trimb[1]
port 44 nsew signal output
rlabel metal3 s 0 10976 400 11032 6 trimb[2]
port 45 nsew signal output
rlabel metal3 s 0 11984 400 12040 6 trimb[3]
port 46 nsew signal output
rlabel metal3 s 0 7952 400 8008 6 trimb[4]
port 47 nsew signal output
rlabel metal3 s 17600 3696 18000 3752 6 valid
port 48 nsew signal output
rlabel metal4 s 2671 1538 2831 11398 6 vdd
port 49 nsew power bidirectional
rlabel metal4 s 6829 1538 6989 11398 6 vdd
port 49 nsew power bidirectional
rlabel metal4 s 10987 1538 11147 11398 6 vdd
port 49 nsew power bidirectional
rlabel metal4 s 15145 1538 15305 11398 6 vdd
port 49 nsew power bidirectional
rlabel metal4 s 4750 1538 4910 11398 6 vss
port 50 nsew ground bidirectional
rlabel metal4 s 8908 1538 9068 11398 6 vss
port 50 nsew ground bidirectional
rlabel metal4 s 13066 1538 13226 11398 6 vss
port 50 nsew ground bidirectional
rlabel metal4 s 17224 1538 17384 11398 6 vss
port 50 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 13000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 764234
string GDS_FILE /home/oe23ranan/gf_analog/openlane/sarlogic/runs/23_11_29_12_37/results/signoff/sarlogic.magic.gds
string GDS_START 214126
<< end >>

