* NGSPICE file created from comparator.ext - technology: gf180mcuD

.subckt XM3$2 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n640_n791# a_n336_n791# 0.040052f
C1 a_n176_n791# a_n80_n571# 0.005902f
C2 a_n176_n791# a_n336_n791# 0.131547f
C3 a_n80_n571# a_n16_n791# 0.005902f
C4 a_n496_n791# a_n400_n571# 0.005902f
C5 a_n176_n791# a_n16_n791# 0.131547f
C6 a_n336_n791# a_n16_n791# 0.040052f
C7 a_n496_n791# a_n640_n791# 0.131547f
C8 a_n400_n571# a_n240_n571# 0.043712f
C9 a_n496_n791# a_n560_n571# 0.005902f
C10 a_n80_n571# a_n240_n571# 0.043712f
C11 a_n496_n791# a_n336_n791# 0.131547f
C12 a_n176_n791# a_n240_n571# 0.005902f
C13 a_n400_n571# a_n560_n571# 0.043712f
C14 a_n336_n791# a_n240_n571# 0.005902f
C15 a_n336_n791# a_n400_n571# 0.005902f
C16 a_n640_n791# a_n560_n571# 0.005902f
C17 a_n16_n791# a_n778_n975# 0.182857f
C18 a_n176_n791# a_n778_n975# 0.043869f
C19 a_n336_n791# a_n778_n975# 0.097543f
C20 a_n496_n791# a_n778_n975# 0.043869f
C21 a_n640_n791# a_n778_n975# 0.277121f
C22 a_n80_n571# a_n778_n975# 0.191307f
C23 a_n240_n571# a_n778_n975# 0.164084f
C24 a_n400_n571# a_n778_n975# 0.16416f
C25 a_n560_n571# a_n778_n975# 0.198604f
.ends

.subckt XM2$2 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n157_n712# a_n237_n932# 0.005902f
C1 a_3_n712# a_67_n932# 0.005902f
C2 a_n93_n932# a_n237_n932# 0.131547f
C3 a_n93_n932# a_67_n932# 0.131547f
C4 a_n237_n932# a_67_n932# 0.040052f
C5 a_3_n712# a_n157_n712# 0.043712f
C6 a_n93_n932# a_3_n712# 0.005902f
C7 a_n93_n932# a_n157_n712# 0.005902f
C8 a_67_n932# a_n375_n1116# 0.182823f
C9 a_n93_n932# a_n375_n1116# 0.043869f
C10 a_n237_n932# a_n375_n1116# 0.182332f
C11 a_3_n712# a_n375_n1116# 0.191252f
C12 a_n157_n712# a_n375_n1116# 0.191252f
.ends

.subckt XM0$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n266_803# a_n202_583# 0.005902f
C1 a_n346_583# a_n266_803# 0.011845f
C2 a_n346_583# a_n202_583# 0.14243f
C3 a_n202_583# a_n484_399# 0.098801f
C4 a_n346_583# a_n484_399# 0.215099f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM1$2 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n266_803# a_n202_583# 0.011845f
C1 a_n346_583# a_n266_803# 0.001764f
C2 a_n346_583# a_n202_583# 0.075352f
C3 a_n202_583# a_n484_399# 0.24117f
C4 a_n346_583# a_n484_399# 0.057381f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM4$2 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_2250_n696# a_2090_n696# 0.043712f
C1 a_1610_n696# a_1514_n916# 0.005902f
C2 a_1930_n696# a_1834_n916# 0.005902f
C3 a_1674_n916# a_1994_n916# 0.040052f
C4 a_2154_n916# a_1994_n916# 0.131547f
C5 a_1834_n916# a_1770_n696# 0.005902f
C6 a_2250_n696# a_2410_n696# 0.043712f
C7 a_2154_n916# a_2090_n696# 0.005902f
C8 a_1674_n916# a_1514_n916# 0.131547f
C9 a_1930_n696# a_1770_n696# 0.043712f
C10 a_1514_n916# a_1354_n916# 0.131547f
C11 a_2474_n916# a_2410_n696# 0.005902f
C12 a_1994_n916# a_2314_n916# 0.040052f
C13 a_1450_n696# a_1514_n916# 0.005902f
C14 a_2250_n696# a_2154_n916# 0.005902f
C15 a_1210_n916# a_1354_n916# 0.131547f
C16 a_1610_n696# a_1674_n916# 0.005902f
C17 a_1834_n916# a_1994_n916# 0.131547f
C18 a_1930_n696# a_1994_n916# 0.005902f
C19 a_1930_n696# a_2090_n696# 0.043712f
C20 a_2410_n696# a_2314_n916# 0.005902f
C21 a_2250_n696# a_2314_n916# 0.005902f
C22 a_1610_n696# a_1450_n696# 0.043712f
C23 a_1674_n916# a_1354_n916# 0.040052f
C24 a_1290_n696# a_1210_n916# 0.005902f
C25 a_2474_n916# a_2314_n916# 0.131547f
C26 a_1450_n696# a_1354_n916# 0.005902f
C27 a_2154_n916# a_2314_n916# 0.131547f
C28 a_1290_n696# a_1354_n916# 0.005902f
C29 a_1610_n696# a_1770_n696# 0.043712f
C30 a_1834_n916# a_1674_n916# 0.131547f
C31 a_1994_n916# a_2090_n696# 0.005902f
C32 a_1450_n696# a_1290_n696# 0.043712f
C33 a_1770_n696# a_1674_n916# 0.005902f
C34 a_2474_n916# a_1072_n1100# 0.19427f
C35 a_2314_n916# a_1072_n1100# 0.126868f
C36 a_2154_n916# a_1072_n1100# 0.043869f
C37 a_1994_n916# a_1072_n1100# 0.097543f
C38 a_1834_n916# a_1072_n1100# 0.043869f
C39 a_1674_n916# a_1072_n1100# 0.097543f
C40 a_1514_n916# a_1072_n1100# 0.043869f
C41 a_1354_n916# a_1072_n1100# 0.126868f
C42 a_1210_n916# a_1072_n1100# 0.099481f
C43 a_2410_n696# a_1072_n1100# 0.198604f
C44 a_2250_n696# a_1072_n1100# 0.16416f
C45 a_2090_n696# a_1072_n1100# 0.164084f
C46 a_1930_n696# a_1072_n1100# 0.164049f
C47 a_1770_n696# a_1072_n1100# 0.164031f
C48 a_1610_n696# a_1072_n1100# 0.16402f
C49 a_1450_n696# a_1072_n1100# 0.164014f
C50 a_1290_n696# a_1072_n1100# 0.191268f
.ends

.subckt trim_switch$1 m1_n149_n1117# m1_n1378_n1819# m1_711_n1117# m1_n2738_n1819#
+ m1_n447_n1117# m1_n2669_n1117# XM1$2_0/a_n202_583# XM0$1_0/a_n346_583# m1_n1309_n1117#
+ m1_802_n1819# VSUBS
XXM3$2_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$2
XXM2$2_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$2
XXM0$1_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0$1_0/a_n346_583# XM0$1
XXM1$2_0 VSUBS XM1$2_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$2
XXM4$2_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$2
C0 m1_n1309_n1117# m1_n1378_n1819# 0.014034f
C1 m1_n447_n1117# m1_n1309_n1117# 0.041018f
C2 XM1$2_0/a_n202_583# XM0$1_0/a_n346_583# 0.027386f
C3 m1_n447_n1117# m1_n149_n1117# 0.123582f
C4 m1_n2738_n1819# m1_n1378_n1819# 0.040124f
C5 m1_n1309_n1117# m1_n2669_n1117# 0.027949f
C6 m1_n149_n1117# m1_711_n1117# 0.02663f
C7 m1_802_n1819# m1_711_n1117# 0.272119f
C8 XM0$1_0/a_n346_583# m1_n1378_n1819# 0.039382f
C9 m1_n2669_n1117# m1_n2738_n1819# 0.092062f
C10 m1_n447_n1117# XM0$1_0/a_n346_583# 0.07096f
C11 m1_n149_n1117# XM1$2_0/a_n202_583# 0.07096f
C12 m1_802_n1819# XM1$2_0/a_n202_583# 0.00859f
C13 m1_802_n1819# VSUBS 1.278621f
C14 m1_711_n1117# VSUBS 1.959711f
C15 XM1$2_0/a_n202_583# VSUBS 0.42776f
C16 m1_n149_n1117# VSUBS 0.407201f
C17 XM0$1_0/a_n346_583# VSUBS 0.314559f
C18 m1_n447_n1117# VSUBS 0.388025f
C19 m1_n1378_n1819# VSUBS 0.604021f
C20 m1_n1309_n1117# VSUBS 0.637566f
C21 m1_n2738_n1819# VSUBS 1.12292f
C22 m1_n2669_n1117# VSUBS 1.128649f
.ends

.subckt trim$1 n4 n1 n0 n2 n3 drain d_4 d_1 d_0 d_2 d_3 VSUBS
Xtrim_switch$1_0 d_1 n2 d_4 n3 d_0 d_3 n1 n0 d_2 n4 VSUBS trim_switch$1
C0 n0 n4 0.166348f
C1 d_4 n2 0.00312f
C2 n1 d_1 0.003099f
C3 d_1 n2 0.003137f
C4 n1 n2 0.081094f
C5 drain n1 1.60623f
C6 n3 n1 0.087807f
C7 drain n2 3.213024f
C8 n3 n2 0.58337f
C9 n0 n1 0.520979f
C10 n3 drain 6.427485f
C11 n0 n2 0.103368f
C12 n0 drain 1.60623f
C13 d_0 n2 0.002632f
C14 n3 n0 0.087807f
C15 n0 d_0 0.004139f
C16 n4 n1 0.169398f
C17 n4 n2 0.596682f
C18 n4 drain 12.877382f
C19 n3 n4 1.600479f
C20 n2 VSUBS 2.03715f
C21 n4 VSUBS 4.367046f
C22 drain VSUBS -5.906306f
C23 n3 VSUBS 3.463842f
C24 n0 VSUBS 0.689164f
C25 n1 VSUBS 0.727243f
C26 d_4 VSUBS 1.64786f
C27 d_1 VSUBS 0.345562f
C28 d_0 VSUBS 0.33412f
C29 d_2 VSUBS 0.513348f
C30 d_3 VSUBS 0.927186f
.ends

.subckt XM3 a_n71_n882# a_73_n882# a_9_n662# w_n509_n1092# VSUBS
X0 a_73_n882# a_9_n662# a_n71_n882# w_n509_n1092# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n71_n882# a_73_n882# 0.06854f
C1 w_n509_n1092# a_73_n882# 0.008358f
C2 w_n509_n1092# a_n71_n882# 0.010275f
C3 a_9_n662# a_73_n882# 0.001764f
C4 a_9_n662# a_n71_n882# 0.001764f
C5 w_n509_n1092# a_9_n662# 0.131025f
C6 a_73_n882# VSUBS 0.049403f
C7 a_n71_n882# VSUBS 0.047486f
C8 a_9_n662# VSUBS 0.087507f
C9 w_n509_n1092# VSUBS 1.54752f
.ends

.subckt XMinn a_719_n1284# a_937_n880# a_857_n1100# a_719_n788# a_1001_n1100#
X0 a_1001_n1100# a_937_n880# a_857_n1100# a_719_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_857_n1100# a_1001_n1100# 0.06854f
C1 a_937_n880# a_1001_n1100# 0.001764f
C2 a_937_n880# a_857_n1100# 0.001764f
C3 a_1001_n1100# a_719_n1284# 0.057707f
C4 a_857_n1100# a_719_n1284# 0.057707f
C5 a_937_n880# a_719_n1284# 0.21851f
.ends

.subckt XM1 a_n1416_1000# a_n1336_908# a_n1272_1000# w_n1578_790# VSUBS
X0 a_n1272_1000# a_n1336_908# a_n1416_1000# w_n1578_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n1416_1000# a_n1272_1000# 0.06854f
C1 w_n1578_790# a_n1272_1000# 0.021497f
C2 w_n1578_790# a_n1416_1000# 0.022441f
C3 a_n1336_908# a_n1272_1000# 0.001764f
C4 a_n1336_908# a_n1416_1000# 0.001764f
C5 w_n1578_790# a_n1336_908# 0.132558f
C6 a_n1272_1000# VSUBS 0.043675f
C7 a_n1416_1000# VSUBS 0.043675f
C8 a_n1336_908# VSUBS 0.08816f
C9 w_n1578_790# VSUBS 1.17557f
.ends

.subckt XM2$1 a_3_n712# a_n375_n620# a_n157_n712# a_n375_n1116# a_n237_n932# a_67_n932#
+ a_n93_n932#
X0 a_67_n932# a_3_n712# a_n93_n932# a_n375_n1116# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n93_n932# a_n157_n712# a_n237_n932# a_n375_n1116# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n93_n932# a_3_n712# 0.005902f
C1 a_n157_n712# a_n93_n932# 0.005902f
C2 a_n157_n712# a_n237_n932# 0.005902f
C3 a_n157_n712# a_3_n712# 0.043712f
C4 a_n93_n932# a_67_n932# 0.131547f
C5 a_n237_n932# a_67_n932# 0.040052f
C6 a_3_n712# a_67_n932# 0.005902f
C7 a_n93_n932# a_n237_n932# 0.131547f
C8 a_67_n932# a_n375_n1116# 0.182823f
C9 a_n93_n932# a_n375_n1116# 0.043869f
C10 a_n237_n932# a_n375_n1116# 0.182332f
C11 a_3_n712# a_n375_n1116# 0.191252f
C12 a_n157_n712# a_n375_n1116# 0.191252f
.ends

.subckt XM1$1 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n346_583# a_n202_583# 0.075352f
C1 a_n266_803# a_n202_583# 0.011845f
C2 a_n266_803# a_n346_583# 0.001764f
C3 a_n202_583# a_n484_399# 0.24117f
C4 a_n346_583# a_n484_399# 0.057381f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt XM4$1 a_1930_n696# a_2474_n916# a_1514_n916# a_2250_n696# a_1290_n696# a_1210_n916#
+ a_1674_n916# a_1450_n696# a_2410_n696# a_1072_n1100# a_1834_n916# a_1610_n696# a_2154_n916#
+ a_1994_n916# a_1770_n696# a_2314_n916# a_1354_n916# a_2090_n696#
X0 a_1834_n916# a_1770_n696# a_1674_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_2154_n916# a_2090_n696# a_1994_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_1674_n916# a_1610_n696# a_1514_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_1514_n916# a_1450_n696# a_1354_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_2474_n916# a_2410_n696# a_2314_n916# a_1072_n1100# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_1354_n916# a_1290_n696# a_1210_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_1994_n916# a_1930_n696# a_1834_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_2314_n916# a_2250_n696# a_2154_n916# a_1072_n1100# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_1450_n696# a_1514_n916# 0.005902f
C1 a_1834_n916# a_1674_n916# 0.131547f
C2 a_2250_n696# a_2410_n696# 0.043712f
C3 a_1610_n696# a_1770_n696# 0.043712f
C4 a_1834_n916# a_1994_n916# 0.131547f
C5 a_1994_n916# a_2314_n916# 0.040052f
C6 a_1514_n916# a_1674_n916# 0.131547f
C7 a_2314_n916# a_2154_n916# 0.131547f
C8 a_1994_n916# a_1674_n916# 0.040052f
C9 a_1994_n916# a_2154_n916# 0.131547f
C10 a_1994_n916# a_2090_n696# 0.005902f
C11 a_2474_n916# a_2410_n696# 0.005902f
C12 a_2154_n916# a_2090_n696# 0.005902f
C13 a_1834_n916# a_1930_n696# 0.005902f
C14 a_1290_n696# a_1354_n916# 0.005902f
C15 a_1834_n916# a_1770_n696# 0.005902f
C16 a_1450_n696# a_1610_n696# 0.043712f
C17 a_2410_n696# a_2314_n916# 0.005902f
C18 a_1770_n696# a_1674_n916# 0.005902f
C19 a_1290_n696# a_1450_n696# 0.043712f
C20 a_2250_n696# a_2314_n916# 0.005902f
C21 a_1994_n916# a_1930_n696# 0.005902f
C22 a_1450_n696# a_1354_n916# 0.005902f
C23 a_1610_n696# a_1674_n916# 0.005902f
C24 a_1930_n696# a_2090_n696# 0.043712f
C25 a_2250_n696# a_2154_n916# 0.005902f
C26 a_1610_n696# a_1514_n916# 0.005902f
C27 a_2250_n696# a_2090_n696# 0.043712f
C28 a_1290_n696# a_1210_n916# 0.005902f
C29 a_1354_n916# a_1674_n916# 0.040052f
C30 a_1930_n696# a_1770_n696# 0.043712f
C31 a_1210_n916# a_1354_n916# 0.131547f
C32 a_1354_n916# a_1514_n916# 0.131547f
C33 a_2474_n916# a_2314_n916# 0.131547f
C34 a_2474_n916# a_1072_n1100# 0.19427f
C35 a_2314_n916# a_1072_n1100# 0.126868f
C36 a_2154_n916# a_1072_n1100# 0.043869f
C37 a_1994_n916# a_1072_n1100# 0.097543f
C38 a_1834_n916# a_1072_n1100# 0.043869f
C39 a_1674_n916# a_1072_n1100# 0.097543f
C40 a_1514_n916# a_1072_n1100# 0.043869f
C41 a_1354_n916# a_1072_n1100# 0.126868f
C42 a_1210_n916# a_1072_n1100# 0.099481f
C43 a_2410_n696# a_1072_n1100# 0.198604f
C44 a_2250_n696# a_1072_n1100# 0.16416f
C45 a_2090_n696# a_1072_n1100# 0.164084f
C46 a_1930_n696# a_1072_n1100# 0.164049f
C47 a_1770_n696# a_1072_n1100# 0.164031f
C48 a_1610_n696# a_1072_n1100# 0.16402f
C49 a_1450_n696# a_1072_n1100# 0.164014f
C50 a_1290_n696# a_1072_n1100# 0.191268f
.ends

.subckt XM3$1 a_n16_n791# a_n778_n975# a_n80_n571# a_n176_n791# a_n240_n571# a_n336_n791#
+ a_n400_n571# a_n496_n791# a_n560_n571# a_n640_n791#
X0 a_n336_n791# a_n400_n571# a_n496_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n176_n791# a_n240_n571# a_n336_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n16_n791# a_n80_n571# a_n176_n791# a_n778_n975# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n496_n791# a_n560_n571# a_n640_n791# a_n778_n975# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n560_n571# a_n400_n571# 0.043712f
C1 a_n496_n791# a_n336_n791# 0.131547f
C2 a_n560_n571# a_n640_n791# 0.005902f
C3 a_n80_n571# a_n176_n791# 0.005902f
C4 a_n240_n571# a_n400_n571# 0.043712f
C5 a_n240_n571# a_n176_n791# 0.005902f
C6 a_n400_n571# a_n336_n791# 0.005902f
C7 a_n16_n791# a_n176_n791# 0.131547f
C8 a_n176_n791# a_n336_n791# 0.131547f
C9 a_n80_n571# a_n240_n571# 0.043712f
C10 a_n640_n791# a_n336_n791# 0.040052f
C11 a_n560_n571# a_n496_n791# 0.005902f
C12 a_n16_n791# a_n80_n571# 0.005902f
C13 a_n240_n571# a_n336_n791# 0.005902f
C14 a_n16_n791# a_n336_n791# 0.040052f
C15 a_n496_n791# a_n400_n571# 0.005902f
C16 a_n496_n791# a_n640_n791# 0.131547f
C17 a_n16_n791# a_n778_n975# 0.182857f
C18 a_n176_n791# a_n778_n975# 0.043869f
C19 a_n336_n791# a_n778_n975# 0.097543f
C20 a_n496_n791# a_n778_n975# 0.043869f
C21 a_n640_n791# a_n778_n975# 0.277121f
C22 a_n80_n571# a_n778_n975# 0.191307f
C23 a_n240_n571# a_n778_n975# 0.164084f
C24 a_n400_n571# a_n778_n975# 0.16416f
C25 a_n560_n571# a_n778_n975# 0.198604f
.ends

.subckt XM0 a_n484_399# a_n202_583# a_n266_803# a_n484_895# a_n346_583#
X0 a_n202_583# a_n266_803# a_n346_583# a_n484_399# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n202_583# a_n266_803# 0.005902f
C1 a_n346_583# a_n266_803# 0.011845f
C2 a_n346_583# a_n202_583# 0.14243f
C3 a_n202_583# a_n484_399# 0.098801f
C4 a_n346_583# a_n484_399# 0.215099f
C5 a_n266_803# a_n484_399# 0.21851f
.ends

.subckt trim_switch m1_n149_n1117# XM0_0/a_n346_583# m1_711_n1117# XM1$1_0/a_n202_583#
+ m1_n447_n1117# m1_n2669_n1117# m1_802_n1819# m1_n1309_n1117# m1_n1378_n1819# m1_n2738_n1819#
+ VSUBS
XXM2$1_0 m1_n1309_n1117# VSUBS m1_n1309_n1117# VSUBS m1_n1378_n1819# m1_n1378_n1819#
+ VSUBS XM2$1
XXM1$1_0 VSUBS XM1$1_0/a_n202_583# m1_n149_n1117# VSUBS VSUBS XM1$1
XXM4$1_0 m1_711_n1117# VSUBS VSUBS m1_711_n1117# m1_711_n1117# VSUBS m1_802_n1819#
+ m1_711_n1117# m1_711_n1117# VSUBS VSUBS m1_711_n1117# VSUBS m1_802_n1819# m1_711_n1117#
+ m1_802_n1819# m1_802_n1819# m1_711_n1117# XM4$1
XXM3$1_0 m1_n2738_n1819# VSUBS m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819#
+ m1_n2669_n1117# VSUBS m1_n2669_n1117# m1_n2738_n1819# XM3$1
XXM0_0 VSUBS VSUBS m1_n447_n1117# VSUBS XM0_0/a_n346_583# XM0
C0 XM0_0/a_n346_583# XM1$1_0/a_n202_583# 0.027386f
C1 m1_n149_n1117# XM1$1_0/a_n202_583# 0.07096f
C2 m1_n2669_n1117# m1_n2738_n1819# 0.092062f
C3 m1_711_n1117# m1_802_n1819# 0.272119f
C4 m1_n1378_n1819# m1_n1309_n1117# 0.014034f
C5 m1_711_n1117# m1_n149_n1117# 0.02663f
C6 m1_n447_n1117# m1_n1309_n1117# 0.041018f
C7 XM0_0/a_n346_583# m1_n1378_n1819# 0.039382f
C8 XM0_0/a_n346_583# m1_n447_n1117# 0.07096f
C9 m1_n2669_n1117# m1_n1309_n1117# 0.027949f
C10 m1_n447_n1117# m1_n149_n1117# 0.123582f
C11 XM1$1_0/a_n202_583# m1_802_n1819# 0.00859f
C12 m1_n1378_n1819# m1_n2738_n1819# 0.040124f
C13 XM0_0/a_n346_583# VSUBS 0.314559f
C14 m1_n447_n1117# VSUBS 0.388025f
C15 m1_n2738_n1819# VSUBS 1.12292f
C16 m1_n2669_n1117# VSUBS 1.128649f
C17 m1_802_n1819# VSUBS 1.278621f
C18 m1_711_n1117# VSUBS 1.959711f
C19 XM1$1_0/a_n202_583# VSUBS 0.42776f
C20 m1_n149_n1117# VSUBS 0.407201f
C21 m1_n1378_n1819# VSUBS 0.604021f
C22 m1_n1309_n1117# VSUBS 0.637566f
.ends

.subckt trim n1 n0 n3 d_4 d_1 d_0 d_2 d_3 n4 drain n2 VSUBS
Xtrim_switch_0 d_1 n0 d_4 n1 d_0 d_3 n4 d_2 n2 n3 VSUBS trim_switch
C0 d_0 n0 0.004139f
C1 d_1 n2 0.003137f
C2 d_0 n2 0.002632f
C3 n4 n1 0.169398f
C4 n4 drain 12.877382f
C5 drain n1 1.60623f
C6 n4 n3 1.600479f
C7 n3 n1 0.087807f
C8 drain n3 6.427485f
C9 d_4 n2 0.00312f
C10 n4 n0 0.166348f
C11 n4 n2 0.596682f
C12 n0 n1 0.520979f
C13 n2 n1 0.081094f
C14 drain n0 1.60623f
C15 drain n2 3.213024f
C16 n3 n0 0.087807f
C17 n2 n3 0.58337f
C18 d_1 n1 0.003099f
C19 n2 n0 0.103368f
C20 n0 VSUBS 0.689164f
C21 n1 VSUBS 0.727243f
C22 n4 VSUBS 4.367046f
C23 drain VSUBS -5.906306f
C24 n2 VSUBS 2.03715f
C25 n3 VSUBS 3.463842f
C26 d_0 VSUBS 0.33412f
C27 d_3 VSUBS 0.927186f
C28 d_4 VSUBS 1.64786f
C29 d_1 VSUBS 0.345562f
C30 d_2 VSUBS 0.513348f
.ends

.subckt XMl4 a_44_908# a_108_1000# a_n36_1000# w_n198_790# VSUBS
X0 a_108_1000# a_44_908# a_n36_1000# w_n198_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_44_908# w_n198_790# 0.131025f
C1 a_n36_1000# a_44_908# 0.001764f
C2 a_n36_1000# w_n198_790# 0.008358f
C3 a_108_1000# a_44_908# 0.001764f
C4 a_108_1000# w_n198_790# 0.010275f
C5 a_n36_1000# a_108_1000# 0.06854f
C6 a_108_1000# VSUBS 0.047486f
C7 a_n36_1000# VSUBS 0.049403f
C8 a_44_908# VSUBS 0.087507f
C9 w_n198_790# VSUBS 1.54752f
.ends

.subckt XMl2 a_33_n1100# a_n111_n1100# a_n31_n880# a_n249_n1284#
X0 a_33_n1100# a_n31_n880# a_n111_n1100# a_n249_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n111_n1100# a_n31_n880# 0.001764f
C1 a_33_n1100# a_n111_n1100# 0.06854f
C2 a_33_n1100# a_n31_n880# 0.001764f
C3 a_33_n1100# a_n249_n1284# 0.066395f
C4 a_n111_n1100# a_n249_n1284# 0.057707f
C5 a_n31_n880# a_n249_n1284# 0.218606f
.ends

.subckt XM4 a_1264_908# a_1328_1000# w_1022_790# a_1184_1000# VSUBS
X0 a_1328_1000# a_1264_908# a_1184_1000# w_1022_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_1264_908# w_1022_790# 0.132558f
C1 a_1184_1000# a_1264_908# 0.001764f
C2 a_1184_1000# w_1022_790# 0.021497f
C3 a_1328_1000# a_1264_908# 0.001764f
C4 a_1328_1000# w_1022_790# 0.022441f
C5 a_1184_1000# a_1328_1000# 0.06854f
C6 a_1328_1000# VSUBS 0.043675f
C7 a_1184_1000# VSUBS 0.043675f
C8 a_1264_908# VSUBS 0.08816f
C9 w_1022_790# VSUBS 1.17557f
.ends

.subckt XM2 a_69_n911# w_n237_n1121# a_5_n691# a_n75_n911# VSUBS
X0 a_69_n911# a_5_n691# a_n75_n911# w_n237_n1121# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_5_n691# w_n237_n1121# 0.131025f
C1 a_n75_n911# a_5_n691# 0.001764f
C2 a_n75_n911# w_n237_n1121# 0.008358f
C3 a_69_n911# a_5_n691# 0.001764f
C4 a_69_n911# w_n237_n1121# 0.010275f
C5 a_n75_n911# a_69_n911# 0.06854f
C6 a_69_n911# VSUBS 0.047486f
C7 a_n75_n911# VSUBS 0.049403f
C8 a_5_n691# VSUBS 0.087507f
C9 w_n237_n1121# VSUBS 1.54752f
.ends

.subckt XMdiff a_721_n1097# a_817_n1189# a_439_n1281# a_657_n1189# a_577_n1097# a_881_n1097#
X0 a_721_n1097# a_657_n1189# a_577_n1097# a_439_n1281# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_881_n1097# a_817_n1189# a_721_n1097# a_439_n1281# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
C0 a_721_n1097# a_881_n1097# 0.06854f
C1 a_817_n1189# a_657_n1189# 0.043712f
C2 a_577_n1097# a_657_n1189# 0.001764f
C3 a_721_n1097# a_817_n1189# 0.001764f
C4 a_721_n1097# a_657_n1189# 0.001764f
C5 a_577_n1097# a_721_n1097# 0.06854f
C6 a_817_n1189# a_881_n1097# 0.001764f
C7 a_881_n1097# a_439_n1281# 0.115307f
C8 a_721_n1097# a_439_n1281# 0.02923f
C9 a_577_n1097# a_439_n1281# 0.115307f
C10 a_817_n1189# a_439_n1281# 0.191347f
C11 a_657_n1189# a_439_n1281# 0.191347f
.ends

.subckt XMl3 a_n116_908# w_n634_790# a_n196_1000# a_n52_1000# VSUBS
X0 a_n52_1000# a_n116_908# a_n196_1000# w_n634_790# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_n116_908# w_n634_790# 0.139286f
C1 a_n196_1000# a_n116_908# 0.001764f
C2 a_n196_1000# w_n634_790# 0.024248f
C3 a_n52_1000# a_n116_908# 0.001764f
C4 a_n52_1000# w_n634_790# 0.021497f
C5 a_n196_1000# a_n52_1000# 0.06854f
C6 a_n52_1000# VSUBS 0.043675f
C7 a_n196_1000# VSUBS 0.041759f
C8 a_n116_908# VSUBS 0.081314f
C9 w_n634_790# VSUBS 1.68331f
.ends

.subckt XMl1 a_1362_n1100# a_1442_n880# a_1506_n1100# a_1224_n1284#
X0 a_1506_n1100# a_1442_n880# a_1362_n1100# a_1224_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_1362_n1100# a_1442_n880# 0.001764f
C1 a_1506_n1100# a_1362_n1100# 0.06854f
C2 a_1506_n1100# a_1442_n880# 0.001764f
C3 a_1506_n1100# a_1224_n1284# 0.057707f
C4 a_1362_n1100# a_1224_n1284# 0.066395f
C5 a_1442_n880# a_1224_n1284# 0.218606f
.ends

.subckt XMinp a_251_n1284# a_389_n1100# a_251_n788# a_469_n880# a_533_n1100#
X0 a_533_n1100# a_469_n880# a_389_n1100# a_251_n1284# nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 a_389_n1100# a_469_n880# 0.001764f
C1 a_533_n1100# a_469_n880# 0.001764f
C2 a_389_n1100# a_533_n1100# 0.06854f
C3 a_533_n1100# a_251_n1284# 0.057707f
C4 a_389_n1100# a_251_n1284# 0.057707f
C5 a_469_n880# a_251_n1284# 0.21851f
.ends

.subckt comparator diff ip in clkc vss vdd outp outn vp vn trim4 trim1 trim0 trim2
+ trim3 trimb4 trimb1 trimb0 trimb2 trimb3
Xtrim$1_0 trim$1_0/n4 trim$1_0/n1 trim$1_0/n0 trim$1_0/n2 trim$1_0/n3 in trim4 trim1
+ trim0 trim2 trim3 vss trim$1
XXM3_0 outp vdd clkc vdd vss XM3
XXMinn_0 vss vn in vss diff XMinn
XXM1_0 in clkc vdd vdd vss XM1
Xtrim_0 trim_0/n1 trim_0/n0 trim_0/n3 trimb4 trimb1 trimb0 trimb2 trimb3 trim_0/n4
+ ip trim_0/n2 vss trim
XXMl4_0 outn outp vdd vdd vss XMl4
XXMl2_0 outp ip outn vss XMl2
XXM4_0 clkc ip vdd vdd vss XM4
XXM2_0 outn vdd clkc vdd vss XM2
XXMdiff_0 diff clkc vss clkc vss vss XMdiff
XXMl3_0 outp vdd outn vdd vss XMl3
XXMl1_0 outn outp in vss XMl1
XXMinp_0 vss diff vss vp ip XMinp
C0 vn vdd 0.059928f
C1 trim4 trim0 0.001193f
C2 trim0 trim2 0.78245f
C3 trim$1_0/n2 trim$1_0/n4 0.128631f
C4 trim_0/n2 trim_0/n4 0.128631f
C5 trim$1_0/n4 trim$1_0/n0 0.032158f
C6 trimb2 trimb3 0.919951f
C7 outp vdd 0.441033f
C8 in outn 0.120156f
C9 trim$1_0/n1 trim$1_0/n0 0.032158f
C10 trim_0/n1 trim_0/n0 0.032158f
C11 clkc in 0.467511f
C12 ip trim_0/n1 1.606993f
C13 clkc outn 0.223756f
C14 ip outn 0.016739f
C15 vp outn 0.197573f
C16 trimb4 trimb0 0.001193f
C17 ip trim_0/n0 1.606993f
C18 ip clkc 0.46748f
C19 clkc vp 0.104841f
C20 ip vp 0.542294f
C21 diff in 0.133902f
C22 trim$1_0/n1 trim$1_0/n4 0.032158f
C23 trimb0 trimb1 0.720503f
C24 trim_0/n1 trim_0/n4 0.032158f
C25 trim1 trim4 0.420884f
C26 diff outn 0.003297f
C27 trim$1_0/n2 in 3.21681f
C28 diff clkc 0.071648f
C29 ip diff 0.133902f
C30 diff vp 0.004194f
C31 trim_0/n0 trim_0/n4 0.032158f
C32 in vn 0.542295f
C33 trim$1_0/n0 in 1.606993f
C34 ip trim_0/n4 12.853658f
C35 trim$1_0/n4 trim$1_0/n3 0.241184f
C36 outn vn 0.196568f
C37 trim3 trim2 0.919951f
C38 outp in 0.016739f
C39 in vdd 0.088929f
C40 clkc vn 0.104842f
C41 ip trim_0/n3 6.427209f
C42 vp vn 0.180638f
C43 trimb4 trim_0/n4 0.002224f
C44 trimb2 trimb0 0.78245f
C45 outp outn 1.248977f
C46 trim$1_0/n4 in 12.853658f
C47 outn vdd 0.464524f
C48 trimb4 trimb1 0.420884f
C49 outp clkc 0.22388f
C50 trim$1_0/n1 in 1.606993f
C51 outp ip 0.120151f
C52 clkc vdd 0.233505f
C53 outp vp 0.243335f
C54 trim_0/n4 trimb1 0.001374f
C55 ip vdd 0.088929f
C56 vp vdd 0.059928f
C57 trim1 trim$1_0/n4 0.001374f
C58 diff vn 0.004194f
C59 trim_0/n3 trim_0/n4 0.241184f
C60 trim1 trim0 0.720503f
C61 outp diff 0.006112f
C62 in trim$1_0/n3 6.427209f
C63 ip trim_0/n2 3.21681f
C64 trim$1_0/n4 trim4 0.002224f
C65 outp vn 0.223138f
C66 vp vss 1.116181f
C67 outn vss 2.443821f
C68 clkc vss 4.180552f
C69 vdd vss 7.878819f
C70 outp vss 2.478554f
C71 trim_0/n0 vss 0.677622f
C72 trim_0/n1 vss 0.716105f
C73 trim_0/n4 vss 4.199544f
C74 ip vss -4.381578f
C75 trim_0/n2 vss 1.980196f
C76 trim_0/n3 vss 3.31053f
C77 trimb0 vss 0.985146f
C78 trimb3 vss 2.983196f
C79 trimb4 vss 2.263372f
C80 trimb1 vss 0.99849f
C81 trimb2 vss 1.41065f
C82 diff vss 0.21339f
C83 vn vss 1.131981f
C84 trim$1_0/n2 vss 1.980196f
C85 trim$1_0/n4 vss 4.199544f
C86 in vss -4.381556f
C87 trim$1_0/n3 vss 3.31053f
C88 trim$1_0/n0 vss 0.677622f
C89 trim$1_0/n1 vss 0.716105f
C90 trim4 vss 2.263372f
C91 trim1 vss 0.99849f
C92 trim0 vss 0.985146f
C93 trim2 vss 1.41065f
C94 trim3 vss 2.983196f
.ends

