VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO saradc
  CLASS BLOCK ;
  FOREIGN saradc ;
  ORIGIN 838.480 1163.700 ;
  SIZE 1679.800 BY 2327.400 ;
  PIN vss
    ANTENNADIFFAREA 703.663269 ;
    PORT
      LAYER Pwell ;
        RECT -494.560 94.725 -491.460 97.505 ;
        RECT -495.535 80.535 -491.455 87.615 ;
        RECT 145.205 59.240 147.395 102.660 ;
        RECT 295.490 43.000 462.670 46.520 ;
        RECT 364.880 42.865 367.795 43.000 ;
        RECT 403.520 42.865 406.435 43.000 ;
        RECT 431.245 42.865 434.160 43.000 ;
        RECT 327.920 38.680 330.835 38.815 ;
        RECT 448.605 38.680 451.520 38.815 ;
        RECT 295.490 35.160 462.670 38.680 ;
        RECT 351.440 35.025 354.355 35.160 ;
        RECT 399.600 35.025 402.515 35.160 ;
        RECT 440.205 35.025 443.120 35.160 ;
        RECT 165.715 31.815 190.995 34.895 ;
        RECT 326.240 30.840 329.155 30.975 ;
        RECT 372.720 30.840 375.635 30.975 ;
        RECT 440.765 30.840 443.680 30.975 ;
        RECT 295.490 27.320 462.670 30.840 ;
        RECT 348.640 27.185 351.555 27.320 ;
        RECT 448.605 23.000 451.520 23.135 ;
        RECT 295.490 19.480 462.670 23.000 ;
        RECT 302.035 19.355 308.065 19.480 ;
        RECT 398.480 19.345 401.395 19.480 ;
        RECT 372.720 15.160 375.635 15.295 ;
        RECT 413.600 15.160 416.515 15.295 ;
        RECT 448.605 15.160 451.520 15.295 ;
        RECT 295.490 11.640 462.670 15.160 ;
        RECT 180.815 -2.590 183.895 2.590 ;
        RECT 184.815 -1.790 187.895 1.790 ;
        RECT 229.175 -2.120 232.275 11.560 ;
        RECT 321.830 11.515 322.930 11.640 ;
        RECT 345.715 11.515 351.745 11.640 ;
        RECT 377.760 7.320 380.675 7.455 ;
        RECT 418.080 7.320 420.995 7.455 ;
        RECT 295.490 3.800 462.670 7.320 ;
        RECT 364.880 3.665 367.795 3.800 ;
        RECT 337.440 -0.520 340.355 -0.385 ;
        RECT 448.605 -0.520 451.520 -0.385 ;
        RECT 295.490 -4.040 462.670 -0.520 ;
        RECT 306.175 -4.165 312.205 -4.040 ;
        RECT 330.160 -8.360 333.075 -8.225 ;
        RECT 451.680 -8.360 454.595 -8.225 ;
        RECT 229.550 -12.550 232.330 -9.450 ;
        RECT 233.065 -12.550 235.845 -9.450 ;
        RECT 295.490 -11.880 462.670 -8.360 ;
        RECT 432.365 -12.015 435.280 -11.880 ;
        RECT 341.360 -16.200 344.275 -16.065 ;
        RECT 295.490 -19.720 462.670 -16.200 ;
        RECT 312.800 -19.855 315.715 -19.720 ;
        RECT 443.280 -19.855 446.195 -19.720 ;
        RECT 409.120 -24.040 412.035 -23.905 ;
        RECT 295.490 -27.560 462.670 -24.040 ;
        RECT 307.760 -27.695 310.675 -27.560 ;
        RECT 165.715 -34.895 190.995 -31.815 ;
        RECT 337.440 -31.880 340.355 -31.745 ;
        RECT 451.680 -31.880 454.595 -31.745 ;
        RECT 295.490 -35.400 462.670 -31.880 ;
        RECT 310.000 -35.535 312.915 -35.400 ;
        RECT 438.810 -35.525 442.590 -35.400 ;
        RECT 338.560 -39.720 341.475 -39.585 ;
        RECT 378.880 -39.720 381.795 -39.585 ;
        RECT 409.120 -39.720 412.035 -39.585 ;
        RECT 295.490 -43.240 462.670 -39.720 ;
        RECT 325.680 -43.375 328.595 -43.240 ;
        RECT 361.245 -43.375 364.160 -43.240 ;
        RECT 388.685 -43.375 391.600 -43.240 ;
        RECT 429.840 -43.375 432.755 -43.240 ;
        RECT 295.490 -49.750 462.670 -47.560 ;
        RECT -495.535 -87.615 -491.455 -80.535 ;
        RECT -494.560 -97.505 -491.460 -94.725 ;
        RECT 145.205 -102.660 147.395 -59.240 ;
      LAYER Metal1 ;
        RECT 146.625 127.660 147.865 132.620 ;
        RECT 146.665 101.860 147.825 127.660 ;
        RECT 145.775 101.520 147.825 101.860 ;
        RECT 146.665 98.815 147.825 101.520 ;
        RECT 146.015 98.585 147.825 98.815 ;
        RECT -494.375 96.630 -494.145 97.115 ;
        RECT -494.375 96.565 -492.575 96.630 ;
        RECT -494.525 96.400 -492.575 96.565 ;
        RECT 146.665 96.545 147.825 98.585 ;
        RECT -494.525 95.665 -494.145 96.400 ;
        RECT 146.015 96.315 147.825 96.545 ;
        RECT -494.375 95.115 -494.145 95.665 ;
        RECT 146.665 95.455 147.825 96.315 ;
        RECT 146.015 95.225 147.825 95.455 ;
        RECT 146.665 93.185 147.825 95.225 ;
        RECT 146.015 92.955 147.825 93.185 ;
        RECT 146.665 92.095 147.825 92.955 ;
        RECT 146.015 91.865 147.825 92.095 ;
        RECT 146.665 89.825 147.825 91.865 ;
        RECT 146.015 89.595 147.825 89.825 ;
        RECT 146.665 88.735 147.825 89.595 ;
        RECT 146.015 88.505 147.825 88.735 ;
        RECT -496.745 84.700 -496.365 85.370 ;
        RECT -495.350 84.700 -495.120 87.115 ;
        RECT 146.665 86.465 147.825 88.505 ;
        RECT 146.015 86.235 147.825 86.465 ;
        RECT 146.665 85.375 147.825 86.235 ;
        RECT 146.015 85.145 147.825 85.375 ;
        RECT -496.745 84.470 -492.560 84.700 ;
        RECT 146.665 83.105 147.825 85.145 ;
        RECT 146.015 82.875 147.825 83.105 ;
        RECT 146.665 82.015 147.825 82.875 ;
        RECT 146.015 81.785 147.825 82.015 ;
        RECT 146.665 79.745 147.825 81.785 ;
        RECT 146.015 79.515 147.825 79.745 ;
        RECT 146.665 78.655 147.825 79.515 ;
        RECT 146.015 78.425 147.825 78.655 ;
        RECT 146.665 76.385 147.825 78.425 ;
        RECT 146.015 76.155 147.825 76.385 ;
        RECT 146.665 75.295 147.825 76.155 ;
        RECT 146.015 75.065 147.825 75.295 ;
        RECT 146.665 73.025 147.825 75.065 ;
        RECT 146.015 72.795 147.825 73.025 ;
        RECT 146.665 71.935 147.825 72.795 ;
        RECT 146.015 71.705 147.825 71.935 ;
        RECT 146.665 69.665 147.825 71.705 ;
        RECT 146.015 69.435 147.825 69.665 ;
        RECT 146.665 68.575 147.825 69.435 ;
        RECT 146.015 68.345 147.825 68.575 ;
        RECT 146.665 66.305 147.825 68.345 ;
        RECT 146.015 66.075 147.825 66.305 ;
        RECT 146.665 65.215 147.825 66.075 ;
        RECT 146.015 64.985 147.825 65.215 ;
        RECT 146.665 62.945 147.825 64.985 ;
        RECT 146.015 62.715 147.825 62.945 ;
        RECT 146.665 60.380 147.825 62.715 ;
        RECT 145.775 60.040 147.825 60.380 ;
        RECT 146.665 59.670 147.825 60.040 ;
        RECT 296.290 45.060 296.630 45.950 ;
        RECT 299.310 45.060 299.650 45.525 ;
        RECT 301.550 45.060 301.890 45.525 ;
        RECT 303.790 45.060 304.130 45.525 ;
        RECT 306.030 45.060 306.370 45.525 ;
        RECT 308.270 45.060 308.610 45.525 ;
        RECT 310.510 45.060 310.850 45.525 ;
        RECT 312.750 45.060 313.090 45.525 ;
        RECT 315.350 45.060 315.690 45.945 ;
        RECT 316.830 45.060 317.170 45.525 ;
        RECT 319.070 45.060 319.410 45.525 ;
        RECT 321.310 45.060 321.650 45.525 ;
        RECT 323.550 45.060 323.890 45.525 ;
        RECT 325.790 45.060 326.130 45.525 ;
        RECT 328.030 45.060 328.370 45.525 ;
        RECT 330.270 45.060 330.610 45.525 ;
        RECT 331.445 45.060 331.675 45.855 ;
        RECT 334.390 45.060 334.730 45.945 ;
        RECT 335.710 45.060 336.050 45.525 ;
        RECT 337.950 45.060 338.290 45.525 ;
        RECT 340.190 45.060 340.530 45.525 ;
        RECT 342.430 45.060 342.770 45.525 ;
        RECT 344.670 45.060 345.010 45.525 ;
        RECT 346.910 45.060 347.250 45.525 ;
        RECT 349.150 45.060 349.490 45.525 ;
        RECT 349.925 45.060 350.155 45.855 ;
        RECT 353.430 45.060 353.770 45.945 ;
        RECT 354.350 45.060 354.690 45.525 ;
        RECT 356.590 45.060 356.930 45.525 ;
        RECT 358.830 45.060 359.170 45.525 ;
        RECT 361.070 45.060 361.410 45.525 ;
        RECT 363.310 45.060 363.650 45.525 ;
        RECT 365.550 45.060 365.890 45.525 ;
        RECT 367.790 45.060 368.130 45.525 ;
        RECT 368.965 45.060 369.195 45.855 ;
        RECT 372.470 45.060 372.810 45.945 ;
        RECT 373.790 45.060 374.130 45.525 ;
        RECT 376.030 45.060 376.370 45.525 ;
        RECT 378.270 45.060 378.610 45.525 ;
        RECT 380.510 45.060 380.850 45.525 ;
        RECT 382.750 45.060 383.090 45.525 ;
        RECT 384.990 45.060 385.330 45.525 ;
        RECT 387.230 45.060 387.570 45.525 ;
        RECT 391.510 45.060 391.850 45.945 ;
        RECT 392.830 45.060 393.170 45.525 ;
        RECT 395.070 45.060 395.410 45.525 ;
        RECT 397.310 45.060 397.650 45.525 ;
        RECT 399.550 45.060 399.890 45.525 ;
        RECT 401.790 45.060 402.130 45.525 ;
        RECT 404.030 45.060 404.370 45.525 ;
        RECT 406.270 45.060 406.610 45.525 ;
        RECT 410.550 45.060 410.890 45.945 ;
        RECT 411.470 45.060 411.810 45.525 ;
        RECT 413.710 45.060 414.050 45.525 ;
        RECT 415.950 45.060 416.290 45.525 ;
        RECT 418.190 45.060 418.530 45.525 ;
        RECT 420.430 45.060 420.770 45.525 ;
        RECT 422.670 45.060 423.010 45.525 ;
        RECT 424.910 45.060 425.250 45.525 ;
        RECT 426.085 45.060 426.315 45.705 ;
        RECT 428.325 45.060 428.555 45.850 ;
        RECT 429.590 45.060 429.930 45.945 ;
        RECT 430.910 45.060 431.250 45.525 ;
        RECT 433.150 45.060 433.490 45.525 ;
        RECT 435.390 45.060 435.730 45.525 ;
        RECT 437.630 45.060 437.970 45.525 ;
        RECT 439.870 45.060 440.210 45.525 ;
        RECT 442.110 45.060 442.450 45.525 ;
        RECT 444.350 45.060 444.690 45.525 ;
        RECT 448.630 45.060 448.970 45.945 ;
        RECT 449.605 45.060 449.835 45.830 ;
        RECT 451.845 45.060 452.075 45.830 ;
        RECT 454.085 45.060 454.315 45.830 ;
        RECT 456.325 45.060 456.555 45.830 ;
        RECT 458.565 45.060 458.795 45.855 ;
        RECT 461.530 45.060 461.870 45.950 ;
        RECT 295.920 44.460 463.040 45.060 ;
        RECT 296.290 43.570 296.630 44.460 ;
        RECT 297.630 43.995 297.970 44.460 ;
        RECT 299.870 43.995 300.210 44.460 ;
        RECT 302.110 43.995 302.450 44.460 ;
        RECT 304.350 43.995 304.690 44.460 ;
        RECT 306.590 43.995 306.930 44.460 ;
        RECT 308.830 43.995 309.170 44.460 ;
        RECT 311.070 43.995 311.410 44.460 ;
        RECT 313.365 43.720 313.595 44.460 ;
        RECT 315.605 43.720 315.835 44.460 ;
        RECT 320.805 43.690 321.035 44.460 ;
        RECT 323.045 43.690 323.275 44.460 ;
        RECT 325.285 43.690 325.515 44.460 ;
        RECT 327.525 43.690 327.755 44.460 ;
        RECT 329.765 43.665 329.995 44.460 ;
        RECT 334.645 43.600 334.875 44.460 ;
        RECT 335.510 43.575 335.850 44.460 ;
        RECT 337.660 43.935 337.890 44.460 ;
        RECT 340.140 43.910 340.370 44.460 ;
        RECT 343.425 43.895 343.655 44.460 ;
        RECT 345.445 43.665 345.675 44.460 ;
        RECT 349.365 43.600 349.595 44.460 ;
        RECT 352.905 43.895 353.135 44.460 ;
        RECT 356.590 43.710 356.935 44.460 ;
        RECT 358.450 43.685 358.790 44.460 ;
        RECT 363.710 43.845 364.050 44.460 ;
        RECT 369.350 43.630 369.580 44.460 ;
        RECT 372.595 43.885 372.935 44.460 ;
        RECT 374.710 43.575 375.050 44.460 ;
        RECT 376.910 43.910 377.140 44.460 ;
        RECT 379.390 43.935 379.620 44.460 ;
        RECT 380.890 43.710 381.230 44.460 ;
        RECT 383.130 43.665 383.470 44.460 ;
        RECT 385.270 44.035 385.500 44.460 ;
        RECT 389.350 43.855 389.580 44.460 ;
        RECT 391.365 43.720 391.595 44.460 ;
        RECT 395.230 43.710 395.575 44.460 ;
        RECT 397.090 43.685 397.430 44.460 ;
        RECT 402.350 43.845 402.690 44.460 ;
        RECT 407.990 43.630 408.220 44.460 ;
        RECT 411.235 43.885 411.575 44.460 ;
        RECT 413.910 43.575 414.250 44.460 ;
        RECT 415.265 43.995 415.495 44.460 ;
        RECT 418.645 43.995 418.875 44.460 ;
        RECT 419.745 43.995 419.975 44.460 ;
        RECT 423.125 43.995 423.355 44.460 ;
        RECT 426.105 43.885 426.445 44.460 ;
        RECT 429.460 43.630 429.690 44.460 ;
        RECT 434.990 43.845 435.330 44.460 ;
        RECT 440.250 43.685 440.590 44.460 ;
        RECT 442.105 43.710 442.450 44.460 ;
        RECT 444.005 43.815 444.235 44.460 ;
        RECT 446.245 43.670 446.475 44.460 ;
        RECT 449.605 43.665 449.835 44.460 ;
        RECT 453.110 43.575 453.450 44.460 ;
        RECT 454.085 43.675 454.315 44.460 ;
        RECT 456.325 43.675 456.555 44.460 ;
        RECT 458.565 43.665 458.795 44.460 ;
        RECT 461.530 43.570 461.870 44.460 ;
        RECT 296.290 37.220 296.630 38.110 ;
        RECT 297.630 37.220 297.970 37.685 ;
        RECT 299.870 37.220 300.210 37.685 ;
        RECT 302.110 37.220 302.450 37.685 ;
        RECT 304.350 37.220 304.690 37.685 ;
        RECT 306.590 37.220 306.930 37.685 ;
        RECT 308.830 37.220 309.170 37.685 ;
        RECT 311.070 37.220 311.410 37.685 ;
        RECT 315.910 37.220 316.250 38.105 ;
        RECT 319.630 37.220 319.975 37.970 ;
        RECT 321.490 37.220 321.830 37.995 ;
        RECT 326.750 37.220 327.090 37.835 ;
        RECT 332.390 37.220 332.620 38.050 ;
        RECT 335.635 37.220 335.975 37.795 ;
        RECT 337.985 37.220 338.215 37.685 ;
        RECT 341.365 37.220 341.595 37.685 ;
        RECT 344.325 37.220 344.555 37.990 ;
        RECT 346.565 37.220 346.795 37.990 ;
        RECT 348.805 37.220 349.035 37.990 ;
        RECT 351.045 37.220 351.275 37.990 ;
        RECT 355.110 37.220 355.450 38.105 ;
        RECT 356.085 37.220 356.315 38.005 ;
        RECT 358.325 37.220 358.555 38.005 ;
        RECT 362.085 37.220 362.315 37.960 ;
        RECT 362.870 37.220 363.100 37.645 ;
        RECT 366.950 37.220 367.180 37.825 ;
        RECT 367.845 37.220 368.075 37.965 ;
        RECT 370.085 37.220 370.315 37.965 ;
        RECT 372.325 37.220 372.555 37.965 ;
        RECT 374.565 37.220 374.795 37.965 ;
        RECT 376.805 37.220 377.035 37.965 ;
        RECT 379.045 37.220 379.275 37.965 ;
        RECT 381.285 37.220 381.515 37.965 ;
        RECT 383.525 37.220 383.755 37.965 ;
        RECT 386.990 37.220 387.220 37.770 ;
        RECT 389.470 37.220 389.700 37.745 ;
        RECT 390.245 37.220 390.475 37.960 ;
        RECT 394.310 37.220 394.650 38.105 ;
        RECT 395.285 37.220 395.515 37.990 ;
        RECT 397.525 37.220 397.755 37.990 ;
        RECT 399.765 37.220 399.995 37.990 ;
        RECT 402.005 37.220 402.235 37.990 ;
        RECT 404.190 37.220 404.530 37.685 ;
        RECT 406.430 37.220 406.770 37.685 ;
        RECT 408.670 37.220 409.010 37.685 ;
        RECT 410.910 37.220 411.250 37.685 ;
        RECT 413.150 37.220 413.490 37.685 ;
        RECT 415.390 37.220 415.730 37.685 ;
        RECT 417.630 37.220 417.970 37.685 ;
        RECT 419.150 37.220 419.490 37.685 ;
        RECT 421.390 37.220 421.730 37.685 ;
        RECT 423.630 37.220 423.970 37.685 ;
        RECT 425.870 37.220 426.210 37.685 ;
        RECT 428.110 37.220 428.450 37.685 ;
        RECT 430.350 37.220 430.690 37.685 ;
        RECT 432.590 37.220 432.930 37.685 ;
        RECT 433.510 37.220 433.850 38.105 ;
        RECT 434.865 37.220 435.095 37.685 ;
        RECT 438.245 37.220 438.475 37.685 ;
        RECT 438.965 37.220 439.195 37.865 ;
        RECT 441.205 37.220 441.435 38.010 ;
        RECT 443.465 37.220 443.805 37.795 ;
        RECT 446.820 37.220 447.050 38.050 ;
        RECT 452.350 37.220 452.690 37.835 ;
        RECT 457.610 37.220 457.950 37.995 ;
        RECT 459.465 37.220 459.810 37.970 ;
        RECT 461.530 37.220 461.870 38.110 ;
        RECT 295.920 36.620 463.040 37.220 ;
        RECT 296.290 35.730 296.630 36.620 ;
        RECT 297.630 36.155 297.970 36.620 ;
        RECT 299.870 36.155 300.210 36.620 ;
        RECT 302.110 36.155 302.450 36.620 ;
        RECT 304.350 36.155 304.690 36.620 ;
        RECT 306.590 36.155 306.930 36.620 ;
        RECT 308.830 36.155 309.170 36.620 ;
        RECT 311.070 36.155 311.410 36.620 ;
        RECT 311.845 35.875 312.075 36.620 ;
        RECT 314.085 35.875 314.315 36.620 ;
        RECT 316.325 35.875 316.555 36.620 ;
        RECT 318.565 35.875 318.795 36.620 ;
        RECT 320.805 35.875 321.035 36.620 ;
        RECT 323.045 35.875 323.275 36.620 ;
        RECT 325.285 35.875 325.515 36.620 ;
        RECT 327.525 35.875 327.755 36.620 ;
        RECT 329.765 35.835 329.995 36.620 ;
        RECT 332.005 35.835 332.235 36.620 ;
        RECT 335.510 35.735 335.850 36.620 ;
        RECT 336.885 35.830 337.115 36.620 ;
        RECT 339.125 35.975 339.355 36.620 ;
        RECT 343.150 35.870 343.495 36.620 ;
        RECT 345.010 35.845 345.350 36.620 ;
        RECT 350.270 36.005 350.610 36.620 ;
        RECT 355.910 35.790 356.140 36.620 ;
        RECT 359.155 36.045 359.495 36.620 ;
        RECT 361.190 36.195 361.420 36.620 ;
        RECT 365.270 36.015 365.500 36.620 ;
        RECT 366.165 35.835 366.395 36.620 ;
        RECT 368.405 35.835 368.635 36.620 ;
        RECT 370.645 35.825 370.875 36.620 ;
        RECT 374.710 35.735 375.050 36.620 ;
        RECT 375.685 35.835 375.915 36.620 ;
        RECT 377.925 35.835 378.155 36.620 ;
        RECT 380.165 35.825 380.395 36.620 ;
        RECT 384.260 36.015 384.490 36.620 ;
        RECT 388.340 36.195 388.570 36.620 ;
        RECT 391.310 35.870 391.655 36.620 ;
        RECT 393.170 35.845 393.510 36.620 ;
        RECT 398.430 36.005 398.770 36.620 ;
        RECT 404.070 35.790 404.300 36.620 ;
        RECT 407.315 36.045 407.655 36.620 ;
        RECT 411.525 35.825 411.755 36.620 ;
        RECT 413.910 35.735 414.250 36.620 ;
        RECT 416.110 36.070 416.340 36.620 ;
        RECT 418.590 36.095 418.820 36.620 ;
        RECT 419.310 36.155 419.650 36.620 ;
        RECT 421.550 36.155 421.890 36.620 ;
        RECT 423.790 36.155 424.130 36.620 ;
        RECT 426.030 36.155 426.370 36.620 ;
        RECT 428.270 36.155 428.610 36.620 ;
        RECT 430.510 36.155 430.850 36.620 ;
        RECT 432.750 36.155 433.090 36.620 ;
        RECT 435.065 36.045 435.405 36.620 ;
        RECT 438.420 35.790 438.650 36.620 ;
        RECT 443.950 36.005 444.290 36.620 ;
        RECT 449.210 35.845 449.550 36.620 ;
        RECT 451.065 35.870 451.410 36.620 ;
        RECT 453.110 35.735 453.450 36.620 ;
        RECT 456.325 35.835 456.555 36.620 ;
        RECT 458.565 35.835 458.795 36.620 ;
        RECT 461.530 35.730 461.870 36.620 ;
        RECT 165.900 33.805 166.130 34.355 ;
        RECT 190.580 33.805 190.810 34.355 ;
        RECT 165.825 32.905 166.205 33.805 ;
        RECT 165.900 32.355 166.130 32.905 ;
        RECT 167.390 32.555 167.620 33.790 ;
        RECT 168.990 32.555 169.220 33.790 ;
        RECT 174.190 32.555 174.420 33.790 ;
        RECT 179.190 32.555 179.420 33.790 ;
        RECT 183.490 32.555 183.720 33.790 ;
        RECT 185.090 32.555 185.320 33.790 ;
        RECT 186.690 32.555 186.920 33.790 ;
        RECT 188.290 32.555 188.520 33.790 ;
        RECT 189.890 32.555 190.120 33.790 ;
        RECT 190.505 32.905 190.885 33.805 ;
        RECT 167.315 31.655 167.695 32.555 ;
        RECT 168.915 31.655 169.295 32.555 ;
        RECT 174.115 31.655 174.495 32.555 ;
        RECT 179.115 31.655 179.495 32.555 ;
        RECT 183.415 31.655 183.795 32.555 ;
        RECT 185.015 31.655 185.395 32.555 ;
        RECT 186.615 31.655 186.995 32.555 ;
        RECT 188.215 31.655 188.595 32.555 ;
        RECT 189.815 31.655 190.195 32.555 ;
        RECT 190.580 32.355 190.810 32.905 ;
        RECT 296.290 29.380 296.630 30.270 ;
        RECT 297.285 29.380 297.515 30.165 ;
        RECT 299.525 29.380 299.755 30.165 ;
        RECT 303.845 29.380 304.075 30.120 ;
        RECT 304.565 29.380 304.795 30.150 ;
        RECT 306.805 29.380 307.035 30.150 ;
        RECT 309.045 29.380 309.275 30.150 ;
        RECT 311.285 29.380 311.515 30.150 ;
        RECT 313.525 29.380 313.755 30.175 ;
        RECT 315.910 29.380 316.250 30.265 ;
        RECT 317.950 29.380 318.295 30.130 ;
        RECT 319.810 29.380 320.150 30.155 ;
        RECT 325.070 29.380 325.410 29.995 ;
        RECT 330.710 29.380 330.940 30.210 ;
        RECT 333.955 29.380 334.295 29.955 ;
        RECT 336.305 29.380 336.535 29.845 ;
        RECT 339.685 29.380 339.915 29.845 ;
        RECT 344.885 29.380 345.115 30.175 ;
        RECT 350.325 29.380 350.555 30.120 ;
        RECT 351.045 29.380 351.275 30.175 ;
        RECT 355.110 29.380 355.450 30.265 ;
        RECT 356.085 29.380 356.315 30.175 ;
        RECT 361.470 29.380 361.810 30.005 ;
        RECT 364.430 29.380 364.775 30.130 ;
        RECT 366.290 29.380 366.630 30.155 ;
        RECT 371.550 29.380 371.890 29.995 ;
        RECT 377.190 29.380 377.420 30.210 ;
        RECT 380.435 29.380 380.775 29.955 ;
        RECT 382.580 29.380 382.810 29.985 ;
        RECT 386.660 29.380 386.890 29.805 ;
        RECT 388.745 29.380 388.975 29.945 ;
        RECT 390.805 29.380 391.035 30.175 ;
        RECT 394.310 29.380 394.650 30.265 ;
        RECT 395.285 29.380 395.515 30.150 ;
        RECT 397.525 29.380 397.755 30.150 ;
        RECT 399.765 29.380 399.995 30.150 ;
        RECT 402.005 29.380 402.235 30.150 ;
        RECT 404.245 29.380 404.475 30.165 ;
        RECT 406.485 29.380 406.715 30.165 ;
        RECT 410.570 29.380 410.910 30.130 ;
        RECT 412.810 29.380 413.150 30.175 ;
        RECT 416.785 29.380 417.015 29.945 ;
        RECT 419.150 29.380 419.490 29.845 ;
        RECT 421.390 29.380 421.730 29.845 ;
        RECT 423.630 29.380 423.970 29.845 ;
        RECT 425.870 29.380 426.210 29.845 ;
        RECT 428.110 29.380 428.450 29.845 ;
        RECT 430.350 29.380 430.690 29.845 ;
        RECT 432.590 29.380 432.930 29.845 ;
        RECT 433.510 29.380 433.850 30.265 ;
        RECT 435.625 29.380 435.965 29.955 ;
        RECT 438.980 29.380 439.210 30.210 ;
        RECT 444.510 29.380 444.850 29.995 ;
        RECT 449.770 29.380 450.110 30.155 ;
        RECT 451.625 29.380 451.970 30.130 ;
        RECT 454.990 29.380 455.330 30.005 ;
        RECT 459.470 29.380 459.810 30.005 ;
        RECT 461.530 29.380 461.870 30.270 ;
        RECT 295.920 28.780 463.040 29.380 ;
        RECT 296.290 27.890 296.630 28.780 ;
        RECT 297.230 28.315 297.570 28.780 ;
        RECT 299.470 28.315 299.810 28.780 ;
        RECT 301.710 28.315 302.050 28.780 ;
        RECT 303.950 28.315 304.290 28.780 ;
        RECT 306.190 28.315 306.530 28.780 ;
        RECT 308.430 28.315 308.770 28.780 ;
        RECT 310.670 28.315 311.010 28.780 ;
        RECT 311.845 27.995 312.075 28.780 ;
        RECT 314.085 27.995 314.315 28.780 ;
        RECT 318.225 28.215 318.455 28.780 ;
        RECT 321.765 27.920 321.995 28.780 ;
        RECT 322.485 27.995 322.715 28.780 ;
        RECT 324.725 27.995 324.955 28.780 ;
        RECT 326.965 27.985 327.195 28.780 ;
        RECT 332.110 28.230 332.340 28.780 ;
        RECT 334.590 28.255 334.820 28.780 ;
        RECT 335.510 27.895 335.850 28.780 ;
        RECT 340.350 28.030 340.695 28.780 ;
        RECT 342.210 28.005 342.550 28.780 ;
        RECT 347.470 28.165 347.810 28.780 ;
        RECT 353.110 27.950 353.340 28.780 ;
        RECT 356.355 28.205 356.695 28.780 ;
        RECT 358.325 27.995 358.555 28.780 ;
        RECT 360.565 27.995 360.795 28.780 ;
        RECT 364.145 28.215 364.375 28.780 ;
        RECT 366.165 27.985 366.395 28.780 ;
        RECT 370.485 28.040 370.715 28.780 ;
        RECT 371.205 27.985 371.435 28.780 ;
        RECT 374.710 27.895 375.050 28.780 ;
        RECT 375.685 27.985 375.915 28.780 ;
        RECT 378.650 28.030 378.990 28.780 ;
        RECT 380.890 27.985 381.230 28.780 ;
        RECT 382.965 27.995 383.195 28.780 ;
        RECT 385.205 27.995 385.435 28.780 ;
        RECT 389.865 28.215 390.095 28.780 ;
        RECT 391.925 28.010 392.155 28.780 ;
        RECT 394.165 28.010 394.395 28.780 ;
        RECT 396.405 28.010 396.635 28.780 ;
        RECT 398.645 28.010 398.875 28.780 ;
        RECT 400.885 27.995 401.115 28.780 ;
        RECT 403.125 27.995 403.355 28.780 ;
        RECT 405.365 27.985 405.595 28.780 ;
        RECT 408.330 28.030 408.670 28.780 ;
        RECT 410.570 27.985 410.910 28.780 ;
        RECT 413.910 27.895 414.250 28.780 ;
        RECT 416.110 28.230 416.340 28.780 ;
        RECT 418.590 28.255 418.820 28.780 ;
        RECT 419.745 28.315 419.975 28.780 ;
        RECT 423.125 28.315 423.355 28.780 ;
        RECT 423.790 28.315 424.130 28.780 ;
        RECT 426.030 28.315 426.370 28.780 ;
        RECT 428.270 28.315 428.610 28.780 ;
        RECT 430.510 28.315 430.850 28.780 ;
        RECT 432.750 28.315 433.090 28.780 ;
        RECT 434.990 28.315 435.330 28.780 ;
        RECT 437.230 28.315 437.570 28.780 ;
        RECT 438.350 28.315 438.690 28.780 ;
        RECT 440.590 28.315 440.930 28.780 ;
        RECT 442.830 28.315 443.170 28.780 ;
        RECT 445.070 28.315 445.410 28.780 ;
        RECT 447.310 28.315 447.650 28.780 ;
        RECT 449.550 28.315 449.890 28.780 ;
        RECT 451.790 28.315 452.130 28.780 ;
        RECT 453.110 27.895 453.450 28.780 ;
        RECT 454.085 28.135 454.315 28.780 ;
        RECT 456.325 27.990 456.555 28.780 ;
        RECT 458.910 28.155 459.250 28.780 ;
        RECT 461.530 27.890 461.870 28.780 ;
        RECT 296.290 21.540 296.630 22.430 ;
        RECT 297.285 21.540 297.515 22.285 ;
        RECT 299.525 21.540 299.755 22.285 ;
        RECT 301.765 21.540 301.995 22.285 ;
        RECT 304.005 21.540 304.235 22.285 ;
        RECT 306.245 21.540 306.475 22.285 ;
        RECT 308.485 21.540 308.715 22.285 ;
        RECT 310.725 21.540 310.955 22.285 ;
        RECT 312.965 21.540 313.195 22.285 ;
        RECT 315.910 21.540 316.250 22.425 ;
        RECT 316.885 21.540 317.115 22.310 ;
        RECT 319.125 21.540 319.355 22.310 ;
        RECT 321.365 21.540 321.595 22.310 ;
        RECT 323.605 21.540 323.835 22.310 ;
        RECT 325.845 21.540 326.075 22.325 ;
        RECT 328.085 21.540 328.315 22.325 ;
        RECT 330.325 21.540 330.555 22.335 ;
        RECT 333.525 21.540 333.755 22.330 ;
        RECT 335.765 21.540 335.995 22.185 ;
        RECT 338.725 21.540 338.955 22.325 ;
        RECT 340.965 21.540 341.195 22.325 ;
        RECT 344.725 21.540 344.955 22.280 ;
        RECT 345.825 21.540 346.055 22.005 ;
        RECT 349.205 21.540 349.435 22.005 ;
        RECT 352.165 21.540 352.395 22.335 ;
        RECT 355.110 21.540 355.450 22.425 ;
        RECT 356.085 21.540 356.315 22.285 ;
        RECT 358.325 21.540 358.555 22.285 ;
        RECT 360.565 21.540 360.795 22.285 ;
        RECT 362.805 21.540 363.035 22.285 ;
        RECT 365.045 21.540 365.275 22.285 ;
        RECT 367.285 21.540 367.515 22.285 ;
        RECT 369.525 21.540 369.755 22.285 ;
        RECT 371.765 21.540 371.995 22.285 ;
        RECT 374.005 21.540 374.235 22.310 ;
        RECT 376.245 21.540 376.475 22.310 ;
        RECT 378.485 21.540 378.715 22.310 ;
        RECT 380.725 21.540 380.955 22.310 ;
        RECT 384.710 21.540 384.940 21.965 ;
        RECT 388.790 21.540 389.020 22.145 ;
        RECT 389.685 21.540 389.915 22.280 ;
        RECT 391.925 21.540 392.155 22.335 ;
        RECT 394.310 21.540 394.650 22.425 ;
        RECT 395.285 21.540 395.515 22.285 ;
        RECT 397.525 21.540 397.755 22.285 ;
        RECT 399.765 21.540 399.995 22.285 ;
        RECT 402.005 21.540 402.235 22.285 ;
        RECT 404.245 21.540 404.475 22.285 ;
        RECT 406.485 21.540 406.715 22.285 ;
        RECT 408.725 21.540 408.955 22.285 ;
        RECT 410.965 21.540 411.195 22.285 ;
        RECT 413.205 21.540 413.435 22.325 ;
        RECT 415.445 21.540 415.675 22.325 ;
        RECT 419.545 21.540 419.775 22.105 ;
        RECT 422.945 21.540 423.175 22.105 ;
        RECT 426.250 21.540 426.590 22.290 ;
        RECT 428.490 21.540 428.830 22.335 ;
        RECT 433.510 21.540 433.850 22.425 ;
        RECT 435.825 21.540 436.055 22.105 ;
        RECT 438.405 21.540 438.635 22.185 ;
        RECT 440.645 21.540 440.875 22.330 ;
        RECT 443.465 21.540 443.805 22.115 ;
        RECT 446.820 21.540 447.050 22.370 ;
        RECT 452.350 21.540 452.690 22.155 ;
        RECT 457.610 21.540 457.950 22.315 ;
        RECT 459.465 21.540 459.810 22.290 ;
        RECT 461.530 21.540 461.870 22.430 ;
        RECT 295.920 20.940 463.040 21.540 ;
        RECT 296.290 20.050 296.630 20.940 ;
        RECT 298.520 20.475 298.750 20.940 ;
        RECT 300.305 20.190 300.645 20.940 ;
        RECT 309.405 20.165 309.745 20.940 ;
        RECT 313.710 20.165 314.050 20.940 ;
        RECT 315.550 20.190 315.890 20.940 ;
        RECT 317.445 20.155 317.675 20.940 ;
        RECT 319.685 20.155 319.915 20.940 ;
        RECT 323.045 20.475 323.275 20.940 ;
        RECT 326.425 20.475 326.655 20.940 ;
        RECT 327.525 20.155 327.755 20.940 ;
        RECT 329.765 20.155 329.995 20.940 ;
        RECT 332.005 20.145 332.235 20.940 ;
        RECT 335.510 20.055 335.850 20.940 ;
        RECT 336.485 20.195 336.715 20.940 ;
        RECT 338.725 20.195 338.955 20.940 ;
        RECT 340.965 20.195 341.195 20.940 ;
        RECT 343.205 20.195 343.435 20.940 ;
        RECT 345.445 20.195 345.675 20.940 ;
        RECT 347.685 20.195 347.915 20.940 ;
        RECT 349.925 20.195 350.155 20.940 ;
        RECT 352.165 20.195 352.395 20.940 ;
        RECT 354.405 20.170 354.635 20.940 ;
        RECT 356.645 20.170 356.875 20.940 ;
        RECT 358.885 20.170 359.115 20.940 ;
        RECT 361.125 20.170 361.355 20.940 ;
        RECT 366.385 20.375 366.615 20.940 ;
        RECT 369.925 20.200 370.155 20.940 ;
        RECT 370.645 20.145 370.875 20.940 ;
        RECT 374.710 20.055 375.050 20.940 ;
        RECT 375.685 20.155 375.915 20.940 ;
        RECT 377.925 20.155 378.155 20.940 ;
        RECT 381.460 20.335 381.690 20.940 ;
        RECT 385.540 20.515 385.770 20.940 ;
        RECT 386.325 20.145 386.555 20.940 ;
        RECT 390.190 20.190 390.535 20.940 ;
        RECT 392.050 20.165 392.390 20.940 ;
        RECT 397.310 20.325 397.650 20.940 ;
        RECT 402.950 20.110 403.180 20.940 ;
        RECT 406.195 20.365 406.535 20.940 ;
        RECT 408.165 20.155 408.395 20.940 ;
        RECT 410.405 20.155 410.635 20.940 ;
        RECT 413.910 20.055 414.250 20.940 ;
        RECT 415.285 20.150 415.515 20.940 ;
        RECT 417.525 20.295 417.755 20.940 ;
        RECT 418.245 20.155 418.475 20.940 ;
        RECT 420.485 20.155 420.715 20.940 ;
        RECT 422.725 20.145 422.955 20.940 ;
        RECT 425.525 20.295 425.755 20.940 ;
        RECT 427.765 20.150 427.995 20.940 ;
        RECT 430.670 20.390 430.900 20.940 ;
        RECT 433.150 20.415 433.380 20.940 ;
        RECT 433.925 20.475 434.155 20.940 ;
        RECT 437.305 20.475 437.535 20.940 ;
        RECT 438.350 20.475 438.690 20.940 ;
        RECT 440.590 20.475 440.930 20.940 ;
        RECT 442.830 20.475 443.170 20.940 ;
        RECT 445.070 20.475 445.410 20.940 ;
        RECT 447.310 20.475 447.650 20.940 ;
        RECT 449.550 20.475 449.890 20.940 ;
        RECT 451.790 20.475 452.130 20.940 ;
        RECT 453.110 20.055 453.450 20.940 ;
        RECT 454.085 20.145 454.315 20.940 ;
        RECT 457.050 20.190 457.390 20.940 ;
        RECT 459.290 20.145 459.630 20.940 ;
        RECT 461.530 20.050 461.870 20.940 ;
        RECT 296.290 13.700 296.630 14.590 ;
        RECT 297.630 13.700 297.970 14.165 ;
        RECT 299.870 13.700 300.210 14.165 ;
        RECT 302.110 13.700 302.450 14.165 ;
        RECT 304.350 13.700 304.690 14.165 ;
        RECT 306.590 13.700 306.930 14.165 ;
        RECT 308.830 13.700 309.170 14.165 ;
        RECT 311.070 13.700 311.410 14.165 ;
        RECT 315.910 13.700 316.250 14.585 ;
        RECT 316.885 13.700 317.115 14.495 ;
        RECT 319.685 13.700 319.915 14.345 ;
        RECT 321.925 13.700 322.155 14.490 ;
        RECT 325.125 13.700 325.355 14.490 ;
        RECT 327.365 13.700 327.595 14.345 ;
        RECT 328.085 13.700 328.315 14.470 ;
        RECT 330.325 13.700 330.555 14.470 ;
        RECT 332.565 13.700 332.795 14.470 ;
        RECT 334.805 13.700 335.035 14.470 ;
        RECT 337.045 13.700 337.275 14.485 ;
        RECT 339.285 13.700 339.515 14.485 ;
        RECT 341.525 13.700 341.755 14.165 ;
        RECT 344.905 13.700 345.135 14.165 ;
        RECT 346.005 13.700 346.235 14.470 ;
        RECT 348.245 13.700 348.475 14.470 ;
        RECT 350.485 13.700 350.715 14.470 ;
        RECT 352.725 13.700 352.955 14.470 ;
        RECT 355.110 13.700 355.450 14.585 ;
        RECT 356.085 13.700 356.315 14.485 ;
        RECT 358.325 13.700 358.555 14.485 ;
        RECT 360.565 13.700 360.795 14.495 ;
        RECT 364.430 13.700 364.775 14.450 ;
        RECT 366.290 13.700 366.630 14.475 ;
        RECT 371.550 13.700 371.890 14.315 ;
        RECT 377.190 13.700 377.420 14.530 ;
        RECT 380.435 13.700 380.775 14.275 ;
        RECT 382.405 13.700 382.635 14.470 ;
        RECT 384.645 13.700 384.875 14.470 ;
        RECT 386.885 13.700 387.115 14.470 ;
        RECT 389.125 13.700 389.355 14.470 ;
        RECT 394.310 13.700 394.650 14.585 ;
        RECT 396.625 13.700 396.855 14.265 ;
        RECT 398.710 13.700 398.940 14.125 ;
        RECT 402.790 13.700 403.020 14.305 ;
        RECT 405.310 13.700 405.655 14.450 ;
        RECT 407.170 13.700 407.510 14.475 ;
        RECT 412.430 13.700 412.770 14.315 ;
        RECT 418.070 13.700 418.300 14.530 ;
        RECT 421.315 13.700 421.655 14.275 ;
        RECT 423.450 13.700 423.790 14.450 ;
        RECT 425.690 13.700 426.030 14.495 ;
        RECT 429.105 13.700 429.335 14.265 ;
        RECT 431.125 13.700 431.355 14.495 ;
        RECT 433.510 13.700 433.850 14.585 ;
        RECT 434.485 13.700 434.715 14.165 ;
        RECT 437.865 13.700 438.095 14.165 ;
        RECT 438.965 13.700 439.195 14.495 ;
        RECT 443.465 13.700 443.805 14.275 ;
        RECT 446.820 13.700 447.050 14.530 ;
        RECT 452.350 13.700 452.690 14.315 ;
        RECT 457.610 13.700 457.950 14.475 ;
        RECT 459.465 13.700 459.810 14.450 ;
        RECT 461.530 13.700 461.870 14.590 ;
        RECT 295.920 13.100 463.040 13.700 ;
        RECT 296.290 12.210 296.630 13.100 ;
        RECT 297.285 12.315 297.515 13.100 ;
        RECT 299.525 12.315 299.755 13.100 ;
        RECT 301.765 12.305 301.995 13.100 ;
        RECT 309.065 12.635 309.295 13.100 ;
        RECT 311.230 12.640 311.570 13.100 ;
        RECT 313.470 12.640 313.810 13.100 ;
        RECT 316.810 12.640 317.150 13.100 ;
        RECT 319.570 12.640 319.910 13.100 ;
        RECT 328.085 12.470 328.315 13.100 ;
        RECT 329.205 12.315 329.435 13.100 ;
        RECT 331.445 12.315 331.675 13.100 ;
        RECT 335.510 12.215 335.850 13.100 ;
        RECT 336.485 12.315 336.715 13.100 ;
        RECT 338.725 12.315 338.955 13.100 ;
        RECT 342.200 12.635 342.430 13.100 ;
        RECT 343.985 12.350 344.325 13.100 ;
        RECT 353.085 12.325 353.425 13.100 ;
        RECT 357.390 12.325 357.730 13.100 ;
        RECT 359.230 12.350 359.570 13.100 ;
        RECT 361.125 12.315 361.355 13.100 ;
        RECT 363.365 12.315 363.595 13.100 ;
        RECT 368.190 12.475 368.530 13.100 ;
        RECT 371.550 12.475 371.890 13.100 ;
        RECT 374.710 12.215 375.050 13.100 ;
        RECT 375.685 12.315 375.915 13.100 ;
        RECT 377.925 12.315 378.155 13.100 ;
        RECT 380.165 12.305 380.395 13.100 ;
        RECT 383.690 12.350 384.030 13.100 ;
        RECT 385.930 12.305 386.270 13.100 ;
        RECT 389.470 12.475 389.810 13.100 ;
        RECT 391.300 12.580 391.660 13.100 ;
        RECT 393.540 12.580 393.900 13.100 ;
        RECT 395.780 12.580 396.140 13.100 ;
        RECT 396.965 12.315 397.195 13.100 ;
        RECT 399.205 12.315 399.435 13.100 ;
        RECT 403.125 12.360 403.355 13.100 ;
        RECT 406.830 12.475 407.170 13.100 ;
        RECT 410.965 12.305 411.195 13.100 ;
        RECT 413.910 12.215 414.250 13.100 ;
        RECT 414.885 12.330 415.115 13.100 ;
        RECT 417.125 12.330 417.355 13.100 ;
        RECT 419.365 12.330 419.595 13.100 ;
        RECT 421.605 12.330 421.835 13.100 ;
        RECT 423.845 12.305 424.075 13.100 ;
        RECT 427.765 12.315 427.995 13.100 ;
        RECT 430.005 12.315 430.235 13.100 ;
        RECT 433.980 12.575 434.210 13.100 ;
        RECT 436.460 12.550 436.690 13.100 ;
        RECT 438.350 12.635 438.690 13.100 ;
        RECT 440.590 12.635 440.930 13.100 ;
        RECT 442.830 12.635 443.170 13.100 ;
        RECT 445.070 12.635 445.410 13.100 ;
        RECT 447.310 12.635 447.650 13.100 ;
        RECT 449.550 12.635 449.890 13.100 ;
        RECT 451.790 12.635 452.130 13.100 ;
        RECT 453.110 12.215 453.450 13.100 ;
        RECT 454.085 12.315 454.315 13.100 ;
        RECT 456.325 12.315 456.555 13.100 ;
        RECT 458.565 12.305 458.795 13.100 ;
        RECT 461.530 12.210 461.870 13.100 ;
        RECT 229.360 10.685 229.590 11.170 ;
        RECT 229.360 10.620 231.160 10.685 ;
        RECT 229.210 10.455 231.160 10.620 ;
        RECT 229.210 9.720 229.590 10.455 ;
        RECT 229.360 6.325 229.590 9.720 ;
        RECT 229.360 6.260 231.160 6.325 ;
        RECT 229.210 6.095 231.160 6.260 ;
        RECT 229.210 5.360 229.590 6.095 ;
        RECT 296.290 5.860 296.630 6.750 ;
        RECT 298.350 5.860 298.690 6.485 ;
        RECT 302.830 5.860 303.170 6.485 ;
        RECT 306.370 5.860 306.710 6.655 ;
        RECT 308.610 5.860 308.950 6.610 ;
        RECT 309.660 5.860 309.890 6.385 ;
        RECT 312.140 5.860 312.370 6.410 ;
        RECT 315.910 5.860 316.250 6.745 ;
        RECT 316.885 5.860 317.115 6.325 ;
        RECT 320.265 5.860 320.495 6.325 ;
        RECT 321.370 5.860 321.600 6.365 ;
        RECT 324.165 5.860 324.395 6.655 ;
        RECT 328.590 5.860 328.930 6.320 ;
        RECT 330.830 5.860 331.170 6.320 ;
        RECT 334.170 5.860 335.250 6.320 ;
        RECT 337.315 5.860 337.675 6.320 ;
        RECT 340.485 5.860 340.825 6.195 ;
        RECT 341.525 5.860 341.755 6.655 ;
        RECT 344.165 5.860 344.395 6.650 ;
        RECT 346.405 5.860 346.635 6.505 ;
        RECT 347.125 5.860 347.355 6.645 ;
        RECT 349.365 5.860 349.595 6.645 ;
        RECT 351.605 5.860 351.835 6.655 ;
        RECT 355.110 5.860 355.450 6.745 ;
        RECT 356.085 5.860 356.315 6.630 ;
        RECT 358.325 5.860 358.555 6.630 ;
        RECT 360.565 5.860 360.795 6.630 ;
        RECT 362.805 5.860 363.035 6.630 ;
        RECT 365.045 5.860 365.275 6.655 ;
        RECT 369.470 5.860 369.815 6.610 ;
        RECT 371.330 5.860 371.670 6.635 ;
        RECT 376.590 5.860 376.930 6.475 ;
        RECT 382.230 5.860 382.460 6.690 ;
        RECT 385.475 5.860 385.815 6.350 ;
        RECT 387.715 5.860 388.055 6.350 ;
        RECT 390.645 5.860 390.875 6.650 ;
        RECT 392.885 5.860 393.115 6.505 ;
        RECT 394.310 5.860 394.650 6.745 ;
        RECT 397.525 5.860 397.755 6.655 ;
        RECT 400.390 5.860 400.620 6.285 ;
        RECT 404.470 5.860 404.700 6.465 ;
        RECT 406.485 5.860 406.715 6.600 ;
        RECT 409.790 5.860 410.135 6.610 ;
        RECT 411.650 5.860 411.990 6.635 ;
        RECT 416.910 5.860 417.250 6.475 ;
        RECT 422.550 5.860 422.780 6.690 ;
        RECT 425.795 5.860 426.135 6.435 ;
        RECT 427.765 5.860 427.995 6.645 ;
        RECT 430.005 5.860 430.235 6.645 ;
        RECT 433.510 5.860 433.850 6.745 ;
        RECT 434.485 5.860 434.715 6.325 ;
        RECT 437.865 5.860 438.095 6.325 ;
        RECT 440.210 5.860 440.550 6.655 ;
        RECT 442.450 5.860 442.790 6.610 ;
        RECT 443.445 5.860 443.675 6.655 ;
        RECT 446.750 5.860 447.090 6.325 ;
        RECT 448.990 5.860 449.330 6.325 ;
        RECT 451.230 5.860 451.570 6.325 ;
        RECT 453.470 5.860 453.810 6.325 ;
        RECT 455.710 5.860 456.050 6.325 ;
        RECT 457.950 5.860 458.290 6.325 ;
        RECT 460.190 5.860 460.530 6.325 ;
        RECT 461.530 5.860 461.870 6.750 ;
        RECT 229.360 4.080 229.590 5.360 ;
        RECT 295.920 5.260 463.040 5.860 ;
        RECT 296.290 4.370 296.630 5.260 ;
        RECT 300.810 4.510 301.150 5.260 ;
        RECT 303.050 4.465 303.390 5.260 ;
        RECT 307.310 4.800 307.650 5.260 ;
        RECT 309.550 4.800 309.890 5.260 ;
        RECT 312.890 4.800 313.970 5.260 ;
        RECT 316.035 4.800 316.395 5.260 ;
        RECT 319.205 4.925 319.545 5.260 ;
        RECT 320.805 4.520 321.035 5.260 ;
        RECT 330.670 4.635 331.010 5.260 ;
        RECT 332.565 4.465 332.795 5.260 ;
        RECT 335.510 4.375 335.850 5.260 ;
        RECT 336.485 4.475 336.715 5.260 ;
        RECT 338.725 4.475 338.955 5.260 ;
        RECT 340.965 4.465 341.195 5.260 ;
        RECT 343.370 4.510 343.710 5.260 ;
        RECT 345.610 4.465 345.950 5.260 ;
        RECT 349.205 4.520 349.435 5.260 ;
        RECT 352.165 4.465 352.395 5.260 ;
        RECT 356.590 4.510 356.935 5.260 ;
        RECT 358.450 4.485 358.790 5.260 ;
        RECT 363.710 4.645 364.050 5.260 ;
        RECT 369.350 4.430 369.580 5.260 ;
        RECT 372.595 4.685 372.935 5.260 ;
        RECT 374.710 4.375 375.050 5.260 ;
        RECT 375.685 4.490 375.915 5.260 ;
        RECT 377.925 4.490 378.155 5.260 ;
        RECT 380.165 4.490 380.395 5.260 ;
        RECT 382.405 4.490 382.635 5.260 ;
        RECT 387.665 4.695 387.895 5.260 ;
        RECT 391.700 4.740 392.060 5.260 ;
        RECT 393.940 4.740 394.300 5.260 ;
        RECT 396.180 4.740 396.540 5.260 ;
        RECT 396.910 4.905 397.250 5.260 ;
        RECT 399.150 4.905 399.490 5.260 ;
        RECT 401.390 4.905 401.730 5.260 ;
        RECT 403.630 4.905 403.970 5.260 ;
        RECT 405.870 4.905 406.210 5.260 ;
        RECT 408.110 4.905 408.450 5.260 ;
        RECT 410.350 4.905 410.690 5.260 ;
        RECT 411.525 4.465 411.755 5.260 ;
        RECT 413.910 4.375 414.250 5.260 ;
        RECT 414.885 4.490 415.115 5.260 ;
        RECT 417.125 4.490 417.355 5.260 ;
        RECT 419.365 4.490 419.595 5.260 ;
        RECT 421.605 4.490 421.835 5.260 ;
        RECT 423.845 4.465 424.075 5.260 ;
        RECT 427.310 4.710 427.540 5.260 ;
        RECT 429.790 4.735 430.020 5.260 ;
        RECT 430.945 4.795 431.175 5.260 ;
        RECT 434.325 4.795 434.555 5.260 ;
        RECT 435.045 4.615 435.275 5.260 ;
        RECT 437.285 4.470 437.515 5.260 ;
        RECT 438.350 4.795 438.690 5.260 ;
        RECT 440.590 4.795 440.930 5.260 ;
        RECT 442.830 4.795 443.170 5.260 ;
        RECT 445.070 4.795 445.410 5.260 ;
        RECT 447.310 4.795 447.650 5.260 ;
        RECT 449.550 4.795 449.890 5.260 ;
        RECT 451.790 4.795 452.130 5.260 ;
        RECT 453.110 4.375 453.450 5.260 ;
        RECT 455.330 4.465 455.670 5.260 ;
        RECT 457.570 4.510 457.910 5.260 ;
        RECT 458.565 4.465 458.795 5.260 ;
        RECT 461.530 4.370 461.870 5.260 ;
        RECT 229.210 3.345 229.590 4.080 ;
        RECT 229.210 3.180 231.160 3.345 ;
        RECT 229.360 3.115 231.160 3.180 ;
        RECT 183.415 1.385 183.795 2.285 ;
        RECT 185.905 1.310 186.805 1.690 ;
        RECT 185.920 0.685 186.790 1.310 ;
        RECT 229.360 -0.280 229.590 3.115 ;
        RECT 185.920 -1.310 186.790 -0.685 ;
        RECT 229.210 -1.015 229.590 -0.280 ;
        RECT 229.210 -1.180 231.160 -1.015 ;
        RECT 229.360 -1.245 231.160 -1.180 ;
        RECT 183.415 -2.285 183.795 -1.385 ;
        RECT 185.905 -1.690 186.805 -1.310 ;
        RECT 229.360 -1.730 229.590 -1.245 ;
        RECT 296.290 -1.980 296.630 -1.090 ;
        RECT 297.285 -1.980 297.515 -1.195 ;
        RECT 299.525 -1.980 299.755 -1.195 ;
        RECT 302.100 -1.980 302.460 -1.460 ;
        RECT 304.340 -1.980 304.700 -1.460 ;
        RECT 306.580 -1.980 306.940 -1.460 ;
        RECT 307.365 -1.980 307.595 -1.195 ;
        RECT 309.605 -1.980 309.835 -1.195 ;
        RECT 311.845 -1.980 312.075 -1.185 ;
        RECT 315.910 -1.980 316.250 -1.095 ;
        RECT 317.845 -1.980 318.075 -1.350 ;
        RECT 324.165 -1.980 324.395 -1.185 ;
        RECT 329.150 -1.980 329.495 -1.230 ;
        RECT 331.010 -1.980 331.350 -1.205 ;
        RECT 336.270 -1.980 336.610 -1.365 ;
        RECT 341.910 -1.980 342.140 -1.150 ;
        RECT 345.155 -1.980 345.495 -1.405 ;
        RECT 348.190 -1.980 348.530 -1.645 ;
        RECT 355.110 -1.980 355.450 -1.095 ;
        RECT 357.150 -1.980 357.490 -1.355 ;
        RECT 361.125 -1.980 361.355 -1.515 ;
        RECT 364.505 -1.980 364.735 -1.515 ;
        RECT 365.605 -1.980 365.835 -1.185 ;
        RECT 368.225 -1.980 368.455 -1.515 ;
        RECT 371.605 -1.980 371.835 -1.515 ;
        RECT 372.325 -1.980 372.555 -1.210 ;
        RECT 374.565 -1.980 374.795 -1.210 ;
        RECT 376.805 -1.980 377.035 -1.210 ;
        RECT 379.045 -1.980 379.275 -1.210 ;
        RECT 381.845 -1.980 382.075 -1.120 ;
        RECT 385.245 -1.980 385.585 -1.515 ;
        RECT 387.580 -1.980 387.920 -1.515 ;
        RECT 390.845 -1.980 391.185 -1.515 ;
        RECT 393.180 -1.980 393.520 -1.515 ;
        RECT 394.310 -1.980 394.650 -1.095 ;
        RECT 395.685 -1.980 395.915 -1.240 ;
        RECT 397.925 -1.980 398.155 -1.240 ;
        RECT 398.820 -1.980 399.180 -1.645 ;
        RECT 402.965 -1.980 403.195 -1.375 ;
        RECT 405.925 -1.980 406.155 -1.185 ;
        RECT 408.165 -1.980 408.395 -1.330 ;
        RECT 410.435 -1.980 410.665 -1.330 ;
        RECT 413.045 -1.980 413.275 -1.120 ;
        RECT 416.045 -1.980 416.385 -1.515 ;
        RECT 418.380 -1.980 418.720 -1.515 ;
        RECT 419.365 -1.980 419.595 -1.210 ;
        RECT 421.605 -1.980 421.835 -1.210 ;
        RECT 423.845 -1.980 424.075 -1.210 ;
        RECT 426.085 -1.980 426.315 -1.210 ;
        RECT 428.325 -1.980 428.555 -1.195 ;
        RECT 430.565 -1.980 430.795 -1.195 ;
        RECT 433.510 -1.980 433.850 -1.095 ;
        RECT 434.485 -1.980 434.715 -1.335 ;
        RECT 436.725 -1.980 436.955 -1.190 ;
        RECT 437.900 -1.980 438.130 -1.455 ;
        RECT 440.380 -1.980 440.610 -1.430 ;
        RECT 443.465 -1.980 443.805 -1.405 ;
        RECT 446.820 -1.980 447.050 -1.150 ;
        RECT 452.350 -1.980 452.690 -1.365 ;
        RECT 457.610 -1.980 457.950 -1.205 ;
        RECT 459.465 -1.980 459.810 -1.230 ;
        RECT 461.530 -1.980 461.870 -1.090 ;
        RECT 295.920 -2.580 463.040 -1.980 ;
        RECT 296.290 -3.470 296.630 -2.580 ;
        RECT 298.350 -3.330 298.690 -2.580 ;
        RECT 300.190 -3.355 300.530 -2.580 ;
        RECT 304.495 -3.355 304.835 -2.580 ;
        RECT 313.595 -3.330 313.935 -2.580 ;
        RECT 315.490 -3.045 315.720 -2.580 ;
        RECT 319.520 -3.085 319.750 -2.580 ;
        RECT 323.605 -3.210 323.835 -2.580 ;
        RECT 326.800 -3.085 327.030 -2.580 ;
        RECT 332.005 -3.375 332.235 -2.580 ;
        RECT 335.510 -3.465 335.850 -2.580 ;
        RECT 337.950 -3.205 338.290 -2.580 ;
        RECT 339.845 -3.365 340.075 -2.580 ;
        RECT 342.085 -3.365 342.315 -2.580 ;
        RECT 348.285 -3.370 348.515 -2.580 ;
        RECT 352.005 -3.320 352.235 -2.580 ;
        RECT 352.725 -3.365 352.955 -2.580 ;
        RECT 354.965 -3.365 355.195 -2.580 ;
        RECT 357.205 -3.375 357.435 -2.580 ;
        RECT 361.070 -3.100 361.410 -2.580 ;
        RECT 363.310 -3.100 363.650 -2.580 ;
        RECT 365.605 -3.375 365.835 -2.580 ;
        RECT 368.805 -3.370 369.035 -2.580 ;
        RECT 371.045 -3.225 371.275 -2.580 ;
        RECT 371.765 -3.375 371.995 -2.580 ;
        RECT 374.710 -3.465 375.050 -2.580 ;
        RECT 375.685 -3.365 375.915 -2.580 ;
        RECT 377.925 -3.365 378.155 -2.580 ;
        RECT 381.845 -3.225 382.075 -2.580 ;
        RECT 384.085 -3.370 384.315 -2.580 ;
        RECT 385.150 -2.935 385.490 -2.580 ;
        RECT 387.390 -2.935 387.730 -2.580 ;
        RECT 389.630 -2.935 389.970 -2.580 ;
        RECT 391.870 -2.935 392.210 -2.580 ;
        RECT 394.110 -2.935 394.450 -2.580 ;
        RECT 396.350 -2.935 396.690 -2.580 ;
        RECT 398.590 -2.935 398.930 -2.580 ;
        RECT 399.845 -3.110 400.075 -2.580 ;
        RECT 408.005 -3.110 408.235 -2.580 ;
        RECT 409.885 -3.045 410.225 -2.580 ;
        RECT 412.220 -3.045 412.560 -2.580 ;
        RECT 413.910 -3.465 414.250 -2.580 ;
        RECT 416.970 -2.915 417.310 -2.580 ;
        RECT 421.050 -2.915 421.390 -2.580 ;
        RECT 436.345 -3.145 436.575 -2.580 ;
        RECT 438.350 -3.045 438.690 -2.580 ;
        RECT 440.590 -3.045 440.930 -2.580 ;
        RECT 442.830 -3.045 443.170 -2.580 ;
        RECT 445.070 -3.045 445.410 -2.580 ;
        RECT 447.310 -3.045 447.650 -2.580 ;
        RECT 449.550 -3.045 449.890 -2.580 ;
        RECT 451.790 -3.045 452.130 -2.580 ;
        RECT 453.110 -3.465 453.450 -2.580 ;
        RECT 454.085 -3.375 454.315 -2.580 ;
        RECT 458.130 -3.375 458.470 -2.580 ;
        RECT 460.370 -3.330 460.710 -2.580 ;
        RECT 461.530 -3.470 461.870 -2.580 ;
        RECT 296.290 -9.820 296.630 -8.930 ;
        RECT 297.630 -9.820 297.970 -9.355 ;
        RECT 299.870 -9.820 300.210 -9.355 ;
        RECT 302.110 -9.820 302.450 -9.355 ;
        RECT 304.350 -9.820 304.690 -9.355 ;
        RECT 306.590 -9.820 306.930 -9.355 ;
        RECT 308.830 -9.820 309.170 -9.355 ;
        RECT 311.070 -9.820 311.410 -9.355 ;
        RECT 311.845 -9.820 312.075 -9.025 ;
        RECT 315.910 -9.820 316.250 -8.935 ;
        RECT 316.885 -9.820 317.115 -9.025 ;
        RECT 321.870 -9.820 322.215 -9.070 ;
        RECT 323.730 -9.820 324.070 -9.045 ;
        RECT 328.990 -9.820 329.330 -9.205 ;
        RECT 334.630 -9.820 334.860 -8.990 ;
        RECT 337.875 -9.820 338.215 -9.245 ;
        RECT 339.845 -9.820 340.075 -9.050 ;
        RECT 342.085 -9.820 342.315 -9.050 ;
        RECT 344.325 -9.820 344.555 -9.050 ;
        RECT 346.565 -9.820 346.795 -9.050 ;
        RECT 348.805 -9.820 349.035 -9.035 ;
        RECT 351.045 -9.820 351.275 -9.035 ;
        RECT 355.110 -9.820 355.450 -8.935 ;
        RECT 356.085 -9.820 356.315 -9.035 ;
        RECT 358.325 -9.820 358.555 -9.035 ;
        RECT 361.525 -9.820 361.755 -9.030 ;
        RECT 363.765 -9.820 363.995 -9.175 ;
        RECT 364.595 -9.820 364.825 -9.060 ;
        RECT 367.000 -9.820 367.340 -9.355 ;
        RECT 369.680 -9.820 370.020 -9.355 ;
        RECT 372.360 -9.820 372.700 -9.410 ;
        RECT 375.040 -9.820 375.380 -9.355 ;
        RECT 379.120 -9.820 379.460 -9.480 ;
        RECT 383.440 -9.820 383.780 -9.410 ;
        RECT 384.865 -9.820 385.095 -9.425 ;
        RECT 387.050 -9.820 387.390 -9.480 ;
        RECT 389.525 -9.820 389.755 -9.430 ;
        RECT 393.445 -9.820 393.675 -9.210 ;
        RECT 394.310 -9.820 394.650 -8.935 ;
        RECT 398.150 -9.820 398.380 -9.355 ;
        RECT 400.335 -9.820 400.675 -9.480 ;
        RECT 404.490 -9.820 404.720 -9.355 ;
        RECT 405.540 -9.820 405.900 -9.485 ;
        RECT 409.685 -9.820 409.915 -9.215 ;
        RECT 412.770 -9.820 413.110 -9.025 ;
        RECT 415.010 -9.820 415.350 -9.070 ;
        RECT 416.005 -9.820 416.235 -9.025 ;
        RECT 419.520 -9.820 419.860 -9.355 ;
        RECT 421.855 -9.820 422.195 -9.355 ;
        RECT 424.010 -9.820 424.350 -9.070 ;
        RECT 426.250 -9.820 426.590 -9.025 ;
        RECT 429.390 -9.820 429.730 -9.195 ;
        RECT 433.510 -9.820 433.850 -8.935 ;
        RECT 434.485 -9.820 434.715 -9.025 ;
        RECT 439.525 -9.820 439.755 -9.025 ;
        RECT 443.390 -9.820 443.735 -9.070 ;
        RECT 445.250 -9.820 445.590 -9.045 ;
        RECT 450.510 -9.820 450.850 -9.205 ;
        RECT 456.150 -9.820 456.380 -8.990 ;
        RECT 459.395 -9.820 459.735 -9.245 ;
        RECT 461.530 -9.820 461.870 -8.930 ;
        RECT 295.920 -10.420 463.040 -9.820 ;
        RECT 231.225 -12.135 231.455 -10.565 ;
        RECT 234.740 -12.135 234.970 -10.565 ;
        RECT 296.290 -11.310 296.630 -10.420 ;
        RECT 297.630 -10.885 297.970 -10.420 ;
        RECT 299.870 -10.885 300.210 -10.420 ;
        RECT 302.110 -10.885 302.450 -10.420 ;
        RECT 304.350 -10.885 304.690 -10.420 ;
        RECT 306.590 -10.885 306.930 -10.420 ;
        RECT 308.830 -10.885 309.170 -10.420 ;
        RECT 311.070 -10.885 311.410 -10.420 ;
        RECT 311.845 -11.165 312.075 -10.420 ;
        RECT 314.085 -11.165 314.315 -10.420 ;
        RECT 316.325 -11.165 316.555 -10.420 ;
        RECT 318.565 -11.165 318.795 -10.420 ;
        RECT 320.805 -11.165 321.035 -10.420 ;
        RECT 323.045 -11.165 323.275 -10.420 ;
        RECT 325.285 -11.165 325.515 -10.420 ;
        RECT 327.525 -11.165 327.755 -10.420 ;
        RECT 329.765 -11.205 329.995 -10.420 ;
        RECT 332.005 -11.205 332.235 -10.420 ;
        RECT 335.510 -11.305 335.850 -10.420 ;
        RECT 336.485 -11.190 336.715 -10.420 ;
        RECT 338.725 -11.190 338.955 -10.420 ;
        RECT 340.965 -11.190 341.195 -10.420 ;
        RECT 343.205 -11.190 343.435 -10.420 ;
        RECT 346.565 -10.955 346.795 -10.420 ;
        RECT 348.805 -10.955 349.035 -10.420 ;
        RECT 352.965 -10.955 353.195 -10.420 ;
        RECT 354.965 -11.205 355.195 -10.420 ;
        RECT 357.205 -11.205 357.435 -10.420 ;
        RECT 360.170 -11.170 360.510 -10.420 ;
        RECT 362.410 -11.215 362.750 -10.420 ;
        RECT 365.605 -10.955 365.835 -10.420 ;
        RECT 367.845 -10.955 368.075 -10.420 ;
        RECT 372.005 -10.955 372.235 -10.420 ;
        RECT 374.710 -11.305 375.050 -10.420 ;
        RECT 375.685 -11.215 375.915 -10.420 ;
        RECT 384.935 -10.755 385.275 -10.420 ;
        RECT 389.680 -10.880 390.020 -10.420 ;
        RECT 392.190 -10.880 392.530 -10.420 ;
        RECT 394.790 -10.880 395.130 -10.420 ;
        RECT 397.380 -10.880 397.720 -10.420 ;
        RECT 399.985 -10.880 400.325 -10.420 ;
        RECT 402.500 -10.880 402.840 -10.420 ;
        RECT 404.920 -10.880 405.260 -10.420 ;
        RECT 407.340 -10.880 407.680 -10.420 ;
        RECT 409.580 -10.880 409.920 -10.420 ;
        RECT 410.405 -11.065 410.635 -10.420 ;
        RECT 412.645 -11.210 412.875 -10.420 ;
        RECT 413.910 -11.305 414.250 -10.420 ;
        RECT 417.725 -10.885 418.065 -10.420 ;
        RECT 420.060 -10.885 420.400 -10.420 ;
        RECT 421.045 -11.205 421.275 -10.420 ;
        RECT 423.285 -11.205 423.515 -10.420 ;
        RECT 427.225 -10.995 427.565 -10.420 ;
        RECT 430.580 -11.250 430.810 -10.420 ;
        RECT 436.110 -11.035 436.450 -10.420 ;
        RECT 441.370 -11.195 441.710 -10.420 ;
        RECT 443.225 -11.170 443.570 -10.420 ;
        RECT 447.365 -11.205 447.595 -10.420 ;
        RECT 449.605 -11.205 449.835 -10.420 ;
        RECT 453.110 -11.305 453.450 -10.420 ;
        RECT 454.085 -11.205 454.315 -10.420 ;
        RECT 456.325 -11.205 456.555 -10.420 ;
        RECT 458.565 -11.215 458.795 -10.420 ;
        RECT 461.530 -11.310 461.870 -10.420 ;
        RECT 229.940 -12.365 231.940 -12.135 ;
        RECT 233.455 -12.365 235.455 -12.135 ;
        RECT 230.490 -12.515 231.390 -12.365 ;
        RECT 234.005 -12.515 234.905 -12.365 ;
        RECT 296.290 -17.660 296.630 -16.770 ;
        RECT 297.285 -17.660 297.515 -16.865 ;
        RECT 301.045 -17.660 301.275 -16.800 ;
        RECT 303.105 -17.660 303.335 -17.095 ;
        RECT 305.125 -17.660 305.355 -16.920 ;
        RECT 309.605 -17.660 309.835 -16.875 ;
        RECT 311.845 -17.660 312.075 -16.875 ;
        RECT 315.910 -17.660 316.250 -16.775 ;
        RECT 316.885 -17.660 317.115 -16.875 ;
        RECT 319.125 -17.660 319.355 -16.875 ;
        RECT 322.590 -17.660 322.820 -17.110 ;
        RECT 325.070 -17.660 325.300 -17.135 ;
        RECT 329.985 -17.660 330.215 -17.095 ;
        RECT 333.070 -17.660 333.415 -16.910 ;
        RECT 334.930 -17.660 335.270 -16.885 ;
        RECT 340.190 -17.660 340.530 -17.045 ;
        RECT 345.830 -17.660 346.060 -16.830 ;
        RECT 349.075 -17.660 349.415 -17.085 ;
        RECT 352.385 -17.660 352.615 -17.095 ;
        RECT 355.110 -17.660 355.450 -16.775 ;
        RECT 356.085 -17.660 356.315 -16.865 ;
        RECT 358.725 -17.660 358.955 -16.870 ;
        RECT 360.965 -17.660 361.195 -17.015 ;
        RECT 362.020 -17.660 362.380 -17.140 ;
        RECT 364.260 -17.660 364.620 -17.140 ;
        RECT 366.500 -17.660 366.860 -17.140 ;
        RECT 367.285 -17.660 367.515 -16.865 ;
        RECT 370.085 -17.660 370.315 -17.015 ;
        RECT 372.325 -17.660 372.555 -16.870 ;
        RECT 373.445 -17.660 373.675 -16.865 ;
        RECT 376.910 -17.660 377.140 -17.110 ;
        RECT 379.390 -17.660 379.620 -17.135 ;
        RECT 381.505 -17.660 381.735 -17.095 ;
        RECT 383.525 -17.660 383.755 -16.875 ;
        RECT 385.765 -17.660 385.995 -16.875 ;
        RECT 390.085 -17.660 390.315 -17.030 ;
        RECT 394.310 -17.660 394.650 -16.775 ;
        RECT 395.450 -17.660 395.790 -16.975 ;
        RECT 397.690 -17.660 398.030 -16.975 ;
        RECT 399.930 -17.660 400.270 -16.975 ;
        RECT 402.350 -17.660 402.690 -16.975 ;
        RECT 403.230 -17.660 403.570 -17.325 ;
        RECT 409.265 -17.660 409.495 -17.060 ;
        RECT 413.610 -17.660 413.950 -17.325 ;
        RECT 417.690 -17.660 418.030 -17.325 ;
        RECT 430.005 -17.660 430.235 -16.865 ;
        RECT 433.510 -17.660 433.850 -16.775 ;
        RECT 434.485 -17.660 434.715 -16.890 ;
        RECT 436.725 -17.660 436.955 -16.890 ;
        RECT 438.965 -17.660 439.195 -16.890 ;
        RECT 441.205 -17.660 441.435 -16.890 ;
        RECT 443.445 -17.660 443.675 -16.865 ;
        RECT 446.750 -17.660 447.090 -17.195 ;
        RECT 448.990 -17.660 449.330 -17.195 ;
        RECT 451.230 -17.660 451.570 -17.195 ;
        RECT 453.470 -17.660 453.810 -17.195 ;
        RECT 455.710 -17.660 456.050 -17.195 ;
        RECT 457.950 -17.660 458.290 -17.195 ;
        RECT 460.190 -17.660 460.530 -17.195 ;
        RECT 461.530 -17.660 461.870 -16.770 ;
        RECT 295.920 -18.260 463.040 -17.660 ;
        RECT 296.290 -19.150 296.630 -18.260 ;
        RECT 297.450 -19.010 297.790 -18.260 ;
        RECT 299.690 -19.055 300.030 -18.260 ;
        RECT 304.510 -19.010 304.855 -18.260 ;
        RECT 306.370 -19.035 306.710 -18.260 ;
        RECT 311.630 -18.875 311.970 -18.260 ;
        RECT 317.270 -19.090 317.500 -18.260 ;
        RECT 320.515 -18.835 320.855 -18.260 ;
        RECT 322.485 -18.725 322.715 -18.260 ;
        RECT 325.865 -18.725 326.095 -18.260 ;
        RECT 329.205 -19.045 329.435 -18.260 ;
        RECT 331.445 -19.045 331.675 -18.260 ;
        RECT 335.510 -19.145 335.850 -18.260 ;
        RECT 336.485 -19.005 336.715 -18.260 ;
        RECT 338.725 -19.005 338.955 -18.260 ;
        RECT 340.965 -19.005 341.195 -18.260 ;
        RECT 343.205 -19.005 343.435 -18.260 ;
        RECT 345.445 -19.005 345.675 -18.260 ;
        RECT 347.685 -19.005 347.915 -18.260 ;
        RECT 349.925 -19.005 350.155 -18.260 ;
        RECT 352.165 -19.005 352.395 -18.260 ;
        RECT 354.405 -19.030 354.635 -18.260 ;
        RECT 356.645 -19.030 356.875 -18.260 ;
        RECT 358.885 -19.030 359.115 -18.260 ;
        RECT 361.125 -19.030 361.355 -18.260 ;
        RECT 365.265 -18.655 365.495 -18.260 ;
        RECT 367.450 -18.600 367.790 -18.260 ;
        RECT 369.925 -18.650 370.155 -18.260 ;
        RECT 373.845 -18.870 374.075 -18.260 ;
        RECT 374.710 -19.145 375.050 -18.260 ;
        RECT 377.205 -19.120 377.435 -18.260 ;
        RECT 377.925 -19.055 378.155 -18.260 ;
        RECT 381.845 -18.865 382.075 -18.260 ;
        RECT 385.860 -18.595 386.220 -18.260 ;
        RECT 386.885 -19.055 387.115 -18.260 ;
        RECT 389.460 -18.780 389.820 -18.260 ;
        RECT 391.700 -18.780 392.060 -18.260 ;
        RECT 393.940 -18.780 394.300 -18.260 ;
        RECT 395.790 -18.595 396.130 -18.260 ;
        RECT 405.365 -19.055 405.595 -18.260 ;
        RECT 409.230 -18.780 409.570 -18.260 ;
        RECT 411.470 -18.780 411.810 -18.260 ;
        RECT 413.910 -19.145 414.250 -18.260 ;
        RECT 418.020 -18.615 418.380 -18.260 ;
        RECT 420.260 -18.615 420.620 -18.260 ;
        RECT 422.500 -18.615 422.860 -18.260 ;
        RECT 426.645 -19.055 426.875 -18.260 ;
        RECT 431.630 -18.885 431.970 -18.260 ;
        RECT 434.990 -19.010 435.335 -18.260 ;
        RECT 436.850 -19.035 437.190 -18.260 ;
        RECT 442.110 -18.875 442.450 -18.260 ;
        RECT 447.750 -19.090 447.980 -18.260 ;
        RECT 450.995 -18.835 451.335 -18.260 ;
        RECT 453.110 -19.145 453.450 -18.260 ;
        RECT 455.945 -18.825 456.175 -18.260 ;
        RECT 459.470 -18.885 459.810 -18.260 ;
        RECT 461.530 -19.150 461.870 -18.260 ;
        RECT 296.290 -25.500 296.630 -24.610 ;
        RECT 297.630 -25.500 297.970 -25.035 ;
        RECT 299.870 -25.500 300.210 -25.035 ;
        RECT 302.110 -25.500 302.450 -25.035 ;
        RECT 304.350 -25.500 304.690 -25.035 ;
        RECT 306.590 -25.500 306.930 -25.035 ;
        RECT 308.830 -25.500 309.170 -25.035 ;
        RECT 311.070 -25.500 311.410 -25.035 ;
        RECT 313.145 -25.500 313.375 -24.935 ;
        RECT 315.910 -25.500 316.250 -24.615 ;
        RECT 316.885 -25.500 317.115 -24.705 ;
        RECT 319.525 -25.500 319.755 -24.710 ;
        RECT 321.765 -25.500 321.995 -24.855 ;
        RECT 322.485 -25.500 322.715 -24.755 ;
        RECT 324.725 -25.500 324.955 -24.755 ;
        RECT 326.965 -25.500 327.195 -24.755 ;
        RECT 329.205 -25.500 329.435 -24.755 ;
        RECT 331.445 -25.500 331.675 -24.755 ;
        RECT 333.685 -25.500 333.915 -24.755 ;
        RECT 335.925 -25.500 336.155 -24.755 ;
        RECT 338.165 -25.500 338.395 -24.755 ;
        RECT 340.405 -25.500 340.635 -24.705 ;
        RECT 344.505 -25.500 344.735 -24.935 ;
        RECT 346.565 -25.500 346.795 -24.715 ;
        RECT 348.805 -25.500 349.035 -24.715 ;
        RECT 352.725 -25.500 352.955 -24.760 ;
        RECT 355.110 -25.500 355.450 -24.615 ;
        RECT 357.150 -25.500 357.490 -25.165 ;
        RECT 363.760 -25.500 363.990 -24.995 ;
        RECT 364.860 -25.500 365.200 -25.090 ;
        RECT 369.180 -25.500 369.520 -25.160 ;
        RECT 373.260 -25.500 373.600 -25.035 ;
        RECT 375.940 -25.500 376.280 -25.090 ;
        RECT 378.620 -25.500 378.960 -25.035 ;
        RECT 381.300 -25.500 381.640 -25.035 ;
        RECT 383.815 -25.500 384.045 -24.740 ;
        RECT 385.045 -25.500 385.275 -24.870 ;
        RECT 394.310 -25.500 394.650 -24.615 ;
        RECT 395.285 -25.500 395.515 -24.715 ;
        RECT 397.525 -25.500 397.755 -24.715 ;
        RECT 400.830 -25.500 401.175 -24.750 ;
        RECT 402.690 -25.500 403.030 -24.725 ;
        RECT 407.950 -25.500 408.290 -24.885 ;
        RECT 413.590 -25.500 413.820 -24.670 ;
        RECT 416.835 -25.500 417.175 -24.925 ;
        RECT 418.805 -25.500 419.035 -25.035 ;
        RECT 422.185 -25.500 422.415 -25.035 ;
        RECT 425.525 -25.500 425.755 -24.715 ;
        RECT 427.765 -25.500 427.995 -24.715 ;
        RECT 430.005 -25.500 430.235 -24.705 ;
        RECT 433.510 -25.500 433.850 -24.615 ;
        RECT 434.485 -25.500 434.715 -24.965 ;
        RECT 436.725 -25.500 436.955 -24.965 ;
        RECT 440.885 -25.500 441.115 -24.965 ;
        RECT 444.910 -25.500 445.250 -24.875 ;
        RECT 446.750 -25.500 447.090 -25.035 ;
        RECT 448.990 -25.500 449.330 -25.035 ;
        RECT 451.230 -25.500 451.570 -25.035 ;
        RECT 453.470 -25.500 453.810 -25.035 ;
        RECT 455.710 -25.500 456.050 -25.035 ;
        RECT 457.950 -25.500 458.290 -25.035 ;
        RECT 460.190 -25.500 460.530 -25.035 ;
        RECT 461.530 -25.500 461.870 -24.610 ;
        RECT 295.920 -26.100 463.040 -25.500 ;
        RECT 296.290 -26.990 296.630 -26.100 ;
        RECT 299.470 -26.850 299.815 -26.100 ;
        RECT 301.330 -26.875 301.670 -26.100 ;
        RECT 306.590 -26.715 306.930 -26.100 ;
        RECT 312.230 -26.930 312.460 -26.100 ;
        RECT 315.475 -26.675 315.815 -26.100 ;
        RECT 317.825 -26.565 318.055 -26.100 ;
        RECT 321.205 -26.565 321.435 -26.100 ;
        RECT 323.150 -26.650 323.380 -26.100 ;
        RECT 325.630 -26.625 325.860 -26.100 ;
        RECT 326.405 -26.870 326.635 -26.100 ;
        RECT 328.645 -26.870 328.875 -26.100 ;
        RECT 330.885 -26.870 331.115 -26.100 ;
        RECT 333.125 -26.870 333.355 -26.100 ;
        RECT 335.510 -26.985 335.850 -26.100 ;
        RECT 336.485 -26.870 336.715 -26.100 ;
        RECT 338.725 -26.870 338.955 -26.100 ;
        RECT 340.965 -26.870 341.195 -26.100 ;
        RECT 343.205 -26.870 343.435 -26.100 ;
        RECT 345.445 -26.895 345.675 -26.100 ;
        RECT 348.805 -26.840 349.035 -26.100 ;
        RECT 352.670 -26.435 353.010 -26.100 ;
        RECT 357.205 -26.885 357.435 -26.100 ;
        RECT 359.445 -26.885 359.675 -26.100 ;
        RECT 361.685 -26.895 361.915 -26.100 ;
        RECT 365.785 -26.665 366.015 -26.100 ;
        RECT 367.845 -26.885 368.075 -26.100 ;
        RECT 370.085 -26.885 370.315 -26.100 ;
        RECT 372.325 -26.895 372.555 -26.100 ;
        RECT 374.710 -26.985 375.050 -26.100 ;
        RECT 376.985 -26.665 377.215 -26.100 ;
        RECT 379.045 -26.885 379.275 -26.100 ;
        RECT 381.285 -26.885 381.515 -26.100 ;
        RECT 383.690 -26.850 384.030 -26.100 ;
        RECT 385.930 -26.895 386.270 -26.100 ;
        RECT 388.005 -26.885 388.235 -26.100 ;
        RECT 390.245 -26.885 390.475 -26.100 ;
        RECT 392.485 -26.895 392.715 -26.100 ;
        RECT 394.730 -26.605 394.960 -26.100 ;
        RECT 397.525 -26.895 397.755 -26.100 ;
        RECT 400.325 -26.565 400.555 -26.100 ;
        RECT 403.705 -26.565 403.935 -26.100 ;
        RECT 406.325 -26.840 406.555 -26.100 ;
        RECT 407.045 -26.885 407.275 -26.100 ;
        RECT 409.285 -26.885 409.515 -26.100 ;
        RECT 411.525 -26.895 411.755 -26.100 ;
        RECT 413.910 -26.985 414.250 -26.100 ;
        RECT 414.885 -26.895 415.115 -26.100 ;
        RECT 421.740 -26.605 421.970 -26.100 ;
        RECT 426.865 -26.665 427.095 -26.100 ;
        RECT 431.630 -26.725 431.970 -26.100 ;
        RECT 436.185 -26.565 436.415 -26.100 ;
        RECT 438.350 -26.565 438.690 -26.100 ;
        RECT 440.590 -26.565 440.930 -26.100 ;
        RECT 442.830 -26.565 443.170 -26.100 ;
        RECT 445.070 -26.565 445.410 -26.100 ;
        RECT 447.310 -26.565 447.650 -26.100 ;
        RECT 449.550 -26.565 449.890 -26.100 ;
        RECT 451.790 -26.565 452.130 -26.100 ;
        RECT 453.110 -26.985 453.450 -26.100 ;
        RECT 458.130 -26.895 458.470 -26.100 ;
        RECT 460.370 -26.850 460.710 -26.100 ;
        RECT 461.530 -26.990 461.870 -26.100 ;
        RECT 165.900 -32.905 166.130 -32.355 ;
        RECT 167.315 -32.555 167.695 -31.655 ;
        RECT 168.915 -32.555 169.295 -31.655 ;
        RECT 174.115 -32.555 174.495 -31.655 ;
        RECT 179.115 -32.555 179.495 -31.655 ;
        RECT 183.415 -32.555 183.795 -31.655 ;
        RECT 185.015 -32.555 185.395 -31.655 ;
        RECT 186.615 -32.555 186.995 -31.655 ;
        RECT 188.215 -32.555 188.595 -31.655 ;
        RECT 189.815 -32.555 190.195 -31.655 ;
        RECT 165.825 -33.805 166.205 -32.905 ;
        RECT 167.390 -33.790 167.620 -32.555 ;
        RECT 168.990 -33.790 169.220 -32.555 ;
        RECT 174.190 -33.790 174.420 -32.555 ;
        RECT 179.190 -33.790 179.420 -32.555 ;
        RECT 183.490 -33.790 183.720 -32.555 ;
        RECT 185.090 -33.790 185.320 -32.555 ;
        RECT 186.690 -33.790 186.920 -32.555 ;
        RECT 188.290 -33.790 188.520 -32.555 ;
        RECT 189.890 -33.790 190.120 -32.555 ;
        RECT 190.580 -32.905 190.810 -32.355 ;
        RECT 190.505 -33.805 190.885 -32.905 ;
        RECT 296.290 -33.340 296.630 -32.450 ;
        RECT 297.630 -33.340 297.970 -32.875 ;
        RECT 299.870 -33.340 300.210 -32.875 ;
        RECT 302.110 -33.340 302.450 -32.875 ;
        RECT 304.350 -33.340 304.690 -32.875 ;
        RECT 306.590 -33.340 306.930 -32.875 ;
        RECT 308.830 -33.340 309.170 -32.875 ;
        RECT 311.070 -33.340 311.410 -32.875 ;
        RECT 315.910 -33.340 316.250 -32.455 ;
        RECT 317.285 -33.340 317.515 -32.550 ;
        RECT 319.525 -33.340 319.755 -32.695 ;
        RECT 320.645 -33.340 320.875 -32.550 ;
        RECT 322.885 -33.340 323.115 -32.695 ;
        RECT 323.605 -33.340 323.835 -32.555 ;
        RECT 325.845 -33.340 326.075 -32.555 ;
        RECT 329.150 -33.340 329.495 -32.590 ;
        RECT 331.010 -33.340 331.350 -32.565 ;
        RECT 336.270 -33.340 336.610 -32.725 ;
        RECT 341.910 -33.340 342.140 -32.510 ;
        RECT 345.155 -33.340 345.495 -32.765 ;
        RECT 347.125 -33.340 347.355 -32.555 ;
        RECT 349.365 -33.340 349.595 -32.555 ;
        RECT 351.605 -33.340 351.835 -32.545 ;
        RECT 355.110 -33.340 355.450 -32.455 ;
        RECT 356.085 -33.340 356.315 -32.570 ;
        RECT 358.325 -33.340 358.555 -32.570 ;
        RECT 360.565 -33.340 360.795 -32.570 ;
        RECT 362.805 -33.340 363.035 -32.570 ;
        RECT 365.045 -33.340 365.275 -32.545 ;
        RECT 368.405 -33.340 368.635 -32.805 ;
        RECT 370.645 -33.340 370.875 -32.805 ;
        RECT 374.805 -33.340 375.035 -32.805 ;
        RECT 376.805 -33.340 377.035 -32.555 ;
        RECT 379.045 -33.340 379.275 -32.555 ;
        RECT 381.285 -33.340 381.515 -32.545 ;
        RECT 384.085 -33.340 384.315 -32.805 ;
        RECT 386.325 -33.340 386.555 -32.805 ;
        RECT 390.485 -33.340 390.715 -32.805 ;
        RECT 394.310 -33.340 394.650 -32.455 ;
        RECT 395.285 -33.340 395.515 -32.555 ;
        RECT 397.525 -33.340 397.755 -32.555 ;
        RECT 399.765 -33.340 399.995 -32.545 ;
        RECT 402.005 -33.340 402.235 -32.875 ;
        RECT 405.385 -33.340 405.615 -32.875 ;
        RECT 406.485 -33.340 406.715 -32.570 ;
        RECT 408.725 -33.340 408.955 -32.570 ;
        RECT 410.965 -33.340 411.195 -32.570 ;
        RECT 413.205 -33.340 413.435 -32.570 ;
        RECT 415.445 -33.340 415.675 -32.555 ;
        RECT 417.685 -33.340 417.915 -32.555 ;
        RECT 421.045 -33.340 421.275 -32.875 ;
        RECT 424.425 -33.340 424.655 -32.875 ;
        RECT 425.925 -33.340 426.155 -32.710 ;
        RECT 430.405 -33.340 430.635 -32.550 ;
        RECT 432.645 -33.340 432.875 -32.695 ;
        RECT 433.510 -33.340 433.850 -32.455 ;
        RECT 435.605 -33.340 435.835 -32.725 ;
        RECT 437.845 -33.340 438.075 -32.725 ;
        RECT 443.390 -33.340 443.735 -32.590 ;
        RECT 445.250 -33.340 445.590 -32.565 ;
        RECT 450.510 -33.340 450.850 -32.725 ;
        RECT 456.150 -33.340 456.380 -32.510 ;
        RECT 459.395 -33.340 459.735 -32.765 ;
        RECT 461.530 -33.340 461.870 -32.450 ;
        RECT 165.900 -34.355 166.130 -33.805 ;
        RECT 190.580 -34.355 190.810 -33.805 ;
        RECT 295.920 -33.940 463.040 -33.340 ;
        RECT 296.290 -34.830 296.630 -33.940 ;
        RECT 297.285 -34.735 297.515 -33.940 ;
        RECT 301.710 -34.690 302.055 -33.940 ;
        RECT 303.570 -34.715 303.910 -33.940 ;
        RECT 308.830 -34.555 309.170 -33.940 ;
        RECT 314.470 -34.770 314.700 -33.940 ;
        RECT 317.715 -34.515 318.055 -33.940 ;
        RECT 320.065 -34.405 320.295 -33.940 ;
        RECT 323.445 -34.405 323.675 -33.940 ;
        RECT 326.405 -34.735 326.635 -33.940 ;
        RECT 331.790 -34.565 332.130 -33.940 ;
        RECT 335.510 -34.825 335.850 -33.940 ;
        RECT 336.885 -34.730 337.115 -33.940 ;
        RECT 339.125 -34.585 339.355 -33.940 ;
        RECT 339.845 -34.725 340.075 -33.940 ;
        RECT 342.085 -34.725 342.315 -33.940 ;
        RECT 344.490 -34.690 344.830 -33.940 ;
        RECT 346.730 -34.735 347.070 -33.940 ;
        RECT 348.805 -34.680 349.035 -33.940 ;
        RECT 354.750 -34.275 355.090 -33.940 ;
        RECT 360.350 -34.275 360.690 -33.940 ;
        RECT 363.765 -34.680 363.995 -33.940 ;
        RECT 365.950 -34.565 366.290 -33.940 ;
        RECT 368.910 -34.565 369.250 -33.940 ;
        RECT 372.670 -34.565 373.010 -33.940 ;
        RECT 374.710 -34.825 375.050 -33.940 ;
        RECT 375.685 -34.735 375.915 -33.940 ;
        RECT 382.530 -34.735 382.870 -33.940 ;
        RECT 384.770 -34.690 385.110 -33.940 ;
        RECT 386.165 -34.730 386.395 -33.940 ;
        RECT 388.405 -34.585 388.635 -33.940 ;
        RECT 390.590 -34.565 390.930 -33.940 ;
        RECT 392.485 -34.685 392.715 -33.940 ;
        RECT 394.725 -34.685 394.955 -33.940 ;
        RECT 396.965 -34.685 397.195 -33.940 ;
        RECT 399.205 -34.685 399.435 -33.940 ;
        RECT 401.445 -34.685 401.675 -33.940 ;
        RECT 403.685 -34.685 403.915 -33.940 ;
        RECT 405.925 -34.685 406.155 -33.940 ;
        RECT 408.165 -34.685 408.395 -33.940 ;
        RECT 410.405 -34.735 410.635 -33.940 ;
        RECT 413.910 -34.825 414.250 -33.940 ;
        RECT 414.885 -34.735 415.115 -33.940 ;
        RECT 419.925 -34.710 420.155 -33.940 ;
        RECT 422.165 -34.710 422.395 -33.940 ;
        RECT 424.405 -34.710 424.635 -33.940 ;
        RECT 426.645 -34.710 426.875 -33.940 ;
        RECT 431.520 -34.275 431.880 -33.940 ;
        RECT 435.800 -34.275 436.160 -33.940 ;
        RECT 445.525 -34.680 445.755 -33.940 ;
        RECT 447.585 -34.505 447.815 -33.940 ;
        RECT 450.905 -34.505 451.135 -33.940 ;
        RECT 453.110 -34.825 453.450 -33.940 ;
        RECT 457.050 -34.690 457.390 -33.940 ;
        RECT 459.290 -34.735 459.630 -33.940 ;
        RECT 461.530 -34.830 461.870 -33.940 ;
        RECT 296.290 -41.180 296.630 -40.290 ;
        RECT 297.630 -41.180 297.970 -40.715 ;
        RECT 299.870 -41.180 300.210 -40.715 ;
        RECT 302.110 -41.180 302.450 -40.715 ;
        RECT 304.350 -41.180 304.690 -40.715 ;
        RECT 306.590 -41.180 306.930 -40.715 ;
        RECT 308.830 -41.180 309.170 -40.715 ;
        RECT 311.070 -41.180 311.410 -40.715 ;
        RECT 313.365 -41.180 313.595 -40.440 ;
        RECT 315.910 -41.180 316.250 -40.295 ;
        RECT 318.670 -41.180 318.900 -40.630 ;
        RECT 321.150 -41.180 321.380 -40.655 ;
        RECT 327.310 -41.180 327.650 -40.555 ;
        RECT 330.270 -41.180 330.615 -40.430 ;
        RECT 332.130 -41.180 332.470 -40.405 ;
        RECT 337.390 -41.180 337.730 -40.565 ;
        RECT 343.030 -41.180 343.260 -40.350 ;
        RECT 346.275 -41.180 346.615 -40.605 ;
        RECT 348.245 -41.180 348.475 -40.395 ;
        RECT 350.485 -41.180 350.715 -40.395 ;
        RECT 352.725 -41.180 352.955 -40.385 ;
        RECT 355.110 -41.180 355.450 -40.295 ;
        RECT 356.085 -41.180 356.315 -40.440 ;
        RECT 358.325 -41.180 358.555 -40.410 ;
        RECT 360.565 -41.180 360.795 -40.410 ;
        RECT 362.805 -41.180 363.035 -40.410 ;
        RECT 365.045 -41.180 365.275 -40.410 ;
        RECT 367.285 -41.180 367.515 -40.385 ;
        RECT 370.590 -41.180 370.935 -40.430 ;
        RECT 372.450 -41.180 372.790 -40.405 ;
        RECT 377.710 -41.180 378.050 -40.565 ;
        RECT 383.350 -41.180 383.580 -40.350 ;
        RECT 386.595 -41.180 386.935 -40.605 ;
        RECT 388.565 -41.180 388.795 -40.385 ;
        RECT 391.925 -41.180 392.155 -40.385 ;
        RECT 394.310 -41.180 394.650 -40.295 ;
        RECT 395.285 -41.180 395.515 -40.395 ;
        RECT 397.525 -41.180 397.755 -40.395 ;
        RECT 400.830 -41.180 401.175 -40.430 ;
        RECT 402.690 -41.180 403.030 -40.405 ;
        RECT 407.950 -41.180 408.290 -40.565 ;
        RECT 413.590 -41.180 413.820 -40.350 ;
        RECT 416.835 -41.180 417.175 -40.605 ;
        RECT 419.150 -41.180 419.490 -40.715 ;
        RECT 421.390 -41.180 421.730 -40.715 ;
        RECT 423.630 -41.180 423.970 -40.715 ;
        RECT 425.870 -41.180 426.210 -40.715 ;
        RECT 428.110 -41.180 428.450 -40.715 ;
        RECT 430.350 -41.180 430.690 -40.715 ;
        RECT 432.590 -41.180 432.930 -40.715 ;
        RECT 433.510 -41.180 433.850 -40.295 ;
        RECT 435.045 -41.180 435.275 -40.535 ;
        RECT 437.285 -41.180 437.515 -40.390 ;
        RECT 439.925 -41.180 440.155 -40.440 ;
        RECT 442.270 -41.180 442.610 -40.715 ;
        RECT 444.510 -41.180 444.850 -40.715 ;
        RECT 446.750 -41.180 447.090 -40.715 ;
        RECT 448.990 -41.180 449.330 -40.715 ;
        RECT 451.230 -41.180 451.570 -40.715 ;
        RECT 453.470 -41.180 453.810 -40.715 ;
        RECT 455.710 -41.180 456.050 -40.715 ;
        RECT 457.040 -41.180 457.380 -40.715 ;
        RECT 459.375 -41.180 459.715 -40.715 ;
        RECT 461.530 -41.180 461.870 -40.290 ;
        RECT 295.920 -41.780 463.040 -41.180 ;
        RECT 296.290 -42.670 296.630 -41.780 ;
        RECT 297.630 -42.245 297.970 -41.780 ;
        RECT 299.870 -42.245 300.210 -41.780 ;
        RECT 302.110 -42.245 302.450 -41.780 ;
        RECT 304.350 -42.245 304.690 -41.780 ;
        RECT 306.590 -42.245 306.930 -41.780 ;
        RECT 308.830 -42.245 309.170 -41.780 ;
        RECT 311.070 -42.245 311.410 -41.780 ;
        RECT 312.010 -42.530 312.350 -41.780 ;
        RECT 314.250 -42.575 314.590 -41.780 ;
        RECT 317.390 -42.530 317.735 -41.780 ;
        RECT 319.250 -42.555 319.590 -41.780 ;
        RECT 324.510 -42.395 324.850 -41.780 ;
        RECT 330.150 -42.610 330.380 -41.780 ;
        RECT 333.395 -42.355 333.735 -41.780 ;
        RECT 335.510 -42.665 335.850 -41.780 ;
        RECT 337.770 -42.530 338.110 -41.780 ;
        RECT 340.010 -42.575 340.350 -41.780 ;
        RECT 342.085 -42.245 342.315 -41.780 ;
        RECT 345.465 -42.245 345.695 -41.780 ;
        RECT 347.790 -42.330 348.020 -41.780 ;
        RECT 350.270 -42.305 350.500 -41.780 ;
        RECT 351.045 -42.575 351.275 -41.780 ;
        RECT 356.105 -42.355 356.445 -41.780 ;
        RECT 359.460 -42.610 359.690 -41.780 ;
        RECT 364.990 -42.395 365.330 -41.780 ;
        RECT 370.250 -42.555 370.590 -41.780 ;
        RECT 372.105 -42.530 372.450 -41.780 ;
        RECT 374.710 -42.665 375.050 -41.780 ;
        RECT 377.205 -42.520 377.435 -41.780 ;
        RECT 380.110 -42.405 380.450 -41.780 ;
        RECT 383.545 -42.355 383.885 -41.780 ;
        RECT 386.900 -42.610 387.130 -41.780 ;
        RECT 392.430 -42.395 392.770 -41.780 ;
        RECT 397.690 -42.555 398.030 -41.780 ;
        RECT 399.545 -42.530 399.890 -41.780 ;
        RECT 403.685 -42.575 403.915 -41.780 ;
        RECT 405.925 -42.520 406.155 -41.780 ;
        RECT 410.405 -42.575 410.635 -41.780 ;
        RECT 413.910 -42.665 414.250 -41.780 ;
        RECT 414.885 -42.575 415.115 -41.780 ;
        RECT 418.245 -42.520 418.475 -41.780 ;
        RECT 421.550 -42.530 421.895 -41.780 ;
        RECT 423.410 -42.555 423.750 -41.780 ;
        RECT 428.670 -42.395 429.010 -41.780 ;
        RECT 434.310 -42.610 434.540 -41.780 ;
        RECT 437.555 -42.355 437.895 -41.780 ;
        RECT 440.645 -42.520 440.875 -41.780 ;
        RECT 445.125 -42.565 445.355 -41.780 ;
        RECT 447.365 -42.565 447.595 -41.780 ;
        RECT 453.110 -42.665 453.450 -41.780 ;
        RECT 455.605 -42.640 455.835 -41.780 ;
        RECT 459.470 -42.405 459.810 -41.780 ;
        RECT 461.530 -42.670 461.870 -41.780 ;
        RECT 296.290 -49.020 296.630 -48.130 ;
        RECT 299.310 -49.020 299.650 -48.555 ;
        RECT 301.550 -49.020 301.890 -48.555 ;
        RECT 303.790 -49.020 304.130 -48.555 ;
        RECT 306.030 -49.020 306.370 -48.555 ;
        RECT 308.270 -49.020 308.610 -48.555 ;
        RECT 310.510 -49.020 310.850 -48.555 ;
        RECT 312.750 -49.020 313.090 -48.555 ;
        RECT 315.350 -49.020 315.690 -48.135 ;
        RECT 316.830 -49.020 317.170 -48.555 ;
        RECT 319.070 -49.020 319.410 -48.555 ;
        RECT 321.310 -49.020 321.650 -48.555 ;
        RECT 323.550 -49.020 323.890 -48.555 ;
        RECT 325.790 -49.020 326.130 -48.555 ;
        RECT 328.030 -49.020 328.370 -48.555 ;
        RECT 330.270 -49.020 330.610 -48.555 ;
        RECT 334.390 -49.020 334.730 -48.135 ;
        RECT 335.310 -49.020 335.650 -48.555 ;
        RECT 337.550 -49.020 337.890 -48.555 ;
        RECT 339.790 -49.020 340.130 -48.555 ;
        RECT 342.030 -49.020 342.370 -48.555 ;
        RECT 344.270 -49.020 344.610 -48.555 ;
        RECT 346.510 -49.020 346.850 -48.555 ;
        RECT 348.750 -49.020 349.090 -48.555 ;
        RECT 349.925 -49.020 350.155 -48.225 ;
        RECT 353.430 -49.020 353.770 -48.135 ;
        RECT 354.350 -49.020 354.690 -48.555 ;
        RECT 356.590 -49.020 356.930 -48.555 ;
        RECT 358.830 -49.020 359.170 -48.555 ;
        RECT 361.070 -49.020 361.410 -48.555 ;
        RECT 363.310 -49.020 363.650 -48.555 ;
        RECT 365.550 -49.020 365.890 -48.555 ;
        RECT 367.790 -49.020 368.130 -48.555 ;
        RECT 368.965 -49.020 369.195 -48.225 ;
        RECT 372.470 -49.020 372.810 -48.135 ;
        RECT 373.390 -49.020 373.730 -48.555 ;
        RECT 375.630 -49.020 375.970 -48.555 ;
        RECT 377.870 -49.020 378.210 -48.555 ;
        RECT 380.110 -49.020 380.450 -48.555 ;
        RECT 382.350 -49.020 382.690 -48.555 ;
        RECT 384.590 -49.020 384.930 -48.555 ;
        RECT 386.830 -49.020 387.170 -48.555 ;
        RECT 388.565 -49.020 388.795 -48.280 ;
        RECT 391.510 -49.020 391.850 -48.135 ;
        RECT 392.430 -49.020 392.770 -48.555 ;
        RECT 394.670 -49.020 395.010 -48.555 ;
        RECT 396.910 -49.020 397.250 -48.555 ;
        RECT 399.150 -49.020 399.490 -48.555 ;
        RECT 401.390 -49.020 401.730 -48.555 ;
        RECT 403.630 -49.020 403.970 -48.555 ;
        RECT 405.870 -49.020 406.210 -48.555 ;
        RECT 407.045 -49.020 407.275 -48.225 ;
        RECT 410.550 -49.020 410.890 -48.135 ;
        RECT 411.470 -49.020 411.810 -48.555 ;
        RECT 413.710 -49.020 414.050 -48.555 ;
        RECT 415.950 -49.020 416.290 -48.555 ;
        RECT 418.190 -49.020 418.530 -48.555 ;
        RECT 420.430 -49.020 420.770 -48.555 ;
        RECT 422.670 -49.020 423.010 -48.555 ;
        RECT 424.910 -49.020 425.250 -48.555 ;
        RECT 426.085 -49.020 426.315 -48.225 ;
        RECT 429.590 -49.020 429.930 -48.135 ;
        RECT 430.510 -49.020 430.850 -48.555 ;
        RECT 432.750 -49.020 433.090 -48.555 ;
        RECT 434.990 -49.020 435.330 -48.555 ;
        RECT 437.230 -49.020 437.570 -48.555 ;
        RECT 439.470 -49.020 439.810 -48.555 ;
        RECT 441.710 -49.020 442.050 -48.555 ;
        RECT 443.950 -49.020 444.290 -48.555 ;
        RECT 445.125 -49.020 445.355 -48.225 ;
        RECT 448.630 -49.020 448.970 -48.135 ;
        RECT 455.710 -49.020 456.050 -48.395 ;
        RECT 459.470 -49.020 459.810 -48.395 ;
        RECT 461.530 -49.020 461.870 -48.130 ;
        RECT 295.920 -49.620 463.040 -49.020 ;
        RECT 146.665 -60.040 147.825 -59.670 ;
        RECT 145.775 -60.380 147.825 -60.040 ;
        RECT 146.665 -62.715 147.825 -60.380 ;
        RECT 146.015 -62.945 147.825 -62.715 ;
        RECT 146.665 -64.985 147.825 -62.945 ;
        RECT 146.015 -65.215 147.825 -64.985 ;
        RECT 146.665 -66.075 147.825 -65.215 ;
        RECT 146.015 -66.305 147.825 -66.075 ;
        RECT 146.665 -68.345 147.825 -66.305 ;
        RECT 146.015 -68.575 147.825 -68.345 ;
        RECT 146.665 -69.435 147.825 -68.575 ;
        RECT 146.015 -69.665 147.825 -69.435 ;
        RECT 146.665 -71.705 147.825 -69.665 ;
        RECT 146.015 -71.935 147.825 -71.705 ;
        RECT 146.665 -72.795 147.825 -71.935 ;
        RECT 146.015 -73.025 147.825 -72.795 ;
        RECT 146.665 -75.065 147.825 -73.025 ;
        RECT 146.015 -75.295 147.825 -75.065 ;
        RECT 146.665 -76.155 147.825 -75.295 ;
        RECT 146.015 -76.385 147.825 -76.155 ;
        RECT 146.665 -78.425 147.825 -76.385 ;
        RECT 146.015 -78.655 147.825 -78.425 ;
        RECT 146.665 -79.515 147.825 -78.655 ;
        RECT 146.015 -79.745 147.825 -79.515 ;
        RECT 146.665 -81.785 147.825 -79.745 ;
        RECT 146.015 -82.015 147.825 -81.785 ;
        RECT 146.665 -82.875 147.825 -82.015 ;
        RECT 146.015 -83.105 147.825 -82.875 ;
        RECT -496.745 -84.700 -492.560 -84.470 ;
        RECT -496.745 -85.370 -496.365 -84.700 ;
        RECT -495.350 -87.115 -495.120 -84.700 ;
        RECT 146.665 -85.145 147.825 -83.105 ;
        RECT 146.015 -85.375 147.825 -85.145 ;
        RECT 146.665 -86.235 147.825 -85.375 ;
        RECT 146.015 -86.465 147.825 -86.235 ;
        RECT 146.665 -88.505 147.825 -86.465 ;
        RECT 146.015 -88.735 147.825 -88.505 ;
        RECT 146.665 -89.595 147.825 -88.735 ;
        RECT 146.015 -89.825 147.825 -89.595 ;
        RECT 146.665 -91.865 147.825 -89.825 ;
        RECT 146.015 -92.095 147.825 -91.865 ;
        RECT 146.665 -92.955 147.825 -92.095 ;
        RECT 146.015 -93.185 147.825 -92.955 ;
        RECT -494.375 -95.665 -494.145 -95.115 ;
        RECT 146.665 -95.225 147.825 -93.185 ;
        RECT 146.015 -95.455 147.825 -95.225 ;
        RECT -494.525 -96.400 -494.145 -95.665 ;
        RECT 146.665 -96.315 147.825 -95.455 ;
        RECT -494.525 -96.565 -492.575 -96.400 ;
        RECT 146.015 -96.545 147.825 -96.315 ;
        RECT -494.375 -96.630 -492.575 -96.565 ;
        RECT -494.375 -97.115 -494.145 -96.630 ;
        RECT 146.665 -98.585 147.825 -96.545 ;
        RECT 146.015 -98.815 147.825 -98.585 ;
        RECT 146.665 -101.520 147.825 -98.815 ;
        RECT 145.775 -101.860 147.825 -101.520 ;
        RECT 146.665 -127.660 147.825 -101.860 ;
        RECT 146.625 -132.620 147.865 -127.660 ;
      LAYER Via1 ;
        RECT 146.805 132.180 147.065 132.440 ;
        RECT 147.425 132.180 147.685 132.440 ;
        RECT 146.805 131.560 147.065 131.820 ;
        RECT 147.425 131.560 147.685 131.820 ;
        RECT 146.805 130.940 147.065 131.200 ;
        RECT 147.425 130.940 147.685 131.200 ;
        RECT 146.805 130.320 147.065 130.580 ;
        RECT 147.425 130.320 147.685 130.580 ;
        RECT 146.805 129.700 147.065 129.960 ;
        RECT 147.425 129.700 147.685 129.960 ;
        RECT 146.805 129.080 147.065 129.340 ;
        RECT 147.425 129.080 147.685 129.340 ;
        RECT 146.805 128.460 147.065 128.720 ;
        RECT 147.425 128.460 147.685 128.720 ;
        RECT 146.805 127.840 147.065 128.100 ;
        RECT 147.425 127.840 147.685 128.100 ;
        RECT -494.465 95.725 -494.205 96.505 ;
        RECT -496.685 84.530 -496.425 85.310 ;
        RECT 336.850 44.630 338.150 44.890 ;
        RECT 378.430 44.630 379.730 44.890 ;
        RECT 420.010 44.630 421.310 44.890 ;
        RECT 461.590 44.630 462.890 44.890 ;
        RECT 336.850 36.790 338.150 37.050 ;
        RECT 378.430 36.790 379.730 37.050 ;
        RECT 420.010 36.790 421.310 37.050 ;
        RECT 461.590 36.790 462.890 37.050 ;
        RECT 165.885 32.965 166.145 33.745 ;
        RECT 190.565 32.965 190.825 33.745 ;
        RECT 167.375 31.715 167.635 32.495 ;
        RECT 168.975 31.715 169.235 32.495 ;
        RECT 174.175 31.715 174.435 32.495 ;
        RECT 179.175 31.715 179.435 32.495 ;
        RECT 183.475 31.715 183.735 32.495 ;
        RECT 185.075 31.715 185.335 32.495 ;
        RECT 186.675 31.715 186.935 32.495 ;
        RECT 188.275 31.715 188.535 32.495 ;
        RECT 189.875 31.715 190.135 32.495 ;
        RECT 336.850 28.950 338.150 29.210 ;
        RECT 378.430 28.950 379.730 29.210 ;
        RECT 420.010 28.950 421.310 29.210 ;
        RECT 461.590 28.950 462.890 29.210 ;
        RECT 336.850 21.110 338.150 21.370 ;
        RECT 378.430 21.110 379.730 21.370 ;
        RECT 420.010 21.110 421.310 21.370 ;
        RECT 461.590 21.110 462.890 21.370 ;
        RECT 336.850 13.270 338.150 13.530 ;
        RECT 378.430 13.270 379.730 13.530 ;
        RECT 420.010 13.270 421.310 13.530 ;
        RECT 461.590 13.270 462.890 13.530 ;
        RECT 229.270 9.780 229.530 10.560 ;
        RECT 229.270 5.420 229.530 6.200 ;
        RECT 336.850 5.430 338.150 5.690 ;
        RECT 378.430 5.430 379.730 5.690 ;
        RECT 420.010 5.430 421.310 5.690 ;
        RECT 461.590 5.430 462.890 5.690 ;
        RECT 229.270 3.240 229.530 4.020 ;
        RECT 183.475 1.445 183.735 2.225 ;
        RECT 185.965 1.370 186.745 1.630 ;
        RECT 229.270 -1.120 229.530 -0.340 ;
        RECT 183.475 -2.225 183.735 -1.445 ;
        RECT 185.965 -1.630 186.745 -1.370 ;
        RECT 336.850 -2.410 338.150 -2.150 ;
        RECT 378.430 -2.410 379.730 -2.150 ;
        RECT 420.010 -2.410 421.310 -2.150 ;
        RECT 461.590 -2.410 462.890 -2.150 ;
        RECT 336.850 -10.250 338.150 -9.990 ;
        RECT 378.430 -10.250 379.730 -9.990 ;
        RECT 420.010 -10.250 421.310 -9.990 ;
        RECT 461.590 -10.250 462.890 -9.990 ;
        RECT 230.550 -12.455 231.330 -12.195 ;
        RECT 234.065 -12.455 234.845 -12.195 ;
        RECT 336.850 -18.090 338.150 -17.830 ;
        RECT 378.430 -18.090 379.730 -17.830 ;
        RECT 420.010 -18.090 421.310 -17.830 ;
        RECT 461.590 -18.090 462.890 -17.830 ;
        RECT 336.850 -25.930 338.150 -25.670 ;
        RECT 378.430 -25.930 379.730 -25.670 ;
        RECT 420.010 -25.930 421.310 -25.670 ;
        RECT 461.590 -25.930 462.890 -25.670 ;
        RECT 167.375 -32.495 167.635 -31.715 ;
        RECT 168.975 -32.495 169.235 -31.715 ;
        RECT 174.175 -32.495 174.435 -31.715 ;
        RECT 179.175 -32.495 179.435 -31.715 ;
        RECT 183.475 -32.495 183.735 -31.715 ;
        RECT 185.075 -32.495 185.335 -31.715 ;
        RECT 186.675 -32.495 186.935 -31.715 ;
        RECT 188.275 -32.495 188.535 -31.715 ;
        RECT 189.875 -32.495 190.135 -31.715 ;
        RECT 165.885 -33.745 166.145 -32.965 ;
        RECT 190.565 -33.745 190.825 -32.965 ;
        RECT 336.850 -33.770 338.150 -33.510 ;
        RECT 378.430 -33.770 379.730 -33.510 ;
        RECT 420.010 -33.770 421.310 -33.510 ;
        RECT 461.590 -33.770 462.890 -33.510 ;
        RECT 336.850 -41.610 338.150 -41.350 ;
        RECT 378.430 -41.610 379.730 -41.350 ;
        RECT 420.010 -41.610 421.310 -41.350 ;
        RECT 461.590 -41.610 462.890 -41.350 ;
        RECT 336.850 -49.450 338.150 -49.190 ;
        RECT 378.430 -49.450 379.730 -49.190 ;
        RECT 420.010 -49.450 421.310 -49.190 ;
        RECT 461.590 -49.450 462.890 -49.190 ;
        RECT -496.685 -85.310 -496.425 -84.530 ;
        RECT -494.465 -96.505 -494.205 -95.725 ;
        RECT 146.805 -128.100 147.065 -127.840 ;
        RECT 147.425 -128.100 147.685 -127.840 ;
        RECT 146.805 -128.720 147.065 -128.460 ;
        RECT 147.425 -128.720 147.685 -128.460 ;
        RECT 146.805 -129.340 147.065 -129.080 ;
        RECT 147.425 -129.340 147.685 -129.080 ;
        RECT 146.805 -129.960 147.065 -129.700 ;
        RECT 147.425 -129.960 147.685 -129.700 ;
        RECT 146.805 -130.580 147.065 -130.320 ;
        RECT 147.425 -130.580 147.685 -130.320 ;
        RECT 146.805 -131.200 147.065 -130.940 ;
        RECT 147.425 -131.200 147.685 -130.940 ;
        RECT 146.805 -131.820 147.065 -131.560 ;
        RECT 147.425 -131.820 147.685 -131.560 ;
        RECT 146.805 -132.440 147.065 -132.180 ;
        RECT 147.425 -132.440 147.685 -132.180 ;
      LAYER Metal2 ;
        RECT -499.655 127.660 -493.455 132.620 ;
        RECT 146.625 127.660 147.865 132.620 ;
        RECT -496.745 96.315 -496.365 127.660 ;
        RECT -494.525 96.315 -494.145 97.615 ;
        RECT -496.745 95.915 -494.145 96.315 ;
        RECT -496.745 84.470 -496.365 95.915 ;
        RECT -494.525 94.615 -494.145 95.915 ;
        RECT 336.840 44.570 338.160 44.950 ;
        RECT 378.420 44.570 379.740 44.950 ;
        RECT 420.000 44.570 421.320 44.950 ;
        RECT 461.580 44.570 462.900 44.950 ;
        RECT 336.840 36.730 338.160 37.110 ;
        RECT 378.420 36.730 379.740 37.110 ;
        RECT 420.000 36.730 421.320 37.110 ;
        RECT 461.580 36.730 462.900 37.110 ;
        RECT 165.825 33.355 166.215 33.805 ;
        RECT 165.815 32.325 166.215 33.355 ;
        RECT 190.495 33.355 190.885 33.805 ;
        RECT 167.315 32.325 167.695 32.555 ;
        RECT 168.915 32.325 169.295 32.555 ;
        RECT 174.115 32.325 174.495 32.555 ;
        RECT 179.115 32.325 179.495 32.555 ;
        RECT 183.415 32.325 183.795 32.555 ;
        RECT 185.015 32.325 185.395 32.555 ;
        RECT 186.615 32.325 186.995 32.555 ;
        RECT 188.215 32.325 188.595 32.555 ;
        RECT 189.815 32.325 190.195 32.555 ;
        RECT 190.495 32.325 190.895 33.355 ;
        RECT 194.795 32.325 195.915 32.635 ;
        RECT 165.815 31.925 195.915 32.325 ;
        RECT 165.825 22.350 166.215 31.925 ;
        RECT 167.315 31.655 167.695 31.925 ;
        RECT 168.915 31.655 169.295 31.925 ;
        RECT 174.115 31.655 174.495 31.925 ;
        RECT 179.115 31.655 179.495 31.925 ;
        RECT 183.415 31.655 183.795 31.925 ;
        RECT 185.015 31.655 185.395 31.925 ;
        RECT 186.615 31.655 186.995 31.925 ;
        RECT 188.215 31.655 188.595 31.925 ;
        RECT 189.815 31.655 190.195 31.925 ;
        RECT 190.495 22.350 190.885 31.925 ;
        RECT 194.795 31.615 195.915 31.925 ;
        RECT 336.840 28.890 338.160 29.270 ;
        RECT 378.420 28.890 379.740 29.270 ;
        RECT 420.000 28.890 421.320 29.270 ;
        RECT 461.580 28.890 462.900 29.270 ;
        RECT 165.825 21.950 170.020 22.350 ;
        RECT 169.620 21.240 170.020 21.950 ;
        RECT 188.660 21.950 190.885 22.350 ;
        RECT 188.660 21.240 189.060 21.950 ;
        RECT 169.680 11.625 169.960 21.240 ;
        RECT 188.720 11.625 189.000 21.240 ;
        RECT 336.840 21.050 338.160 21.430 ;
        RECT 378.420 21.050 379.740 21.430 ;
        RECT 420.000 21.050 421.320 21.430 ;
        RECT 461.580 21.050 462.900 21.430 ;
        RECT 336.840 13.210 338.160 13.590 ;
        RECT 378.420 13.210 379.740 13.590 ;
        RECT 420.000 13.210 421.320 13.590 ;
        RECT 461.580 13.210 462.900 13.590 ;
        RECT 229.210 9.220 229.590 11.670 ;
        RECT 183.415 1.690 183.795 2.285 ;
        RECT 183.415 1.310 187.785 1.690 ;
        RECT 187.405 0.220 187.785 1.310 ;
        RECT 194.795 0.220 195.915 0.510 ;
        RECT 227.990 0.220 229.590 9.220 ;
        RECT 336.840 5.370 338.160 5.750 ;
        RECT 378.420 5.370 379.740 5.750 ;
        RECT 420.000 5.370 421.320 5.750 ;
        RECT 461.580 5.370 462.900 5.750 ;
        RECT 187.405 -0.220 195.915 0.220 ;
        RECT 187.405 -1.310 187.785 -0.220 ;
        RECT 194.795 -0.510 195.915 -0.220 ;
        RECT 183.415 -1.690 187.785 -1.310 ;
        RECT 183.415 -2.285 183.795 -1.690 ;
        RECT 229.210 -2.230 229.590 0.220 ;
        RECT 336.840 -2.470 338.160 -2.090 ;
        RECT 378.420 -2.470 379.740 -2.090 ;
        RECT 420.000 -2.470 421.320 -2.090 ;
        RECT 461.580 -2.470 462.900 -2.090 ;
        RECT 336.840 -10.310 338.160 -9.930 ;
        RECT 378.420 -10.310 379.740 -9.930 ;
        RECT 420.000 -10.310 421.320 -9.930 ;
        RECT 461.580 -10.310 462.900 -9.930 ;
        RECT 169.680 -21.240 169.960 -11.625 ;
        RECT 188.720 -21.240 189.000 -11.625 ;
        RECT 229.440 -12.515 235.960 -12.135 ;
        RECT 229.700 -13.735 235.700 -12.515 ;
        RECT 336.840 -18.150 338.160 -17.770 ;
        RECT 378.420 -18.150 379.740 -17.770 ;
        RECT 420.000 -18.150 421.320 -17.770 ;
        RECT 461.580 -18.150 462.900 -17.770 ;
        RECT 169.620 -21.950 170.020 -21.240 ;
        RECT 165.825 -22.350 170.020 -21.950 ;
        RECT 188.660 -21.950 189.060 -21.240 ;
        RECT 188.660 -22.350 190.885 -21.950 ;
        RECT 165.825 -31.925 166.215 -22.350 ;
        RECT 167.315 -31.925 167.695 -31.655 ;
        RECT 168.915 -31.925 169.295 -31.655 ;
        RECT 174.115 -31.925 174.495 -31.655 ;
        RECT 179.115 -31.925 179.495 -31.655 ;
        RECT 183.415 -31.925 183.795 -31.655 ;
        RECT 185.015 -31.925 185.395 -31.655 ;
        RECT 186.615 -31.925 186.995 -31.655 ;
        RECT 188.215 -31.925 188.595 -31.655 ;
        RECT 189.815 -31.925 190.195 -31.655 ;
        RECT 190.495 -31.925 190.885 -22.350 ;
        RECT 336.840 -25.990 338.160 -25.610 ;
        RECT 378.420 -25.990 379.740 -25.610 ;
        RECT 420.000 -25.990 421.320 -25.610 ;
        RECT 461.580 -25.990 462.900 -25.610 ;
        RECT 194.795 -31.925 195.915 -31.615 ;
        RECT 165.815 -32.325 195.915 -31.925 ;
        RECT 165.815 -33.355 166.215 -32.325 ;
        RECT 167.315 -32.555 167.695 -32.325 ;
        RECT 168.915 -32.555 169.295 -32.325 ;
        RECT 174.115 -32.555 174.495 -32.325 ;
        RECT 179.115 -32.555 179.495 -32.325 ;
        RECT 183.415 -32.555 183.795 -32.325 ;
        RECT 185.015 -32.555 185.395 -32.325 ;
        RECT 186.615 -32.555 186.995 -32.325 ;
        RECT 188.215 -32.555 188.595 -32.325 ;
        RECT 189.815 -32.555 190.195 -32.325 ;
        RECT 165.825 -33.805 166.215 -33.355 ;
        RECT 190.495 -33.355 190.895 -32.325 ;
        RECT 194.795 -32.635 195.915 -32.325 ;
        RECT 190.495 -33.805 190.885 -33.355 ;
        RECT 336.840 -33.830 338.160 -33.450 ;
        RECT 378.420 -33.830 379.740 -33.450 ;
        RECT 420.000 -33.830 421.320 -33.450 ;
        RECT 461.580 -33.830 462.900 -33.450 ;
        RECT 336.840 -41.670 338.160 -41.290 ;
        RECT 378.420 -41.670 379.740 -41.290 ;
        RECT 420.000 -41.670 421.320 -41.290 ;
        RECT 461.580 -41.670 462.900 -41.290 ;
        RECT 336.840 -49.510 338.160 -49.130 ;
        RECT 378.420 -49.510 379.740 -49.130 ;
        RECT 420.000 -49.510 421.320 -49.130 ;
        RECT 461.580 -49.510 462.900 -49.130 ;
        RECT -496.745 -95.915 -496.365 -84.470 ;
        RECT -494.525 -95.915 -494.145 -94.615 ;
        RECT -496.745 -96.315 -494.145 -95.915 ;
        RECT -496.745 -127.660 -496.365 -96.315 ;
        RECT -494.525 -97.615 -494.145 -96.315 ;
        RECT -499.655 -132.620 -493.455 -127.660 ;
        RECT 146.625 -132.620 147.865 -127.660 ;
      LAYER Via2 ;
        RECT -499.485 132.170 -499.205 132.450 ;
        RECT -498.865 132.170 -498.585 132.450 ;
        RECT -498.245 132.170 -497.965 132.450 ;
        RECT -497.625 132.170 -497.345 132.450 ;
        RECT -497.005 132.170 -496.725 132.450 ;
        RECT -496.385 132.170 -496.105 132.450 ;
        RECT -495.765 132.170 -495.485 132.450 ;
        RECT -495.145 132.170 -494.865 132.450 ;
        RECT -494.525 132.170 -494.245 132.450 ;
        RECT -493.905 132.170 -493.625 132.450 ;
        RECT -499.485 131.550 -499.205 131.830 ;
        RECT -498.865 131.550 -498.585 131.830 ;
        RECT -498.245 131.550 -497.965 131.830 ;
        RECT -497.625 131.550 -497.345 131.830 ;
        RECT -497.005 131.550 -496.725 131.830 ;
        RECT -496.385 131.550 -496.105 131.830 ;
        RECT -495.765 131.550 -495.485 131.830 ;
        RECT -495.145 131.550 -494.865 131.830 ;
        RECT -494.525 131.550 -494.245 131.830 ;
        RECT -493.905 131.550 -493.625 131.830 ;
        RECT -499.485 130.930 -499.205 131.210 ;
        RECT -498.865 130.930 -498.585 131.210 ;
        RECT -498.245 130.930 -497.965 131.210 ;
        RECT -497.625 130.930 -497.345 131.210 ;
        RECT -497.005 130.930 -496.725 131.210 ;
        RECT -496.385 130.930 -496.105 131.210 ;
        RECT -495.765 130.930 -495.485 131.210 ;
        RECT -495.145 130.930 -494.865 131.210 ;
        RECT -494.525 130.930 -494.245 131.210 ;
        RECT -493.905 130.930 -493.625 131.210 ;
        RECT -499.485 130.310 -499.205 130.590 ;
        RECT -498.865 130.310 -498.585 130.590 ;
        RECT -498.245 130.310 -497.965 130.590 ;
        RECT -497.625 130.310 -497.345 130.590 ;
        RECT -497.005 130.310 -496.725 130.590 ;
        RECT -496.385 130.310 -496.105 130.590 ;
        RECT -495.765 130.310 -495.485 130.590 ;
        RECT -495.145 130.310 -494.865 130.590 ;
        RECT -494.525 130.310 -494.245 130.590 ;
        RECT -493.905 130.310 -493.625 130.590 ;
        RECT -499.485 129.690 -499.205 129.970 ;
        RECT -498.865 129.690 -498.585 129.970 ;
        RECT -498.245 129.690 -497.965 129.970 ;
        RECT -497.625 129.690 -497.345 129.970 ;
        RECT -497.005 129.690 -496.725 129.970 ;
        RECT -496.385 129.690 -496.105 129.970 ;
        RECT -495.765 129.690 -495.485 129.970 ;
        RECT -495.145 129.690 -494.865 129.970 ;
        RECT -494.525 129.690 -494.245 129.970 ;
        RECT -493.905 129.690 -493.625 129.970 ;
        RECT -499.485 129.070 -499.205 129.350 ;
        RECT -498.865 129.070 -498.585 129.350 ;
        RECT -498.245 129.070 -497.965 129.350 ;
        RECT -497.625 129.070 -497.345 129.350 ;
        RECT -497.005 129.070 -496.725 129.350 ;
        RECT -496.385 129.070 -496.105 129.350 ;
        RECT -495.765 129.070 -495.485 129.350 ;
        RECT -495.145 129.070 -494.865 129.350 ;
        RECT -494.525 129.070 -494.245 129.350 ;
        RECT -493.905 129.070 -493.625 129.350 ;
        RECT -499.485 128.450 -499.205 128.730 ;
        RECT -498.865 128.450 -498.585 128.730 ;
        RECT -498.245 128.450 -497.965 128.730 ;
        RECT -497.625 128.450 -497.345 128.730 ;
        RECT -497.005 128.450 -496.725 128.730 ;
        RECT -496.385 128.450 -496.105 128.730 ;
        RECT -495.765 128.450 -495.485 128.730 ;
        RECT -495.145 128.450 -494.865 128.730 ;
        RECT -494.525 128.450 -494.245 128.730 ;
        RECT -493.905 128.450 -493.625 128.730 ;
        RECT -499.485 127.830 -499.205 128.110 ;
        RECT -498.865 127.830 -498.585 128.110 ;
        RECT -498.245 127.830 -497.965 128.110 ;
        RECT -497.625 127.830 -497.345 128.110 ;
        RECT -497.005 127.830 -496.725 128.110 ;
        RECT -496.385 127.830 -496.105 128.110 ;
        RECT -495.765 127.830 -495.485 128.110 ;
        RECT -495.145 127.830 -494.865 128.110 ;
        RECT -494.525 127.830 -494.245 128.110 ;
        RECT -493.905 127.830 -493.625 128.110 ;
        RECT 146.795 132.170 147.075 132.450 ;
        RECT 147.415 132.170 147.695 132.450 ;
        RECT 146.795 131.550 147.075 131.830 ;
        RECT 147.415 131.550 147.695 131.830 ;
        RECT 146.795 130.930 147.075 131.210 ;
        RECT 147.415 130.930 147.695 131.210 ;
        RECT 146.795 130.310 147.075 130.590 ;
        RECT 147.415 130.310 147.695 130.590 ;
        RECT 146.795 129.690 147.075 129.970 ;
        RECT 147.415 129.690 147.695 129.970 ;
        RECT 146.795 129.070 147.075 129.350 ;
        RECT 147.415 129.070 147.695 129.350 ;
        RECT 146.795 128.450 147.075 128.730 ;
        RECT 147.415 128.450 147.695 128.730 ;
        RECT 146.795 127.830 147.075 128.110 ;
        RECT 147.415 127.830 147.695 128.110 ;
        RECT 336.840 44.620 338.160 44.900 ;
        RECT 378.420 44.620 379.740 44.900 ;
        RECT 420.000 44.620 421.320 44.900 ;
        RECT 461.580 44.620 462.900 44.900 ;
        RECT 336.840 36.780 338.160 37.060 ;
        RECT 378.420 36.780 379.740 37.060 ;
        RECT 420.000 36.780 421.320 37.060 ;
        RECT 461.580 36.780 462.900 37.060 ;
        RECT 194.935 31.725 195.215 32.525 ;
        RECT 195.495 31.725 195.775 32.525 ;
        RECT 336.840 28.940 338.160 29.220 ;
        RECT 378.420 28.940 379.740 29.220 ;
        RECT 420.000 28.940 421.320 29.220 ;
        RECT 461.580 28.940 462.900 29.220 ;
        RECT 336.840 21.100 338.160 21.380 ;
        RECT 378.420 21.100 379.740 21.380 ;
        RECT 420.000 21.100 421.320 21.380 ;
        RECT 461.580 21.100 462.900 21.380 ;
        RECT 336.840 13.260 338.160 13.540 ;
        RECT 378.420 13.260 379.740 13.540 ;
        RECT 420.000 13.260 421.320 13.540 ;
        RECT 461.580 13.260 462.900 13.540 ;
        RECT 228.130 6.540 229.450 8.900 ;
        RECT 228.130 3.540 229.450 5.900 ;
        RECT 336.840 5.420 338.160 5.700 ;
        RECT 378.420 5.420 379.740 5.700 ;
        RECT 420.000 5.420 421.320 5.700 ;
        RECT 461.580 5.420 462.900 5.700 ;
        RECT 228.130 0.540 229.450 2.900 ;
        RECT 194.935 -0.400 195.215 0.400 ;
        RECT 195.495 -0.400 195.775 0.400 ;
        RECT 336.840 -2.420 338.160 -2.140 ;
        RECT 378.420 -2.420 379.740 -2.140 ;
        RECT 420.000 -2.420 421.320 -2.140 ;
        RECT 461.580 -2.420 462.900 -2.140 ;
        RECT 336.840 -10.260 338.160 -9.980 ;
        RECT 378.420 -10.260 379.740 -9.980 ;
        RECT 420.000 -10.260 421.320 -9.980 ;
        RECT 461.580 -10.260 462.900 -9.980 ;
        RECT 230.020 -13.595 232.380 -12.275 ;
        RECT 233.020 -13.595 235.380 -12.275 ;
        RECT 336.840 -18.100 338.160 -17.820 ;
        RECT 378.420 -18.100 379.740 -17.820 ;
        RECT 420.000 -18.100 421.320 -17.820 ;
        RECT 461.580 -18.100 462.900 -17.820 ;
        RECT 336.840 -25.940 338.160 -25.660 ;
        RECT 378.420 -25.940 379.740 -25.660 ;
        RECT 420.000 -25.940 421.320 -25.660 ;
        RECT 461.580 -25.940 462.900 -25.660 ;
        RECT 194.935 -32.525 195.215 -31.725 ;
        RECT 195.495 -32.525 195.775 -31.725 ;
        RECT 336.840 -33.780 338.160 -33.500 ;
        RECT 378.420 -33.780 379.740 -33.500 ;
        RECT 420.000 -33.780 421.320 -33.500 ;
        RECT 461.580 -33.780 462.900 -33.500 ;
        RECT 336.840 -41.620 338.160 -41.340 ;
        RECT 378.420 -41.620 379.740 -41.340 ;
        RECT 420.000 -41.620 421.320 -41.340 ;
        RECT 461.580 -41.620 462.900 -41.340 ;
        RECT 336.840 -49.460 338.160 -49.180 ;
        RECT 378.420 -49.460 379.740 -49.180 ;
        RECT 420.000 -49.460 421.320 -49.180 ;
        RECT 461.580 -49.460 462.900 -49.180 ;
        RECT -499.485 -128.110 -499.205 -127.830 ;
        RECT -498.865 -128.110 -498.585 -127.830 ;
        RECT -498.245 -128.110 -497.965 -127.830 ;
        RECT -497.625 -128.110 -497.345 -127.830 ;
        RECT -497.005 -128.110 -496.725 -127.830 ;
        RECT -496.385 -128.110 -496.105 -127.830 ;
        RECT -495.765 -128.110 -495.485 -127.830 ;
        RECT -495.145 -128.110 -494.865 -127.830 ;
        RECT -494.525 -128.110 -494.245 -127.830 ;
        RECT -493.905 -128.110 -493.625 -127.830 ;
        RECT -499.485 -128.730 -499.205 -128.450 ;
        RECT -498.865 -128.730 -498.585 -128.450 ;
        RECT -498.245 -128.730 -497.965 -128.450 ;
        RECT -497.625 -128.730 -497.345 -128.450 ;
        RECT -497.005 -128.730 -496.725 -128.450 ;
        RECT -496.385 -128.730 -496.105 -128.450 ;
        RECT -495.765 -128.730 -495.485 -128.450 ;
        RECT -495.145 -128.730 -494.865 -128.450 ;
        RECT -494.525 -128.730 -494.245 -128.450 ;
        RECT -493.905 -128.730 -493.625 -128.450 ;
        RECT -499.485 -129.350 -499.205 -129.070 ;
        RECT -498.865 -129.350 -498.585 -129.070 ;
        RECT -498.245 -129.350 -497.965 -129.070 ;
        RECT -497.625 -129.350 -497.345 -129.070 ;
        RECT -497.005 -129.350 -496.725 -129.070 ;
        RECT -496.385 -129.350 -496.105 -129.070 ;
        RECT -495.765 -129.350 -495.485 -129.070 ;
        RECT -495.145 -129.350 -494.865 -129.070 ;
        RECT -494.525 -129.350 -494.245 -129.070 ;
        RECT -493.905 -129.350 -493.625 -129.070 ;
        RECT -499.485 -129.970 -499.205 -129.690 ;
        RECT -498.865 -129.970 -498.585 -129.690 ;
        RECT -498.245 -129.970 -497.965 -129.690 ;
        RECT -497.625 -129.970 -497.345 -129.690 ;
        RECT -497.005 -129.970 -496.725 -129.690 ;
        RECT -496.385 -129.970 -496.105 -129.690 ;
        RECT -495.765 -129.970 -495.485 -129.690 ;
        RECT -495.145 -129.970 -494.865 -129.690 ;
        RECT -494.525 -129.970 -494.245 -129.690 ;
        RECT -493.905 -129.970 -493.625 -129.690 ;
        RECT -499.485 -130.590 -499.205 -130.310 ;
        RECT -498.865 -130.590 -498.585 -130.310 ;
        RECT -498.245 -130.590 -497.965 -130.310 ;
        RECT -497.625 -130.590 -497.345 -130.310 ;
        RECT -497.005 -130.590 -496.725 -130.310 ;
        RECT -496.385 -130.590 -496.105 -130.310 ;
        RECT -495.765 -130.590 -495.485 -130.310 ;
        RECT -495.145 -130.590 -494.865 -130.310 ;
        RECT -494.525 -130.590 -494.245 -130.310 ;
        RECT -493.905 -130.590 -493.625 -130.310 ;
        RECT -499.485 -131.210 -499.205 -130.930 ;
        RECT -498.865 -131.210 -498.585 -130.930 ;
        RECT -498.245 -131.210 -497.965 -130.930 ;
        RECT -497.625 -131.210 -497.345 -130.930 ;
        RECT -497.005 -131.210 -496.725 -130.930 ;
        RECT -496.385 -131.210 -496.105 -130.930 ;
        RECT -495.765 -131.210 -495.485 -130.930 ;
        RECT -495.145 -131.210 -494.865 -130.930 ;
        RECT -494.525 -131.210 -494.245 -130.930 ;
        RECT -493.905 -131.210 -493.625 -130.930 ;
        RECT -499.485 -131.830 -499.205 -131.550 ;
        RECT -498.865 -131.830 -498.585 -131.550 ;
        RECT -498.245 -131.830 -497.965 -131.550 ;
        RECT -497.625 -131.830 -497.345 -131.550 ;
        RECT -497.005 -131.830 -496.725 -131.550 ;
        RECT -496.385 -131.830 -496.105 -131.550 ;
        RECT -495.765 -131.830 -495.485 -131.550 ;
        RECT -495.145 -131.830 -494.865 -131.550 ;
        RECT -494.525 -131.830 -494.245 -131.550 ;
        RECT -493.905 -131.830 -493.625 -131.550 ;
        RECT -499.485 -132.450 -499.205 -132.170 ;
        RECT -498.865 -132.450 -498.585 -132.170 ;
        RECT -498.245 -132.450 -497.965 -132.170 ;
        RECT -497.625 -132.450 -497.345 -132.170 ;
        RECT -497.005 -132.450 -496.725 -132.170 ;
        RECT -496.385 -132.450 -496.105 -132.170 ;
        RECT -495.765 -132.450 -495.485 -132.170 ;
        RECT -495.145 -132.450 -494.865 -132.170 ;
        RECT -494.525 -132.450 -494.245 -132.170 ;
        RECT -493.905 -132.450 -493.625 -132.170 ;
        RECT 146.795 -128.110 147.075 -127.830 ;
        RECT 147.415 -128.110 147.695 -127.830 ;
        RECT 146.795 -128.730 147.075 -128.450 ;
        RECT 147.415 -128.730 147.695 -128.450 ;
        RECT 146.795 -129.350 147.075 -129.070 ;
        RECT 147.415 -129.350 147.695 -129.070 ;
        RECT 146.795 -129.970 147.075 -129.690 ;
        RECT 147.415 -129.970 147.695 -129.690 ;
        RECT 146.795 -130.590 147.075 -130.310 ;
        RECT 147.415 -130.590 147.695 -130.310 ;
        RECT 146.795 -131.210 147.075 -130.930 ;
        RECT 147.415 -131.210 147.695 -130.930 ;
        RECT 146.795 -131.830 147.075 -131.550 ;
        RECT 147.415 -131.830 147.695 -131.550 ;
        RECT 146.795 -132.450 147.075 -132.170 ;
        RECT 147.415 -132.450 147.695 -132.170 ;
      LAYER Metal3 ;
        RECT -499.655 127.660 -493.455 132.620 ;
        RECT 146.625 127.660 147.865 132.620 ;
        RECT 336.790 44.620 338.210 44.900 ;
        RECT 378.370 44.620 379.790 44.900 ;
        RECT 419.950 44.620 421.370 44.900 ;
        RECT 461.530 44.620 462.950 44.900 ;
        RECT 336.790 36.780 338.210 37.060 ;
        RECT 378.370 36.780 379.790 37.060 ;
        RECT 419.950 36.780 421.370 37.060 ;
        RECT 461.530 36.780 462.950 37.060 ;
        RECT 194.795 31.615 195.915 32.635 ;
        RECT 336.790 28.940 338.210 29.220 ;
        RECT 378.370 28.940 379.790 29.220 ;
        RECT 419.950 28.940 421.370 29.220 ;
        RECT 461.530 28.940 462.950 29.220 ;
        RECT 336.790 21.100 338.210 21.380 ;
        RECT 378.370 21.100 379.790 21.380 ;
        RECT 419.950 21.100 421.370 21.380 ;
        RECT 461.530 21.100 462.950 21.380 ;
        RECT 336.790 13.260 338.210 13.540 ;
        RECT 378.370 13.260 379.790 13.540 ;
        RECT 419.950 13.260 421.370 13.540 ;
        RECT 461.530 13.260 462.950 13.540 ;
        RECT 194.795 -0.510 195.915 0.510 ;
        RECT 227.990 0.220 229.590 9.220 ;
        RECT 336.790 5.420 338.210 5.700 ;
        RECT 378.370 5.420 379.790 5.700 ;
        RECT 419.950 5.420 421.370 5.700 ;
        RECT 461.530 5.420 462.950 5.700 ;
        RECT 336.790 -2.420 338.210 -2.140 ;
        RECT 378.370 -2.420 379.790 -2.140 ;
        RECT 419.950 -2.420 421.370 -2.140 ;
        RECT 461.530 -2.420 462.950 -2.140 ;
        RECT 336.790 -10.260 338.210 -9.980 ;
        RECT 378.370 -10.260 379.790 -9.980 ;
        RECT 419.950 -10.260 421.370 -9.980 ;
        RECT 461.530 -10.260 462.950 -9.980 ;
        RECT 229.700 -13.735 235.700 -12.135 ;
        RECT 336.790 -18.100 338.210 -17.820 ;
        RECT 378.370 -18.100 379.790 -17.820 ;
        RECT 419.950 -18.100 421.370 -17.820 ;
        RECT 461.530 -18.100 462.950 -17.820 ;
        RECT 336.790 -25.940 338.210 -25.660 ;
        RECT 378.370 -25.940 379.790 -25.660 ;
        RECT 419.950 -25.940 421.370 -25.660 ;
        RECT 461.530 -25.940 462.950 -25.660 ;
        RECT 194.795 -32.635 195.915 -31.615 ;
        RECT 336.790 -33.780 338.210 -33.500 ;
        RECT 378.370 -33.780 379.790 -33.500 ;
        RECT 419.950 -33.780 421.370 -33.500 ;
        RECT 461.530 -33.780 462.950 -33.500 ;
        RECT 336.790 -41.620 338.210 -41.340 ;
        RECT 378.370 -41.620 379.790 -41.340 ;
        RECT 419.950 -41.620 421.370 -41.340 ;
        RECT 461.530 -41.620 462.950 -41.340 ;
        RECT 336.790 -49.460 338.210 -49.180 ;
        RECT 378.370 -49.460 379.790 -49.180 ;
        RECT 419.950 -49.460 421.370 -49.180 ;
        RECT 461.530 -49.460 462.950 -49.180 ;
        RECT -499.655 -132.620 -493.455 -127.660 ;
        RECT 146.625 -132.620 147.865 -127.660 ;
      LAYER Via3 ;
        RECT -499.485 132.170 -499.205 132.450 ;
        RECT -498.865 132.170 -498.585 132.450 ;
        RECT -498.245 132.170 -497.965 132.450 ;
        RECT -497.625 132.170 -497.345 132.450 ;
        RECT -497.005 132.170 -496.725 132.450 ;
        RECT -496.385 132.170 -496.105 132.450 ;
        RECT -495.765 132.170 -495.485 132.450 ;
        RECT -495.145 132.170 -494.865 132.450 ;
        RECT -494.525 132.170 -494.245 132.450 ;
        RECT -493.905 132.170 -493.625 132.450 ;
        RECT -499.485 131.550 -499.205 131.830 ;
        RECT -498.865 131.550 -498.585 131.830 ;
        RECT -498.245 131.550 -497.965 131.830 ;
        RECT -497.625 131.550 -497.345 131.830 ;
        RECT -497.005 131.550 -496.725 131.830 ;
        RECT -496.385 131.550 -496.105 131.830 ;
        RECT -495.765 131.550 -495.485 131.830 ;
        RECT -495.145 131.550 -494.865 131.830 ;
        RECT -494.525 131.550 -494.245 131.830 ;
        RECT -493.905 131.550 -493.625 131.830 ;
        RECT -499.485 130.930 -499.205 131.210 ;
        RECT -498.865 130.930 -498.585 131.210 ;
        RECT -498.245 130.930 -497.965 131.210 ;
        RECT -497.625 130.930 -497.345 131.210 ;
        RECT -497.005 130.930 -496.725 131.210 ;
        RECT -496.385 130.930 -496.105 131.210 ;
        RECT -495.765 130.930 -495.485 131.210 ;
        RECT -495.145 130.930 -494.865 131.210 ;
        RECT -494.525 130.930 -494.245 131.210 ;
        RECT -493.905 130.930 -493.625 131.210 ;
        RECT -499.485 130.310 -499.205 130.590 ;
        RECT -498.865 130.310 -498.585 130.590 ;
        RECT -498.245 130.310 -497.965 130.590 ;
        RECT -497.625 130.310 -497.345 130.590 ;
        RECT -497.005 130.310 -496.725 130.590 ;
        RECT -496.385 130.310 -496.105 130.590 ;
        RECT -495.765 130.310 -495.485 130.590 ;
        RECT -495.145 130.310 -494.865 130.590 ;
        RECT -494.525 130.310 -494.245 130.590 ;
        RECT -493.905 130.310 -493.625 130.590 ;
        RECT -499.485 129.690 -499.205 129.970 ;
        RECT -498.865 129.690 -498.585 129.970 ;
        RECT -498.245 129.690 -497.965 129.970 ;
        RECT -497.625 129.690 -497.345 129.970 ;
        RECT -497.005 129.690 -496.725 129.970 ;
        RECT -496.385 129.690 -496.105 129.970 ;
        RECT -495.765 129.690 -495.485 129.970 ;
        RECT -495.145 129.690 -494.865 129.970 ;
        RECT -494.525 129.690 -494.245 129.970 ;
        RECT -493.905 129.690 -493.625 129.970 ;
        RECT -499.485 129.070 -499.205 129.350 ;
        RECT -498.865 129.070 -498.585 129.350 ;
        RECT -498.245 129.070 -497.965 129.350 ;
        RECT -497.625 129.070 -497.345 129.350 ;
        RECT -497.005 129.070 -496.725 129.350 ;
        RECT -496.385 129.070 -496.105 129.350 ;
        RECT -495.765 129.070 -495.485 129.350 ;
        RECT -495.145 129.070 -494.865 129.350 ;
        RECT -494.525 129.070 -494.245 129.350 ;
        RECT -493.905 129.070 -493.625 129.350 ;
        RECT -499.485 128.450 -499.205 128.730 ;
        RECT -498.865 128.450 -498.585 128.730 ;
        RECT -498.245 128.450 -497.965 128.730 ;
        RECT -497.625 128.450 -497.345 128.730 ;
        RECT -497.005 128.450 -496.725 128.730 ;
        RECT -496.385 128.450 -496.105 128.730 ;
        RECT -495.765 128.450 -495.485 128.730 ;
        RECT -495.145 128.450 -494.865 128.730 ;
        RECT -494.525 128.450 -494.245 128.730 ;
        RECT -493.905 128.450 -493.625 128.730 ;
        RECT -499.485 127.830 -499.205 128.110 ;
        RECT -498.865 127.830 -498.585 128.110 ;
        RECT -498.245 127.830 -497.965 128.110 ;
        RECT -497.625 127.830 -497.345 128.110 ;
        RECT -497.005 127.830 -496.725 128.110 ;
        RECT -496.385 127.830 -496.105 128.110 ;
        RECT -495.765 127.830 -495.485 128.110 ;
        RECT -495.145 127.830 -494.865 128.110 ;
        RECT -494.525 127.830 -494.245 128.110 ;
        RECT -493.905 127.830 -493.625 128.110 ;
        RECT 146.795 132.170 147.075 132.450 ;
        RECT 147.415 132.170 147.695 132.450 ;
        RECT 146.795 131.550 147.075 131.830 ;
        RECT 147.415 131.550 147.695 131.830 ;
        RECT 146.795 130.930 147.075 131.210 ;
        RECT 147.415 130.930 147.695 131.210 ;
        RECT 146.795 130.310 147.075 130.590 ;
        RECT 147.415 130.310 147.695 130.590 ;
        RECT 146.795 129.690 147.075 129.970 ;
        RECT 147.415 129.690 147.695 129.970 ;
        RECT 146.795 129.070 147.075 129.350 ;
        RECT 147.415 129.070 147.695 129.350 ;
        RECT 146.795 128.450 147.075 128.730 ;
        RECT 147.415 128.450 147.695 128.730 ;
        RECT 146.795 127.830 147.075 128.110 ;
        RECT 147.415 127.830 147.695 128.110 ;
        RECT 336.840 44.620 338.160 44.900 ;
        RECT 378.420 44.620 379.740 44.900 ;
        RECT 420.000 44.620 421.320 44.900 ;
        RECT 461.580 44.620 462.900 44.900 ;
        RECT 336.840 36.780 338.160 37.060 ;
        RECT 378.420 36.780 379.740 37.060 ;
        RECT 420.000 36.780 421.320 37.060 ;
        RECT 461.580 36.780 462.900 37.060 ;
        RECT 194.935 31.725 195.215 32.525 ;
        RECT 195.495 31.725 195.775 32.525 ;
        RECT 336.840 28.940 338.160 29.220 ;
        RECT 378.420 28.940 379.740 29.220 ;
        RECT 420.000 28.940 421.320 29.220 ;
        RECT 461.580 28.940 462.900 29.220 ;
        RECT 336.840 21.100 338.160 21.380 ;
        RECT 378.420 21.100 379.740 21.380 ;
        RECT 420.000 21.100 421.320 21.380 ;
        RECT 461.580 21.100 462.900 21.380 ;
        RECT 336.840 13.260 338.160 13.540 ;
        RECT 378.420 13.260 379.740 13.540 ;
        RECT 420.000 13.260 421.320 13.540 ;
        RECT 461.580 13.260 462.900 13.540 ;
        RECT 228.130 6.540 229.450 8.900 ;
        RECT 228.130 3.540 229.450 5.900 ;
        RECT 336.840 5.420 338.160 5.700 ;
        RECT 378.420 5.420 379.740 5.700 ;
        RECT 420.000 5.420 421.320 5.700 ;
        RECT 461.580 5.420 462.900 5.700 ;
        RECT 228.130 0.540 229.450 2.900 ;
        RECT 194.935 -0.400 195.215 0.400 ;
        RECT 195.495 -0.400 195.775 0.400 ;
        RECT 336.840 -2.420 338.160 -2.140 ;
        RECT 378.420 -2.420 379.740 -2.140 ;
        RECT 420.000 -2.420 421.320 -2.140 ;
        RECT 461.580 -2.420 462.900 -2.140 ;
        RECT 336.840 -10.260 338.160 -9.980 ;
        RECT 378.420 -10.260 379.740 -9.980 ;
        RECT 420.000 -10.260 421.320 -9.980 ;
        RECT 461.580 -10.260 462.900 -9.980 ;
        RECT 230.020 -13.595 232.380 -12.275 ;
        RECT 233.020 -13.595 235.380 -12.275 ;
        RECT 336.840 -18.100 338.160 -17.820 ;
        RECT 378.420 -18.100 379.740 -17.820 ;
        RECT 420.000 -18.100 421.320 -17.820 ;
        RECT 461.580 -18.100 462.900 -17.820 ;
        RECT 336.840 -25.940 338.160 -25.660 ;
        RECT 378.420 -25.940 379.740 -25.660 ;
        RECT 420.000 -25.940 421.320 -25.660 ;
        RECT 461.580 -25.940 462.900 -25.660 ;
        RECT 194.935 -32.525 195.215 -31.725 ;
        RECT 195.495 -32.525 195.775 -31.725 ;
        RECT 336.840 -33.780 338.160 -33.500 ;
        RECT 378.420 -33.780 379.740 -33.500 ;
        RECT 420.000 -33.780 421.320 -33.500 ;
        RECT 461.580 -33.780 462.900 -33.500 ;
        RECT 336.840 -41.620 338.160 -41.340 ;
        RECT 378.420 -41.620 379.740 -41.340 ;
        RECT 420.000 -41.620 421.320 -41.340 ;
        RECT 461.580 -41.620 462.900 -41.340 ;
        RECT 336.840 -49.460 338.160 -49.180 ;
        RECT 378.420 -49.460 379.740 -49.180 ;
        RECT 420.000 -49.460 421.320 -49.180 ;
        RECT 461.580 -49.460 462.900 -49.180 ;
        RECT -499.485 -128.110 -499.205 -127.830 ;
        RECT -498.865 -128.110 -498.585 -127.830 ;
        RECT -498.245 -128.110 -497.965 -127.830 ;
        RECT -497.625 -128.110 -497.345 -127.830 ;
        RECT -497.005 -128.110 -496.725 -127.830 ;
        RECT -496.385 -128.110 -496.105 -127.830 ;
        RECT -495.765 -128.110 -495.485 -127.830 ;
        RECT -495.145 -128.110 -494.865 -127.830 ;
        RECT -494.525 -128.110 -494.245 -127.830 ;
        RECT -493.905 -128.110 -493.625 -127.830 ;
        RECT -499.485 -128.730 -499.205 -128.450 ;
        RECT -498.865 -128.730 -498.585 -128.450 ;
        RECT -498.245 -128.730 -497.965 -128.450 ;
        RECT -497.625 -128.730 -497.345 -128.450 ;
        RECT -497.005 -128.730 -496.725 -128.450 ;
        RECT -496.385 -128.730 -496.105 -128.450 ;
        RECT -495.765 -128.730 -495.485 -128.450 ;
        RECT -495.145 -128.730 -494.865 -128.450 ;
        RECT -494.525 -128.730 -494.245 -128.450 ;
        RECT -493.905 -128.730 -493.625 -128.450 ;
        RECT -499.485 -129.350 -499.205 -129.070 ;
        RECT -498.865 -129.350 -498.585 -129.070 ;
        RECT -498.245 -129.350 -497.965 -129.070 ;
        RECT -497.625 -129.350 -497.345 -129.070 ;
        RECT -497.005 -129.350 -496.725 -129.070 ;
        RECT -496.385 -129.350 -496.105 -129.070 ;
        RECT -495.765 -129.350 -495.485 -129.070 ;
        RECT -495.145 -129.350 -494.865 -129.070 ;
        RECT -494.525 -129.350 -494.245 -129.070 ;
        RECT -493.905 -129.350 -493.625 -129.070 ;
        RECT -499.485 -129.970 -499.205 -129.690 ;
        RECT -498.865 -129.970 -498.585 -129.690 ;
        RECT -498.245 -129.970 -497.965 -129.690 ;
        RECT -497.625 -129.970 -497.345 -129.690 ;
        RECT -497.005 -129.970 -496.725 -129.690 ;
        RECT -496.385 -129.970 -496.105 -129.690 ;
        RECT -495.765 -129.970 -495.485 -129.690 ;
        RECT -495.145 -129.970 -494.865 -129.690 ;
        RECT -494.525 -129.970 -494.245 -129.690 ;
        RECT -493.905 -129.970 -493.625 -129.690 ;
        RECT -499.485 -130.590 -499.205 -130.310 ;
        RECT -498.865 -130.590 -498.585 -130.310 ;
        RECT -498.245 -130.590 -497.965 -130.310 ;
        RECT -497.625 -130.590 -497.345 -130.310 ;
        RECT -497.005 -130.590 -496.725 -130.310 ;
        RECT -496.385 -130.590 -496.105 -130.310 ;
        RECT -495.765 -130.590 -495.485 -130.310 ;
        RECT -495.145 -130.590 -494.865 -130.310 ;
        RECT -494.525 -130.590 -494.245 -130.310 ;
        RECT -493.905 -130.590 -493.625 -130.310 ;
        RECT -499.485 -131.210 -499.205 -130.930 ;
        RECT -498.865 -131.210 -498.585 -130.930 ;
        RECT -498.245 -131.210 -497.965 -130.930 ;
        RECT -497.625 -131.210 -497.345 -130.930 ;
        RECT -497.005 -131.210 -496.725 -130.930 ;
        RECT -496.385 -131.210 -496.105 -130.930 ;
        RECT -495.765 -131.210 -495.485 -130.930 ;
        RECT -495.145 -131.210 -494.865 -130.930 ;
        RECT -494.525 -131.210 -494.245 -130.930 ;
        RECT -493.905 -131.210 -493.625 -130.930 ;
        RECT -499.485 -131.830 -499.205 -131.550 ;
        RECT -498.865 -131.830 -498.585 -131.550 ;
        RECT -498.245 -131.830 -497.965 -131.550 ;
        RECT -497.625 -131.830 -497.345 -131.550 ;
        RECT -497.005 -131.830 -496.725 -131.550 ;
        RECT -496.385 -131.830 -496.105 -131.550 ;
        RECT -495.765 -131.830 -495.485 -131.550 ;
        RECT -495.145 -131.830 -494.865 -131.550 ;
        RECT -494.525 -131.830 -494.245 -131.550 ;
        RECT -493.905 -131.830 -493.625 -131.550 ;
        RECT -499.485 -132.450 -499.205 -132.170 ;
        RECT -498.865 -132.450 -498.585 -132.170 ;
        RECT -498.245 -132.450 -497.965 -132.170 ;
        RECT -497.625 -132.450 -497.345 -132.170 ;
        RECT -497.005 -132.450 -496.725 -132.170 ;
        RECT -496.385 -132.450 -496.105 -132.170 ;
        RECT -495.765 -132.450 -495.485 -132.170 ;
        RECT -495.145 -132.450 -494.865 -132.170 ;
        RECT -494.525 -132.450 -494.245 -132.170 ;
        RECT -493.905 -132.450 -493.625 -132.170 ;
        RECT 146.795 -128.110 147.075 -127.830 ;
        RECT 147.415 -128.110 147.695 -127.830 ;
        RECT 146.795 -128.730 147.075 -128.450 ;
        RECT 147.415 -128.730 147.695 -128.450 ;
        RECT 146.795 -129.350 147.075 -129.070 ;
        RECT 147.415 -129.350 147.695 -129.070 ;
        RECT 146.795 -129.970 147.075 -129.690 ;
        RECT 147.415 -129.970 147.695 -129.690 ;
        RECT 146.795 -130.590 147.075 -130.310 ;
        RECT 147.415 -130.590 147.695 -130.310 ;
        RECT 146.795 -131.210 147.075 -130.930 ;
        RECT 147.415 -131.210 147.695 -130.930 ;
        RECT 146.795 -131.830 147.075 -131.550 ;
        RECT 147.415 -131.830 147.695 -131.550 ;
        RECT 146.795 -132.450 147.075 -132.170 ;
        RECT 147.415 -132.450 147.695 -132.170 ;
      LAYER Metal4 ;
        RECT -838.480 1085.700 841.320 1163.700 ;
        RECT -838.480 352.720 -760.480 1085.700 ;
        RECT -557.530 945.220 -525.130 945.820 ;
        RECT -557.530 915.220 -556.930 945.220 ;
        RECT -526.930 915.220 -525.130 945.220 ;
        RECT -557.530 914.620 -525.130 915.220 ;
        RECT -521.830 945.220 -489.430 945.820 ;
        RECT -521.830 915.220 -520.030 945.220 ;
        RECT -490.030 915.220 -489.430 945.220 ;
        RECT -521.830 914.620 -489.430 915.220 ;
        RECT -482.530 945.220 -450.130 945.820 ;
        RECT -482.530 915.220 -481.930 945.220 ;
        RECT -451.930 915.220 -450.130 945.220 ;
        RECT -482.530 914.620 -450.130 915.220 ;
        RECT -446.830 945.220 -414.430 945.820 ;
        RECT -446.830 915.220 -445.030 945.220 ;
        RECT -415.030 915.220 -414.430 945.220 ;
        RECT -446.830 914.620 -414.430 915.220 ;
        RECT -407.530 945.220 -375.130 945.820 ;
        RECT -407.530 915.220 -406.930 945.220 ;
        RECT -376.930 915.220 -375.130 945.220 ;
        RECT -407.530 914.620 -375.130 915.220 ;
        RECT -371.830 945.220 -339.430 945.820 ;
        RECT -371.830 915.220 -370.030 945.220 ;
        RECT -340.030 915.220 -339.430 945.220 ;
        RECT -371.830 914.620 -339.430 915.220 ;
        RECT -332.530 945.220 -300.130 945.820 ;
        RECT -332.530 915.220 -331.930 945.220 ;
        RECT -301.930 915.220 -300.130 945.220 ;
        RECT -332.530 914.620 -300.130 915.220 ;
        RECT -296.830 945.220 -264.430 945.820 ;
        RECT -296.830 915.220 -295.030 945.220 ;
        RECT -265.030 915.220 -264.430 945.220 ;
        RECT -296.830 914.620 -264.430 915.220 ;
        RECT -257.530 945.220 -225.130 945.820 ;
        RECT -257.530 915.220 -256.930 945.220 ;
        RECT -226.930 915.220 -225.130 945.220 ;
        RECT -257.530 914.620 -225.130 915.220 ;
        RECT -221.830 945.220 -189.430 945.820 ;
        RECT -221.830 915.220 -220.030 945.220 ;
        RECT -190.030 915.220 -189.430 945.220 ;
        RECT -221.830 914.620 -189.430 915.220 ;
        RECT -182.530 945.220 -150.130 945.820 ;
        RECT -182.530 915.220 -181.930 945.220 ;
        RECT -151.930 915.220 -150.130 945.220 ;
        RECT -182.530 914.620 -150.130 915.220 ;
        RECT -146.830 945.220 -114.430 945.820 ;
        RECT -146.830 915.220 -145.030 945.220 ;
        RECT -115.030 915.220 -114.430 945.220 ;
        RECT -146.830 914.620 -114.430 915.220 ;
        RECT -107.530 945.220 -75.130 945.820 ;
        RECT -107.530 915.220 -106.930 945.220 ;
        RECT -76.930 915.220 -75.130 945.220 ;
        RECT -107.530 914.620 -75.130 915.220 ;
        RECT -71.830 945.220 -39.430 945.820 ;
        RECT -71.830 915.220 -70.030 945.220 ;
        RECT -40.030 915.220 -39.430 945.220 ;
        RECT -71.830 914.620 -39.430 915.220 ;
        RECT -32.530 945.220 -0.130 945.820 ;
        RECT -32.530 915.220 -31.930 945.220 ;
        RECT -1.930 915.220 -0.130 945.220 ;
        RECT -32.530 914.620 -0.130 915.220 ;
        RECT 3.170 945.220 35.570 945.820 ;
        RECT 3.170 915.220 4.970 945.220 ;
        RECT 34.970 915.220 35.570 945.220 ;
        RECT 3.170 914.620 35.570 915.220 ;
        RECT 42.470 945.220 74.870 945.820 ;
        RECT 42.470 915.220 43.070 945.220 ;
        RECT 73.070 915.220 74.870 945.220 ;
        RECT 42.470 914.620 74.870 915.220 ;
        RECT 78.170 945.220 110.570 945.820 ;
        RECT 78.170 915.220 79.970 945.220 ;
        RECT 109.970 915.220 110.570 945.220 ;
        RECT 78.170 914.620 110.570 915.220 ;
        RECT 117.470 945.220 149.870 945.820 ;
        RECT 117.470 915.220 118.070 945.220 ;
        RECT 148.070 915.220 149.870 945.220 ;
        RECT 117.470 914.620 149.870 915.220 ;
        RECT 153.170 945.220 185.570 945.820 ;
        RECT 153.170 915.220 154.970 945.220 ;
        RECT 184.970 915.220 185.570 945.220 ;
        RECT 153.170 914.620 185.570 915.220 ;
        RECT 192.470 945.220 224.870 945.820 ;
        RECT 192.470 915.220 193.070 945.220 ;
        RECT 223.070 915.220 224.870 945.220 ;
        RECT 192.470 914.620 224.870 915.220 ;
        RECT 228.170 945.220 260.570 945.820 ;
        RECT 228.170 915.220 229.970 945.220 ;
        RECT 259.970 915.220 260.570 945.220 ;
        RECT 228.170 914.620 260.570 915.220 ;
        RECT 267.470 945.220 299.870 945.820 ;
        RECT 267.470 915.220 268.070 945.220 ;
        RECT 298.070 915.220 299.870 945.220 ;
        RECT 267.470 914.620 299.870 915.220 ;
        RECT 303.170 945.220 335.570 945.820 ;
        RECT 303.170 915.220 304.970 945.220 ;
        RECT 334.970 915.220 335.570 945.220 ;
        RECT 303.170 914.620 335.570 915.220 ;
        RECT 342.470 945.220 374.870 945.820 ;
        RECT 342.470 915.220 343.070 945.220 ;
        RECT 373.070 915.220 374.870 945.220 ;
        RECT 342.470 914.620 374.870 915.220 ;
        RECT 378.170 945.220 410.570 945.820 ;
        RECT 378.170 915.220 379.970 945.220 ;
        RECT 409.970 915.220 410.570 945.220 ;
        RECT 378.170 914.620 410.570 915.220 ;
        RECT 417.470 945.220 449.870 945.820 ;
        RECT 417.470 915.220 418.070 945.220 ;
        RECT 448.070 915.220 449.870 945.220 ;
        RECT 417.470 914.620 449.870 915.220 ;
        RECT 453.170 945.220 485.570 945.820 ;
        RECT 453.170 915.220 454.970 945.220 ;
        RECT 484.970 915.220 485.570 945.220 ;
        RECT 453.170 914.620 485.570 915.220 ;
        RECT 492.470 945.220 524.870 945.820 ;
        RECT 492.470 915.220 493.070 945.220 ;
        RECT 523.070 915.220 524.870 945.220 ;
        RECT 492.470 914.620 524.870 915.220 ;
        RECT 528.170 945.220 560.570 945.820 ;
        RECT 528.170 915.220 529.970 945.220 ;
        RECT 559.970 915.220 560.570 945.220 ;
        RECT 528.170 914.620 560.570 915.220 ;
        RECT -557.530 910.220 -525.130 910.820 ;
        RECT -557.530 880.220 -556.930 910.220 ;
        RECT -526.930 880.220 -525.130 910.220 ;
        RECT -557.530 879.620 -525.130 880.220 ;
        RECT -521.830 910.220 -489.430 910.820 ;
        RECT -521.830 880.220 -520.030 910.220 ;
        RECT -490.030 880.220 -489.430 910.220 ;
        RECT -521.830 879.620 -489.430 880.220 ;
        RECT -482.530 910.220 -450.130 910.820 ;
        RECT -482.530 880.220 -481.930 910.220 ;
        RECT -451.930 880.220 -450.130 910.220 ;
        RECT -482.530 879.620 -450.130 880.220 ;
        RECT -446.830 910.220 -414.430 910.820 ;
        RECT -446.830 880.220 -445.030 910.220 ;
        RECT -415.030 880.220 -414.430 910.220 ;
        RECT -446.830 879.620 -414.430 880.220 ;
        RECT -407.530 910.220 -375.130 910.820 ;
        RECT -407.530 880.220 -406.930 910.220 ;
        RECT -376.930 880.220 -375.130 910.220 ;
        RECT -407.530 879.620 -375.130 880.220 ;
        RECT -371.830 910.220 -339.430 910.820 ;
        RECT -371.830 880.220 -370.030 910.220 ;
        RECT -340.030 880.220 -339.430 910.220 ;
        RECT -371.830 879.620 -339.430 880.220 ;
        RECT -332.530 910.220 -300.130 910.820 ;
        RECT -332.530 880.220 -331.930 910.220 ;
        RECT -301.930 880.220 -300.130 910.220 ;
        RECT -332.530 879.620 -300.130 880.220 ;
        RECT -296.830 910.220 -264.430 910.820 ;
        RECT -296.830 880.220 -295.030 910.220 ;
        RECT -265.030 880.220 -264.430 910.220 ;
        RECT -296.830 879.620 -264.430 880.220 ;
        RECT -257.530 910.220 -225.130 910.820 ;
        RECT -257.530 880.220 -256.930 910.220 ;
        RECT -226.930 880.220 -225.130 910.220 ;
        RECT -257.530 879.620 -225.130 880.220 ;
        RECT -221.830 910.220 -189.430 910.820 ;
        RECT -221.830 880.220 -220.030 910.220 ;
        RECT -190.030 880.220 -189.430 910.220 ;
        RECT -221.830 879.620 -189.430 880.220 ;
        RECT -182.530 910.220 -150.130 910.820 ;
        RECT -182.530 880.220 -181.930 910.220 ;
        RECT -151.930 880.220 -150.130 910.220 ;
        RECT -182.530 879.620 -150.130 880.220 ;
        RECT -146.830 910.220 -114.430 910.820 ;
        RECT -146.830 880.220 -145.030 910.220 ;
        RECT -115.030 880.220 -114.430 910.220 ;
        RECT -146.830 879.620 -114.430 880.220 ;
        RECT -107.530 910.220 -75.130 910.820 ;
        RECT -107.530 880.220 -106.930 910.220 ;
        RECT -76.930 880.220 -75.130 910.220 ;
        RECT -107.530 879.620 -75.130 880.220 ;
        RECT -71.830 910.220 -39.430 910.820 ;
        RECT -71.830 880.220 -70.030 910.220 ;
        RECT -40.030 880.220 -39.430 910.220 ;
        RECT -71.830 879.620 -39.430 880.220 ;
        RECT -32.530 910.220 -0.130 910.820 ;
        RECT -32.530 880.220 -31.930 910.220 ;
        RECT -1.930 880.220 -0.130 910.220 ;
        RECT -32.530 879.620 -0.130 880.220 ;
        RECT 3.170 910.220 35.570 910.820 ;
        RECT 3.170 880.220 4.970 910.220 ;
        RECT 34.970 880.220 35.570 910.220 ;
        RECT 3.170 879.620 35.570 880.220 ;
        RECT 42.470 910.220 74.870 910.820 ;
        RECT 42.470 880.220 43.070 910.220 ;
        RECT 73.070 880.220 74.870 910.220 ;
        RECT 42.470 879.620 74.870 880.220 ;
        RECT 78.170 910.220 110.570 910.820 ;
        RECT 78.170 880.220 79.970 910.220 ;
        RECT 109.970 880.220 110.570 910.220 ;
        RECT 78.170 879.620 110.570 880.220 ;
        RECT 117.470 910.220 149.870 910.820 ;
        RECT 117.470 880.220 118.070 910.220 ;
        RECT 148.070 880.220 149.870 910.220 ;
        RECT 117.470 879.620 149.870 880.220 ;
        RECT 153.170 910.220 185.570 910.820 ;
        RECT 153.170 880.220 154.970 910.220 ;
        RECT 184.970 880.220 185.570 910.220 ;
        RECT 153.170 879.620 185.570 880.220 ;
        RECT 192.470 910.220 224.870 910.820 ;
        RECT 192.470 880.220 193.070 910.220 ;
        RECT 223.070 880.220 224.870 910.220 ;
        RECT 192.470 879.620 224.870 880.220 ;
        RECT 228.170 910.220 260.570 910.820 ;
        RECT 228.170 880.220 229.970 910.220 ;
        RECT 259.970 880.220 260.570 910.220 ;
        RECT 228.170 879.620 260.570 880.220 ;
        RECT 267.470 910.220 299.870 910.820 ;
        RECT 267.470 880.220 268.070 910.220 ;
        RECT 298.070 880.220 299.870 910.220 ;
        RECT 267.470 879.620 299.870 880.220 ;
        RECT 303.170 910.220 335.570 910.820 ;
        RECT 303.170 880.220 304.970 910.220 ;
        RECT 334.970 880.220 335.570 910.220 ;
        RECT 303.170 879.620 335.570 880.220 ;
        RECT 342.470 910.220 374.870 910.820 ;
        RECT 342.470 880.220 343.070 910.220 ;
        RECT 373.070 880.220 374.870 910.220 ;
        RECT 342.470 879.620 374.870 880.220 ;
        RECT 378.170 910.220 410.570 910.820 ;
        RECT 378.170 880.220 379.970 910.220 ;
        RECT 409.970 880.220 410.570 910.220 ;
        RECT 378.170 879.620 410.570 880.220 ;
        RECT 417.470 910.220 449.870 910.820 ;
        RECT 417.470 880.220 418.070 910.220 ;
        RECT 448.070 880.220 449.870 910.220 ;
        RECT 417.470 879.620 449.870 880.220 ;
        RECT 453.170 910.220 485.570 910.820 ;
        RECT 453.170 880.220 454.970 910.220 ;
        RECT 484.970 880.220 485.570 910.220 ;
        RECT 453.170 879.620 485.570 880.220 ;
        RECT 492.470 910.220 524.870 910.820 ;
        RECT 492.470 880.220 493.070 910.220 ;
        RECT 523.070 880.220 524.870 910.220 ;
        RECT 492.470 879.620 524.870 880.220 ;
        RECT 528.170 910.220 560.570 910.820 ;
        RECT 528.170 880.220 529.970 910.220 ;
        RECT 559.970 880.220 560.570 910.220 ;
        RECT 528.170 879.620 560.570 880.220 ;
        RECT -557.530 875.220 -525.130 875.820 ;
        RECT -557.530 845.220 -556.930 875.220 ;
        RECT -526.930 845.220 -525.130 875.220 ;
        RECT -557.530 844.620 -525.130 845.220 ;
        RECT -521.830 875.220 -489.430 875.820 ;
        RECT -521.830 845.220 -520.030 875.220 ;
        RECT -490.030 845.220 -489.430 875.220 ;
        RECT -521.830 844.620 -489.430 845.220 ;
        RECT -482.530 875.220 -450.130 875.820 ;
        RECT -482.530 845.220 -481.930 875.220 ;
        RECT -451.930 845.220 -450.130 875.220 ;
        RECT -482.530 844.620 -450.130 845.220 ;
        RECT -446.830 875.220 -414.430 875.820 ;
        RECT -446.830 845.220 -445.030 875.220 ;
        RECT -415.030 845.220 -414.430 875.220 ;
        RECT -446.830 844.620 -414.430 845.220 ;
        RECT -407.530 875.220 -375.130 875.820 ;
        RECT -407.530 845.220 -406.930 875.220 ;
        RECT -376.930 845.220 -375.130 875.220 ;
        RECT -407.530 844.620 -375.130 845.220 ;
        RECT -371.830 875.220 -339.430 875.820 ;
        RECT -371.830 845.220 -370.030 875.220 ;
        RECT -340.030 845.220 -339.430 875.220 ;
        RECT -371.830 844.620 -339.430 845.220 ;
        RECT -332.530 875.220 -300.130 875.820 ;
        RECT -332.530 845.220 -331.930 875.220 ;
        RECT -301.930 845.220 -300.130 875.220 ;
        RECT -332.530 844.620 -300.130 845.220 ;
        RECT -296.830 875.220 -264.430 875.820 ;
        RECT -296.830 845.220 -295.030 875.220 ;
        RECT -265.030 845.220 -264.430 875.220 ;
        RECT -296.830 844.620 -264.430 845.220 ;
        RECT -257.530 875.220 -225.130 875.820 ;
        RECT -257.530 845.220 -256.930 875.220 ;
        RECT -226.930 845.220 -225.130 875.220 ;
        RECT -257.530 844.620 -225.130 845.220 ;
        RECT -221.830 875.220 -189.430 875.820 ;
        RECT -221.830 845.220 -220.030 875.220 ;
        RECT -190.030 845.220 -189.430 875.220 ;
        RECT -221.830 844.620 -189.430 845.220 ;
        RECT -182.530 875.220 -150.130 875.820 ;
        RECT -182.530 845.220 -181.930 875.220 ;
        RECT -151.930 845.220 -150.130 875.220 ;
        RECT -182.530 844.620 -150.130 845.220 ;
        RECT -146.830 875.220 -114.430 875.820 ;
        RECT -146.830 845.220 -145.030 875.220 ;
        RECT -115.030 845.220 -114.430 875.220 ;
        RECT -146.830 844.620 -114.430 845.220 ;
        RECT -107.530 875.220 -75.130 875.820 ;
        RECT -107.530 845.220 -106.930 875.220 ;
        RECT -76.930 845.220 -75.130 875.220 ;
        RECT -107.530 844.620 -75.130 845.220 ;
        RECT -71.830 875.220 -39.430 875.820 ;
        RECT -71.830 845.220 -70.030 875.220 ;
        RECT -40.030 845.220 -39.430 875.220 ;
        RECT -71.830 844.620 -39.430 845.220 ;
        RECT -32.530 875.220 -0.130 875.820 ;
        RECT -32.530 845.220 -31.930 875.220 ;
        RECT -1.930 845.220 -0.130 875.220 ;
        RECT -32.530 844.620 -0.130 845.220 ;
        RECT 3.170 875.220 35.570 875.820 ;
        RECT 3.170 845.220 4.970 875.220 ;
        RECT 34.970 845.220 35.570 875.220 ;
        RECT 3.170 844.620 35.570 845.220 ;
        RECT 42.470 875.220 74.870 875.820 ;
        RECT 42.470 845.220 43.070 875.220 ;
        RECT 73.070 845.220 74.870 875.220 ;
        RECT 42.470 844.620 74.870 845.220 ;
        RECT 78.170 875.220 110.570 875.820 ;
        RECT 78.170 845.220 79.970 875.220 ;
        RECT 109.970 845.220 110.570 875.220 ;
        RECT 78.170 844.620 110.570 845.220 ;
        RECT 117.470 875.220 149.870 875.820 ;
        RECT 117.470 845.220 118.070 875.220 ;
        RECT 148.070 845.220 149.870 875.220 ;
        RECT 117.470 844.620 149.870 845.220 ;
        RECT 153.170 875.220 185.570 875.820 ;
        RECT 153.170 845.220 154.970 875.220 ;
        RECT 184.970 845.220 185.570 875.220 ;
        RECT 153.170 844.620 185.570 845.220 ;
        RECT 192.470 875.220 224.870 875.820 ;
        RECT 192.470 845.220 193.070 875.220 ;
        RECT 223.070 845.220 224.870 875.220 ;
        RECT 192.470 844.620 224.870 845.220 ;
        RECT 228.170 875.220 260.570 875.820 ;
        RECT 228.170 845.220 229.970 875.220 ;
        RECT 259.970 845.220 260.570 875.220 ;
        RECT 228.170 844.620 260.570 845.220 ;
        RECT 267.470 875.220 299.870 875.820 ;
        RECT 267.470 845.220 268.070 875.220 ;
        RECT 298.070 845.220 299.870 875.220 ;
        RECT 267.470 844.620 299.870 845.220 ;
        RECT 303.170 875.220 335.570 875.820 ;
        RECT 303.170 845.220 304.970 875.220 ;
        RECT 334.970 845.220 335.570 875.220 ;
        RECT 303.170 844.620 335.570 845.220 ;
        RECT 342.470 875.220 374.870 875.820 ;
        RECT 342.470 845.220 343.070 875.220 ;
        RECT 373.070 845.220 374.870 875.220 ;
        RECT 342.470 844.620 374.870 845.220 ;
        RECT 378.170 875.220 410.570 875.820 ;
        RECT 378.170 845.220 379.970 875.220 ;
        RECT 409.970 845.220 410.570 875.220 ;
        RECT 378.170 844.620 410.570 845.220 ;
        RECT 417.470 875.220 449.870 875.820 ;
        RECT 417.470 845.220 418.070 875.220 ;
        RECT 448.070 845.220 449.870 875.220 ;
        RECT 417.470 844.620 449.870 845.220 ;
        RECT 453.170 875.220 485.570 875.820 ;
        RECT 453.170 845.220 454.970 875.220 ;
        RECT 484.970 845.220 485.570 875.220 ;
        RECT 453.170 844.620 485.570 845.220 ;
        RECT 492.470 875.220 524.870 875.820 ;
        RECT 492.470 845.220 493.070 875.220 ;
        RECT 523.070 845.220 524.870 875.220 ;
        RECT 492.470 844.620 524.870 845.220 ;
        RECT 528.170 875.220 560.570 875.820 ;
        RECT 528.170 845.220 529.970 875.220 ;
        RECT 559.970 845.220 560.570 875.220 ;
        RECT 528.170 844.620 560.570 845.220 ;
        RECT -557.530 840.220 -525.130 840.820 ;
        RECT -557.530 810.220 -556.930 840.220 ;
        RECT -526.930 810.220 -525.130 840.220 ;
        RECT -557.530 809.620 -525.130 810.220 ;
        RECT -521.830 840.220 -489.430 840.820 ;
        RECT -521.830 810.220 -520.030 840.220 ;
        RECT -490.030 810.220 -489.430 840.220 ;
        RECT -521.830 809.620 -489.430 810.220 ;
        RECT -482.530 840.220 -450.130 840.820 ;
        RECT -482.530 810.220 -481.930 840.220 ;
        RECT -451.930 810.220 -450.130 840.220 ;
        RECT -482.530 809.620 -450.130 810.220 ;
        RECT -446.830 840.220 -414.430 840.820 ;
        RECT -446.830 810.220 -445.030 840.220 ;
        RECT -415.030 810.220 -414.430 840.220 ;
        RECT -446.830 809.620 -414.430 810.220 ;
        RECT -407.530 840.220 -375.130 840.820 ;
        RECT -407.530 810.220 -406.930 840.220 ;
        RECT -376.930 810.220 -375.130 840.220 ;
        RECT -407.530 809.620 -375.130 810.220 ;
        RECT -371.830 840.220 -339.430 840.820 ;
        RECT -371.830 810.220 -370.030 840.220 ;
        RECT -340.030 810.220 -339.430 840.220 ;
        RECT -371.830 809.620 -339.430 810.220 ;
        RECT -332.530 840.220 -300.130 840.820 ;
        RECT -332.530 810.220 -331.930 840.220 ;
        RECT -301.930 810.220 -300.130 840.220 ;
        RECT -332.530 809.620 -300.130 810.220 ;
        RECT -296.830 840.220 -264.430 840.820 ;
        RECT -296.830 810.220 -295.030 840.220 ;
        RECT -265.030 810.220 -264.430 840.220 ;
        RECT -296.830 809.620 -264.430 810.220 ;
        RECT -257.530 840.220 -225.130 840.820 ;
        RECT -257.530 810.220 -256.930 840.220 ;
        RECT -226.930 810.220 -225.130 840.220 ;
        RECT -257.530 809.620 -225.130 810.220 ;
        RECT -221.830 840.220 -189.430 840.820 ;
        RECT -221.830 810.220 -220.030 840.220 ;
        RECT -190.030 810.220 -189.430 840.220 ;
        RECT -221.830 809.620 -189.430 810.220 ;
        RECT -182.530 840.220 -150.130 840.820 ;
        RECT -182.530 810.220 -181.930 840.220 ;
        RECT -151.930 810.220 -150.130 840.220 ;
        RECT -182.530 809.620 -150.130 810.220 ;
        RECT -146.830 840.220 -114.430 840.820 ;
        RECT -146.830 810.220 -145.030 840.220 ;
        RECT -115.030 810.220 -114.430 840.220 ;
        RECT -146.830 809.620 -114.430 810.220 ;
        RECT -107.530 840.220 -75.130 840.820 ;
        RECT -107.530 810.220 -106.930 840.220 ;
        RECT -76.930 810.220 -75.130 840.220 ;
        RECT -107.530 809.620 -75.130 810.220 ;
        RECT -71.830 840.220 -39.430 840.820 ;
        RECT -71.830 810.220 -70.030 840.220 ;
        RECT -40.030 810.220 -39.430 840.220 ;
        RECT -71.830 809.620 -39.430 810.220 ;
        RECT -32.530 840.220 -0.130 840.820 ;
        RECT -32.530 810.220 -31.930 840.220 ;
        RECT -1.930 810.220 -0.130 840.220 ;
        RECT -32.530 809.620 -0.130 810.220 ;
        RECT 3.170 840.220 35.570 840.820 ;
        RECT 3.170 810.220 4.970 840.220 ;
        RECT 34.970 810.220 35.570 840.220 ;
        RECT 3.170 809.620 35.570 810.220 ;
        RECT 42.470 840.220 74.870 840.820 ;
        RECT 42.470 810.220 43.070 840.220 ;
        RECT 73.070 810.220 74.870 840.220 ;
        RECT 42.470 809.620 74.870 810.220 ;
        RECT 78.170 840.220 110.570 840.820 ;
        RECT 78.170 810.220 79.970 840.220 ;
        RECT 109.970 810.220 110.570 840.220 ;
        RECT 78.170 809.620 110.570 810.220 ;
        RECT 117.470 840.220 149.870 840.820 ;
        RECT 117.470 810.220 118.070 840.220 ;
        RECT 148.070 810.220 149.870 840.220 ;
        RECT 117.470 809.620 149.870 810.220 ;
        RECT 153.170 840.220 185.570 840.820 ;
        RECT 153.170 810.220 154.970 840.220 ;
        RECT 184.970 810.220 185.570 840.220 ;
        RECT 153.170 809.620 185.570 810.220 ;
        RECT 192.470 840.220 224.870 840.820 ;
        RECT 192.470 810.220 193.070 840.220 ;
        RECT 223.070 810.220 224.870 840.220 ;
        RECT 192.470 809.620 224.870 810.220 ;
        RECT 228.170 840.220 260.570 840.820 ;
        RECT 228.170 810.220 229.970 840.220 ;
        RECT 259.970 810.220 260.570 840.220 ;
        RECT 228.170 809.620 260.570 810.220 ;
        RECT 267.470 840.220 299.870 840.820 ;
        RECT 267.470 810.220 268.070 840.220 ;
        RECT 298.070 810.220 299.870 840.220 ;
        RECT 267.470 809.620 299.870 810.220 ;
        RECT 303.170 840.220 335.570 840.820 ;
        RECT 303.170 810.220 304.970 840.220 ;
        RECT 334.970 810.220 335.570 840.220 ;
        RECT 303.170 809.620 335.570 810.220 ;
        RECT 342.470 840.220 374.870 840.820 ;
        RECT 342.470 810.220 343.070 840.220 ;
        RECT 373.070 810.220 374.870 840.220 ;
        RECT 342.470 809.620 374.870 810.220 ;
        RECT 378.170 840.220 410.570 840.820 ;
        RECT 378.170 810.220 379.970 840.220 ;
        RECT 409.970 810.220 410.570 840.220 ;
        RECT 378.170 809.620 410.570 810.220 ;
        RECT 417.470 840.220 449.870 840.820 ;
        RECT 417.470 810.220 418.070 840.220 ;
        RECT 448.070 810.220 449.870 840.220 ;
        RECT 417.470 809.620 449.870 810.220 ;
        RECT 453.170 840.220 485.570 840.820 ;
        RECT 453.170 810.220 454.970 840.220 ;
        RECT 484.970 810.220 485.570 840.220 ;
        RECT 453.170 809.620 485.570 810.220 ;
        RECT 492.470 840.220 524.870 840.820 ;
        RECT 492.470 810.220 493.070 840.220 ;
        RECT 523.070 810.220 524.870 840.220 ;
        RECT 492.470 809.620 524.870 810.220 ;
        RECT 528.170 840.220 560.570 840.820 ;
        RECT 528.170 810.220 529.970 840.220 ;
        RECT 559.970 810.220 560.570 840.220 ;
        RECT 528.170 809.620 560.570 810.220 ;
        RECT -557.530 805.220 -525.130 805.820 ;
        RECT -557.530 775.220 -556.930 805.220 ;
        RECT -526.930 775.220 -525.130 805.220 ;
        RECT -557.530 774.620 -525.130 775.220 ;
        RECT -521.830 805.220 -489.430 805.820 ;
        RECT -521.830 775.220 -520.030 805.220 ;
        RECT -490.030 775.220 -489.430 805.220 ;
        RECT -521.830 774.620 -489.430 775.220 ;
        RECT -482.530 805.220 -450.130 805.820 ;
        RECT -482.530 775.220 -481.930 805.220 ;
        RECT -451.930 775.220 -450.130 805.220 ;
        RECT -482.530 774.620 -450.130 775.220 ;
        RECT -446.830 805.220 -414.430 805.820 ;
        RECT -446.830 775.220 -445.030 805.220 ;
        RECT -415.030 775.220 -414.430 805.220 ;
        RECT -446.830 774.620 -414.430 775.220 ;
        RECT -407.530 805.220 -375.130 805.820 ;
        RECT -407.530 775.220 -406.930 805.220 ;
        RECT -376.930 775.220 -375.130 805.220 ;
        RECT -407.530 774.620 -375.130 775.220 ;
        RECT -371.830 805.220 -339.430 805.820 ;
        RECT -371.830 775.220 -370.030 805.220 ;
        RECT -340.030 775.220 -339.430 805.220 ;
        RECT -371.830 774.620 -339.430 775.220 ;
        RECT -332.530 805.220 -300.130 805.820 ;
        RECT -332.530 775.220 -331.930 805.220 ;
        RECT -301.930 775.220 -300.130 805.220 ;
        RECT -332.530 774.620 -300.130 775.220 ;
        RECT -296.830 805.220 -264.430 805.820 ;
        RECT -296.830 775.220 -295.030 805.220 ;
        RECT -265.030 775.220 -264.430 805.220 ;
        RECT -296.830 774.620 -264.430 775.220 ;
        RECT -257.530 805.220 -225.130 805.820 ;
        RECT -257.530 775.220 -256.930 805.220 ;
        RECT -226.930 775.220 -225.130 805.220 ;
        RECT -257.530 774.620 -225.130 775.220 ;
        RECT -221.830 805.220 -189.430 805.820 ;
        RECT -221.830 775.220 -220.030 805.220 ;
        RECT -190.030 775.220 -189.430 805.220 ;
        RECT -221.830 774.620 -189.430 775.220 ;
        RECT -182.530 805.220 -150.130 805.820 ;
        RECT -182.530 775.220 -181.930 805.220 ;
        RECT -151.930 775.220 -150.130 805.220 ;
        RECT -182.530 774.620 -150.130 775.220 ;
        RECT -146.830 805.220 -114.430 805.820 ;
        RECT -146.830 775.220 -145.030 805.220 ;
        RECT -115.030 775.220 -114.430 805.220 ;
        RECT -146.830 774.620 -114.430 775.220 ;
        RECT -107.530 805.220 -75.130 805.820 ;
        RECT -107.530 775.220 -106.930 805.220 ;
        RECT -76.930 775.220 -75.130 805.220 ;
        RECT -107.530 774.620 -75.130 775.220 ;
        RECT -71.830 805.220 -39.430 805.820 ;
        RECT -71.830 775.220 -70.030 805.220 ;
        RECT -40.030 775.220 -39.430 805.220 ;
        RECT -71.830 774.620 -39.430 775.220 ;
        RECT -32.530 805.220 -0.130 805.820 ;
        RECT -32.530 775.220 -31.930 805.220 ;
        RECT -1.930 775.220 -0.130 805.220 ;
        RECT -32.530 774.620 -0.130 775.220 ;
        RECT 3.170 805.220 35.570 805.820 ;
        RECT 3.170 775.220 4.970 805.220 ;
        RECT 34.970 775.220 35.570 805.220 ;
        RECT 3.170 774.620 35.570 775.220 ;
        RECT 42.470 805.220 74.870 805.820 ;
        RECT 42.470 775.220 43.070 805.220 ;
        RECT 73.070 775.220 74.870 805.220 ;
        RECT 42.470 774.620 74.870 775.220 ;
        RECT 78.170 805.220 110.570 805.820 ;
        RECT 78.170 775.220 79.970 805.220 ;
        RECT 109.970 775.220 110.570 805.220 ;
        RECT 78.170 774.620 110.570 775.220 ;
        RECT 117.470 805.220 149.870 805.820 ;
        RECT 117.470 775.220 118.070 805.220 ;
        RECT 148.070 775.220 149.870 805.220 ;
        RECT 117.470 774.620 149.870 775.220 ;
        RECT 153.170 805.220 185.570 805.820 ;
        RECT 153.170 775.220 154.970 805.220 ;
        RECT 184.970 775.220 185.570 805.220 ;
        RECT 153.170 774.620 185.570 775.220 ;
        RECT 192.470 805.220 224.870 805.820 ;
        RECT 192.470 775.220 193.070 805.220 ;
        RECT 223.070 775.220 224.870 805.220 ;
        RECT 192.470 774.620 224.870 775.220 ;
        RECT 228.170 805.220 260.570 805.820 ;
        RECT 228.170 775.220 229.970 805.220 ;
        RECT 259.970 775.220 260.570 805.220 ;
        RECT 228.170 774.620 260.570 775.220 ;
        RECT 267.470 805.220 299.870 805.820 ;
        RECT 267.470 775.220 268.070 805.220 ;
        RECT 298.070 775.220 299.870 805.220 ;
        RECT 267.470 774.620 299.870 775.220 ;
        RECT 303.170 805.220 335.570 805.820 ;
        RECT 303.170 775.220 304.970 805.220 ;
        RECT 334.970 775.220 335.570 805.220 ;
        RECT 303.170 774.620 335.570 775.220 ;
        RECT 342.470 805.220 374.870 805.820 ;
        RECT 342.470 775.220 343.070 805.220 ;
        RECT 373.070 775.220 374.870 805.220 ;
        RECT 342.470 774.620 374.870 775.220 ;
        RECT 378.170 805.220 410.570 805.820 ;
        RECT 378.170 775.220 379.970 805.220 ;
        RECT 409.970 775.220 410.570 805.220 ;
        RECT 378.170 774.620 410.570 775.220 ;
        RECT 417.470 805.220 449.870 805.820 ;
        RECT 417.470 775.220 418.070 805.220 ;
        RECT 448.070 775.220 449.870 805.220 ;
        RECT 417.470 774.620 449.870 775.220 ;
        RECT 453.170 805.220 485.570 805.820 ;
        RECT 453.170 775.220 454.970 805.220 ;
        RECT 484.970 775.220 485.570 805.220 ;
        RECT 453.170 774.620 485.570 775.220 ;
        RECT 492.470 805.220 524.870 805.820 ;
        RECT 492.470 775.220 493.070 805.220 ;
        RECT 523.070 775.220 524.870 805.220 ;
        RECT 492.470 774.620 524.870 775.220 ;
        RECT 528.170 805.220 560.570 805.820 ;
        RECT 528.170 775.220 529.970 805.220 ;
        RECT 559.970 775.220 560.570 805.220 ;
        RECT 528.170 774.620 560.570 775.220 ;
        RECT -557.530 770.220 -525.130 770.820 ;
        RECT -557.530 740.220 -556.930 770.220 ;
        RECT -526.930 740.220 -525.130 770.220 ;
        RECT -557.530 739.620 -525.130 740.220 ;
        RECT -521.830 770.220 -489.430 770.820 ;
        RECT -521.830 740.220 -520.030 770.220 ;
        RECT -490.030 740.220 -489.430 770.220 ;
        RECT -521.830 739.620 -489.430 740.220 ;
        RECT -482.530 770.220 -450.130 770.820 ;
        RECT -482.530 740.220 -481.930 770.220 ;
        RECT -451.930 740.220 -450.130 770.220 ;
        RECT -482.530 739.620 -450.130 740.220 ;
        RECT -446.830 770.220 -414.430 770.820 ;
        RECT -446.830 740.220 -445.030 770.220 ;
        RECT -415.030 740.220 -414.430 770.220 ;
        RECT -446.830 739.620 -414.430 740.220 ;
        RECT -407.530 770.220 -375.130 770.820 ;
        RECT -407.530 740.220 -406.930 770.220 ;
        RECT -376.930 740.220 -375.130 770.220 ;
        RECT -407.530 739.620 -375.130 740.220 ;
        RECT -371.830 770.220 -339.430 770.820 ;
        RECT -371.830 740.220 -370.030 770.220 ;
        RECT -340.030 740.220 -339.430 770.220 ;
        RECT -371.830 739.620 -339.430 740.220 ;
        RECT -332.530 770.220 -300.130 770.820 ;
        RECT -332.530 740.220 -331.930 770.220 ;
        RECT -301.930 740.220 -300.130 770.220 ;
        RECT -332.530 739.620 -300.130 740.220 ;
        RECT -296.830 770.220 -264.430 770.820 ;
        RECT -296.830 740.220 -295.030 770.220 ;
        RECT -265.030 740.220 -264.430 770.220 ;
        RECT -296.830 739.620 -264.430 740.220 ;
        RECT -257.530 770.220 -225.130 770.820 ;
        RECT -257.530 740.220 -256.930 770.220 ;
        RECT -226.930 740.220 -225.130 770.220 ;
        RECT -257.530 739.620 -225.130 740.220 ;
        RECT -221.830 770.220 -189.430 770.820 ;
        RECT -221.830 740.220 -220.030 770.220 ;
        RECT -190.030 740.220 -189.430 770.220 ;
        RECT -221.830 739.620 -189.430 740.220 ;
        RECT -182.530 770.220 -150.130 770.820 ;
        RECT -182.530 740.220 -181.930 770.220 ;
        RECT -151.930 740.220 -150.130 770.220 ;
        RECT -182.530 739.620 -150.130 740.220 ;
        RECT -146.830 770.220 -114.430 770.820 ;
        RECT -146.830 740.220 -145.030 770.220 ;
        RECT -115.030 740.220 -114.430 770.220 ;
        RECT -146.830 739.620 -114.430 740.220 ;
        RECT -107.530 770.220 -75.130 770.820 ;
        RECT -107.530 740.220 -106.930 770.220 ;
        RECT -76.930 740.220 -75.130 770.220 ;
        RECT -107.530 739.620 -75.130 740.220 ;
        RECT -71.830 770.220 -39.430 770.820 ;
        RECT -71.830 740.220 -70.030 770.220 ;
        RECT -40.030 740.220 -39.430 770.220 ;
        RECT -71.830 739.620 -39.430 740.220 ;
        RECT -32.530 770.220 -0.130 770.820 ;
        RECT -32.530 740.220 -31.930 770.220 ;
        RECT -1.930 740.220 -0.130 770.220 ;
        RECT -32.530 739.620 -0.130 740.220 ;
        RECT 3.170 770.220 35.570 770.820 ;
        RECT 3.170 740.220 4.970 770.220 ;
        RECT 34.970 740.220 35.570 770.220 ;
        RECT 3.170 739.620 35.570 740.220 ;
        RECT 42.470 770.220 74.870 770.820 ;
        RECT 42.470 740.220 43.070 770.220 ;
        RECT 73.070 740.220 74.870 770.220 ;
        RECT 42.470 739.620 74.870 740.220 ;
        RECT 78.170 770.220 110.570 770.820 ;
        RECT 78.170 740.220 79.970 770.220 ;
        RECT 109.970 740.220 110.570 770.220 ;
        RECT 78.170 739.620 110.570 740.220 ;
        RECT 117.470 770.220 149.870 770.820 ;
        RECT 117.470 740.220 118.070 770.220 ;
        RECT 148.070 740.220 149.870 770.220 ;
        RECT 117.470 739.620 149.870 740.220 ;
        RECT 153.170 770.220 185.570 770.820 ;
        RECT 153.170 740.220 154.970 770.220 ;
        RECT 184.970 740.220 185.570 770.220 ;
        RECT 153.170 739.620 185.570 740.220 ;
        RECT 192.470 770.220 224.870 770.820 ;
        RECT 192.470 740.220 193.070 770.220 ;
        RECT 223.070 740.220 224.870 770.220 ;
        RECT 192.470 739.620 224.870 740.220 ;
        RECT 228.170 770.220 260.570 770.820 ;
        RECT 228.170 740.220 229.970 770.220 ;
        RECT 259.970 740.220 260.570 770.220 ;
        RECT 228.170 739.620 260.570 740.220 ;
        RECT 267.470 770.220 299.870 770.820 ;
        RECT 267.470 740.220 268.070 770.220 ;
        RECT 298.070 740.220 299.870 770.220 ;
        RECT 267.470 739.620 299.870 740.220 ;
        RECT 303.170 770.220 335.570 770.820 ;
        RECT 303.170 740.220 304.970 770.220 ;
        RECT 334.970 740.220 335.570 770.220 ;
        RECT 303.170 739.620 335.570 740.220 ;
        RECT 342.470 770.220 374.870 770.820 ;
        RECT 342.470 740.220 343.070 770.220 ;
        RECT 373.070 740.220 374.870 770.220 ;
        RECT 342.470 739.620 374.870 740.220 ;
        RECT 378.170 770.220 410.570 770.820 ;
        RECT 378.170 740.220 379.970 770.220 ;
        RECT 409.970 740.220 410.570 770.220 ;
        RECT 378.170 739.620 410.570 740.220 ;
        RECT 417.470 770.220 449.870 770.820 ;
        RECT 417.470 740.220 418.070 770.220 ;
        RECT 448.070 740.220 449.870 770.220 ;
        RECT 417.470 739.620 449.870 740.220 ;
        RECT 453.170 770.220 485.570 770.820 ;
        RECT 453.170 740.220 454.970 770.220 ;
        RECT 484.970 740.220 485.570 770.220 ;
        RECT 453.170 739.620 485.570 740.220 ;
        RECT 492.470 770.220 524.870 770.820 ;
        RECT 492.470 740.220 493.070 770.220 ;
        RECT 523.070 740.220 524.870 770.220 ;
        RECT 492.470 739.620 524.870 740.220 ;
        RECT 528.170 770.220 560.570 770.820 ;
        RECT 528.170 740.220 529.970 770.220 ;
        RECT 559.970 740.220 560.570 770.220 ;
        RECT 528.170 739.620 560.570 740.220 ;
        RECT -557.530 735.220 -525.130 735.820 ;
        RECT -557.530 705.220 -556.930 735.220 ;
        RECT -526.930 705.220 -525.130 735.220 ;
        RECT -557.530 704.620 -525.130 705.220 ;
        RECT -521.830 735.220 -489.430 735.820 ;
        RECT -521.830 705.220 -520.030 735.220 ;
        RECT -490.030 705.220 -489.430 735.220 ;
        RECT -521.830 704.620 -489.430 705.220 ;
        RECT -482.530 735.220 -450.130 735.820 ;
        RECT -482.530 705.220 -481.930 735.220 ;
        RECT -451.930 705.220 -450.130 735.220 ;
        RECT -482.530 704.620 -450.130 705.220 ;
        RECT -446.830 735.220 -414.430 735.820 ;
        RECT -446.830 705.220 -445.030 735.220 ;
        RECT -415.030 705.220 -414.430 735.220 ;
        RECT -446.830 704.620 -414.430 705.220 ;
        RECT -407.530 735.220 -375.130 735.820 ;
        RECT -407.530 705.220 -406.930 735.220 ;
        RECT -376.930 705.220 -375.130 735.220 ;
        RECT -407.530 704.620 -375.130 705.220 ;
        RECT -371.830 735.220 -339.430 735.820 ;
        RECT -371.830 705.220 -370.030 735.220 ;
        RECT -340.030 705.220 -339.430 735.220 ;
        RECT -371.830 704.620 -339.430 705.220 ;
        RECT -332.530 735.220 -300.130 735.820 ;
        RECT -332.530 705.220 -331.930 735.220 ;
        RECT -301.930 705.220 -300.130 735.220 ;
        RECT -332.530 704.620 -300.130 705.220 ;
        RECT -296.830 735.220 -264.430 735.820 ;
        RECT -296.830 705.220 -295.030 735.220 ;
        RECT -265.030 705.220 -264.430 735.220 ;
        RECT -296.830 704.620 -264.430 705.220 ;
        RECT -257.530 735.220 -225.130 735.820 ;
        RECT -257.530 705.220 -256.930 735.220 ;
        RECT -226.930 705.220 -225.130 735.220 ;
        RECT -257.530 704.620 -225.130 705.220 ;
        RECT -221.830 735.220 -189.430 735.820 ;
        RECT -221.830 705.220 -220.030 735.220 ;
        RECT -190.030 705.220 -189.430 735.220 ;
        RECT -221.830 704.620 -189.430 705.220 ;
        RECT -182.530 735.220 -150.130 735.820 ;
        RECT -182.530 705.220 -181.930 735.220 ;
        RECT -151.930 705.220 -150.130 735.220 ;
        RECT -182.530 704.620 -150.130 705.220 ;
        RECT -146.830 735.220 -114.430 735.820 ;
        RECT -146.830 705.220 -145.030 735.220 ;
        RECT -115.030 705.220 -114.430 735.220 ;
        RECT -146.830 704.620 -114.430 705.220 ;
        RECT -107.530 735.220 -75.130 735.820 ;
        RECT -107.530 705.220 -106.930 735.220 ;
        RECT -76.930 705.220 -75.130 735.220 ;
        RECT -107.530 704.620 -75.130 705.220 ;
        RECT -71.830 735.220 -39.430 735.820 ;
        RECT -71.830 705.220 -70.030 735.220 ;
        RECT -40.030 705.220 -39.430 735.220 ;
        RECT -71.830 704.620 -39.430 705.220 ;
        RECT -32.530 735.220 -0.130 735.820 ;
        RECT -32.530 705.220 -31.930 735.220 ;
        RECT -1.930 705.220 -0.130 735.220 ;
        RECT -32.530 704.620 -0.130 705.220 ;
        RECT 3.170 735.220 35.570 735.820 ;
        RECT 3.170 705.220 4.970 735.220 ;
        RECT 34.970 705.220 35.570 735.220 ;
        RECT 3.170 704.620 35.570 705.220 ;
        RECT 42.470 735.220 74.870 735.820 ;
        RECT 42.470 705.220 43.070 735.220 ;
        RECT 73.070 705.220 74.870 735.220 ;
        RECT 42.470 704.620 74.870 705.220 ;
        RECT 78.170 735.220 110.570 735.820 ;
        RECT 78.170 705.220 79.970 735.220 ;
        RECT 109.970 705.220 110.570 735.220 ;
        RECT 78.170 704.620 110.570 705.220 ;
        RECT 117.470 735.220 149.870 735.820 ;
        RECT 117.470 705.220 118.070 735.220 ;
        RECT 148.070 705.220 149.870 735.220 ;
        RECT 117.470 704.620 149.870 705.220 ;
        RECT 153.170 735.220 185.570 735.820 ;
        RECT 153.170 705.220 154.970 735.220 ;
        RECT 184.970 705.220 185.570 735.220 ;
        RECT 153.170 704.620 185.570 705.220 ;
        RECT 192.470 735.220 224.870 735.820 ;
        RECT 192.470 705.220 193.070 735.220 ;
        RECT 223.070 705.220 224.870 735.220 ;
        RECT 192.470 704.620 224.870 705.220 ;
        RECT 228.170 735.220 260.570 735.820 ;
        RECT 228.170 705.220 229.970 735.220 ;
        RECT 259.970 705.220 260.570 735.220 ;
        RECT 228.170 704.620 260.570 705.220 ;
        RECT 267.470 735.220 299.870 735.820 ;
        RECT 267.470 705.220 268.070 735.220 ;
        RECT 298.070 705.220 299.870 735.220 ;
        RECT 267.470 704.620 299.870 705.220 ;
        RECT 303.170 735.220 335.570 735.820 ;
        RECT 303.170 705.220 304.970 735.220 ;
        RECT 334.970 705.220 335.570 735.220 ;
        RECT 303.170 704.620 335.570 705.220 ;
        RECT 342.470 735.220 374.870 735.820 ;
        RECT 342.470 705.220 343.070 735.220 ;
        RECT 373.070 705.220 374.870 735.220 ;
        RECT 342.470 704.620 374.870 705.220 ;
        RECT 378.170 735.220 410.570 735.820 ;
        RECT 378.170 705.220 379.970 735.220 ;
        RECT 409.970 705.220 410.570 735.220 ;
        RECT 378.170 704.620 410.570 705.220 ;
        RECT 417.470 735.220 449.870 735.820 ;
        RECT 417.470 705.220 418.070 735.220 ;
        RECT 448.070 705.220 449.870 735.220 ;
        RECT 417.470 704.620 449.870 705.220 ;
        RECT 453.170 735.220 485.570 735.820 ;
        RECT 453.170 705.220 454.970 735.220 ;
        RECT 484.970 705.220 485.570 735.220 ;
        RECT 453.170 704.620 485.570 705.220 ;
        RECT 492.470 735.220 524.870 735.820 ;
        RECT 492.470 705.220 493.070 735.220 ;
        RECT 523.070 705.220 524.870 735.220 ;
        RECT 492.470 704.620 524.870 705.220 ;
        RECT 528.170 735.220 560.570 735.820 ;
        RECT 528.170 705.220 529.970 735.220 ;
        RECT 559.970 705.220 560.570 735.220 ;
        RECT 528.170 704.620 560.570 705.220 ;
        RECT -557.530 700.220 -525.130 700.820 ;
        RECT -557.530 670.220 -556.930 700.220 ;
        RECT -526.930 670.220 -525.130 700.220 ;
        RECT -557.530 669.620 -525.130 670.220 ;
        RECT -521.830 700.220 -489.430 700.820 ;
        RECT -521.830 670.220 -520.030 700.220 ;
        RECT -490.030 670.220 -489.430 700.220 ;
        RECT -521.830 669.620 -489.430 670.220 ;
        RECT -482.530 700.220 -450.130 700.820 ;
        RECT -482.530 670.220 -481.930 700.220 ;
        RECT -451.930 670.220 -450.130 700.220 ;
        RECT -482.530 669.620 -450.130 670.220 ;
        RECT -446.830 700.220 -414.430 700.820 ;
        RECT -446.830 670.220 -445.030 700.220 ;
        RECT -415.030 670.220 -414.430 700.220 ;
        RECT -446.830 669.620 -414.430 670.220 ;
        RECT -407.530 700.220 -375.130 700.820 ;
        RECT -407.530 670.220 -406.930 700.220 ;
        RECT -376.930 670.220 -375.130 700.220 ;
        RECT -407.530 669.620 -375.130 670.220 ;
        RECT -371.830 700.220 -339.430 700.820 ;
        RECT -371.830 670.220 -370.030 700.220 ;
        RECT -340.030 670.220 -339.430 700.220 ;
        RECT -371.830 669.620 -339.430 670.220 ;
        RECT -332.530 700.220 -300.130 700.820 ;
        RECT -332.530 670.220 -331.930 700.220 ;
        RECT -301.930 670.220 -300.130 700.220 ;
        RECT -332.530 669.620 -300.130 670.220 ;
        RECT -296.830 700.220 -264.430 700.820 ;
        RECT -296.830 670.220 -295.030 700.220 ;
        RECT -265.030 670.220 -264.430 700.220 ;
        RECT -296.830 669.620 -264.430 670.220 ;
        RECT -257.530 700.220 -225.130 700.820 ;
        RECT -257.530 670.220 -256.930 700.220 ;
        RECT -226.930 670.220 -225.130 700.220 ;
        RECT -257.530 669.620 -225.130 670.220 ;
        RECT -221.830 700.220 -189.430 700.820 ;
        RECT -221.830 670.220 -220.030 700.220 ;
        RECT -190.030 670.220 -189.430 700.220 ;
        RECT -221.830 669.620 -189.430 670.220 ;
        RECT -182.530 700.220 -150.130 700.820 ;
        RECT -182.530 670.220 -181.930 700.220 ;
        RECT -151.930 670.220 -150.130 700.220 ;
        RECT -182.530 669.620 -150.130 670.220 ;
        RECT -146.830 700.220 -114.430 700.820 ;
        RECT -146.830 670.220 -145.030 700.220 ;
        RECT -115.030 670.220 -114.430 700.220 ;
        RECT -146.830 669.620 -114.430 670.220 ;
        RECT -107.530 700.220 -75.130 700.820 ;
        RECT -107.530 670.220 -106.930 700.220 ;
        RECT -76.930 670.220 -75.130 700.220 ;
        RECT -107.530 669.620 -75.130 670.220 ;
        RECT -71.830 700.220 -39.430 700.820 ;
        RECT -71.830 670.220 -70.030 700.220 ;
        RECT -40.030 670.220 -39.430 700.220 ;
        RECT -71.830 669.620 -39.430 670.220 ;
        RECT -32.530 700.220 -0.130 700.820 ;
        RECT -32.530 670.220 -31.930 700.220 ;
        RECT -1.930 670.220 -0.130 700.220 ;
        RECT -32.530 669.620 -0.130 670.220 ;
        RECT 3.170 700.220 35.570 700.820 ;
        RECT 3.170 670.220 4.970 700.220 ;
        RECT 34.970 670.220 35.570 700.220 ;
        RECT 3.170 669.620 35.570 670.220 ;
        RECT 42.470 700.220 74.870 700.820 ;
        RECT 42.470 670.220 43.070 700.220 ;
        RECT 73.070 670.220 74.870 700.220 ;
        RECT 42.470 669.620 74.870 670.220 ;
        RECT 78.170 700.220 110.570 700.820 ;
        RECT 78.170 670.220 79.970 700.220 ;
        RECT 109.970 670.220 110.570 700.220 ;
        RECT 78.170 669.620 110.570 670.220 ;
        RECT 117.470 700.220 149.870 700.820 ;
        RECT 117.470 670.220 118.070 700.220 ;
        RECT 148.070 670.220 149.870 700.220 ;
        RECT 117.470 669.620 149.870 670.220 ;
        RECT 153.170 700.220 185.570 700.820 ;
        RECT 153.170 670.220 154.970 700.220 ;
        RECT 184.970 670.220 185.570 700.220 ;
        RECT 153.170 669.620 185.570 670.220 ;
        RECT 192.470 700.220 224.870 700.820 ;
        RECT 192.470 670.220 193.070 700.220 ;
        RECT 223.070 670.220 224.870 700.220 ;
        RECT 192.470 669.620 224.870 670.220 ;
        RECT 228.170 700.220 260.570 700.820 ;
        RECT 228.170 670.220 229.970 700.220 ;
        RECT 259.970 670.220 260.570 700.220 ;
        RECT 228.170 669.620 260.570 670.220 ;
        RECT 267.470 700.220 299.870 700.820 ;
        RECT 267.470 670.220 268.070 700.220 ;
        RECT 298.070 670.220 299.870 700.220 ;
        RECT 267.470 669.620 299.870 670.220 ;
        RECT 303.170 700.220 335.570 700.820 ;
        RECT 303.170 670.220 304.970 700.220 ;
        RECT 334.970 670.220 335.570 700.220 ;
        RECT 303.170 669.620 335.570 670.220 ;
        RECT 342.470 700.220 374.870 700.820 ;
        RECT 342.470 670.220 343.070 700.220 ;
        RECT 373.070 670.220 374.870 700.220 ;
        RECT 342.470 669.620 374.870 670.220 ;
        RECT 378.170 700.220 410.570 700.820 ;
        RECT 378.170 670.220 379.970 700.220 ;
        RECT 409.970 670.220 410.570 700.220 ;
        RECT 378.170 669.620 410.570 670.220 ;
        RECT 417.470 700.220 449.870 700.820 ;
        RECT 417.470 670.220 418.070 700.220 ;
        RECT 448.070 670.220 449.870 700.220 ;
        RECT 417.470 669.620 449.870 670.220 ;
        RECT 453.170 700.220 485.570 700.820 ;
        RECT 453.170 670.220 454.970 700.220 ;
        RECT 484.970 670.220 485.570 700.220 ;
        RECT 453.170 669.620 485.570 670.220 ;
        RECT 492.470 700.220 524.870 700.820 ;
        RECT 492.470 670.220 493.070 700.220 ;
        RECT 523.070 670.220 524.870 700.220 ;
        RECT 492.470 669.620 524.870 670.220 ;
        RECT 528.170 700.220 560.570 700.820 ;
        RECT 528.170 670.220 529.970 700.220 ;
        RECT 559.970 670.220 560.570 700.220 ;
        RECT 528.170 669.620 560.570 670.220 ;
        RECT -557.530 665.220 -525.130 665.820 ;
        RECT -557.530 635.220 -556.930 665.220 ;
        RECT -526.930 635.220 -525.130 665.220 ;
        RECT -557.530 634.620 -525.130 635.220 ;
        RECT -521.830 665.220 -489.430 665.820 ;
        RECT -521.830 635.220 -520.030 665.220 ;
        RECT -490.030 635.220 -489.430 665.220 ;
        RECT -521.830 634.620 -489.430 635.220 ;
        RECT -482.530 665.220 -450.130 665.820 ;
        RECT -482.530 635.220 -481.930 665.220 ;
        RECT -451.930 635.220 -450.130 665.220 ;
        RECT -482.530 634.620 -450.130 635.220 ;
        RECT -446.830 665.220 -414.430 665.820 ;
        RECT -446.830 635.220 -445.030 665.220 ;
        RECT -415.030 635.220 -414.430 665.220 ;
        RECT -446.830 634.620 -414.430 635.220 ;
        RECT -407.530 665.220 -375.130 665.820 ;
        RECT -407.530 635.220 -406.930 665.220 ;
        RECT -376.930 635.220 -375.130 665.220 ;
        RECT -407.530 634.620 -375.130 635.220 ;
        RECT -371.830 665.220 -339.430 665.820 ;
        RECT -371.830 635.220 -370.030 665.220 ;
        RECT -340.030 635.220 -339.430 665.220 ;
        RECT -371.830 634.620 -339.430 635.220 ;
        RECT -332.530 665.220 -300.130 665.820 ;
        RECT -332.530 635.220 -331.930 665.220 ;
        RECT -301.930 635.220 -300.130 665.220 ;
        RECT -332.530 634.620 -300.130 635.220 ;
        RECT -296.830 665.220 -264.430 665.820 ;
        RECT -296.830 635.220 -295.030 665.220 ;
        RECT -265.030 635.220 -264.430 665.220 ;
        RECT -296.830 634.620 -264.430 635.220 ;
        RECT -257.530 665.220 -225.130 665.820 ;
        RECT -257.530 635.220 -256.930 665.220 ;
        RECT -226.930 635.220 -225.130 665.220 ;
        RECT -257.530 634.620 -225.130 635.220 ;
        RECT -221.830 665.220 -189.430 665.820 ;
        RECT -221.830 635.220 -220.030 665.220 ;
        RECT -190.030 635.220 -189.430 665.220 ;
        RECT -221.830 634.620 -189.430 635.220 ;
        RECT -182.530 665.220 -150.130 665.820 ;
        RECT -182.530 635.220 -181.930 665.220 ;
        RECT -151.930 635.220 -150.130 665.220 ;
        RECT -182.530 634.620 -150.130 635.220 ;
        RECT -146.830 665.220 -114.430 665.820 ;
        RECT -146.830 635.220 -145.030 665.220 ;
        RECT -115.030 635.220 -114.430 665.220 ;
        RECT -146.830 634.620 -114.430 635.220 ;
        RECT -107.530 665.220 -75.130 665.820 ;
        RECT -107.530 635.220 -106.930 665.220 ;
        RECT -76.930 635.220 -75.130 665.220 ;
        RECT -107.530 634.620 -75.130 635.220 ;
        RECT -71.830 665.220 -39.430 665.820 ;
        RECT -71.830 635.220 -70.030 665.220 ;
        RECT -40.030 635.220 -39.430 665.220 ;
        RECT -71.830 634.620 -39.430 635.220 ;
        RECT -32.530 665.220 -0.130 665.820 ;
        RECT -32.530 635.220 -31.930 665.220 ;
        RECT -1.930 635.220 -0.130 665.220 ;
        RECT -32.530 634.620 -0.130 635.220 ;
        RECT 3.170 665.220 35.570 665.820 ;
        RECT 3.170 635.220 4.970 665.220 ;
        RECT 34.970 635.220 35.570 665.220 ;
        RECT 3.170 634.620 35.570 635.220 ;
        RECT 42.470 665.220 74.870 665.820 ;
        RECT 42.470 635.220 43.070 665.220 ;
        RECT 73.070 635.220 74.870 665.220 ;
        RECT 42.470 634.620 74.870 635.220 ;
        RECT 78.170 665.220 110.570 665.820 ;
        RECT 78.170 635.220 79.970 665.220 ;
        RECT 109.970 635.220 110.570 665.220 ;
        RECT 78.170 634.620 110.570 635.220 ;
        RECT 117.470 665.220 149.870 665.820 ;
        RECT 117.470 635.220 118.070 665.220 ;
        RECT 148.070 635.220 149.870 665.220 ;
        RECT 117.470 634.620 149.870 635.220 ;
        RECT 153.170 665.220 185.570 665.820 ;
        RECT 153.170 635.220 154.970 665.220 ;
        RECT 184.970 635.220 185.570 665.220 ;
        RECT 153.170 634.620 185.570 635.220 ;
        RECT 192.470 665.220 224.870 665.820 ;
        RECT 192.470 635.220 193.070 665.220 ;
        RECT 223.070 635.220 224.870 665.220 ;
        RECT 192.470 634.620 224.870 635.220 ;
        RECT 228.170 665.220 260.570 665.820 ;
        RECT 228.170 635.220 229.970 665.220 ;
        RECT 259.970 635.220 260.570 665.220 ;
        RECT 228.170 634.620 260.570 635.220 ;
        RECT 267.470 665.220 299.870 665.820 ;
        RECT 267.470 635.220 268.070 665.220 ;
        RECT 298.070 635.220 299.870 665.220 ;
        RECT 267.470 634.620 299.870 635.220 ;
        RECT 303.170 665.220 335.570 665.820 ;
        RECT 303.170 635.220 304.970 665.220 ;
        RECT 334.970 635.220 335.570 665.220 ;
        RECT 303.170 634.620 335.570 635.220 ;
        RECT 342.470 665.220 374.870 665.820 ;
        RECT 342.470 635.220 343.070 665.220 ;
        RECT 373.070 635.220 374.870 665.220 ;
        RECT 342.470 634.620 374.870 635.220 ;
        RECT 378.170 665.220 410.570 665.820 ;
        RECT 378.170 635.220 379.970 665.220 ;
        RECT 409.970 635.220 410.570 665.220 ;
        RECT 378.170 634.620 410.570 635.220 ;
        RECT 417.470 665.220 449.870 665.820 ;
        RECT 417.470 635.220 418.070 665.220 ;
        RECT 448.070 635.220 449.870 665.220 ;
        RECT 417.470 634.620 449.870 635.220 ;
        RECT 453.170 665.220 485.570 665.820 ;
        RECT 453.170 635.220 454.970 665.220 ;
        RECT 484.970 635.220 485.570 665.220 ;
        RECT 453.170 634.620 485.570 635.220 ;
        RECT 492.470 665.220 524.870 665.820 ;
        RECT 492.470 635.220 493.070 665.220 ;
        RECT 523.070 635.220 524.870 665.220 ;
        RECT 492.470 634.620 524.870 635.220 ;
        RECT 528.170 665.220 560.570 665.820 ;
        RECT 528.170 635.220 529.970 665.220 ;
        RECT 559.970 635.220 560.570 665.220 ;
        RECT 528.170 634.620 560.570 635.220 ;
        RECT -557.530 630.220 -525.130 630.820 ;
        RECT -557.530 600.220 -556.930 630.220 ;
        RECT -526.930 600.220 -525.130 630.220 ;
        RECT -557.530 599.620 -525.130 600.220 ;
        RECT -521.830 630.220 -489.430 630.820 ;
        RECT -521.830 600.220 -520.030 630.220 ;
        RECT -490.030 600.220 -489.430 630.220 ;
        RECT -521.830 599.620 -489.430 600.220 ;
        RECT -482.530 630.220 -450.130 630.820 ;
        RECT -482.530 600.220 -481.930 630.220 ;
        RECT -451.930 600.220 -450.130 630.220 ;
        RECT -482.530 599.620 -450.130 600.220 ;
        RECT -446.830 630.220 -414.430 630.820 ;
        RECT -446.830 600.220 -445.030 630.220 ;
        RECT -415.030 600.220 -414.430 630.220 ;
        RECT -446.830 599.620 -414.430 600.220 ;
        RECT -407.530 630.220 -375.130 630.820 ;
        RECT -407.530 600.220 -406.930 630.220 ;
        RECT -376.930 600.220 -375.130 630.220 ;
        RECT -407.530 599.620 -375.130 600.220 ;
        RECT -371.830 630.220 -339.430 630.820 ;
        RECT -371.830 600.220 -370.030 630.220 ;
        RECT -340.030 600.220 -339.430 630.220 ;
        RECT -371.830 599.620 -339.430 600.220 ;
        RECT -332.530 630.220 -300.130 630.820 ;
        RECT -332.530 600.220 -331.930 630.220 ;
        RECT -301.930 600.220 -300.130 630.220 ;
        RECT -332.530 599.620 -300.130 600.220 ;
        RECT -296.830 630.220 -264.430 630.820 ;
        RECT -296.830 600.220 -295.030 630.220 ;
        RECT -265.030 600.220 -264.430 630.220 ;
        RECT -296.830 599.620 -264.430 600.220 ;
        RECT -257.530 630.220 -225.130 630.820 ;
        RECT -257.530 600.220 -256.930 630.220 ;
        RECT -226.930 600.220 -225.130 630.220 ;
        RECT -257.530 599.620 -225.130 600.220 ;
        RECT -221.830 630.220 -189.430 630.820 ;
        RECT -221.830 600.220 -220.030 630.220 ;
        RECT -190.030 600.220 -189.430 630.220 ;
        RECT -221.830 599.620 -189.430 600.220 ;
        RECT -182.530 630.220 -150.130 630.820 ;
        RECT -182.530 600.220 -181.930 630.220 ;
        RECT -151.930 600.220 -150.130 630.220 ;
        RECT -182.530 599.620 -150.130 600.220 ;
        RECT -146.830 630.220 -114.430 630.820 ;
        RECT -146.830 600.220 -145.030 630.220 ;
        RECT -115.030 600.220 -114.430 630.220 ;
        RECT -146.830 599.620 -114.430 600.220 ;
        RECT -107.530 630.220 -75.130 630.820 ;
        RECT -107.530 600.220 -106.930 630.220 ;
        RECT -76.930 600.220 -75.130 630.220 ;
        RECT -107.530 599.620 -75.130 600.220 ;
        RECT -71.830 630.220 -39.430 630.820 ;
        RECT -71.830 600.220 -70.030 630.220 ;
        RECT -40.030 600.220 -39.430 630.220 ;
        RECT -71.830 599.620 -39.430 600.220 ;
        RECT -32.530 630.220 -0.130 630.820 ;
        RECT -32.530 600.220 -31.930 630.220 ;
        RECT -1.930 600.220 -0.130 630.220 ;
        RECT -32.530 599.620 -0.130 600.220 ;
        RECT 3.170 630.220 35.570 630.820 ;
        RECT 3.170 600.220 4.970 630.220 ;
        RECT 34.970 600.220 35.570 630.220 ;
        RECT 3.170 599.620 35.570 600.220 ;
        RECT 42.470 630.220 74.870 630.820 ;
        RECT 42.470 600.220 43.070 630.220 ;
        RECT 73.070 600.220 74.870 630.220 ;
        RECT 42.470 599.620 74.870 600.220 ;
        RECT 78.170 630.220 110.570 630.820 ;
        RECT 78.170 600.220 79.970 630.220 ;
        RECT 109.970 600.220 110.570 630.220 ;
        RECT 78.170 599.620 110.570 600.220 ;
        RECT 117.470 630.220 149.870 630.820 ;
        RECT 117.470 600.220 118.070 630.220 ;
        RECT 148.070 600.220 149.870 630.220 ;
        RECT 117.470 599.620 149.870 600.220 ;
        RECT 153.170 630.220 185.570 630.820 ;
        RECT 153.170 600.220 154.970 630.220 ;
        RECT 184.970 600.220 185.570 630.220 ;
        RECT 153.170 599.620 185.570 600.220 ;
        RECT 192.470 630.220 224.870 630.820 ;
        RECT 192.470 600.220 193.070 630.220 ;
        RECT 223.070 600.220 224.870 630.220 ;
        RECT 192.470 599.620 224.870 600.220 ;
        RECT 228.170 630.220 260.570 630.820 ;
        RECT 228.170 600.220 229.970 630.220 ;
        RECT 259.970 600.220 260.570 630.220 ;
        RECT 228.170 599.620 260.570 600.220 ;
        RECT 267.470 630.220 299.870 630.820 ;
        RECT 267.470 600.220 268.070 630.220 ;
        RECT 298.070 600.220 299.870 630.220 ;
        RECT 267.470 599.620 299.870 600.220 ;
        RECT 303.170 630.220 335.570 630.820 ;
        RECT 303.170 600.220 304.970 630.220 ;
        RECT 334.970 600.220 335.570 630.220 ;
        RECT 303.170 599.620 335.570 600.220 ;
        RECT 342.470 630.220 374.870 630.820 ;
        RECT 342.470 600.220 343.070 630.220 ;
        RECT 373.070 600.220 374.870 630.220 ;
        RECT 342.470 599.620 374.870 600.220 ;
        RECT 378.170 630.220 410.570 630.820 ;
        RECT 378.170 600.220 379.970 630.220 ;
        RECT 409.970 600.220 410.570 630.220 ;
        RECT 378.170 599.620 410.570 600.220 ;
        RECT 417.470 630.220 449.870 630.820 ;
        RECT 417.470 600.220 418.070 630.220 ;
        RECT 448.070 600.220 449.870 630.220 ;
        RECT 417.470 599.620 449.870 600.220 ;
        RECT 453.170 630.220 485.570 630.820 ;
        RECT 453.170 600.220 454.970 630.220 ;
        RECT 484.970 600.220 485.570 630.220 ;
        RECT 453.170 599.620 485.570 600.220 ;
        RECT 492.470 630.220 524.870 630.820 ;
        RECT 492.470 600.220 493.070 630.220 ;
        RECT 523.070 600.220 524.870 630.220 ;
        RECT 492.470 599.620 524.870 600.220 ;
        RECT 528.170 630.220 560.570 630.820 ;
        RECT 528.170 600.220 529.970 630.220 ;
        RECT 559.970 600.220 560.570 630.220 ;
        RECT 528.170 599.620 560.570 600.220 ;
        RECT -557.530 595.220 -525.130 595.820 ;
        RECT -557.530 565.220 -556.930 595.220 ;
        RECT -526.930 565.220 -525.130 595.220 ;
        RECT -557.530 564.620 -525.130 565.220 ;
        RECT -521.830 595.220 -489.430 595.820 ;
        RECT -521.830 565.220 -520.030 595.220 ;
        RECT -490.030 565.220 -489.430 595.220 ;
        RECT -521.830 564.620 -489.430 565.220 ;
        RECT -482.530 595.220 -450.130 595.820 ;
        RECT -482.530 565.220 -481.930 595.220 ;
        RECT -451.930 565.220 -450.130 595.220 ;
        RECT -482.530 564.620 -450.130 565.220 ;
        RECT -446.830 595.220 -414.430 595.820 ;
        RECT -446.830 565.220 -445.030 595.220 ;
        RECT -415.030 565.220 -414.430 595.220 ;
        RECT -446.830 564.620 -414.430 565.220 ;
        RECT -407.530 595.220 -375.130 595.820 ;
        RECT -407.530 565.220 -406.930 595.220 ;
        RECT -376.930 565.220 -375.130 595.220 ;
        RECT -407.530 564.620 -375.130 565.220 ;
        RECT -371.830 595.220 -339.430 595.820 ;
        RECT -371.830 565.220 -370.030 595.220 ;
        RECT -340.030 565.220 -339.430 595.220 ;
        RECT -371.830 564.620 -339.430 565.220 ;
        RECT -332.530 595.220 -300.130 595.820 ;
        RECT -332.530 565.220 -331.930 595.220 ;
        RECT -301.930 565.220 -300.130 595.220 ;
        RECT -332.530 564.620 -300.130 565.220 ;
        RECT -296.830 595.220 -264.430 595.820 ;
        RECT -296.830 565.220 -295.030 595.220 ;
        RECT -265.030 565.220 -264.430 595.220 ;
        RECT -296.830 564.620 -264.430 565.220 ;
        RECT -257.530 595.220 -225.130 595.820 ;
        RECT -257.530 565.220 -256.930 595.220 ;
        RECT -226.930 565.220 -225.130 595.220 ;
        RECT -257.530 564.620 -225.130 565.220 ;
        RECT -221.830 595.220 -189.430 595.820 ;
        RECT -221.830 565.220 -220.030 595.220 ;
        RECT -190.030 565.220 -189.430 595.220 ;
        RECT -221.830 564.620 -189.430 565.220 ;
        RECT -182.530 595.220 -150.130 595.820 ;
        RECT -182.530 565.220 -181.930 595.220 ;
        RECT -151.930 565.220 -150.130 595.220 ;
        RECT -182.530 564.620 -150.130 565.220 ;
        RECT -146.830 595.220 -114.430 595.820 ;
        RECT -146.830 565.220 -145.030 595.220 ;
        RECT -115.030 565.220 -114.430 595.220 ;
        RECT -146.830 564.620 -114.430 565.220 ;
        RECT -107.530 595.220 -75.130 595.820 ;
        RECT -107.530 565.220 -106.930 595.220 ;
        RECT -76.930 565.220 -75.130 595.220 ;
        RECT -107.530 564.620 -75.130 565.220 ;
        RECT -71.830 595.220 -39.430 595.820 ;
        RECT -71.830 565.220 -70.030 595.220 ;
        RECT -40.030 565.220 -39.430 595.220 ;
        RECT -71.830 564.620 -39.430 565.220 ;
        RECT -32.530 595.220 -0.130 595.820 ;
        RECT -32.530 565.220 -31.930 595.220 ;
        RECT -1.930 565.220 -0.130 595.220 ;
        RECT -32.530 564.620 -0.130 565.220 ;
        RECT 3.170 595.220 35.570 595.820 ;
        RECT 3.170 565.220 4.970 595.220 ;
        RECT 34.970 565.220 35.570 595.220 ;
        RECT 3.170 564.620 35.570 565.220 ;
        RECT 42.470 595.220 74.870 595.820 ;
        RECT 42.470 565.220 43.070 595.220 ;
        RECT 73.070 565.220 74.870 595.220 ;
        RECT 42.470 564.620 74.870 565.220 ;
        RECT 78.170 595.220 110.570 595.820 ;
        RECT 78.170 565.220 79.970 595.220 ;
        RECT 109.970 565.220 110.570 595.220 ;
        RECT 78.170 564.620 110.570 565.220 ;
        RECT 117.470 595.220 149.870 595.820 ;
        RECT 117.470 565.220 118.070 595.220 ;
        RECT 148.070 565.220 149.870 595.220 ;
        RECT 117.470 564.620 149.870 565.220 ;
        RECT 153.170 595.220 185.570 595.820 ;
        RECT 153.170 565.220 154.970 595.220 ;
        RECT 184.970 565.220 185.570 595.220 ;
        RECT 153.170 564.620 185.570 565.220 ;
        RECT 192.470 595.220 224.870 595.820 ;
        RECT 192.470 565.220 193.070 595.220 ;
        RECT 223.070 565.220 224.870 595.220 ;
        RECT 192.470 564.620 224.870 565.220 ;
        RECT 228.170 595.220 260.570 595.820 ;
        RECT 228.170 565.220 229.970 595.220 ;
        RECT 259.970 565.220 260.570 595.220 ;
        RECT 228.170 564.620 260.570 565.220 ;
        RECT 267.470 595.220 299.870 595.820 ;
        RECT 267.470 565.220 268.070 595.220 ;
        RECT 298.070 565.220 299.870 595.220 ;
        RECT 267.470 564.620 299.870 565.220 ;
        RECT 303.170 595.220 335.570 595.820 ;
        RECT 303.170 565.220 304.970 595.220 ;
        RECT 334.970 565.220 335.570 595.220 ;
        RECT 303.170 564.620 335.570 565.220 ;
        RECT 342.470 595.220 374.870 595.820 ;
        RECT 342.470 565.220 343.070 595.220 ;
        RECT 373.070 565.220 374.870 595.220 ;
        RECT 342.470 564.620 374.870 565.220 ;
        RECT 378.170 595.220 410.570 595.820 ;
        RECT 378.170 565.220 379.970 595.220 ;
        RECT 409.970 565.220 410.570 595.220 ;
        RECT 378.170 564.620 410.570 565.220 ;
        RECT 417.470 595.220 449.870 595.820 ;
        RECT 417.470 565.220 418.070 595.220 ;
        RECT 448.070 565.220 449.870 595.220 ;
        RECT 417.470 564.620 449.870 565.220 ;
        RECT 453.170 595.220 485.570 595.820 ;
        RECT 453.170 565.220 454.970 595.220 ;
        RECT 484.970 565.220 485.570 595.220 ;
        RECT 453.170 564.620 485.570 565.220 ;
        RECT 492.470 595.220 524.870 595.820 ;
        RECT 492.470 565.220 493.070 595.220 ;
        RECT 523.070 565.220 524.870 595.220 ;
        RECT 492.470 564.620 524.870 565.220 ;
        RECT 528.170 595.220 560.570 595.820 ;
        RECT 528.170 565.220 529.970 595.220 ;
        RECT 559.970 565.220 560.570 595.220 ;
        RECT 528.170 564.620 560.570 565.220 ;
        RECT -557.530 560.220 -525.130 560.820 ;
        RECT -557.530 530.220 -556.930 560.220 ;
        RECT -526.930 530.220 -525.130 560.220 ;
        RECT -557.530 529.620 -525.130 530.220 ;
        RECT -521.830 560.220 -489.430 560.820 ;
        RECT -521.830 530.220 -520.030 560.220 ;
        RECT -490.030 530.220 -489.430 560.220 ;
        RECT -521.830 529.620 -489.430 530.220 ;
        RECT -482.530 560.220 -450.130 560.820 ;
        RECT -482.530 530.220 -481.930 560.220 ;
        RECT -451.930 530.220 -450.130 560.220 ;
        RECT -482.530 529.620 -450.130 530.220 ;
        RECT -446.830 560.220 -414.430 560.820 ;
        RECT -446.830 530.220 -445.030 560.220 ;
        RECT -415.030 530.220 -414.430 560.220 ;
        RECT -446.830 529.620 -414.430 530.220 ;
        RECT -407.530 560.220 -375.130 560.820 ;
        RECT -407.530 530.220 -406.930 560.220 ;
        RECT -376.930 530.220 -375.130 560.220 ;
        RECT -407.530 529.620 -375.130 530.220 ;
        RECT -371.830 560.220 -339.430 560.820 ;
        RECT -371.830 530.220 -370.030 560.220 ;
        RECT -340.030 530.220 -339.430 560.220 ;
        RECT -371.830 529.620 -339.430 530.220 ;
        RECT -332.530 560.220 -300.130 560.820 ;
        RECT -332.530 530.220 -331.930 560.220 ;
        RECT -301.930 530.220 -300.130 560.220 ;
        RECT -332.530 529.620 -300.130 530.220 ;
        RECT -296.830 560.220 -264.430 560.820 ;
        RECT -296.830 530.220 -295.030 560.220 ;
        RECT -265.030 530.220 -264.430 560.220 ;
        RECT -296.830 529.620 -264.430 530.220 ;
        RECT -257.530 560.220 -225.130 560.820 ;
        RECT -257.530 530.220 -256.930 560.220 ;
        RECT -226.930 530.220 -225.130 560.220 ;
        RECT -257.530 529.620 -225.130 530.220 ;
        RECT -221.830 560.220 -189.430 560.820 ;
        RECT -221.830 530.220 -220.030 560.220 ;
        RECT -190.030 530.220 -189.430 560.220 ;
        RECT -221.830 529.620 -189.430 530.220 ;
        RECT -182.530 560.220 -150.130 560.820 ;
        RECT -182.530 530.220 -181.930 560.220 ;
        RECT -151.930 530.220 -150.130 560.220 ;
        RECT -182.530 529.620 -150.130 530.220 ;
        RECT -146.830 560.220 -114.430 560.820 ;
        RECT -146.830 530.220 -145.030 560.220 ;
        RECT -115.030 530.220 -114.430 560.220 ;
        RECT -146.830 529.620 -114.430 530.220 ;
        RECT -107.530 560.220 -75.130 560.820 ;
        RECT -107.530 530.220 -106.930 560.220 ;
        RECT -76.930 530.220 -75.130 560.220 ;
        RECT -107.530 529.620 -75.130 530.220 ;
        RECT -71.830 560.220 -39.430 560.820 ;
        RECT -71.830 530.220 -70.030 560.220 ;
        RECT -40.030 530.220 -39.430 560.220 ;
        RECT -71.830 529.620 -39.430 530.220 ;
        RECT -32.530 560.220 -0.130 560.820 ;
        RECT -32.530 530.220 -31.930 560.220 ;
        RECT -1.930 530.220 -0.130 560.220 ;
        RECT -32.530 529.620 -0.130 530.220 ;
        RECT 3.170 560.220 35.570 560.820 ;
        RECT 3.170 530.220 4.970 560.220 ;
        RECT 34.970 530.220 35.570 560.220 ;
        RECT 3.170 529.620 35.570 530.220 ;
        RECT 42.470 560.220 74.870 560.820 ;
        RECT 42.470 530.220 43.070 560.220 ;
        RECT 73.070 530.220 74.870 560.220 ;
        RECT 42.470 529.620 74.870 530.220 ;
        RECT 78.170 560.220 110.570 560.820 ;
        RECT 78.170 530.220 79.970 560.220 ;
        RECT 109.970 530.220 110.570 560.220 ;
        RECT 78.170 529.620 110.570 530.220 ;
        RECT 117.470 560.220 149.870 560.820 ;
        RECT 117.470 530.220 118.070 560.220 ;
        RECT 148.070 530.220 149.870 560.220 ;
        RECT 117.470 529.620 149.870 530.220 ;
        RECT 153.170 560.220 185.570 560.820 ;
        RECT 153.170 530.220 154.970 560.220 ;
        RECT 184.970 530.220 185.570 560.220 ;
        RECT 153.170 529.620 185.570 530.220 ;
        RECT 192.470 560.220 224.870 560.820 ;
        RECT 192.470 530.220 193.070 560.220 ;
        RECT 223.070 530.220 224.870 560.220 ;
        RECT 192.470 529.620 224.870 530.220 ;
        RECT 228.170 560.220 260.570 560.820 ;
        RECT 228.170 530.220 229.970 560.220 ;
        RECT 259.970 530.220 260.570 560.220 ;
        RECT 228.170 529.620 260.570 530.220 ;
        RECT 267.470 560.220 299.870 560.820 ;
        RECT 267.470 530.220 268.070 560.220 ;
        RECT 298.070 530.220 299.870 560.220 ;
        RECT 267.470 529.620 299.870 530.220 ;
        RECT 303.170 560.220 335.570 560.820 ;
        RECT 303.170 530.220 304.970 560.220 ;
        RECT 334.970 530.220 335.570 560.220 ;
        RECT 303.170 529.620 335.570 530.220 ;
        RECT 342.470 560.220 374.870 560.820 ;
        RECT 342.470 530.220 343.070 560.220 ;
        RECT 373.070 530.220 374.870 560.220 ;
        RECT 342.470 529.620 374.870 530.220 ;
        RECT 378.170 560.220 410.570 560.820 ;
        RECT 378.170 530.220 379.970 560.220 ;
        RECT 409.970 530.220 410.570 560.220 ;
        RECT 378.170 529.620 410.570 530.220 ;
        RECT 417.470 560.220 449.870 560.820 ;
        RECT 417.470 530.220 418.070 560.220 ;
        RECT 448.070 530.220 449.870 560.220 ;
        RECT 417.470 529.620 449.870 530.220 ;
        RECT 453.170 560.220 485.570 560.820 ;
        RECT 453.170 530.220 454.970 560.220 ;
        RECT 484.970 530.220 485.570 560.220 ;
        RECT 453.170 529.620 485.570 530.220 ;
        RECT 492.470 560.220 524.870 560.820 ;
        RECT 492.470 530.220 493.070 560.220 ;
        RECT 523.070 530.220 524.870 560.220 ;
        RECT 492.470 529.620 524.870 530.220 ;
        RECT 528.170 560.220 560.570 560.820 ;
        RECT 528.170 530.220 529.970 560.220 ;
        RECT 559.970 530.220 560.570 560.220 ;
        RECT 528.170 529.620 560.570 530.220 ;
        RECT -557.530 525.220 -525.130 525.820 ;
        RECT -557.530 495.220 -556.930 525.220 ;
        RECT -526.930 495.220 -525.130 525.220 ;
        RECT -557.530 494.620 -525.130 495.220 ;
        RECT -521.830 525.220 -489.430 525.820 ;
        RECT -521.830 495.220 -520.030 525.220 ;
        RECT -490.030 495.220 -489.430 525.220 ;
        RECT -521.830 494.620 -489.430 495.220 ;
        RECT -482.530 525.220 -450.130 525.820 ;
        RECT -482.530 495.220 -481.930 525.220 ;
        RECT -451.930 495.220 -450.130 525.220 ;
        RECT -482.530 494.620 -450.130 495.220 ;
        RECT -446.830 525.220 -414.430 525.820 ;
        RECT -446.830 495.220 -445.030 525.220 ;
        RECT -415.030 495.220 -414.430 525.220 ;
        RECT -446.830 494.620 -414.430 495.220 ;
        RECT -407.530 525.220 -375.130 525.820 ;
        RECT -407.530 495.220 -406.930 525.220 ;
        RECT -376.930 495.220 -375.130 525.220 ;
        RECT -407.530 494.620 -375.130 495.220 ;
        RECT -371.830 525.220 -339.430 525.820 ;
        RECT -371.830 495.220 -370.030 525.220 ;
        RECT -340.030 495.220 -339.430 525.220 ;
        RECT -371.830 494.620 -339.430 495.220 ;
        RECT -332.530 525.220 -300.130 525.820 ;
        RECT -332.530 495.220 -331.930 525.220 ;
        RECT -301.930 495.220 -300.130 525.220 ;
        RECT -332.530 494.620 -300.130 495.220 ;
        RECT -296.830 525.220 -264.430 525.820 ;
        RECT -296.830 495.220 -295.030 525.220 ;
        RECT -265.030 495.220 -264.430 525.220 ;
        RECT -296.830 494.620 -264.430 495.220 ;
        RECT -257.530 525.220 -225.130 525.820 ;
        RECT -257.530 495.220 -256.930 525.220 ;
        RECT -226.930 495.220 -225.130 525.220 ;
        RECT -257.530 494.620 -225.130 495.220 ;
        RECT -221.830 525.220 -189.430 525.820 ;
        RECT -221.830 495.220 -220.030 525.220 ;
        RECT -190.030 495.220 -189.430 525.220 ;
        RECT -221.830 494.620 -189.430 495.220 ;
        RECT -182.530 525.220 -150.130 525.820 ;
        RECT -182.530 495.220 -181.930 525.220 ;
        RECT -151.930 495.220 -150.130 525.220 ;
        RECT -182.530 494.620 -150.130 495.220 ;
        RECT -146.830 525.220 -114.430 525.820 ;
        RECT -146.830 495.220 -145.030 525.220 ;
        RECT -115.030 495.220 -114.430 525.220 ;
        RECT -146.830 494.620 -114.430 495.220 ;
        RECT -107.530 525.220 -75.130 525.820 ;
        RECT -107.530 495.220 -106.930 525.220 ;
        RECT -76.930 495.220 -75.130 525.220 ;
        RECT -107.530 494.620 -75.130 495.220 ;
        RECT -71.830 525.220 -39.430 525.820 ;
        RECT -71.830 495.220 -70.030 525.220 ;
        RECT -40.030 495.220 -39.430 525.220 ;
        RECT -71.830 494.620 -39.430 495.220 ;
        RECT -32.530 525.220 -0.130 525.820 ;
        RECT -32.530 495.220 -31.930 525.220 ;
        RECT -1.930 495.220 -0.130 525.220 ;
        RECT -32.530 494.620 -0.130 495.220 ;
        RECT 3.170 525.220 35.570 525.820 ;
        RECT 3.170 495.220 4.970 525.220 ;
        RECT 34.970 495.220 35.570 525.220 ;
        RECT 3.170 494.620 35.570 495.220 ;
        RECT 42.470 525.220 74.870 525.820 ;
        RECT 42.470 495.220 43.070 525.220 ;
        RECT 73.070 495.220 74.870 525.220 ;
        RECT 42.470 494.620 74.870 495.220 ;
        RECT 78.170 525.220 110.570 525.820 ;
        RECT 78.170 495.220 79.970 525.220 ;
        RECT 109.970 495.220 110.570 525.220 ;
        RECT 78.170 494.620 110.570 495.220 ;
        RECT 117.470 525.220 149.870 525.820 ;
        RECT 117.470 495.220 118.070 525.220 ;
        RECT 148.070 495.220 149.870 525.220 ;
        RECT 117.470 494.620 149.870 495.220 ;
        RECT 153.170 525.220 185.570 525.820 ;
        RECT 153.170 495.220 154.970 525.220 ;
        RECT 184.970 495.220 185.570 525.220 ;
        RECT 153.170 494.620 185.570 495.220 ;
        RECT 192.470 525.220 224.870 525.820 ;
        RECT 192.470 495.220 193.070 525.220 ;
        RECT 223.070 495.220 224.870 525.220 ;
        RECT 192.470 494.620 224.870 495.220 ;
        RECT 228.170 525.220 260.570 525.820 ;
        RECT 228.170 495.220 229.970 525.220 ;
        RECT 259.970 495.220 260.570 525.220 ;
        RECT 228.170 494.620 260.570 495.220 ;
        RECT 267.470 525.220 299.870 525.820 ;
        RECT 267.470 495.220 268.070 525.220 ;
        RECT 298.070 495.220 299.870 525.220 ;
        RECT 267.470 494.620 299.870 495.220 ;
        RECT 303.170 525.220 335.570 525.820 ;
        RECT 303.170 495.220 304.970 525.220 ;
        RECT 334.970 495.220 335.570 525.220 ;
        RECT 303.170 494.620 335.570 495.220 ;
        RECT 342.470 525.220 374.870 525.820 ;
        RECT 342.470 495.220 343.070 525.220 ;
        RECT 373.070 495.220 374.870 525.220 ;
        RECT 342.470 494.620 374.870 495.220 ;
        RECT 378.170 525.220 410.570 525.820 ;
        RECT 378.170 495.220 379.970 525.220 ;
        RECT 409.970 495.220 410.570 525.220 ;
        RECT 378.170 494.620 410.570 495.220 ;
        RECT 417.470 525.220 449.870 525.820 ;
        RECT 417.470 495.220 418.070 525.220 ;
        RECT 448.070 495.220 449.870 525.220 ;
        RECT 417.470 494.620 449.870 495.220 ;
        RECT 453.170 525.220 485.570 525.820 ;
        RECT 453.170 495.220 454.970 525.220 ;
        RECT 484.970 495.220 485.570 525.220 ;
        RECT 453.170 494.620 485.570 495.220 ;
        RECT 492.470 525.220 524.870 525.820 ;
        RECT 492.470 495.220 493.070 525.220 ;
        RECT 523.070 495.220 524.870 525.220 ;
        RECT 492.470 494.620 524.870 495.220 ;
        RECT 528.170 525.220 560.570 525.820 ;
        RECT 528.170 495.220 529.970 525.220 ;
        RECT 559.970 495.220 560.570 525.220 ;
        RECT 528.170 494.620 560.570 495.220 ;
        RECT -557.530 490.220 -525.130 490.820 ;
        RECT -557.530 460.220 -556.930 490.220 ;
        RECT -526.930 460.220 -525.130 490.220 ;
        RECT -557.530 459.620 -525.130 460.220 ;
        RECT -521.830 490.220 -489.430 490.820 ;
        RECT -521.830 460.220 -520.030 490.220 ;
        RECT -490.030 460.220 -489.430 490.220 ;
        RECT -521.830 459.620 -489.430 460.220 ;
        RECT -482.530 490.220 -450.130 490.820 ;
        RECT -482.530 460.220 -481.930 490.220 ;
        RECT -451.930 460.220 -450.130 490.220 ;
        RECT -482.530 459.620 -450.130 460.220 ;
        RECT -446.830 490.220 -414.430 490.820 ;
        RECT -446.830 460.220 -445.030 490.220 ;
        RECT -415.030 460.220 -414.430 490.220 ;
        RECT -446.830 459.620 -414.430 460.220 ;
        RECT -407.530 490.220 -375.130 490.820 ;
        RECT -407.530 460.220 -406.930 490.220 ;
        RECT -376.930 460.220 -375.130 490.220 ;
        RECT -407.530 459.620 -375.130 460.220 ;
        RECT -371.830 490.220 -339.430 490.820 ;
        RECT -371.830 460.220 -370.030 490.220 ;
        RECT -340.030 460.220 -339.430 490.220 ;
        RECT -371.830 459.620 -339.430 460.220 ;
        RECT -332.530 490.220 -300.130 490.820 ;
        RECT -332.530 460.220 -331.930 490.220 ;
        RECT -301.930 460.220 -300.130 490.220 ;
        RECT -332.530 459.620 -300.130 460.220 ;
        RECT -296.830 490.220 -264.430 490.820 ;
        RECT -296.830 460.220 -295.030 490.220 ;
        RECT -265.030 460.220 -264.430 490.220 ;
        RECT -296.830 459.620 -264.430 460.220 ;
        RECT -257.530 490.220 -225.130 490.820 ;
        RECT -257.530 460.220 -256.930 490.220 ;
        RECT -226.930 460.220 -225.130 490.220 ;
        RECT -257.530 459.620 -225.130 460.220 ;
        RECT -221.830 490.220 -189.430 490.820 ;
        RECT -221.830 460.220 -220.030 490.220 ;
        RECT -190.030 460.220 -189.430 490.220 ;
        RECT -221.830 459.620 -189.430 460.220 ;
        RECT -182.530 490.220 -150.130 490.820 ;
        RECT -182.530 460.220 -181.930 490.220 ;
        RECT -151.930 460.220 -150.130 490.220 ;
        RECT -182.530 459.620 -150.130 460.220 ;
        RECT -146.830 490.220 -114.430 490.820 ;
        RECT -146.830 460.220 -145.030 490.220 ;
        RECT -115.030 460.220 -114.430 490.220 ;
        RECT -146.830 459.620 -114.430 460.220 ;
        RECT -107.530 490.220 -75.130 490.820 ;
        RECT -107.530 460.220 -106.930 490.220 ;
        RECT -76.930 460.220 -75.130 490.220 ;
        RECT -107.530 459.620 -75.130 460.220 ;
        RECT -71.830 490.220 -39.430 490.820 ;
        RECT -71.830 460.220 -70.030 490.220 ;
        RECT -40.030 460.220 -39.430 490.220 ;
        RECT -71.830 459.620 -39.430 460.220 ;
        RECT -32.530 490.220 -0.130 490.820 ;
        RECT -32.530 460.220 -31.930 490.220 ;
        RECT -1.930 460.220 -0.130 490.220 ;
        RECT -32.530 459.620 -0.130 460.220 ;
        RECT 3.170 490.220 35.570 490.820 ;
        RECT 3.170 460.220 4.970 490.220 ;
        RECT 34.970 460.220 35.570 490.220 ;
        RECT 3.170 459.620 35.570 460.220 ;
        RECT 42.470 490.220 74.870 490.820 ;
        RECT 42.470 460.220 43.070 490.220 ;
        RECT 73.070 460.220 74.870 490.220 ;
        RECT 42.470 459.620 74.870 460.220 ;
        RECT 78.170 490.220 110.570 490.820 ;
        RECT 78.170 460.220 79.970 490.220 ;
        RECT 109.970 460.220 110.570 490.220 ;
        RECT 78.170 459.620 110.570 460.220 ;
        RECT 117.470 490.220 149.870 490.820 ;
        RECT 117.470 460.220 118.070 490.220 ;
        RECT 148.070 460.220 149.870 490.220 ;
        RECT 117.470 459.620 149.870 460.220 ;
        RECT 153.170 490.220 185.570 490.820 ;
        RECT 153.170 460.220 154.970 490.220 ;
        RECT 184.970 460.220 185.570 490.220 ;
        RECT 153.170 459.620 185.570 460.220 ;
        RECT 192.470 490.220 224.870 490.820 ;
        RECT 192.470 460.220 193.070 490.220 ;
        RECT 223.070 460.220 224.870 490.220 ;
        RECT 192.470 459.620 224.870 460.220 ;
        RECT 228.170 490.220 260.570 490.820 ;
        RECT 228.170 460.220 229.970 490.220 ;
        RECT 259.970 460.220 260.570 490.220 ;
        RECT 228.170 459.620 260.570 460.220 ;
        RECT 267.470 490.220 299.870 490.820 ;
        RECT 267.470 460.220 268.070 490.220 ;
        RECT 298.070 460.220 299.870 490.220 ;
        RECT 267.470 459.620 299.870 460.220 ;
        RECT 303.170 490.220 335.570 490.820 ;
        RECT 303.170 460.220 304.970 490.220 ;
        RECT 334.970 460.220 335.570 490.220 ;
        RECT 303.170 459.620 335.570 460.220 ;
        RECT 342.470 490.220 374.870 490.820 ;
        RECT 342.470 460.220 343.070 490.220 ;
        RECT 373.070 460.220 374.870 490.220 ;
        RECT 342.470 459.620 374.870 460.220 ;
        RECT 378.170 490.220 410.570 490.820 ;
        RECT 378.170 460.220 379.970 490.220 ;
        RECT 409.970 460.220 410.570 490.220 ;
        RECT 378.170 459.620 410.570 460.220 ;
        RECT 417.470 490.220 449.870 490.820 ;
        RECT 417.470 460.220 418.070 490.220 ;
        RECT 448.070 460.220 449.870 490.220 ;
        RECT 417.470 459.620 449.870 460.220 ;
        RECT 453.170 490.220 485.570 490.820 ;
        RECT 453.170 460.220 454.970 490.220 ;
        RECT 484.970 460.220 485.570 490.220 ;
        RECT 453.170 459.620 485.570 460.220 ;
        RECT 492.470 490.220 524.870 490.820 ;
        RECT 492.470 460.220 493.070 490.220 ;
        RECT 523.070 460.220 524.870 490.220 ;
        RECT 492.470 459.620 524.870 460.220 ;
        RECT 528.170 490.220 560.570 490.820 ;
        RECT 528.170 460.220 529.970 490.220 ;
        RECT 559.970 460.220 560.570 490.220 ;
        RECT 528.170 459.620 560.570 460.220 ;
        RECT -557.530 455.220 -525.130 455.820 ;
        RECT -557.530 425.220 -556.930 455.220 ;
        RECT -526.930 425.220 -525.130 455.220 ;
        RECT -557.530 424.620 -525.130 425.220 ;
        RECT -521.830 455.220 -489.430 455.820 ;
        RECT -521.830 425.220 -520.030 455.220 ;
        RECT -490.030 425.220 -489.430 455.220 ;
        RECT -521.830 424.620 -489.430 425.220 ;
        RECT -482.530 455.220 -450.130 455.820 ;
        RECT -482.530 425.220 -481.930 455.220 ;
        RECT -451.930 425.220 -450.130 455.220 ;
        RECT -482.530 424.620 -450.130 425.220 ;
        RECT -446.830 455.220 -414.430 455.820 ;
        RECT -446.830 425.220 -445.030 455.220 ;
        RECT -415.030 425.220 -414.430 455.220 ;
        RECT -446.830 424.620 -414.430 425.220 ;
        RECT -407.530 455.220 -375.130 455.820 ;
        RECT -407.530 425.220 -406.930 455.220 ;
        RECT -376.930 425.220 -375.130 455.220 ;
        RECT -407.530 424.620 -375.130 425.220 ;
        RECT -371.830 455.220 -339.430 455.820 ;
        RECT -371.830 425.220 -370.030 455.220 ;
        RECT -340.030 425.220 -339.430 455.220 ;
        RECT -371.830 424.620 -339.430 425.220 ;
        RECT -332.530 455.220 -300.130 455.820 ;
        RECT -332.530 425.220 -331.930 455.220 ;
        RECT -301.930 425.220 -300.130 455.220 ;
        RECT -332.530 424.620 -300.130 425.220 ;
        RECT -296.830 455.220 -264.430 455.820 ;
        RECT -296.830 425.220 -295.030 455.220 ;
        RECT -265.030 425.220 -264.430 455.220 ;
        RECT -296.830 424.620 -264.430 425.220 ;
        RECT -257.530 455.220 -225.130 455.820 ;
        RECT -257.530 425.220 -256.930 455.220 ;
        RECT -226.930 425.220 -225.130 455.220 ;
        RECT -257.530 424.620 -225.130 425.220 ;
        RECT -221.830 455.220 -189.430 455.820 ;
        RECT -221.830 425.220 -220.030 455.220 ;
        RECT -190.030 425.220 -189.430 455.220 ;
        RECT -221.830 424.620 -189.430 425.220 ;
        RECT -182.530 455.220 -150.130 455.820 ;
        RECT -182.530 425.220 -181.930 455.220 ;
        RECT -151.930 425.220 -150.130 455.220 ;
        RECT -182.530 424.620 -150.130 425.220 ;
        RECT -146.830 455.220 -114.430 455.820 ;
        RECT -146.830 425.220 -145.030 455.220 ;
        RECT -115.030 425.220 -114.430 455.220 ;
        RECT -146.830 424.620 -114.430 425.220 ;
        RECT -107.530 455.220 -75.130 455.820 ;
        RECT -107.530 425.220 -106.930 455.220 ;
        RECT -76.930 425.220 -75.130 455.220 ;
        RECT -107.530 424.620 -75.130 425.220 ;
        RECT -71.830 455.220 -39.430 455.820 ;
        RECT -71.830 425.220 -70.030 455.220 ;
        RECT -40.030 425.220 -39.430 455.220 ;
        RECT -71.830 424.620 -39.430 425.220 ;
        RECT -32.530 455.220 -0.130 455.820 ;
        RECT -32.530 425.220 -31.930 455.220 ;
        RECT -1.930 425.220 -0.130 455.220 ;
        RECT -32.530 424.620 -0.130 425.220 ;
        RECT 3.170 455.220 35.570 455.820 ;
        RECT 3.170 425.220 4.970 455.220 ;
        RECT 34.970 425.220 35.570 455.220 ;
        RECT 3.170 424.620 35.570 425.220 ;
        RECT 42.470 455.220 74.870 455.820 ;
        RECT 42.470 425.220 43.070 455.220 ;
        RECT 73.070 425.220 74.870 455.220 ;
        RECT 42.470 424.620 74.870 425.220 ;
        RECT 78.170 455.220 110.570 455.820 ;
        RECT 78.170 425.220 79.970 455.220 ;
        RECT 109.970 425.220 110.570 455.220 ;
        RECT 78.170 424.620 110.570 425.220 ;
        RECT 117.470 455.220 149.870 455.820 ;
        RECT 117.470 425.220 118.070 455.220 ;
        RECT 148.070 425.220 149.870 455.220 ;
        RECT 117.470 424.620 149.870 425.220 ;
        RECT 153.170 455.220 185.570 455.820 ;
        RECT 153.170 425.220 154.970 455.220 ;
        RECT 184.970 425.220 185.570 455.220 ;
        RECT 153.170 424.620 185.570 425.220 ;
        RECT 192.470 455.220 224.870 455.820 ;
        RECT 192.470 425.220 193.070 455.220 ;
        RECT 223.070 425.220 224.870 455.220 ;
        RECT 192.470 424.620 224.870 425.220 ;
        RECT 228.170 455.220 260.570 455.820 ;
        RECT 228.170 425.220 229.970 455.220 ;
        RECT 259.970 425.220 260.570 455.220 ;
        RECT 228.170 424.620 260.570 425.220 ;
        RECT 267.470 455.220 299.870 455.820 ;
        RECT 267.470 425.220 268.070 455.220 ;
        RECT 298.070 425.220 299.870 455.220 ;
        RECT 267.470 424.620 299.870 425.220 ;
        RECT 303.170 455.220 335.570 455.820 ;
        RECT 303.170 425.220 304.970 455.220 ;
        RECT 334.970 425.220 335.570 455.220 ;
        RECT 303.170 424.620 335.570 425.220 ;
        RECT 342.470 455.220 374.870 455.820 ;
        RECT 342.470 425.220 343.070 455.220 ;
        RECT 373.070 425.220 374.870 455.220 ;
        RECT 342.470 424.620 374.870 425.220 ;
        RECT 378.170 455.220 410.570 455.820 ;
        RECT 378.170 425.220 379.970 455.220 ;
        RECT 409.970 425.220 410.570 455.220 ;
        RECT 378.170 424.620 410.570 425.220 ;
        RECT 417.470 455.220 449.870 455.820 ;
        RECT 417.470 425.220 418.070 455.220 ;
        RECT 448.070 425.220 449.870 455.220 ;
        RECT 417.470 424.620 449.870 425.220 ;
        RECT 453.170 455.220 485.570 455.820 ;
        RECT 453.170 425.220 454.970 455.220 ;
        RECT 484.970 425.220 485.570 455.220 ;
        RECT 453.170 424.620 485.570 425.220 ;
        RECT 492.470 455.220 524.870 455.820 ;
        RECT 492.470 425.220 493.070 455.220 ;
        RECT 523.070 425.220 524.870 455.220 ;
        RECT 492.470 424.620 524.870 425.220 ;
        RECT 528.170 455.220 560.570 455.820 ;
        RECT 528.170 425.220 529.970 455.220 ;
        RECT 559.970 425.220 560.570 455.220 ;
        RECT 528.170 424.620 560.570 425.220 ;
        RECT -557.530 420.220 -525.130 420.820 ;
        RECT -557.530 390.220 -556.930 420.220 ;
        RECT -526.930 390.220 -525.130 420.220 ;
        RECT -557.530 389.620 -525.130 390.220 ;
        RECT -521.830 420.220 -489.430 420.820 ;
        RECT -521.830 390.220 -520.030 420.220 ;
        RECT -490.030 390.220 -489.430 420.220 ;
        RECT -521.830 389.620 -489.430 390.220 ;
        RECT -482.530 420.220 -450.130 420.820 ;
        RECT -482.530 390.220 -481.930 420.220 ;
        RECT -451.930 390.220 -450.130 420.220 ;
        RECT -482.530 389.620 -450.130 390.220 ;
        RECT -446.830 420.220 -414.430 420.820 ;
        RECT -446.830 390.220 -445.030 420.220 ;
        RECT -415.030 390.220 -414.430 420.220 ;
        RECT -446.830 389.620 -414.430 390.220 ;
        RECT -407.530 420.220 -375.130 420.820 ;
        RECT -407.530 390.220 -406.930 420.220 ;
        RECT -376.930 390.220 -375.130 420.220 ;
        RECT -407.530 389.620 -375.130 390.220 ;
        RECT -371.830 420.220 -339.430 420.820 ;
        RECT -371.830 390.220 -370.030 420.220 ;
        RECT -340.030 390.220 -339.430 420.220 ;
        RECT -371.830 389.620 -339.430 390.220 ;
        RECT -332.530 420.220 -300.130 420.820 ;
        RECT -332.530 390.220 -331.930 420.220 ;
        RECT -301.930 390.220 -300.130 420.220 ;
        RECT -332.530 389.620 -300.130 390.220 ;
        RECT -296.830 420.220 -264.430 420.820 ;
        RECT -296.830 390.220 -295.030 420.220 ;
        RECT -265.030 390.220 -264.430 420.220 ;
        RECT -296.830 389.620 -264.430 390.220 ;
        RECT -257.530 420.220 -225.130 420.820 ;
        RECT -257.530 390.220 -256.930 420.220 ;
        RECT -226.930 390.220 -225.130 420.220 ;
        RECT -257.530 389.620 -225.130 390.220 ;
        RECT -221.830 420.220 -189.430 420.820 ;
        RECT -221.830 390.220 -220.030 420.220 ;
        RECT -190.030 390.220 -189.430 420.220 ;
        RECT -221.830 389.620 -189.430 390.220 ;
        RECT -182.530 420.220 -150.130 420.820 ;
        RECT -182.530 390.220 -181.930 420.220 ;
        RECT -151.930 390.220 -150.130 420.220 ;
        RECT -182.530 389.620 -150.130 390.220 ;
        RECT -146.830 420.220 -114.430 420.820 ;
        RECT -146.830 390.220 -145.030 420.220 ;
        RECT -115.030 390.220 -114.430 420.220 ;
        RECT -146.830 389.620 -114.430 390.220 ;
        RECT -107.530 420.220 -75.130 420.820 ;
        RECT -107.530 390.220 -106.930 420.220 ;
        RECT -76.930 390.220 -75.130 420.220 ;
        RECT -107.530 389.620 -75.130 390.220 ;
        RECT -71.830 420.220 -39.430 420.820 ;
        RECT -71.830 390.220 -70.030 420.220 ;
        RECT -40.030 390.220 -39.430 420.220 ;
        RECT -71.830 389.620 -39.430 390.220 ;
        RECT -32.530 420.220 -0.130 420.820 ;
        RECT -32.530 390.220 -31.930 420.220 ;
        RECT -1.930 390.220 -0.130 420.220 ;
        RECT -32.530 389.620 -0.130 390.220 ;
        RECT 3.170 420.220 35.570 420.820 ;
        RECT 3.170 390.220 4.970 420.220 ;
        RECT 34.970 390.220 35.570 420.220 ;
        RECT 3.170 389.620 35.570 390.220 ;
        RECT 42.470 420.220 74.870 420.820 ;
        RECT 42.470 390.220 43.070 420.220 ;
        RECT 73.070 390.220 74.870 420.220 ;
        RECT 42.470 389.620 74.870 390.220 ;
        RECT 78.170 420.220 110.570 420.820 ;
        RECT 78.170 390.220 79.970 420.220 ;
        RECT 109.970 390.220 110.570 420.220 ;
        RECT 78.170 389.620 110.570 390.220 ;
        RECT 117.470 420.220 149.870 420.820 ;
        RECT 117.470 390.220 118.070 420.220 ;
        RECT 148.070 390.220 149.870 420.220 ;
        RECT 117.470 389.620 149.870 390.220 ;
        RECT 153.170 420.220 185.570 420.820 ;
        RECT 153.170 390.220 154.970 420.220 ;
        RECT 184.970 390.220 185.570 420.220 ;
        RECT 153.170 389.620 185.570 390.220 ;
        RECT 192.470 420.220 224.870 420.820 ;
        RECT 192.470 390.220 193.070 420.220 ;
        RECT 223.070 390.220 224.870 420.220 ;
        RECT 192.470 389.620 224.870 390.220 ;
        RECT 228.170 420.220 260.570 420.820 ;
        RECT 228.170 390.220 229.970 420.220 ;
        RECT 259.970 390.220 260.570 420.220 ;
        RECT 228.170 389.620 260.570 390.220 ;
        RECT 267.470 420.220 299.870 420.820 ;
        RECT 267.470 390.220 268.070 420.220 ;
        RECT 298.070 390.220 299.870 420.220 ;
        RECT 267.470 389.620 299.870 390.220 ;
        RECT 303.170 420.220 335.570 420.820 ;
        RECT 303.170 390.220 304.970 420.220 ;
        RECT 334.970 390.220 335.570 420.220 ;
        RECT 303.170 389.620 335.570 390.220 ;
        RECT 342.470 420.220 374.870 420.820 ;
        RECT 342.470 390.220 343.070 420.220 ;
        RECT 373.070 390.220 374.870 420.220 ;
        RECT 342.470 389.620 374.870 390.220 ;
        RECT 378.170 420.220 410.570 420.820 ;
        RECT 378.170 390.220 379.970 420.220 ;
        RECT 409.970 390.220 410.570 420.220 ;
        RECT 378.170 389.620 410.570 390.220 ;
        RECT 417.470 420.220 449.870 420.820 ;
        RECT 417.470 390.220 418.070 420.220 ;
        RECT 448.070 390.220 449.870 420.220 ;
        RECT 417.470 389.620 449.870 390.220 ;
        RECT 453.170 420.220 485.570 420.820 ;
        RECT 453.170 390.220 454.970 420.220 ;
        RECT 484.970 390.220 485.570 420.220 ;
        RECT 453.170 389.620 485.570 390.220 ;
        RECT 492.470 420.220 524.870 420.820 ;
        RECT 492.470 390.220 493.070 420.220 ;
        RECT 523.070 390.220 524.870 420.220 ;
        RECT 492.470 389.620 524.870 390.220 ;
        RECT 528.170 420.220 560.570 420.820 ;
        RECT 528.170 390.220 529.970 420.220 ;
        RECT 559.970 390.220 560.570 420.220 ;
        RECT 528.170 389.620 560.570 390.220 ;
        RECT 763.320 352.720 841.320 1085.700 ;
        RECT -838.480 172.480 -543.480 352.720 ;
        RECT -533.380 320.920 -430.980 321.520 ;
        RECT -533.380 220.920 -532.780 320.920 ;
        RECT -432.780 220.920 -430.980 320.920 ;
        RECT -533.380 220.320 -430.980 220.920 ;
        RECT -425.980 320.920 -323.580 321.520 ;
        RECT -425.980 220.920 -424.180 320.920 ;
        RECT -324.180 220.920 -323.580 320.920 ;
        RECT -425.980 220.320 -323.580 220.920 ;
        RECT -318.380 320.920 -215.980 321.520 ;
        RECT -318.380 220.920 -317.780 320.920 ;
        RECT -217.780 220.920 -215.980 320.920 ;
        RECT -318.380 220.320 -215.980 220.920 ;
        RECT -210.980 320.920 -108.580 321.520 ;
        RECT -210.980 220.920 -209.180 320.920 ;
        RECT -109.180 220.920 -108.580 320.920 ;
        RECT -210.980 220.320 -108.580 220.920 ;
        RECT -103.380 320.920 -0.980 321.520 ;
        RECT -103.380 220.920 -102.780 320.920 ;
        RECT -2.780 220.920 -0.980 320.920 ;
        RECT -103.380 220.320 -0.980 220.920 ;
        RECT 4.020 320.920 106.420 321.520 ;
        RECT 4.020 220.920 5.820 320.920 ;
        RECT 105.820 220.920 106.420 320.920 ;
        RECT 4.020 220.320 106.420 220.920 ;
        RECT 111.620 320.920 214.020 321.520 ;
        RECT 111.620 220.920 112.220 320.920 ;
        RECT 212.220 220.920 214.020 320.920 ;
        RECT 111.620 220.320 214.020 220.920 ;
        RECT 219.020 320.920 321.420 321.520 ;
        RECT 219.020 220.920 220.820 320.920 ;
        RECT 320.820 220.920 321.420 320.920 ;
        RECT 219.020 220.320 321.420 220.920 ;
        RECT 326.620 320.920 429.020 321.520 ;
        RECT 326.620 220.920 327.220 320.920 ;
        RECT 427.220 220.920 429.020 320.920 ;
        RECT 326.620 220.320 429.020 220.920 ;
        RECT 434.020 320.920 536.420 321.520 ;
        RECT 434.020 220.920 435.820 320.920 ;
        RECT 535.820 220.920 536.420 320.920 ;
        RECT 434.020 220.320 536.420 220.920 ;
        RECT -838.480 132.620 -760.480 172.480 ;
        RECT -509.680 171.430 -478.480 173.230 ;
        RECT -509.680 141.430 -509.080 171.430 ;
        RECT -479.080 141.430 -478.480 171.430 ;
        RECT -509.680 140.830 -478.480 141.430 ;
        RECT -469.680 171.430 -438.480 173.230 ;
        RECT -469.680 141.430 -469.080 171.430 ;
        RECT -439.080 141.430 -438.480 171.430 ;
        RECT -469.680 140.830 -438.480 141.430 ;
        RECT -429.680 171.430 -398.480 173.230 ;
        RECT -429.680 141.430 -429.080 171.430 ;
        RECT -399.080 141.430 -398.480 171.430 ;
        RECT -429.680 140.830 -398.480 141.430 ;
        RECT -389.680 171.430 -358.480 173.230 ;
        RECT -389.680 141.430 -389.080 171.430 ;
        RECT -359.080 141.430 -358.480 171.430 ;
        RECT -389.680 140.830 -358.480 141.430 ;
        RECT -349.680 171.430 -318.480 173.230 ;
        RECT -349.680 141.430 -349.080 171.430 ;
        RECT -319.080 141.430 -318.480 171.430 ;
        RECT -349.680 140.830 -318.480 141.430 ;
        RECT -309.680 171.430 -278.480 173.230 ;
        RECT -309.680 141.430 -309.080 171.430 ;
        RECT -279.080 141.430 -278.480 171.430 ;
        RECT -309.680 140.830 -278.480 141.430 ;
        RECT -269.680 171.430 -238.480 173.230 ;
        RECT -269.680 141.430 -269.080 171.430 ;
        RECT -239.080 141.430 -238.480 171.430 ;
        RECT -269.680 140.830 -238.480 141.430 ;
        RECT -229.680 171.430 -198.480 173.230 ;
        RECT -229.680 141.430 -229.080 171.430 ;
        RECT -199.080 141.430 -198.480 171.430 ;
        RECT -229.680 140.830 -198.480 141.430 ;
        RECT -189.680 171.430 -158.480 173.230 ;
        RECT -189.680 141.430 -189.080 171.430 ;
        RECT -159.080 141.430 -158.480 171.430 ;
        RECT -189.680 140.830 -158.480 141.430 ;
        RECT -149.680 171.430 -118.480 173.230 ;
        RECT -149.680 141.430 -149.080 171.430 ;
        RECT -119.080 141.430 -118.480 171.430 ;
        RECT -149.680 140.830 -118.480 141.430 ;
        RECT -109.680 171.430 -78.480 173.230 ;
        RECT -109.680 141.430 -109.080 171.430 ;
        RECT -79.080 141.430 -78.480 171.430 ;
        RECT -109.680 140.830 -78.480 141.430 ;
        RECT -69.680 171.430 -38.480 173.230 ;
        RECT -69.680 141.430 -69.080 171.430 ;
        RECT -39.080 141.430 -38.480 171.430 ;
        RECT -69.680 140.830 -38.480 141.430 ;
        RECT -29.680 171.430 1.520 173.230 ;
        RECT -29.680 141.430 -29.080 171.430 ;
        RECT 0.920 141.430 1.520 171.430 ;
        RECT -29.680 140.830 1.520 141.430 ;
        RECT 10.320 171.430 41.520 173.230 ;
        RECT 10.320 141.430 10.920 171.430 ;
        RECT 40.920 141.430 41.520 171.430 ;
        RECT 10.320 140.830 41.520 141.430 ;
        RECT 50.320 171.430 81.520 173.230 ;
        RECT 50.320 141.430 50.920 171.430 ;
        RECT 80.920 141.430 81.520 171.430 ;
        RECT 50.320 140.830 81.520 141.430 ;
        RECT 90.320 171.430 121.520 173.230 ;
        RECT 90.320 141.430 90.920 171.430 ;
        RECT 120.920 141.430 121.520 171.430 ;
        RECT 90.320 140.830 121.520 141.430 ;
        RECT 130.320 171.430 161.520 173.230 ;
        RECT 130.320 141.430 130.920 171.430 ;
        RECT 160.920 141.430 161.520 171.430 ;
        RECT 130.320 140.830 161.520 141.430 ;
        RECT 170.320 171.430 201.520 173.230 ;
        RECT 170.320 141.430 170.920 171.430 ;
        RECT 200.920 141.430 201.520 171.430 ;
        RECT 170.320 140.830 201.520 141.430 ;
        RECT 225.920 171.430 257.120 173.230 ;
        RECT 225.920 141.430 226.520 171.430 ;
        RECT 256.520 141.430 257.120 171.430 ;
        RECT 225.920 140.830 257.120 141.430 ;
        RECT 265.920 171.430 297.120 173.230 ;
        RECT 265.920 141.430 266.520 171.430 ;
        RECT 296.520 141.430 297.120 171.430 ;
        RECT 265.920 140.830 297.120 141.430 ;
        RECT 305.920 171.430 337.120 173.230 ;
        RECT 305.920 141.430 306.520 171.430 ;
        RECT 336.520 141.430 337.120 171.430 ;
        RECT 305.920 140.830 337.120 141.430 ;
        RECT 345.920 171.430 377.120 173.230 ;
        RECT 345.920 141.430 346.520 171.430 ;
        RECT 376.520 141.430 377.120 171.430 ;
        RECT 345.920 140.830 377.120 141.430 ;
        RECT 385.920 171.430 417.120 173.230 ;
        RECT 385.920 141.430 386.520 171.430 ;
        RECT 416.520 141.430 417.120 171.430 ;
        RECT 385.920 140.830 417.120 141.430 ;
        RECT 425.920 171.430 457.120 173.230 ;
        RECT 425.920 141.430 426.520 171.430 ;
        RECT 456.520 141.430 457.120 171.430 ;
        RECT 425.920 140.830 457.120 141.430 ;
        RECT 465.920 171.430 497.120 173.230 ;
        RECT 546.520 172.480 841.320 352.720 ;
        RECT 465.920 141.430 466.520 171.430 ;
        RECT 496.520 141.430 497.120 171.430 ;
        RECT 465.920 140.830 497.120 141.430 ;
        RECT 763.320 132.620 841.320 172.480 ;
        RECT -839.240 127.660 841.320 132.620 ;
        RECT -839.240 -127.660 -760.480 127.660 ;
        RECT 194.795 9.220 228.000 127.660 ;
        RECT 194.795 0.220 229.590 9.220 ;
        RECT 194.795 -12.135 228.000 0.220 ;
        RECT 194.795 -13.735 235.700 -12.135 ;
        RECT 194.795 -127.660 228.000 -13.735 ;
        RECT 336.700 -127.660 338.300 127.660 ;
        RECT 378.280 -127.660 379.880 127.660 ;
        RECT 419.860 -127.660 421.460 127.660 ;
        RECT 461.440 -127.660 463.040 127.660 ;
        RECT 763.320 -127.660 841.320 127.660 ;
        RECT -839.240 -132.620 841.320 -127.660 ;
        RECT -838.480 -172.480 -760.480 -132.620 ;
        RECT -509.680 -141.430 -478.480 -140.830 ;
        RECT -509.680 -171.430 -509.080 -141.430 ;
        RECT -479.080 -171.430 -478.480 -141.430 ;
        RECT -838.480 -352.720 -543.480 -172.480 ;
        RECT -509.680 -173.230 -478.480 -171.430 ;
        RECT -469.680 -141.430 -438.480 -140.830 ;
        RECT -469.680 -171.430 -469.080 -141.430 ;
        RECT -439.080 -171.430 -438.480 -141.430 ;
        RECT -469.680 -173.230 -438.480 -171.430 ;
        RECT -429.680 -141.430 -398.480 -140.830 ;
        RECT -429.680 -171.430 -429.080 -141.430 ;
        RECT -399.080 -171.430 -398.480 -141.430 ;
        RECT -429.680 -173.230 -398.480 -171.430 ;
        RECT -389.680 -141.430 -358.480 -140.830 ;
        RECT -389.680 -171.430 -389.080 -141.430 ;
        RECT -359.080 -171.430 -358.480 -141.430 ;
        RECT -389.680 -173.230 -358.480 -171.430 ;
        RECT -349.680 -141.430 -318.480 -140.830 ;
        RECT -349.680 -171.430 -349.080 -141.430 ;
        RECT -319.080 -171.430 -318.480 -141.430 ;
        RECT -349.680 -173.230 -318.480 -171.430 ;
        RECT -309.680 -141.430 -278.480 -140.830 ;
        RECT -309.680 -171.430 -309.080 -141.430 ;
        RECT -279.080 -171.430 -278.480 -141.430 ;
        RECT -309.680 -173.230 -278.480 -171.430 ;
        RECT -269.680 -141.430 -238.480 -140.830 ;
        RECT -269.680 -171.430 -269.080 -141.430 ;
        RECT -239.080 -171.430 -238.480 -141.430 ;
        RECT -269.680 -173.230 -238.480 -171.430 ;
        RECT -229.680 -141.430 -198.480 -140.830 ;
        RECT -229.680 -171.430 -229.080 -141.430 ;
        RECT -199.080 -171.430 -198.480 -141.430 ;
        RECT -229.680 -173.230 -198.480 -171.430 ;
        RECT -189.680 -141.430 -158.480 -140.830 ;
        RECT -189.680 -171.430 -189.080 -141.430 ;
        RECT -159.080 -171.430 -158.480 -141.430 ;
        RECT -189.680 -173.230 -158.480 -171.430 ;
        RECT -149.680 -141.430 -118.480 -140.830 ;
        RECT -149.680 -171.430 -149.080 -141.430 ;
        RECT -119.080 -171.430 -118.480 -141.430 ;
        RECT -149.680 -173.230 -118.480 -171.430 ;
        RECT -109.680 -141.430 -78.480 -140.830 ;
        RECT -109.680 -171.430 -109.080 -141.430 ;
        RECT -79.080 -171.430 -78.480 -141.430 ;
        RECT -109.680 -173.230 -78.480 -171.430 ;
        RECT -69.680 -141.430 -38.480 -140.830 ;
        RECT -69.680 -171.430 -69.080 -141.430 ;
        RECT -39.080 -171.430 -38.480 -141.430 ;
        RECT -69.680 -173.230 -38.480 -171.430 ;
        RECT -29.680 -141.430 1.520 -140.830 ;
        RECT -29.680 -171.430 -29.080 -141.430 ;
        RECT 0.920 -171.430 1.520 -141.430 ;
        RECT -29.680 -173.230 1.520 -171.430 ;
        RECT 10.320 -141.430 41.520 -140.830 ;
        RECT 10.320 -171.430 10.920 -141.430 ;
        RECT 40.920 -171.430 41.520 -141.430 ;
        RECT 10.320 -173.230 41.520 -171.430 ;
        RECT 50.320 -141.430 81.520 -140.830 ;
        RECT 50.320 -171.430 50.920 -141.430 ;
        RECT 80.920 -171.430 81.520 -141.430 ;
        RECT 50.320 -173.230 81.520 -171.430 ;
        RECT 90.320 -141.430 121.520 -140.830 ;
        RECT 90.320 -171.430 90.920 -141.430 ;
        RECT 120.920 -171.430 121.520 -141.430 ;
        RECT 90.320 -173.230 121.520 -171.430 ;
        RECT 130.320 -141.430 161.520 -140.830 ;
        RECT 130.320 -171.430 130.920 -141.430 ;
        RECT 160.920 -171.430 161.520 -141.430 ;
        RECT 130.320 -173.230 161.520 -171.430 ;
        RECT 170.320 -141.430 201.520 -140.830 ;
        RECT 170.320 -171.430 170.920 -141.430 ;
        RECT 200.920 -171.430 201.520 -141.430 ;
        RECT 170.320 -173.230 201.520 -171.430 ;
        RECT 225.920 -141.430 257.120 -140.830 ;
        RECT 225.920 -171.430 226.520 -141.430 ;
        RECT 256.520 -171.430 257.120 -141.430 ;
        RECT 225.920 -173.230 257.120 -171.430 ;
        RECT 265.920 -141.430 297.120 -140.830 ;
        RECT 265.920 -171.430 266.520 -141.430 ;
        RECT 296.520 -171.430 297.120 -141.430 ;
        RECT 265.920 -173.230 297.120 -171.430 ;
        RECT 305.920 -141.430 337.120 -140.830 ;
        RECT 305.920 -171.430 306.520 -141.430 ;
        RECT 336.520 -171.430 337.120 -141.430 ;
        RECT 305.920 -173.230 337.120 -171.430 ;
        RECT 345.920 -141.430 377.120 -140.830 ;
        RECT 345.920 -171.430 346.520 -141.430 ;
        RECT 376.520 -171.430 377.120 -141.430 ;
        RECT 345.920 -173.230 377.120 -171.430 ;
        RECT 385.920 -141.430 417.120 -140.830 ;
        RECT 385.920 -171.430 386.520 -141.430 ;
        RECT 416.520 -171.430 417.120 -141.430 ;
        RECT 385.920 -173.230 417.120 -171.430 ;
        RECT 425.920 -141.430 457.120 -140.830 ;
        RECT 425.920 -171.430 426.520 -141.430 ;
        RECT 456.520 -171.430 457.120 -141.430 ;
        RECT 425.920 -173.230 457.120 -171.430 ;
        RECT 465.920 -141.430 497.120 -140.830 ;
        RECT 465.920 -171.430 466.520 -141.430 ;
        RECT 496.520 -171.430 497.120 -141.430 ;
        RECT 465.920 -173.230 497.120 -171.430 ;
        RECT 763.320 -172.480 841.320 -132.620 ;
        RECT -533.380 -220.920 -430.980 -220.320 ;
        RECT -533.380 -320.920 -532.780 -220.920 ;
        RECT -432.780 -320.920 -430.980 -220.920 ;
        RECT -533.380 -321.520 -430.980 -320.920 ;
        RECT -425.980 -220.920 -323.580 -220.320 ;
        RECT -425.980 -320.920 -424.180 -220.920 ;
        RECT -324.180 -320.920 -323.580 -220.920 ;
        RECT -425.980 -321.520 -323.580 -320.920 ;
        RECT -318.380 -220.920 -215.980 -220.320 ;
        RECT -318.380 -320.920 -317.780 -220.920 ;
        RECT -217.780 -320.920 -215.980 -220.920 ;
        RECT -318.380 -321.520 -215.980 -320.920 ;
        RECT -210.980 -220.920 -108.580 -220.320 ;
        RECT -210.980 -320.920 -209.180 -220.920 ;
        RECT -109.180 -320.920 -108.580 -220.920 ;
        RECT -210.980 -321.520 -108.580 -320.920 ;
        RECT -103.380 -220.920 -0.980 -220.320 ;
        RECT -103.380 -320.920 -102.780 -220.920 ;
        RECT -2.780 -320.920 -0.980 -220.920 ;
        RECT -103.380 -321.520 -0.980 -320.920 ;
        RECT 4.020 -220.920 106.420 -220.320 ;
        RECT 4.020 -320.920 5.820 -220.920 ;
        RECT 105.820 -320.920 106.420 -220.920 ;
        RECT 4.020 -321.520 106.420 -320.920 ;
        RECT 111.620 -220.920 214.020 -220.320 ;
        RECT 111.620 -320.920 112.220 -220.920 ;
        RECT 212.220 -320.920 214.020 -220.920 ;
        RECT 111.620 -321.520 214.020 -320.920 ;
        RECT 219.020 -220.920 321.420 -220.320 ;
        RECT 219.020 -320.920 220.820 -220.920 ;
        RECT 320.820 -320.920 321.420 -220.920 ;
        RECT 219.020 -321.520 321.420 -320.920 ;
        RECT 326.620 -220.920 429.020 -220.320 ;
        RECT 326.620 -320.920 327.220 -220.920 ;
        RECT 427.220 -320.920 429.020 -220.920 ;
        RECT 326.620 -321.520 429.020 -320.920 ;
        RECT 434.020 -220.920 536.420 -220.320 ;
        RECT 434.020 -320.920 435.820 -220.920 ;
        RECT 535.820 -320.920 536.420 -220.920 ;
        RECT 434.020 -321.520 536.420 -320.920 ;
        RECT 546.520 -352.720 841.320 -172.480 ;
        RECT -838.480 -1085.700 -760.480 -352.720 ;
        RECT -557.530 -390.220 -525.130 -389.620 ;
        RECT -557.530 -420.220 -556.930 -390.220 ;
        RECT -526.930 -420.220 -525.130 -390.220 ;
        RECT -557.530 -420.820 -525.130 -420.220 ;
        RECT -521.830 -390.220 -489.430 -389.620 ;
        RECT -521.830 -420.220 -520.030 -390.220 ;
        RECT -490.030 -420.220 -489.430 -390.220 ;
        RECT -521.830 -420.820 -489.430 -420.220 ;
        RECT -482.530 -390.220 -450.130 -389.620 ;
        RECT -482.530 -420.220 -481.930 -390.220 ;
        RECT -451.930 -420.220 -450.130 -390.220 ;
        RECT -482.530 -420.820 -450.130 -420.220 ;
        RECT -446.830 -390.220 -414.430 -389.620 ;
        RECT -446.830 -420.220 -445.030 -390.220 ;
        RECT -415.030 -420.220 -414.430 -390.220 ;
        RECT -446.830 -420.820 -414.430 -420.220 ;
        RECT -407.530 -390.220 -375.130 -389.620 ;
        RECT -407.530 -420.220 -406.930 -390.220 ;
        RECT -376.930 -420.220 -375.130 -390.220 ;
        RECT -407.530 -420.820 -375.130 -420.220 ;
        RECT -371.830 -390.220 -339.430 -389.620 ;
        RECT -371.830 -420.220 -370.030 -390.220 ;
        RECT -340.030 -420.220 -339.430 -390.220 ;
        RECT -371.830 -420.820 -339.430 -420.220 ;
        RECT -332.530 -390.220 -300.130 -389.620 ;
        RECT -332.530 -420.220 -331.930 -390.220 ;
        RECT -301.930 -420.220 -300.130 -390.220 ;
        RECT -332.530 -420.820 -300.130 -420.220 ;
        RECT -296.830 -390.220 -264.430 -389.620 ;
        RECT -296.830 -420.220 -295.030 -390.220 ;
        RECT -265.030 -420.220 -264.430 -390.220 ;
        RECT -296.830 -420.820 -264.430 -420.220 ;
        RECT -257.530 -390.220 -225.130 -389.620 ;
        RECT -257.530 -420.220 -256.930 -390.220 ;
        RECT -226.930 -420.220 -225.130 -390.220 ;
        RECT -257.530 -420.820 -225.130 -420.220 ;
        RECT -221.830 -390.220 -189.430 -389.620 ;
        RECT -221.830 -420.220 -220.030 -390.220 ;
        RECT -190.030 -420.220 -189.430 -390.220 ;
        RECT -221.830 -420.820 -189.430 -420.220 ;
        RECT -182.530 -390.220 -150.130 -389.620 ;
        RECT -182.530 -420.220 -181.930 -390.220 ;
        RECT -151.930 -420.220 -150.130 -390.220 ;
        RECT -182.530 -420.820 -150.130 -420.220 ;
        RECT -146.830 -390.220 -114.430 -389.620 ;
        RECT -146.830 -420.220 -145.030 -390.220 ;
        RECT -115.030 -420.220 -114.430 -390.220 ;
        RECT -146.830 -420.820 -114.430 -420.220 ;
        RECT -107.530 -390.220 -75.130 -389.620 ;
        RECT -107.530 -420.220 -106.930 -390.220 ;
        RECT -76.930 -420.220 -75.130 -390.220 ;
        RECT -107.530 -420.820 -75.130 -420.220 ;
        RECT -71.830 -390.220 -39.430 -389.620 ;
        RECT -71.830 -420.220 -70.030 -390.220 ;
        RECT -40.030 -420.220 -39.430 -390.220 ;
        RECT -71.830 -420.820 -39.430 -420.220 ;
        RECT -32.530 -390.220 -0.130 -389.620 ;
        RECT -32.530 -420.220 -31.930 -390.220 ;
        RECT -1.930 -420.220 -0.130 -390.220 ;
        RECT -32.530 -420.820 -0.130 -420.220 ;
        RECT 3.170 -390.220 35.570 -389.620 ;
        RECT 3.170 -420.220 4.970 -390.220 ;
        RECT 34.970 -420.220 35.570 -390.220 ;
        RECT 3.170 -420.820 35.570 -420.220 ;
        RECT 42.470 -390.220 74.870 -389.620 ;
        RECT 42.470 -420.220 43.070 -390.220 ;
        RECT 73.070 -420.220 74.870 -390.220 ;
        RECT 42.470 -420.820 74.870 -420.220 ;
        RECT 78.170 -390.220 110.570 -389.620 ;
        RECT 78.170 -420.220 79.970 -390.220 ;
        RECT 109.970 -420.220 110.570 -390.220 ;
        RECT 78.170 -420.820 110.570 -420.220 ;
        RECT 117.470 -390.220 149.870 -389.620 ;
        RECT 117.470 -420.220 118.070 -390.220 ;
        RECT 148.070 -420.220 149.870 -390.220 ;
        RECT 117.470 -420.820 149.870 -420.220 ;
        RECT 153.170 -390.220 185.570 -389.620 ;
        RECT 153.170 -420.220 154.970 -390.220 ;
        RECT 184.970 -420.220 185.570 -390.220 ;
        RECT 153.170 -420.820 185.570 -420.220 ;
        RECT 192.470 -390.220 224.870 -389.620 ;
        RECT 192.470 -420.220 193.070 -390.220 ;
        RECT 223.070 -420.220 224.870 -390.220 ;
        RECT 192.470 -420.820 224.870 -420.220 ;
        RECT 228.170 -390.220 260.570 -389.620 ;
        RECT 228.170 -420.220 229.970 -390.220 ;
        RECT 259.970 -420.220 260.570 -390.220 ;
        RECT 228.170 -420.820 260.570 -420.220 ;
        RECT 267.470 -390.220 299.870 -389.620 ;
        RECT 267.470 -420.220 268.070 -390.220 ;
        RECT 298.070 -420.220 299.870 -390.220 ;
        RECT 267.470 -420.820 299.870 -420.220 ;
        RECT 303.170 -390.220 335.570 -389.620 ;
        RECT 303.170 -420.220 304.970 -390.220 ;
        RECT 334.970 -420.220 335.570 -390.220 ;
        RECT 303.170 -420.820 335.570 -420.220 ;
        RECT 342.470 -390.220 374.870 -389.620 ;
        RECT 342.470 -420.220 343.070 -390.220 ;
        RECT 373.070 -420.220 374.870 -390.220 ;
        RECT 342.470 -420.820 374.870 -420.220 ;
        RECT 378.170 -390.220 410.570 -389.620 ;
        RECT 378.170 -420.220 379.970 -390.220 ;
        RECT 409.970 -420.220 410.570 -390.220 ;
        RECT 378.170 -420.820 410.570 -420.220 ;
        RECT 417.470 -390.220 449.870 -389.620 ;
        RECT 417.470 -420.220 418.070 -390.220 ;
        RECT 448.070 -420.220 449.870 -390.220 ;
        RECT 417.470 -420.820 449.870 -420.220 ;
        RECT 453.170 -390.220 485.570 -389.620 ;
        RECT 453.170 -420.220 454.970 -390.220 ;
        RECT 484.970 -420.220 485.570 -390.220 ;
        RECT 453.170 -420.820 485.570 -420.220 ;
        RECT 492.470 -390.220 524.870 -389.620 ;
        RECT 492.470 -420.220 493.070 -390.220 ;
        RECT 523.070 -420.220 524.870 -390.220 ;
        RECT 492.470 -420.820 524.870 -420.220 ;
        RECT 528.170 -390.220 560.570 -389.620 ;
        RECT 528.170 -420.220 529.970 -390.220 ;
        RECT 559.970 -420.220 560.570 -390.220 ;
        RECT 528.170 -420.820 560.570 -420.220 ;
        RECT -557.530 -425.220 -525.130 -424.620 ;
        RECT -557.530 -455.220 -556.930 -425.220 ;
        RECT -526.930 -455.220 -525.130 -425.220 ;
        RECT -557.530 -455.820 -525.130 -455.220 ;
        RECT -521.830 -425.220 -489.430 -424.620 ;
        RECT -521.830 -455.220 -520.030 -425.220 ;
        RECT -490.030 -455.220 -489.430 -425.220 ;
        RECT -521.830 -455.820 -489.430 -455.220 ;
        RECT -482.530 -425.220 -450.130 -424.620 ;
        RECT -482.530 -455.220 -481.930 -425.220 ;
        RECT -451.930 -455.220 -450.130 -425.220 ;
        RECT -482.530 -455.820 -450.130 -455.220 ;
        RECT -446.830 -425.220 -414.430 -424.620 ;
        RECT -446.830 -455.220 -445.030 -425.220 ;
        RECT -415.030 -455.220 -414.430 -425.220 ;
        RECT -446.830 -455.820 -414.430 -455.220 ;
        RECT -407.530 -425.220 -375.130 -424.620 ;
        RECT -407.530 -455.220 -406.930 -425.220 ;
        RECT -376.930 -455.220 -375.130 -425.220 ;
        RECT -407.530 -455.820 -375.130 -455.220 ;
        RECT -371.830 -425.220 -339.430 -424.620 ;
        RECT -371.830 -455.220 -370.030 -425.220 ;
        RECT -340.030 -455.220 -339.430 -425.220 ;
        RECT -371.830 -455.820 -339.430 -455.220 ;
        RECT -332.530 -425.220 -300.130 -424.620 ;
        RECT -332.530 -455.220 -331.930 -425.220 ;
        RECT -301.930 -455.220 -300.130 -425.220 ;
        RECT -332.530 -455.820 -300.130 -455.220 ;
        RECT -296.830 -425.220 -264.430 -424.620 ;
        RECT -296.830 -455.220 -295.030 -425.220 ;
        RECT -265.030 -455.220 -264.430 -425.220 ;
        RECT -296.830 -455.820 -264.430 -455.220 ;
        RECT -257.530 -425.220 -225.130 -424.620 ;
        RECT -257.530 -455.220 -256.930 -425.220 ;
        RECT -226.930 -455.220 -225.130 -425.220 ;
        RECT -257.530 -455.820 -225.130 -455.220 ;
        RECT -221.830 -425.220 -189.430 -424.620 ;
        RECT -221.830 -455.220 -220.030 -425.220 ;
        RECT -190.030 -455.220 -189.430 -425.220 ;
        RECT -221.830 -455.820 -189.430 -455.220 ;
        RECT -182.530 -425.220 -150.130 -424.620 ;
        RECT -182.530 -455.220 -181.930 -425.220 ;
        RECT -151.930 -455.220 -150.130 -425.220 ;
        RECT -182.530 -455.820 -150.130 -455.220 ;
        RECT -146.830 -425.220 -114.430 -424.620 ;
        RECT -146.830 -455.220 -145.030 -425.220 ;
        RECT -115.030 -455.220 -114.430 -425.220 ;
        RECT -146.830 -455.820 -114.430 -455.220 ;
        RECT -107.530 -425.220 -75.130 -424.620 ;
        RECT -107.530 -455.220 -106.930 -425.220 ;
        RECT -76.930 -455.220 -75.130 -425.220 ;
        RECT -107.530 -455.820 -75.130 -455.220 ;
        RECT -71.830 -425.220 -39.430 -424.620 ;
        RECT -71.830 -455.220 -70.030 -425.220 ;
        RECT -40.030 -455.220 -39.430 -425.220 ;
        RECT -71.830 -455.820 -39.430 -455.220 ;
        RECT -32.530 -425.220 -0.130 -424.620 ;
        RECT -32.530 -455.220 -31.930 -425.220 ;
        RECT -1.930 -455.220 -0.130 -425.220 ;
        RECT -32.530 -455.820 -0.130 -455.220 ;
        RECT 3.170 -425.220 35.570 -424.620 ;
        RECT 3.170 -455.220 4.970 -425.220 ;
        RECT 34.970 -455.220 35.570 -425.220 ;
        RECT 3.170 -455.820 35.570 -455.220 ;
        RECT 42.470 -425.220 74.870 -424.620 ;
        RECT 42.470 -455.220 43.070 -425.220 ;
        RECT 73.070 -455.220 74.870 -425.220 ;
        RECT 42.470 -455.820 74.870 -455.220 ;
        RECT 78.170 -425.220 110.570 -424.620 ;
        RECT 78.170 -455.220 79.970 -425.220 ;
        RECT 109.970 -455.220 110.570 -425.220 ;
        RECT 78.170 -455.820 110.570 -455.220 ;
        RECT 117.470 -425.220 149.870 -424.620 ;
        RECT 117.470 -455.220 118.070 -425.220 ;
        RECT 148.070 -455.220 149.870 -425.220 ;
        RECT 117.470 -455.820 149.870 -455.220 ;
        RECT 153.170 -425.220 185.570 -424.620 ;
        RECT 153.170 -455.220 154.970 -425.220 ;
        RECT 184.970 -455.220 185.570 -425.220 ;
        RECT 153.170 -455.820 185.570 -455.220 ;
        RECT 192.470 -425.220 224.870 -424.620 ;
        RECT 192.470 -455.220 193.070 -425.220 ;
        RECT 223.070 -455.220 224.870 -425.220 ;
        RECT 192.470 -455.820 224.870 -455.220 ;
        RECT 228.170 -425.220 260.570 -424.620 ;
        RECT 228.170 -455.220 229.970 -425.220 ;
        RECT 259.970 -455.220 260.570 -425.220 ;
        RECT 228.170 -455.820 260.570 -455.220 ;
        RECT 267.470 -425.220 299.870 -424.620 ;
        RECT 267.470 -455.220 268.070 -425.220 ;
        RECT 298.070 -455.220 299.870 -425.220 ;
        RECT 267.470 -455.820 299.870 -455.220 ;
        RECT 303.170 -425.220 335.570 -424.620 ;
        RECT 303.170 -455.220 304.970 -425.220 ;
        RECT 334.970 -455.220 335.570 -425.220 ;
        RECT 303.170 -455.820 335.570 -455.220 ;
        RECT 342.470 -425.220 374.870 -424.620 ;
        RECT 342.470 -455.220 343.070 -425.220 ;
        RECT 373.070 -455.220 374.870 -425.220 ;
        RECT 342.470 -455.820 374.870 -455.220 ;
        RECT 378.170 -425.220 410.570 -424.620 ;
        RECT 378.170 -455.220 379.970 -425.220 ;
        RECT 409.970 -455.220 410.570 -425.220 ;
        RECT 378.170 -455.820 410.570 -455.220 ;
        RECT 417.470 -425.220 449.870 -424.620 ;
        RECT 417.470 -455.220 418.070 -425.220 ;
        RECT 448.070 -455.220 449.870 -425.220 ;
        RECT 417.470 -455.820 449.870 -455.220 ;
        RECT 453.170 -425.220 485.570 -424.620 ;
        RECT 453.170 -455.220 454.970 -425.220 ;
        RECT 484.970 -455.220 485.570 -425.220 ;
        RECT 453.170 -455.820 485.570 -455.220 ;
        RECT 492.470 -425.220 524.870 -424.620 ;
        RECT 492.470 -455.220 493.070 -425.220 ;
        RECT 523.070 -455.220 524.870 -425.220 ;
        RECT 492.470 -455.820 524.870 -455.220 ;
        RECT 528.170 -425.220 560.570 -424.620 ;
        RECT 528.170 -455.220 529.970 -425.220 ;
        RECT 559.970 -455.220 560.570 -425.220 ;
        RECT 528.170 -455.820 560.570 -455.220 ;
        RECT -557.530 -460.220 -525.130 -459.620 ;
        RECT -557.530 -490.220 -556.930 -460.220 ;
        RECT -526.930 -490.220 -525.130 -460.220 ;
        RECT -557.530 -490.820 -525.130 -490.220 ;
        RECT -521.830 -460.220 -489.430 -459.620 ;
        RECT -521.830 -490.220 -520.030 -460.220 ;
        RECT -490.030 -490.220 -489.430 -460.220 ;
        RECT -521.830 -490.820 -489.430 -490.220 ;
        RECT -482.530 -460.220 -450.130 -459.620 ;
        RECT -482.530 -490.220 -481.930 -460.220 ;
        RECT -451.930 -490.220 -450.130 -460.220 ;
        RECT -482.530 -490.820 -450.130 -490.220 ;
        RECT -446.830 -460.220 -414.430 -459.620 ;
        RECT -446.830 -490.220 -445.030 -460.220 ;
        RECT -415.030 -490.220 -414.430 -460.220 ;
        RECT -446.830 -490.820 -414.430 -490.220 ;
        RECT -407.530 -460.220 -375.130 -459.620 ;
        RECT -407.530 -490.220 -406.930 -460.220 ;
        RECT -376.930 -490.220 -375.130 -460.220 ;
        RECT -407.530 -490.820 -375.130 -490.220 ;
        RECT -371.830 -460.220 -339.430 -459.620 ;
        RECT -371.830 -490.220 -370.030 -460.220 ;
        RECT -340.030 -490.220 -339.430 -460.220 ;
        RECT -371.830 -490.820 -339.430 -490.220 ;
        RECT -332.530 -460.220 -300.130 -459.620 ;
        RECT -332.530 -490.220 -331.930 -460.220 ;
        RECT -301.930 -490.220 -300.130 -460.220 ;
        RECT -332.530 -490.820 -300.130 -490.220 ;
        RECT -296.830 -460.220 -264.430 -459.620 ;
        RECT -296.830 -490.220 -295.030 -460.220 ;
        RECT -265.030 -490.220 -264.430 -460.220 ;
        RECT -296.830 -490.820 -264.430 -490.220 ;
        RECT -257.530 -460.220 -225.130 -459.620 ;
        RECT -257.530 -490.220 -256.930 -460.220 ;
        RECT -226.930 -490.220 -225.130 -460.220 ;
        RECT -257.530 -490.820 -225.130 -490.220 ;
        RECT -221.830 -460.220 -189.430 -459.620 ;
        RECT -221.830 -490.220 -220.030 -460.220 ;
        RECT -190.030 -490.220 -189.430 -460.220 ;
        RECT -221.830 -490.820 -189.430 -490.220 ;
        RECT -182.530 -460.220 -150.130 -459.620 ;
        RECT -182.530 -490.220 -181.930 -460.220 ;
        RECT -151.930 -490.220 -150.130 -460.220 ;
        RECT -182.530 -490.820 -150.130 -490.220 ;
        RECT -146.830 -460.220 -114.430 -459.620 ;
        RECT -146.830 -490.220 -145.030 -460.220 ;
        RECT -115.030 -490.220 -114.430 -460.220 ;
        RECT -146.830 -490.820 -114.430 -490.220 ;
        RECT -107.530 -460.220 -75.130 -459.620 ;
        RECT -107.530 -490.220 -106.930 -460.220 ;
        RECT -76.930 -490.220 -75.130 -460.220 ;
        RECT -107.530 -490.820 -75.130 -490.220 ;
        RECT -71.830 -460.220 -39.430 -459.620 ;
        RECT -71.830 -490.220 -70.030 -460.220 ;
        RECT -40.030 -490.220 -39.430 -460.220 ;
        RECT -71.830 -490.820 -39.430 -490.220 ;
        RECT -32.530 -460.220 -0.130 -459.620 ;
        RECT -32.530 -490.220 -31.930 -460.220 ;
        RECT -1.930 -490.220 -0.130 -460.220 ;
        RECT -32.530 -490.820 -0.130 -490.220 ;
        RECT 3.170 -460.220 35.570 -459.620 ;
        RECT 3.170 -490.220 4.970 -460.220 ;
        RECT 34.970 -490.220 35.570 -460.220 ;
        RECT 3.170 -490.820 35.570 -490.220 ;
        RECT 42.470 -460.220 74.870 -459.620 ;
        RECT 42.470 -490.220 43.070 -460.220 ;
        RECT 73.070 -490.220 74.870 -460.220 ;
        RECT 42.470 -490.820 74.870 -490.220 ;
        RECT 78.170 -460.220 110.570 -459.620 ;
        RECT 78.170 -490.220 79.970 -460.220 ;
        RECT 109.970 -490.220 110.570 -460.220 ;
        RECT 78.170 -490.820 110.570 -490.220 ;
        RECT 117.470 -460.220 149.870 -459.620 ;
        RECT 117.470 -490.220 118.070 -460.220 ;
        RECT 148.070 -490.220 149.870 -460.220 ;
        RECT 117.470 -490.820 149.870 -490.220 ;
        RECT 153.170 -460.220 185.570 -459.620 ;
        RECT 153.170 -490.220 154.970 -460.220 ;
        RECT 184.970 -490.220 185.570 -460.220 ;
        RECT 153.170 -490.820 185.570 -490.220 ;
        RECT 192.470 -460.220 224.870 -459.620 ;
        RECT 192.470 -490.220 193.070 -460.220 ;
        RECT 223.070 -490.220 224.870 -460.220 ;
        RECT 192.470 -490.820 224.870 -490.220 ;
        RECT 228.170 -460.220 260.570 -459.620 ;
        RECT 228.170 -490.220 229.970 -460.220 ;
        RECT 259.970 -490.220 260.570 -460.220 ;
        RECT 228.170 -490.820 260.570 -490.220 ;
        RECT 267.470 -460.220 299.870 -459.620 ;
        RECT 267.470 -490.220 268.070 -460.220 ;
        RECT 298.070 -490.220 299.870 -460.220 ;
        RECT 267.470 -490.820 299.870 -490.220 ;
        RECT 303.170 -460.220 335.570 -459.620 ;
        RECT 303.170 -490.220 304.970 -460.220 ;
        RECT 334.970 -490.220 335.570 -460.220 ;
        RECT 303.170 -490.820 335.570 -490.220 ;
        RECT 342.470 -460.220 374.870 -459.620 ;
        RECT 342.470 -490.220 343.070 -460.220 ;
        RECT 373.070 -490.220 374.870 -460.220 ;
        RECT 342.470 -490.820 374.870 -490.220 ;
        RECT 378.170 -460.220 410.570 -459.620 ;
        RECT 378.170 -490.220 379.970 -460.220 ;
        RECT 409.970 -490.220 410.570 -460.220 ;
        RECT 378.170 -490.820 410.570 -490.220 ;
        RECT 417.470 -460.220 449.870 -459.620 ;
        RECT 417.470 -490.220 418.070 -460.220 ;
        RECT 448.070 -490.220 449.870 -460.220 ;
        RECT 417.470 -490.820 449.870 -490.220 ;
        RECT 453.170 -460.220 485.570 -459.620 ;
        RECT 453.170 -490.220 454.970 -460.220 ;
        RECT 484.970 -490.220 485.570 -460.220 ;
        RECT 453.170 -490.820 485.570 -490.220 ;
        RECT 492.470 -460.220 524.870 -459.620 ;
        RECT 492.470 -490.220 493.070 -460.220 ;
        RECT 523.070 -490.220 524.870 -460.220 ;
        RECT 492.470 -490.820 524.870 -490.220 ;
        RECT 528.170 -460.220 560.570 -459.620 ;
        RECT 528.170 -490.220 529.970 -460.220 ;
        RECT 559.970 -490.220 560.570 -460.220 ;
        RECT 528.170 -490.820 560.570 -490.220 ;
        RECT -557.530 -495.220 -525.130 -494.620 ;
        RECT -557.530 -525.220 -556.930 -495.220 ;
        RECT -526.930 -525.220 -525.130 -495.220 ;
        RECT -557.530 -525.820 -525.130 -525.220 ;
        RECT -521.830 -495.220 -489.430 -494.620 ;
        RECT -521.830 -525.220 -520.030 -495.220 ;
        RECT -490.030 -525.220 -489.430 -495.220 ;
        RECT -521.830 -525.820 -489.430 -525.220 ;
        RECT -482.530 -495.220 -450.130 -494.620 ;
        RECT -482.530 -525.220 -481.930 -495.220 ;
        RECT -451.930 -525.220 -450.130 -495.220 ;
        RECT -482.530 -525.820 -450.130 -525.220 ;
        RECT -446.830 -495.220 -414.430 -494.620 ;
        RECT -446.830 -525.220 -445.030 -495.220 ;
        RECT -415.030 -525.220 -414.430 -495.220 ;
        RECT -446.830 -525.820 -414.430 -525.220 ;
        RECT -407.530 -495.220 -375.130 -494.620 ;
        RECT -407.530 -525.220 -406.930 -495.220 ;
        RECT -376.930 -525.220 -375.130 -495.220 ;
        RECT -407.530 -525.820 -375.130 -525.220 ;
        RECT -371.830 -495.220 -339.430 -494.620 ;
        RECT -371.830 -525.220 -370.030 -495.220 ;
        RECT -340.030 -525.220 -339.430 -495.220 ;
        RECT -371.830 -525.820 -339.430 -525.220 ;
        RECT -332.530 -495.220 -300.130 -494.620 ;
        RECT -332.530 -525.220 -331.930 -495.220 ;
        RECT -301.930 -525.220 -300.130 -495.220 ;
        RECT -332.530 -525.820 -300.130 -525.220 ;
        RECT -296.830 -495.220 -264.430 -494.620 ;
        RECT -296.830 -525.220 -295.030 -495.220 ;
        RECT -265.030 -525.220 -264.430 -495.220 ;
        RECT -296.830 -525.820 -264.430 -525.220 ;
        RECT -257.530 -495.220 -225.130 -494.620 ;
        RECT -257.530 -525.220 -256.930 -495.220 ;
        RECT -226.930 -525.220 -225.130 -495.220 ;
        RECT -257.530 -525.820 -225.130 -525.220 ;
        RECT -221.830 -495.220 -189.430 -494.620 ;
        RECT -221.830 -525.220 -220.030 -495.220 ;
        RECT -190.030 -525.220 -189.430 -495.220 ;
        RECT -221.830 -525.820 -189.430 -525.220 ;
        RECT -182.530 -495.220 -150.130 -494.620 ;
        RECT -182.530 -525.220 -181.930 -495.220 ;
        RECT -151.930 -525.220 -150.130 -495.220 ;
        RECT -182.530 -525.820 -150.130 -525.220 ;
        RECT -146.830 -495.220 -114.430 -494.620 ;
        RECT -146.830 -525.220 -145.030 -495.220 ;
        RECT -115.030 -525.220 -114.430 -495.220 ;
        RECT -146.830 -525.820 -114.430 -525.220 ;
        RECT -107.530 -495.220 -75.130 -494.620 ;
        RECT -107.530 -525.220 -106.930 -495.220 ;
        RECT -76.930 -525.220 -75.130 -495.220 ;
        RECT -107.530 -525.820 -75.130 -525.220 ;
        RECT -71.830 -495.220 -39.430 -494.620 ;
        RECT -71.830 -525.220 -70.030 -495.220 ;
        RECT -40.030 -525.220 -39.430 -495.220 ;
        RECT -71.830 -525.820 -39.430 -525.220 ;
        RECT -32.530 -495.220 -0.130 -494.620 ;
        RECT -32.530 -525.220 -31.930 -495.220 ;
        RECT -1.930 -525.220 -0.130 -495.220 ;
        RECT -32.530 -525.820 -0.130 -525.220 ;
        RECT 3.170 -495.220 35.570 -494.620 ;
        RECT 3.170 -525.220 4.970 -495.220 ;
        RECT 34.970 -525.220 35.570 -495.220 ;
        RECT 3.170 -525.820 35.570 -525.220 ;
        RECT 42.470 -495.220 74.870 -494.620 ;
        RECT 42.470 -525.220 43.070 -495.220 ;
        RECT 73.070 -525.220 74.870 -495.220 ;
        RECT 42.470 -525.820 74.870 -525.220 ;
        RECT 78.170 -495.220 110.570 -494.620 ;
        RECT 78.170 -525.220 79.970 -495.220 ;
        RECT 109.970 -525.220 110.570 -495.220 ;
        RECT 78.170 -525.820 110.570 -525.220 ;
        RECT 117.470 -495.220 149.870 -494.620 ;
        RECT 117.470 -525.220 118.070 -495.220 ;
        RECT 148.070 -525.220 149.870 -495.220 ;
        RECT 117.470 -525.820 149.870 -525.220 ;
        RECT 153.170 -495.220 185.570 -494.620 ;
        RECT 153.170 -525.220 154.970 -495.220 ;
        RECT 184.970 -525.220 185.570 -495.220 ;
        RECT 153.170 -525.820 185.570 -525.220 ;
        RECT 192.470 -495.220 224.870 -494.620 ;
        RECT 192.470 -525.220 193.070 -495.220 ;
        RECT 223.070 -525.220 224.870 -495.220 ;
        RECT 192.470 -525.820 224.870 -525.220 ;
        RECT 228.170 -495.220 260.570 -494.620 ;
        RECT 228.170 -525.220 229.970 -495.220 ;
        RECT 259.970 -525.220 260.570 -495.220 ;
        RECT 228.170 -525.820 260.570 -525.220 ;
        RECT 267.470 -495.220 299.870 -494.620 ;
        RECT 267.470 -525.220 268.070 -495.220 ;
        RECT 298.070 -525.220 299.870 -495.220 ;
        RECT 267.470 -525.820 299.870 -525.220 ;
        RECT 303.170 -495.220 335.570 -494.620 ;
        RECT 303.170 -525.220 304.970 -495.220 ;
        RECT 334.970 -525.220 335.570 -495.220 ;
        RECT 303.170 -525.820 335.570 -525.220 ;
        RECT 342.470 -495.220 374.870 -494.620 ;
        RECT 342.470 -525.220 343.070 -495.220 ;
        RECT 373.070 -525.220 374.870 -495.220 ;
        RECT 342.470 -525.820 374.870 -525.220 ;
        RECT 378.170 -495.220 410.570 -494.620 ;
        RECT 378.170 -525.220 379.970 -495.220 ;
        RECT 409.970 -525.220 410.570 -495.220 ;
        RECT 378.170 -525.820 410.570 -525.220 ;
        RECT 417.470 -495.220 449.870 -494.620 ;
        RECT 417.470 -525.220 418.070 -495.220 ;
        RECT 448.070 -525.220 449.870 -495.220 ;
        RECT 417.470 -525.820 449.870 -525.220 ;
        RECT 453.170 -495.220 485.570 -494.620 ;
        RECT 453.170 -525.220 454.970 -495.220 ;
        RECT 484.970 -525.220 485.570 -495.220 ;
        RECT 453.170 -525.820 485.570 -525.220 ;
        RECT 492.470 -495.220 524.870 -494.620 ;
        RECT 492.470 -525.220 493.070 -495.220 ;
        RECT 523.070 -525.220 524.870 -495.220 ;
        RECT 492.470 -525.820 524.870 -525.220 ;
        RECT 528.170 -495.220 560.570 -494.620 ;
        RECT 528.170 -525.220 529.970 -495.220 ;
        RECT 559.970 -525.220 560.570 -495.220 ;
        RECT 528.170 -525.820 560.570 -525.220 ;
        RECT -557.530 -530.220 -525.130 -529.620 ;
        RECT -557.530 -560.220 -556.930 -530.220 ;
        RECT -526.930 -560.220 -525.130 -530.220 ;
        RECT -557.530 -560.820 -525.130 -560.220 ;
        RECT -521.830 -530.220 -489.430 -529.620 ;
        RECT -521.830 -560.220 -520.030 -530.220 ;
        RECT -490.030 -560.220 -489.430 -530.220 ;
        RECT -521.830 -560.820 -489.430 -560.220 ;
        RECT -482.530 -530.220 -450.130 -529.620 ;
        RECT -482.530 -560.220 -481.930 -530.220 ;
        RECT -451.930 -560.220 -450.130 -530.220 ;
        RECT -482.530 -560.820 -450.130 -560.220 ;
        RECT -446.830 -530.220 -414.430 -529.620 ;
        RECT -446.830 -560.220 -445.030 -530.220 ;
        RECT -415.030 -560.220 -414.430 -530.220 ;
        RECT -446.830 -560.820 -414.430 -560.220 ;
        RECT -407.530 -530.220 -375.130 -529.620 ;
        RECT -407.530 -560.220 -406.930 -530.220 ;
        RECT -376.930 -560.220 -375.130 -530.220 ;
        RECT -407.530 -560.820 -375.130 -560.220 ;
        RECT -371.830 -530.220 -339.430 -529.620 ;
        RECT -371.830 -560.220 -370.030 -530.220 ;
        RECT -340.030 -560.220 -339.430 -530.220 ;
        RECT -371.830 -560.820 -339.430 -560.220 ;
        RECT -332.530 -530.220 -300.130 -529.620 ;
        RECT -332.530 -560.220 -331.930 -530.220 ;
        RECT -301.930 -560.220 -300.130 -530.220 ;
        RECT -332.530 -560.820 -300.130 -560.220 ;
        RECT -296.830 -530.220 -264.430 -529.620 ;
        RECT -296.830 -560.220 -295.030 -530.220 ;
        RECT -265.030 -560.220 -264.430 -530.220 ;
        RECT -296.830 -560.820 -264.430 -560.220 ;
        RECT -257.530 -530.220 -225.130 -529.620 ;
        RECT -257.530 -560.220 -256.930 -530.220 ;
        RECT -226.930 -560.220 -225.130 -530.220 ;
        RECT -257.530 -560.820 -225.130 -560.220 ;
        RECT -221.830 -530.220 -189.430 -529.620 ;
        RECT -221.830 -560.220 -220.030 -530.220 ;
        RECT -190.030 -560.220 -189.430 -530.220 ;
        RECT -221.830 -560.820 -189.430 -560.220 ;
        RECT -182.530 -530.220 -150.130 -529.620 ;
        RECT -182.530 -560.220 -181.930 -530.220 ;
        RECT -151.930 -560.220 -150.130 -530.220 ;
        RECT -182.530 -560.820 -150.130 -560.220 ;
        RECT -146.830 -530.220 -114.430 -529.620 ;
        RECT -146.830 -560.220 -145.030 -530.220 ;
        RECT -115.030 -560.220 -114.430 -530.220 ;
        RECT -146.830 -560.820 -114.430 -560.220 ;
        RECT -107.530 -530.220 -75.130 -529.620 ;
        RECT -107.530 -560.220 -106.930 -530.220 ;
        RECT -76.930 -560.220 -75.130 -530.220 ;
        RECT -107.530 -560.820 -75.130 -560.220 ;
        RECT -71.830 -530.220 -39.430 -529.620 ;
        RECT -71.830 -560.220 -70.030 -530.220 ;
        RECT -40.030 -560.220 -39.430 -530.220 ;
        RECT -71.830 -560.820 -39.430 -560.220 ;
        RECT -32.530 -530.220 -0.130 -529.620 ;
        RECT -32.530 -560.220 -31.930 -530.220 ;
        RECT -1.930 -560.220 -0.130 -530.220 ;
        RECT -32.530 -560.820 -0.130 -560.220 ;
        RECT 3.170 -530.220 35.570 -529.620 ;
        RECT 3.170 -560.220 4.970 -530.220 ;
        RECT 34.970 -560.220 35.570 -530.220 ;
        RECT 3.170 -560.820 35.570 -560.220 ;
        RECT 42.470 -530.220 74.870 -529.620 ;
        RECT 42.470 -560.220 43.070 -530.220 ;
        RECT 73.070 -560.220 74.870 -530.220 ;
        RECT 42.470 -560.820 74.870 -560.220 ;
        RECT 78.170 -530.220 110.570 -529.620 ;
        RECT 78.170 -560.220 79.970 -530.220 ;
        RECT 109.970 -560.220 110.570 -530.220 ;
        RECT 78.170 -560.820 110.570 -560.220 ;
        RECT 117.470 -530.220 149.870 -529.620 ;
        RECT 117.470 -560.220 118.070 -530.220 ;
        RECT 148.070 -560.220 149.870 -530.220 ;
        RECT 117.470 -560.820 149.870 -560.220 ;
        RECT 153.170 -530.220 185.570 -529.620 ;
        RECT 153.170 -560.220 154.970 -530.220 ;
        RECT 184.970 -560.220 185.570 -530.220 ;
        RECT 153.170 -560.820 185.570 -560.220 ;
        RECT 192.470 -530.220 224.870 -529.620 ;
        RECT 192.470 -560.220 193.070 -530.220 ;
        RECT 223.070 -560.220 224.870 -530.220 ;
        RECT 192.470 -560.820 224.870 -560.220 ;
        RECT 228.170 -530.220 260.570 -529.620 ;
        RECT 228.170 -560.220 229.970 -530.220 ;
        RECT 259.970 -560.220 260.570 -530.220 ;
        RECT 228.170 -560.820 260.570 -560.220 ;
        RECT 267.470 -530.220 299.870 -529.620 ;
        RECT 267.470 -560.220 268.070 -530.220 ;
        RECT 298.070 -560.220 299.870 -530.220 ;
        RECT 267.470 -560.820 299.870 -560.220 ;
        RECT 303.170 -530.220 335.570 -529.620 ;
        RECT 303.170 -560.220 304.970 -530.220 ;
        RECT 334.970 -560.220 335.570 -530.220 ;
        RECT 303.170 -560.820 335.570 -560.220 ;
        RECT 342.470 -530.220 374.870 -529.620 ;
        RECT 342.470 -560.220 343.070 -530.220 ;
        RECT 373.070 -560.220 374.870 -530.220 ;
        RECT 342.470 -560.820 374.870 -560.220 ;
        RECT 378.170 -530.220 410.570 -529.620 ;
        RECT 378.170 -560.220 379.970 -530.220 ;
        RECT 409.970 -560.220 410.570 -530.220 ;
        RECT 378.170 -560.820 410.570 -560.220 ;
        RECT 417.470 -530.220 449.870 -529.620 ;
        RECT 417.470 -560.220 418.070 -530.220 ;
        RECT 448.070 -560.220 449.870 -530.220 ;
        RECT 417.470 -560.820 449.870 -560.220 ;
        RECT 453.170 -530.220 485.570 -529.620 ;
        RECT 453.170 -560.220 454.970 -530.220 ;
        RECT 484.970 -560.220 485.570 -530.220 ;
        RECT 453.170 -560.820 485.570 -560.220 ;
        RECT 492.470 -530.220 524.870 -529.620 ;
        RECT 492.470 -560.220 493.070 -530.220 ;
        RECT 523.070 -560.220 524.870 -530.220 ;
        RECT 492.470 -560.820 524.870 -560.220 ;
        RECT 528.170 -530.220 560.570 -529.620 ;
        RECT 528.170 -560.220 529.970 -530.220 ;
        RECT 559.970 -560.220 560.570 -530.220 ;
        RECT 528.170 -560.820 560.570 -560.220 ;
        RECT -557.530 -565.220 -525.130 -564.620 ;
        RECT -557.530 -595.220 -556.930 -565.220 ;
        RECT -526.930 -595.220 -525.130 -565.220 ;
        RECT -557.530 -595.820 -525.130 -595.220 ;
        RECT -521.830 -565.220 -489.430 -564.620 ;
        RECT -521.830 -595.220 -520.030 -565.220 ;
        RECT -490.030 -595.220 -489.430 -565.220 ;
        RECT -521.830 -595.820 -489.430 -595.220 ;
        RECT -482.530 -565.220 -450.130 -564.620 ;
        RECT -482.530 -595.220 -481.930 -565.220 ;
        RECT -451.930 -595.220 -450.130 -565.220 ;
        RECT -482.530 -595.820 -450.130 -595.220 ;
        RECT -446.830 -565.220 -414.430 -564.620 ;
        RECT -446.830 -595.220 -445.030 -565.220 ;
        RECT -415.030 -595.220 -414.430 -565.220 ;
        RECT -446.830 -595.820 -414.430 -595.220 ;
        RECT -407.530 -565.220 -375.130 -564.620 ;
        RECT -407.530 -595.220 -406.930 -565.220 ;
        RECT -376.930 -595.220 -375.130 -565.220 ;
        RECT -407.530 -595.820 -375.130 -595.220 ;
        RECT -371.830 -565.220 -339.430 -564.620 ;
        RECT -371.830 -595.220 -370.030 -565.220 ;
        RECT -340.030 -595.220 -339.430 -565.220 ;
        RECT -371.830 -595.820 -339.430 -595.220 ;
        RECT -332.530 -565.220 -300.130 -564.620 ;
        RECT -332.530 -595.220 -331.930 -565.220 ;
        RECT -301.930 -595.220 -300.130 -565.220 ;
        RECT -332.530 -595.820 -300.130 -595.220 ;
        RECT -296.830 -565.220 -264.430 -564.620 ;
        RECT -296.830 -595.220 -295.030 -565.220 ;
        RECT -265.030 -595.220 -264.430 -565.220 ;
        RECT -296.830 -595.820 -264.430 -595.220 ;
        RECT -257.530 -565.220 -225.130 -564.620 ;
        RECT -257.530 -595.220 -256.930 -565.220 ;
        RECT -226.930 -595.220 -225.130 -565.220 ;
        RECT -257.530 -595.820 -225.130 -595.220 ;
        RECT -221.830 -565.220 -189.430 -564.620 ;
        RECT -221.830 -595.220 -220.030 -565.220 ;
        RECT -190.030 -595.220 -189.430 -565.220 ;
        RECT -221.830 -595.820 -189.430 -595.220 ;
        RECT -182.530 -565.220 -150.130 -564.620 ;
        RECT -182.530 -595.220 -181.930 -565.220 ;
        RECT -151.930 -595.220 -150.130 -565.220 ;
        RECT -182.530 -595.820 -150.130 -595.220 ;
        RECT -146.830 -565.220 -114.430 -564.620 ;
        RECT -146.830 -595.220 -145.030 -565.220 ;
        RECT -115.030 -595.220 -114.430 -565.220 ;
        RECT -146.830 -595.820 -114.430 -595.220 ;
        RECT -107.530 -565.220 -75.130 -564.620 ;
        RECT -107.530 -595.220 -106.930 -565.220 ;
        RECT -76.930 -595.220 -75.130 -565.220 ;
        RECT -107.530 -595.820 -75.130 -595.220 ;
        RECT -71.830 -565.220 -39.430 -564.620 ;
        RECT -71.830 -595.220 -70.030 -565.220 ;
        RECT -40.030 -595.220 -39.430 -565.220 ;
        RECT -71.830 -595.820 -39.430 -595.220 ;
        RECT -32.530 -565.220 -0.130 -564.620 ;
        RECT -32.530 -595.220 -31.930 -565.220 ;
        RECT -1.930 -595.220 -0.130 -565.220 ;
        RECT -32.530 -595.820 -0.130 -595.220 ;
        RECT 3.170 -565.220 35.570 -564.620 ;
        RECT 3.170 -595.220 4.970 -565.220 ;
        RECT 34.970 -595.220 35.570 -565.220 ;
        RECT 3.170 -595.820 35.570 -595.220 ;
        RECT 42.470 -565.220 74.870 -564.620 ;
        RECT 42.470 -595.220 43.070 -565.220 ;
        RECT 73.070 -595.220 74.870 -565.220 ;
        RECT 42.470 -595.820 74.870 -595.220 ;
        RECT 78.170 -565.220 110.570 -564.620 ;
        RECT 78.170 -595.220 79.970 -565.220 ;
        RECT 109.970 -595.220 110.570 -565.220 ;
        RECT 78.170 -595.820 110.570 -595.220 ;
        RECT 117.470 -565.220 149.870 -564.620 ;
        RECT 117.470 -595.220 118.070 -565.220 ;
        RECT 148.070 -595.220 149.870 -565.220 ;
        RECT 117.470 -595.820 149.870 -595.220 ;
        RECT 153.170 -565.220 185.570 -564.620 ;
        RECT 153.170 -595.220 154.970 -565.220 ;
        RECT 184.970 -595.220 185.570 -565.220 ;
        RECT 153.170 -595.820 185.570 -595.220 ;
        RECT 192.470 -565.220 224.870 -564.620 ;
        RECT 192.470 -595.220 193.070 -565.220 ;
        RECT 223.070 -595.220 224.870 -565.220 ;
        RECT 192.470 -595.820 224.870 -595.220 ;
        RECT 228.170 -565.220 260.570 -564.620 ;
        RECT 228.170 -595.220 229.970 -565.220 ;
        RECT 259.970 -595.220 260.570 -565.220 ;
        RECT 228.170 -595.820 260.570 -595.220 ;
        RECT 267.470 -565.220 299.870 -564.620 ;
        RECT 267.470 -595.220 268.070 -565.220 ;
        RECT 298.070 -595.220 299.870 -565.220 ;
        RECT 267.470 -595.820 299.870 -595.220 ;
        RECT 303.170 -565.220 335.570 -564.620 ;
        RECT 303.170 -595.220 304.970 -565.220 ;
        RECT 334.970 -595.220 335.570 -565.220 ;
        RECT 303.170 -595.820 335.570 -595.220 ;
        RECT 342.470 -565.220 374.870 -564.620 ;
        RECT 342.470 -595.220 343.070 -565.220 ;
        RECT 373.070 -595.220 374.870 -565.220 ;
        RECT 342.470 -595.820 374.870 -595.220 ;
        RECT 378.170 -565.220 410.570 -564.620 ;
        RECT 378.170 -595.220 379.970 -565.220 ;
        RECT 409.970 -595.220 410.570 -565.220 ;
        RECT 378.170 -595.820 410.570 -595.220 ;
        RECT 417.470 -565.220 449.870 -564.620 ;
        RECT 417.470 -595.220 418.070 -565.220 ;
        RECT 448.070 -595.220 449.870 -565.220 ;
        RECT 417.470 -595.820 449.870 -595.220 ;
        RECT 453.170 -565.220 485.570 -564.620 ;
        RECT 453.170 -595.220 454.970 -565.220 ;
        RECT 484.970 -595.220 485.570 -565.220 ;
        RECT 453.170 -595.820 485.570 -595.220 ;
        RECT 492.470 -565.220 524.870 -564.620 ;
        RECT 492.470 -595.220 493.070 -565.220 ;
        RECT 523.070 -595.220 524.870 -565.220 ;
        RECT 492.470 -595.820 524.870 -595.220 ;
        RECT 528.170 -565.220 560.570 -564.620 ;
        RECT 528.170 -595.220 529.970 -565.220 ;
        RECT 559.970 -595.220 560.570 -565.220 ;
        RECT 528.170 -595.820 560.570 -595.220 ;
        RECT -557.530 -600.220 -525.130 -599.620 ;
        RECT -557.530 -630.220 -556.930 -600.220 ;
        RECT -526.930 -630.220 -525.130 -600.220 ;
        RECT -557.530 -630.820 -525.130 -630.220 ;
        RECT -521.830 -600.220 -489.430 -599.620 ;
        RECT -521.830 -630.220 -520.030 -600.220 ;
        RECT -490.030 -630.220 -489.430 -600.220 ;
        RECT -521.830 -630.820 -489.430 -630.220 ;
        RECT -482.530 -600.220 -450.130 -599.620 ;
        RECT -482.530 -630.220 -481.930 -600.220 ;
        RECT -451.930 -630.220 -450.130 -600.220 ;
        RECT -482.530 -630.820 -450.130 -630.220 ;
        RECT -446.830 -600.220 -414.430 -599.620 ;
        RECT -446.830 -630.220 -445.030 -600.220 ;
        RECT -415.030 -630.220 -414.430 -600.220 ;
        RECT -446.830 -630.820 -414.430 -630.220 ;
        RECT -407.530 -600.220 -375.130 -599.620 ;
        RECT -407.530 -630.220 -406.930 -600.220 ;
        RECT -376.930 -630.220 -375.130 -600.220 ;
        RECT -407.530 -630.820 -375.130 -630.220 ;
        RECT -371.830 -600.220 -339.430 -599.620 ;
        RECT -371.830 -630.220 -370.030 -600.220 ;
        RECT -340.030 -630.220 -339.430 -600.220 ;
        RECT -371.830 -630.820 -339.430 -630.220 ;
        RECT -332.530 -600.220 -300.130 -599.620 ;
        RECT -332.530 -630.220 -331.930 -600.220 ;
        RECT -301.930 -630.220 -300.130 -600.220 ;
        RECT -332.530 -630.820 -300.130 -630.220 ;
        RECT -296.830 -600.220 -264.430 -599.620 ;
        RECT -296.830 -630.220 -295.030 -600.220 ;
        RECT -265.030 -630.220 -264.430 -600.220 ;
        RECT -296.830 -630.820 -264.430 -630.220 ;
        RECT -257.530 -600.220 -225.130 -599.620 ;
        RECT -257.530 -630.220 -256.930 -600.220 ;
        RECT -226.930 -630.220 -225.130 -600.220 ;
        RECT -257.530 -630.820 -225.130 -630.220 ;
        RECT -221.830 -600.220 -189.430 -599.620 ;
        RECT -221.830 -630.220 -220.030 -600.220 ;
        RECT -190.030 -630.220 -189.430 -600.220 ;
        RECT -221.830 -630.820 -189.430 -630.220 ;
        RECT -182.530 -600.220 -150.130 -599.620 ;
        RECT -182.530 -630.220 -181.930 -600.220 ;
        RECT -151.930 -630.220 -150.130 -600.220 ;
        RECT -182.530 -630.820 -150.130 -630.220 ;
        RECT -146.830 -600.220 -114.430 -599.620 ;
        RECT -146.830 -630.220 -145.030 -600.220 ;
        RECT -115.030 -630.220 -114.430 -600.220 ;
        RECT -146.830 -630.820 -114.430 -630.220 ;
        RECT -107.530 -600.220 -75.130 -599.620 ;
        RECT -107.530 -630.220 -106.930 -600.220 ;
        RECT -76.930 -630.220 -75.130 -600.220 ;
        RECT -107.530 -630.820 -75.130 -630.220 ;
        RECT -71.830 -600.220 -39.430 -599.620 ;
        RECT -71.830 -630.220 -70.030 -600.220 ;
        RECT -40.030 -630.220 -39.430 -600.220 ;
        RECT -71.830 -630.820 -39.430 -630.220 ;
        RECT -32.530 -600.220 -0.130 -599.620 ;
        RECT -32.530 -630.220 -31.930 -600.220 ;
        RECT -1.930 -630.220 -0.130 -600.220 ;
        RECT -32.530 -630.820 -0.130 -630.220 ;
        RECT 3.170 -600.220 35.570 -599.620 ;
        RECT 3.170 -630.220 4.970 -600.220 ;
        RECT 34.970 -630.220 35.570 -600.220 ;
        RECT 3.170 -630.820 35.570 -630.220 ;
        RECT 42.470 -600.220 74.870 -599.620 ;
        RECT 42.470 -630.220 43.070 -600.220 ;
        RECT 73.070 -630.220 74.870 -600.220 ;
        RECT 42.470 -630.820 74.870 -630.220 ;
        RECT 78.170 -600.220 110.570 -599.620 ;
        RECT 78.170 -630.220 79.970 -600.220 ;
        RECT 109.970 -630.220 110.570 -600.220 ;
        RECT 78.170 -630.820 110.570 -630.220 ;
        RECT 117.470 -600.220 149.870 -599.620 ;
        RECT 117.470 -630.220 118.070 -600.220 ;
        RECT 148.070 -630.220 149.870 -600.220 ;
        RECT 117.470 -630.820 149.870 -630.220 ;
        RECT 153.170 -600.220 185.570 -599.620 ;
        RECT 153.170 -630.220 154.970 -600.220 ;
        RECT 184.970 -630.220 185.570 -600.220 ;
        RECT 153.170 -630.820 185.570 -630.220 ;
        RECT 192.470 -600.220 224.870 -599.620 ;
        RECT 192.470 -630.220 193.070 -600.220 ;
        RECT 223.070 -630.220 224.870 -600.220 ;
        RECT 192.470 -630.820 224.870 -630.220 ;
        RECT 228.170 -600.220 260.570 -599.620 ;
        RECT 228.170 -630.220 229.970 -600.220 ;
        RECT 259.970 -630.220 260.570 -600.220 ;
        RECT 228.170 -630.820 260.570 -630.220 ;
        RECT 267.470 -600.220 299.870 -599.620 ;
        RECT 267.470 -630.220 268.070 -600.220 ;
        RECT 298.070 -630.220 299.870 -600.220 ;
        RECT 267.470 -630.820 299.870 -630.220 ;
        RECT 303.170 -600.220 335.570 -599.620 ;
        RECT 303.170 -630.220 304.970 -600.220 ;
        RECT 334.970 -630.220 335.570 -600.220 ;
        RECT 303.170 -630.820 335.570 -630.220 ;
        RECT 342.470 -600.220 374.870 -599.620 ;
        RECT 342.470 -630.220 343.070 -600.220 ;
        RECT 373.070 -630.220 374.870 -600.220 ;
        RECT 342.470 -630.820 374.870 -630.220 ;
        RECT 378.170 -600.220 410.570 -599.620 ;
        RECT 378.170 -630.220 379.970 -600.220 ;
        RECT 409.970 -630.220 410.570 -600.220 ;
        RECT 378.170 -630.820 410.570 -630.220 ;
        RECT 417.470 -600.220 449.870 -599.620 ;
        RECT 417.470 -630.220 418.070 -600.220 ;
        RECT 448.070 -630.220 449.870 -600.220 ;
        RECT 417.470 -630.820 449.870 -630.220 ;
        RECT 453.170 -600.220 485.570 -599.620 ;
        RECT 453.170 -630.220 454.970 -600.220 ;
        RECT 484.970 -630.220 485.570 -600.220 ;
        RECT 453.170 -630.820 485.570 -630.220 ;
        RECT 492.470 -600.220 524.870 -599.620 ;
        RECT 492.470 -630.220 493.070 -600.220 ;
        RECT 523.070 -630.220 524.870 -600.220 ;
        RECT 492.470 -630.820 524.870 -630.220 ;
        RECT 528.170 -600.220 560.570 -599.620 ;
        RECT 528.170 -630.220 529.970 -600.220 ;
        RECT 559.970 -630.220 560.570 -600.220 ;
        RECT 528.170 -630.820 560.570 -630.220 ;
        RECT -557.530 -635.220 -525.130 -634.620 ;
        RECT -557.530 -665.220 -556.930 -635.220 ;
        RECT -526.930 -665.220 -525.130 -635.220 ;
        RECT -557.530 -665.820 -525.130 -665.220 ;
        RECT -521.830 -635.220 -489.430 -634.620 ;
        RECT -521.830 -665.220 -520.030 -635.220 ;
        RECT -490.030 -665.220 -489.430 -635.220 ;
        RECT -521.830 -665.820 -489.430 -665.220 ;
        RECT -482.530 -635.220 -450.130 -634.620 ;
        RECT -482.530 -665.220 -481.930 -635.220 ;
        RECT -451.930 -665.220 -450.130 -635.220 ;
        RECT -482.530 -665.820 -450.130 -665.220 ;
        RECT -446.830 -635.220 -414.430 -634.620 ;
        RECT -446.830 -665.220 -445.030 -635.220 ;
        RECT -415.030 -665.220 -414.430 -635.220 ;
        RECT -446.830 -665.820 -414.430 -665.220 ;
        RECT -407.530 -635.220 -375.130 -634.620 ;
        RECT -407.530 -665.220 -406.930 -635.220 ;
        RECT -376.930 -665.220 -375.130 -635.220 ;
        RECT -407.530 -665.820 -375.130 -665.220 ;
        RECT -371.830 -635.220 -339.430 -634.620 ;
        RECT -371.830 -665.220 -370.030 -635.220 ;
        RECT -340.030 -665.220 -339.430 -635.220 ;
        RECT -371.830 -665.820 -339.430 -665.220 ;
        RECT -332.530 -635.220 -300.130 -634.620 ;
        RECT -332.530 -665.220 -331.930 -635.220 ;
        RECT -301.930 -665.220 -300.130 -635.220 ;
        RECT -332.530 -665.820 -300.130 -665.220 ;
        RECT -296.830 -635.220 -264.430 -634.620 ;
        RECT -296.830 -665.220 -295.030 -635.220 ;
        RECT -265.030 -665.220 -264.430 -635.220 ;
        RECT -296.830 -665.820 -264.430 -665.220 ;
        RECT -257.530 -635.220 -225.130 -634.620 ;
        RECT -257.530 -665.220 -256.930 -635.220 ;
        RECT -226.930 -665.220 -225.130 -635.220 ;
        RECT -257.530 -665.820 -225.130 -665.220 ;
        RECT -221.830 -635.220 -189.430 -634.620 ;
        RECT -221.830 -665.220 -220.030 -635.220 ;
        RECT -190.030 -665.220 -189.430 -635.220 ;
        RECT -221.830 -665.820 -189.430 -665.220 ;
        RECT -182.530 -635.220 -150.130 -634.620 ;
        RECT -182.530 -665.220 -181.930 -635.220 ;
        RECT -151.930 -665.220 -150.130 -635.220 ;
        RECT -182.530 -665.820 -150.130 -665.220 ;
        RECT -146.830 -635.220 -114.430 -634.620 ;
        RECT -146.830 -665.220 -145.030 -635.220 ;
        RECT -115.030 -665.220 -114.430 -635.220 ;
        RECT -146.830 -665.820 -114.430 -665.220 ;
        RECT -107.530 -635.220 -75.130 -634.620 ;
        RECT -107.530 -665.220 -106.930 -635.220 ;
        RECT -76.930 -665.220 -75.130 -635.220 ;
        RECT -107.530 -665.820 -75.130 -665.220 ;
        RECT -71.830 -635.220 -39.430 -634.620 ;
        RECT -71.830 -665.220 -70.030 -635.220 ;
        RECT -40.030 -665.220 -39.430 -635.220 ;
        RECT -71.830 -665.820 -39.430 -665.220 ;
        RECT -32.530 -635.220 -0.130 -634.620 ;
        RECT -32.530 -665.220 -31.930 -635.220 ;
        RECT -1.930 -665.220 -0.130 -635.220 ;
        RECT -32.530 -665.820 -0.130 -665.220 ;
        RECT 3.170 -635.220 35.570 -634.620 ;
        RECT 3.170 -665.220 4.970 -635.220 ;
        RECT 34.970 -665.220 35.570 -635.220 ;
        RECT 3.170 -665.820 35.570 -665.220 ;
        RECT 42.470 -635.220 74.870 -634.620 ;
        RECT 42.470 -665.220 43.070 -635.220 ;
        RECT 73.070 -665.220 74.870 -635.220 ;
        RECT 42.470 -665.820 74.870 -665.220 ;
        RECT 78.170 -635.220 110.570 -634.620 ;
        RECT 78.170 -665.220 79.970 -635.220 ;
        RECT 109.970 -665.220 110.570 -635.220 ;
        RECT 78.170 -665.820 110.570 -665.220 ;
        RECT 117.470 -635.220 149.870 -634.620 ;
        RECT 117.470 -665.220 118.070 -635.220 ;
        RECT 148.070 -665.220 149.870 -635.220 ;
        RECT 117.470 -665.820 149.870 -665.220 ;
        RECT 153.170 -635.220 185.570 -634.620 ;
        RECT 153.170 -665.220 154.970 -635.220 ;
        RECT 184.970 -665.220 185.570 -635.220 ;
        RECT 153.170 -665.820 185.570 -665.220 ;
        RECT 192.470 -635.220 224.870 -634.620 ;
        RECT 192.470 -665.220 193.070 -635.220 ;
        RECT 223.070 -665.220 224.870 -635.220 ;
        RECT 192.470 -665.820 224.870 -665.220 ;
        RECT 228.170 -635.220 260.570 -634.620 ;
        RECT 228.170 -665.220 229.970 -635.220 ;
        RECT 259.970 -665.220 260.570 -635.220 ;
        RECT 228.170 -665.820 260.570 -665.220 ;
        RECT 267.470 -635.220 299.870 -634.620 ;
        RECT 267.470 -665.220 268.070 -635.220 ;
        RECT 298.070 -665.220 299.870 -635.220 ;
        RECT 267.470 -665.820 299.870 -665.220 ;
        RECT 303.170 -635.220 335.570 -634.620 ;
        RECT 303.170 -665.220 304.970 -635.220 ;
        RECT 334.970 -665.220 335.570 -635.220 ;
        RECT 303.170 -665.820 335.570 -665.220 ;
        RECT 342.470 -635.220 374.870 -634.620 ;
        RECT 342.470 -665.220 343.070 -635.220 ;
        RECT 373.070 -665.220 374.870 -635.220 ;
        RECT 342.470 -665.820 374.870 -665.220 ;
        RECT 378.170 -635.220 410.570 -634.620 ;
        RECT 378.170 -665.220 379.970 -635.220 ;
        RECT 409.970 -665.220 410.570 -635.220 ;
        RECT 378.170 -665.820 410.570 -665.220 ;
        RECT 417.470 -635.220 449.870 -634.620 ;
        RECT 417.470 -665.220 418.070 -635.220 ;
        RECT 448.070 -665.220 449.870 -635.220 ;
        RECT 417.470 -665.820 449.870 -665.220 ;
        RECT 453.170 -635.220 485.570 -634.620 ;
        RECT 453.170 -665.220 454.970 -635.220 ;
        RECT 484.970 -665.220 485.570 -635.220 ;
        RECT 453.170 -665.820 485.570 -665.220 ;
        RECT 492.470 -635.220 524.870 -634.620 ;
        RECT 492.470 -665.220 493.070 -635.220 ;
        RECT 523.070 -665.220 524.870 -635.220 ;
        RECT 492.470 -665.820 524.870 -665.220 ;
        RECT 528.170 -635.220 560.570 -634.620 ;
        RECT 528.170 -665.220 529.970 -635.220 ;
        RECT 559.970 -665.220 560.570 -635.220 ;
        RECT 528.170 -665.820 560.570 -665.220 ;
        RECT -557.530 -670.220 -525.130 -669.620 ;
        RECT -557.530 -700.220 -556.930 -670.220 ;
        RECT -526.930 -700.220 -525.130 -670.220 ;
        RECT -557.530 -700.820 -525.130 -700.220 ;
        RECT -521.830 -670.220 -489.430 -669.620 ;
        RECT -521.830 -700.220 -520.030 -670.220 ;
        RECT -490.030 -700.220 -489.430 -670.220 ;
        RECT -521.830 -700.820 -489.430 -700.220 ;
        RECT -482.530 -670.220 -450.130 -669.620 ;
        RECT -482.530 -700.220 -481.930 -670.220 ;
        RECT -451.930 -700.220 -450.130 -670.220 ;
        RECT -482.530 -700.820 -450.130 -700.220 ;
        RECT -446.830 -670.220 -414.430 -669.620 ;
        RECT -446.830 -700.220 -445.030 -670.220 ;
        RECT -415.030 -700.220 -414.430 -670.220 ;
        RECT -446.830 -700.820 -414.430 -700.220 ;
        RECT -407.530 -670.220 -375.130 -669.620 ;
        RECT -407.530 -700.220 -406.930 -670.220 ;
        RECT -376.930 -700.220 -375.130 -670.220 ;
        RECT -407.530 -700.820 -375.130 -700.220 ;
        RECT -371.830 -670.220 -339.430 -669.620 ;
        RECT -371.830 -700.220 -370.030 -670.220 ;
        RECT -340.030 -700.220 -339.430 -670.220 ;
        RECT -371.830 -700.820 -339.430 -700.220 ;
        RECT -332.530 -670.220 -300.130 -669.620 ;
        RECT -332.530 -700.220 -331.930 -670.220 ;
        RECT -301.930 -700.220 -300.130 -670.220 ;
        RECT -332.530 -700.820 -300.130 -700.220 ;
        RECT -296.830 -670.220 -264.430 -669.620 ;
        RECT -296.830 -700.220 -295.030 -670.220 ;
        RECT -265.030 -700.220 -264.430 -670.220 ;
        RECT -296.830 -700.820 -264.430 -700.220 ;
        RECT -257.530 -670.220 -225.130 -669.620 ;
        RECT -257.530 -700.220 -256.930 -670.220 ;
        RECT -226.930 -700.220 -225.130 -670.220 ;
        RECT -257.530 -700.820 -225.130 -700.220 ;
        RECT -221.830 -670.220 -189.430 -669.620 ;
        RECT -221.830 -700.220 -220.030 -670.220 ;
        RECT -190.030 -700.220 -189.430 -670.220 ;
        RECT -221.830 -700.820 -189.430 -700.220 ;
        RECT -182.530 -670.220 -150.130 -669.620 ;
        RECT -182.530 -700.220 -181.930 -670.220 ;
        RECT -151.930 -700.220 -150.130 -670.220 ;
        RECT -182.530 -700.820 -150.130 -700.220 ;
        RECT -146.830 -670.220 -114.430 -669.620 ;
        RECT -146.830 -700.220 -145.030 -670.220 ;
        RECT -115.030 -700.220 -114.430 -670.220 ;
        RECT -146.830 -700.820 -114.430 -700.220 ;
        RECT -107.530 -670.220 -75.130 -669.620 ;
        RECT -107.530 -700.220 -106.930 -670.220 ;
        RECT -76.930 -700.220 -75.130 -670.220 ;
        RECT -107.530 -700.820 -75.130 -700.220 ;
        RECT -71.830 -670.220 -39.430 -669.620 ;
        RECT -71.830 -700.220 -70.030 -670.220 ;
        RECT -40.030 -700.220 -39.430 -670.220 ;
        RECT -71.830 -700.820 -39.430 -700.220 ;
        RECT -32.530 -670.220 -0.130 -669.620 ;
        RECT -32.530 -700.220 -31.930 -670.220 ;
        RECT -1.930 -700.220 -0.130 -670.220 ;
        RECT -32.530 -700.820 -0.130 -700.220 ;
        RECT 3.170 -670.220 35.570 -669.620 ;
        RECT 3.170 -700.220 4.970 -670.220 ;
        RECT 34.970 -700.220 35.570 -670.220 ;
        RECT 3.170 -700.820 35.570 -700.220 ;
        RECT 42.470 -670.220 74.870 -669.620 ;
        RECT 42.470 -700.220 43.070 -670.220 ;
        RECT 73.070 -700.220 74.870 -670.220 ;
        RECT 42.470 -700.820 74.870 -700.220 ;
        RECT 78.170 -670.220 110.570 -669.620 ;
        RECT 78.170 -700.220 79.970 -670.220 ;
        RECT 109.970 -700.220 110.570 -670.220 ;
        RECT 78.170 -700.820 110.570 -700.220 ;
        RECT 117.470 -670.220 149.870 -669.620 ;
        RECT 117.470 -700.220 118.070 -670.220 ;
        RECT 148.070 -700.220 149.870 -670.220 ;
        RECT 117.470 -700.820 149.870 -700.220 ;
        RECT 153.170 -670.220 185.570 -669.620 ;
        RECT 153.170 -700.220 154.970 -670.220 ;
        RECT 184.970 -700.220 185.570 -670.220 ;
        RECT 153.170 -700.820 185.570 -700.220 ;
        RECT 192.470 -670.220 224.870 -669.620 ;
        RECT 192.470 -700.220 193.070 -670.220 ;
        RECT 223.070 -700.220 224.870 -670.220 ;
        RECT 192.470 -700.820 224.870 -700.220 ;
        RECT 228.170 -670.220 260.570 -669.620 ;
        RECT 228.170 -700.220 229.970 -670.220 ;
        RECT 259.970 -700.220 260.570 -670.220 ;
        RECT 228.170 -700.820 260.570 -700.220 ;
        RECT 267.470 -670.220 299.870 -669.620 ;
        RECT 267.470 -700.220 268.070 -670.220 ;
        RECT 298.070 -700.220 299.870 -670.220 ;
        RECT 267.470 -700.820 299.870 -700.220 ;
        RECT 303.170 -670.220 335.570 -669.620 ;
        RECT 303.170 -700.220 304.970 -670.220 ;
        RECT 334.970 -700.220 335.570 -670.220 ;
        RECT 303.170 -700.820 335.570 -700.220 ;
        RECT 342.470 -670.220 374.870 -669.620 ;
        RECT 342.470 -700.220 343.070 -670.220 ;
        RECT 373.070 -700.220 374.870 -670.220 ;
        RECT 342.470 -700.820 374.870 -700.220 ;
        RECT 378.170 -670.220 410.570 -669.620 ;
        RECT 378.170 -700.220 379.970 -670.220 ;
        RECT 409.970 -700.220 410.570 -670.220 ;
        RECT 378.170 -700.820 410.570 -700.220 ;
        RECT 417.470 -670.220 449.870 -669.620 ;
        RECT 417.470 -700.220 418.070 -670.220 ;
        RECT 448.070 -700.220 449.870 -670.220 ;
        RECT 417.470 -700.820 449.870 -700.220 ;
        RECT 453.170 -670.220 485.570 -669.620 ;
        RECT 453.170 -700.220 454.970 -670.220 ;
        RECT 484.970 -700.220 485.570 -670.220 ;
        RECT 453.170 -700.820 485.570 -700.220 ;
        RECT 492.470 -670.220 524.870 -669.620 ;
        RECT 492.470 -700.220 493.070 -670.220 ;
        RECT 523.070 -700.220 524.870 -670.220 ;
        RECT 492.470 -700.820 524.870 -700.220 ;
        RECT 528.170 -670.220 560.570 -669.620 ;
        RECT 528.170 -700.220 529.970 -670.220 ;
        RECT 559.970 -700.220 560.570 -670.220 ;
        RECT 528.170 -700.820 560.570 -700.220 ;
        RECT -557.530 -705.220 -525.130 -704.620 ;
        RECT -557.530 -735.220 -556.930 -705.220 ;
        RECT -526.930 -735.220 -525.130 -705.220 ;
        RECT -557.530 -735.820 -525.130 -735.220 ;
        RECT -521.830 -705.220 -489.430 -704.620 ;
        RECT -521.830 -735.220 -520.030 -705.220 ;
        RECT -490.030 -735.220 -489.430 -705.220 ;
        RECT -521.830 -735.820 -489.430 -735.220 ;
        RECT -482.530 -705.220 -450.130 -704.620 ;
        RECT -482.530 -735.220 -481.930 -705.220 ;
        RECT -451.930 -735.220 -450.130 -705.220 ;
        RECT -482.530 -735.820 -450.130 -735.220 ;
        RECT -446.830 -705.220 -414.430 -704.620 ;
        RECT -446.830 -735.220 -445.030 -705.220 ;
        RECT -415.030 -735.220 -414.430 -705.220 ;
        RECT -446.830 -735.820 -414.430 -735.220 ;
        RECT -407.530 -705.220 -375.130 -704.620 ;
        RECT -407.530 -735.220 -406.930 -705.220 ;
        RECT -376.930 -735.220 -375.130 -705.220 ;
        RECT -407.530 -735.820 -375.130 -735.220 ;
        RECT -371.830 -705.220 -339.430 -704.620 ;
        RECT -371.830 -735.220 -370.030 -705.220 ;
        RECT -340.030 -735.220 -339.430 -705.220 ;
        RECT -371.830 -735.820 -339.430 -735.220 ;
        RECT -332.530 -705.220 -300.130 -704.620 ;
        RECT -332.530 -735.220 -331.930 -705.220 ;
        RECT -301.930 -735.220 -300.130 -705.220 ;
        RECT -332.530 -735.820 -300.130 -735.220 ;
        RECT -296.830 -705.220 -264.430 -704.620 ;
        RECT -296.830 -735.220 -295.030 -705.220 ;
        RECT -265.030 -735.220 -264.430 -705.220 ;
        RECT -296.830 -735.820 -264.430 -735.220 ;
        RECT -257.530 -705.220 -225.130 -704.620 ;
        RECT -257.530 -735.220 -256.930 -705.220 ;
        RECT -226.930 -735.220 -225.130 -705.220 ;
        RECT -257.530 -735.820 -225.130 -735.220 ;
        RECT -221.830 -705.220 -189.430 -704.620 ;
        RECT -221.830 -735.220 -220.030 -705.220 ;
        RECT -190.030 -735.220 -189.430 -705.220 ;
        RECT -221.830 -735.820 -189.430 -735.220 ;
        RECT -182.530 -705.220 -150.130 -704.620 ;
        RECT -182.530 -735.220 -181.930 -705.220 ;
        RECT -151.930 -735.220 -150.130 -705.220 ;
        RECT -182.530 -735.820 -150.130 -735.220 ;
        RECT -146.830 -705.220 -114.430 -704.620 ;
        RECT -146.830 -735.220 -145.030 -705.220 ;
        RECT -115.030 -735.220 -114.430 -705.220 ;
        RECT -146.830 -735.820 -114.430 -735.220 ;
        RECT -107.530 -705.220 -75.130 -704.620 ;
        RECT -107.530 -735.220 -106.930 -705.220 ;
        RECT -76.930 -735.220 -75.130 -705.220 ;
        RECT -107.530 -735.820 -75.130 -735.220 ;
        RECT -71.830 -705.220 -39.430 -704.620 ;
        RECT -71.830 -735.220 -70.030 -705.220 ;
        RECT -40.030 -735.220 -39.430 -705.220 ;
        RECT -71.830 -735.820 -39.430 -735.220 ;
        RECT -32.530 -705.220 -0.130 -704.620 ;
        RECT -32.530 -735.220 -31.930 -705.220 ;
        RECT -1.930 -735.220 -0.130 -705.220 ;
        RECT -32.530 -735.820 -0.130 -735.220 ;
        RECT 3.170 -705.220 35.570 -704.620 ;
        RECT 3.170 -735.220 4.970 -705.220 ;
        RECT 34.970 -735.220 35.570 -705.220 ;
        RECT 3.170 -735.820 35.570 -735.220 ;
        RECT 42.470 -705.220 74.870 -704.620 ;
        RECT 42.470 -735.220 43.070 -705.220 ;
        RECT 73.070 -735.220 74.870 -705.220 ;
        RECT 42.470 -735.820 74.870 -735.220 ;
        RECT 78.170 -705.220 110.570 -704.620 ;
        RECT 78.170 -735.220 79.970 -705.220 ;
        RECT 109.970 -735.220 110.570 -705.220 ;
        RECT 78.170 -735.820 110.570 -735.220 ;
        RECT 117.470 -705.220 149.870 -704.620 ;
        RECT 117.470 -735.220 118.070 -705.220 ;
        RECT 148.070 -735.220 149.870 -705.220 ;
        RECT 117.470 -735.820 149.870 -735.220 ;
        RECT 153.170 -705.220 185.570 -704.620 ;
        RECT 153.170 -735.220 154.970 -705.220 ;
        RECT 184.970 -735.220 185.570 -705.220 ;
        RECT 153.170 -735.820 185.570 -735.220 ;
        RECT 192.470 -705.220 224.870 -704.620 ;
        RECT 192.470 -735.220 193.070 -705.220 ;
        RECT 223.070 -735.220 224.870 -705.220 ;
        RECT 192.470 -735.820 224.870 -735.220 ;
        RECT 228.170 -705.220 260.570 -704.620 ;
        RECT 228.170 -735.220 229.970 -705.220 ;
        RECT 259.970 -735.220 260.570 -705.220 ;
        RECT 228.170 -735.820 260.570 -735.220 ;
        RECT 267.470 -705.220 299.870 -704.620 ;
        RECT 267.470 -735.220 268.070 -705.220 ;
        RECT 298.070 -735.220 299.870 -705.220 ;
        RECT 267.470 -735.820 299.870 -735.220 ;
        RECT 303.170 -705.220 335.570 -704.620 ;
        RECT 303.170 -735.220 304.970 -705.220 ;
        RECT 334.970 -735.220 335.570 -705.220 ;
        RECT 303.170 -735.820 335.570 -735.220 ;
        RECT 342.470 -705.220 374.870 -704.620 ;
        RECT 342.470 -735.220 343.070 -705.220 ;
        RECT 373.070 -735.220 374.870 -705.220 ;
        RECT 342.470 -735.820 374.870 -735.220 ;
        RECT 378.170 -705.220 410.570 -704.620 ;
        RECT 378.170 -735.220 379.970 -705.220 ;
        RECT 409.970 -735.220 410.570 -705.220 ;
        RECT 378.170 -735.820 410.570 -735.220 ;
        RECT 417.470 -705.220 449.870 -704.620 ;
        RECT 417.470 -735.220 418.070 -705.220 ;
        RECT 448.070 -735.220 449.870 -705.220 ;
        RECT 417.470 -735.820 449.870 -735.220 ;
        RECT 453.170 -705.220 485.570 -704.620 ;
        RECT 453.170 -735.220 454.970 -705.220 ;
        RECT 484.970 -735.220 485.570 -705.220 ;
        RECT 453.170 -735.820 485.570 -735.220 ;
        RECT 492.470 -705.220 524.870 -704.620 ;
        RECT 492.470 -735.220 493.070 -705.220 ;
        RECT 523.070 -735.220 524.870 -705.220 ;
        RECT 492.470 -735.820 524.870 -735.220 ;
        RECT 528.170 -705.220 560.570 -704.620 ;
        RECT 528.170 -735.220 529.970 -705.220 ;
        RECT 559.970 -735.220 560.570 -705.220 ;
        RECT 528.170 -735.820 560.570 -735.220 ;
        RECT -557.530 -740.220 -525.130 -739.620 ;
        RECT -557.530 -770.220 -556.930 -740.220 ;
        RECT -526.930 -770.220 -525.130 -740.220 ;
        RECT -557.530 -770.820 -525.130 -770.220 ;
        RECT -521.830 -740.220 -489.430 -739.620 ;
        RECT -521.830 -770.220 -520.030 -740.220 ;
        RECT -490.030 -770.220 -489.430 -740.220 ;
        RECT -521.830 -770.820 -489.430 -770.220 ;
        RECT -482.530 -740.220 -450.130 -739.620 ;
        RECT -482.530 -770.220 -481.930 -740.220 ;
        RECT -451.930 -770.220 -450.130 -740.220 ;
        RECT -482.530 -770.820 -450.130 -770.220 ;
        RECT -446.830 -740.220 -414.430 -739.620 ;
        RECT -446.830 -770.220 -445.030 -740.220 ;
        RECT -415.030 -770.220 -414.430 -740.220 ;
        RECT -446.830 -770.820 -414.430 -770.220 ;
        RECT -407.530 -740.220 -375.130 -739.620 ;
        RECT -407.530 -770.220 -406.930 -740.220 ;
        RECT -376.930 -770.220 -375.130 -740.220 ;
        RECT -407.530 -770.820 -375.130 -770.220 ;
        RECT -371.830 -740.220 -339.430 -739.620 ;
        RECT -371.830 -770.220 -370.030 -740.220 ;
        RECT -340.030 -770.220 -339.430 -740.220 ;
        RECT -371.830 -770.820 -339.430 -770.220 ;
        RECT -332.530 -740.220 -300.130 -739.620 ;
        RECT -332.530 -770.220 -331.930 -740.220 ;
        RECT -301.930 -770.220 -300.130 -740.220 ;
        RECT -332.530 -770.820 -300.130 -770.220 ;
        RECT -296.830 -740.220 -264.430 -739.620 ;
        RECT -296.830 -770.220 -295.030 -740.220 ;
        RECT -265.030 -770.220 -264.430 -740.220 ;
        RECT -296.830 -770.820 -264.430 -770.220 ;
        RECT -257.530 -740.220 -225.130 -739.620 ;
        RECT -257.530 -770.220 -256.930 -740.220 ;
        RECT -226.930 -770.220 -225.130 -740.220 ;
        RECT -257.530 -770.820 -225.130 -770.220 ;
        RECT -221.830 -740.220 -189.430 -739.620 ;
        RECT -221.830 -770.220 -220.030 -740.220 ;
        RECT -190.030 -770.220 -189.430 -740.220 ;
        RECT -221.830 -770.820 -189.430 -770.220 ;
        RECT -182.530 -740.220 -150.130 -739.620 ;
        RECT -182.530 -770.220 -181.930 -740.220 ;
        RECT -151.930 -770.220 -150.130 -740.220 ;
        RECT -182.530 -770.820 -150.130 -770.220 ;
        RECT -146.830 -740.220 -114.430 -739.620 ;
        RECT -146.830 -770.220 -145.030 -740.220 ;
        RECT -115.030 -770.220 -114.430 -740.220 ;
        RECT -146.830 -770.820 -114.430 -770.220 ;
        RECT -107.530 -740.220 -75.130 -739.620 ;
        RECT -107.530 -770.220 -106.930 -740.220 ;
        RECT -76.930 -770.220 -75.130 -740.220 ;
        RECT -107.530 -770.820 -75.130 -770.220 ;
        RECT -71.830 -740.220 -39.430 -739.620 ;
        RECT -71.830 -770.220 -70.030 -740.220 ;
        RECT -40.030 -770.220 -39.430 -740.220 ;
        RECT -71.830 -770.820 -39.430 -770.220 ;
        RECT -32.530 -740.220 -0.130 -739.620 ;
        RECT -32.530 -770.220 -31.930 -740.220 ;
        RECT -1.930 -770.220 -0.130 -740.220 ;
        RECT -32.530 -770.820 -0.130 -770.220 ;
        RECT 3.170 -740.220 35.570 -739.620 ;
        RECT 3.170 -770.220 4.970 -740.220 ;
        RECT 34.970 -770.220 35.570 -740.220 ;
        RECT 3.170 -770.820 35.570 -770.220 ;
        RECT 42.470 -740.220 74.870 -739.620 ;
        RECT 42.470 -770.220 43.070 -740.220 ;
        RECT 73.070 -770.220 74.870 -740.220 ;
        RECT 42.470 -770.820 74.870 -770.220 ;
        RECT 78.170 -740.220 110.570 -739.620 ;
        RECT 78.170 -770.220 79.970 -740.220 ;
        RECT 109.970 -770.220 110.570 -740.220 ;
        RECT 78.170 -770.820 110.570 -770.220 ;
        RECT 117.470 -740.220 149.870 -739.620 ;
        RECT 117.470 -770.220 118.070 -740.220 ;
        RECT 148.070 -770.220 149.870 -740.220 ;
        RECT 117.470 -770.820 149.870 -770.220 ;
        RECT 153.170 -740.220 185.570 -739.620 ;
        RECT 153.170 -770.220 154.970 -740.220 ;
        RECT 184.970 -770.220 185.570 -740.220 ;
        RECT 153.170 -770.820 185.570 -770.220 ;
        RECT 192.470 -740.220 224.870 -739.620 ;
        RECT 192.470 -770.220 193.070 -740.220 ;
        RECT 223.070 -770.220 224.870 -740.220 ;
        RECT 192.470 -770.820 224.870 -770.220 ;
        RECT 228.170 -740.220 260.570 -739.620 ;
        RECT 228.170 -770.220 229.970 -740.220 ;
        RECT 259.970 -770.220 260.570 -740.220 ;
        RECT 228.170 -770.820 260.570 -770.220 ;
        RECT 267.470 -740.220 299.870 -739.620 ;
        RECT 267.470 -770.220 268.070 -740.220 ;
        RECT 298.070 -770.220 299.870 -740.220 ;
        RECT 267.470 -770.820 299.870 -770.220 ;
        RECT 303.170 -740.220 335.570 -739.620 ;
        RECT 303.170 -770.220 304.970 -740.220 ;
        RECT 334.970 -770.220 335.570 -740.220 ;
        RECT 303.170 -770.820 335.570 -770.220 ;
        RECT 342.470 -740.220 374.870 -739.620 ;
        RECT 342.470 -770.220 343.070 -740.220 ;
        RECT 373.070 -770.220 374.870 -740.220 ;
        RECT 342.470 -770.820 374.870 -770.220 ;
        RECT 378.170 -740.220 410.570 -739.620 ;
        RECT 378.170 -770.220 379.970 -740.220 ;
        RECT 409.970 -770.220 410.570 -740.220 ;
        RECT 378.170 -770.820 410.570 -770.220 ;
        RECT 417.470 -740.220 449.870 -739.620 ;
        RECT 417.470 -770.220 418.070 -740.220 ;
        RECT 448.070 -770.220 449.870 -740.220 ;
        RECT 417.470 -770.820 449.870 -770.220 ;
        RECT 453.170 -740.220 485.570 -739.620 ;
        RECT 453.170 -770.220 454.970 -740.220 ;
        RECT 484.970 -770.220 485.570 -740.220 ;
        RECT 453.170 -770.820 485.570 -770.220 ;
        RECT 492.470 -740.220 524.870 -739.620 ;
        RECT 492.470 -770.220 493.070 -740.220 ;
        RECT 523.070 -770.220 524.870 -740.220 ;
        RECT 492.470 -770.820 524.870 -770.220 ;
        RECT 528.170 -740.220 560.570 -739.620 ;
        RECT 528.170 -770.220 529.970 -740.220 ;
        RECT 559.970 -770.220 560.570 -740.220 ;
        RECT 528.170 -770.820 560.570 -770.220 ;
        RECT -557.530 -775.220 -525.130 -774.620 ;
        RECT -557.530 -805.220 -556.930 -775.220 ;
        RECT -526.930 -805.220 -525.130 -775.220 ;
        RECT -557.530 -805.820 -525.130 -805.220 ;
        RECT -521.830 -775.220 -489.430 -774.620 ;
        RECT -521.830 -805.220 -520.030 -775.220 ;
        RECT -490.030 -805.220 -489.430 -775.220 ;
        RECT -521.830 -805.820 -489.430 -805.220 ;
        RECT -482.530 -775.220 -450.130 -774.620 ;
        RECT -482.530 -805.220 -481.930 -775.220 ;
        RECT -451.930 -805.220 -450.130 -775.220 ;
        RECT -482.530 -805.820 -450.130 -805.220 ;
        RECT -446.830 -775.220 -414.430 -774.620 ;
        RECT -446.830 -805.220 -445.030 -775.220 ;
        RECT -415.030 -805.220 -414.430 -775.220 ;
        RECT -446.830 -805.820 -414.430 -805.220 ;
        RECT -407.530 -775.220 -375.130 -774.620 ;
        RECT -407.530 -805.220 -406.930 -775.220 ;
        RECT -376.930 -805.220 -375.130 -775.220 ;
        RECT -407.530 -805.820 -375.130 -805.220 ;
        RECT -371.830 -775.220 -339.430 -774.620 ;
        RECT -371.830 -805.220 -370.030 -775.220 ;
        RECT -340.030 -805.220 -339.430 -775.220 ;
        RECT -371.830 -805.820 -339.430 -805.220 ;
        RECT -332.530 -775.220 -300.130 -774.620 ;
        RECT -332.530 -805.220 -331.930 -775.220 ;
        RECT -301.930 -805.220 -300.130 -775.220 ;
        RECT -332.530 -805.820 -300.130 -805.220 ;
        RECT -296.830 -775.220 -264.430 -774.620 ;
        RECT -296.830 -805.220 -295.030 -775.220 ;
        RECT -265.030 -805.220 -264.430 -775.220 ;
        RECT -296.830 -805.820 -264.430 -805.220 ;
        RECT -257.530 -775.220 -225.130 -774.620 ;
        RECT -257.530 -805.220 -256.930 -775.220 ;
        RECT -226.930 -805.220 -225.130 -775.220 ;
        RECT -257.530 -805.820 -225.130 -805.220 ;
        RECT -221.830 -775.220 -189.430 -774.620 ;
        RECT -221.830 -805.220 -220.030 -775.220 ;
        RECT -190.030 -805.220 -189.430 -775.220 ;
        RECT -221.830 -805.820 -189.430 -805.220 ;
        RECT -182.530 -775.220 -150.130 -774.620 ;
        RECT -182.530 -805.220 -181.930 -775.220 ;
        RECT -151.930 -805.220 -150.130 -775.220 ;
        RECT -182.530 -805.820 -150.130 -805.220 ;
        RECT -146.830 -775.220 -114.430 -774.620 ;
        RECT -146.830 -805.220 -145.030 -775.220 ;
        RECT -115.030 -805.220 -114.430 -775.220 ;
        RECT -146.830 -805.820 -114.430 -805.220 ;
        RECT -107.530 -775.220 -75.130 -774.620 ;
        RECT -107.530 -805.220 -106.930 -775.220 ;
        RECT -76.930 -805.220 -75.130 -775.220 ;
        RECT -107.530 -805.820 -75.130 -805.220 ;
        RECT -71.830 -775.220 -39.430 -774.620 ;
        RECT -71.830 -805.220 -70.030 -775.220 ;
        RECT -40.030 -805.220 -39.430 -775.220 ;
        RECT -71.830 -805.820 -39.430 -805.220 ;
        RECT -32.530 -775.220 -0.130 -774.620 ;
        RECT -32.530 -805.220 -31.930 -775.220 ;
        RECT -1.930 -805.220 -0.130 -775.220 ;
        RECT -32.530 -805.820 -0.130 -805.220 ;
        RECT 3.170 -775.220 35.570 -774.620 ;
        RECT 3.170 -805.220 4.970 -775.220 ;
        RECT 34.970 -805.220 35.570 -775.220 ;
        RECT 3.170 -805.820 35.570 -805.220 ;
        RECT 42.470 -775.220 74.870 -774.620 ;
        RECT 42.470 -805.220 43.070 -775.220 ;
        RECT 73.070 -805.220 74.870 -775.220 ;
        RECT 42.470 -805.820 74.870 -805.220 ;
        RECT 78.170 -775.220 110.570 -774.620 ;
        RECT 78.170 -805.220 79.970 -775.220 ;
        RECT 109.970 -805.220 110.570 -775.220 ;
        RECT 78.170 -805.820 110.570 -805.220 ;
        RECT 117.470 -775.220 149.870 -774.620 ;
        RECT 117.470 -805.220 118.070 -775.220 ;
        RECT 148.070 -805.220 149.870 -775.220 ;
        RECT 117.470 -805.820 149.870 -805.220 ;
        RECT 153.170 -775.220 185.570 -774.620 ;
        RECT 153.170 -805.220 154.970 -775.220 ;
        RECT 184.970 -805.220 185.570 -775.220 ;
        RECT 153.170 -805.820 185.570 -805.220 ;
        RECT 192.470 -775.220 224.870 -774.620 ;
        RECT 192.470 -805.220 193.070 -775.220 ;
        RECT 223.070 -805.220 224.870 -775.220 ;
        RECT 192.470 -805.820 224.870 -805.220 ;
        RECT 228.170 -775.220 260.570 -774.620 ;
        RECT 228.170 -805.220 229.970 -775.220 ;
        RECT 259.970 -805.220 260.570 -775.220 ;
        RECT 228.170 -805.820 260.570 -805.220 ;
        RECT 267.470 -775.220 299.870 -774.620 ;
        RECT 267.470 -805.220 268.070 -775.220 ;
        RECT 298.070 -805.220 299.870 -775.220 ;
        RECT 267.470 -805.820 299.870 -805.220 ;
        RECT 303.170 -775.220 335.570 -774.620 ;
        RECT 303.170 -805.220 304.970 -775.220 ;
        RECT 334.970 -805.220 335.570 -775.220 ;
        RECT 303.170 -805.820 335.570 -805.220 ;
        RECT 342.470 -775.220 374.870 -774.620 ;
        RECT 342.470 -805.220 343.070 -775.220 ;
        RECT 373.070 -805.220 374.870 -775.220 ;
        RECT 342.470 -805.820 374.870 -805.220 ;
        RECT 378.170 -775.220 410.570 -774.620 ;
        RECT 378.170 -805.220 379.970 -775.220 ;
        RECT 409.970 -805.220 410.570 -775.220 ;
        RECT 378.170 -805.820 410.570 -805.220 ;
        RECT 417.470 -775.220 449.870 -774.620 ;
        RECT 417.470 -805.220 418.070 -775.220 ;
        RECT 448.070 -805.220 449.870 -775.220 ;
        RECT 417.470 -805.820 449.870 -805.220 ;
        RECT 453.170 -775.220 485.570 -774.620 ;
        RECT 453.170 -805.220 454.970 -775.220 ;
        RECT 484.970 -805.220 485.570 -775.220 ;
        RECT 453.170 -805.820 485.570 -805.220 ;
        RECT 492.470 -775.220 524.870 -774.620 ;
        RECT 492.470 -805.220 493.070 -775.220 ;
        RECT 523.070 -805.220 524.870 -775.220 ;
        RECT 492.470 -805.820 524.870 -805.220 ;
        RECT 528.170 -775.220 560.570 -774.620 ;
        RECT 528.170 -805.220 529.970 -775.220 ;
        RECT 559.970 -805.220 560.570 -775.220 ;
        RECT 528.170 -805.820 560.570 -805.220 ;
        RECT -557.530 -810.220 -525.130 -809.620 ;
        RECT -557.530 -840.220 -556.930 -810.220 ;
        RECT -526.930 -840.220 -525.130 -810.220 ;
        RECT -557.530 -840.820 -525.130 -840.220 ;
        RECT -521.830 -810.220 -489.430 -809.620 ;
        RECT -521.830 -840.220 -520.030 -810.220 ;
        RECT -490.030 -840.220 -489.430 -810.220 ;
        RECT -521.830 -840.820 -489.430 -840.220 ;
        RECT -482.530 -810.220 -450.130 -809.620 ;
        RECT -482.530 -840.220 -481.930 -810.220 ;
        RECT -451.930 -840.220 -450.130 -810.220 ;
        RECT -482.530 -840.820 -450.130 -840.220 ;
        RECT -446.830 -810.220 -414.430 -809.620 ;
        RECT -446.830 -840.220 -445.030 -810.220 ;
        RECT -415.030 -840.220 -414.430 -810.220 ;
        RECT -446.830 -840.820 -414.430 -840.220 ;
        RECT -407.530 -810.220 -375.130 -809.620 ;
        RECT -407.530 -840.220 -406.930 -810.220 ;
        RECT -376.930 -840.220 -375.130 -810.220 ;
        RECT -407.530 -840.820 -375.130 -840.220 ;
        RECT -371.830 -810.220 -339.430 -809.620 ;
        RECT -371.830 -840.220 -370.030 -810.220 ;
        RECT -340.030 -840.220 -339.430 -810.220 ;
        RECT -371.830 -840.820 -339.430 -840.220 ;
        RECT -332.530 -810.220 -300.130 -809.620 ;
        RECT -332.530 -840.220 -331.930 -810.220 ;
        RECT -301.930 -840.220 -300.130 -810.220 ;
        RECT -332.530 -840.820 -300.130 -840.220 ;
        RECT -296.830 -810.220 -264.430 -809.620 ;
        RECT -296.830 -840.220 -295.030 -810.220 ;
        RECT -265.030 -840.220 -264.430 -810.220 ;
        RECT -296.830 -840.820 -264.430 -840.220 ;
        RECT -257.530 -810.220 -225.130 -809.620 ;
        RECT -257.530 -840.220 -256.930 -810.220 ;
        RECT -226.930 -840.220 -225.130 -810.220 ;
        RECT -257.530 -840.820 -225.130 -840.220 ;
        RECT -221.830 -810.220 -189.430 -809.620 ;
        RECT -221.830 -840.220 -220.030 -810.220 ;
        RECT -190.030 -840.220 -189.430 -810.220 ;
        RECT -221.830 -840.820 -189.430 -840.220 ;
        RECT -182.530 -810.220 -150.130 -809.620 ;
        RECT -182.530 -840.220 -181.930 -810.220 ;
        RECT -151.930 -840.220 -150.130 -810.220 ;
        RECT -182.530 -840.820 -150.130 -840.220 ;
        RECT -146.830 -810.220 -114.430 -809.620 ;
        RECT -146.830 -840.220 -145.030 -810.220 ;
        RECT -115.030 -840.220 -114.430 -810.220 ;
        RECT -146.830 -840.820 -114.430 -840.220 ;
        RECT -107.530 -810.220 -75.130 -809.620 ;
        RECT -107.530 -840.220 -106.930 -810.220 ;
        RECT -76.930 -840.220 -75.130 -810.220 ;
        RECT -107.530 -840.820 -75.130 -840.220 ;
        RECT -71.830 -810.220 -39.430 -809.620 ;
        RECT -71.830 -840.220 -70.030 -810.220 ;
        RECT -40.030 -840.220 -39.430 -810.220 ;
        RECT -71.830 -840.820 -39.430 -840.220 ;
        RECT -32.530 -810.220 -0.130 -809.620 ;
        RECT -32.530 -840.220 -31.930 -810.220 ;
        RECT -1.930 -840.220 -0.130 -810.220 ;
        RECT -32.530 -840.820 -0.130 -840.220 ;
        RECT 3.170 -810.220 35.570 -809.620 ;
        RECT 3.170 -840.220 4.970 -810.220 ;
        RECT 34.970 -840.220 35.570 -810.220 ;
        RECT 3.170 -840.820 35.570 -840.220 ;
        RECT 42.470 -810.220 74.870 -809.620 ;
        RECT 42.470 -840.220 43.070 -810.220 ;
        RECT 73.070 -840.220 74.870 -810.220 ;
        RECT 42.470 -840.820 74.870 -840.220 ;
        RECT 78.170 -810.220 110.570 -809.620 ;
        RECT 78.170 -840.220 79.970 -810.220 ;
        RECT 109.970 -840.220 110.570 -810.220 ;
        RECT 78.170 -840.820 110.570 -840.220 ;
        RECT 117.470 -810.220 149.870 -809.620 ;
        RECT 117.470 -840.220 118.070 -810.220 ;
        RECT 148.070 -840.220 149.870 -810.220 ;
        RECT 117.470 -840.820 149.870 -840.220 ;
        RECT 153.170 -810.220 185.570 -809.620 ;
        RECT 153.170 -840.220 154.970 -810.220 ;
        RECT 184.970 -840.220 185.570 -810.220 ;
        RECT 153.170 -840.820 185.570 -840.220 ;
        RECT 192.470 -810.220 224.870 -809.620 ;
        RECT 192.470 -840.220 193.070 -810.220 ;
        RECT 223.070 -840.220 224.870 -810.220 ;
        RECT 192.470 -840.820 224.870 -840.220 ;
        RECT 228.170 -810.220 260.570 -809.620 ;
        RECT 228.170 -840.220 229.970 -810.220 ;
        RECT 259.970 -840.220 260.570 -810.220 ;
        RECT 228.170 -840.820 260.570 -840.220 ;
        RECT 267.470 -810.220 299.870 -809.620 ;
        RECT 267.470 -840.220 268.070 -810.220 ;
        RECT 298.070 -840.220 299.870 -810.220 ;
        RECT 267.470 -840.820 299.870 -840.220 ;
        RECT 303.170 -810.220 335.570 -809.620 ;
        RECT 303.170 -840.220 304.970 -810.220 ;
        RECT 334.970 -840.220 335.570 -810.220 ;
        RECT 303.170 -840.820 335.570 -840.220 ;
        RECT 342.470 -810.220 374.870 -809.620 ;
        RECT 342.470 -840.220 343.070 -810.220 ;
        RECT 373.070 -840.220 374.870 -810.220 ;
        RECT 342.470 -840.820 374.870 -840.220 ;
        RECT 378.170 -810.220 410.570 -809.620 ;
        RECT 378.170 -840.220 379.970 -810.220 ;
        RECT 409.970 -840.220 410.570 -810.220 ;
        RECT 378.170 -840.820 410.570 -840.220 ;
        RECT 417.470 -810.220 449.870 -809.620 ;
        RECT 417.470 -840.220 418.070 -810.220 ;
        RECT 448.070 -840.220 449.870 -810.220 ;
        RECT 417.470 -840.820 449.870 -840.220 ;
        RECT 453.170 -810.220 485.570 -809.620 ;
        RECT 453.170 -840.220 454.970 -810.220 ;
        RECT 484.970 -840.220 485.570 -810.220 ;
        RECT 453.170 -840.820 485.570 -840.220 ;
        RECT 492.470 -810.220 524.870 -809.620 ;
        RECT 492.470 -840.220 493.070 -810.220 ;
        RECT 523.070 -840.220 524.870 -810.220 ;
        RECT 492.470 -840.820 524.870 -840.220 ;
        RECT 528.170 -810.220 560.570 -809.620 ;
        RECT 528.170 -840.220 529.970 -810.220 ;
        RECT 559.970 -840.220 560.570 -810.220 ;
        RECT 528.170 -840.820 560.570 -840.220 ;
        RECT -557.530 -845.220 -525.130 -844.620 ;
        RECT -557.530 -875.220 -556.930 -845.220 ;
        RECT -526.930 -875.220 -525.130 -845.220 ;
        RECT -557.530 -875.820 -525.130 -875.220 ;
        RECT -521.830 -845.220 -489.430 -844.620 ;
        RECT -521.830 -875.220 -520.030 -845.220 ;
        RECT -490.030 -875.220 -489.430 -845.220 ;
        RECT -521.830 -875.820 -489.430 -875.220 ;
        RECT -482.530 -845.220 -450.130 -844.620 ;
        RECT -482.530 -875.220 -481.930 -845.220 ;
        RECT -451.930 -875.220 -450.130 -845.220 ;
        RECT -482.530 -875.820 -450.130 -875.220 ;
        RECT -446.830 -845.220 -414.430 -844.620 ;
        RECT -446.830 -875.220 -445.030 -845.220 ;
        RECT -415.030 -875.220 -414.430 -845.220 ;
        RECT -446.830 -875.820 -414.430 -875.220 ;
        RECT -407.530 -845.220 -375.130 -844.620 ;
        RECT -407.530 -875.220 -406.930 -845.220 ;
        RECT -376.930 -875.220 -375.130 -845.220 ;
        RECT -407.530 -875.820 -375.130 -875.220 ;
        RECT -371.830 -845.220 -339.430 -844.620 ;
        RECT -371.830 -875.220 -370.030 -845.220 ;
        RECT -340.030 -875.220 -339.430 -845.220 ;
        RECT -371.830 -875.820 -339.430 -875.220 ;
        RECT -332.530 -845.220 -300.130 -844.620 ;
        RECT -332.530 -875.220 -331.930 -845.220 ;
        RECT -301.930 -875.220 -300.130 -845.220 ;
        RECT -332.530 -875.820 -300.130 -875.220 ;
        RECT -296.830 -845.220 -264.430 -844.620 ;
        RECT -296.830 -875.220 -295.030 -845.220 ;
        RECT -265.030 -875.220 -264.430 -845.220 ;
        RECT -296.830 -875.820 -264.430 -875.220 ;
        RECT -257.530 -845.220 -225.130 -844.620 ;
        RECT -257.530 -875.220 -256.930 -845.220 ;
        RECT -226.930 -875.220 -225.130 -845.220 ;
        RECT -257.530 -875.820 -225.130 -875.220 ;
        RECT -221.830 -845.220 -189.430 -844.620 ;
        RECT -221.830 -875.220 -220.030 -845.220 ;
        RECT -190.030 -875.220 -189.430 -845.220 ;
        RECT -221.830 -875.820 -189.430 -875.220 ;
        RECT -182.530 -845.220 -150.130 -844.620 ;
        RECT -182.530 -875.220 -181.930 -845.220 ;
        RECT -151.930 -875.220 -150.130 -845.220 ;
        RECT -182.530 -875.820 -150.130 -875.220 ;
        RECT -146.830 -845.220 -114.430 -844.620 ;
        RECT -146.830 -875.220 -145.030 -845.220 ;
        RECT -115.030 -875.220 -114.430 -845.220 ;
        RECT -146.830 -875.820 -114.430 -875.220 ;
        RECT -107.530 -845.220 -75.130 -844.620 ;
        RECT -107.530 -875.220 -106.930 -845.220 ;
        RECT -76.930 -875.220 -75.130 -845.220 ;
        RECT -107.530 -875.820 -75.130 -875.220 ;
        RECT -71.830 -845.220 -39.430 -844.620 ;
        RECT -71.830 -875.220 -70.030 -845.220 ;
        RECT -40.030 -875.220 -39.430 -845.220 ;
        RECT -71.830 -875.820 -39.430 -875.220 ;
        RECT -32.530 -845.220 -0.130 -844.620 ;
        RECT -32.530 -875.220 -31.930 -845.220 ;
        RECT -1.930 -875.220 -0.130 -845.220 ;
        RECT -32.530 -875.820 -0.130 -875.220 ;
        RECT 3.170 -845.220 35.570 -844.620 ;
        RECT 3.170 -875.220 4.970 -845.220 ;
        RECT 34.970 -875.220 35.570 -845.220 ;
        RECT 3.170 -875.820 35.570 -875.220 ;
        RECT 42.470 -845.220 74.870 -844.620 ;
        RECT 42.470 -875.220 43.070 -845.220 ;
        RECT 73.070 -875.220 74.870 -845.220 ;
        RECT 42.470 -875.820 74.870 -875.220 ;
        RECT 78.170 -845.220 110.570 -844.620 ;
        RECT 78.170 -875.220 79.970 -845.220 ;
        RECT 109.970 -875.220 110.570 -845.220 ;
        RECT 78.170 -875.820 110.570 -875.220 ;
        RECT 117.470 -845.220 149.870 -844.620 ;
        RECT 117.470 -875.220 118.070 -845.220 ;
        RECT 148.070 -875.220 149.870 -845.220 ;
        RECT 117.470 -875.820 149.870 -875.220 ;
        RECT 153.170 -845.220 185.570 -844.620 ;
        RECT 153.170 -875.220 154.970 -845.220 ;
        RECT 184.970 -875.220 185.570 -845.220 ;
        RECT 153.170 -875.820 185.570 -875.220 ;
        RECT 192.470 -845.220 224.870 -844.620 ;
        RECT 192.470 -875.220 193.070 -845.220 ;
        RECT 223.070 -875.220 224.870 -845.220 ;
        RECT 192.470 -875.820 224.870 -875.220 ;
        RECT 228.170 -845.220 260.570 -844.620 ;
        RECT 228.170 -875.220 229.970 -845.220 ;
        RECT 259.970 -875.220 260.570 -845.220 ;
        RECT 228.170 -875.820 260.570 -875.220 ;
        RECT 267.470 -845.220 299.870 -844.620 ;
        RECT 267.470 -875.220 268.070 -845.220 ;
        RECT 298.070 -875.220 299.870 -845.220 ;
        RECT 267.470 -875.820 299.870 -875.220 ;
        RECT 303.170 -845.220 335.570 -844.620 ;
        RECT 303.170 -875.220 304.970 -845.220 ;
        RECT 334.970 -875.220 335.570 -845.220 ;
        RECT 303.170 -875.820 335.570 -875.220 ;
        RECT 342.470 -845.220 374.870 -844.620 ;
        RECT 342.470 -875.220 343.070 -845.220 ;
        RECT 373.070 -875.220 374.870 -845.220 ;
        RECT 342.470 -875.820 374.870 -875.220 ;
        RECT 378.170 -845.220 410.570 -844.620 ;
        RECT 378.170 -875.220 379.970 -845.220 ;
        RECT 409.970 -875.220 410.570 -845.220 ;
        RECT 378.170 -875.820 410.570 -875.220 ;
        RECT 417.470 -845.220 449.870 -844.620 ;
        RECT 417.470 -875.220 418.070 -845.220 ;
        RECT 448.070 -875.220 449.870 -845.220 ;
        RECT 417.470 -875.820 449.870 -875.220 ;
        RECT 453.170 -845.220 485.570 -844.620 ;
        RECT 453.170 -875.220 454.970 -845.220 ;
        RECT 484.970 -875.220 485.570 -845.220 ;
        RECT 453.170 -875.820 485.570 -875.220 ;
        RECT 492.470 -845.220 524.870 -844.620 ;
        RECT 492.470 -875.220 493.070 -845.220 ;
        RECT 523.070 -875.220 524.870 -845.220 ;
        RECT 492.470 -875.820 524.870 -875.220 ;
        RECT 528.170 -845.220 560.570 -844.620 ;
        RECT 528.170 -875.220 529.970 -845.220 ;
        RECT 559.970 -875.220 560.570 -845.220 ;
        RECT 528.170 -875.820 560.570 -875.220 ;
        RECT -557.530 -880.220 -525.130 -879.620 ;
        RECT -557.530 -910.220 -556.930 -880.220 ;
        RECT -526.930 -910.220 -525.130 -880.220 ;
        RECT -557.530 -910.820 -525.130 -910.220 ;
        RECT -521.830 -880.220 -489.430 -879.620 ;
        RECT -521.830 -910.220 -520.030 -880.220 ;
        RECT -490.030 -910.220 -489.430 -880.220 ;
        RECT -521.830 -910.820 -489.430 -910.220 ;
        RECT -482.530 -880.220 -450.130 -879.620 ;
        RECT -482.530 -910.220 -481.930 -880.220 ;
        RECT -451.930 -910.220 -450.130 -880.220 ;
        RECT -482.530 -910.820 -450.130 -910.220 ;
        RECT -446.830 -880.220 -414.430 -879.620 ;
        RECT -446.830 -910.220 -445.030 -880.220 ;
        RECT -415.030 -910.220 -414.430 -880.220 ;
        RECT -446.830 -910.820 -414.430 -910.220 ;
        RECT -407.530 -880.220 -375.130 -879.620 ;
        RECT -407.530 -910.220 -406.930 -880.220 ;
        RECT -376.930 -910.220 -375.130 -880.220 ;
        RECT -407.530 -910.820 -375.130 -910.220 ;
        RECT -371.830 -880.220 -339.430 -879.620 ;
        RECT -371.830 -910.220 -370.030 -880.220 ;
        RECT -340.030 -910.220 -339.430 -880.220 ;
        RECT -371.830 -910.820 -339.430 -910.220 ;
        RECT -332.530 -880.220 -300.130 -879.620 ;
        RECT -332.530 -910.220 -331.930 -880.220 ;
        RECT -301.930 -910.220 -300.130 -880.220 ;
        RECT -332.530 -910.820 -300.130 -910.220 ;
        RECT -296.830 -880.220 -264.430 -879.620 ;
        RECT -296.830 -910.220 -295.030 -880.220 ;
        RECT -265.030 -910.220 -264.430 -880.220 ;
        RECT -296.830 -910.820 -264.430 -910.220 ;
        RECT -257.530 -880.220 -225.130 -879.620 ;
        RECT -257.530 -910.220 -256.930 -880.220 ;
        RECT -226.930 -910.220 -225.130 -880.220 ;
        RECT -257.530 -910.820 -225.130 -910.220 ;
        RECT -221.830 -880.220 -189.430 -879.620 ;
        RECT -221.830 -910.220 -220.030 -880.220 ;
        RECT -190.030 -910.220 -189.430 -880.220 ;
        RECT -221.830 -910.820 -189.430 -910.220 ;
        RECT -182.530 -880.220 -150.130 -879.620 ;
        RECT -182.530 -910.220 -181.930 -880.220 ;
        RECT -151.930 -910.220 -150.130 -880.220 ;
        RECT -182.530 -910.820 -150.130 -910.220 ;
        RECT -146.830 -880.220 -114.430 -879.620 ;
        RECT -146.830 -910.220 -145.030 -880.220 ;
        RECT -115.030 -910.220 -114.430 -880.220 ;
        RECT -146.830 -910.820 -114.430 -910.220 ;
        RECT -107.530 -880.220 -75.130 -879.620 ;
        RECT -107.530 -910.220 -106.930 -880.220 ;
        RECT -76.930 -910.220 -75.130 -880.220 ;
        RECT -107.530 -910.820 -75.130 -910.220 ;
        RECT -71.830 -880.220 -39.430 -879.620 ;
        RECT -71.830 -910.220 -70.030 -880.220 ;
        RECT -40.030 -910.220 -39.430 -880.220 ;
        RECT -71.830 -910.820 -39.430 -910.220 ;
        RECT -32.530 -880.220 -0.130 -879.620 ;
        RECT -32.530 -910.220 -31.930 -880.220 ;
        RECT -1.930 -910.220 -0.130 -880.220 ;
        RECT -32.530 -910.820 -0.130 -910.220 ;
        RECT 3.170 -880.220 35.570 -879.620 ;
        RECT 3.170 -910.220 4.970 -880.220 ;
        RECT 34.970 -910.220 35.570 -880.220 ;
        RECT 3.170 -910.820 35.570 -910.220 ;
        RECT 42.470 -880.220 74.870 -879.620 ;
        RECT 42.470 -910.220 43.070 -880.220 ;
        RECT 73.070 -910.220 74.870 -880.220 ;
        RECT 42.470 -910.820 74.870 -910.220 ;
        RECT 78.170 -880.220 110.570 -879.620 ;
        RECT 78.170 -910.220 79.970 -880.220 ;
        RECT 109.970 -910.220 110.570 -880.220 ;
        RECT 78.170 -910.820 110.570 -910.220 ;
        RECT 117.470 -880.220 149.870 -879.620 ;
        RECT 117.470 -910.220 118.070 -880.220 ;
        RECT 148.070 -910.220 149.870 -880.220 ;
        RECT 117.470 -910.820 149.870 -910.220 ;
        RECT 153.170 -880.220 185.570 -879.620 ;
        RECT 153.170 -910.220 154.970 -880.220 ;
        RECT 184.970 -910.220 185.570 -880.220 ;
        RECT 153.170 -910.820 185.570 -910.220 ;
        RECT 192.470 -880.220 224.870 -879.620 ;
        RECT 192.470 -910.220 193.070 -880.220 ;
        RECT 223.070 -910.220 224.870 -880.220 ;
        RECT 192.470 -910.820 224.870 -910.220 ;
        RECT 228.170 -880.220 260.570 -879.620 ;
        RECT 228.170 -910.220 229.970 -880.220 ;
        RECT 259.970 -910.220 260.570 -880.220 ;
        RECT 228.170 -910.820 260.570 -910.220 ;
        RECT 267.470 -880.220 299.870 -879.620 ;
        RECT 267.470 -910.220 268.070 -880.220 ;
        RECT 298.070 -910.220 299.870 -880.220 ;
        RECT 267.470 -910.820 299.870 -910.220 ;
        RECT 303.170 -880.220 335.570 -879.620 ;
        RECT 303.170 -910.220 304.970 -880.220 ;
        RECT 334.970 -910.220 335.570 -880.220 ;
        RECT 303.170 -910.820 335.570 -910.220 ;
        RECT 342.470 -880.220 374.870 -879.620 ;
        RECT 342.470 -910.220 343.070 -880.220 ;
        RECT 373.070 -910.220 374.870 -880.220 ;
        RECT 342.470 -910.820 374.870 -910.220 ;
        RECT 378.170 -880.220 410.570 -879.620 ;
        RECT 378.170 -910.220 379.970 -880.220 ;
        RECT 409.970 -910.220 410.570 -880.220 ;
        RECT 378.170 -910.820 410.570 -910.220 ;
        RECT 417.470 -880.220 449.870 -879.620 ;
        RECT 417.470 -910.220 418.070 -880.220 ;
        RECT 448.070 -910.220 449.870 -880.220 ;
        RECT 417.470 -910.820 449.870 -910.220 ;
        RECT 453.170 -880.220 485.570 -879.620 ;
        RECT 453.170 -910.220 454.970 -880.220 ;
        RECT 484.970 -910.220 485.570 -880.220 ;
        RECT 453.170 -910.820 485.570 -910.220 ;
        RECT 492.470 -880.220 524.870 -879.620 ;
        RECT 492.470 -910.220 493.070 -880.220 ;
        RECT 523.070 -910.220 524.870 -880.220 ;
        RECT 492.470 -910.820 524.870 -910.220 ;
        RECT 528.170 -880.220 560.570 -879.620 ;
        RECT 528.170 -910.220 529.970 -880.220 ;
        RECT 559.970 -910.220 560.570 -880.220 ;
        RECT 528.170 -910.820 560.570 -910.220 ;
        RECT -557.530 -915.220 -525.130 -914.620 ;
        RECT -557.530 -945.220 -556.930 -915.220 ;
        RECT -526.930 -945.220 -525.130 -915.220 ;
        RECT -557.530 -945.820 -525.130 -945.220 ;
        RECT -521.830 -915.220 -489.430 -914.620 ;
        RECT -521.830 -945.220 -520.030 -915.220 ;
        RECT -490.030 -945.220 -489.430 -915.220 ;
        RECT -521.830 -945.820 -489.430 -945.220 ;
        RECT -482.530 -915.220 -450.130 -914.620 ;
        RECT -482.530 -945.220 -481.930 -915.220 ;
        RECT -451.930 -945.220 -450.130 -915.220 ;
        RECT -482.530 -945.820 -450.130 -945.220 ;
        RECT -446.830 -915.220 -414.430 -914.620 ;
        RECT -446.830 -945.220 -445.030 -915.220 ;
        RECT -415.030 -945.220 -414.430 -915.220 ;
        RECT -446.830 -945.820 -414.430 -945.220 ;
        RECT -407.530 -915.220 -375.130 -914.620 ;
        RECT -407.530 -945.220 -406.930 -915.220 ;
        RECT -376.930 -945.220 -375.130 -915.220 ;
        RECT -407.530 -945.820 -375.130 -945.220 ;
        RECT -371.830 -915.220 -339.430 -914.620 ;
        RECT -371.830 -945.220 -370.030 -915.220 ;
        RECT -340.030 -945.220 -339.430 -915.220 ;
        RECT -371.830 -945.820 -339.430 -945.220 ;
        RECT -332.530 -915.220 -300.130 -914.620 ;
        RECT -332.530 -945.220 -331.930 -915.220 ;
        RECT -301.930 -945.220 -300.130 -915.220 ;
        RECT -332.530 -945.820 -300.130 -945.220 ;
        RECT -296.830 -915.220 -264.430 -914.620 ;
        RECT -296.830 -945.220 -295.030 -915.220 ;
        RECT -265.030 -945.220 -264.430 -915.220 ;
        RECT -296.830 -945.820 -264.430 -945.220 ;
        RECT -257.530 -915.220 -225.130 -914.620 ;
        RECT -257.530 -945.220 -256.930 -915.220 ;
        RECT -226.930 -945.220 -225.130 -915.220 ;
        RECT -257.530 -945.820 -225.130 -945.220 ;
        RECT -221.830 -915.220 -189.430 -914.620 ;
        RECT -221.830 -945.220 -220.030 -915.220 ;
        RECT -190.030 -945.220 -189.430 -915.220 ;
        RECT -221.830 -945.820 -189.430 -945.220 ;
        RECT -182.530 -915.220 -150.130 -914.620 ;
        RECT -182.530 -945.220 -181.930 -915.220 ;
        RECT -151.930 -945.220 -150.130 -915.220 ;
        RECT -182.530 -945.820 -150.130 -945.220 ;
        RECT -146.830 -915.220 -114.430 -914.620 ;
        RECT -146.830 -945.220 -145.030 -915.220 ;
        RECT -115.030 -945.220 -114.430 -915.220 ;
        RECT -146.830 -945.820 -114.430 -945.220 ;
        RECT -107.530 -915.220 -75.130 -914.620 ;
        RECT -107.530 -945.220 -106.930 -915.220 ;
        RECT -76.930 -945.220 -75.130 -915.220 ;
        RECT -107.530 -945.820 -75.130 -945.220 ;
        RECT -71.830 -915.220 -39.430 -914.620 ;
        RECT -71.830 -945.220 -70.030 -915.220 ;
        RECT -40.030 -945.220 -39.430 -915.220 ;
        RECT -71.830 -945.820 -39.430 -945.220 ;
        RECT -32.530 -915.220 -0.130 -914.620 ;
        RECT -32.530 -945.220 -31.930 -915.220 ;
        RECT -1.930 -945.220 -0.130 -915.220 ;
        RECT -32.530 -945.820 -0.130 -945.220 ;
        RECT 3.170 -915.220 35.570 -914.620 ;
        RECT 3.170 -945.220 4.970 -915.220 ;
        RECT 34.970 -945.220 35.570 -915.220 ;
        RECT 3.170 -945.820 35.570 -945.220 ;
        RECT 42.470 -915.220 74.870 -914.620 ;
        RECT 42.470 -945.220 43.070 -915.220 ;
        RECT 73.070 -945.220 74.870 -915.220 ;
        RECT 42.470 -945.820 74.870 -945.220 ;
        RECT 78.170 -915.220 110.570 -914.620 ;
        RECT 78.170 -945.220 79.970 -915.220 ;
        RECT 109.970 -945.220 110.570 -915.220 ;
        RECT 78.170 -945.820 110.570 -945.220 ;
        RECT 117.470 -915.220 149.870 -914.620 ;
        RECT 117.470 -945.220 118.070 -915.220 ;
        RECT 148.070 -945.220 149.870 -915.220 ;
        RECT 117.470 -945.820 149.870 -945.220 ;
        RECT 153.170 -915.220 185.570 -914.620 ;
        RECT 153.170 -945.220 154.970 -915.220 ;
        RECT 184.970 -945.220 185.570 -915.220 ;
        RECT 153.170 -945.820 185.570 -945.220 ;
        RECT 192.470 -915.220 224.870 -914.620 ;
        RECT 192.470 -945.220 193.070 -915.220 ;
        RECT 223.070 -945.220 224.870 -915.220 ;
        RECT 192.470 -945.820 224.870 -945.220 ;
        RECT 228.170 -915.220 260.570 -914.620 ;
        RECT 228.170 -945.220 229.970 -915.220 ;
        RECT 259.970 -945.220 260.570 -915.220 ;
        RECT 228.170 -945.820 260.570 -945.220 ;
        RECT 267.470 -915.220 299.870 -914.620 ;
        RECT 267.470 -945.220 268.070 -915.220 ;
        RECT 298.070 -945.220 299.870 -915.220 ;
        RECT 267.470 -945.820 299.870 -945.220 ;
        RECT 303.170 -915.220 335.570 -914.620 ;
        RECT 303.170 -945.220 304.970 -915.220 ;
        RECT 334.970 -945.220 335.570 -915.220 ;
        RECT 303.170 -945.820 335.570 -945.220 ;
        RECT 342.470 -915.220 374.870 -914.620 ;
        RECT 342.470 -945.220 343.070 -915.220 ;
        RECT 373.070 -945.220 374.870 -915.220 ;
        RECT 342.470 -945.820 374.870 -945.220 ;
        RECT 378.170 -915.220 410.570 -914.620 ;
        RECT 378.170 -945.220 379.970 -915.220 ;
        RECT 409.970 -945.220 410.570 -915.220 ;
        RECT 378.170 -945.820 410.570 -945.220 ;
        RECT 417.470 -915.220 449.870 -914.620 ;
        RECT 417.470 -945.220 418.070 -915.220 ;
        RECT 448.070 -945.220 449.870 -915.220 ;
        RECT 417.470 -945.820 449.870 -945.220 ;
        RECT 453.170 -915.220 485.570 -914.620 ;
        RECT 453.170 -945.220 454.970 -915.220 ;
        RECT 484.970 -945.220 485.570 -915.220 ;
        RECT 453.170 -945.820 485.570 -945.220 ;
        RECT 492.470 -915.220 524.870 -914.620 ;
        RECT 492.470 -945.220 493.070 -915.220 ;
        RECT 523.070 -945.220 524.870 -915.220 ;
        RECT 492.470 -945.820 524.870 -945.220 ;
        RECT 528.170 -915.220 560.570 -914.620 ;
        RECT 528.170 -945.220 529.970 -915.220 ;
        RECT 559.970 -945.220 560.570 -915.220 ;
        RECT 528.170 -945.820 560.570 -945.220 ;
        RECT 763.320 -1085.700 841.320 -352.720 ;
        RECT -838.480 -1163.700 841.320 -1085.700 ;
      LAYER Via4 ;
        RECT -525.800 915.000 -525.520 945.440 ;
        RECT -521.440 915.000 -521.160 945.440 ;
        RECT -450.800 915.000 -450.520 945.440 ;
        RECT -446.440 915.000 -446.160 945.440 ;
        RECT -375.800 915.000 -375.520 945.440 ;
        RECT -371.440 915.000 -371.160 945.440 ;
        RECT -300.800 915.000 -300.520 945.440 ;
        RECT -296.440 915.000 -296.160 945.440 ;
        RECT -225.800 915.000 -225.520 945.440 ;
        RECT -221.440 915.000 -221.160 945.440 ;
        RECT -150.800 915.000 -150.520 945.440 ;
        RECT -146.440 915.000 -146.160 945.440 ;
        RECT -75.800 915.000 -75.520 945.440 ;
        RECT -71.440 915.000 -71.160 945.440 ;
        RECT -0.800 915.000 -0.520 945.440 ;
        RECT 3.560 915.000 3.840 945.440 ;
        RECT 74.200 915.000 74.480 945.440 ;
        RECT 78.560 915.000 78.840 945.440 ;
        RECT 149.200 915.000 149.480 945.440 ;
        RECT 153.560 915.000 153.840 945.440 ;
        RECT 224.200 915.000 224.480 945.440 ;
        RECT 228.560 915.000 228.840 945.440 ;
        RECT 299.200 915.000 299.480 945.440 ;
        RECT 303.560 915.000 303.840 945.440 ;
        RECT 374.200 915.000 374.480 945.440 ;
        RECT 378.560 915.000 378.840 945.440 ;
        RECT 449.200 915.000 449.480 945.440 ;
        RECT 453.560 915.000 453.840 945.440 ;
        RECT 524.200 915.000 524.480 945.440 ;
        RECT 528.560 915.000 528.840 945.440 ;
        RECT -525.800 880.000 -525.520 910.440 ;
        RECT -521.440 880.000 -521.160 910.440 ;
        RECT -450.800 880.000 -450.520 910.440 ;
        RECT -446.440 880.000 -446.160 910.440 ;
        RECT -375.800 880.000 -375.520 910.440 ;
        RECT -371.440 880.000 -371.160 910.440 ;
        RECT -300.800 880.000 -300.520 910.440 ;
        RECT -296.440 880.000 -296.160 910.440 ;
        RECT -225.800 880.000 -225.520 910.440 ;
        RECT -221.440 880.000 -221.160 910.440 ;
        RECT -150.800 880.000 -150.520 910.440 ;
        RECT -146.440 880.000 -146.160 910.440 ;
        RECT -75.800 880.000 -75.520 910.440 ;
        RECT -71.440 880.000 -71.160 910.440 ;
        RECT -0.800 880.000 -0.520 910.440 ;
        RECT 3.560 880.000 3.840 910.440 ;
        RECT 74.200 880.000 74.480 910.440 ;
        RECT 78.560 880.000 78.840 910.440 ;
        RECT 149.200 880.000 149.480 910.440 ;
        RECT 153.560 880.000 153.840 910.440 ;
        RECT 224.200 880.000 224.480 910.440 ;
        RECT 228.560 880.000 228.840 910.440 ;
        RECT 299.200 880.000 299.480 910.440 ;
        RECT 303.560 880.000 303.840 910.440 ;
        RECT 374.200 880.000 374.480 910.440 ;
        RECT 378.560 880.000 378.840 910.440 ;
        RECT 449.200 880.000 449.480 910.440 ;
        RECT 453.560 880.000 453.840 910.440 ;
        RECT 524.200 880.000 524.480 910.440 ;
        RECT 528.560 880.000 528.840 910.440 ;
        RECT -525.800 845.000 -525.520 875.440 ;
        RECT -521.440 845.000 -521.160 875.440 ;
        RECT -450.800 845.000 -450.520 875.440 ;
        RECT -446.440 845.000 -446.160 875.440 ;
        RECT -375.800 845.000 -375.520 875.440 ;
        RECT -371.440 845.000 -371.160 875.440 ;
        RECT -300.800 845.000 -300.520 875.440 ;
        RECT -296.440 845.000 -296.160 875.440 ;
        RECT -225.800 845.000 -225.520 875.440 ;
        RECT -221.440 845.000 -221.160 875.440 ;
        RECT -150.800 845.000 -150.520 875.440 ;
        RECT -146.440 845.000 -146.160 875.440 ;
        RECT -75.800 845.000 -75.520 875.440 ;
        RECT -71.440 845.000 -71.160 875.440 ;
        RECT -0.800 845.000 -0.520 875.440 ;
        RECT 3.560 845.000 3.840 875.440 ;
        RECT 74.200 845.000 74.480 875.440 ;
        RECT 78.560 845.000 78.840 875.440 ;
        RECT 149.200 845.000 149.480 875.440 ;
        RECT 153.560 845.000 153.840 875.440 ;
        RECT 224.200 845.000 224.480 875.440 ;
        RECT 228.560 845.000 228.840 875.440 ;
        RECT 299.200 845.000 299.480 875.440 ;
        RECT 303.560 845.000 303.840 875.440 ;
        RECT 374.200 845.000 374.480 875.440 ;
        RECT 378.560 845.000 378.840 875.440 ;
        RECT 449.200 845.000 449.480 875.440 ;
        RECT 453.560 845.000 453.840 875.440 ;
        RECT 524.200 845.000 524.480 875.440 ;
        RECT 528.560 845.000 528.840 875.440 ;
        RECT -525.800 810.000 -525.520 840.440 ;
        RECT -521.440 810.000 -521.160 840.440 ;
        RECT -450.800 810.000 -450.520 840.440 ;
        RECT -446.440 810.000 -446.160 840.440 ;
        RECT -375.800 810.000 -375.520 840.440 ;
        RECT -371.440 810.000 -371.160 840.440 ;
        RECT -300.800 810.000 -300.520 840.440 ;
        RECT -296.440 810.000 -296.160 840.440 ;
        RECT -225.800 810.000 -225.520 840.440 ;
        RECT -221.440 810.000 -221.160 840.440 ;
        RECT -150.800 810.000 -150.520 840.440 ;
        RECT -146.440 810.000 -146.160 840.440 ;
        RECT -75.800 810.000 -75.520 840.440 ;
        RECT -71.440 810.000 -71.160 840.440 ;
        RECT -0.800 810.000 -0.520 840.440 ;
        RECT 3.560 810.000 3.840 840.440 ;
        RECT 74.200 810.000 74.480 840.440 ;
        RECT 78.560 810.000 78.840 840.440 ;
        RECT 149.200 810.000 149.480 840.440 ;
        RECT 153.560 810.000 153.840 840.440 ;
        RECT 224.200 810.000 224.480 840.440 ;
        RECT 228.560 810.000 228.840 840.440 ;
        RECT 299.200 810.000 299.480 840.440 ;
        RECT 303.560 810.000 303.840 840.440 ;
        RECT 374.200 810.000 374.480 840.440 ;
        RECT 378.560 810.000 378.840 840.440 ;
        RECT 449.200 810.000 449.480 840.440 ;
        RECT 453.560 810.000 453.840 840.440 ;
        RECT 524.200 810.000 524.480 840.440 ;
        RECT 528.560 810.000 528.840 840.440 ;
        RECT -525.800 775.000 -525.520 805.440 ;
        RECT -521.440 775.000 -521.160 805.440 ;
        RECT -450.800 775.000 -450.520 805.440 ;
        RECT -446.440 775.000 -446.160 805.440 ;
        RECT -375.800 775.000 -375.520 805.440 ;
        RECT -371.440 775.000 -371.160 805.440 ;
        RECT -300.800 775.000 -300.520 805.440 ;
        RECT -296.440 775.000 -296.160 805.440 ;
        RECT -225.800 775.000 -225.520 805.440 ;
        RECT -221.440 775.000 -221.160 805.440 ;
        RECT -150.800 775.000 -150.520 805.440 ;
        RECT -146.440 775.000 -146.160 805.440 ;
        RECT -75.800 775.000 -75.520 805.440 ;
        RECT -71.440 775.000 -71.160 805.440 ;
        RECT -0.800 775.000 -0.520 805.440 ;
        RECT 3.560 775.000 3.840 805.440 ;
        RECT 74.200 775.000 74.480 805.440 ;
        RECT 78.560 775.000 78.840 805.440 ;
        RECT 149.200 775.000 149.480 805.440 ;
        RECT 153.560 775.000 153.840 805.440 ;
        RECT 224.200 775.000 224.480 805.440 ;
        RECT 228.560 775.000 228.840 805.440 ;
        RECT 299.200 775.000 299.480 805.440 ;
        RECT 303.560 775.000 303.840 805.440 ;
        RECT 374.200 775.000 374.480 805.440 ;
        RECT 378.560 775.000 378.840 805.440 ;
        RECT 449.200 775.000 449.480 805.440 ;
        RECT 453.560 775.000 453.840 805.440 ;
        RECT 524.200 775.000 524.480 805.440 ;
        RECT 528.560 775.000 528.840 805.440 ;
        RECT -525.800 740.000 -525.520 770.440 ;
        RECT -521.440 740.000 -521.160 770.440 ;
        RECT -450.800 740.000 -450.520 770.440 ;
        RECT -446.440 740.000 -446.160 770.440 ;
        RECT -375.800 740.000 -375.520 770.440 ;
        RECT -371.440 740.000 -371.160 770.440 ;
        RECT -300.800 740.000 -300.520 770.440 ;
        RECT -296.440 740.000 -296.160 770.440 ;
        RECT -225.800 740.000 -225.520 770.440 ;
        RECT -221.440 740.000 -221.160 770.440 ;
        RECT -150.800 740.000 -150.520 770.440 ;
        RECT -146.440 740.000 -146.160 770.440 ;
        RECT -75.800 740.000 -75.520 770.440 ;
        RECT -71.440 740.000 -71.160 770.440 ;
        RECT -0.800 740.000 -0.520 770.440 ;
        RECT 3.560 740.000 3.840 770.440 ;
        RECT 74.200 740.000 74.480 770.440 ;
        RECT 78.560 740.000 78.840 770.440 ;
        RECT 149.200 740.000 149.480 770.440 ;
        RECT 153.560 740.000 153.840 770.440 ;
        RECT 224.200 740.000 224.480 770.440 ;
        RECT 228.560 740.000 228.840 770.440 ;
        RECT 299.200 740.000 299.480 770.440 ;
        RECT 303.560 740.000 303.840 770.440 ;
        RECT 374.200 740.000 374.480 770.440 ;
        RECT 378.560 740.000 378.840 770.440 ;
        RECT 449.200 740.000 449.480 770.440 ;
        RECT 453.560 740.000 453.840 770.440 ;
        RECT 524.200 740.000 524.480 770.440 ;
        RECT 528.560 740.000 528.840 770.440 ;
        RECT -525.800 705.000 -525.520 735.440 ;
        RECT -521.440 705.000 -521.160 735.440 ;
        RECT -450.800 705.000 -450.520 735.440 ;
        RECT -446.440 705.000 -446.160 735.440 ;
        RECT -375.800 705.000 -375.520 735.440 ;
        RECT -371.440 705.000 -371.160 735.440 ;
        RECT -300.800 705.000 -300.520 735.440 ;
        RECT -296.440 705.000 -296.160 735.440 ;
        RECT -225.800 705.000 -225.520 735.440 ;
        RECT -221.440 705.000 -221.160 735.440 ;
        RECT -150.800 705.000 -150.520 735.440 ;
        RECT -146.440 705.000 -146.160 735.440 ;
        RECT -75.800 705.000 -75.520 735.440 ;
        RECT -71.440 705.000 -71.160 735.440 ;
        RECT -0.800 705.000 -0.520 735.440 ;
        RECT 3.560 705.000 3.840 735.440 ;
        RECT 74.200 705.000 74.480 735.440 ;
        RECT 78.560 705.000 78.840 735.440 ;
        RECT 149.200 705.000 149.480 735.440 ;
        RECT 153.560 705.000 153.840 735.440 ;
        RECT 224.200 705.000 224.480 735.440 ;
        RECT 228.560 705.000 228.840 735.440 ;
        RECT 299.200 705.000 299.480 735.440 ;
        RECT 303.560 705.000 303.840 735.440 ;
        RECT 374.200 705.000 374.480 735.440 ;
        RECT 378.560 705.000 378.840 735.440 ;
        RECT 449.200 705.000 449.480 735.440 ;
        RECT 453.560 705.000 453.840 735.440 ;
        RECT 524.200 705.000 524.480 735.440 ;
        RECT 528.560 705.000 528.840 735.440 ;
        RECT -525.800 670.000 -525.520 700.440 ;
        RECT -521.440 670.000 -521.160 700.440 ;
        RECT -450.800 670.000 -450.520 700.440 ;
        RECT -446.440 670.000 -446.160 700.440 ;
        RECT -375.800 670.000 -375.520 700.440 ;
        RECT -371.440 670.000 -371.160 700.440 ;
        RECT -300.800 670.000 -300.520 700.440 ;
        RECT -296.440 670.000 -296.160 700.440 ;
        RECT -225.800 670.000 -225.520 700.440 ;
        RECT -221.440 670.000 -221.160 700.440 ;
        RECT -150.800 670.000 -150.520 700.440 ;
        RECT -146.440 670.000 -146.160 700.440 ;
        RECT -75.800 670.000 -75.520 700.440 ;
        RECT -71.440 670.000 -71.160 700.440 ;
        RECT -0.800 670.000 -0.520 700.440 ;
        RECT 3.560 670.000 3.840 700.440 ;
        RECT 74.200 670.000 74.480 700.440 ;
        RECT 78.560 670.000 78.840 700.440 ;
        RECT 149.200 670.000 149.480 700.440 ;
        RECT 153.560 670.000 153.840 700.440 ;
        RECT 224.200 670.000 224.480 700.440 ;
        RECT 228.560 670.000 228.840 700.440 ;
        RECT 299.200 670.000 299.480 700.440 ;
        RECT 303.560 670.000 303.840 700.440 ;
        RECT 374.200 670.000 374.480 700.440 ;
        RECT 378.560 670.000 378.840 700.440 ;
        RECT 449.200 670.000 449.480 700.440 ;
        RECT 453.560 670.000 453.840 700.440 ;
        RECT 524.200 670.000 524.480 700.440 ;
        RECT 528.560 670.000 528.840 700.440 ;
        RECT -525.800 635.000 -525.520 665.440 ;
        RECT -521.440 635.000 -521.160 665.440 ;
        RECT -450.800 635.000 -450.520 665.440 ;
        RECT -446.440 635.000 -446.160 665.440 ;
        RECT -375.800 635.000 -375.520 665.440 ;
        RECT -371.440 635.000 -371.160 665.440 ;
        RECT -300.800 635.000 -300.520 665.440 ;
        RECT -296.440 635.000 -296.160 665.440 ;
        RECT -225.800 635.000 -225.520 665.440 ;
        RECT -221.440 635.000 -221.160 665.440 ;
        RECT -150.800 635.000 -150.520 665.440 ;
        RECT -146.440 635.000 -146.160 665.440 ;
        RECT -75.800 635.000 -75.520 665.440 ;
        RECT -71.440 635.000 -71.160 665.440 ;
        RECT -0.800 635.000 -0.520 665.440 ;
        RECT 3.560 635.000 3.840 665.440 ;
        RECT 74.200 635.000 74.480 665.440 ;
        RECT 78.560 635.000 78.840 665.440 ;
        RECT 149.200 635.000 149.480 665.440 ;
        RECT 153.560 635.000 153.840 665.440 ;
        RECT 224.200 635.000 224.480 665.440 ;
        RECT 228.560 635.000 228.840 665.440 ;
        RECT 299.200 635.000 299.480 665.440 ;
        RECT 303.560 635.000 303.840 665.440 ;
        RECT 374.200 635.000 374.480 665.440 ;
        RECT 378.560 635.000 378.840 665.440 ;
        RECT 449.200 635.000 449.480 665.440 ;
        RECT 453.560 635.000 453.840 665.440 ;
        RECT 524.200 635.000 524.480 665.440 ;
        RECT 528.560 635.000 528.840 665.440 ;
        RECT -525.800 600.000 -525.520 630.440 ;
        RECT -521.440 600.000 -521.160 630.440 ;
        RECT -450.800 600.000 -450.520 630.440 ;
        RECT -446.440 600.000 -446.160 630.440 ;
        RECT -375.800 600.000 -375.520 630.440 ;
        RECT -371.440 600.000 -371.160 630.440 ;
        RECT -300.800 600.000 -300.520 630.440 ;
        RECT -296.440 600.000 -296.160 630.440 ;
        RECT -225.800 600.000 -225.520 630.440 ;
        RECT -221.440 600.000 -221.160 630.440 ;
        RECT -150.800 600.000 -150.520 630.440 ;
        RECT -146.440 600.000 -146.160 630.440 ;
        RECT -75.800 600.000 -75.520 630.440 ;
        RECT -71.440 600.000 -71.160 630.440 ;
        RECT -0.800 600.000 -0.520 630.440 ;
        RECT 3.560 600.000 3.840 630.440 ;
        RECT 74.200 600.000 74.480 630.440 ;
        RECT 78.560 600.000 78.840 630.440 ;
        RECT 149.200 600.000 149.480 630.440 ;
        RECT 153.560 600.000 153.840 630.440 ;
        RECT 224.200 600.000 224.480 630.440 ;
        RECT 228.560 600.000 228.840 630.440 ;
        RECT 299.200 600.000 299.480 630.440 ;
        RECT 303.560 600.000 303.840 630.440 ;
        RECT 374.200 600.000 374.480 630.440 ;
        RECT 378.560 600.000 378.840 630.440 ;
        RECT 449.200 600.000 449.480 630.440 ;
        RECT 453.560 600.000 453.840 630.440 ;
        RECT 524.200 600.000 524.480 630.440 ;
        RECT 528.560 600.000 528.840 630.440 ;
        RECT -525.800 565.000 -525.520 595.440 ;
        RECT -521.440 565.000 -521.160 595.440 ;
        RECT -450.800 565.000 -450.520 595.440 ;
        RECT -446.440 565.000 -446.160 595.440 ;
        RECT -375.800 565.000 -375.520 595.440 ;
        RECT -371.440 565.000 -371.160 595.440 ;
        RECT -300.800 565.000 -300.520 595.440 ;
        RECT -296.440 565.000 -296.160 595.440 ;
        RECT -225.800 565.000 -225.520 595.440 ;
        RECT -221.440 565.000 -221.160 595.440 ;
        RECT -150.800 565.000 -150.520 595.440 ;
        RECT -146.440 565.000 -146.160 595.440 ;
        RECT -75.800 565.000 -75.520 595.440 ;
        RECT -71.440 565.000 -71.160 595.440 ;
        RECT -0.800 565.000 -0.520 595.440 ;
        RECT 3.560 565.000 3.840 595.440 ;
        RECT 74.200 565.000 74.480 595.440 ;
        RECT 78.560 565.000 78.840 595.440 ;
        RECT 149.200 565.000 149.480 595.440 ;
        RECT 153.560 565.000 153.840 595.440 ;
        RECT 224.200 565.000 224.480 595.440 ;
        RECT 228.560 565.000 228.840 595.440 ;
        RECT 299.200 565.000 299.480 595.440 ;
        RECT 303.560 565.000 303.840 595.440 ;
        RECT 374.200 565.000 374.480 595.440 ;
        RECT 378.560 565.000 378.840 595.440 ;
        RECT 449.200 565.000 449.480 595.440 ;
        RECT 453.560 565.000 453.840 595.440 ;
        RECT 524.200 565.000 524.480 595.440 ;
        RECT 528.560 565.000 528.840 595.440 ;
        RECT -525.800 530.000 -525.520 560.440 ;
        RECT -521.440 530.000 -521.160 560.440 ;
        RECT -450.800 530.000 -450.520 560.440 ;
        RECT -446.440 530.000 -446.160 560.440 ;
        RECT -375.800 530.000 -375.520 560.440 ;
        RECT -371.440 530.000 -371.160 560.440 ;
        RECT -300.800 530.000 -300.520 560.440 ;
        RECT -296.440 530.000 -296.160 560.440 ;
        RECT -225.800 530.000 -225.520 560.440 ;
        RECT -221.440 530.000 -221.160 560.440 ;
        RECT -150.800 530.000 -150.520 560.440 ;
        RECT -146.440 530.000 -146.160 560.440 ;
        RECT -75.800 530.000 -75.520 560.440 ;
        RECT -71.440 530.000 -71.160 560.440 ;
        RECT -0.800 530.000 -0.520 560.440 ;
        RECT 3.560 530.000 3.840 560.440 ;
        RECT 74.200 530.000 74.480 560.440 ;
        RECT 78.560 530.000 78.840 560.440 ;
        RECT 149.200 530.000 149.480 560.440 ;
        RECT 153.560 530.000 153.840 560.440 ;
        RECT 224.200 530.000 224.480 560.440 ;
        RECT 228.560 530.000 228.840 560.440 ;
        RECT 299.200 530.000 299.480 560.440 ;
        RECT 303.560 530.000 303.840 560.440 ;
        RECT 374.200 530.000 374.480 560.440 ;
        RECT 378.560 530.000 378.840 560.440 ;
        RECT 449.200 530.000 449.480 560.440 ;
        RECT 453.560 530.000 453.840 560.440 ;
        RECT 524.200 530.000 524.480 560.440 ;
        RECT 528.560 530.000 528.840 560.440 ;
        RECT -525.800 495.000 -525.520 525.440 ;
        RECT -521.440 495.000 -521.160 525.440 ;
        RECT -450.800 495.000 -450.520 525.440 ;
        RECT -446.440 495.000 -446.160 525.440 ;
        RECT -375.800 495.000 -375.520 525.440 ;
        RECT -371.440 495.000 -371.160 525.440 ;
        RECT -300.800 495.000 -300.520 525.440 ;
        RECT -296.440 495.000 -296.160 525.440 ;
        RECT -225.800 495.000 -225.520 525.440 ;
        RECT -221.440 495.000 -221.160 525.440 ;
        RECT -150.800 495.000 -150.520 525.440 ;
        RECT -146.440 495.000 -146.160 525.440 ;
        RECT -75.800 495.000 -75.520 525.440 ;
        RECT -71.440 495.000 -71.160 525.440 ;
        RECT -0.800 495.000 -0.520 525.440 ;
        RECT 3.560 495.000 3.840 525.440 ;
        RECT 74.200 495.000 74.480 525.440 ;
        RECT 78.560 495.000 78.840 525.440 ;
        RECT 149.200 495.000 149.480 525.440 ;
        RECT 153.560 495.000 153.840 525.440 ;
        RECT 224.200 495.000 224.480 525.440 ;
        RECT 228.560 495.000 228.840 525.440 ;
        RECT 299.200 495.000 299.480 525.440 ;
        RECT 303.560 495.000 303.840 525.440 ;
        RECT 374.200 495.000 374.480 525.440 ;
        RECT 378.560 495.000 378.840 525.440 ;
        RECT 449.200 495.000 449.480 525.440 ;
        RECT 453.560 495.000 453.840 525.440 ;
        RECT 524.200 495.000 524.480 525.440 ;
        RECT 528.560 495.000 528.840 525.440 ;
        RECT -525.800 460.000 -525.520 490.440 ;
        RECT -521.440 460.000 -521.160 490.440 ;
        RECT -450.800 460.000 -450.520 490.440 ;
        RECT -446.440 460.000 -446.160 490.440 ;
        RECT -375.800 460.000 -375.520 490.440 ;
        RECT -371.440 460.000 -371.160 490.440 ;
        RECT -300.800 460.000 -300.520 490.440 ;
        RECT -296.440 460.000 -296.160 490.440 ;
        RECT -225.800 460.000 -225.520 490.440 ;
        RECT -221.440 460.000 -221.160 490.440 ;
        RECT -150.800 460.000 -150.520 490.440 ;
        RECT -146.440 460.000 -146.160 490.440 ;
        RECT -75.800 460.000 -75.520 490.440 ;
        RECT -71.440 460.000 -71.160 490.440 ;
        RECT -0.800 460.000 -0.520 490.440 ;
        RECT 3.560 460.000 3.840 490.440 ;
        RECT 74.200 460.000 74.480 490.440 ;
        RECT 78.560 460.000 78.840 490.440 ;
        RECT 149.200 460.000 149.480 490.440 ;
        RECT 153.560 460.000 153.840 490.440 ;
        RECT 224.200 460.000 224.480 490.440 ;
        RECT 228.560 460.000 228.840 490.440 ;
        RECT 299.200 460.000 299.480 490.440 ;
        RECT 303.560 460.000 303.840 490.440 ;
        RECT 374.200 460.000 374.480 490.440 ;
        RECT 378.560 460.000 378.840 490.440 ;
        RECT 449.200 460.000 449.480 490.440 ;
        RECT 453.560 460.000 453.840 490.440 ;
        RECT 524.200 460.000 524.480 490.440 ;
        RECT 528.560 460.000 528.840 490.440 ;
        RECT -525.800 425.000 -525.520 455.440 ;
        RECT -521.440 425.000 -521.160 455.440 ;
        RECT -450.800 425.000 -450.520 455.440 ;
        RECT -446.440 425.000 -446.160 455.440 ;
        RECT -375.800 425.000 -375.520 455.440 ;
        RECT -371.440 425.000 -371.160 455.440 ;
        RECT -300.800 425.000 -300.520 455.440 ;
        RECT -296.440 425.000 -296.160 455.440 ;
        RECT -225.800 425.000 -225.520 455.440 ;
        RECT -221.440 425.000 -221.160 455.440 ;
        RECT -150.800 425.000 -150.520 455.440 ;
        RECT -146.440 425.000 -146.160 455.440 ;
        RECT -75.800 425.000 -75.520 455.440 ;
        RECT -71.440 425.000 -71.160 455.440 ;
        RECT -0.800 425.000 -0.520 455.440 ;
        RECT 3.560 425.000 3.840 455.440 ;
        RECT 74.200 425.000 74.480 455.440 ;
        RECT 78.560 425.000 78.840 455.440 ;
        RECT 149.200 425.000 149.480 455.440 ;
        RECT 153.560 425.000 153.840 455.440 ;
        RECT 224.200 425.000 224.480 455.440 ;
        RECT 228.560 425.000 228.840 455.440 ;
        RECT 299.200 425.000 299.480 455.440 ;
        RECT 303.560 425.000 303.840 455.440 ;
        RECT 374.200 425.000 374.480 455.440 ;
        RECT 378.560 425.000 378.840 455.440 ;
        RECT 449.200 425.000 449.480 455.440 ;
        RECT 453.560 425.000 453.840 455.440 ;
        RECT 524.200 425.000 524.480 455.440 ;
        RECT 528.560 425.000 528.840 455.440 ;
        RECT -525.800 390.000 -525.520 420.440 ;
        RECT -521.440 390.000 -521.160 420.440 ;
        RECT -450.800 390.000 -450.520 420.440 ;
        RECT -446.440 390.000 -446.160 420.440 ;
        RECT -375.800 390.000 -375.520 420.440 ;
        RECT -371.440 390.000 -371.160 420.440 ;
        RECT -300.800 390.000 -300.520 420.440 ;
        RECT -296.440 390.000 -296.160 420.440 ;
        RECT -225.800 390.000 -225.520 420.440 ;
        RECT -221.440 390.000 -221.160 420.440 ;
        RECT -150.800 390.000 -150.520 420.440 ;
        RECT -146.440 390.000 -146.160 420.440 ;
        RECT -75.800 390.000 -75.520 420.440 ;
        RECT -71.440 390.000 -71.160 420.440 ;
        RECT -0.800 390.000 -0.520 420.440 ;
        RECT 3.560 390.000 3.840 420.440 ;
        RECT 74.200 390.000 74.480 420.440 ;
        RECT 78.560 390.000 78.840 420.440 ;
        RECT 149.200 390.000 149.480 420.440 ;
        RECT 153.560 390.000 153.840 420.440 ;
        RECT 224.200 390.000 224.480 420.440 ;
        RECT 228.560 390.000 228.840 420.440 ;
        RECT 299.200 390.000 299.480 420.440 ;
        RECT 303.560 390.000 303.840 420.440 ;
        RECT 374.200 390.000 374.480 420.440 ;
        RECT 378.560 390.000 378.840 420.440 ;
        RECT 449.200 390.000 449.480 420.440 ;
        RECT 453.560 390.000 453.840 420.440 ;
        RECT 524.200 390.000 524.480 420.440 ;
        RECT 528.560 390.000 528.840 420.440 ;
        RECT -573.280 321.640 -572.480 352.600 ;
        RECT -572.080 321.640 -571.280 352.600 ;
        RECT -570.880 321.640 -570.080 352.600 ;
        RECT -569.680 321.640 -568.880 352.600 ;
        RECT -568.480 321.640 -567.680 352.600 ;
        RECT -567.280 321.640 -566.480 352.600 ;
        RECT -566.080 321.640 -565.280 352.600 ;
        RECT -564.880 321.640 -564.080 352.600 ;
        RECT -563.680 321.640 -562.880 352.600 ;
        RECT -562.480 321.640 -561.680 352.600 ;
        RECT -561.280 321.640 -560.480 352.600 ;
        RECT -560.080 321.640 -559.280 352.600 ;
        RECT -558.880 321.640 -558.080 352.600 ;
        RECT -557.680 321.640 -556.880 352.600 ;
        RECT -556.480 321.640 -555.680 352.600 ;
        RECT -555.280 321.640 -554.480 352.600 ;
        RECT -554.080 321.640 -553.280 352.600 ;
        RECT -552.880 321.640 -552.080 352.600 ;
        RECT -551.680 321.640 -550.880 352.600 ;
        RECT -550.480 321.640 -549.680 352.600 ;
        RECT -549.280 321.640 -548.480 352.600 ;
        RECT -548.080 321.640 -547.280 352.600 ;
        RECT -546.880 321.640 -546.080 352.600 ;
        RECT -545.680 321.640 -544.880 352.600 ;
        RECT -544.480 321.640 -543.680 352.600 ;
        RECT 546.720 321.640 547.520 352.600 ;
        RECT 547.920 321.640 548.720 352.600 ;
        RECT 549.120 321.640 549.920 352.600 ;
        RECT 550.320 321.640 551.120 352.600 ;
        RECT 551.520 321.640 552.320 352.600 ;
        RECT 552.720 321.640 553.520 352.600 ;
        RECT 553.920 321.640 554.720 352.600 ;
        RECT 555.120 321.640 555.920 352.600 ;
        RECT 556.320 321.640 557.120 352.600 ;
        RECT 557.520 321.640 558.320 352.600 ;
        RECT 558.720 321.640 559.520 352.600 ;
        RECT 559.920 321.640 560.720 352.600 ;
        RECT 561.120 321.640 561.920 352.600 ;
        RECT 562.320 321.640 563.120 352.600 ;
        RECT 563.520 321.640 564.320 352.600 ;
        RECT 564.720 321.640 565.520 352.600 ;
        RECT 565.920 321.640 566.720 352.600 ;
        RECT 567.120 321.640 567.920 352.600 ;
        RECT 568.320 321.640 569.120 352.600 ;
        RECT 569.520 321.640 570.320 352.600 ;
        RECT 570.720 321.640 571.520 352.600 ;
        RECT 571.920 321.640 572.720 352.600 ;
        RECT 573.120 321.640 573.920 352.600 ;
        RECT 574.320 321.640 575.120 352.600 ;
        RECT 575.520 321.640 576.320 352.600 ;
        RECT -431.650 220.860 -431.370 320.980 ;
        RECT -425.590 220.860 -425.310 320.980 ;
        RECT -216.650 220.860 -216.370 320.980 ;
        RECT -210.590 220.860 -210.310 320.980 ;
        RECT -1.650 220.860 -1.370 320.980 ;
        RECT 4.410 220.860 4.690 320.980 ;
        RECT 213.350 220.860 213.630 320.980 ;
        RECT 219.410 220.860 219.690 320.980 ;
        RECT 428.350 220.860 428.630 320.980 ;
        RECT 434.410 220.860 434.690 320.980 ;
        RECT -573.280 172.600 -572.480 192.640 ;
        RECT -572.080 172.600 -571.280 192.640 ;
        RECT -570.880 172.600 -570.080 192.640 ;
        RECT -569.680 172.600 -568.880 192.640 ;
        RECT -568.480 172.600 -567.680 192.640 ;
        RECT -567.280 172.600 -566.480 192.640 ;
        RECT -566.080 172.600 -565.280 192.640 ;
        RECT -564.880 172.600 -564.080 192.640 ;
        RECT -563.680 172.600 -562.880 192.640 ;
        RECT -562.480 172.600 -561.680 192.640 ;
        RECT -561.280 172.600 -560.480 192.640 ;
        RECT -560.080 172.600 -559.280 192.640 ;
        RECT -558.880 172.600 -558.080 192.640 ;
        RECT -557.680 172.600 -556.880 192.640 ;
        RECT -556.480 172.600 -555.680 192.640 ;
        RECT -555.280 172.600 -554.480 192.640 ;
        RECT -554.080 172.600 -553.280 192.640 ;
        RECT -552.880 172.600 -552.080 192.640 ;
        RECT -551.680 172.600 -550.880 192.640 ;
        RECT -550.480 172.600 -549.680 192.640 ;
        RECT -549.280 172.600 -548.480 192.640 ;
        RECT -548.080 172.600 -547.280 192.640 ;
        RECT -546.880 172.600 -546.080 192.640 ;
        RECT -545.680 172.600 -544.880 192.640 ;
        RECT -544.480 172.600 -543.680 192.640 ;
        RECT -509.300 172.560 -478.860 172.840 ;
        RECT -469.300 172.560 -438.860 172.840 ;
        RECT -429.300 172.560 -398.860 172.840 ;
        RECT -389.300 172.560 -358.860 172.840 ;
        RECT -349.300 172.560 -318.860 172.840 ;
        RECT -309.300 172.560 -278.860 172.840 ;
        RECT -269.300 172.560 -238.860 172.840 ;
        RECT -229.300 172.560 -198.860 172.840 ;
        RECT -189.300 172.560 -158.860 172.840 ;
        RECT -149.300 172.560 -118.860 172.840 ;
        RECT -109.300 172.560 -78.860 172.840 ;
        RECT -69.300 172.560 -38.860 172.840 ;
        RECT -29.300 172.560 1.140 172.840 ;
        RECT 10.700 172.560 41.140 172.840 ;
        RECT 50.700 172.560 81.140 172.840 ;
        RECT 90.700 172.560 121.140 172.840 ;
        RECT 130.700 172.560 161.140 172.840 ;
        RECT 170.700 172.560 201.140 172.840 ;
        RECT 226.300 172.560 256.740 172.840 ;
        RECT 266.300 172.560 296.740 172.840 ;
        RECT 306.300 172.560 336.740 172.840 ;
        RECT 346.300 172.560 376.740 172.840 ;
        RECT 386.300 172.560 416.740 172.840 ;
        RECT 426.300 172.560 456.740 172.840 ;
        RECT 466.300 172.560 496.740 172.840 ;
        RECT 546.720 172.600 547.520 192.640 ;
        RECT 547.920 172.600 548.720 192.640 ;
        RECT 549.120 172.600 549.920 192.640 ;
        RECT 550.320 172.600 551.120 192.640 ;
        RECT 551.520 172.600 552.320 192.640 ;
        RECT 552.720 172.600 553.520 192.640 ;
        RECT 553.920 172.600 554.720 192.640 ;
        RECT 555.120 172.600 555.920 192.640 ;
        RECT 556.320 172.600 557.120 192.640 ;
        RECT 557.520 172.600 558.320 192.640 ;
        RECT 558.720 172.600 559.520 192.640 ;
        RECT 559.920 172.600 560.720 192.640 ;
        RECT 561.120 172.600 561.920 192.640 ;
        RECT 562.320 172.600 563.120 192.640 ;
        RECT 563.520 172.600 564.320 192.640 ;
        RECT 564.720 172.600 565.520 192.640 ;
        RECT 565.920 172.600 566.720 192.640 ;
        RECT 567.120 172.600 567.920 192.640 ;
        RECT 568.320 172.600 569.120 192.640 ;
        RECT 569.520 172.600 570.320 192.640 ;
        RECT 570.720 172.600 571.520 192.640 ;
        RECT 571.920 172.600 572.720 192.640 ;
        RECT 573.120 172.600 573.920 192.640 ;
        RECT 574.320 172.600 575.120 192.640 ;
        RECT 575.520 172.600 576.320 192.640 ;
        RECT -573.280 -192.640 -572.480 -172.600 ;
        RECT -572.080 -192.640 -571.280 -172.600 ;
        RECT -570.880 -192.640 -570.080 -172.600 ;
        RECT -569.680 -192.640 -568.880 -172.600 ;
        RECT -568.480 -192.640 -567.680 -172.600 ;
        RECT -567.280 -192.640 -566.480 -172.600 ;
        RECT -566.080 -192.640 -565.280 -172.600 ;
        RECT -564.880 -192.640 -564.080 -172.600 ;
        RECT -563.680 -192.640 -562.880 -172.600 ;
        RECT -562.480 -192.640 -561.680 -172.600 ;
        RECT -561.280 -192.640 -560.480 -172.600 ;
        RECT -560.080 -192.640 -559.280 -172.600 ;
        RECT -558.880 -192.640 -558.080 -172.600 ;
        RECT -557.680 -192.640 -556.880 -172.600 ;
        RECT -556.480 -192.640 -555.680 -172.600 ;
        RECT -555.280 -192.640 -554.480 -172.600 ;
        RECT -554.080 -192.640 -553.280 -172.600 ;
        RECT -552.880 -192.640 -552.080 -172.600 ;
        RECT -551.680 -192.640 -550.880 -172.600 ;
        RECT -550.480 -192.640 -549.680 -172.600 ;
        RECT -549.280 -192.640 -548.480 -172.600 ;
        RECT -548.080 -192.640 -547.280 -172.600 ;
        RECT -546.880 -192.640 -546.080 -172.600 ;
        RECT -545.680 -192.640 -544.880 -172.600 ;
        RECT -544.480 -192.640 -543.680 -172.600 ;
        RECT -509.300 -172.840 -478.860 -172.560 ;
        RECT -469.300 -172.840 -438.860 -172.560 ;
        RECT -429.300 -172.840 -398.860 -172.560 ;
        RECT -389.300 -172.840 -358.860 -172.560 ;
        RECT -349.300 -172.840 -318.860 -172.560 ;
        RECT -309.300 -172.840 -278.860 -172.560 ;
        RECT -269.300 -172.840 -238.860 -172.560 ;
        RECT -229.300 -172.840 -198.860 -172.560 ;
        RECT -189.300 -172.840 -158.860 -172.560 ;
        RECT -149.300 -172.840 -118.860 -172.560 ;
        RECT -109.300 -172.840 -78.860 -172.560 ;
        RECT -69.300 -172.840 -38.860 -172.560 ;
        RECT -29.300 -172.840 1.140 -172.560 ;
        RECT 10.700 -172.840 41.140 -172.560 ;
        RECT 50.700 -172.840 81.140 -172.560 ;
        RECT 90.700 -172.840 121.140 -172.560 ;
        RECT 130.700 -172.840 161.140 -172.560 ;
        RECT 170.700 -172.840 201.140 -172.560 ;
        RECT 226.300 -172.840 256.740 -172.560 ;
        RECT 266.300 -172.840 296.740 -172.560 ;
        RECT 306.300 -172.840 336.740 -172.560 ;
        RECT 346.300 -172.840 376.740 -172.560 ;
        RECT 386.300 -172.840 416.740 -172.560 ;
        RECT 426.300 -172.840 456.740 -172.560 ;
        RECT 466.300 -172.840 496.740 -172.560 ;
        RECT 546.720 -192.640 547.520 -172.600 ;
        RECT 547.920 -192.640 548.720 -172.600 ;
        RECT 549.120 -192.640 549.920 -172.600 ;
        RECT 550.320 -192.640 551.120 -172.600 ;
        RECT 551.520 -192.640 552.320 -172.600 ;
        RECT 552.720 -192.640 553.520 -172.600 ;
        RECT 553.920 -192.640 554.720 -172.600 ;
        RECT 555.120 -192.640 555.920 -172.600 ;
        RECT 556.320 -192.640 557.120 -172.600 ;
        RECT 557.520 -192.640 558.320 -172.600 ;
        RECT 558.720 -192.640 559.520 -172.600 ;
        RECT 559.920 -192.640 560.720 -172.600 ;
        RECT 561.120 -192.640 561.920 -172.600 ;
        RECT 562.320 -192.640 563.120 -172.600 ;
        RECT 563.520 -192.640 564.320 -172.600 ;
        RECT 564.720 -192.640 565.520 -172.600 ;
        RECT 565.920 -192.640 566.720 -172.600 ;
        RECT 567.120 -192.640 567.920 -172.600 ;
        RECT 568.320 -192.640 569.120 -172.600 ;
        RECT 569.520 -192.640 570.320 -172.600 ;
        RECT 570.720 -192.640 571.520 -172.600 ;
        RECT 571.920 -192.640 572.720 -172.600 ;
        RECT 573.120 -192.640 573.920 -172.600 ;
        RECT 574.320 -192.640 575.120 -172.600 ;
        RECT 575.520 -192.640 576.320 -172.600 ;
        RECT -431.650 -320.980 -431.370 -220.860 ;
        RECT -425.590 -320.980 -425.310 -220.860 ;
        RECT -216.650 -320.980 -216.370 -220.860 ;
        RECT -210.590 -320.980 -210.310 -220.860 ;
        RECT -1.650 -320.980 -1.370 -220.860 ;
        RECT 4.410 -320.980 4.690 -220.860 ;
        RECT 213.350 -320.980 213.630 -220.860 ;
        RECT 219.410 -320.980 219.690 -220.860 ;
        RECT 428.350 -320.980 428.630 -220.860 ;
        RECT 434.410 -320.980 434.690 -220.860 ;
        RECT -573.280 -352.600 -572.480 -321.640 ;
        RECT -572.080 -352.600 -571.280 -321.640 ;
        RECT -570.880 -352.600 -570.080 -321.640 ;
        RECT -569.680 -352.600 -568.880 -321.640 ;
        RECT -568.480 -352.600 -567.680 -321.640 ;
        RECT -567.280 -352.600 -566.480 -321.640 ;
        RECT -566.080 -352.600 -565.280 -321.640 ;
        RECT -564.880 -352.600 -564.080 -321.640 ;
        RECT -563.680 -352.600 -562.880 -321.640 ;
        RECT -562.480 -352.600 -561.680 -321.640 ;
        RECT -561.280 -352.600 -560.480 -321.640 ;
        RECT -560.080 -352.600 -559.280 -321.640 ;
        RECT -558.880 -352.600 -558.080 -321.640 ;
        RECT -557.680 -352.600 -556.880 -321.640 ;
        RECT -556.480 -352.600 -555.680 -321.640 ;
        RECT -555.280 -352.600 -554.480 -321.640 ;
        RECT -554.080 -352.600 -553.280 -321.640 ;
        RECT -552.880 -352.600 -552.080 -321.640 ;
        RECT -551.680 -352.600 -550.880 -321.640 ;
        RECT -550.480 -352.600 -549.680 -321.640 ;
        RECT -549.280 -352.600 -548.480 -321.640 ;
        RECT -548.080 -352.600 -547.280 -321.640 ;
        RECT -546.880 -352.600 -546.080 -321.640 ;
        RECT -545.680 -352.600 -544.880 -321.640 ;
        RECT -544.480 -352.600 -543.680 -321.640 ;
        RECT 546.720 -352.600 547.520 -321.640 ;
        RECT 547.920 -352.600 548.720 -321.640 ;
        RECT 549.120 -352.600 549.920 -321.640 ;
        RECT 550.320 -352.600 551.120 -321.640 ;
        RECT 551.520 -352.600 552.320 -321.640 ;
        RECT 552.720 -352.600 553.520 -321.640 ;
        RECT 553.920 -352.600 554.720 -321.640 ;
        RECT 555.120 -352.600 555.920 -321.640 ;
        RECT 556.320 -352.600 557.120 -321.640 ;
        RECT 557.520 -352.600 558.320 -321.640 ;
        RECT 558.720 -352.600 559.520 -321.640 ;
        RECT 559.920 -352.600 560.720 -321.640 ;
        RECT 561.120 -352.600 561.920 -321.640 ;
        RECT 562.320 -352.600 563.120 -321.640 ;
        RECT 563.520 -352.600 564.320 -321.640 ;
        RECT 564.720 -352.600 565.520 -321.640 ;
        RECT 565.920 -352.600 566.720 -321.640 ;
        RECT 567.120 -352.600 567.920 -321.640 ;
        RECT 568.320 -352.600 569.120 -321.640 ;
        RECT 569.520 -352.600 570.320 -321.640 ;
        RECT 570.720 -352.600 571.520 -321.640 ;
        RECT 571.920 -352.600 572.720 -321.640 ;
        RECT 573.120 -352.600 573.920 -321.640 ;
        RECT 574.320 -352.600 575.120 -321.640 ;
        RECT 575.520 -352.600 576.320 -321.640 ;
        RECT -525.800 -420.440 -525.520 -390.000 ;
        RECT -521.440 -420.440 -521.160 -390.000 ;
        RECT -450.800 -420.440 -450.520 -390.000 ;
        RECT -446.440 -420.440 -446.160 -390.000 ;
        RECT -375.800 -420.440 -375.520 -390.000 ;
        RECT -371.440 -420.440 -371.160 -390.000 ;
        RECT -300.800 -420.440 -300.520 -390.000 ;
        RECT -296.440 -420.440 -296.160 -390.000 ;
        RECT -225.800 -420.440 -225.520 -390.000 ;
        RECT -221.440 -420.440 -221.160 -390.000 ;
        RECT -150.800 -420.440 -150.520 -390.000 ;
        RECT -146.440 -420.440 -146.160 -390.000 ;
        RECT -75.800 -420.440 -75.520 -390.000 ;
        RECT -71.440 -420.440 -71.160 -390.000 ;
        RECT -0.800 -420.440 -0.520 -390.000 ;
        RECT 3.560 -420.440 3.840 -390.000 ;
        RECT 74.200 -420.440 74.480 -390.000 ;
        RECT 78.560 -420.440 78.840 -390.000 ;
        RECT 149.200 -420.440 149.480 -390.000 ;
        RECT 153.560 -420.440 153.840 -390.000 ;
        RECT 224.200 -420.440 224.480 -390.000 ;
        RECT 228.560 -420.440 228.840 -390.000 ;
        RECT 299.200 -420.440 299.480 -390.000 ;
        RECT 303.560 -420.440 303.840 -390.000 ;
        RECT 374.200 -420.440 374.480 -390.000 ;
        RECT 378.560 -420.440 378.840 -390.000 ;
        RECT 449.200 -420.440 449.480 -390.000 ;
        RECT 453.560 -420.440 453.840 -390.000 ;
        RECT 524.200 -420.440 524.480 -390.000 ;
        RECT 528.560 -420.440 528.840 -390.000 ;
        RECT -525.800 -455.440 -525.520 -425.000 ;
        RECT -521.440 -455.440 -521.160 -425.000 ;
        RECT -450.800 -455.440 -450.520 -425.000 ;
        RECT -446.440 -455.440 -446.160 -425.000 ;
        RECT -375.800 -455.440 -375.520 -425.000 ;
        RECT -371.440 -455.440 -371.160 -425.000 ;
        RECT -300.800 -455.440 -300.520 -425.000 ;
        RECT -296.440 -455.440 -296.160 -425.000 ;
        RECT -225.800 -455.440 -225.520 -425.000 ;
        RECT -221.440 -455.440 -221.160 -425.000 ;
        RECT -150.800 -455.440 -150.520 -425.000 ;
        RECT -146.440 -455.440 -146.160 -425.000 ;
        RECT -75.800 -455.440 -75.520 -425.000 ;
        RECT -71.440 -455.440 -71.160 -425.000 ;
        RECT -0.800 -455.440 -0.520 -425.000 ;
        RECT 3.560 -455.440 3.840 -425.000 ;
        RECT 74.200 -455.440 74.480 -425.000 ;
        RECT 78.560 -455.440 78.840 -425.000 ;
        RECT 149.200 -455.440 149.480 -425.000 ;
        RECT 153.560 -455.440 153.840 -425.000 ;
        RECT 224.200 -455.440 224.480 -425.000 ;
        RECT 228.560 -455.440 228.840 -425.000 ;
        RECT 299.200 -455.440 299.480 -425.000 ;
        RECT 303.560 -455.440 303.840 -425.000 ;
        RECT 374.200 -455.440 374.480 -425.000 ;
        RECT 378.560 -455.440 378.840 -425.000 ;
        RECT 449.200 -455.440 449.480 -425.000 ;
        RECT 453.560 -455.440 453.840 -425.000 ;
        RECT 524.200 -455.440 524.480 -425.000 ;
        RECT 528.560 -455.440 528.840 -425.000 ;
        RECT -525.800 -490.440 -525.520 -460.000 ;
        RECT -521.440 -490.440 -521.160 -460.000 ;
        RECT -450.800 -490.440 -450.520 -460.000 ;
        RECT -446.440 -490.440 -446.160 -460.000 ;
        RECT -375.800 -490.440 -375.520 -460.000 ;
        RECT -371.440 -490.440 -371.160 -460.000 ;
        RECT -300.800 -490.440 -300.520 -460.000 ;
        RECT -296.440 -490.440 -296.160 -460.000 ;
        RECT -225.800 -490.440 -225.520 -460.000 ;
        RECT -221.440 -490.440 -221.160 -460.000 ;
        RECT -150.800 -490.440 -150.520 -460.000 ;
        RECT -146.440 -490.440 -146.160 -460.000 ;
        RECT -75.800 -490.440 -75.520 -460.000 ;
        RECT -71.440 -490.440 -71.160 -460.000 ;
        RECT -0.800 -490.440 -0.520 -460.000 ;
        RECT 3.560 -490.440 3.840 -460.000 ;
        RECT 74.200 -490.440 74.480 -460.000 ;
        RECT 78.560 -490.440 78.840 -460.000 ;
        RECT 149.200 -490.440 149.480 -460.000 ;
        RECT 153.560 -490.440 153.840 -460.000 ;
        RECT 224.200 -490.440 224.480 -460.000 ;
        RECT 228.560 -490.440 228.840 -460.000 ;
        RECT 299.200 -490.440 299.480 -460.000 ;
        RECT 303.560 -490.440 303.840 -460.000 ;
        RECT 374.200 -490.440 374.480 -460.000 ;
        RECT 378.560 -490.440 378.840 -460.000 ;
        RECT 449.200 -490.440 449.480 -460.000 ;
        RECT 453.560 -490.440 453.840 -460.000 ;
        RECT 524.200 -490.440 524.480 -460.000 ;
        RECT 528.560 -490.440 528.840 -460.000 ;
        RECT -525.800 -525.440 -525.520 -495.000 ;
        RECT -521.440 -525.440 -521.160 -495.000 ;
        RECT -450.800 -525.440 -450.520 -495.000 ;
        RECT -446.440 -525.440 -446.160 -495.000 ;
        RECT -375.800 -525.440 -375.520 -495.000 ;
        RECT -371.440 -525.440 -371.160 -495.000 ;
        RECT -300.800 -525.440 -300.520 -495.000 ;
        RECT -296.440 -525.440 -296.160 -495.000 ;
        RECT -225.800 -525.440 -225.520 -495.000 ;
        RECT -221.440 -525.440 -221.160 -495.000 ;
        RECT -150.800 -525.440 -150.520 -495.000 ;
        RECT -146.440 -525.440 -146.160 -495.000 ;
        RECT -75.800 -525.440 -75.520 -495.000 ;
        RECT -71.440 -525.440 -71.160 -495.000 ;
        RECT -0.800 -525.440 -0.520 -495.000 ;
        RECT 3.560 -525.440 3.840 -495.000 ;
        RECT 74.200 -525.440 74.480 -495.000 ;
        RECT 78.560 -525.440 78.840 -495.000 ;
        RECT 149.200 -525.440 149.480 -495.000 ;
        RECT 153.560 -525.440 153.840 -495.000 ;
        RECT 224.200 -525.440 224.480 -495.000 ;
        RECT 228.560 -525.440 228.840 -495.000 ;
        RECT 299.200 -525.440 299.480 -495.000 ;
        RECT 303.560 -525.440 303.840 -495.000 ;
        RECT 374.200 -525.440 374.480 -495.000 ;
        RECT 378.560 -525.440 378.840 -495.000 ;
        RECT 449.200 -525.440 449.480 -495.000 ;
        RECT 453.560 -525.440 453.840 -495.000 ;
        RECT 524.200 -525.440 524.480 -495.000 ;
        RECT 528.560 -525.440 528.840 -495.000 ;
        RECT -525.800 -560.440 -525.520 -530.000 ;
        RECT -521.440 -560.440 -521.160 -530.000 ;
        RECT -450.800 -560.440 -450.520 -530.000 ;
        RECT -446.440 -560.440 -446.160 -530.000 ;
        RECT -375.800 -560.440 -375.520 -530.000 ;
        RECT -371.440 -560.440 -371.160 -530.000 ;
        RECT -300.800 -560.440 -300.520 -530.000 ;
        RECT -296.440 -560.440 -296.160 -530.000 ;
        RECT -225.800 -560.440 -225.520 -530.000 ;
        RECT -221.440 -560.440 -221.160 -530.000 ;
        RECT -150.800 -560.440 -150.520 -530.000 ;
        RECT -146.440 -560.440 -146.160 -530.000 ;
        RECT -75.800 -560.440 -75.520 -530.000 ;
        RECT -71.440 -560.440 -71.160 -530.000 ;
        RECT -0.800 -560.440 -0.520 -530.000 ;
        RECT 3.560 -560.440 3.840 -530.000 ;
        RECT 74.200 -560.440 74.480 -530.000 ;
        RECT 78.560 -560.440 78.840 -530.000 ;
        RECT 149.200 -560.440 149.480 -530.000 ;
        RECT 153.560 -560.440 153.840 -530.000 ;
        RECT 224.200 -560.440 224.480 -530.000 ;
        RECT 228.560 -560.440 228.840 -530.000 ;
        RECT 299.200 -560.440 299.480 -530.000 ;
        RECT 303.560 -560.440 303.840 -530.000 ;
        RECT 374.200 -560.440 374.480 -530.000 ;
        RECT 378.560 -560.440 378.840 -530.000 ;
        RECT 449.200 -560.440 449.480 -530.000 ;
        RECT 453.560 -560.440 453.840 -530.000 ;
        RECT 524.200 -560.440 524.480 -530.000 ;
        RECT 528.560 -560.440 528.840 -530.000 ;
        RECT -525.800 -595.440 -525.520 -565.000 ;
        RECT -521.440 -595.440 -521.160 -565.000 ;
        RECT -450.800 -595.440 -450.520 -565.000 ;
        RECT -446.440 -595.440 -446.160 -565.000 ;
        RECT -375.800 -595.440 -375.520 -565.000 ;
        RECT -371.440 -595.440 -371.160 -565.000 ;
        RECT -300.800 -595.440 -300.520 -565.000 ;
        RECT -296.440 -595.440 -296.160 -565.000 ;
        RECT -225.800 -595.440 -225.520 -565.000 ;
        RECT -221.440 -595.440 -221.160 -565.000 ;
        RECT -150.800 -595.440 -150.520 -565.000 ;
        RECT -146.440 -595.440 -146.160 -565.000 ;
        RECT -75.800 -595.440 -75.520 -565.000 ;
        RECT -71.440 -595.440 -71.160 -565.000 ;
        RECT -0.800 -595.440 -0.520 -565.000 ;
        RECT 3.560 -595.440 3.840 -565.000 ;
        RECT 74.200 -595.440 74.480 -565.000 ;
        RECT 78.560 -595.440 78.840 -565.000 ;
        RECT 149.200 -595.440 149.480 -565.000 ;
        RECT 153.560 -595.440 153.840 -565.000 ;
        RECT 224.200 -595.440 224.480 -565.000 ;
        RECT 228.560 -595.440 228.840 -565.000 ;
        RECT 299.200 -595.440 299.480 -565.000 ;
        RECT 303.560 -595.440 303.840 -565.000 ;
        RECT 374.200 -595.440 374.480 -565.000 ;
        RECT 378.560 -595.440 378.840 -565.000 ;
        RECT 449.200 -595.440 449.480 -565.000 ;
        RECT 453.560 -595.440 453.840 -565.000 ;
        RECT 524.200 -595.440 524.480 -565.000 ;
        RECT 528.560 -595.440 528.840 -565.000 ;
        RECT -525.800 -630.440 -525.520 -600.000 ;
        RECT -521.440 -630.440 -521.160 -600.000 ;
        RECT -450.800 -630.440 -450.520 -600.000 ;
        RECT -446.440 -630.440 -446.160 -600.000 ;
        RECT -375.800 -630.440 -375.520 -600.000 ;
        RECT -371.440 -630.440 -371.160 -600.000 ;
        RECT -300.800 -630.440 -300.520 -600.000 ;
        RECT -296.440 -630.440 -296.160 -600.000 ;
        RECT -225.800 -630.440 -225.520 -600.000 ;
        RECT -221.440 -630.440 -221.160 -600.000 ;
        RECT -150.800 -630.440 -150.520 -600.000 ;
        RECT -146.440 -630.440 -146.160 -600.000 ;
        RECT -75.800 -630.440 -75.520 -600.000 ;
        RECT -71.440 -630.440 -71.160 -600.000 ;
        RECT -0.800 -630.440 -0.520 -600.000 ;
        RECT 3.560 -630.440 3.840 -600.000 ;
        RECT 74.200 -630.440 74.480 -600.000 ;
        RECT 78.560 -630.440 78.840 -600.000 ;
        RECT 149.200 -630.440 149.480 -600.000 ;
        RECT 153.560 -630.440 153.840 -600.000 ;
        RECT 224.200 -630.440 224.480 -600.000 ;
        RECT 228.560 -630.440 228.840 -600.000 ;
        RECT 299.200 -630.440 299.480 -600.000 ;
        RECT 303.560 -630.440 303.840 -600.000 ;
        RECT 374.200 -630.440 374.480 -600.000 ;
        RECT 378.560 -630.440 378.840 -600.000 ;
        RECT 449.200 -630.440 449.480 -600.000 ;
        RECT 453.560 -630.440 453.840 -600.000 ;
        RECT 524.200 -630.440 524.480 -600.000 ;
        RECT 528.560 -630.440 528.840 -600.000 ;
        RECT -525.800 -665.440 -525.520 -635.000 ;
        RECT -521.440 -665.440 -521.160 -635.000 ;
        RECT -450.800 -665.440 -450.520 -635.000 ;
        RECT -446.440 -665.440 -446.160 -635.000 ;
        RECT -375.800 -665.440 -375.520 -635.000 ;
        RECT -371.440 -665.440 -371.160 -635.000 ;
        RECT -300.800 -665.440 -300.520 -635.000 ;
        RECT -296.440 -665.440 -296.160 -635.000 ;
        RECT -225.800 -665.440 -225.520 -635.000 ;
        RECT -221.440 -665.440 -221.160 -635.000 ;
        RECT -150.800 -665.440 -150.520 -635.000 ;
        RECT -146.440 -665.440 -146.160 -635.000 ;
        RECT -75.800 -665.440 -75.520 -635.000 ;
        RECT -71.440 -665.440 -71.160 -635.000 ;
        RECT -0.800 -665.440 -0.520 -635.000 ;
        RECT 3.560 -665.440 3.840 -635.000 ;
        RECT 74.200 -665.440 74.480 -635.000 ;
        RECT 78.560 -665.440 78.840 -635.000 ;
        RECT 149.200 -665.440 149.480 -635.000 ;
        RECT 153.560 -665.440 153.840 -635.000 ;
        RECT 224.200 -665.440 224.480 -635.000 ;
        RECT 228.560 -665.440 228.840 -635.000 ;
        RECT 299.200 -665.440 299.480 -635.000 ;
        RECT 303.560 -665.440 303.840 -635.000 ;
        RECT 374.200 -665.440 374.480 -635.000 ;
        RECT 378.560 -665.440 378.840 -635.000 ;
        RECT 449.200 -665.440 449.480 -635.000 ;
        RECT 453.560 -665.440 453.840 -635.000 ;
        RECT 524.200 -665.440 524.480 -635.000 ;
        RECT 528.560 -665.440 528.840 -635.000 ;
        RECT -525.800 -700.440 -525.520 -670.000 ;
        RECT -521.440 -700.440 -521.160 -670.000 ;
        RECT -450.800 -700.440 -450.520 -670.000 ;
        RECT -446.440 -700.440 -446.160 -670.000 ;
        RECT -375.800 -700.440 -375.520 -670.000 ;
        RECT -371.440 -700.440 -371.160 -670.000 ;
        RECT -300.800 -700.440 -300.520 -670.000 ;
        RECT -296.440 -700.440 -296.160 -670.000 ;
        RECT -225.800 -700.440 -225.520 -670.000 ;
        RECT -221.440 -700.440 -221.160 -670.000 ;
        RECT -150.800 -700.440 -150.520 -670.000 ;
        RECT -146.440 -700.440 -146.160 -670.000 ;
        RECT -75.800 -700.440 -75.520 -670.000 ;
        RECT -71.440 -700.440 -71.160 -670.000 ;
        RECT -0.800 -700.440 -0.520 -670.000 ;
        RECT 3.560 -700.440 3.840 -670.000 ;
        RECT 74.200 -700.440 74.480 -670.000 ;
        RECT 78.560 -700.440 78.840 -670.000 ;
        RECT 149.200 -700.440 149.480 -670.000 ;
        RECT 153.560 -700.440 153.840 -670.000 ;
        RECT 224.200 -700.440 224.480 -670.000 ;
        RECT 228.560 -700.440 228.840 -670.000 ;
        RECT 299.200 -700.440 299.480 -670.000 ;
        RECT 303.560 -700.440 303.840 -670.000 ;
        RECT 374.200 -700.440 374.480 -670.000 ;
        RECT 378.560 -700.440 378.840 -670.000 ;
        RECT 449.200 -700.440 449.480 -670.000 ;
        RECT 453.560 -700.440 453.840 -670.000 ;
        RECT 524.200 -700.440 524.480 -670.000 ;
        RECT 528.560 -700.440 528.840 -670.000 ;
        RECT -525.800 -735.440 -525.520 -705.000 ;
        RECT -521.440 -735.440 -521.160 -705.000 ;
        RECT -450.800 -735.440 -450.520 -705.000 ;
        RECT -446.440 -735.440 -446.160 -705.000 ;
        RECT -375.800 -735.440 -375.520 -705.000 ;
        RECT -371.440 -735.440 -371.160 -705.000 ;
        RECT -300.800 -735.440 -300.520 -705.000 ;
        RECT -296.440 -735.440 -296.160 -705.000 ;
        RECT -225.800 -735.440 -225.520 -705.000 ;
        RECT -221.440 -735.440 -221.160 -705.000 ;
        RECT -150.800 -735.440 -150.520 -705.000 ;
        RECT -146.440 -735.440 -146.160 -705.000 ;
        RECT -75.800 -735.440 -75.520 -705.000 ;
        RECT -71.440 -735.440 -71.160 -705.000 ;
        RECT -0.800 -735.440 -0.520 -705.000 ;
        RECT 3.560 -735.440 3.840 -705.000 ;
        RECT 74.200 -735.440 74.480 -705.000 ;
        RECT 78.560 -735.440 78.840 -705.000 ;
        RECT 149.200 -735.440 149.480 -705.000 ;
        RECT 153.560 -735.440 153.840 -705.000 ;
        RECT 224.200 -735.440 224.480 -705.000 ;
        RECT 228.560 -735.440 228.840 -705.000 ;
        RECT 299.200 -735.440 299.480 -705.000 ;
        RECT 303.560 -735.440 303.840 -705.000 ;
        RECT 374.200 -735.440 374.480 -705.000 ;
        RECT 378.560 -735.440 378.840 -705.000 ;
        RECT 449.200 -735.440 449.480 -705.000 ;
        RECT 453.560 -735.440 453.840 -705.000 ;
        RECT 524.200 -735.440 524.480 -705.000 ;
        RECT 528.560 -735.440 528.840 -705.000 ;
        RECT -525.800 -770.440 -525.520 -740.000 ;
        RECT -521.440 -770.440 -521.160 -740.000 ;
        RECT -450.800 -770.440 -450.520 -740.000 ;
        RECT -446.440 -770.440 -446.160 -740.000 ;
        RECT -375.800 -770.440 -375.520 -740.000 ;
        RECT -371.440 -770.440 -371.160 -740.000 ;
        RECT -300.800 -770.440 -300.520 -740.000 ;
        RECT -296.440 -770.440 -296.160 -740.000 ;
        RECT -225.800 -770.440 -225.520 -740.000 ;
        RECT -221.440 -770.440 -221.160 -740.000 ;
        RECT -150.800 -770.440 -150.520 -740.000 ;
        RECT -146.440 -770.440 -146.160 -740.000 ;
        RECT -75.800 -770.440 -75.520 -740.000 ;
        RECT -71.440 -770.440 -71.160 -740.000 ;
        RECT -0.800 -770.440 -0.520 -740.000 ;
        RECT 3.560 -770.440 3.840 -740.000 ;
        RECT 74.200 -770.440 74.480 -740.000 ;
        RECT 78.560 -770.440 78.840 -740.000 ;
        RECT 149.200 -770.440 149.480 -740.000 ;
        RECT 153.560 -770.440 153.840 -740.000 ;
        RECT 224.200 -770.440 224.480 -740.000 ;
        RECT 228.560 -770.440 228.840 -740.000 ;
        RECT 299.200 -770.440 299.480 -740.000 ;
        RECT 303.560 -770.440 303.840 -740.000 ;
        RECT 374.200 -770.440 374.480 -740.000 ;
        RECT 378.560 -770.440 378.840 -740.000 ;
        RECT 449.200 -770.440 449.480 -740.000 ;
        RECT 453.560 -770.440 453.840 -740.000 ;
        RECT 524.200 -770.440 524.480 -740.000 ;
        RECT 528.560 -770.440 528.840 -740.000 ;
        RECT -525.800 -805.440 -525.520 -775.000 ;
        RECT -521.440 -805.440 -521.160 -775.000 ;
        RECT -450.800 -805.440 -450.520 -775.000 ;
        RECT -446.440 -805.440 -446.160 -775.000 ;
        RECT -375.800 -805.440 -375.520 -775.000 ;
        RECT -371.440 -805.440 -371.160 -775.000 ;
        RECT -300.800 -805.440 -300.520 -775.000 ;
        RECT -296.440 -805.440 -296.160 -775.000 ;
        RECT -225.800 -805.440 -225.520 -775.000 ;
        RECT -221.440 -805.440 -221.160 -775.000 ;
        RECT -150.800 -805.440 -150.520 -775.000 ;
        RECT -146.440 -805.440 -146.160 -775.000 ;
        RECT -75.800 -805.440 -75.520 -775.000 ;
        RECT -71.440 -805.440 -71.160 -775.000 ;
        RECT -0.800 -805.440 -0.520 -775.000 ;
        RECT 3.560 -805.440 3.840 -775.000 ;
        RECT 74.200 -805.440 74.480 -775.000 ;
        RECT 78.560 -805.440 78.840 -775.000 ;
        RECT 149.200 -805.440 149.480 -775.000 ;
        RECT 153.560 -805.440 153.840 -775.000 ;
        RECT 224.200 -805.440 224.480 -775.000 ;
        RECT 228.560 -805.440 228.840 -775.000 ;
        RECT 299.200 -805.440 299.480 -775.000 ;
        RECT 303.560 -805.440 303.840 -775.000 ;
        RECT 374.200 -805.440 374.480 -775.000 ;
        RECT 378.560 -805.440 378.840 -775.000 ;
        RECT 449.200 -805.440 449.480 -775.000 ;
        RECT 453.560 -805.440 453.840 -775.000 ;
        RECT 524.200 -805.440 524.480 -775.000 ;
        RECT 528.560 -805.440 528.840 -775.000 ;
        RECT -525.800 -840.440 -525.520 -810.000 ;
        RECT -521.440 -840.440 -521.160 -810.000 ;
        RECT -450.800 -840.440 -450.520 -810.000 ;
        RECT -446.440 -840.440 -446.160 -810.000 ;
        RECT -375.800 -840.440 -375.520 -810.000 ;
        RECT -371.440 -840.440 -371.160 -810.000 ;
        RECT -300.800 -840.440 -300.520 -810.000 ;
        RECT -296.440 -840.440 -296.160 -810.000 ;
        RECT -225.800 -840.440 -225.520 -810.000 ;
        RECT -221.440 -840.440 -221.160 -810.000 ;
        RECT -150.800 -840.440 -150.520 -810.000 ;
        RECT -146.440 -840.440 -146.160 -810.000 ;
        RECT -75.800 -840.440 -75.520 -810.000 ;
        RECT -71.440 -840.440 -71.160 -810.000 ;
        RECT -0.800 -840.440 -0.520 -810.000 ;
        RECT 3.560 -840.440 3.840 -810.000 ;
        RECT 74.200 -840.440 74.480 -810.000 ;
        RECT 78.560 -840.440 78.840 -810.000 ;
        RECT 149.200 -840.440 149.480 -810.000 ;
        RECT 153.560 -840.440 153.840 -810.000 ;
        RECT 224.200 -840.440 224.480 -810.000 ;
        RECT 228.560 -840.440 228.840 -810.000 ;
        RECT 299.200 -840.440 299.480 -810.000 ;
        RECT 303.560 -840.440 303.840 -810.000 ;
        RECT 374.200 -840.440 374.480 -810.000 ;
        RECT 378.560 -840.440 378.840 -810.000 ;
        RECT 449.200 -840.440 449.480 -810.000 ;
        RECT 453.560 -840.440 453.840 -810.000 ;
        RECT 524.200 -840.440 524.480 -810.000 ;
        RECT 528.560 -840.440 528.840 -810.000 ;
        RECT -525.800 -875.440 -525.520 -845.000 ;
        RECT -521.440 -875.440 -521.160 -845.000 ;
        RECT -450.800 -875.440 -450.520 -845.000 ;
        RECT -446.440 -875.440 -446.160 -845.000 ;
        RECT -375.800 -875.440 -375.520 -845.000 ;
        RECT -371.440 -875.440 -371.160 -845.000 ;
        RECT -300.800 -875.440 -300.520 -845.000 ;
        RECT -296.440 -875.440 -296.160 -845.000 ;
        RECT -225.800 -875.440 -225.520 -845.000 ;
        RECT -221.440 -875.440 -221.160 -845.000 ;
        RECT -150.800 -875.440 -150.520 -845.000 ;
        RECT -146.440 -875.440 -146.160 -845.000 ;
        RECT -75.800 -875.440 -75.520 -845.000 ;
        RECT -71.440 -875.440 -71.160 -845.000 ;
        RECT -0.800 -875.440 -0.520 -845.000 ;
        RECT 3.560 -875.440 3.840 -845.000 ;
        RECT 74.200 -875.440 74.480 -845.000 ;
        RECT 78.560 -875.440 78.840 -845.000 ;
        RECT 149.200 -875.440 149.480 -845.000 ;
        RECT 153.560 -875.440 153.840 -845.000 ;
        RECT 224.200 -875.440 224.480 -845.000 ;
        RECT 228.560 -875.440 228.840 -845.000 ;
        RECT 299.200 -875.440 299.480 -845.000 ;
        RECT 303.560 -875.440 303.840 -845.000 ;
        RECT 374.200 -875.440 374.480 -845.000 ;
        RECT 378.560 -875.440 378.840 -845.000 ;
        RECT 449.200 -875.440 449.480 -845.000 ;
        RECT 453.560 -875.440 453.840 -845.000 ;
        RECT 524.200 -875.440 524.480 -845.000 ;
        RECT 528.560 -875.440 528.840 -845.000 ;
        RECT -525.800 -910.440 -525.520 -880.000 ;
        RECT -521.440 -910.440 -521.160 -880.000 ;
        RECT -450.800 -910.440 -450.520 -880.000 ;
        RECT -446.440 -910.440 -446.160 -880.000 ;
        RECT -375.800 -910.440 -375.520 -880.000 ;
        RECT -371.440 -910.440 -371.160 -880.000 ;
        RECT -300.800 -910.440 -300.520 -880.000 ;
        RECT -296.440 -910.440 -296.160 -880.000 ;
        RECT -225.800 -910.440 -225.520 -880.000 ;
        RECT -221.440 -910.440 -221.160 -880.000 ;
        RECT -150.800 -910.440 -150.520 -880.000 ;
        RECT -146.440 -910.440 -146.160 -880.000 ;
        RECT -75.800 -910.440 -75.520 -880.000 ;
        RECT -71.440 -910.440 -71.160 -880.000 ;
        RECT -0.800 -910.440 -0.520 -880.000 ;
        RECT 3.560 -910.440 3.840 -880.000 ;
        RECT 74.200 -910.440 74.480 -880.000 ;
        RECT 78.560 -910.440 78.840 -880.000 ;
        RECT 149.200 -910.440 149.480 -880.000 ;
        RECT 153.560 -910.440 153.840 -880.000 ;
        RECT 224.200 -910.440 224.480 -880.000 ;
        RECT 228.560 -910.440 228.840 -880.000 ;
        RECT 299.200 -910.440 299.480 -880.000 ;
        RECT 303.560 -910.440 303.840 -880.000 ;
        RECT 374.200 -910.440 374.480 -880.000 ;
        RECT 378.560 -910.440 378.840 -880.000 ;
        RECT 449.200 -910.440 449.480 -880.000 ;
        RECT 453.560 -910.440 453.840 -880.000 ;
        RECT 524.200 -910.440 524.480 -880.000 ;
        RECT 528.560 -910.440 528.840 -880.000 ;
        RECT -525.800 -945.440 -525.520 -915.000 ;
        RECT -521.440 -945.440 -521.160 -915.000 ;
        RECT -450.800 -945.440 -450.520 -915.000 ;
        RECT -446.440 -945.440 -446.160 -915.000 ;
        RECT -375.800 -945.440 -375.520 -915.000 ;
        RECT -371.440 -945.440 -371.160 -915.000 ;
        RECT -300.800 -945.440 -300.520 -915.000 ;
        RECT -296.440 -945.440 -296.160 -915.000 ;
        RECT -225.800 -945.440 -225.520 -915.000 ;
        RECT -221.440 -945.440 -221.160 -915.000 ;
        RECT -150.800 -945.440 -150.520 -915.000 ;
        RECT -146.440 -945.440 -146.160 -915.000 ;
        RECT -75.800 -945.440 -75.520 -915.000 ;
        RECT -71.440 -945.440 -71.160 -915.000 ;
        RECT -0.800 -945.440 -0.520 -915.000 ;
        RECT 3.560 -945.440 3.840 -915.000 ;
        RECT 74.200 -945.440 74.480 -915.000 ;
        RECT 78.560 -945.440 78.840 -915.000 ;
        RECT 149.200 -945.440 149.480 -915.000 ;
        RECT 153.560 -945.440 153.840 -915.000 ;
        RECT 224.200 -945.440 224.480 -915.000 ;
        RECT 228.560 -945.440 228.840 -915.000 ;
        RECT 299.200 -945.440 299.480 -915.000 ;
        RECT 303.560 -945.440 303.840 -915.000 ;
        RECT 374.200 -945.440 374.480 -915.000 ;
        RECT 378.560 -945.440 378.840 -915.000 ;
        RECT 449.200 -945.440 449.480 -915.000 ;
        RECT 453.560 -945.440 453.840 -915.000 ;
        RECT 524.200 -945.440 524.480 -915.000 ;
        RECT 528.560 -945.440 528.840 -915.000 ;
    END
  END vss
  PIN vdd
    ANTENNAGATEAREA 6.408000 ;
    ANTENNADIFFAREA 1005.486084 ;
    PORT
      LAYER Nwell ;
        RECT -490.560 94.725 -487.460 97.505 ;
        RECT 142.615 59.240 145.205 102.660 ;
        RECT 295.490 46.520 462.670 49.110 ;
        RECT 295.490 42.865 364.880 43.000 ;
        RECT 367.795 42.865 403.520 43.000 ;
        RECT 406.435 42.865 431.245 43.000 ;
        RECT 434.160 42.865 462.670 43.000 ;
        RECT 295.490 38.815 462.670 42.865 ;
        RECT 295.490 38.680 327.920 38.815 ;
        RECT 330.835 38.680 448.605 38.815 ;
        RECT 451.520 38.680 462.670 38.815 ;
        RECT 295.490 35.025 351.440 35.160 ;
        RECT 354.355 35.025 399.600 35.160 ;
        RECT 402.515 35.025 440.205 35.160 ;
        RECT 443.120 35.025 462.670 35.160 ;
        RECT 295.490 30.975 462.670 35.025 ;
        RECT 295.490 30.840 326.240 30.975 ;
        RECT 329.155 30.840 372.720 30.975 ;
        RECT 375.635 30.840 440.765 30.975 ;
        RECT 443.680 30.840 462.670 30.975 ;
        RECT 295.490 27.185 348.640 27.320 ;
        RECT 351.555 27.185 462.670 27.320 ;
        RECT 295.490 23.135 462.670 27.185 ;
        RECT 295.490 23.000 448.605 23.135 ;
        RECT 451.520 23.000 462.670 23.135 ;
        RECT 295.490 19.355 302.035 19.480 ;
        RECT 308.065 19.355 398.480 19.480 ;
        RECT 295.490 19.345 398.480 19.355 ;
        RECT 401.395 19.345 462.670 19.480 ;
        RECT 295.490 15.295 462.670 19.345 ;
        RECT 295.490 15.160 372.720 15.295 ;
        RECT 375.635 15.160 413.600 15.295 ;
        RECT 416.515 15.160 448.605 15.295 ;
        RECT 451.520 15.160 462.670 15.295 ;
        RECT 295.490 11.515 321.830 11.640 ;
        RECT 322.930 11.515 345.715 11.640 ;
        RECT 351.745 11.515 462.670 11.640 ;
        RECT 170.305 -7.890 173.405 7.890 ;
        RECT 295.490 7.455 462.670 11.515 ;
        RECT 295.490 7.320 377.760 7.455 ;
        RECT 380.675 7.320 418.080 7.455 ;
        RECT 420.995 7.320 462.670 7.455 ;
        RECT 295.490 3.665 364.880 3.800 ;
        RECT 367.795 3.665 462.670 3.800 ;
        RECT 295.490 -0.385 462.670 3.665 ;
        RECT 295.490 -0.520 337.440 -0.385 ;
        RECT 340.355 -0.520 448.605 -0.385 ;
        RECT 451.520 -0.520 462.670 -0.385 ;
        RECT 295.490 -4.165 306.175 -4.040 ;
        RECT 312.205 -4.165 424.125 -4.040 ;
        RECT 431.985 -4.165 462.670 -4.040 ;
        RECT 295.490 -8.225 462.670 -4.165 ;
        RECT 295.490 -8.360 330.160 -8.225 ;
        RECT 333.075 -8.360 451.680 -8.225 ;
        RECT 454.595 -8.360 462.670 -8.225 ;
        RECT 295.490 -12.005 378.755 -11.880 ;
        RECT 382.295 -12.005 432.365 -11.880 ;
        RECT 295.490 -12.015 432.365 -12.005 ;
        RECT 435.280 -12.015 462.670 -11.880 ;
        RECT 295.490 -16.065 462.670 -12.015 ;
        RECT 295.490 -16.200 341.360 -16.065 ;
        RECT 344.275 -16.075 462.670 -16.065 ;
        RECT 344.275 -16.200 420.765 -16.075 ;
        RECT 428.625 -16.200 462.670 -16.075 ;
        RECT 295.490 -19.855 312.800 -19.720 ;
        RECT 315.715 -19.845 397.820 -19.720 ;
        RECT 403.550 -19.845 443.280 -19.720 ;
        RECT 315.715 -19.855 443.280 -19.845 ;
        RECT 446.195 -19.855 462.670 -19.720 ;
        RECT 295.490 -23.905 462.670 -19.855 ;
        RECT 295.490 -24.040 409.120 -23.905 ;
        RECT 412.035 -24.040 462.670 -23.905 ;
        RECT 295.490 -27.695 307.760 -27.560 ;
        RECT 310.675 -27.695 462.670 -27.560 ;
        RECT 295.490 -31.745 462.670 -27.695 ;
        RECT 295.490 -31.880 337.440 -31.745 ;
        RECT 340.355 -31.880 451.680 -31.745 ;
        RECT 454.595 -31.880 462.670 -31.745 ;
        RECT 295.490 -35.535 310.000 -35.400 ;
        RECT 312.915 -35.525 438.810 -35.400 ;
        RECT 442.590 -35.525 462.670 -35.400 ;
        RECT 312.915 -35.535 462.670 -35.525 ;
        RECT 295.490 -39.585 462.670 -35.535 ;
        RECT 295.490 -39.720 338.560 -39.585 ;
        RECT 341.475 -39.720 378.880 -39.585 ;
        RECT 381.795 -39.720 409.120 -39.585 ;
        RECT 412.035 -39.720 462.670 -39.585 ;
        RECT 295.490 -43.375 325.680 -43.240 ;
        RECT 328.595 -43.375 361.245 -43.240 ;
        RECT 364.160 -43.375 388.685 -43.240 ;
        RECT 391.600 -43.375 429.840 -43.240 ;
        RECT 432.755 -43.375 462.670 -43.240 ;
        RECT 295.490 -47.560 462.670 -43.375 ;
        RECT -490.560 -97.505 -487.460 -94.725 ;
        RECT 142.615 -102.660 145.205 -59.240 ;
      LAYER Metal1 ;
        RECT 142.145 117.620 143.385 122.580 ;
        RECT 142.185 101.860 143.345 117.620 ;
        RECT 142.185 101.520 145.045 101.860 ;
        RECT 142.185 98.815 143.345 101.520 ;
        RECT 142.185 98.585 144.035 98.815 ;
        RECT -487.875 96.630 -487.645 97.140 ;
        RECT -489.445 96.565 -487.645 96.630 ;
        RECT -489.445 96.400 -487.495 96.565 ;
        RECT -487.875 95.665 -487.495 96.400 ;
        RECT 142.185 96.545 143.345 98.585 ;
        RECT 144.845 96.700 145.260 98.220 ;
        RECT 142.185 96.315 144.325 96.545 ;
        RECT -487.875 95.115 -487.645 95.665 ;
        RECT 142.185 95.455 143.345 96.315 ;
        RECT 142.185 95.225 144.035 95.455 ;
        RECT 142.185 93.185 143.345 95.225 ;
        RECT 142.185 92.955 144.325 93.185 ;
        RECT 142.185 92.095 143.345 92.955 ;
        RECT 142.185 91.865 144.035 92.095 ;
        RECT 142.185 89.825 143.345 91.865 ;
        RECT 142.185 89.595 144.325 89.825 ;
        RECT -491.830 88.695 -491.430 89.085 ;
        RECT -485.890 88.695 -485.490 89.085 ;
        RECT -491.830 88.435 -485.490 88.695 ;
        RECT -491.830 88.045 -491.430 88.435 ;
        RECT -485.890 88.045 -485.490 88.435 ;
        RECT 142.185 88.735 143.345 89.595 ;
        RECT 142.185 88.505 144.035 88.735 ;
        RECT 142.185 86.465 143.345 88.505 ;
        RECT -492.330 86.305 -492.100 86.355 ;
        RECT -492.340 85.925 -491.440 86.305 ;
        RECT 142.185 86.235 144.325 86.465 ;
        RECT -492.330 85.875 -492.100 85.925 ;
        RECT 142.185 85.375 143.345 86.235 ;
        RECT 142.185 85.145 144.035 85.375 ;
        RECT -488.460 84.700 -487.560 84.775 ;
        RECT -489.430 84.470 -487.560 84.700 ;
        RECT -488.460 84.395 -487.560 84.470 ;
        RECT 142.185 83.105 143.345 85.145 ;
        RECT 142.185 82.875 144.325 83.105 ;
        RECT 142.185 82.015 143.345 82.875 ;
        RECT 142.185 81.785 144.035 82.015 ;
        RECT 142.185 79.745 143.345 81.785 ;
        RECT 142.185 79.515 144.325 79.745 ;
        RECT 142.185 78.655 143.345 79.515 ;
        RECT 142.185 78.425 144.035 78.655 ;
        RECT 142.185 76.385 143.345 78.425 ;
        RECT 142.185 76.155 144.325 76.385 ;
        RECT 142.185 75.295 143.345 76.155 ;
        RECT 142.185 75.065 144.035 75.295 ;
        RECT 142.185 73.025 143.345 75.065 ;
        RECT 142.185 72.795 144.325 73.025 ;
        RECT 142.185 71.935 143.345 72.795 ;
        RECT 142.185 71.705 144.035 71.935 ;
        RECT 142.185 69.665 143.345 71.705 ;
        RECT 142.185 69.435 144.325 69.665 ;
        RECT 142.185 68.575 143.345 69.435 ;
        RECT 142.185 68.345 144.035 68.575 ;
        RECT 142.185 66.305 143.345 68.345 ;
        RECT 142.185 66.075 144.325 66.305 ;
        RECT 142.185 65.215 143.345 66.075 ;
        RECT 142.185 64.985 144.035 65.215 ;
        RECT 142.185 62.945 143.345 64.985 ;
        RECT 142.185 62.715 144.325 62.945 ;
        RECT 142.185 60.380 143.345 62.715 ;
        RECT 142.185 60.040 145.045 60.380 ;
        RECT 142.185 59.670 143.345 60.040 ;
        RECT 295.920 48.380 462.240 48.980 ;
        RECT 296.290 46.680 296.630 48.380 ;
        RECT 299.465 47.330 299.695 48.380 ;
        RECT 301.705 47.800 301.935 48.380 ;
        RECT 303.945 47.800 304.175 48.380 ;
        RECT 306.185 47.800 306.415 48.380 ;
        RECT 308.425 47.330 308.655 48.380 ;
        RECT 310.665 47.800 310.895 48.380 ;
        RECT 312.805 47.330 313.035 48.380 ;
        RECT 315.350 46.690 315.690 48.380 ;
        RECT 316.885 47.330 317.115 48.380 ;
        RECT 319.025 47.800 319.255 48.380 ;
        RECT 321.265 47.330 321.495 48.380 ;
        RECT 323.505 47.800 323.735 48.380 ;
        RECT 325.745 47.800 325.975 48.380 ;
        RECT 327.985 47.800 328.215 48.380 ;
        RECT 330.225 47.330 330.455 48.380 ;
        RECT 332.965 47.250 333.195 48.380 ;
        RECT 334.390 46.690 334.730 48.380 ;
        RECT 335.865 47.330 336.095 48.380 ;
        RECT 338.105 47.800 338.335 48.380 ;
        RECT 340.345 47.800 340.575 48.380 ;
        RECT 342.585 47.800 342.815 48.380 ;
        RECT 344.825 47.330 345.055 48.380 ;
        RECT 347.065 47.800 347.295 48.380 ;
        RECT 349.205 47.330 349.435 48.380 ;
        RECT 351.445 47.250 351.675 48.380 ;
        RECT 353.430 46.690 353.770 48.380 ;
        RECT 354.405 47.330 354.635 48.380 ;
        RECT 356.545 47.800 356.775 48.380 ;
        RECT 358.785 47.330 359.015 48.380 ;
        RECT 361.025 47.800 361.255 48.380 ;
        RECT 363.265 47.800 363.495 48.380 ;
        RECT 365.505 47.800 365.735 48.380 ;
        RECT 367.745 47.330 367.975 48.380 ;
        RECT 370.485 47.250 370.715 48.380 ;
        RECT 372.470 46.690 372.810 48.380 ;
        RECT 373.945 47.330 374.175 48.380 ;
        RECT 376.185 47.800 376.415 48.380 ;
        RECT 378.425 47.800 378.655 48.380 ;
        RECT 380.665 47.800 380.895 48.380 ;
        RECT 382.905 47.330 383.135 48.380 ;
        RECT 385.145 47.800 385.375 48.380 ;
        RECT 387.285 47.330 387.515 48.380 ;
        RECT 391.510 46.690 391.850 48.380 ;
        RECT 392.985 47.330 393.215 48.380 ;
        RECT 395.225 47.800 395.455 48.380 ;
        RECT 397.465 47.800 397.695 48.380 ;
        RECT 399.705 47.800 399.935 48.380 ;
        RECT 401.945 47.330 402.175 48.380 ;
        RECT 404.185 47.800 404.415 48.380 ;
        RECT 406.325 47.330 406.555 48.380 ;
        RECT 410.550 46.690 410.890 48.380 ;
        RECT 411.525 47.330 411.755 48.380 ;
        RECT 413.665 47.800 413.895 48.380 ;
        RECT 415.905 47.330 416.135 48.380 ;
        RECT 418.145 47.800 418.375 48.380 ;
        RECT 420.385 47.800 420.615 48.380 ;
        RECT 422.625 47.800 422.855 48.380 ;
        RECT 424.865 47.330 425.095 48.380 ;
        RECT 426.085 47.290 426.315 48.380 ;
        RECT 429.590 46.690 429.930 48.380 ;
        RECT 431.065 47.330 431.295 48.380 ;
        RECT 433.305 47.800 433.535 48.380 ;
        RECT 435.545 47.800 435.775 48.380 ;
        RECT 437.785 47.800 438.015 48.380 ;
        RECT 440.025 47.330 440.255 48.380 ;
        RECT 442.265 47.800 442.495 48.380 ;
        RECT 444.405 47.330 444.635 48.380 ;
        RECT 448.630 46.690 448.970 48.380 ;
        RECT 451.125 47.250 451.355 48.380 ;
        RECT 453.365 47.250 453.595 48.380 ;
        RECT 455.605 47.250 455.835 48.380 ;
        RECT 457.845 47.250 458.075 48.380 ;
        RECT 460.085 47.250 460.315 48.380 ;
        RECT 461.530 46.680 461.870 48.380 ;
        RECT 296.290 41.140 296.630 42.840 ;
        RECT 297.785 41.140 298.015 42.190 ;
        RECT 300.025 41.140 300.255 41.720 ;
        RECT 302.265 41.140 302.495 41.720 ;
        RECT 304.505 41.140 304.735 41.720 ;
        RECT 306.745 41.140 306.975 42.190 ;
        RECT 308.985 41.140 309.215 41.720 ;
        RECT 311.125 41.140 311.355 42.190 ;
        RECT 313.365 41.140 313.595 42.280 ;
        RECT 315.605 41.140 315.835 42.280 ;
        RECT 322.325 41.140 322.555 42.270 ;
        RECT 324.565 41.140 324.795 42.270 ;
        RECT 326.805 41.140 327.035 42.270 ;
        RECT 329.045 41.140 329.275 42.270 ;
        RECT 331.285 41.140 331.515 42.270 ;
        RECT 334.545 41.140 334.775 42.230 ;
        RECT 335.510 41.140 335.850 42.830 ;
        RECT 340.140 41.140 340.370 42.230 ;
        RECT 343.370 41.140 343.710 41.630 ;
        RECT 346.965 41.140 347.195 42.270 ;
        RECT 349.465 41.140 349.695 42.230 ;
        RECT 352.850 41.140 353.190 41.630 ;
        RECT 356.590 41.140 356.930 41.895 ;
        RECT 358.330 41.140 358.670 41.915 ;
        RECT 362.630 41.140 362.970 41.770 ;
        RECT 364.765 41.140 364.995 41.970 ;
        RECT 369.935 41.140 370.275 41.480 ;
        RECT 372.030 41.140 372.260 42.170 ;
        RECT 372.750 41.140 372.980 42.230 ;
        RECT 374.710 41.140 375.050 42.830 ;
        RECT 376.910 41.140 377.140 42.230 ;
        RECT 381.045 41.140 381.275 41.710 ;
        RECT 383.260 41.140 383.600 41.710 ;
        RECT 386.290 41.140 386.520 41.720 ;
        RECT 391.365 41.140 391.595 42.280 ;
        RECT 395.230 41.140 395.570 41.895 ;
        RECT 396.970 41.140 397.310 41.915 ;
        RECT 401.270 41.140 401.610 41.770 ;
        RECT 403.405 41.140 403.635 41.970 ;
        RECT 408.575 41.140 408.915 41.480 ;
        RECT 410.670 41.140 410.900 42.170 ;
        RECT 411.390 41.140 411.620 42.230 ;
        RECT 413.910 41.140 414.250 42.830 ;
        RECT 415.365 41.140 415.595 42.070 ;
        RECT 419.845 41.140 420.075 42.070 ;
        RECT 426.060 41.140 426.290 42.230 ;
        RECT 426.780 41.140 427.010 42.170 ;
        RECT 428.765 41.140 429.105 41.480 ;
        RECT 434.045 41.140 434.275 41.970 ;
        RECT 436.070 41.140 436.410 41.770 ;
        RECT 440.370 41.140 440.710 41.915 ;
        RECT 442.110 41.140 442.450 41.895 ;
        RECT 444.005 41.140 444.235 42.230 ;
        RECT 451.125 41.140 451.355 42.270 ;
        RECT 453.110 41.140 453.450 42.830 ;
        RECT 455.605 41.140 455.835 42.270 ;
        RECT 457.845 41.140 458.075 42.270 ;
        RECT 460.085 41.140 460.315 42.270 ;
        RECT 461.530 41.140 461.870 42.840 ;
        RECT 295.920 40.540 462.240 41.140 ;
        RECT 296.290 38.840 296.630 40.540 ;
        RECT 297.785 39.490 298.015 40.540 ;
        RECT 300.025 39.960 300.255 40.540 ;
        RECT 302.265 39.960 302.495 40.540 ;
        RECT 304.505 39.960 304.735 40.540 ;
        RECT 306.745 39.490 306.975 40.540 ;
        RECT 308.985 39.960 309.215 40.540 ;
        RECT 311.125 39.490 311.355 40.540 ;
        RECT 315.910 38.850 316.250 40.540 ;
        RECT 319.630 39.785 319.970 40.540 ;
        RECT 321.370 39.765 321.710 40.540 ;
        RECT 325.670 39.910 326.010 40.540 ;
        RECT 327.805 39.710 328.035 40.540 ;
        RECT 332.975 40.200 333.315 40.540 ;
        RECT 335.070 39.510 335.300 40.540 ;
        RECT 335.790 39.450 336.020 40.540 ;
        RECT 338.085 39.610 338.315 40.540 ;
        RECT 345.845 39.410 346.075 40.540 ;
        RECT 348.085 39.410 348.315 40.540 ;
        RECT 350.325 39.410 350.555 40.540 ;
        RECT 352.565 39.410 352.795 40.540 ;
        RECT 355.110 38.850 355.450 40.540 ;
        RECT 357.605 39.410 357.835 40.540 ;
        RECT 359.845 39.410 360.075 40.540 ;
        RECT 362.085 39.400 362.315 40.540 ;
        RECT 363.890 39.960 364.120 40.540 ;
        RECT 369.365 39.410 369.595 40.540 ;
        RECT 371.605 39.410 371.835 40.540 ;
        RECT 373.845 39.410 374.075 40.540 ;
        RECT 376.085 39.410 376.315 40.540 ;
        RECT 378.325 39.410 378.555 40.540 ;
        RECT 380.565 39.410 380.795 40.540 ;
        RECT 382.805 39.410 383.035 40.540 ;
        RECT 385.045 39.410 385.275 40.540 ;
        RECT 386.990 39.450 387.220 40.540 ;
        RECT 390.245 39.400 390.475 40.540 ;
        RECT 394.310 38.850 394.650 40.540 ;
        RECT 396.805 39.410 397.035 40.540 ;
        RECT 399.045 39.410 399.275 40.540 ;
        RECT 401.285 39.410 401.515 40.540 ;
        RECT 403.525 39.410 403.755 40.540 ;
        RECT 404.245 39.490 404.475 40.540 ;
        RECT 406.385 39.960 406.615 40.540 ;
        RECT 408.625 39.490 408.855 40.540 ;
        RECT 410.865 39.960 411.095 40.540 ;
        RECT 413.105 39.960 413.335 40.540 ;
        RECT 415.345 39.960 415.575 40.540 ;
        RECT 417.585 39.490 417.815 40.540 ;
        RECT 419.305 39.490 419.535 40.540 ;
        RECT 421.545 39.960 421.775 40.540 ;
        RECT 423.785 39.960 424.015 40.540 ;
        RECT 426.025 39.960 426.255 40.540 ;
        RECT 428.265 39.490 428.495 40.540 ;
        RECT 430.505 39.960 430.735 40.540 ;
        RECT 432.645 39.490 432.875 40.540 ;
        RECT 433.510 38.850 433.850 40.540 ;
        RECT 434.965 39.610 435.195 40.540 ;
        RECT 438.965 39.450 439.195 40.540 ;
        RECT 443.420 39.450 443.650 40.540 ;
        RECT 444.140 39.510 444.370 40.540 ;
        RECT 446.125 40.200 446.465 40.540 ;
        RECT 451.405 39.710 451.635 40.540 ;
        RECT 453.430 39.910 453.770 40.540 ;
        RECT 457.730 39.765 458.070 40.540 ;
        RECT 459.470 39.785 459.810 40.540 ;
        RECT 461.530 38.840 461.870 40.540 ;
        RECT 296.290 33.300 296.630 35.000 ;
        RECT 297.785 33.300 298.015 34.350 ;
        RECT 300.025 33.300 300.255 33.880 ;
        RECT 302.265 33.300 302.495 33.880 ;
        RECT 304.505 33.300 304.735 33.880 ;
        RECT 306.745 33.300 306.975 34.350 ;
        RECT 308.985 33.300 309.215 33.880 ;
        RECT 311.125 33.300 311.355 34.350 ;
        RECT 313.365 33.300 313.595 34.430 ;
        RECT 315.605 33.300 315.835 34.430 ;
        RECT 317.845 33.300 318.075 34.430 ;
        RECT 320.085 33.300 320.315 34.430 ;
        RECT 322.325 33.300 322.555 34.430 ;
        RECT 324.565 33.300 324.795 34.430 ;
        RECT 326.805 33.300 327.035 34.430 ;
        RECT 329.045 33.300 329.275 34.430 ;
        RECT 331.285 33.300 331.515 34.430 ;
        RECT 333.525 33.300 333.755 34.430 ;
        RECT 335.510 33.300 335.850 34.990 ;
        RECT 339.125 33.300 339.355 34.390 ;
        RECT 343.150 33.300 343.490 34.055 ;
        RECT 344.890 33.300 345.230 34.075 ;
        RECT 349.190 33.300 349.530 33.930 ;
        RECT 351.325 33.300 351.555 34.130 ;
        RECT 356.495 33.300 356.835 33.640 ;
        RECT 358.590 33.300 358.820 34.330 ;
        RECT 359.310 33.300 359.540 34.390 ;
        RECT 362.210 33.300 362.440 33.880 ;
        RECT 367.685 33.300 367.915 34.430 ;
        RECT 369.925 33.300 370.155 34.430 ;
        RECT 372.165 33.300 372.395 34.430 ;
        RECT 374.710 33.300 375.050 34.990 ;
        RECT 377.205 33.300 377.435 34.430 ;
        RECT 379.445 33.300 379.675 34.430 ;
        RECT 381.685 33.300 381.915 34.430 ;
        RECT 387.320 33.300 387.550 33.880 ;
        RECT 391.310 33.300 391.650 34.055 ;
        RECT 393.050 33.300 393.390 34.075 ;
        RECT 397.350 33.300 397.690 33.930 ;
        RECT 399.485 33.300 399.715 34.130 ;
        RECT 404.655 33.300 404.995 33.640 ;
        RECT 406.750 33.300 406.980 34.330 ;
        RECT 407.470 33.300 407.700 34.390 ;
        RECT 413.045 33.300 413.275 34.430 ;
        RECT 413.910 33.300 414.250 34.990 ;
        RECT 416.110 33.300 416.340 34.390 ;
        RECT 419.365 33.300 419.595 34.350 ;
        RECT 421.505 33.300 421.735 33.880 ;
        RECT 423.745 33.300 423.975 34.350 ;
        RECT 425.985 33.300 426.215 33.880 ;
        RECT 428.225 33.300 428.455 33.880 ;
        RECT 430.465 33.300 430.695 33.880 ;
        RECT 432.705 33.300 432.935 34.350 ;
        RECT 435.020 33.300 435.250 34.390 ;
        RECT 435.740 33.300 435.970 34.330 ;
        RECT 437.725 33.300 438.065 33.640 ;
        RECT 443.005 33.300 443.235 34.130 ;
        RECT 445.030 33.300 445.370 33.930 ;
        RECT 449.330 33.300 449.670 34.075 ;
        RECT 451.070 33.300 451.410 34.055 ;
        RECT 453.110 33.300 453.450 34.990 ;
        RECT 457.845 33.300 458.075 34.430 ;
        RECT 460.085 33.300 460.315 34.430 ;
        RECT 461.530 33.300 461.870 35.000 ;
        RECT 295.920 32.700 462.240 33.300 ;
        RECT 296.290 31.000 296.630 32.700 ;
        RECT 298.805 31.570 299.035 32.700 ;
        RECT 301.045 31.570 301.275 32.700 ;
        RECT 303.845 31.560 304.075 32.700 ;
        RECT 306.085 31.570 306.315 32.700 ;
        RECT 308.325 31.570 308.555 32.700 ;
        RECT 310.565 31.570 310.795 32.700 ;
        RECT 312.805 31.570 313.035 32.700 ;
        RECT 315.045 31.570 315.275 32.700 ;
        RECT 315.910 31.010 316.250 32.700 ;
        RECT 317.950 31.945 318.290 32.700 ;
        RECT 319.690 31.925 320.030 32.700 ;
        RECT 323.990 32.070 324.330 32.700 ;
        RECT 326.125 31.870 326.355 32.700 ;
        RECT 331.295 32.360 331.635 32.700 ;
        RECT 333.390 31.670 333.620 32.700 ;
        RECT 334.110 31.610 334.340 32.700 ;
        RECT 336.405 31.770 336.635 32.700 ;
        RECT 346.405 31.570 346.635 32.700 ;
        RECT 350.325 31.560 350.555 32.700 ;
        RECT 352.565 31.570 352.795 32.700 ;
        RECT 355.110 31.010 355.450 32.700 ;
        RECT 357.605 31.570 357.835 32.700 ;
        RECT 361.470 32.095 361.810 32.700 ;
        RECT 364.430 31.945 364.770 32.700 ;
        RECT 366.170 31.925 366.510 32.700 ;
        RECT 370.470 32.070 370.810 32.700 ;
        RECT 372.605 31.870 372.835 32.700 ;
        RECT 377.775 32.360 378.115 32.700 ;
        RECT 379.870 31.670 380.100 32.700 ;
        RECT 380.590 31.610 380.820 32.700 ;
        RECT 385.640 32.120 385.870 32.700 ;
        RECT 388.690 32.210 389.030 32.700 ;
        RECT 392.325 31.570 392.555 32.700 ;
        RECT 394.310 31.010 394.650 32.700 ;
        RECT 396.805 31.570 397.035 32.700 ;
        RECT 399.045 31.570 399.275 32.700 ;
        RECT 401.285 31.570 401.515 32.700 ;
        RECT 403.525 31.570 403.755 32.700 ;
        RECT 405.765 31.570 405.995 32.700 ;
        RECT 408.005 31.570 408.235 32.700 ;
        RECT 410.725 32.130 410.955 32.700 ;
        RECT 412.940 32.130 413.280 32.700 ;
        RECT 416.730 32.210 417.070 32.700 ;
        RECT 419.305 31.650 419.535 32.700 ;
        RECT 421.545 32.120 421.775 32.700 ;
        RECT 423.785 32.120 424.015 32.700 ;
        RECT 426.025 32.120 426.255 32.700 ;
        RECT 428.265 31.650 428.495 32.700 ;
        RECT 430.505 32.120 430.735 32.700 ;
        RECT 432.645 31.650 432.875 32.700 ;
        RECT 433.510 31.010 433.850 32.700 ;
        RECT 435.580 31.610 435.810 32.700 ;
        RECT 436.300 31.670 436.530 32.700 ;
        RECT 438.285 32.360 438.625 32.700 ;
        RECT 443.565 31.870 443.795 32.700 ;
        RECT 445.590 32.070 445.930 32.700 ;
        RECT 449.890 31.925 450.230 32.700 ;
        RECT 451.630 31.945 451.970 32.700 ;
        RECT 454.990 32.095 455.330 32.700 ;
        RECT 459.470 32.095 459.810 32.700 ;
        RECT 461.530 31.000 461.870 32.700 ;
        RECT 296.290 25.460 296.630 27.160 ;
        RECT 297.285 25.460 297.515 26.510 ;
        RECT 299.425 25.460 299.655 26.040 ;
        RECT 301.665 25.460 301.895 26.510 ;
        RECT 303.905 25.460 304.135 26.040 ;
        RECT 306.145 25.460 306.375 26.040 ;
        RECT 308.385 25.460 308.615 26.040 ;
        RECT 310.625 25.460 310.855 26.510 ;
        RECT 313.365 25.460 313.595 26.590 ;
        RECT 315.605 25.460 315.835 26.590 ;
        RECT 318.170 25.460 318.510 25.950 ;
        RECT 321.665 25.460 321.895 26.550 ;
        RECT 324.005 25.460 324.235 26.590 ;
        RECT 326.245 25.460 326.475 26.590 ;
        RECT 328.485 25.460 328.715 26.590 ;
        RECT 332.110 25.460 332.340 26.550 ;
        RECT 335.510 25.460 335.850 27.150 ;
        RECT 340.350 25.460 340.690 26.215 ;
        RECT 342.090 25.460 342.430 26.235 ;
        RECT 346.390 25.460 346.730 26.090 ;
        RECT 348.525 25.460 348.755 26.290 ;
        RECT 353.695 25.460 354.035 25.800 ;
        RECT 355.790 25.460 356.020 26.490 ;
        RECT 356.510 25.460 356.740 26.550 ;
        RECT 359.845 25.460 360.075 26.590 ;
        RECT 362.085 25.460 362.315 26.590 ;
        RECT 364.090 25.460 364.430 25.950 ;
        RECT 367.685 25.460 367.915 26.590 ;
        RECT 370.485 25.460 370.715 26.600 ;
        RECT 372.725 25.460 372.955 26.590 ;
        RECT 374.710 25.460 375.050 27.150 ;
        RECT 377.205 25.460 377.435 26.590 ;
        RECT 378.805 25.460 379.035 26.030 ;
        RECT 381.020 25.460 381.360 26.030 ;
        RECT 384.485 25.460 384.715 26.590 ;
        RECT 386.725 25.460 386.955 26.590 ;
        RECT 389.810 25.460 390.150 25.950 ;
        RECT 393.445 25.460 393.675 26.590 ;
        RECT 395.685 25.460 395.915 26.590 ;
        RECT 397.925 25.460 398.155 26.590 ;
        RECT 400.165 25.460 400.395 26.590 ;
        RECT 402.405 25.460 402.635 26.590 ;
        RECT 404.645 25.460 404.875 26.590 ;
        RECT 406.885 25.460 407.115 26.590 ;
        RECT 408.485 25.460 408.715 26.030 ;
        RECT 410.700 25.460 411.040 26.030 ;
        RECT 413.910 25.460 414.250 27.150 ;
        RECT 416.110 25.460 416.340 26.550 ;
        RECT 419.845 25.460 420.075 26.390 ;
        RECT 423.845 25.460 424.075 26.510 ;
        RECT 425.985 25.460 426.215 26.040 ;
        RECT 428.225 25.460 428.455 26.510 ;
        RECT 430.465 25.460 430.695 26.040 ;
        RECT 432.705 25.460 432.935 26.040 ;
        RECT 434.945 25.460 435.175 26.040 ;
        RECT 437.185 25.460 437.415 26.510 ;
        RECT 438.405 25.460 438.635 26.510 ;
        RECT 440.545 25.460 440.775 26.040 ;
        RECT 442.785 25.460 443.015 26.510 ;
        RECT 445.025 25.460 445.255 26.040 ;
        RECT 447.265 25.460 447.495 26.040 ;
        RECT 449.505 25.460 449.735 26.040 ;
        RECT 451.745 25.460 451.975 26.510 ;
        RECT 453.110 25.460 453.450 27.150 ;
        RECT 454.085 25.460 454.315 26.550 ;
        RECT 458.910 25.460 459.250 26.065 ;
        RECT 461.530 25.460 461.870 27.160 ;
        RECT 295.920 24.860 462.240 25.460 ;
        RECT 296.290 23.160 296.630 24.860 ;
        RECT 298.805 23.730 299.035 24.860 ;
        RECT 301.045 23.730 301.275 24.860 ;
        RECT 303.285 23.730 303.515 24.860 ;
        RECT 305.525 23.730 305.755 24.860 ;
        RECT 307.765 23.730 307.995 24.860 ;
        RECT 310.005 23.730 310.235 24.860 ;
        RECT 312.245 23.730 312.475 24.860 ;
        RECT 314.485 23.730 314.715 24.860 ;
        RECT 315.910 23.170 316.250 24.860 ;
        RECT 318.405 23.730 318.635 24.860 ;
        RECT 320.645 23.730 320.875 24.860 ;
        RECT 322.885 23.730 323.115 24.860 ;
        RECT 325.125 23.730 325.355 24.860 ;
        RECT 327.365 23.730 327.595 24.860 ;
        RECT 329.605 23.730 329.835 24.860 ;
        RECT 331.845 23.730 332.075 24.860 ;
        RECT 335.765 23.770 335.995 24.860 ;
        RECT 340.245 23.730 340.475 24.860 ;
        RECT 342.485 23.730 342.715 24.860 ;
        RECT 344.725 23.720 344.955 24.860 ;
        RECT 345.925 23.930 346.155 24.860 ;
        RECT 353.685 23.730 353.915 24.860 ;
        RECT 355.110 23.170 355.450 24.860 ;
        RECT 357.605 23.730 357.835 24.860 ;
        RECT 359.845 23.730 360.075 24.860 ;
        RECT 362.085 23.730 362.315 24.860 ;
        RECT 364.325 23.730 364.555 24.860 ;
        RECT 366.565 23.730 366.795 24.860 ;
        RECT 368.805 23.730 369.035 24.860 ;
        RECT 371.045 23.730 371.275 24.860 ;
        RECT 373.285 23.730 373.515 24.860 ;
        RECT 375.525 23.730 375.755 24.860 ;
        RECT 377.765 23.730 377.995 24.860 ;
        RECT 380.005 23.730 380.235 24.860 ;
        RECT 382.245 23.730 382.475 24.860 ;
        RECT 385.730 24.280 385.960 24.860 ;
        RECT 389.685 23.720 389.915 24.860 ;
        RECT 393.445 23.730 393.675 24.860 ;
        RECT 394.310 23.170 394.650 24.860 ;
        RECT 396.805 23.730 397.035 24.860 ;
        RECT 399.045 23.730 399.275 24.860 ;
        RECT 401.285 23.730 401.515 24.860 ;
        RECT 403.525 23.730 403.755 24.860 ;
        RECT 405.765 23.730 405.995 24.860 ;
        RECT 408.005 23.730 408.235 24.860 ;
        RECT 410.245 23.730 410.475 24.860 ;
        RECT 412.485 23.730 412.715 24.860 ;
        RECT 414.725 23.730 414.955 24.860 ;
        RECT 416.965 23.730 417.195 24.860 ;
        RECT 419.490 24.370 419.830 24.860 ;
        RECT 422.890 24.370 423.230 24.860 ;
        RECT 426.405 24.290 426.635 24.860 ;
        RECT 428.620 24.290 428.960 24.860 ;
        RECT 433.510 23.170 433.850 24.860 ;
        RECT 435.770 24.370 436.110 24.860 ;
        RECT 438.405 23.770 438.635 24.860 ;
        RECT 443.420 23.770 443.650 24.860 ;
        RECT 444.140 23.830 444.370 24.860 ;
        RECT 446.125 24.520 446.465 24.860 ;
        RECT 451.405 24.030 451.635 24.860 ;
        RECT 453.430 24.230 453.770 24.860 ;
        RECT 457.730 24.085 458.070 24.860 ;
        RECT 459.470 24.105 459.810 24.860 ;
        RECT 461.530 23.160 461.870 24.860 ;
        RECT 296.290 17.620 296.630 19.320 ;
        RECT 298.520 17.620 298.750 18.710 ;
        RECT 300.260 17.620 300.490 18.710 ;
        RECT 302.565 17.620 302.905 18.235 ;
        RECT 306.585 17.620 306.925 18.235 ;
        RECT 309.185 17.620 309.525 17.795 ;
        RECT 313.620 17.620 313.960 18.395 ;
        RECT 315.550 17.620 315.890 18.310 ;
        RECT 318.965 17.620 319.195 18.750 ;
        RECT 321.205 17.620 321.435 18.750 ;
        RECT 326.325 17.620 326.555 18.550 ;
        RECT 329.045 17.620 329.275 18.750 ;
        RECT 331.285 17.620 331.515 18.750 ;
        RECT 333.525 17.620 333.755 18.750 ;
        RECT 335.510 17.620 335.850 19.310 ;
        RECT 338.005 17.620 338.235 18.750 ;
        RECT 340.245 17.620 340.475 18.750 ;
        RECT 342.485 17.620 342.715 18.750 ;
        RECT 344.725 17.620 344.955 18.750 ;
        RECT 346.965 17.620 347.195 18.750 ;
        RECT 349.205 17.620 349.435 18.750 ;
        RECT 351.445 17.620 351.675 18.750 ;
        RECT 353.685 17.620 353.915 18.750 ;
        RECT 355.925 17.620 356.155 18.750 ;
        RECT 358.165 17.620 358.395 18.750 ;
        RECT 360.405 17.620 360.635 18.750 ;
        RECT 362.645 17.620 362.875 18.750 ;
        RECT 366.330 17.620 366.670 18.110 ;
        RECT 369.925 17.620 370.155 18.760 ;
        RECT 372.165 17.620 372.395 18.750 ;
        RECT 374.710 17.620 375.050 19.310 ;
        RECT 377.205 17.620 377.435 18.750 ;
        RECT 379.445 17.620 379.675 18.750 ;
        RECT 384.520 17.620 384.750 18.200 ;
        RECT 387.845 17.620 388.075 18.750 ;
        RECT 390.190 17.620 390.530 18.375 ;
        RECT 391.930 17.620 392.270 18.395 ;
        RECT 396.230 17.620 396.570 18.250 ;
        RECT 398.365 17.620 398.595 18.450 ;
        RECT 403.535 17.620 403.875 17.960 ;
        RECT 405.630 17.620 405.860 18.650 ;
        RECT 406.350 17.620 406.580 18.710 ;
        RECT 409.685 17.620 409.915 18.750 ;
        RECT 411.925 17.620 412.155 18.750 ;
        RECT 413.910 17.620 414.250 19.310 ;
        RECT 417.525 17.620 417.755 18.710 ;
        RECT 419.765 17.620 419.995 18.750 ;
        RECT 422.005 17.620 422.235 18.750 ;
        RECT 424.245 17.620 424.475 18.750 ;
        RECT 425.525 17.620 425.755 18.710 ;
        RECT 430.670 17.620 430.900 18.710 ;
        RECT 437.205 17.620 437.435 18.550 ;
        RECT 438.405 17.620 438.635 18.670 ;
        RECT 440.545 17.620 440.775 18.200 ;
        RECT 442.785 17.620 443.015 18.670 ;
        RECT 445.025 17.620 445.255 18.200 ;
        RECT 447.265 17.620 447.495 18.200 ;
        RECT 449.505 17.620 449.735 18.200 ;
        RECT 451.745 17.620 451.975 18.670 ;
        RECT 453.110 17.620 453.450 19.310 ;
        RECT 455.605 17.620 455.835 18.750 ;
        RECT 457.205 17.620 457.435 18.190 ;
        RECT 459.420 17.620 459.760 18.190 ;
        RECT 461.530 17.620 461.870 19.320 ;
        RECT 295.920 17.020 462.240 17.620 ;
        RECT 296.290 15.320 296.630 17.020 ;
        RECT 297.785 15.970 298.015 17.020 ;
        RECT 300.025 16.440 300.255 17.020 ;
        RECT 302.265 16.440 302.495 17.020 ;
        RECT 304.505 16.440 304.735 17.020 ;
        RECT 306.745 15.970 306.975 17.020 ;
        RECT 308.985 16.440 309.215 17.020 ;
        RECT 311.125 15.970 311.355 17.020 ;
        RECT 315.910 15.330 316.250 17.020 ;
        RECT 318.405 15.890 318.635 17.020 ;
        RECT 319.685 15.930 319.915 17.020 ;
        RECT 327.365 15.930 327.595 17.020 ;
        RECT 329.605 15.890 329.835 17.020 ;
        RECT 331.845 15.890 332.075 17.020 ;
        RECT 334.085 15.890 334.315 17.020 ;
        RECT 336.325 15.890 336.555 17.020 ;
        RECT 338.565 15.890 338.795 17.020 ;
        RECT 340.805 15.890 341.035 17.020 ;
        RECT 344.805 16.090 345.035 17.020 ;
        RECT 347.525 15.890 347.755 17.020 ;
        RECT 349.765 15.890 349.995 17.020 ;
        RECT 352.005 15.890 352.235 17.020 ;
        RECT 354.245 15.890 354.475 17.020 ;
        RECT 355.110 15.330 355.450 17.020 ;
        RECT 357.605 15.890 357.835 17.020 ;
        RECT 359.845 15.890 360.075 17.020 ;
        RECT 362.085 15.890 362.315 17.020 ;
        RECT 364.430 16.265 364.770 17.020 ;
        RECT 366.170 16.245 366.510 17.020 ;
        RECT 370.470 16.390 370.810 17.020 ;
        RECT 372.605 16.190 372.835 17.020 ;
        RECT 377.775 16.680 378.115 17.020 ;
        RECT 379.870 15.990 380.100 17.020 ;
        RECT 380.590 15.930 380.820 17.020 ;
        RECT 383.925 15.890 384.155 17.020 ;
        RECT 386.165 15.890 386.395 17.020 ;
        RECT 388.405 15.890 388.635 17.020 ;
        RECT 390.645 15.890 390.875 17.020 ;
        RECT 394.310 15.330 394.650 17.020 ;
        RECT 396.570 16.530 396.910 17.020 ;
        RECT 399.730 16.440 399.960 17.020 ;
        RECT 405.310 16.265 405.650 17.020 ;
        RECT 407.050 16.245 407.390 17.020 ;
        RECT 411.350 16.390 411.690 17.020 ;
        RECT 413.485 16.190 413.715 17.020 ;
        RECT 418.655 16.680 418.995 17.020 ;
        RECT 420.750 15.990 420.980 17.020 ;
        RECT 421.470 15.930 421.700 17.020 ;
        RECT 423.605 16.450 423.835 17.020 ;
        RECT 425.820 16.450 426.160 17.020 ;
        RECT 429.050 16.530 429.390 17.020 ;
        RECT 432.645 15.890 432.875 17.020 ;
        RECT 433.510 15.330 433.850 17.020 ;
        RECT 437.765 16.090 437.995 17.020 ;
        RECT 440.485 15.890 440.715 17.020 ;
        RECT 443.420 15.930 443.650 17.020 ;
        RECT 444.140 15.990 444.370 17.020 ;
        RECT 446.125 16.680 446.465 17.020 ;
        RECT 451.405 16.190 451.635 17.020 ;
        RECT 453.430 16.390 453.770 17.020 ;
        RECT 457.730 16.245 458.070 17.020 ;
        RECT 459.470 16.265 459.810 17.020 ;
        RECT 461.530 15.320 461.870 17.020 ;
        RECT 296.290 9.780 296.630 11.480 ;
        RECT 298.805 9.780 299.035 10.910 ;
        RECT 301.045 9.780 301.275 10.910 ;
        RECT 303.285 9.780 303.515 10.910 ;
        RECT 306.805 9.780 307.035 10.175 ;
        RECT 309.165 9.780 309.395 10.870 ;
        RECT 313.410 9.780 313.770 10.500 ;
        RECT 317.585 9.780 317.815 10.560 ;
        RECT 319.800 9.780 320.140 10.585 ;
        RECT 323.505 9.780 323.735 10.385 ;
        RECT 324.775 9.780 325.005 10.480 ;
        RECT 328.085 9.780 328.315 10.480 ;
        RECT 330.725 9.780 330.955 10.910 ;
        RECT 332.965 9.780 333.195 10.910 ;
        RECT 335.510 9.780 335.850 11.470 ;
        RECT 338.005 9.780 338.235 10.910 ;
        RECT 340.245 9.780 340.475 10.910 ;
        RECT 342.200 9.780 342.430 10.870 ;
        RECT 343.940 9.780 344.170 10.870 ;
        RECT 346.245 9.780 346.585 10.395 ;
        RECT 350.265 9.780 350.605 10.395 ;
        RECT 352.865 9.780 353.205 9.955 ;
        RECT 357.300 9.780 357.640 10.555 ;
        RECT 359.230 9.780 359.570 10.470 ;
        RECT 362.645 9.780 362.875 10.910 ;
        RECT 364.885 9.780 365.115 10.910 ;
        RECT 368.190 9.780 368.530 10.385 ;
        RECT 371.550 9.780 371.890 10.385 ;
        RECT 374.710 9.780 375.050 11.470 ;
        RECT 377.205 9.780 377.435 10.910 ;
        RECT 379.445 9.780 379.675 10.910 ;
        RECT 381.685 9.780 381.915 10.910 ;
        RECT 383.845 9.780 384.075 10.350 ;
        RECT 386.060 9.780 386.400 10.350 ;
        RECT 389.470 9.780 389.810 10.385 ;
        RECT 391.415 9.780 391.645 10.775 ;
        RECT 395.730 9.780 396.090 10.115 ;
        RECT 398.485 9.780 398.715 10.910 ;
        RECT 400.725 9.780 400.955 10.910 ;
        RECT 403.125 9.780 403.355 10.920 ;
        RECT 406.830 9.780 407.170 10.385 ;
        RECT 412.485 9.780 412.715 10.910 ;
        RECT 413.910 9.780 414.250 11.470 ;
        RECT 416.405 9.780 416.635 10.910 ;
        RECT 418.645 9.780 418.875 10.910 ;
        RECT 420.885 9.780 421.115 10.910 ;
        RECT 423.125 9.780 423.355 10.910 ;
        RECT 425.365 9.780 425.595 10.910 ;
        RECT 429.285 9.780 429.515 10.910 ;
        RECT 431.525 9.780 431.755 10.910 ;
        RECT 436.460 9.780 436.690 10.870 ;
        RECT 438.405 9.780 438.635 10.830 ;
        RECT 440.545 9.780 440.775 10.360 ;
        RECT 442.785 9.780 443.015 10.830 ;
        RECT 445.025 9.780 445.255 10.360 ;
        RECT 447.265 9.780 447.495 10.360 ;
        RECT 449.505 9.780 449.735 10.360 ;
        RECT 451.745 9.780 451.975 10.830 ;
        RECT 453.110 9.780 453.450 11.470 ;
        RECT 455.605 9.780 455.835 10.910 ;
        RECT 457.845 9.780 458.075 10.910 ;
        RECT 460.085 9.780 460.315 10.910 ;
        RECT 461.530 9.780 461.870 11.480 ;
        RECT 295.920 9.180 462.240 9.780 ;
        RECT 296.290 7.480 296.630 9.180 ;
        RECT 298.350 8.575 298.690 9.180 ;
        RECT 302.830 8.575 303.170 9.180 ;
        RECT 306.240 8.610 306.580 9.180 ;
        RECT 308.565 8.610 308.795 9.180 ;
        RECT 312.140 8.090 312.370 9.180 ;
        RECT 315.910 7.490 316.250 9.180 ;
        RECT 320.165 8.250 320.395 9.180 ;
        RECT 321.370 8.090 321.600 9.180 ;
        RECT 323.410 8.090 323.640 9.180 ;
        RECT 325.685 8.050 325.915 9.180 ;
        RECT 330.730 8.245 331.070 9.180 ;
        RECT 337.150 8.350 337.490 9.180 ;
        RECT 343.045 8.050 343.275 9.180 ;
        RECT 346.405 8.090 346.635 9.180 ;
        RECT 348.645 8.050 348.875 9.180 ;
        RECT 350.885 8.050 351.115 9.180 ;
        RECT 353.125 8.050 353.355 9.180 ;
        RECT 355.110 7.490 355.450 9.180 ;
        RECT 357.605 8.050 357.835 9.180 ;
        RECT 359.845 8.050 360.075 9.180 ;
        RECT 362.085 8.050 362.315 9.180 ;
        RECT 364.325 8.050 364.555 9.180 ;
        RECT 366.565 8.050 366.795 9.180 ;
        RECT 369.470 8.425 369.810 9.180 ;
        RECT 371.210 8.405 371.550 9.180 ;
        RECT 375.510 8.550 375.850 9.180 ;
        RECT 377.645 8.350 377.875 9.180 ;
        RECT 382.815 8.840 383.155 9.180 ;
        RECT 384.910 8.130 385.145 9.180 ;
        RECT 385.625 8.130 385.860 9.180 ;
        RECT 387.615 8.090 387.955 9.180 ;
        RECT 392.885 8.090 393.115 9.180 ;
        RECT 394.310 7.490 394.650 9.180 ;
        RECT 399.045 8.050 399.275 9.180 ;
        RECT 401.410 8.600 401.640 9.180 ;
        RECT 406.485 8.040 406.715 9.180 ;
        RECT 409.790 8.425 410.130 9.180 ;
        RECT 411.530 8.405 411.870 9.180 ;
        RECT 415.830 8.550 416.170 9.180 ;
        RECT 417.965 8.350 418.195 9.180 ;
        RECT 423.135 8.840 423.475 9.180 ;
        RECT 425.230 8.150 425.460 9.180 ;
        RECT 425.950 8.090 426.180 9.180 ;
        RECT 429.285 8.050 429.515 9.180 ;
        RECT 431.525 8.050 431.755 9.180 ;
        RECT 433.510 7.490 433.850 9.180 ;
        RECT 437.765 8.250 437.995 9.180 ;
        RECT 440.080 8.610 440.420 9.180 ;
        RECT 442.405 8.610 442.635 9.180 ;
        RECT 444.965 8.050 445.195 9.180 ;
        RECT 446.805 8.130 447.035 9.180 ;
        RECT 448.945 8.600 449.175 9.180 ;
        RECT 451.185 8.130 451.415 9.180 ;
        RECT 453.425 8.600 453.655 9.180 ;
        RECT 455.665 8.600 455.895 9.180 ;
        RECT 457.905 8.600 458.135 9.180 ;
        RECT 460.145 8.130 460.375 9.180 ;
        RECT 461.530 7.480 461.870 9.180 ;
        RECT 169.355 6.215 169.735 6.550 ;
        RECT 170.490 6.215 170.720 7.100 ;
        RECT 169.355 5.985 172.290 6.215 ;
        RECT 169.355 5.650 169.735 5.985 ;
        RECT 170.490 5.100 170.720 5.985 ;
        RECT 296.290 1.940 296.630 3.640 ;
        RECT 300.965 1.940 301.195 2.510 ;
        RECT 303.180 1.940 303.520 2.510 ;
        RECT 309.450 1.940 309.790 2.875 ;
        RECT 315.870 1.940 316.210 2.770 ;
        RECT 320.805 1.940 321.035 3.080 ;
        RECT 330.670 1.940 331.010 2.545 ;
        RECT 334.085 1.940 334.315 3.070 ;
        RECT 335.510 1.940 335.850 3.630 ;
        RECT 338.005 1.940 338.235 3.070 ;
        RECT 340.245 1.940 340.475 3.070 ;
        RECT 342.485 1.940 342.715 3.070 ;
        RECT 343.525 1.940 343.755 2.510 ;
        RECT 345.740 1.940 346.080 2.510 ;
        RECT 349.205 1.940 349.435 3.080 ;
        RECT 353.685 1.940 353.915 3.070 ;
        RECT 356.590 1.940 356.930 2.695 ;
        RECT 358.330 1.940 358.670 2.715 ;
        RECT 362.630 1.940 362.970 2.570 ;
        RECT 364.765 1.940 364.995 2.770 ;
        RECT 369.935 1.940 370.275 2.280 ;
        RECT 372.030 1.940 372.260 2.970 ;
        RECT 372.750 1.940 372.980 3.030 ;
        RECT 374.710 1.940 375.050 3.630 ;
        RECT 377.205 1.940 377.435 3.070 ;
        RECT 379.445 1.940 379.675 3.070 ;
        RECT 381.685 1.940 381.915 3.070 ;
        RECT 383.925 1.940 384.155 3.070 ;
        RECT 387.610 1.940 387.950 2.430 ;
        RECT 391.750 1.940 392.110 2.275 ;
        RECT 396.195 1.940 396.425 2.935 ;
        RECT 399.105 1.940 399.335 2.405 ;
        RECT 403.585 1.940 403.815 2.405 ;
        RECT 413.045 1.940 413.275 3.070 ;
        RECT 413.910 1.940 414.250 3.630 ;
        RECT 416.405 1.940 416.635 3.070 ;
        RECT 418.645 1.940 418.875 3.070 ;
        RECT 420.885 1.940 421.115 3.070 ;
        RECT 423.125 1.940 423.355 3.070 ;
        RECT 425.365 1.940 425.595 3.070 ;
        RECT 427.310 1.940 427.540 3.030 ;
        RECT 431.045 1.940 431.275 2.870 ;
        RECT 435.045 1.940 435.275 3.030 ;
        RECT 438.405 1.940 438.635 2.990 ;
        RECT 440.545 1.940 440.775 2.520 ;
        RECT 442.785 1.940 443.015 2.990 ;
        RECT 445.025 1.940 445.255 2.520 ;
        RECT 447.265 1.940 447.495 2.520 ;
        RECT 449.505 1.940 449.735 2.520 ;
        RECT 451.745 1.940 451.975 2.990 ;
        RECT 453.110 1.940 453.450 3.630 ;
        RECT 455.200 1.940 455.540 2.510 ;
        RECT 457.525 1.940 457.755 2.510 ;
        RECT 460.085 1.940 460.315 3.070 ;
        RECT 461.530 1.940 461.870 3.640 ;
        RECT 295.920 1.340 462.240 1.940 ;
        RECT 169.355 0.115 169.735 0.450 ;
        RECT 170.490 0.115 170.720 1.000 ;
        RECT 169.355 -0.115 172.290 0.115 ;
        RECT 169.355 -0.450 169.735 -0.115 ;
        RECT 170.490 -1.000 170.720 -0.115 ;
        RECT 296.290 -0.360 296.630 1.340 ;
        RECT 298.805 0.210 299.035 1.340 ;
        RECT 301.045 0.210 301.275 1.340 ;
        RECT 302.150 1.005 302.510 1.340 ;
        RECT 306.595 0.345 306.825 1.340 ;
        RECT 308.885 0.210 309.115 1.340 ;
        RECT 311.125 0.210 311.355 1.340 ;
        RECT 313.365 0.210 313.595 1.340 ;
        RECT 315.910 -0.350 316.250 1.340 ;
        RECT 317.845 0.640 318.075 1.340 ;
        RECT 321.155 0.640 321.385 1.340 ;
        RECT 325.685 0.210 325.915 1.340 ;
        RECT 329.150 0.585 329.490 1.340 ;
        RECT 330.890 0.565 331.230 1.340 ;
        RECT 335.190 0.710 335.530 1.340 ;
        RECT 337.325 0.510 337.555 1.340 ;
        RECT 342.495 1.000 342.835 1.340 ;
        RECT 344.590 0.310 344.820 1.340 ;
        RECT 345.310 0.250 345.540 1.340 ;
        RECT 347.125 0.310 347.355 1.340 ;
        RECT 351.505 0.680 351.735 1.340 ;
        RECT 355.110 -0.350 355.450 1.340 ;
        RECT 357.150 0.735 357.490 1.340 ;
        RECT 364.405 0.410 364.635 1.340 ;
        RECT 367.125 0.210 367.355 1.340 ;
        RECT 368.325 0.410 368.555 1.340 ;
        RECT 373.845 0.210 374.075 1.340 ;
        RECT 376.085 0.210 376.315 1.340 ;
        RECT 378.325 0.210 378.555 1.340 ;
        RECT 380.565 0.210 380.795 1.340 ;
        RECT 381.945 0.250 382.175 1.340 ;
        RECT 385.245 0.730 385.585 1.340 ;
        RECT 387.480 0.730 387.820 1.340 ;
        RECT 390.845 0.730 391.185 1.340 ;
        RECT 393.080 0.730 393.420 1.340 ;
        RECT 394.310 -0.350 394.650 1.340 ;
        RECT 395.730 0.685 396.070 1.340 ;
        RECT 397.925 0.250 398.155 1.340 ;
        RECT 398.885 0.805 399.115 1.340 ;
        RECT 400.925 0.805 401.155 1.340 ;
        RECT 402.965 0.360 403.195 1.340 ;
        RECT 407.445 0.210 407.675 1.340 ;
        RECT 408.165 0.360 408.395 1.340 ;
        RECT 410.435 0.650 410.665 1.340 ;
        RECT 412.945 0.250 413.175 1.340 ;
        RECT 416.045 0.730 416.385 1.340 ;
        RECT 418.280 0.730 418.620 1.340 ;
        RECT 420.885 0.210 421.115 1.340 ;
        RECT 423.125 0.210 423.355 1.340 ;
        RECT 425.365 0.210 425.595 1.340 ;
        RECT 427.605 0.210 427.835 1.340 ;
        RECT 429.845 0.210 430.075 1.340 ;
        RECT 432.085 0.210 432.315 1.340 ;
        RECT 433.510 -0.350 433.850 1.340 ;
        RECT 434.485 0.250 434.715 1.340 ;
        RECT 440.380 0.250 440.610 1.340 ;
        RECT 443.420 0.250 443.650 1.340 ;
        RECT 444.140 0.310 444.370 1.340 ;
        RECT 446.125 1.000 446.465 1.340 ;
        RECT 451.405 0.510 451.635 1.340 ;
        RECT 453.430 0.710 453.770 1.340 ;
        RECT 457.730 0.565 458.070 1.340 ;
        RECT 459.470 0.585 459.810 1.340 ;
        RECT 461.530 -0.360 461.870 1.340 ;
        RECT 169.355 -5.985 169.735 -5.650 ;
        RECT 170.490 -5.985 170.720 -5.100 ;
        RECT 296.290 -5.900 296.630 -4.200 ;
        RECT 298.350 -5.900 298.690 -5.210 ;
        RECT 300.280 -5.900 300.620 -5.125 ;
        RECT 304.715 -5.900 305.055 -5.725 ;
        RECT 307.315 -5.900 307.655 -5.285 ;
        RECT 311.335 -5.900 311.675 -5.285 ;
        RECT 313.750 -5.900 313.980 -4.810 ;
        RECT 315.490 -5.900 315.720 -4.810 ;
        RECT 317.480 -5.900 317.710 -4.810 ;
        RECT 319.520 -5.900 319.750 -4.810 ;
        RECT 320.295 -5.900 320.525 -5.200 ;
        RECT 323.605 -5.900 323.835 -5.200 ;
        RECT 324.760 -5.900 324.990 -4.810 ;
        RECT 326.800 -5.900 327.030 -4.810 ;
        RECT 333.525 -5.900 333.755 -4.770 ;
        RECT 335.510 -5.900 335.850 -4.210 ;
        RECT 337.950 -5.900 338.290 -5.295 ;
        RECT 341.365 -5.900 341.595 -4.770 ;
        RECT 343.605 -5.900 343.835 -4.770 ;
        RECT 345.850 -5.900 346.190 -5.565 ;
        RECT 348.385 -5.900 348.615 -4.810 ;
        RECT 352.005 -5.900 352.235 -4.760 ;
        RECT 354.245 -5.900 354.475 -4.770 ;
        RECT 356.485 -5.900 356.715 -4.770 ;
        RECT 358.725 -5.900 358.955 -4.770 ;
        RECT 361.225 -5.900 361.455 -4.810 ;
        RECT 367.125 -5.900 367.355 -4.770 ;
        RECT 371.045 -5.900 371.275 -4.810 ;
        RECT 373.285 -5.900 373.515 -4.770 ;
        RECT 374.710 -5.900 375.050 -4.210 ;
        RECT 377.205 -5.900 377.435 -4.770 ;
        RECT 379.445 -5.900 379.675 -4.770 ;
        RECT 381.845 -5.900 382.075 -4.810 ;
        RECT 387.345 -5.900 387.575 -5.435 ;
        RECT 391.825 -5.900 392.055 -5.435 ;
        RECT 400.865 -5.900 401.095 -5.280 ;
        RECT 402.850 -5.900 403.190 -5.565 ;
        RECT 404.890 -5.900 405.230 -5.565 ;
        RECT 406.930 -5.900 407.270 -5.565 ;
        RECT 409.885 -5.900 410.225 -5.290 ;
        RECT 412.120 -5.900 412.460 -5.290 ;
        RECT 413.910 -5.900 414.250 -4.210 ;
        RECT 414.985 -5.900 415.215 -4.875 ;
        RECT 416.970 -5.900 417.310 -5.565 ;
        RECT 419.010 -5.900 419.350 -5.565 ;
        RECT 421.050 -5.900 421.390 -5.565 ;
        RECT 423.190 -5.900 423.530 -5.565 ;
        RECT 427.890 -5.900 428.230 -5.565 ;
        RECT 432.545 -5.900 432.775 -4.810 ;
        RECT 436.290 -5.900 436.630 -5.410 ;
        RECT 438.405 -5.900 438.635 -4.850 ;
        RECT 440.545 -5.900 440.775 -5.320 ;
        RECT 442.785 -5.900 443.015 -4.850 ;
        RECT 445.025 -5.900 445.255 -5.320 ;
        RECT 447.265 -5.900 447.495 -5.320 ;
        RECT 449.505 -5.900 449.735 -5.320 ;
        RECT 451.745 -5.900 451.975 -4.850 ;
        RECT 453.110 -5.900 453.450 -4.210 ;
        RECT 455.605 -5.900 455.835 -4.770 ;
        RECT 458.000 -5.900 458.340 -5.330 ;
        RECT 460.325 -5.900 460.555 -5.330 ;
        RECT 461.530 -5.900 461.870 -4.200 ;
        RECT 169.355 -6.215 172.290 -5.985 ;
        RECT 169.355 -6.550 169.735 -6.215 ;
        RECT 170.490 -7.100 170.720 -6.215 ;
        RECT 295.920 -6.500 462.240 -5.900 ;
        RECT 296.290 -8.200 296.630 -6.500 ;
        RECT 297.785 -7.550 298.015 -6.500 ;
        RECT 300.025 -7.080 300.255 -6.500 ;
        RECT 302.265 -7.080 302.495 -6.500 ;
        RECT 304.505 -7.080 304.735 -6.500 ;
        RECT 306.745 -7.550 306.975 -6.500 ;
        RECT 308.985 -7.080 309.215 -6.500 ;
        RECT 311.125 -7.550 311.355 -6.500 ;
        RECT 313.365 -7.630 313.595 -6.500 ;
        RECT 315.910 -8.190 316.250 -6.500 ;
        RECT 318.405 -7.630 318.635 -6.500 ;
        RECT 321.870 -7.255 322.210 -6.500 ;
        RECT 323.610 -7.275 323.950 -6.500 ;
        RECT 327.910 -7.130 328.250 -6.500 ;
        RECT 330.045 -7.330 330.275 -6.500 ;
        RECT 335.215 -6.840 335.555 -6.500 ;
        RECT 337.310 -7.530 337.540 -6.500 ;
        RECT 338.030 -7.590 338.260 -6.500 ;
        RECT 341.365 -7.630 341.595 -6.500 ;
        RECT 343.605 -7.630 343.835 -6.500 ;
        RECT 345.845 -7.630 346.075 -6.500 ;
        RECT 348.085 -7.630 348.315 -6.500 ;
        RECT 350.325 -7.630 350.555 -6.500 ;
        RECT 352.565 -7.630 352.795 -6.500 ;
        RECT 355.110 -8.190 355.450 -6.500 ;
        RECT 357.605 -7.630 357.835 -6.500 ;
        RECT 359.845 -7.630 360.075 -6.500 ;
        RECT 363.765 -7.590 363.995 -6.500 ;
        RECT 367.085 -6.835 367.425 -6.500 ;
        RECT 372.360 -6.835 372.700 -6.500 ;
        RECT 387.130 -6.835 387.470 -6.500 ;
        RECT 394.310 -8.190 394.650 -6.500 ;
        RECT 399.170 -7.080 399.400 -6.500 ;
        RECT 405.605 -7.035 405.835 -6.500 ;
        RECT 407.645 -7.035 407.875 -6.500 ;
        RECT 409.685 -7.480 409.915 -6.500 ;
        RECT 412.640 -7.070 412.980 -6.500 ;
        RECT 414.965 -7.070 415.195 -6.500 ;
        RECT 417.525 -7.630 417.755 -6.500 ;
        RECT 419.620 -7.110 419.960 -6.500 ;
        RECT 421.855 -7.110 422.195 -6.500 ;
        RECT 424.165 -7.070 424.395 -6.500 ;
        RECT 426.380 -7.070 426.720 -6.500 ;
        RECT 429.390 -7.105 429.730 -6.500 ;
        RECT 433.510 -8.190 433.850 -6.500 ;
        RECT 436.005 -7.630 436.235 -6.500 ;
        RECT 441.045 -7.630 441.275 -6.500 ;
        RECT 443.390 -7.255 443.730 -6.500 ;
        RECT 445.130 -7.275 445.470 -6.500 ;
        RECT 449.430 -7.130 449.770 -6.500 ;
        RECT 451.565 -7.330 451.795 -6.500 ;
        RECT 456.735 -6.840 457.075 -6.500 ;
        RECT 458.830 -7.530 459.060 -6.500 ;
        RECT 459.550 -7.590 459.780 -6.500 ;
        RECT 461.530 -8.200 461.870 -6.500 ;
        RECT 296.290 -13.740 296.630 -12.040 ;
        RECT 297.785 -13.740 298.015 -12.690 ;
        RECT 300.025 -13.740 300.255 -13.160 ;
        RECT 302.265 -13.740 302.495 -13.160 ;
        RECT 304.505 -13.740 304.735 -13.160 ;
        RECT 306.745 -13.740 306.975 -12.690 ;
        RECT 308.985 -13.740 309.215 -13.160 ;
        RECT 311.125 -13.740 311.355 -12.690 ;
        RECT 313.365 -13.740 313.595 -12.610 ;
        RECT 315.605 -13.740 315.835 -12.610 ;
        RECT 317.845 -13.740 318.075 -12.610 ;
        RECT 320.085 -13.740 320.315 -12.610 ;
        RECT 322.325 -13.740 322.555 -12.610 ;
        RECT 324.565 -13.740 324.795 -12.610 ;
        RECT 326.805 -13.740 327.035 -12.610 ;
        RECT 329.045 -13.740 329.275 -12.610 ;
        RECT 331.285 -13.740 331.515 -12.610 ;
        RECT 333.525 -13.740 333.755 -12.610 ;
        RECT 335.510 -13.740 335.850 -12.050 ;
        RECT 338.005 -13.740 338.235 -12.610 ;
        RECT 340.245 -13.740 340.475 -12.610 ;
        RECT 342.485 -13.740 342.715 -12.610 ;
        RECT 344.725 -13.740 344.955 -12.610 ;
        RECT 346.615 -13.740 346.845 -12.650 ;
        RECT 348.705 -13.740 348.935 -12.650 ;
        RECT 352.910 -13.740 353.250 -13.085 ;
        RECT 356.485 -13.740 356.715 -12.610 ;
        RECT 358.725 -13.740 358.955 -12.610 ;
        RECT 360.325 -13.740 360.555 -13.170 ;
        RECT 362.540 -13.740 362.880 -13.170 ;
        RECT 365.655 -13.740 365.885 -12.650 ;
        RECT 367.745 -13.740 367.975 -12.650 ;
        RECT 371.950 -13.740 372.290 -13.085 ;
        RECT 374.710 -13.740 375.050 -12.050 ;
        RECT 377.205 -13.740 377.435 -12.610 ;
        RECT 378.025 -13.740 378.255 -12.605 ;
        RECT 382.795 -13.740 383.135 -13.325 ;
        RECT 384.935 -13.740 385.275 -13.325 ;
        RECT 387.030 -13.740 387.260 -12.715 ;
        RECT 402.605 -13.740 402.835 -13.070 ;
        RECT 407.445 -13.740 407.675 -13.070 ;
        RECT 410.405 -13.740 410.635 -12.650 ;
        RECT 413.910 -13.740 414.250 -12.050 ;
        RECT 417.725 -13.740 418.065 -13.130 ;
        RECT 419.960 -13.740 420.300 -13.130 ;
        RECT 422.565 -13.740 422.795 -12.610 ;
        RECT 424.805 -13.740 425.035 -12.610 ;
        RECT 427.180 -13.740 427.410 -12.650 ;
        RECT 427.900 -13.740 428.130 -12.710 ;
        RECT 429.885 -13.740 430.225 -13.400 ;
        RECT 435.165 -13.740 435.395 -12.910 ;
        RECT 437.190 -13.740 437.530 -13.110 ;
        RECT 441.490 -13.740 441.830 -12.965 ;
        RECT 443.230 -13.740 443.570 -12.985 ;
        RECT 448.885 -13.740 449.115 -12.610 ;
        RECT 451.125 -13.740 451.355 -12.610 ;
        RECT 453.110 -13.740 453.450 -12.050 ;
        RECT 455.605 -13.740 455.835 -12.610 ;
        RECT 457.845 -13.740 458.075 -12.610 ;
        RECT 460.085 -13.740 460.315 -12.610 ;
        RECT 461.530 -13.740 461.870 -12.040 ;
        RECT 295.920 -14.340 462.240 -13.740 ;
        RECT 296.290 -16.040 296.630 -14.340 ;
        RECT 298.805 -15.470 299.035 -14.340 ;
        RECT 300.945 -15.430 301.175 -14.340 ;
        RECT 303.050 -14.830 303.390 -14.340 ;
        RECT 305.125 -15.480 305.355 -14.340 ;
        RECT 311.125 -15.470 311.355 -14.340 ;
        RECT 313.365 -15.470 313.595 -14.340 ;
        RECT 315.910 -16.030 316.250 -14.340 ;
        RECT 318.405 -15.470 318.635 -14.340 ;
        RECT 320.645 -15.470 320.875 -14.340 ;
        RECT 322.590 -15.430 322.820 -14.340 ;
        RECT 329.930 -14.830 330.270 -14.340 ;
        RECT 333.070 -15.095 333.410 -14.340 ;
        RECT 334.810 -15.115 335.150 -14.340 ;
        RECT 339.110 -14.970 339.450 -14.340 ;
        RECT 341.245 -15.170 341.475 -14.340 ;
        RECT 346.415 -14.680 346.755 -14.340 ;
        RECT 348.510 -15.370 348.740 -14.340 ;
        RECT 349.230 -15.430 349.460 -14.340 ;
        RECT 352.330 -14.830 352.670 -14.340 ;
        RECT 355.110 -16.030 355.450 -14.340 ;
        RECT 357.605 -15.470 357.835 -14.340 ;
        RECT 360.965 -15.430 361.195 -14.340 ;
        RECT 362.070 -14.675 362.430 -14.340 ;
        RECT 366.515 -15.335 366.745 -14.340 ;
        RECT 368.805 -15.470 369.035 -14.340 ;
        RECT 370.085 -15.430 370.315 -14.340 ;
        RECT 374.965 -15.470 375.195 -14.340 ;
        RECT 376.910 -15.430 377.140 -14.340 ;
        RECT 381.450 -14.830 381.790 -14.340 ;
        RECT 385.045 -15.470 385.275 -14.340 ;
        RECT 387.285 -15.470 387.515 -14.340 ;
        RECT 390.085 -15.040 390.315 -14.340 ;
        RECT 393.395 -15.040 393.625 -14.340 ;
        RECT 394.310 -16.030 394.650 -14.340 ;
        RECT 395.605 -15.230 395.835 -14.340 ;
        RECT 397.845 -14.910 398.075 -14.340 ;
        RECT 400.265 -14.800 400.495 -14.340 ;
        RECT 402.405 -14.760 402.635 -14.340 ;
        RECT 403.145 -14.780 403.375 -14.340 ;
        RECT 405.185 -14.780 405.415 -14.340 ;
        RECT 407.225 -14.780 407.455 -14.340 ;
        RECT 409.265 -15.320 409.495 -14.340 ;
        RECT 411.625 -15.365 411.855 -14.340 ;
        RECT 413.610 -14.675 413.950 -14.340 ;
        RECT 415.650 -14.675 415.990 -14.340 ;
        RECT 417.690 -14.675 418.030 -14.340 ;
        RECT 419.830 -14.675 420.170 -14.340 ;
        RECT 424.530 -14.675 424.870 -14.340 ;
        RECT 429.185 -15.430 429.415 -14.340 ;
        RECT 431.525 -15.470 431.755 -14.340 ;
        RECT 433.510 -16.030 433.850 -14.340 ;
        RECT 436.005 -15.470 436.235 -14.340 ;
        RECT 438.245 -15.470 438.475 -14.340 ;
        RECT 440.485 -15.470 440.715 -14.340 ;
        RECT 442.725 -15.470 442.955 -14.340 ;
        RECT 444.965 -15.470 445.195 -14.340 ;
        RECT 446.805 -15.390 447.035 -14.340 ;
        RECT 448.945 -14.920 449.175 -14.340 ;
        RECT 451.185 -15.390 451.415 -14.340 ;
        RECT 453.425 -14.920 453.655 -14.340 ;
        RECT 455.665 -14.920 455.895 -14.340 ;
        RECT 457.905 -14.920 458.135 -14.340 ;
        RECT 460.145 -15.390 460.375 -14.340 ;
        RECT 461.530 -16.040 461.870 -14.340 ;
        RECT 296.290 -21.580 296.630 -19.880 ;
        RECT 297.605 -21.580 297.835 -21.010 ;
        RECT 299.820 -21.580 300.160 -21.010 ;
        RECT 304.510 -21.580 304.850 -20.825 ;
        RECT 306.250 -21.580 306.590 -20.805 ;
        RECT 310.550 -21.580 310.890 -20.950 ;
        RECT 312.685 -21.580 312.915 -20.750 ;
        RECT 317.855 -21.580 318.195 -21.240 ;
        RECT 319.950 -21.580 320.180 -20.550 ;
        RECT 320.670 -21.580 320.900 -20.490 ;
        RECT 325.765 -21.580 325.995 -20.650 ;
        RECT 330.725 -21.580 330.955 -20.450 ;
        RECT 332.965 -21.580 333.195 -20.450 ;
        RECT 335.510 -21.580 335.850 -19.890 ;
        RECT 338.005 -21.580 338.235 -20.450 ;
        RECT 340.245 -21.580 340.475 -20.450 ;
        RECT 342.485 -21.580 342.715 -20.450 ;
        RECT 344.725 -21.580 344.955 -20.450 ;
        RECT 346.965 -21.580 347.195 -20.450 ;
        RECT 349.205 -21.580 349.435 -20.450 ;
        RECT 351.445 -21.580 351.675 -20.450 ;
        RECT 353.685 -21.580 353.915 -20.450 ;
        RECT 355.925 -21.580 356.155 -20.450 ;
        RECT 358.165 -21.580 358.395 -20.450 ;
        RECT 360.405 -21.580 360.635 -20.450 ;
        RECT 362.645 -21.580 362.875 -20.450 ;
        RECT 367.530 -21.580 367.870 -21.245 ;
        RECT 374.710 -21.580 375.050 -19.890 ;
        RECT 377.105 -21.580 377.335 -20.490 ;
        RECT 379.445 -21.580 379.675 -20.450 ;
        RECT 381.845 -21.580 382.075 -20.600 ;
        RECT 383.885 -21.580 384.115 -21.045 ;
        RECT 385.925 -21.580 386.155 -21.045 ;
        RECT 388.405 -21.580 388.635 -20.450 ;
        RECT 389.510 -21.580 389.870 -21.245 ;
        RECT 393.955 -21.580 394.185 -20.585 ;
        RECT 394.775 -21.580 395.005 -20.490 ;
        RECT 396.810 -21.580 397.150 -20.980 ;
        RECT 403.970 -21.580 404.310 -20.490 ;
        RECT 406.885 -21.580 407.115 -20.450 ;
        RECT 409.385 -21.580 409.615 -20.490 ;
        RECT 413.910 -21.580 414.250 -19.890 ;
        RECT 417.065 -21.580 417.295 -20.590 ;
        RECT 423.585 -21.580 423.815 -20.550 ;
        RECT 428.165 -21.580 428.395 -20.450 ;
        RECT 431.630 -21.580 431.970 -20.975 ;
        RECT 434.990 -21.580 435.330 -20.825 ;
        RECT 436.730 -21.580 437.070 -20.805 ;
        RECT 441.030 -21.580 441.370 -20.950 ;
        RECT 443.165 -21.580 443.395 -20.750 ;
        RECT 448.335 -21.580 448.675 -21.240 ;
        RECT 450.430 -21.580 450.660 -20.550 ;
        RECT 451.150 -21.580 451.380 -20.490 ;
        RECT 453.110 -21.580 453.450 -19.890 ;
        RECT 455.890 -21.580 456.230 -21.090 ;
        RECT 459.470 -21.580 459.810 -20.975 ;
        RECT 461.530 -21.580 461.870 -19.880 ;
        RECT 295.920 -22.180 462.240 -21.580 ;
        RECT 296.290 -23.880 296.630 -22.180 ;
        RECT 297.785 -23.230 298.015 -22.180 ;
        RECT 300.025 -22.760 300.255 -22.180 ;
        RECT 302.265 -22.760 302.495 -22.180 ;
        RECT 304.505 -22.760 304.735 -22.180 ;
        RECT 306.745 -23.230 306.975 -22.180 ;
        RECT 308.985 -22.760 309.215 -22.180 ;
        RECT 311.125 -23.230 311.355 -22.180 ;
        RECT 313.090 -22.670 313.430 -22.180 ;
        RECT 315.910 -23.870 316.250 -22.180 ;
        RECT 318.405 -23.310 318.635 -22.180 ;
        RECT 321.765 -23.270 321.995 -22.180 ;
        RECT 324.005 -23.310 324.235 -22.180 ;
        RECT 326.245 -23.310 326.475 -22.180 ;
        RECT 328.485 -23.310 328.715 -22.180 ;
        RECT 330.725 -23.310 330.955 -22.180 ;
        RECT 332.965 -23.310 333.195 -22.180 ;
        RECT 335.205 -23.310 335.435 -22.180 ;
        RECT 337.445 -23.310 337.675 -22.180 ;
        RECT 339.685 -23.310 339.915 -22.180 ;
        RECT 341.925 -23.310 342.155 -22.180 ;
        RECT 344.450 -22.670 344.790 -22.180 ;
        RECT 348.085 -23.310 348.315 -22.180 ;
        RECT 350.325 -23.310 350.555 -22.180 ;
        RECT 352.725 -23.320 352.955 -22.180 ;
        RECT 355.110 -23.870 355.450 -22.180 ;
        RECT 356.085 -23.210 356.315 -22.180 ;
        RECT 360.465 -22.840 360.695 -22.180 ;
        RECT 361.720 -23.270 361.950 -22.180 ;
        RECT 363.760 -23.270 363.990 -22.180 ;
        RECT 375.940 -22.515 376.280 -22.180 ;
        RECT 381.215 -22.515 381.555 -22.180 ;
        RECT 385.045 -22.880 385.275 -22.180 ;
        RECT 388.355 -22.880 388.585 -22.180 ;
        RECT 394.310 -23.870 394.650 -22.180 ;
        RECT 396.805 -23.310 397.035 -22.180 ;
        RECT 399.045 -23.310 399.275 -22.180 ;
        RECT 400.830 -22.935 401.170 -22.180 ;
        RECT 402.570 -22.955 402.910 -22.180 ;
        RECT 406.870 -22.810 407.210 -22.180 ;
        RECT 409.005 -23.010 409.235 -22.180 ;
        RECT 414.175 -22.520 414.515 -22.180 ;
        RECT 416.270 -23.210 416.500 -22.180 ;
        RECT 416.990 -23.270 417.220 -22.180 ;
        RECT 422.085 -23.110 422.315 -22.180 ;
        RECT 427.045 -23.310 427.275 -22.180 ;
        RECT 429.285 -23.310 429.515 -22.180 ;
        RECT 431.525 -23.310 431.755 -22.180 ;
        RECT 433.510 -23.870 433.850 -22.180 ;
        RECT 434.535 -23.270 434.765 -22.180 ;
        RECT 436.625 -23.270 436.855 -22.180 ;
        RECT 440.830 -22.835 441.170 -22.180 ;
        RECT 444.910 -22.785 445.250 -22.180 ;
        RECT 446.805 -23.230 447.035 -22.180 ;
        RECT 448.945 -22.760 449.175 -22.180 ;
        RECT 451.185 -23.230 451.415 -22.180 ;
        RECT 453.425 -22.760 453.655 -22.180 ;
        RECT 455.665 -22.760 455.895 -22.180 ;
        RECT 457.905 -22.760 458.135 -22.180 ;
        RECT 460.145 -23.230 460.375 -22.180 ;
        RECT 461.530 -23.880 461.870 -22.180 ;
        RECT 296.290 -29.420 296.630 -27.720 ;
        RECT 299.470 -29.420 299.810 -28.665 ;
        RECT 301.210 -29.420 301.550 -28.645 ;
        RECT 305.510 -29.420 305.850 -28.790 ;
        RECT 307.645 -29.420 307.875 -28.590 ;
        RECT 312.815 -29.420 313.155 -29.080 ;
        RECT 314.910 -29.420 315.140 -28.390 ;
        RECT 315.630 -29.420 315.860 -28.330 ;
        RECT 317.925 -29.420 318.155 -28.490 ;
        RECT 323.150 -29.420 323.380 -28.330 ;
        RECT 327.925 -29.420 328.155 -28.290 ;
        RECT 330.165 -29.420 330.395 -28.290 ;
        RECT 332.405 -29.420 332.635 -28.290 ;
        RECT 334.645 -29.420 334.875 -28.290 ;
        RECT 335.510 -29.420 335.850 -27.730 ;
        RECT 338.005 -29.420 338.235 -28.290 ;
        RECT 340.245 -29.420 340.475 -28.290 ;
        RECT 342.485 -29.420 342.715 -28.290 ;
        RECT 344.725 -29.420 344.955 -28.290 ;
        RECT 346.965 -29.420 347.195 -28.290 ;
        RECT 348.805 -29.420 349.035 -28.280 ;
        RECT 351.605 -29.420 351.835 -28.390 ;
        RECT 355.985 -29.420 356.215 -28.760 ;
        RECT 358.725 -29.420 358.955 -28.290 ;
        RECT 360.965 -29.420 361.195 -28.290 ;
        RECT 363.205 -29.420 363.435 -28.290 ;
        RECT 365.730 -29.420 366.070 -28.930 ;
        RECT 369.365 -29.420 369.595 -28.290 ;
        RECT 371.605 -29.420 371.835 -28.290 ;
        RECT 373.845 -29.420 374.075 -28.290 ;
        RECT 374.710 -29.420 375.050 -27.730 ;
        RECT 376.930 -29.420 377.270 -28.930 ;
        RECT 380.565 -29.420 380.795 -28.290 ;
        RECT 382.805 -29.420 383.035 -28.290 ;
        RECT 383.845 -29.420 384.075 -28.850 ;
        RECT 386.060 -29.420 386.400 -28.850 ;
        RECT 389.525 -29.420 389.755 -28.290 ;
        RECT 391.765 -29.420 391.995 -28.290 ;
        RECT 394.005 -29.420 394.235 -28.290 ;
        RECT 394.730 -29.420 394.960 -28.330 ;
        RECT 396.770 -29.420 397.000 -28.330 ;
        RECT 399.045 -29.420 399.275 -28.290 ;
        RECT 403.605 -29.420 403.835 -28.490 ;
        RECT 406.325 -29.420 406.555 -28.280 ;
        RECT 408.565 -29.420 408.795 -28.290 ;
        RECT 410.805 -29.420 411.035 -28.290 ;
        RECT 413.045 -29.420 413.275 -28.290 ;
        RECT 413.910 -29.420 414.250 -27.730 ;
        RECT 416.405 -29.420 416.635 -28.290 ;
        RECT 421.740 -29.420 421.970 -28.330 ;
        RECT 423.725 -29.420 424.065 -28.930 ;
        RECT 426.810 -29.420 427.150 -28.930 ;
        RECT 431.630 -29.420 431.970 -28.815 ;
        RECT 433.925 -29.420 434.155 -29.025 ;
        RECT 436.285 -29.420 436.515 -28.330 ;
        RECT 438.405 -29.420 438.635 -28.370 ;
        RECT 440.545 -29.420 440.775 -28.840 ;
        RECT 442.785 -29.420 443.015 -28.370 ;
        RECT 445.025 -29.420 445.255 -28.840 ;
        RECT 447.265 -29.420 447.495 -28.840 ;
        RECT 449.505 -29.420 449.735 -28.840 ;
        RECT 451.745 -29.420 451.975 -28.370 ;
        RECT 453.110 -29.420 453.450 -27.730 ;
        RECT 458.000 -29.420 458.340 -28.850 ;
        RECT 460.325 -29.420 460.555 -28.850 ;
        RECT 461.530 -29.420 461.870 -27.720 ;
        RECT 295.920 -30.020 462.240 -29.420 ;
        RECT 296.290 -31.720 296.630 -30.020 ;
        RECT 297.785 -31.070 298.015 -30.020 ;
        RECT 300.025 -30.600 300.255 -30.020 ;
        RECT 302.265 -30.600 302.495 -30.020 ;
        RECT 304.505 -30.600 304.735 -30.020 ;
        RECT 306.745 -31.070 306.975 -30.020 ;
        RECT 308.985 -30.600 309.215 -30.020 ;
        RECT 311.125 -31.070 311.355 -30.020 ;
        RECT 315.910 -31.710 316.250 -30.020 ;
        RECT 319.525 -31.110 319.755 -30.020 ;
        RECT 322.885 -31.110 323.115 -30.020 ;
        RECT 325.125 -31.150 325.355 -30.020 ;
        RECT 327.365 -31.150 327.595 -30.020 ;
        RECT 329.150 -30.775 329.490 -30.020 ;
        RECT 330.890 -30.795 331.230 -30.020 ;
        RECT 335.190 -30.650 335.530 -30.020 ;
        RECT 337.325 -30.850 337.555 -30.020 ;
        RECT 342.495 -30.360 342.835 -30.020 ;
        RECT 344.590 -31.050 344.820 -30.020 ;
        RECT 345.310 -31.110 345.540 -30.020 ;
        RECT 348.645 -31.150 348.875 -30.020 ;
        RECT 350.885 -31.150 351.115 -30.020 ;
        RECT 353.125 -31.150 353.355 -30.020 ;
        RECT 355.110 -31.710 355.450 -30.020 ;
        RECT 357.605 -31.150 357.835 -30.020 ;
        RECT 359.845 -31.150 360.075 -30.020 ;
        RECT 362.085 -31.150 362.315 -30.020 ;
        RECT 364.325 -31.150 364.555 -30.020 ;
        RECT 366.565 -31.150 366.795 -30.020 ;
        RECT 368.455 -31.110 368.685 -30.020 ;
        RECT 370.545 -31.110 370.775 -30.020 ;
        RECT 374.750 -30.675 375.090 -30.020 ;
        RECT 378.325 -31.150 378.555 -30.020 ;
        RECT 380.565 -31.150 380.795 -30.020 ;
        RECT 382.805 -31.150 383.035 -30.020 ;
        RECT 384.135 -31.110 384.365 -30.020 ;
        RECT 386.225 -31.110 386.455 -30.020 ;
        RECT 390.430 -30.675 390.770 -30.020 ;
        RECT 394.310 -31.710 394.650 -30.020 ;
        RECT 396.805 -31.150 397.035 -30.020 ;
        RECT 399.045 -31.150 399.275 -30.020 ;
        RECT 401.285 -31.150 401.515 -30.020 ;
        RECT 405.285 -30.950 405.515 -30.020 ;
        RECT 408.005 -31.150 408.235 -30.020 ;
        RECT 410.245 -31.150 410.475 -30.020 ;
        RECT 412.485 -31.150 412.715 -30.020 ;
        RECT 414.725 -31.150 414.955 -30.020 ;
        RECT 416.965 -31.150 417.195 -30.020 ;
        RECT 419.205 -31.150 419.435 -30.020 ;
        RECT 424.325 -30.950 424.555 -30.020 ;
        RECT 425.925 -30.720 426.155 -30.020 ;
        RECT 429.235 -30.720 429.465 -30.020 ;
        RECT 432.645 -31.110 432.875 -30.020 ;
        RECT 433.510 -31.710 433.850 -30.020 ;
        RECT 435.605 -31.050 435.835 -30.020 ;
        RECT 441.105 -30.440 441.335 -30.020 ;
        RECT 443.390 -30.775 443.730 -30.020 ;
        RECT 445.130 -30.795 445.470 -30.020 ;
        RECT 449.430 -30.650 449.770 -30.020 ;
        RECT 451.565 -30.850 451.795 -30.020 ;
        RECT 456.735 -30.360 457.075 -30.020 ;
        RECT 458.830 -31.050 459.060 -30.020 ;
        RECT 459.550 -31.110 459.780 -30.020 ;
        RECT 461.530 -31.720 461.870 -30.020 ;
        RECT 296.290 -37.260 296.630 -35.560 ;
        RECT 298.805 -37.260 299.035 -36.130 ;
        RECT 301.710 -37.260 302.050 -36.505 ;
        RECT 303.450 -37.260 303.790 -36.485 ;
        RECT 307.750 -37.260 308.090 -36.630 ;
        RECT 309.885 -37.260 310.115 -36.430 ;
        RECT 315.055 -37.260 315.395 -36.920 ;
        RECT 317.150 -37.260 317.380 -36.230 ;
        RECT 317.870 -37.260 318.100 -36.170 ;
        RECT 320.165 -37.260 320.395 -36.330 ;
        RECT 327.925 -37.260 328.155 -36.130 ;
        RECT 331.790 -37.260 332.130 -36.655 ;
        RECT 335.510 -37.260 335.850 -35.570 ;
        RECT 339.125 -37.260 339.355 -36.170 ;
        RECT 341.365 -37.260 341.595 -36.130 ;
        RECT 343.605 -37.260 343.835 -36.130 ;
        RECT 344.645 -37.260 344.875 -36.690 ;
        RECT 346.860 -37.260 347.200 -36.690 ;
        RECT 348.805 -37.260 349.035 -36.120 ;
        RECT 351.545 -37.260 351.775 -36.600 ;
        RECT 355.925 -37.260 356.155 -36.230 ;
        RECT 357.145 -37.260 357.375 -36.600 ;
        RECT 361.525 -37.260 361.755 -36.230 ;
        RECT 363.765 -37.260 363.995 -36.120 ;
        RECT 365.950 -37.260 366.290 -36.655 ;
        RECT 368.910 -37.260 369.250 -36.655 ;
        RECT 372.670 -37.260 373.010 -36.655 ;
        RECT 374.710 -37.260 375.050 -35.570 ;
        RECT 377.205 -37.260 377.435 -36.130 ;
        RECT 382.400 -37.260 382.740 -36.690 ;
        RECT 384.725 -37.260 384.955 -36.690 ;
        RECT 388.405 -37.260 388.635 -36.170 ;
        RECT 390.590 -37.260 390.930 -36.655 ;
        RECT 394.005 -37.260 394.235 -36.130 ;
        RECT 396.245 -37.260 396.475 -36.130 ;
        RECT 398.485 -37.260 398.715 -36.130 ;
        RECT 400.725 -37.260 400.955 -36.130 ;
        RECT 402.965 -37.260 403.195 -36.130 ;
        RECT 405.205 -37.260 405.435 -36.130 ;
        RECT 407.445 -37.260 407.675 -36.130 ;
        RECT 409.685 -37.260 409.915 -36.130 ;
        RECT 411.925 -37.260 412.155 -36.130 ;
        RECT 413.910 -37.260 414.250 -35.570 ;
        RECT 416.405 -37.260 416.635 -36.130 ;
        RECT 421.445 -37.260 421.675 -36.130 ;
        RECT 423.685 -37.260 423.915 -36.130 ;
        RECT 425.925 -37.260 426.155 -36.130 ;
        RECT 428.165 -37.260 428.395 -36.130 ;
        RECT 429.445 -37.260 429.675 -36.400 ;
        RECT 431.485 -37.260 431.715 -36.625 ;
        RECT 433.625 -37.260 433.855 -36.625 ;
        RECT 435.765 -37.260 435.995 -36.625 ;
        RECT 437.905 -37.260 438.135 -36.625 ;
        RECT 440.485 -37.260 440.715 -36.625 ;
        RECT 443.165 -37.260 443.395 -36.400 ;
        RECT 445.525 -37.260 445.755 -36.120 ;
        RECT 447.530 -37.260 447.870 -36.770 ;
        RECT 450.850 -37.260 451.190 -36.770 ;
        RECT 453.110 -37.260 453.450 -35.570 ;
        RECT 457.205 -37.260 457.435 -36.690 ;
        RECT 459.420 -37.260 459.760 -36.690 ;
        RECT 461.530 -37.260 461.870 -35.560 ;
        RECT 295.920 -37.860 462.240 -37.260 ;
        RECT 296.290 -39.560 296.630 -37.860 ;
        RECT 297.785 -38.910 298.015 -37.860 ;
        RECT 300.025 -38.440 300.255 -37.860 ;
        RECT 302.265 -38.440 302.495 -37.860 ;
        RECT 304.505 -38.440 304.735 -37.860 ;
        RECT 306.745 -38.910 306.975 -37.860 ;
        RECT 308.985 -38.440 309.215 -37.860 ;
        RECT 311.125 -38.910 311.355 -37.860 ;
        RECT 313.365 -39.000 313.595 -37.860 ;
        RECT 315.910 -39.550 316.250 -37.860 ;
        RECT 318.670 -38.950 318.900 -37.860 ;
        RECT 327.310 -38.465 327.650 -37.860 ;
        RECT 330.270 -38.615 330.610 -37.860 ;
        RECT 332.010 -38.635 332.350 -37.860 ;
        RECT 336.310 -38.490 336.650 -37.860 ;
        RECT 338.445 -38.690 338.675 -37.860 ;
        RECT 343.615 -38.200 343.955 -37.860 ;
        RECT 345.710 -38.890 345.940 -37.860 ;
        RECT 346.430 -38.950 346.660 -37.860 ;
        RECT 349.765 -38.990 349.995 -37.860 ;
        RECT 352.005 -38.990 352.235 -37.860 ;
        RECT 354.245 -38.990 354.475 -37.860 ;
        RECT 355.110 -39.550 355.450 -37.860 ;
        RECT 356.085 -39.000 356.315 -37.860 ;
        RECT 359.845 -38.990 360.075 -37.860 ;
        RECT 362.085 -38.990 362.315 -37.860 ;
        RECT 364.325 -38.990 364.555 -37.860 ;
        RECT 366.565 -38.990 366.795 -37.860 ;
        RECT 368.805 -38.990 369.035 -37.860 ;
        RECT 370.590 -38.615 370.930 -37.860 ;
        RECT 372.330 -38.635 372.670 -37.860 ;
        RECT 376.630 -38.490 376.970 -37.860 ;
        RECT 378.765 -38.690 378.995 -37.860 ;
        RECT 383.935 -38.200 384.275 -37.860 ;
        RECT 386.030 -38.890 386.260 -37.860 ;
        RECT 386.750 -38.950 386.980 -37.860 ;
        RECT 390.085 -38.990 390.315 -37.860 ;
        RECT 393.445 -38.990 393.675 -37.860 ;
        RECT 394.310 -39.550 394.650 -37.860 ;
        RECT 396.805 -38.990 397.035 -37.860 ;
        RECT 399.045 -38.990 399.275 -37.860 ;
        RECT 400.830 -38.615 401.170 -37.860 ;
        RECT 402.570 -38.635 402.910 -37.860 ;
        RECT 406.870 -38.490 407.210 -37.860 ;
        RECT 409.005 -38.690 409.235 -37.860 ;
        RECT 414.175 -38.200 414.515 -37.860 ;
        RECT 416.270 -38.890 416.500 -37.860 ;
        RECT 416.990 -38.950 417.220 -37.860 ;
        RECT 419.305 -38.910 419.535 -37.860 ;
        RECT 421.545 -38.440 421.775 -37.860 ;
        RECT 423.785 -38.440 424.015 -37.860 ;
        RECT 426.025 -38.440 426.255 -37.860 ;
        RECT 428.265 -38.910 428.495 -37.860 ;
        RECT 430.505 -38.440 430.735 -37.860 ;
        RECT 432.645 -38.910 432.875 -37.860 ;
        RECT 433.510 -39.550 433.850 -37.860 ;
        RECT 435.045 -38.950 435.275 -37.860 ;
        RECT 439.925 -39.000 440.155 -37.860 ;
        RECT 442.325 -38.910 442.555 -37.860 ;
        RECT 444.465 -38.440 444.695 -37.860 ;
        RECT 446.705 -38.910 446.935 -37.860 ;
        RECT 448.945 -38.440 449.175 -37.860 ;
        RECT 451.185 -38.440 451.415 -37.860 ;
        RECT 453.425 -38.440 453.655 -37.860 ;
        RECT 455.665 -38.910 455.895 -37.860 ;
        RECT 457.140 -38.470 457.480 -37.860 ;
        RECT 459.375 -38.470 459.715 -37.860 ;
        RECT 461.530 -39.560 461.870 -37.860 ;
        RECT 296.290 -45.100 296.630 -43.400 ;
        RECT 297.785 -45.100 298.015 -44.050 ;
        RECT 300.025 -45.100 300.255 -44.520 ;
        RECT 302.265 -45.100 302.495 -44.520 ;
        RECT 304.505 -45.100 304.735 -44.520 ;
        RECT 306.745 -45.100 306.975 -44.050 ;
        RECT 308.985 -45.100 309.215 -44.520 ;
        RECT 311.125 -45.100 311.355 -44.050 ;
        RECT 312.165 -45.100 312.395 -44.530 ;
        RECT 314.380 -45.100 314.720 -44.530 ;
        RECT 317.390 -45.100 317.730 -44.345 ;
        RECT 319.130 -45.100 319.470 -44.325 ;
        RECT 323.430 -45.100 323.770 -44.470 ;
        RECT 325.565 -45.100 325.795 -44.270 ;
        RECT 330.735 -45.100 331.075 -44.760 ;
        RECT 332.830 -45.100 333.060 -44.070 ;
        RECT 333.550 -45.100 333.780 -44.010 ;
        RECT 335.510 -45.100 335.850 -43.410 ;
        RECT 337.925 -45.100 338.155 -44.530 ;
        RECT 340.140 -45.100 340.480 -44.530 ;
        RECT 345.365 -45.100 345.595 -44.170 ;
        RECT 347.790 -45.100 348.020 -44.010 ;
        RECT 352.565 -45.100 352.795 -43.970 ;
        RECT 356.060 -45.100 356.290 -44.010 ;
        RECT 356.780 -45.100 357.010 -44.070 ;
        RECT 358.765 -45.100 359.105 -44.760 ;
        RECT 364.045 -45.100 364.275 -44.270 ;
        RECT 366.070 -45.100 366.410 -44.470 ;
        RECT 370.370 -45.100 370.710 -44.325 ;
        RECT 372.110 -45.100 372.450 -44.345 ;
        RECT 374.710 -45.100 375.050 -43.410 ;
        RECT 377.205 -45.100 377.435 -43.960 ;
        RECT 380.110 -45.100 380.450 -44.495 ;
        RECT 383.500 -45.100 383.730 -44.010 ;
        RECT 384.220 -45.100 384.450 -44.070 ;
        RECT 386.205 -45.100 386.545 -44.760 ;
        RECT 391.485 -45.100 391.715 -44.270 ;
        RECT 393.510 -45.100 393.850 -44.470 ;
        RECT 397.810 -45.100 398.150 -44.325 ;
        RECT 399.550 -45.100 399.890 -44.345 ;
        RECT 405.205 -45.100 405.435 -43.970 ;
        RECT 405.925 -45.100 406.155 -43.960 ;
        RECT 411.925 -45.100 412.155 -43.970 ;
        RECT 413.910 -45.100 414.250 -43.410 ;
        RECT 416.405 -45.100 416.635 -43.970 ;
        RECT 418.245 -45.100 418.475 -43.960 ;
        RECT 421.550 -45.100 421.890 -44.345 ;
        RECT 423.290 -45.100 423.630 -44.325 ;
        RECT 427.590 -45.100 427.930 -44.470 ;
        RECT 429.725 -45.100 429.955 -44.270 ;
        RECT 434.895 -45.100 435.235 -44.760 ;
        RECT 436.990 -45.100 437.220 -44.070 ;
        RECT 437.710 -45.100 437.940 -44.010 ;
        RECT 440.645 -45.100 440.875 -43.960 ;
        RECT 446.645 -45.100 446.875 -43.970 ;
        RECT 448.885 -45.100 449.115 -43.970 ;
        RECT 453.110 -45.100 453.450 -43.410 ;
        RECT 455.505 -45.100 455.735 -44.010 ;
        RECT 459.470 -45.100 459.810 -44.495 ;
        RECT 461.530 -45.100 461.870 -43.400 ;
        RECT 295.920 -45.700 462.240 -45.100 ;
        RECT 296.290 -47.400 296.630 -45.700 ;
        RECT 299.465 -46.750 299.695 -45.700 ;
        RECT 301.705 -46.280 301.935 -45.700 ;
        RECT 303.945 -46.280 304.175 -45.700 ;
        RECT 306.185 -46.280 306.415 -45.700 ;
        RECT 308.425 -46.750 308.655 -45.700 ;
        RECT 310.665 -46.280 310.895 -45.700 ;
        RECT 312.805 -46.750 313.035 -45.700 ;
        RECT 315.350 -47.390 315.690 -45.700 ;
        RECT 316.885 -46.750 317.115 -45.700 ;
        RECT 319.025 -46.280 319.255 -45.700 ;
        RECT 321.265 -46.750 321.495 -45.700 ;
        RECT 323.505 -46.280 323.735 -45.700 ;
        RECT 325.745 -46.280 325.975 -45.700 ;
        RECT 327.985 -46.280 328.215 -45.700 ;
        RECT 330.225 -46.750 330.455 -45.700 ;
        RECT 334.390 -47.390 334.730 -45.700 ;
        RECT 335.365 -46.750 335.595 -45.700 ;
        RECT 337.505 -46.280 337.735 -45.700 ;
        RECT 339.745 -46.750 339.975 -45.700 ;
        RECT 341.985 -46.280 342.215 -45.700 ;
        RECT 344.225 -46.280 344.455 -45.700 ;
        RECT 346.465 -46.280 346.695 -45.700 ;
        RECT 348.705 -46.750 348.935 -45.700 ;
        RECT 351.445 -46.830 351.675 -45.700 ;
        RECT 353.430 -47.390 353.770 -45.700 ;
        RECT 354.405 -46.750 354.635 -45.700 ;
        RECT 356.545 -46.280 356.775 -45.700 ;
        RECT 358.785 -46.750 359.015 -45.700 ;
        RECT 361.025 -46.280 361.255 -45.700 ;
        RECT 363.265 -46.280 363.495 -45.700 ;
        RECT 365.505 -46.280 365.735 -45.700 ;
        RECT 367.745 -46.750 367.975 -45.700 ;
        RECT 370.485 -46.830 370.715 -45.700 ;
        RECT 372.470 -47.390 372.810 -45.700 ;
        RECT 373.445 -46.750 373.675 -45.700 ;
        RECT 375.585 -46.280 375.815 -45.700 ;
        RECT 377.825 -46.750 378.055 -45.700 ;
        RECT 380.065 -46.280 380.295 -45.700 ;
        RECT 382.305 -46.280 382.535 -45.700 ;
        RECT 384.545 -46.280 384.775 -45.700 ;
        RECT 386.785 -46.750 387.015 -45.700 ;
        RECT 388.565 -46.840 388.795 -45.700 ;
        RECT 391.510 -47.390 391.850 -45.700 ;
        RECT 392.485 -46.750 392.715 -45.700 ;
        RECT 394.625 -46.280 394.855 -45.700 ;
        RECT 396.865 -46.750 397.095 -45.700 ;
        RECT 399.105 -46.280 399.335 -45.700 ;
        RECT 401.345 -46.280 401.575 -45.700 ;
        RECT 403.585 -46.280 403.815 -45.700 ;
        RECT 405.825 -46.750 406.055 -45.700 ;
        RECT 408.565 -46.830 408.795 -45.700 ;
        RECT 410.550 -47.390 410.890 -45.700 ;
        RECT 411.525 -46.750 411.755 -45.700 ;
        RECT 413.665 -46.280 413.895 -45.700 ;
        RECT 415.905 -46.750 416.135 -45.700 ;
        RECT 418.145 -46.280 418.375 -45.700 ;
        RECT 420.385 -46.280 420.615 -45.700 ;
        RECT 422.625 -46.280 422.855 -45.700 ;
        RECT 424.865 -46.750 425.095 -45.700 ;
        RECT 427.605 -46.830 427.835 -45.700 ;
        RECT 429.590 -47.390 429.930 -45.700 ;
        RECT 430.565 -46.750 430.795 -45.700 ;
        RECT 432.705 -46.280 432.935 -45.700 ;
        RECT 434.945 -46.750 435.175 -45.700 ;
        RECT 437.185 -46.280 437.415 -45.700 ;
        RECT 439.425 -46.280 439.655 -45.700 ;
        RECT 441.665 -46.280 441.895 -45.700 ;
        RECT 443.905 -46.750 444.135 -45.700 ;
        RECT 446.645 -46.830 446.875 -45.700 ;
        RECT 448.630 -47.390 448.970 -45.700 ;
        RECT 455.710 -46.305 456.050 -45.700 ;
        RECT 459.470 -46.305 459.810 -45.700 ;
        RECT 461.530 -47.400 461.870 -45.700 ;
        RECT 142.185 -60.040 143.345 -59.670 ;
        RECT 142.185 -60.380 145.045 -60.040 ;
        RECT 142.185 -62.715 143.345 -60.380 ;
        RECT 142.185 -62.945 144.325 -62.715 ;
        RECT 142.185 -64.985 143.345 -62.945 ;
        RECT 142.185 -65.215 144.035 -64.985 ;
        RECT 142.185 -66.075 143.345 -65.215 ;
        RECT 142.185 -66.305 144.325 -66.075 ;
        RECT 142.185 -68.345 143.345 -66.305 ;
        RECT 142.185 -68.575 144.035 -68.345 ;
        RECT 142.185 -69.435 143.345 -68.575 ;
        RECT 142.185 -69.665 144.325 -69.435 ;
        RECT 142.185 -71.705 143.345 -69.665 ;
        RECT 142.185 -71.935 144.035 -71.705 ;
        RECT 142.185 -72.795 143.345 -71.935 ;
        RECT 142.185 -73.025 144.325 -72.795 ;
        RECT 142.185 -75.065 143.345 -73.025 ;
        RECT 142.185 -75.295 144.035 -75.065 ;
        RECT 142.185 -76.155 143.345 -75.295 ;
        RECT 142.185 -76.385 144.325 -76.155 ;
        RECT 142.185 -78.425 143.345 -76.385 ;
        RECT 142.185 -78.655 144.035 -78.425 ;
        RECT 142.185 -79.515 143.345 -78.655 ;
        RECT 142.185 -79.745 144.325 -79.515 ;
        RECT 142.185 -81.785 143.345 -79.745 ;
        RECT 142.185 -82.015 144.035 -81.785 ;
        RECT 142.185 -82.875 143.345 -82.015 ;
        RECT 142.185 -83.105 144.325 -82.875 ;
        RECT -488.460 -84.470 -487.560 -84.395 ;
        RECT -489.430 -84.700 -487.560 -84.470 ;
        RECT -488.460 -84.775 -487.560 -84.700 ;
        RECT 142.185 -85.145 143.345 -83.105 ;
        RECT 142.185 -85.375 144.035 -85.145 ;
        RECT -492.330 -85.925 -492.100 -85.875 ;
        RECT -492.340 -86.305 -491.440 -85.925 ;
        RECT 142.185 -86.235 143.345 -85.375 ;
        RECT -492.330 -86.355 -492.100 -86.305 ;
        RECT 142.185 -86.465 144.325 -86.235 ;
        RECT -491.830 -88.435 -491.430 -88.045 ;
        RECT -485.890 -88.435 -485.490 -88.045 ;
        RECT -491.830 -88.695 -485.490 -88.435 ;
        RECT -491.830 -89.085 -491.430 -88.695 ;
        RECT -485.890 -89.085 -485.490 -88.695 ;
        RECT 142.185 -88.505 143.345 -86.465 ;
        RECT 142.185 -88.735 144.035 -88.505 ;
        RECT 142.185 -89.595 143.345 -88.735 ;
        RECT 142.185 -89.825 144.325 -89.595 ;
        RECT 142.185 -91.865 143.345 -89.825 ;
        RECT 142.185 -92.095 144.035 -91.865 ;
        RECT 142.185 -92.955 143.345 -92.095 ;
        RECT 142.185 -93.185 144.325 -92.955 ;
        RECT -487.875 -95.665 -487.645 -95.115 ;
        RECT 142.185 -95.225 143.345 -93.185 ;
        RECT 142.185 -95.455 144.035 -95.225 ;
        RECT -487.875 -96.400 -487.495 -95.665 ;
        RECT -489.445 -96.565 -487.495 -96.400 ;
        RECT 142.185 -96.315 143.345 -95.455 ;
        RECT 142.185 -96.545 144.325 -96.315 ;
        RECT -489.445 -96.630 -487.645 -96.565 ;
        RECT -487.875 -97.140 -487.645 -96.630 ;
        RECT 142.185 -98.585 143.345 -96.545 ;
        RECT 144.845 -98.220 145.260 -96.700 ;
        RECT 142.185 -98.815 144.035 -98.585 ;
        RECT 142.185 -101.520 143.345 -98.815 ;
        RECT 142.185 -101.860 145.045 -101.520 ;
        RECT 142.185 -117.620 143.345 -101.860 ;
        RECT 142.145 -122.580 143.385 -117.620 ;
      LAYER Via1 ;
        RECT 142.325 122.140 142.585 122.400 ;
        RECT 142.945 122.140 143.205 122.400 ;
        RECT 142.325 121.520 142.585 121.780 ;
        RECT 142.945 121.520 143.205 121.780 ;
        RECT 142.325 120.900 142.585 121.160 ;
        RECT 142.945 120.900 143.205 121.160 ;
        RECT 142.325 120.280 142.585 120.540 ;
        RECT 142.945 120.280 143.205 120.540 ;
        RECT 142.325 119.660 142.585 119.920 ;
        RECT 142.945 119.660 143.205 119.920 ;
        RECT 142.325 119.040 142.585 119.300 ;
        RECT 142.945 119.040 143.205 119.300 ;
        RECT 142.325 118.420 142.585 118.680 ;
        RECT 142.945 118.420 143.205 118.680 ;
        RECT 142.325 117.800 142.585 118.060 ;
        RECT 142.945 117.800 143.205 118.060 ;
        RECT -487.815 95.725 -487.555 96.505 ;
        RECT 144.920 96.860 145.180 97.120 ;
        RECT -491.760 88.175 -491.500 88.955 ;
        RECT -485.820 88.175 -485.560 88.955 ;
        RECT -492.280 85.985 -491.500 86.245 ;
        RECT -488.400 84.455 -487.620 84.715 ;
        RECT 316.060 48.550 317.360 48.810 ;
        RECT 357.640 48.550 358.940 48.810 ;
        RECT 399.220 48.550 400.520 48.810 ;
        RECT 440.800 48.550 442.100 48.810 ;
        RECT 316.060 40.710 317.360 40.970 ;
        RECT 357.640 40.710 358.940 40.970 ;
        RECT 399.220 40.710 400.520 40.970 ;
        RECT 440.800 40.710 442.100 40.970 ;
        RECT 316.060 32.870 317.360 33.130 ;
        RECT 357.640 32.870 358.940 33.130 ;
        RECT 399.220 32.870 400.520 33.130 ;
        RECT 440.800 32.870 442.100 33.130 ;
        RECT 316.060 25.030 317.360 25.290 ;
        RECT 357.640 25.030 358.940 25.290 ;
        RECT 399.220 25.030 400.520 25.290 ;
        RECT 440.800 25.030 442.100 25.290 ;
        RECT 316.060 17.190 317.360 17.450 ;
        RECT 357.640 17.190 358.940 17.450 ;
        RECT 399.220 17.190 400.520 17.450 ;
        RECT 440.800 17.190 442.100 17.450 ;
        RECT 316.060 9.350 317.360 9.610 ;
        RECT 357.640 9.350 358.940 9.610 ;
        RECT 399.220 9.350 400.520 9.610 ;
        RECT 440.800 9.350 442.100 9.610 ;
        RECT 169.415 5.710 169.675 6.490 ;
        RECT 316.060 1.510 317.360 1.770 ;
        RECT 357.640 1.510 358.940 1.770 ;
        RECT 399.220 1.510 400.520 1.770 ;
        RECT 440.800 1.510 442.100 1.770 ;
        RECT 169.415 -0.390 169.675 0.390 ;
        RECT 169.415 -6.490 169.675 -5.710 ;
        RECT 316.060 -6.330 317.360 -6.070 ;
        RECT 357.640 -6.330 358.940 -6.070 ;
        RECT 399.220 -6.330 400.520 -6.070 ;
        RECT 440.800 -6.330 442.100 -6.070 ;
        RECT 316.060 -14.170 317.360 -13.910 ;
        RECT 357.640 -14.170 358.940 -13.910 ;
        RECT 399.220 -14.170 400.520 -13.910 ;
        RECT 440.800 -14.170 442.100 -13.910 ;
        RECT 316.060 -22.010 317.360 -21.750 ;
        RECT 357.640 -22.010 358.940 -21.750 ;
        RECT 399.220 -22.010 400.520 -21.750 ;
        RECT 440.800 -22.010 442.100 -21.750 ;
        RECT 316.060 -29.850 317.360 -29.590 ;
        RECT 357.640 -29.850 358.940 -29.590 ;
        RECT 399.220 -29.850 400.520 -29.590 ;
        RECT 440.800 -29.850 442.100 -29.590 ;
        RECT 316.060 -37.690 317.360 -37.430 ;
        RECT 357.640 -37.690 358.940 -37.430 ;
        RECT 399.220 -37.690 400.520 -37.430 ;
        RECT 440.800 -37.690 442.100 -37.430 ;
        RECT 316.060 -45.530 317.360 -45.270 ;
        RECT 357.640 -45.530 358.940 -45.270 ;
        RECT 399.220 -45.530 400.520 -45.270 ;
        RECT 440.800 -45.530 442.100 -45.270 ;
        RECT -488.400 -84.715 -487.620 -84.455 ;
        RECT -492.280 -86.245 -491.500 -85.985 ;
        RECT -491.760 -88.955 -491.500 -88.175 ;
        RECT -485.820 -88.955 -485.560 -88.175 ;
        RECT -487.815 -96.505 -487.555 -95.725 ;
        RECT 144.920 -97.120 145.180 -96.860 ;
        RECT 142.325 -118.060 142.585 -117.800 ;
        RECT 142.945 -118.060 143.205 -117.800 ;
        RECT 142.325 -118.680 142.585 -118.420 ;
        RECT 142.945 -118.680 143.205 -118.420 ;
        RECT 142.325 -119.300 142.585 -119.040 ;
        RECT 142.945 -119.300 143.205 -119.040 ;
        RECT 142.325 -119.920 142.585 -119.660 ;
        RECT 142.945 -119.920 143.205 -119.660 ;
        RECT 142.325 -120.540 142.585 -120.280 ;
        RECT 142.945 -120.540 143.205 -120.280 ;
        RECT 142.325 -121.160 142.585 -120.900 ;
        RECT 142.945 -121.160 143.205 -120.900 ;
        RECT 142.325 -121.780 142.585 -121.520 ;
        RECT 142.945 -121.780 143.205 -121.520 ;
        RECT 142.325 -122.400 142.585 -122.140 ;
        RECT 142.945 -122.400 143.205 -122.140 ;
      LAYER Metal2 ;
        RECT 142.145 117.620 143.385 122.580 ;
        RECT 164.720 117.620 170.920 122.580 ;
        RECT -487.875 96.315 -487.495 97.615 ;
        RECT -485.885 96.315 -485.495 98.115 ;
        RECT 167.490 97.190 168.150 117.620 ;
        RECT 144.850 96.790 168.150 97.190 ;
        RECT -487.875 95.915 -485.495 96.315 ;
        RECT -487.875 94.615 -487.495 95.915 ;
        RECT -485.885 94.890 -485.495 95.915 ;
        RECT -485.885 89.085 -484.285 94.890 ;
        RECT -491.830 88.045 -491.430 89.085 ;
        RECT -485.890 88.045 -484.285 89.085 ;
        RECT -491.820 86.305 -491.440 88.045 ;
        RECT -492.340 85.925 -491.440 86.305 ;
        RECT -485.885 85.890 -484.285 88.045 ;
        RECT -485.885 84.775 -485.495 85.890 ;
        RECT -488.465 84.395 -485.495 84.775 ;
        RECT 316.050 48.490 317.370 48.870 ;
        RECT 357.630 48.490 358.950 48.870 ;
        RECT 399.210 48.490 400.530 48.870 ;
        RECT 440.790 48.490 442.110 48.870 ;
        RECT 316.050 40.650 317.370 41.030 ;
        RECT 357.630 40.650 358.950 41.030 ;
        RECT 399.210 40.650 400.530 41.030 ;
        RECT 440.790 40.650 442.110 41.030 ;
        RECT 316.050 32.810 317.370 33.190 ;
        RECT 357.630 32.810 358.950 33.190 ;
        RECT 399.210 32.810 400.530 33.190 ;
        RECT 440.790 32.810 442.110 33.190 ;
        RECT 316.050 24.970 317.370 25.350 ;
        RECT 357.630 24.970 358.950 25.350 ;
        RECT 399.210 24.970 400.530 25.350 ;
        RECT 440.790 24.970 442.110 25.350 ;
        RECT 316.050 17.130 317.370 17.510 ;
        RECT 357.630 17.130 358.950 17.510 ;
        RECT 399.210 17.130 400.530 17.510 ;
        RECT 440.790 17.130 442.110 17.510 ;
        RECT 316.050 9.290 317.370 9.670 ;
        RECT 357.630 9.290 358.950 9.670 ;
        RECT 399.210 9.290 400.530 9.670 ;
        RECT 440.790 9.290 442.110 9.670 ;
        RECT 169.295 -7.000 169.795 7.000 ;
        RECT 316.050 1.450 317.370 1.830 ;
        RECT 357.630 1.450 358.950 1.830 ;
        RECT 399.210 1.450 400.530 1.830 ;
        RECT 440.790 1.450 442.110 1.830 ;
        RECT 316.050 -6.390 317.370 -6.010 ;
        RECT 357.630 -6.390 358.950 -6.010 ;
        RECT 399.210 -6.390 400.530 -6.010 ;
        RECT 440.790 -6.390 442.110 -6.010 ;
        RECT 316.050 -14.230 317.370 -13.850 ;
        RECT 357.630 -14.230 358.950 -13.850 ;
        RECT 399.210 -14.230 400.530 -13.850 ;
        RECT 440.790 -14.230 442.110 -13.850 ;
        RECT 316.050 -22.070 317.370 -21.690 ;
        RECT 357.630 -22.070 358.950 -21.690 ;
        RECT 399.210 -22.070 400.530 -21.690 ;
        RECT 440.790 -22.070 442.110 -21.690 ;
        RECT 316.050 -29.910 317.370 -29.530 ;
        RECT 357.630 -29.910 358.950 -29.530 ;
        RECT 399.210 -29.910 400.530 -29.530 ;
        RECT 440.790 -29.910 442.110 -29.530 ;
        RECT 316.050 -37.750 317.370 -37.370 ;
        RECT 357.630 -37.750 358.950 -37.370 ;
        RECT 399.210 -37.750 400.530 -37.370 ;
        RECT 440.790 -37.750 442.110 -37.370 ;
        RECT 316.050 -45.590 317.370 -45.210 ;
        RECT 357.630 -45.590 358.950 -45.210 ;
        RECT 399.210 -45.590 400.530 -45.210 ;
        RECT 440.790 -45.590 442.110 -45.210 ;
        RECT -488.465 -84.775 -485.495 -84.395 ;
        RECT -485.885 -85.890 -485.495 -84.775 ;
        RECT -492.340 -86.305 -491.440 -85.925 ;
        RECT -491.820 -88.045 -491.440 -86.305 ;
        RECT -485.885 -88.045 -484.285 -85.890 ;
        RECT -491.830 -89.085 -491.430 -88.045 ;
        RECT -485.890 -89.085 -484.285 -88.045 ;
        RECT -487.875 -95.915 -487.495 -94.615 ;
        RECT -485.885 -94.890 -484.285 -89.085 ;
        RECT -485.885 -95.915 -485.495 -94.890 ;
        RECT -487.875 -96.315 -485.495 -95.915 ;
        RECT -487.875 -97.615 -487.495 -96.315 ;
        RECT -485.885 -98.115 -485.495 -96.315 ;
        RECT 144.850 -97.190 168.150 -96.790 ;
        RECT 167.490 -117.620 168.150 -97.190 ;
        RECT 142.145 -122.580 143.385 -117.620 ;
        RECT 164.720 -122.580 170.920 -117.620 ;
      LAYER Via2 ;
        RECT 142.315 122.130 142.595 122.410 ;
        RECT 142.935 122.130 143.215 122.410 ;
        RECT 142.315 121.510 142.595 121.790 ;
        RECT 142.935 121.510 143.215 121.790 ;
        RECT 142.315 120.890 142.595 121.170 ;
        RECT 142.935 120.890 143.215 121.170 ;
        RECT 142.315 120.270 142.595 120.550 ;
        RECT 142.935 120.270 143.215 120.550 ;
        RECT 142.315 119.650 142.595 119.930 ;
        RECT 142.935 119.650 143.215 119.930 ;
        RECT 142.315 119.030 142.595 119.310 ;
        RECT 142.935 119.030 143.215 119.310 ;
        RECT 142.315 118.410 142.595 118.690 ;
        RECT 142.935 118.410 143.215 118.690 ;
        RECT 142.315 117.790 142.595 118.070 ;
        RECT 142.935 117.790 143.215 118.070 ;
        RECT 164.890 122.130 165.170 122.410 ;
        RECT 165.510 122.130 165.790 122.410 ;
        RECT 166.130 122.130 166.410 122.410 ;
        RECT 166.750 122.130 167.030 122.410 ;
        RECT 167.370 122.130 167.650 122.410 ;
        RECT 167.990 122.130 168.270 122.410 ;
        RECT 168.610 122.130 168.890 122.410 ;
        RECT 169.230 122.130 169.510 122.410 ;
        RECT 169.850 122.130 170.130 122.410 ;
        RECT 170.470 122.130 170.750 122.410 ;
        RECT 164.890 121.510 165.170 121.790 ;
        RECT 165.510 121.510 165.790 121.790 ;
        RECT 166.130 121.510 166.410 121.790 ;
        RECT 166.750 121.510 167.030 121.790 ;
        RECT 167.370 121.510 167.650 121.790 ;
        RECT 167.990 121.510 168.270 121.790 ;
        RECT 168.610 121.510 168.890 121.790 ;
        RECT 169.230 121.510 169.510 121.790 ;
        RECT 169.850 121.510 170.130 121.790 ;
        RECT 170.470 121.510 170.750 121.790 ;
        RECT 164.890 120.890 165.170 121.170 ;
        RECT 165.510 120.890 165.790 121.170 ;
        RECT 166.130 120.890 166.410 121.170 ;
        RECT 166.750 120.890 167.030 121.170 ;
        RECT 167.370 120.890 167.650 121.170 ;
        RECT 167.990 120.890 168.270 121.170 ;
        RECT 168.610 120.890 168.890 121.170 ;
        RECT 169.230 120.890 169.510 121.170 ;
        RECT 169.850 120.890 170.130 121.170 ;
        RECT 170.470 120.890 170.750 121.170 ;
        RECT 164.890 120.270 165.170 120.550 ;
        RECT 165.510 120.270 165.790 120.550 ;
        RECT 166.130 120.270 166.410 120.550 ;
        RECT 166.750 120.270 167.030 120.550 ;
        RECT 167.370 120.270 167.650 120.550 ;
        RECT 167.990 120.270 168.270 120.550 ;
        RECT 168.610 120.270 168.890 120.550 ;
        RECT 169.230 120.270 169.510 120.550 ;
        RECT 169.850 120.270 170.130 120.550 ;
        RECT 170.470 120.270 170.750 120.550 ;
        RECT 164.890 119.650 165.170 119.930 ;
        RECT 165.510 119.650 165.790 119.930 ;
        RECT 166.130 119.650 166.410 119.930 ;
        RECT 166.750 119.650 167.030 119.930 ;
        RECT 167.370 119.650 167.650 119.930 ;
        RECT 167.990 119.650 168.270 119.930 ;
        RECT 168.610 119.650 168.890 119.930 ;
        RECT 169.230 119.650 169.510 119.930 ;
        RECT 169.850 119.650 170.130 119.930 ;
        RECT 170.470 119.650 170.750 119.930 ;
        RECT 164.890 119.030 165.170 119.310 ;
        RECT 165.510 119.030 165.790 119.310 ;
        RECT 166.130 119.030 166.410 119.310 ;
        RECT 166.750 119.030 167.030 119.310 ;
        RECT 167.370 119.030 167.650 119.310 ;
        RECT 167.990 119.030 168.270 119.310 ;
        RECT 168.610 119.030 168.890 119.310 ;
        RECT 169.230 119.030 169.510 119.310 ;
        RECT 169.850 119.030 170.130 119.310 ;
        RECT 170.470 119.030 170.750 119.310 ;
        RECT 164.890 118.410 165.170 118.690 ;
        RECT 165.510 118.410 165.790 118.690 ;
        RECT 166.130 118.410 166.410 118.690 ;
        RECT 166.750 118.410 167.030 118.690 ;
        RECT 167.370 118.410 167.650 118.690 ;
        RECT 167.990 118.410 168.270 118.690 ;
        RECT 168.610 118.410 168.890 118.690 ;
        RECT 169.230 118.410 169.510 118.690 ;
        RECT 169.850 118.410 170.130 118.690 ;
        RECT 170.470 118.410 170.750 118.690 ;
        RECT 164.890 117.790 165.170 118.070 ;
        RECT 165.510 117.790 165.790 118.070 ;
        RECT 166.130 117.790 166.410 118.070 ;
        RECT 166.750 117.790 167.030 118.070 ;
        RECT 167.370 117.790 167.650 118.070 ;
        RECT 167.990 117.790 168.270 118.070 ;
        RECT 168.610 117.790 168.890 118.070 ;
        RECT 169.230 117.790 169.510 118.070 ;
        RECT 169.850 117.790 170.130 118.070 ;
        RECT 170.470 117.790 170.750 118.070 ;
        RECT -485.745 92.210 -484.425 94.570 ;
        RECT -485.745 89.210 -484.425 91.570 ;
        RECT -485.745 86.210 -484.425 88.570 ;
        RECT 316.050 48.540 317.370 48.820 ;
        RECT 357.630 48.540 358.950 48.820 ;
        RECT 399.210 48.540 400.530 48.820 ;
        RECT 440.790 48.540 442.110 48.820 ;
        RECT 316.050 40.700 317.370 40.980 ;
        RECT 357.630 40.700 358.950 40.980 ;
        RECT 399.210 40.700 400.530 40.980 ;
        RECT 440.790 40.700 442.110 40.980 ;
        RECT 316.050 32.860 317.370 33.140 ;
        RECT 357.630 32.860 358.950 33.140 ;
        RECT 399.210 32.860 400.530 33.140 ;
        RECT 440.790 32.860 442.110 33.140 ;
        RECT 316.050 25.020 317.370 25.300 ;
        RECT 357.630 25.020 358.950 25.300 ;
        RECT 399.210 25.020 400.530 25.300 ;
        RECT 440.790 25.020 442.110 25.300 ;
        RECT 316.050 17.180 317.370 17.460 ;
        RECT 357.630 17.180 358.950 17.460 ;
        RECT 399.210 17.180 400.530 17.460 ;
        RECT 440.790 17.180 442.110 17.460 ;
        RECT 316.050 9.340 317.370 9.620 ;
        RECT 357.630 9.340 358.950 9.620 ;
        RECT 399.210 9.340 400.530 9.620 ;
        RECT 440.790 9.340 442.110 9.620 ;
        RECT 169.405 -6.640 169.685 6.640 ;
        RECT 316.050 1.500 317.370 1.780 ;
        RECT 357.630 1.500 358.950 1.780 ;
        RECT 399.210 1.500 400.530 1.780 ;
        RECT 440.790 1.500 442.110 1.780 ;
        RECT 316.050 -6.340 317.370 -6.060 ;
        RECT 357.630 -6.340 358.950 -6.060 ;
        RECT 399.210 -6.340 400.530 -6.060 ;
        RECT 440.790 -6.340 442.110 -6.060 ;
        RECT 316.050 -14.180 317.370 -13.900 ;
        RECT 357.630 -14.180 358.950 -13.900 ;
        RECT 399.210 -14.180 400.530 -13.900 ;
        RECT 440.790 -14.180 442.110 -13.900 ;
        RECT 316.050 -22.020 317.370 -21.740 ;
        RECT 357.630 -22.020 358.950 -21.740 ;
        RECT 399.210 -22.020 400.530 -21.740 ;
        RECT 440.790 -22.020 442.110 -21.740 ;
        RECT 316.050 -29.860 317.370 -29.580 ;
        RECT 357.630 -29.860 358.950 -29.580 ;
        RECT 399.210 -29.860 400.530 -29.580 ;
        RECT 440.790 -29.860 442.110 -29.580 ;
        RECT 316.050 -37.700 317.370 -37.420 ;
        RECT 357.630 -37.700 358.950 -37.420 ;
        RECT 399.210 -37.700 400.530 -37.420 ;
        RECT 440.790 -37.700 442.110 -37.420 ;
        RECT 316.050 -45.540 317.370 -45.260 ;
        RECT 357.630 -45.540 358.950 -45.260 ;
        RECT 399.210 -45.540 400.530 -45.260 ;
        RECT 440.790 -45.540 442.110 -45.260 ;
        RECT -485.745 -88.570 -484.425 -86.210 ;
        RECT -485.745 -91.570 -484.425 -89.210 ;
        RECT -485.745 -94.570 -484.425 -92.210 ;
        RECT 142.315 -118.070 142.595 -117.790 ;
        RECT 142.935 -118.070 143.215 -117.790 ;
        RECT 142.315 -118.690 142.595 -118.410 ;
        RECT 142.935 -118.690 143.215 -118.410 ;
        RECT 142.315 -119.310 142.595 -119.030 ;
        RECT 142.935 -119.310 143.215 -119.030 ;
        RECT 142.315 -119.930 142.595 -119.650 ;
        RECT 142.935 -119.930 143.215 -119.650 ;
        RECT 142.315 -120.550 142.595 -120.270 ;
        RECT 142.935 -120.550 143.215 -120.270 ;
        RECT 142.315 -121.170 142.595 -120.890 ;
        RECT 142.935 -121.170 143.215 -120.890 ;
        RECT 142.315 -121.790 142.595 -121.510 ;
        RECT 142.935 -121.790 143.215 -121.510 ;
        RECT 142.315 -122.410 142.595 -122.130 ;
        RECT 142.935 -122.410 143.215 -122.130 ;
        RECT 164.890 -118.070 165.170 -117.790 ;
        RECT 165.510 -118.070 165.790 -117.790 ;
        RECT 166.130 -118.070 166.410 -117.790 ;
        RECT 166.750 -118.070 167.030 -117.790 ;
        RECT 167.370 -118.070 167.650 -117.790 ;
        RECT 167.990 -118.070 168.270 -117.790 ;
        RECT 168.610 -118.070 168.890 -117.790 ;
        RECT 169.230 -118.070 169.510 -117.790 ;
        RECT 169.850 -118.070 170.130 -117.790 ;
        RECT 170.470 -118.070 170.750 -117.790 ;
        RECT 164.890 -118.690 165.170 -118.410 ;
        RECT 165.510 -118.690 165.790 -118.410 ;
        RECT 166.130 -118.690 166.410 -118.410 ;
        RECT 166.750 -118.690 167.030 -118.410 ;
        RECT 167.370 -118.690 167.650 -118.410 ;
        RECT 167.990 -118.690 168.270 -118.410 ;
        RECT 168.610 -118.690 168.890 -118.410 ;
        RECT 169.230 -118.690 169.510 -118.410 ;
        RECT 169.850 -118.690 170.130 -118.410 ;
        RECT 170.470 -118.690 170.750 -118.410 ;
        RECT 164.890 -119.310 165.170 -119.030 ;
        RECT 165.510 -119.310 165.790 -119.030 ;
        RECT 166.130 -119.310 166.410 -119.030 ;
        RECT 166.750 -119.310 167.030 -119.030 ;
        RECT 167.370 -119.310 167.650 -119.030 ;
        RECT 167.990 -119.310 168.270 -119.030 ;
        RECT 168.610 -119.310 168.890 -119.030 ;
        RECT 169.230 -119.310 169.510 -119.030 ;
        RECT 169.850 -119.310 170.130 -119.030 ;
        RECT 170.470 -119.310 170.750 -119.030 ;
        RECT 164.890 -119.930 165.170 -119.650 ;
        RECT 165.510 -119.930 165.790 -119.650 ;
        RECT 166.130 -119.930 166.410 -119.650 ;
        RECT 166.750 -119.930 167.030 -119.650 ;
        RECT 167.370 -119.930 167.650 -119.650 ;
        RECT 167.990 -119.930 168.270 -119.650 ;
        RECT 168.610 -119.930 168.890 -119.650 ;
        RECT 169.230 -119.930 169.510 -119.650 ;
        RECT 169.850 -119.930 170.130 -119.650 ;
        RECT 170.470 -119.930 170.750 -119.650 ;
        RECT 164.890 -120.550 165.170 -120.270 ;
        RECT 165.510 -120.550 165.790 -120.270 ;
        RECT 166.130 -120.550 166.410 -120.270 ;
        RECT 166.750 -120.550 167.030 -120.270 ;
        RECT 167.370 -120.550 167.650 -120.270 ;
        RECT 167.990 -120.550 168.270 -120.270 ;
        RECT 168.610 -120.550 168.890 -120.270 ;
        RECT 169.230 -120.550 169.510 -120.270 ;
        RECT 169.850 -120.550 170.130 -120.270 ;
        RECT 170.470 -120.550 170.750 -120.270 ;
        RECT 164.890 -121.170 165.170 -120.890 ;
        RECT 165.510 -121.170 165.790 -120.890 ;
        RECT 166.130 -121.170 166.410 -120.890 ;
        RECT 166.750 -121.170 167.030 -120.890 ;
        RECT 167.370 -121.170 167.650 -120.890 ;
        RECT 167.990 -121.170 168.270 -120.890 ;
        RECT 168.610 -121.170 168.890 -120.890 ;
        RECT 169.230 -121.170 169.510 -120.890 ;
        RECT 169.850 -121.170 170.130 -120.890 ;
        RECT 170.470 -121.170 170.750 -120.890 ;
        RECT 164.890 -121.790 165.170 -121.510 ;
        RECT 165.510 -121.790 165.790 -121.510 ;
        RECT 166.130 -121.790 166.410 -121.510 ;
        RECT 166.750 -121.790 167.030 -121.510 ;
        RECT 167.370 -121.790 167.650 -121.510 ;
        RECT 167.990 -121.790 168.270 -121.510 ;
        RECT 168.610 -121.790 168.890 -121.510 ;
        RECT 169.230 -121.790 169.510 -121.510 ;
        RECT 169.850 -121.790 170.130 -121.510 ;
        RECT 170.470 -121.790 170.750 -121.510 ;
        RECT 164.890 -122.410 165.170 -122.130 ;
        RECT 165.510 -122.410 165.790 -122.130 ;
        RECT 166.130 -122.410 166.410 -122.130 ;
        RECT 166.750 -122.410 167.030 -122.130 ;
        RECT 167.370 -122.410 167.650 -122.130 ;
        RECT 167.990 -122.410 168.270 -122.130 ;
        RECT 168.610 -122.410 168.890 -122.130 ;
        RECT 169.230 -122.410 169.510 -122.130 ;
        RECT 169.850 -122.410 170.130 -122.130 ;
        RECT 170.470 -122.410 170.750 -122.130 ;
      LAYER Metal3 ;
        RECT 142.145 117.620 143.385 122.580 ;
        RECT 164.720 117.620 170.920 122.580 ;
        RECT -485.885 85.890 -484.285 94.890 ;
        RECT 316.000 48.540 317.420 48.820 ;
        RECT 357.580 48.540 359.000 48.820 ;
        RECT 399.160 48.540 400.580 48.820 ;
        RECT 440.740 48.540 442.160 48.820 ;
        RECT 316.000 40.700 317.420 40.980 ;
        RECT 357.580 40.700 359.000 40.980 ;
        RECT 399.160 40.700 400.580 40.980 ;
        RECT 440.740 40.700 442.160 40.980 ;
        RECT 316.000 32.860 317.420 33.140 ;
        RECT 357.580 32.860 359.000 33.140 ;
        RECT 399.160 32.860 400.580 33.140 ;
        RECT 440.740 32.860 442.160 33.140 ;
        RECT 316.000 25.020 317.420 25.300 ;
        RECT 357.580 25.020 359.000 25.300 ;
        RECT 399.160 25.020 400.580 25.300 ;
        RECT 440.740 25.020 442.160 25.300 ;
        RECT 316.000 17.180 317.420 17.460 ;
        RECT 357.580 17.180 359.000 17.460 ;
        RECT 399.160 17.180 400.580 17.460 ;
        RECT 440.740 17.180 442.160 17.460 ;
        RECT 168.220 8.000 169.820 10.500 ;
        RECT 316.000 9.340 317.420 9.620 ;
        RECT 357.580 9.340 359.000 9.620 ;
        RECT 399.160 9.340 400.580 9.620 ;
        RECT 440.740 9.340 442.160 9.620 ;
        RECT 168.220 -8.000 169.825 8.000 ;
        RECT 316.000 1.500 317.420 1.780 ;
        RECT 357.580 1.500 359.000 1.780 ;
        RECT 399.160 1.500 400.580 1.780 ;
        RECT 440.740 1.500 442.160 1.780 ;
        RECT 316.000 -6.340 317.420 -6.060 ;
        RECT 357.580 -6.340 359.000 -6.060 ;
        RECT 399.160 -6.340 400.580 -6.060 ;
        RECT 440.740 -6.340 442.160 -6.060 ;
        RECT 168.220 -10.500 169.820 -8.000 ;
        RECT 316.000 -14.180 317.420 -13.900 ;
        RECT 357.580 -14.180 359.000 -13.900 ;
        RECT 399.160 -14.180 400.580 -13.900 ;
        RECT 440.740 -14.180 442.160 -13.900 ;
        RECT 316.000 -22.020 317.420 -21.740 ;
        RECT 357.580 -22.020 359.000 -21.740 ;
        RECT 399.160 -22.020 400.580 -21.740 ;
        RECT 440.740 -22.020 442.160 -21.740 ;
        RECT 316.000 -29.860 317.420 -29.580 ;
        RECT 357.580 -29.860 359.000 -29.580 ;
        RECT 399.160 -29.860 400.580 -29.580 ;
        RECT 440.740 -29.860 442.160 -29.580 ;
        RECT 316.000 -37.700 317.420 -37.420 ;
        RECT 357.580 -37.700 359.000 -37.420 ;
        RECT 399.160 -37.700 400.580 -37.420 ;
        RECT 440.740 -37.700 442.160 -37.420 ;
        RECT 316.000 -45.540 317.420 -45.260 ;
        RECT 357.580 -45.540 359.000 -45.260 ;
        RECT 399.160 -45.540 400.580 -45.260 ;
        RECT 440.740 -45.540 442.160 -45.260 ;
        RECT -485.885 -94.890 -484.285 -85.890 ;
        RECT 142.145 -122.580 143.385 -117.620 ;
        RECT 164.720 -122.580 170.920 -117.620 ;
      LAYER Via3 ;
        RECT 142.315 122.130 142.595 122.410 ;
        RECT 142.935 122.130 143.215 122.410 ;
        RECT 142.315 121.510 142.595 121.790 ;
        RECT 142.935 121.510 143.215 121.790 ;
        RECT 142.315 120.890 142.595 121.170 ;
        RECT 142.935 120.890 143.215 121.170 ;
        RECT 142.315 120.270 142.595 120.550 ;
        RECT 142.935 120.270 143.215 120.550 ;
        RECT 142.315 119.650 142.595 119.930 ;
        RECT 142.935 119.650 143.215 119.930 ;
        RECT 142.315 119.030 142.595 119.310 ;
        RECT 142.935 119.030 143.215 119.310 ;
        RECT 142.315 118.410 142.595 118.690 ;
        RECT 142.935 118.410 143.215 118.690 ;
        RECT 142.315 117.790 142.595 118.070 ;
        RECT 142.935 117.790 143.215 118.070 ;
        RECT 164.890 122.130 165.170 122.410 ;
        RECT 165.510 122.130 165.790 122.410 ;
        RECT 166.130 122.130 166.410 122.410 ;
        RECT 166.750 122.130 167.030 122.410 ;
        RECT 167.370 122.130 167.650 122.410 ;
        RECT 167.990 122.130 168.270 122.410 ;
        RECT 168.610 122.130 168.890 122.410 ;
        RECT 169.230 122.130 169.510 122.410 ;
        RECT 169.850 122.130 170.130 122.410 ;
        RECT 170.470 122.130 170.750 122.410 ;
        RECT 164.890 121.510 165.170 121.790 ;
        RECT 165.510 121.510 165.790 121.790 ;
        RECT 166.130 121.510 166.410 121.790 ;
        RECT 166.750 121.510 167.030 121.790 ;
        RECT 167.370 121.510 167.650 121.790 ;
        RECT 167.990 121.510 168.270 121.790 ;
        RECT 168.610 121.510 168.890 121.790 ;
        RECT 169.230 121.510 169.510 121.790 ;
        RECT 169.850 121.510 170.130 121.790 ;
        RECT 170.470 121.510 170.750 121.790 ;
        RECT 164.890 120.890 165.170 121.170 ;
        RECT 165.510 120.890 165.790 121.170 ;
        RECT 166.130 120.890 166.410 121.170 ;
        RECT 166.750 120.890 167.030 121.170 ;
        RECT 167.370 120.890 167.650 121.170 ;
        RECT 167.990 120.890 168.270 121.170 ;
        RECT 168.610 120.890 168.890 121.170 ;
        RECT 169.230 120.890 169.510 121.170 ;
        RECT 169.850 120.890 170.130 121.170 ;
        RECT 170.470 120.890 170.750 121.170 ;
        RECT 164.890 120.270 165.170 120.550 ;
        RECT 165.510 120.270 165.790 120.550 ;
        RECT 166.130 120.270 166.410 120.550 ;
        RECT 166.750 120.270 167.030 120.550 ;
        RECT 167.370 120.270 167.650 120.550 ;
        RECT 167.990 120.270 168.270 120.550 ;
        RECT 168.610 120.270 168.890 120.550 ;
        RECT 169.230 120.270 169.510 120.550 ;
        RECT 169.850 120.270 170.130 120.550 ;
        RECT 170.470 120.270 170.750 120.550 ;
        RECT 164.890 119.650 165.170 119.930 ;
        RECT 165.510 119.650 165.790 119.930 ;
        RECT 166.130 119.650 166.410 119.930 ;
        RECT 166.750 119.650 167.030 119.930 ;
        RECT 167.370 119.650 167.650 119.930 ;
        RECT 167.990 119.650 168.270 119.930 ;
        RECT 168.610 119.650 168.890 119.930 ;
        RECT 169.230 119.650 169.510 119.930 ;
        RECT 169.850 119.650 170.130 119.930 ;
        RECT 170.470 119.650 170.750 119.930 ;
        RECT 164.890 119.030 165.170 119.310 ;
        RECT 165.510 119.030 165.790 119.310 ;
        RECT 166.130 119.030 166.410 119.310 ;
        RECT 166.750 119.030 167.030 119.310 ;
        RECT 167.370 119.030 167.650 119.310 ;
        RECT 167.990 119.030 168.270 119.310 ;
        RECT 168.610 119.030 168.890 119.310 ;
        RECT 169.230 119.030 169.510 119.310 ;
        RECT 169.850 119.030 170.130 119.310 ;
        RECT 170.470 119.030 170.750 119.310 ;
        RECT 164.890 118.410 165.170 118.690 ;
        RECT 165.510 118.410 165.790 118.690 ;
        RECT 166.130 118.410 166.410 118.690 ;
        RECT 166.750 118.410 167.030 118.690 ;
        RECT 167.370 118.410 167.650 118.690 ;
        RECT 167.990 118.410 168.270 118.690 ;
        RECT 168.610 118.410 168.890 118.690 ;
        RECT 169.230 118.410 169.510 118.690 ;
        RECT 169.850 118.410 170.130 118.690 ;
        RECT 170.470 118.410 170.750 118.690 ;
        RECT 164.890 117.790 165.170 118.070 ;
        RECT 165.510 117.790 165.790 118.070 ;
        RECT 166.130 117.790 166.410 118.070 ;
        RECT 166.750 117.790 167.030 118.070 ;
        RECT 167.370 117.790 167.650 118.070 ;
        RECT 167.990 117.790 168.270 118.070 ;
        RECT 168.610 117.790 168.890 118.070 ;
        RECT 169.230 117.790 169.510 118.070 ;
        RECT 169.850 117.790 170.130 118.070 ;
        RECT 170.470 117.790 170.750 118.070 ;
        RECT -485.745 92.210 -484.425 94.570 ;
        RECT -485.745 89.210 -484.425 91.570 ;
        RECT -485.745 86.210 -484.425 88.570 ;
        RECT 316.050 48.540 317.370 48.820 ;
        RECT 357.630 48.540 358.950 48.820 ;
        RECT 399.210 48.540 400.530 48.820 ;
        RECT 440.790 48.540 442.110 48.820 ;
        RECT 316.050 40.700 317.370 40.980 ;
        RECT 357.630 40.700 358.950 40.980 ;
        RECT 399.210 40.700 400.530 40.980 ;
        RECT 440.790 40.700 442.110 40.980 ;
        RECT 316.050 32.860 317.370 33.140 ;
        RECT 357.630 32.860 358.950 33.140 ;
        RECT 399.210 32.860 400.530 33.140 ;
        RECT 440.790 32.860 442.110 33.140 ;
        RECT 316.050 25.020 317.370 25.300 ;
        RECT 357.630 25.020 358.950 25.300 ;
        RECT 399.210 25.020 400.530 25.300 ;
        RECT 440.790 25.020 442.110 25.300 ;
        RECT 316.050 17.180 317.370 17.460 ;
        RECT 357.630 17.180 358.950 17.460 ;
        RECT 399.210 17.180 400.530 17.460 ;
        RECT 440.790 17.180 442.110 17.460 ;
        RECT 168.360 7.820 169.680 10.180 ;
        RECT 316.050 9.340 317.370 9.620 ;
        RECT 357.630 9.340 358.950 9.620 ;
        RECT 399.210 9.340 400.530 9.620 ;
        RECT 440.790 9.340 442.110 9.620 ;
        RECT 168.360 4.820 169.680 7.180 ;
        RECT 168.360 1.820 169.680 4.180 ;
        RECT 316.050 1.500 317.370 1.780 ;
        RECT 357.630 1.500 358.950 1.780 ;
        RECT 399.210 1.500 400.530 1.780 ;
        RECT 440.790 1.500 442.110 1.780 ;
        RECT 168.360 -1.180 169.680 1.180 ;
        RECT 168.360 -4.180 169.680 -1.820 ;
        RECT 168.360 -7.180 169.680 -4.820 ;
        RECT 316.050 -6.340 317.370 -6.060 ;
        RECT 357.630 -6.340 358.950 -6.060 ;
        RECT 399.210 -6.340 400.530 -6.060 ;
        RECT 440.790 -6.340 442.110 -6.060 ;
        RECT 168.360 -10.180 169.680 -7.820 ;
        RECT 316.050 -14.180 317.370 -13.900 ;
        RECT 357.630 -14.180 358.950 -13.900 ;
        RECT 399.210 -14.180 400.530 -13.900 ;
        RECT 440.790 -14.180 442.110 -13.900 ;
        RECT 316.050 -22.020 317.370 -21.740 ;
        RECT 357.630 -22.020 358.950 -21.740 ;
        RECT 399.210 -22.020 400.530 -21.740 ;
        RECT 440.790 -22.020 442.110 -21.740 ;
        RECT 316.050 -29.860 317.370 -29.580 ;
        RECT 357.630 -29.860 358.950 -29.580 ;
        RECT 399.210 -29.860 400.530 -29.580 ;
        RECT 440.790 -29.860 442.110 -29.580 ;
        RECT 316.050 -37.700 317.370 -37.420 ;
        RECT 357.630 -37.700 358.950 -37.420 ;
        RECT 399.210 -37.700 400.530 -37.420 ;
        RECT 440.790 -37.700 442.110 -37.420 ;
        RECT 316.050 -45.540 317.370 -45.260 ;
        RECT 357.630 -45.540 358.950 -45.260 ;
        RECT 399.210 -45.540 400.530 -45.260 ;
        RECT 440.790 -45.540 442.110 -45.260 ;
        RECT -485.745 -88.570 -484.425 -86.210 ;
        RECT -485.745 -91.570 -484.425 -89.210 ;
        RECT -485.745 -94.570 -484.425 -92.210 ;
        RECT 142.315 -118.070 142.595 -117.790 ;
        RECT 142.935 -118.070 143.215 -117.790 ;
        RECT 142.315 -118.690 142.595 -118.410 ;
        RECT 142.935 -118.690 143.215 -118.410 ;
        RECT 142.315 -119.310 142.595 -119.030 ;
        RECT 142.935 -119.310 143.215 -119.030 ;
        RECT 142.315 -119.930 142.595 -119.650 ;
        RECT 142.935 -119.930 143.215 -119.650 ;
        RECT 142.315 -120.550 142.595 -120.270 ;
        RECT 142.935 -120.550 143.215 -120.270 ;
        RECT 142.315 -121.170 142.595 -120.890 ;
        RECT 142.935 -121.170 143.215 -120.890 ;
        RECT 142.315 -121.790 142.595 -121.510 ;
        RECT 142.935 -121.790 143.215 -121.510 ;
        RECT 142.315 -122.410 142.595 -122.130 ;
        RECT 142.935 -122.410 143.215 -122.130 ;
        RECT 164.890 -118.070 165.170 -117.790 ;
        RECT 165.510 -118.070 165.790 -117.790 ;
        RECT 166.130 -118.070 166.410 -117.790 ;
        RECT 166.750 -118.070 167.030 -117.790 ;
        RECT 167.370 -118.070 167.650 -117.790 ;
        RECT 167.990 -118.070 168.270 -117.790 ;
        RECT 168.610 -118.070 168.890 -117.790 ;
        RECT 169.230 -118.070 169.510 -117.790 ;
        RECT 169.850 -118.070 170.130 -117.790 ;
        RECT 170.470 -118.070 170.750 -117.790 ;
        RECT 164.890 -118.690 165.170 -118.410 ;
        RECT 165.510 -118.690 165.790 -118.410 ;
        RECT 166.130 -118.690 166.410 -118.410 ;
        RECT 166.750 -118.690 167.030 -118.410 ;
        RECT 167.370 -118.690 167.650 -118.410 ;
        RECT 167.990 -118.690 168.270 -118.410 ;
        RECT 168.610 -118.690 168.890 -118.410 ;
        RECT 169.230 -118.690 169.510 -118.410 ;
        RECT 169.850 -118.690 170.130 -118.410 ;
        RECT 170.470 -118.690 170.750 -118.410 ;
        RECT 164.890 -119.310 165.170 -119.030 ;
        RECT 165.510 -119.310 165.790 -119.030 ;
        RECT 166.130 -119.310 166.410 -119.030 ;
        RECT 166.750 -119.310 167.030 -119.030 ;
        RECT 167.370 -119.310 167.650 -119.030 ;
        RECT 167.990 -119.310 168.270 -119.030 ;
        RECT 168.610 -119.310 168.890 -119.030 ;
        RECT 169.230 -119.310 169.510 -119.030 ;
        RECT 169.850 -119.310 170.130 -119.030 ;
        RECT 170.470 -119.310 170.750 -119.030 ;
        RECT 164.890 -119.930 165.170 -119.650 ;
        RECT 165.510 -119.930 165.790 -119.650 ;
        RECT 166.130 -119.930 166.410 -119.650 ;
        RECT 166.750 -119.930 167.030 -119.650 ;
        RECT 167.370 -119.930 167.650 -119.650 ;
        RECT 167.990 -119.930 168.270 -119.650 ;
        RECT 168.610 -119.930 168.890 -119.650 ;
        RECT 169.230 -119.930 169.510 -119.650 ;
        RECT 169.850 -119.930 170.130 -119.650 ;
        RECT 170.470 -119.930 170.750 -119.650 ;
        RECT 164.890 -120.550 165.170 -120.270 ;
        RECT 165.510 -120.550 165.790 -120.270 ;
        RECT 166.130 -120.550 166.410 -120.270 ;
        RECT 166.750 -120.550 167.030 -120.270 ;
        RECT 167.370 -120.550 167.650 -120.270 ;
        RECT 167.990 -120.550 168.270 -120.270 ;
        RECT 168.610 -120.550 168.890 -120.270 ;
        RECT 169.230 -120.550 169.510 -120.270 ;
        RECT 169.850 -120.550 170.130 -120.270 ;
        RECT 170.470 -120.550 170.750 -120.270 ;
        RECT 164.890 -121.170 165.170 -120.890 ;
        RECT 165.510 -121.170 165.790 -120.890 ;
        RECT 166.130 -121.170 166.410 -120.890 ;
        RECT 166.750 -121.170 167.030 -120.890 ;
        RECT 167.370 -121.170 167.650 -120.890 ;
        RECT 167.990 -121.170 168.270 -120.890 ;
        RECT 168.610 -121.170 168.890 -120.890 ;
        RECT 169.230 -121.170 169.510 -120.890 ;
        RECT 169.850 -121.170 170.130 -120.890 ;
        RECT 170.470 -121.170 170.750 -120.890 ;
        RECT 164.890 -121.790 165.170 -121.510 ;
        RECT 165.510 -121.790 165.790 -121.510 ;
        RECT 166.130 -121.790 166.410 -121.510 ;
        RECT 166.750 -121.790 167.030 -121.510 ;
        RECT 167.370 -121.790 167.650 -121.510 ;
        RECT 167.990 -121.790 168.270 -121.510 ;
        RECT 168.610 -121.790 168.890 -121.510 ;
        RECT 169.230 -121.790 169.510 -121.510 ;
        RECT 169.850 -121.790 170.130 -121.510 ;
        RECT 170.470 -121.790 170.750 -121.510 ;
        RECT 164.890 -122.410 165.170 -122.130 ;
        RECT 165.510 -122.410 165.790 -122.130 ;
        RECT 166.130 -122.410 166.410 -122.130 ;
        RECT 166.750 -122.410 167.030 -122.130 ;
        RECT 167.370 -122.410 167.650 -122.130 ;
        RECT 167.990 -122.410 168.270 -122.130 ;
        RECT 168.610 -122.410 168.890 -122.130 ;
        RECT 169.230 -122.410 169.510 -122.130 ;
        RECT 169.850 -122.410 170.130 -122.130 ;
        RECT 170.470 -122.410 170.750 -122.130 ;
      LAYER Metal4 ;
        RECT -725.980 976.200 729.020 1051.200 ;
        RECT -725.980 414.600 -650.980 976.200 ;
        RECT -542.830 968.335 -539.830 976.200 ;
        RECT -507.130 968.335 -504.130 976.200 ;
        RECT -467.830 968.335 -464.830 976.200 ;
        RECT -432.130 968.335 -429.130 976.200 ;
        RECT -392.830 968.335 -389.830 976.200 ;
        RECT -357.130 968.335 -354.130 976.200 ;
        RECT -317.830 968.335 -314.830 976.200 ;
        RECT -282.130 968.335 -279.130 976.200 ;
        RECT -242.830 968.335 -239.830 976.200 ;
        RECT -207.130 968.335 -204.130 976.200 ;
        RECT -167.830 968.335 -164.830 976.200 ;
        RECT -132.130 968.335 -129.130 976.200 ;
        RECT -92.830 968.335 -89.830 976.200 ;
        RECT -57.130 968.335 -54.130 976.200 ;
        RECT -17.830 968.335 -14.830 976.200 ;
        RECT 17.870 968.335 20.870 976.200 ;
        RECT 57.170 968.335 60.170 976.200 ;
        RECT 92.870 968.335 95.870 976.200 ;
        RECT 132.170 968.335 135.170 976.200 ;
        RECT 167.870 968.335 170.870 976.200 ;
        RECT 207.170 968.335 210.170 976.200 ;
        RECT 242.870 968.335 245.870 976.200 ;
        RECT 282.170 968.335 285.170 976.200 ;
        RECT 317.870 968.335 320.870 976.200 ;
        RECT 357.170 968.335 360.170 976.200 ;
        RECT 392.870 968.335 395.870 976.200 ;
        RECT 432.170 968.335 435.170 976.200 ;
        RECT 467.870 968.335 470.870 976.200 ;
        RECT 507.170 968.335 510.170 976.200 ;
        RECT 542.870 968.335 545.870 976.200 ;
        RECT 654.020 414.600 729.020 976.200 ;
        RECT -486.100 117.620 -479.900 122.580 ;
        RECT 142.145 117.620 143.385 122.580 ;
        RECT 164.720 117.620 170.920 122.580 ;
        RECT -484.695 94.890 -481.305 117.620 ;
        RECT -485.885 85.890 -481.305 94.890 ;
        RECT -484.695 -85.890 -481.305 85.890 ;
        RECT -485.885 -94.890 -481.305 -85.890 ;
        RECT -484.695 -117.620 -481.305 -94.890 ;
        RECT 165.820 -117.620 169.820 117.620 ;
        RECT -486.100 -122.580 -479.900 -117.620 ;
        RECT 142.145 -122.580 143.385 -117.620 ;
        RECT 164.720 -122.580 170.920 -117.620 ;
        RECT 315.910 -120.940 317.510 120.620 ;
        RECT 357.490 -120.940 359.090 120.620 ;
        RECT 399.070 -120.940 400.670 120.620 ;
        RECT 440.650 -120.940 442.250 120.620 ;
        RECT -725.980 -976.200 -650.980 -414.600 ;
        RECT -542.830 -976.200 -539.830 -968.335 ;
        RECT -507.130 -976.200 -504.130 -968.335 ;
        RECT -467.830 -976.200 -464.830 -968.335 ;
        RECT -432.130 -976.200 -429.130 -968.335 ;
        RECT -392.830 -976.200 -389.830 -968.335 ;
        RECT -357.130 -976.200 -354.130 -968.335 ;
        RECT -317.830 -976.200 -314.830 -968.335 ;
        RECT -282.130 -976.200 -279.130 -968.335 ;
        RECT -242.830 -976.200 -239.830 -968.335 ;
        RECT -207.130 -976.200 -204.130 -968.335 ;
        RECT -167.830 -976.200 -164.830 -968.335 ;
        RECT -132.130 -976.200 -129.130 -968.335 ;
        RECT -92.830 -976.200 -89.830 -968.335 ;
        RECT -57.130 -976.200 -54.130 -968.335 ;
        RECT -17.830 -976.200 -14.830 -968.335 ;
        RECT 17.870 -976.200 20.870 -968.335 ;
        RECT 57.170 -976.200 60.170 -968.335 ;
        RECT 92.870 -976.200 95.870 -968.335 ;
        RECT 132.170 -976.200 135.170 -968.335 ;
        RECT 167.870 -976.200 170.870 -968.335 ;
        RECT 207.170 -976.200 210.170 -968.335 ;
        RECT 242.870 -976.200 245.870 -968.335 ;
        RECT 282.170 -976.200 285.170 -968.335 ;
        RECT 317.870 -976.200 320.870 -968.335 ;
        RECT 357.170 -976.200 360.170 -968.335 ;
        RECT 392.870 -976.200 395.870 -968.335 ;
        RECT 432.170 -976.200 435.170 -968.335 ;
        RECT 467.870 -976.200 470.870 -968.335 ;
        RECT 507.170 -976.200 510.170 -968.335 ;
        RECT 542.870 -976.200 545.870 -968.335 ;
        RECT 654.020 -976.200 729.020 -414.600 ;
        RECT -725.980 -1051.200 729.020 -976.200 ;
      LAYER Via4 ;
        RECT -542.230 973.760 -541.950 974.040 ;
        RECT -541.470 973.760 -541.190 974.040 ;
        RECT -540.710 973.760 -540.430 974.040 ;
        RECT -542.230 973.000 -541.950 973.280 ;
        RECT -541.470 973.000 -541.190 973.280 ;
        RECT -540.710 973.000 -540.430 973.280 ;
        RECT -542.230 972.240 -541.950 972.520 ;
        RECT -541.470 972.240 -541.190 972.520 ;
        RECT -540.710 972.240 -540.430 972.520 ;
        RECT -542.230 971.480 -541.950 971.760 ;
        RECT -541.470 971.480 -541.190 971.760 ;
        RECT -540.710 971.480 -540.430 971.760 ;
        RECT -542.230 970.720 -541.950 971.000 ;
        RECT -541.470 970.720 -541.190 971.000 ;
        RECT -540.710 970.720 -540.430 971.000 ;
        RECT -542.230 969.960 -541.950 970.240 ;
        RECT -541.470 969.960 -541.190 970.240 ;
        RECT -540.710 969.960 -540.430 970.240 ;
        RECT -506.530 973.760 -506.250 974.040 ;
        RECT -505.770 973.760 -505.490 974.040 ;
        RECT -505.010 973.760 -504.730 974.040 ;
        RECT -506.530 973.000 -506.250 973.280 ;
        RECT -505.770 973.000 -505.490 973.280 ;
        RECT -505.010 973.000 -504.730 973.280 ;
        RECT -506.530 972.240 -506.250 972.520 ;
        RECT -505.770 972.240 -505.490 972.520 ;
        RECT -505.010 972.240 -504.730 972.520 ;
        RECT -506.530 971.480 -506.250 971.760 ;
        RECT -505.770 971.480 -505.490 971.760 ;
        RECT -505.010 971.480 -504.730 971.760 ;
        RECT -506.530 970.720 -506.250 971.000 ;
        RECT -505.770 970.720 -505.490 971.000 ;
        RECT -505.010 970.720 -504.730 971.000 ;
        RECT -506.530 969.960 -506.250 970.240 ;
        RECT -505.770 969.960 -505.490 970.240 ;
        RECT -505.010 969.960 -504.730 970.240 ;
        RECT -467.230 973.760 -466.950 974.040 ;
        RECT -466.470 973.760 -466.190 974.040 ;
        RECT -465.710 973.760 -465.430 974.040 ;
        RECT -467.230 973.000 -466.950 973.280 ;
        RECT -466.470 973.000 -466.190 973.280 ;
        RECT -465.710 973.000 -465.430 973.280 ;
        RECT -467.230 972.240 -466.950 972.520 ;
        RECT -466.470 972.240 -466.190 972.520 ;
        RECT -465.710 972.240 -465.430 972.520 ;
        RECT -467.230 971.480 -466.950 971.760 ;
        RECT -466.470 971.480 -466.190 971.760 ;
        RECT -465.710 971.480 -465.430 971.760 ;
        RECT -467.230 970.720 -466.950 971.000 ;
        RECT -466.470 970.720 -466.190 971.000 ;
        RECT -465.710 970.720 -465.430 971.000 ;
        RECT -467.230 969.960 -466.950 970.240 ;
        RECT -466.470 969.960 -466.190 970.240 ;
        RECT -465.710 969.960 -465.430 970.240 ;
        RECT -431.530 973.760 -431.250 974.040 ;
        RECT -430.770 973.760 -430.490 974.040 ;
        RECT -430.010 973.760 -429.730 974.040 ;
        RECT -431.530 973.000 -431.250 973.280 ;
        RECT -430.770 973.000 -430.490 973.280 ;
        RECT -430.010 973.000 -429.730 973.280 ;
        RECT -431.530 972.240 -431.250 972.520 ;
        RECT -430.770 972.240 -430.490 972.520 ;
        RECT -430.010 972.240 -429.730 972.520 ;
        RECT -431.530 971.480 -431.250 971.760 ;
        RECT -430.770 971.480 -430.490 971.760 ;
        RECT -430.010 971.480 -429.730 971.760 ;
        RECT -431.530 970.720 -431.250 971.000 ;
        RECT -430.770 970.720 -430.490 971.000 ;
        RECT -430.010 970.720 -429.730 971.000 ;
        RECT -431.530 969.960 -431.250 970.240 ;
        RECT -430.770 969.960 -430.490 970.240 ;
        RECT -430.010 969.960 -429.730 970.240 ;
        RECT -392.230 973.760 -391.950 974.040 ;
        RECT -391.470 973.760 -391.190 974.040 ;
        RECT -390.710 973.760 -390.430 974.040 ;
        RECT -392.230 973.000 -391.950 973.280 ;
        RECT -391.470 973.000 -391.190 973.280 ;
        RECT -390.710 973.000 -390.430 973.280 ;
        RECT -392.230 972.240 -391.950 972.520 ;
        RECT -391.470 972.240 -391.190 972.520 ;
        RECT -390.710 972.240 -390.430 972.520 ;
        RECT -392.230 971.480 -391.950 971.760 ;
        RECT -391.470 971.480 -391.190 971.760 ;
        RECT -390.710 971.480 -390.430 971.760 ;
        RECT -392.230 970.720 -391.950 971.000 ;
        RECT -391.470 970.720 -391.190 971.000 ;
        RECT -390.710 970.720 -390.430 971.000 ;
        RECT -392.230 969.960 -391.950 970.240 ;
        RECT -391.470 969.960 -391.190 970.240 ;
        RECT -390.710 969.960 -390.430 970.240 ;
        RECT -356.530 973.760 -356.250 974.040 ;
        RECT -355.770 973.760 -355.490 974.040 ;
        RECT -355.010 973.760 -354.730 974.040 ;
        RECT -356.530 973.000 -356.250 973.280 ;
        RECT -355.770 973.000 -355.490 973.280 ;
        RECT -355.010 973.000 -354.730 973.280 ;
        RECT -356.530 972.240 -356.250 972.520 ;
        RECT -355.770 972.240 -355.490 972.520 ;
        RECT -355.010 972.240 -354.730 972.520 ;
        RECT -356.530 971.480 -356.250 971.760 ;
        RECT -355.770 971.480 -355.490 971.760 ;
        RECT -355.010 971.480 -354.730 971.760 ;
        RECT -356.530 970.720 -356.250 971.000 ;
        RECT -355.770 970.720 -355.490 971.000 ;
        RECT -355.010 970.720 -354.730 971.000 ;
        RECT -356.530 969.960 -356.250 970.240 ;
        RECT -355.770 969.960 -355.490 970.240 ;
        RECT -355.010 969.960 -354.730 970.240 ;
        RECT -317.230 973.760 -316.950 974.040 ;
        RECT -316.470 973.760 -316.190 974.040 ;
        RECT -315.710 973.760 -315.430 974.040 ;
        RECT -317.230 973.000 -316.950 973.280 ;
        RECT -316.470 973.000 -316.190 973.280 ;
        RECT -315.710 973.000 -315.430 973.280 ;
        RECT -317.230 972.240 -316.950 972.520 ;
        RECT -316.470 972.240 -316.190 972.520 ;
        RECT -315.710 972.240 -315.430 972.520 ;
        RECT -317.230 971.480 -316.950 971.760 ;
        RECT -316.470 971.480 -316.190 971.760 ;
        RECT -315.710 971.480 -315.430 971.760 ;
        RECT -317.230 970.720 -316.950 971.000 ;
        RECT -316.470 970.720 -316.190 971.000 ;
        RECT -315.710 970.720 -315.430 971.000 ;
        RECT -317.230 969.960 -316.950 970.240 ;
        RECT -316.470 969.960 -316.190 970.240 ;
        RECT -315.710 969.960 -315.430 970.240 ;
        RECT -281.530 973.760 -281.250 974.040 ;
        RECT -280.770 973.760 -280.490 974.040 ;
        RECT -280.010 973.760 -279.730 974.040 ;
        RECT -281.530 973.000 -281.250 973.280 ;
        RECT -280.770 973.000 -280.490 973.280 ;
        RECT -280.010 973.000 -279.730 973.280 ;
        RECT -281.530 972.240 -281.250 972.520 ;
        RECT -280.770 972.240 -280.490 972.520 ;
        RECT -280.010 972.240 -279.730 972.520 ;
        RECT -281.530 971.480 -281.250 971.760 ;
        RECT -280.770 971.480 -280.490 971.760 ;
        RECT -280.010 971.480 -279.730 971.760 ;
        RECT -281.530 970.720 -281.250 971.000 ;
        RECT -280.770 970.720 -280.490 971.000 ;
        RECT -280.010 970.720 -279.730 971.000 ;
        RECT -281.530 969.960 -281.250 970.240 ;
        RECT -280.770 969.960 -280.490 970.240 ;
        RECT -280.010 969.960 -279.730 970.240 ;
        RECT -242.230 973.760 -241.950 974.040 ;
        RECT -241.470 973.760 -241.190 974.040 ;
        RECT -240.710 973.760 -240.430 974.040 ;
        RECT -242.230 973.000 -241.950 973.280 ;
        RECT -241.470 973.000 -241.190 973.280 ;
        RECT -240.710 973.000 -240.430 973.280 ;
        RECT -242.230 972.240 -241.950 972.520 ;
        RECT -241.470 972.240 -241.190 972.520 ;
        RECT -240.710 972.240 -240.430 972.520 ;
        RECT -242.230 971.480 -241.950 971.760 ;
        RECT -241.470 971.480 -241.190 971.760 ;
        RECT -240.710 971.480 -240.430 971.760 ;
        RECT -242.230 970.720 -241.950 971.000 ;
        RECT -241.470 970.720 -241.190 971.000 ;
        RECT -240.710 970.720 -240.430 971.000 ;
        RECT -242.230 969.960 -241.950 970.240 ;
        RECT -241.470 969.960 -241.190 970.240 ;
        RECT -240.710 969.960 -240.430 970.240 ;
        RECT -206.530 973.760 -206.250 974.040 ;
        RECT -205.770 973.760 -205.490 974.040 ;
        RECT -205.010 973.760 -204.730 974.040 ;
        RECT -206.530 973.000 -206.250 973.280 ;
        RECT -205.770 973.000 -205.490 973.280 ;
        RECT -205.010 973.000 -204.730 973.280 ;
        RECT -206.530 972.240 -206.250 972.520 ;
        RECT -205.770 972.240 -205.490 972.520 ;
        RECT -205.010 972.240 -204.730 972.520 ;
        RECT -206.530 971.480 -206.250 971.760 ;
        RECT -205.770 971.480 -205.490 971.760 ;
        RECT -205.010 971.480 -204.730 971.760 ;
        RECT -206.530 970.720 -206.250 971.000 ;
        RECT -205.770 970.720 -205.490 971.000 ;
        RECT -205.010 970.720 -204.730 971.000 ;
        RECT -206.530 969.960 -206.250 970.240 ;
        RECT -205.770 969.960 -205.490 970.240 ;
        RECT -205.010 969.960 -204.730 970.240 ;
        RECT -167.230 973.760 -166.950 974.040 ;
        RECT -166.470 973.760 -166.190 974.040 ;
        RECT -165.710 973.760 -165.430 974.040 ;
        RECT -167.230 973.000 -166.950 973.280 ;
        RECT -166.470 973.000 -166.190 973.280 ;
        RECT -165.710 973.000 -165.430 973.280 ;
        RECT -167.230 972.240 -166.950 972.520 ;
        RECT -166.470 972.240 -166.190 972.520 ;
        RECT -165.710 972.240 -165.430 972.520 ;
        RECT -167.230 971.480 -166.950 971.760 ;
        RECT -166.470 971.480 -166.190 971.760 ;
        RECT -165.710 971.480 -165.430 971.760 ;
        RECT -167.230 970.720 -166.950 971.000 ;
        RECT -166.470 970.720 -166.190 971.000 ;
        RECT -165.710 970.720 -165.430 971.000 ;
        RECT -167.230 969.960 -166.950 970.240 ;
        RECT -166.470 969.960 -166.190 970.240 ;
        RECT -165.710 969.960 -165.430 970.240 ;
        RECT -131.530 973.760 -131.250 974.040 ;
        RECT -130.770 973.760 -130.490 974.040 ;
        RECT -130.010 973.760 -129.730 974.040 ;
        RECT -131.530 973.000 -131.250 973.280 ;
        RECT -130.770 973.000 -130.490 973.280 ;
        RECT -130.010 973.000 -129.730 973.280 ;
        RECT -131.530 972.240 -131.250 972.520 ;
        RECT -130.770 972.240 -130.490 972.520 ;
        RECT -130.010 972.240 -129.730 972.520 ;
        RECT -131.530 971.480 -131.250 971.760 ;
        RECT -130.770 971.480 -130.490 971.760 ;
        RECT -130.010 971.480 -129.730 971.760 ;
        RECT -131.530 970.720 -131.250 971.000 ;
        RECT -130.770 970.720 -130.490 971.000 ;
        RECT -130.010 970.720 -129.730 971.000 ;
        RECT -131.530 969.960 -131.250 970.240 ;
        RECT -130.770 969.960 -130.490 970.240 ;
        RECT -130.010 969.960 -129.730 970.240 ;
        RECT -92.230 973.760 -91.950 974.040 ;
        RECT -91.470 973.760 -91.190 974.040 ;
        RECT -90.710 973.760 -90.430 974.040 ;
        RECT -92.230 973.000 -91.950 973.280 ;
        RECT -91.470 973.000 -91.190 973.280 ;
        RECT -90.710 973.000 -90.430 973.280 ;
        RECT -92.230 972.240 -91.950 972.520 ;
        RECT -91.470 972.240 -91.190 972.520 ;
        RECT -90.710 972.240 -90.430 972.520 ;
        RECT -92.230 971.480 -91.950 971.760 ;
        RECT -91.470 971.480 -91.190 971.760 ;
        RECT -90.710 971.480 -90.430 971.760 ;
        RECT -92.230 970.720 -91.950 971.000 ;
        RECT -91.470 970.720 -91.190 971.000 ;
        RECT -90.710 970.720 -90.430 971.000 ;
        RECT -92.230 969.960 -91.950 970.240 ;
        RECT -91.470 969.960 -91.190 970.240 ;
        RECT -90.710 969.960 -90.430 970.240 ;
        RECT -56.530 973.760 -56.250 974.040 ;
        RECT -55.770 973.760 -55.490 974.040 ;
        RECT -55.010 973.760 -54.730 974.040 ;
        RECT -56.530 973.000 -56.250 973.280 ;
        RECT -55.770 973.000 -55.490 973.280 ;
        RECT -55.010 973.000 -54.730 973.280 ;
        RECT -56.530 972.240 -56.250 972.520 ;
        RECT -55.770 972.240 -55.490 972.520 ;
        RECT -55.010 972.240 -54.730 972.520 ;
        RECT -56.530 971.480 -56.250 971.760 ;
        RECT -55.770 971.480 -55.490 971.760 ;
        RECT -55.010 971.480 -54.730 971.760 ;
        RECT -56.530 970.720 -56.250 971.000 ;
        RECT -55.770 970.720 -55.490 971.000 ;
        RECT -55.010 970.720 -54.730 971.000 ;
        RECT -56.530 969.960 -56.250 970.240 ;
        RECT -55.770 969.960 -55.490 970.240 ;
        RECT -55.010 969.960 -54.730 970.240 ;
        RECT -17.230 973.760 -16.950 974.040 ;
        RECT -16.470 973.760 -16.190 974.040 ;
        RECT -15.710 973.760 -15.430 974.040 ;
        RECT -17.230 973.000 -16.950 973.280 ;
        RECT -16.470 973.000 -16.190 973.280 ;
        RECT -15.710 973.000 -15.430 973.280 ;
        RECT -17.230 972.240 -16.950 972.520 ;
        RECT -16.470 972.240 -16.190 972.520 ;
        RECT -15.710 972.240 -15.430 972.520 ;
        RECT -17.230 971.480 -16.950 971.760 ;
        RECT -16.470 971.480 -16.190 971.760 ;
        RECT -15.710 971.480 -15.430 971.760 ;
        RECT -17.230 970.720 -16.950 971.000 ;
        RECT -16.470 970.720 -16.190 971.000 ;
        RECT -15.710 970.720 -15.430 971.000 ;
        RECT -17.230 969.960 -16.950 970.240 ;
        RECT -16.470 969.960 -16.190 970.240 ;
        RECT -15.710 969.960 -15.430 970.240 ;
        RECT 18.470 973.760 18.750 974.040 ;
        RECT 19.230 973.760 19.510 974.040 ;
        RECT 19.990 973.760 20.270 974.040 ;
        RECT 18.470 973.000 18.750 973.280 ;
        RECT 19.230 973.000 19.510 973.280 ;
        RECT 19.990 973.000 20.270 973.280 ;
        RECT 18.470 972.240 18.750 972.520 ;
        RECT 19.230 972.240 19.510 972.520 ;
        RECT 19.990 972.240 20.270 972.520 ;
        RECT 18.470 971.480 18.750 971.760 ;
        RECT 19.230 971.480 19.510 971.760 ;
        RECT 19.990 971.480 20.270 971.760 ;
        RECT 18.470 970.720 18.750 971.000 ;
        RECT 19.230 970.720 19.510 971.000 ;
        RECT 19.990 970.720 20.270 971.000 ;
        RECT 18.470 969.960 18.750 970.240 ;
        RECT 19.230 969.960 19.510 970.240 ;
        RECT 19.990 969.960 20.270 970.240 ;
        RECT 57.770 973.760 58.050 974.040 ;
        RECT 58.530 973.760 58.810 974.040 ;
        RECT 59.290 973.760 59.570 974.040 ;
        RECT 57.770 973.000 58.050 973.280 ;
        RECT 58.530 973.000 58.810 973.280 ;
        RECT 59.290 973.000 59.570 973.280 ;
        RECT 57.770 972.240 58.050 972.520 ;
        RECT 58.530 972.240 58.810 972.520 ;
        RECT 59.290 972.240 59.570 972.520 ;
        RECT 57.770 971.480 58.050 971.760 ;
        RECT 58.530 971.480 58.810 971.760 ;
        RECT 59.290 971.480 59.570 971.760 ;
        RECT 57.770 970.720 58.050 971.000 ;
        RECT 58.530 970.720 58.810 971.000 ;
        RECT 59.290 970.720 59.570 971.000 ;
        RECT 57.770 969.960 58.050 970.240 ;
        RECT 58.530 969.960 58.810 970.240 ;
        RECT 59.290 969.960 59.570 970.240 ;
        RECT 93.470 973.760 93.750 974.040 ;
        RECT 94.230 973.760 94.510 974.040 ;
        RECT 94.990 973.760 95.270 974.040 ;
        RECT 93.470 973.000 93.750 973.280 ;
        RECT 94.230 973.000 94.510 973.280 ;
        RECT 94.990 973.000 95.270 973.280 ;
        RECT 93.470 972.240 93.750 972.520 ;
        RECT 94.230 972.240 94.510 972.520 ;
        RECT 94.990 972.240 95.270 972.520 ;
        RECT 93.470 971.480 93.750 971.760 ;
        RECT 94.230 971.480 94.510 971.760 ;
        RECT 94.990 971.480 95.270 971.760 ;
        RECT 93.470 970.720 93.750 971.000 ;
        RECT 94.230 970.720 94.510 971.000 ;
        RECT 94.990 970.720 95.270 971.000 ;
        RECT 93.470 969.960 93.750 970.240 ;
        RECT 94.230 969.960 94.510 970.240 ;
        RECT 94.990 969.960 95.270 970.240 ;
        RECT 132.770 973.760 133.050 974.040 ;
        RECT 133.530 973.760 133.810 974.040 ;
        RECT 134.290 973.760 134.570 974.040 ;
        RECT 132.770 973.000 133.050 973.280 ;
        RECT 133.530 973.000 133.810 973.280 ;
        RECT 134.290 973.000 134.570 973.280 ;
        RECT 132.770 972.240 133.050 972.520 ;
        RECT 133.530 972.240 133.810 972.520 ;
        RECT 134.290 972.240 134.570 972.520 ;
        RECT 132.770 971.480 133.050 971.760 ;
        RECT 133.530 971.480 133.810 971.760 ;
        RECT 134.290 971.480 134.570 971.760 ;
        RECT 132.770 970.720 133.050 971.000 ;
        RECT 133.530 970.720 133.810 971.000 ;
        RECT 134.290 970.720 134.570 971.000 ;
        RECT 132.770 969.960 133.050 970.240 ;
        RECT 133.530 969.960 133.810 970.240 ;
        RECT 134.290 969.960 134.570 970.240 ;
        RECT 168.470 973.760 168.750 974.040 ;
        RECT 169.230 973.760 169.510 974.040 ;
        RECT 169.990 973.760 170.270 974.040 ;
        RECT 168.470 973.000 168.750 973.280 ;
        RECT 169.230 973.000 169.510 973.280 ;
        RECT 169.990 973.000 170.270 973.280 ;
        RECT 168.470 972.240 168.750 972.520 ;
        RECT 169.230 972.240 169.510 972.520 ;
        RECT 169.990 972.240 170.270 972.520 ;
        RECT 168.470 971.480 168.750 971.760 ;
        RECT 169.230 971.480 169.510 971.760 ;
        RECT 169.990 971.480 170.270 971.760 ;
        RECT 168.470 970.720 168.750 971.000 ;
        RECT 169.230 970.720 169.510 971.000 ;
        RECT 169.990 970.720 170.270 971.000 ;
        RECT 168.470 969.960 168.750 970.240 ;
        RECT 169.230 969.960 169.510 970.240 ;
        RECT 169.990 969.960 170.270 970.240 ;
        RECT 207.770 973.760 208.050 974.040 ;
        RECT 208.530 973.760 208.810 974.040 ;
        RECT 209.290 973.760 209.570 974.040 ;
        RECT 207.770 973.000 208.050 973.280 ;
        RECT 208.530 973.000 208.810 973.280 ;
        RECT 209.290 973.000 209.570 973.280 ;
        RECT 207.770 972.240 208.050 972.520 ;
        RECT 208.530 972.240 208.810 972.520 ;
        RECT 209.290 972.240 209.570 972.520 ;
        RECT 207.770 971.480 208.050 971.760 ;
        RECT 208.530 971.480 208.810 971.760 ;
        RECT 209.290 971.480 209.570 971.760 ;
        RECT 207.770 970.720 208.050 971.000 ;
        RECT 208.530 970.720 208.810 971.000 ;
        RECT 209.290 970.720 209.570 971.000 ;
        RECT 207.770 969.960 208.050 970.240 ;
        RECT 208.530 969.960 208.810 970.240 ;
        RECT 209.290 969.960 209.570 970.240 ;
        RECT 243.470 973.760 243.750 974.040 ;
        RECT 244.230 973.760 244.510 974.040 ;
        RECT 244.990 973.760 245.270 974.040 ;
        RECT 243.470 973.000 243.750 973.280 ;
        RECT 244.230 973.000 244.510 973.280 ;
        RECT 244.990 973.000 245.270 973.280 ;
        RECT 243.470 972.240 243.750 972.520 ;
        RECT 244.230 972.240 244.510 972.520 ;
        RECT 244.990 972.240 245.270 972.520 ;
        RECT 243.470 971.480 243.750 971.760 ;
        RECT 244.230 971.480 244.510 971.760 ;
        RECT 244.990 971.480 245.270 971.760 ;
        RECT 243.470 970.720 243.750 971.000 ;
        RECT 244.230 970.720 244.510 971.000 ;
        RECT 244.990 970.720 245.270 971.000 ;
        RECT 243.470 969.960 243.750 970.240 ;
        RECT 244.230 969.960 244.510 970.240 ;
        RECT 244.990 969.960 245.270 970.240 ;
        RECT 282.770 973.760 283.050 974.040 ;
        RECT 283.530 973.760 283.810 974.040 ;
        RECT 284.290 973.760 284.570 974.040 ;
        RECT 282.770 973.000 283.050 973.280 ;
        RECT 283.530 973.000 283.810 973.280 ;
        RECT 284.290 973.000 284.570 973.280 ;
        RECT 282.770 972.240 283.050 972.520 ;
        RECT 283.530 972.240 283.810 972.520 ;
        RECT 284.290 972.240 284.570 972.520 ;
        RECT 282.770 971.480 283.050 971.760 ;
        RECT 283.530 971.480 283.810 971.760 ;
        RECT 284.290 971.480 284.570 971.760 ;
        RECT 282.770 970.720 283.050 971.000 ;
        RECT 283.530 970.720 283.810 971.000 ;
        RECT 284.290 970.720 284.570 971.000 ;
        RECT 282.770 969.960 283.050 970.240 ;
        RECT 283.530 969.960 283.810 970.240 ;
        RECT 284.290 969.960 284.570 970.240 ;
        RECT 318.470 973.760 318.750 974.040 ;
        RECT 319.230 973.760 319.510 974.040 ;
        RECT 319.990 973.760 320.270 974.040 ;
        RECT 318.470 973.000 318.750 973.280 ;
        RECT 319.230 973.000 319.510 973.280 ;
        RECT 319.990 973.000 320.270 973.280 ;
        RECT 318.470 972.240 318.750 972.520 ;
        RECT 319.230 972.240 319.510 972.520 ;
        RECT 319.990 972.240 320.270 972.520 ;
        RECT 318.470 971.480 318.750 971.760 ;
        RECT 319.230 971.480 319.510 971.760 ;
        RECT 319.990 971.480 320.270 971.760 ;
        RECT 318.470 970.720 318.750 971.000 ;
        RECT 319.230 970.720 319.510 971.000 ;
        RECT 319.990 970.720 320.270 971.000 ;
        RECT 318.470 969.960 318.750 970.240 ;
        RECT 319.230 969.960 319.510 970.240 ;
        RECT 319.990 969.960 320.270 970.240 ;
        RECT 357.770 973.760 358.050 974.040 ;
        RECT 358.530 973.760 358.810 974.040 ;
        RECT 359.290 973.760 359.570 974.040 ;
        RECT 357.770 973.000 358.050 973.280 ;
        RECT 358.530 973.000 358.810 973.280 ;
        RECT 359.290 973.000 359.570 973.280 ;
        RECT 357.770 972.240 358.050 972.520 ;
        RECT 358.530 972.240 358.810 972.520 ;
        RECT 359.290 972.240 359.570 972.520 ;
        RECT 357.770 971.480 358.050 971.760 ;
        RECT 358.530 971.480 358.810 971.760 ;
        RECT 359.290 971.480 359.570 971.760 ;
        RECT 357.770 970.720 358.050 971.000 ;
        RECT 358.530 970.720 358.810 971.000 ;
        RECT 359.290 970.720 359.570 971.000 ;
        RECT 357.770 969.960 358.050 970.240 ;
        RECT 358.530 969.960 358.810 970.240 ;
        RECT 359.290 969.960 359.570 970.240 ;
        RECT 393.470 973.760 393.750 974.040 ;
        RECT 394.230 973.760 394.510 974.040 ;
        RECT 394.990 973.760 395.270 974.040 ;
        RECT 393.470 973.000 393.750 973.280 ;
        RECT 394.230 973.000 394.510 973.280 ;
        RECT 394.990 973.000 395.270 973.280 ;
        RECT 393.470 972.240 393.750 972.520 ;
        RECT 394.230 972.240 394.510 972.520 ;
        RECT 394.990 972.240 395.270 972.520 ;
        RECT 393.470 971.480 393.750 971.760 ;
        RECT 394.230 971.480 394.510 971.760 ;
        RECT 394.990 971.480 395.270 971.760 ;
        RECT 393.470 970.720 393.750 971.000 ;
        RECT 394.230 970.720 394.510 971.000 ;
        RECT 394.990 970.720 395.270 971.000 ;
        RECT 393.470 969.960 393.750 970.240 ;
        RECT 394.230 969.960 394.510 970.240 ;
        RECT 394.990 969.960 395.270 970.240 ;
        RECT 432.770 973.760 433.050 974.040 ;
        RECT 433.530 973.760 433.810 974.040 ;
        RECT 434.290 973.760 434.570 974.040 ;
        RECT 432.770 973.000 433.050 973.280 ;
        RECT 433.530 973.000 433.810 973.280 ;
        RECT 434.290 973.000 434.570 973.280 ;
        RECT 432.770 972.240 433.050 972.520 ;
        RECT 433.530 972.240 433.810 972.520 ;
        RECT 434.290 972.240 434.570 972.520 ;
        RECT 432.770 971.480 433.050 971.760 ;
        RECT 433.530 971.480 433.810 971.760 ;
        RECT 434.290 971.480 434.570 971.760 ;
        RECT 432.770 970.720 433.050 971.000 ;
        RECT 433.530 970.720 433.810 971.000 ;
        RECT 434.290 970.720 434.570 971.000 ;
        RECT 432.770 969.960 433.050 970.240 ;
        RECT 433.530 969.960 433.810 970.240 ;
        RECT 434.290 969.960 434.570 970.240 ;
        RECT 468.470 973.760 468.750 974.040 ;
        RECT 469.230 973.760 469.510 974.040 ;
        RECT 469.990 973.760 470.270 974.040 ;
        RECT 468.470 973.000 468.750 973.280 ;
        RECT 469.230 973.000 469.510 973.280 ;
        RECT 469.990 973.000 470.270 973.280 ;
        RECT 468.470 972.240 468.750 972.520 ;
        RECT 469.230 972.240 469.510 972.520 ;
        RECT 469.990 972.240 470.270 972.520 ;
        RECT 468.470 971.480 468.750 971.760 ;
        RECT 469.230 971.480 469.510 971.760 ;
        RECT 469.990 971.480 470.270 971.760 ;
        RECT 468.470 970.720 468.750 971.000 ;
        RECT 469.230 970.720 469.510 971.000 ;
        RECT 469.990 970.720 470.270 971.000 ;
        RECT 468.470 969.960 468.750 970.240 ;
        RECT 469.230 969.960 469.510 970.240 ;
        RECT 469.990 969.960 470.270 970.240 ;
        RECT 507.770 973.760 508.050 974.040 ;
        RECT 508.530 973.760 508.810 974.040 ;
        RECT 509.290 973.760 509.570 974.040 ;
        RECT 507.770 973.000 508.050 973.280 ;
        RECT 508.530 973.000 508.810 973.280 ;
        RECT 509.290 973.000 509.570 973.280 ;
        RECT 507.770 972.240 508.050 972.520 ;
        RECT 508.530 972.240 508.810 972.520 ;
        RECT 509.290 972.240 509.570 972.520 ;
        RECT 507.770 971.480 508.050 971.760 ;
        RECT 508.530 971.480 508.810 971.760 ;
        RECT 509.290 971.480 509.570 971.760 ;
        RECT 507.770 970.720 508.050 971.000 ;
        RECT 508.530 970.720 508.810 971.000 ;
        RECT 509.290 970.720 509.570 971.000 ;
        RECT 507.770 969.960 508.050 970.240 ;
        RECT 508.530 969.960 508.810 970.240 ;
        RECT 509.290 969.960 509.570 970.240 ;
        RECT 543.470 973.760 543.750 974.040 ;
        RECT 544.230 973.760 544.510 974.040 ;
        RECT 544.990 973.760 545.270 974.040 ;
        RECT 543.470 973.000 543.750 973.280 ;
        RECT 544.230 973.000 544.510 973.280 ;
        RECT 544.990 973.000 545.270 973.280 ;
        RECT 543.470 972.240 543.750 972.520 ;
        RECT 544.230 972.240 544.510 972.520 ;
        RECT 544.990 972.240 545.270 972.520 ;
        RECT 543.470 971.480 543.750 971.760 ;
        RECT 544.230 971.480 544.510 971.760 ;
        RECT 544.990 971.480 545.270 971.760 ;
        RECT 543.470 970.720 543.750 971.000 ;
        RECT 544.230 970.720 544.510 971.000 ;
        RECT 544.990 970.720 545.270 971.000 ;
        RECT 543.470 969.960 543.750 970.240 ;
        RECT 544.230 969.960 544.510 970.240 ;
        RECT 544.990 969.960 545.270 970.240 ;
        RECT -725.780 414.720 -724.980 435.280 ;
        RECT -724.580 414.720 -723.780 435.280 ;
        RECT -723.380 414.720 -722.580 435.280 ;
        RECT -722.180 414.720 -721.380 435.280 ;
        RECT -720.980 414.720 -720.180 435.280 ;
        RECT -719.780 414.720 -718.980 435.280 ;
        RECT -718.580 414.720 -717.780 435.280 ;
        RECT -717.380 414.720 -716.580 435.280 ;
        RECT -716.180 414.720 -715.380 435.280 ;
        RECT -714.980 414.720 -714.180 435.280 ;
        RECT -713.780 414.720 -712.980 435.280 ;
        RECT -712.580 414.720 -711.780 435.280 ;
        RECT -711.380 414.720 -710.580 435.280 ;
        RECT -710.180 414.720 -709.380 435.280 ;
        RECT -708.980 414.720 -708.180 435.280 ;
        RECT -707.780 414.720 -706.980 435.280 ;
        RECT -706.580 414.720 -705.780 435.280 ;
        RECT -705.380 414.720 -704.580 435.280 ;
        RECT -704.180 414.720 -703.380 435.280 ;
        RECT -702.980 414.720 -702.180 435.280 ;
        RECT -701.780 414.720 -700.980 435.280 ;
        RECT -700.580 414.720 -699.780 435.280 ;
        RECT -699.380 414.720 -698.580 435.280 ;
        RECT -698.180 414.720 -697.380 435.280 ;
        RECT -696.980 414.720 -696.180 435.280 ;
        RECT -695.780 414.720 -694.980 435.280 ;
        RECT -694.580 414.720 -693.780 435.280 ;
        RECT -693.380 414.720 -692.580 435.280 ;
        RECT -692.180 414.720 -691.380 435.280 ;
        RECT -690.980 414.720 -690.180 435.280 ;
        RECT -689.780 414.720 -688.980 435.280 ;
        RECT -688.580 414.720 -687.780 435.280 ;
        RECT -687.380 414.720 -686.580 435.280 ;
        RECT -686.180 414.720 -685.380 435.280 ;
        RECT -684.980 414.720 -684.180 435.280 ;
        RECT -683.780 414.720 -682.980 435.280 ;
        RECT -682.580 414.720 -681.780 435.280 ;
        RECT -681.380 414.720 -680.580 435.280 ;
        RECT -680.180 414.720 -679.380 435.280 ;
        RECT -678.980 414.720 -678.180 435.280 ;
        RECT -677.780 414.720 -676.980 435.280 ;
        RECT -676.580 414.720 -675.780 435.280 ;
        RECT -675.380 414.720 -674.580 435.280 ;
        RECT -674.180 414.720 -673.380 435.280 ;
        RECT -672.980 414.720 -672.180 435.280 ;
        RECT -671.780 414.720 -670.980 435.280 ;
        RECT -670.580 414.720 -669.780 435.280 ;
        RECT -669.380 414.720 -668.580 435.280 ;
        RECT -668.180 414.720 -667.380 435.280 ;
        RECT -666.980 414.720 -666.180 435.280 ;
        RECT -665.780 414.720 -664.980 435.280 ;
        RECT -664.580 414.720 -663.780 435.280 ;
        RECT -663.380 414.720 -662.580 435.280 ;
        RECT -662.180 414.720 -661.380 435.280 ;
        RECT -660.980 414.720 -660.180 435.280 ;
        RECT -659.780 414.720 -658.980 435.280 ;
        RECT -658.580 414.720 -657.780 435.280 ;
        RECT -657.380 414.720 -656.580 435.280 ;
        RECT -656.180 414.720 -655.380 435.280 ;
        RECT -654.980 414.720 -654.180 435.280 ;
        RECT -653.780 414.720 -652.980 435.280 ;
        RECT -652.580 414.720 -651.780 435.280 ;
        RECT 654.820 414.720 655.620 435.280 ;
        RECT 656.020 414.720 656.820 435.280 ;
        RECT 657.220 414.720 658.020 435.280 ;
        RECT 658.420 414.720 659.220 435.280 ;
        RECT 659.620 414.720 660.420 435.280 ;
        RECT 660.820 414.720 661.620 435.280 ;
        RECT 662.020 414.720 662.820 435.280 ;
        RECT 663.220 414.720 664.020 435.280 ;
        RECT 664.420 414.720 665.220 435.280 ;
        RECT 665.620 414.720 666.420 435.280 ;
        RECT 666.820 414.720 667.620 435.280 ;
        RECT 668.020 414.720 668.820 435.280 ;
        RECT 669.220 414.720 670.020 435.280 ;
        RECT 670.420 414.720 671.220 435.280 ;
        RECT 671.620 414.720 672.420 435.280 ;
        RECT 672.820 414.720 673.620 435.280 ;
        RECT 674.020 414.720 674.820 435.280 ;
        RECT 675.220 414.720 676.020 435.280 ;
        RECT 676.420 414.720 677.220 435.280 ;
        RECT 677.620 414.720 678.420 435.280 ;
        RECT 678.820 414.720 679.620 435.280 ;
        RECT 680.020 414.720 680.820 435.280 ;
        RECT 681.220 414.720 682.020 435.280 ;
        RECT 682.420 414.720 683.220 435.280 ;
        RECT 683.620 414.720 684.420 435.280 ;
        RECT 684.820 414.720 685.620 435.280 ;
        RECT 686.020 414.720 686.820 435.280 ;
        RECT 687.220 414.720 688.020 435.280 ;
        RECT 688.420 414.720 689.220 435.280 ;
        RECT 689.620 414.720 690.420 435.280 ;
        RECT 690.820 414.720 691.620 435.280 ;
        RECT 692.020 414.720 692.820 435.280 ;
        RECT 693.220 414.720 694.020 435.280 ;
        RECT 694.420 414.720 695.220 435.280 ;
        RECT 695.620 414.720 696.420 435.280 ;
        RECT 696.820 414.720 697.620 435.280 ;
        RECT 698.020 414.720 698.820 435.280 ;
        RECT 699.220 414.720 700.020 435.280 ;
        RECT 700.420 414.720 701.220 435.280 ;
        RECT 701.620 414.720 702.420 435.280 ;
        RECT 702.820 414.720 703.620 435.280 ;
        RECT 704.020 414.720 704.820 435.280 ;
        RECT 705.220 414.720 706.020 435.280 ;
        RECT 706.420 414.720 707.220 435.280 ;
        RECT 707.620 414.720 708.420 435.280 ;
        RECT 708.820 414.720 709.620 435.280 ;
        RECT 710.020 414.720 710.820 435.280 ;
        RECT 711.220 414.720 712.020 435.280 ;
        RECT 712.420 414.720 713.220 435.280 ;
        RECT 713.620 414.720 714.420 435.280 ;
        RECT 714.820 414.720 715.620 435.280 ;
        RECT 716.020 414.720 716.820 435.280 ;
        RECT 717.220 414.720 718.020 435.280 ;
        RECT 718.420 414.720 719.220 435.280 ;
        RECT 719.620 414.720 720.420 435.280 ;
        RECT 720.820 414.720 721.620 435.280 ;
        RECT 722.020 414.720 722.820 435.280 ;
        RECT 723.220 414.720 724.020 435.280 ;
        RECT 724.420 414.720 725.220 435.280 ;
        RECT 725.620 414.720 726.420 435.280 ;
        RECT 726.820 414.720 727.620 435.280 ;
        RECT 728.020 414.720 728.820 435.280 ;
        RECT -485.930 122.130 -485.650 122.410 ;
        RECT -485.310 122.130 -485.030 122.410 ;
        RECT -484.690 122.130 -484.410 122.410 ;
        RECT -484.070 122.130 -483.790 122.410 ;
        RECT -483.450 122.130 -483.170 122.410 ;
        RECT -482.830 122.130 -482.550 122.410 ;
        RECT -482.210 122.130 -481.930 122.410 ;
        RECT -481.590 122.130 -481.310 122.410 ;
        RECT -480.970 122.130 -480.690 122.410 ;
        RECT -480.350 122.130 -480.070 122.410 ;
        RECT -485.930 121.510 -485.650 121.790 ;
        RECT -485.310 121.510 -485.030 121.790 ;
        RECT -484.690 121.510 -484.410 121.790 ;
        RECT -484.070 121.510 -483.790 121.790 ;
        RECT -483.450 121.510 -483.170 121.790 ;
        RECT -482.830 121.510 -482.550 121.790 ;
        RECT -482.210 121.510 -481.930 121.790 ;
        RECT -481.590 121.510 -481.310 121.790 ;
        RECT -480.970 121.510 -480.690 121.790 ;
        RECT -480.350 121.510 -480.070 121.790 ;
        RECT -485.930 120.890 -485.650 121.170 ;
        RECT -485.310 120.890 -485.030 121.170 ;
        RECT -484.690 120.890 -484.410 121.170 ;
        RECT -484.070 120.890 -483.790 121.170 ;
        RECT -483.450 120.890 -483.170 121.170 ;
        RECT -482.830 120.890 -482.550 121.170 ;
        RECT -482.210 120.890 -481.930 121.170 ;
        RECT -481.590 120.890 -481.310 121.170 ;
        RECT -480.970 120.890 -480.690 121.170 ;
        RECT -480.350 120.890 -480.070 121.170 ;
        RECT -485.930 120.270 -485.650 120.550 ;
        RECT -485.310 120.270 -485.030 120.550 ;
        RECT -484.690 120.270 -484.410 120.550 ;
        RECT -484.070 120.270 -483.790 120.550 ;
        RECT -483.450 120.270 -483.170 120.550 ;
        RECT -482.830 120.270 -482.550 120.550 ;
        RECT -482.210 120.270 -481.930 120.550 ;
        RECT -481.590 120.270 -481.310 120.550 ;
        RECT -480.970 120.270 -480.690 120.550 ;
        RECT -480.350 120.270 -480.070 120.550 ;
        RECT -485.930 119.650 -485.650 119.930 ;
        RECT -485.310 119.650 -485.030 119.930 ;
        RECT -484.690 119.650 -484.410 119.930 ;
        RECT -484.070 119.650 -483.790 119.930 ;
        RECT -483.450 119.650 -483.170 119.930 ;
        RECT -482.830 119.650 -482.550 119.930 ;
        RECT -482.210 119.650 -481.930 119.930 ;
        RECT -481.590 119.650 -481.310 119.930 ;
        RECT -480.970 119.650 -480.690 119.930 ;
        RECT -480.350 119.650 -480.070 119.930 ;
        RECT -485.930 119.030 -485.650 119.310 ;
        RECT -485.310 119.030 -485.030 119.310 ;
        RECT -484.690 119.030 -484.410 119.310 ;
        RECT -484.070 119.030 -483.790 119.310 ;
        RECT -483.450 119.030 -483.170 119.310 ;
        RECT -482.830 119.030 -482.550 119.310 ;
        RECT -482.210 119.030 -481.930 119.310 ;
        RECT -481.590 119.030 -481.310 119.310 ;
        RECT -480.970 119.030 -480.690 119.310 ;
        RECT -480.350 119.030 -480.070 119.310 ;
        RECT -485.930 118.410 -485.650 118.690 ;
        RECT -485.310 118.410 -485.030 118.690 ;
        RECT -484.690 118.410 -484.410 118.690 ;
        RECT -484.070 118.410 -483.790 118.690 ;
        RECT -483.450 118.410 -483.170 118.690 ;
        RECT -482.830 118.410 -482.550 118.690 ;
        RECT -482.210 118.410 -481.930 118.690 ;
        RECT -481.590 118.410 -481.310 118.690 ;
        RECT -480.970 118.410 -480.690 118.690 ;
        RECT -480.350 118.410 -480.070 118.690 ;
        RECT -485.930 117.790 -485.650 118.070 ;
        RECT -485.310 117.790 -485.030 118.070 ;
        RECT -484.690 117.790 -484.410 118.070 ;
        RECT -484.070 117.790 -483.790 118.070 ;
        RECT -483.450 117.790 -483.170 118.070 ;
        RECT -482.830 117.790 -482.550 118.070 ;
        RECT -482.210 117.790 -481.930 118.070 ;
        RECT -481.590 117.790 -481.310 118.070 ;
        RECT -480.970 117.790 -480.690 118.070 ;
        RECT -480.350 117.790 -480.070 118.070 ;
        RECT 142.315 122.130 142.595 122.410 ;
        RECT 142.935 122.130 143.215 122.410 ;
        RECT 142.315 121.510 142.595 121.790 ;
        RECT 142.935 121.510 143.215 121.790 ;
        RECT 142.315 120.890 142.595 121.170 ;
        RECT 142.935 120.890 143.215 121.170 ;
        RECT 142.315 120.270 142.595 120.550 ;
        RECT 142.935 120.270 143.215 120.550 ;
        RECT 142.315 119.650 142.595 119.930 ;
        RECT 142.935 119.650 143.215 119.930 ;
        RECT 142.315 119.030 142.595 119.310 ;
        RECT 142.935 119.030 143.215 119.310 ;
        RECT 142.315 118.410 142.595 118.690 ;
        RECT 142.935 118.410 143.215 118.690 ;
        RECT 142.315 117.790 142.595 118.070 ;
        RECT 142.935 117.790 143.215 118.070 ;
        RECT 164.890 122.130 165.170 122.410 ;
        RECT 165.510 122.130 165.790 122.410 ;
        RECT 166.130 122.130 166.410 122.410 ;
        RECT 166.750 122.130 167.030 122.410 ;
        RECT 167.370 122.130 167.650 122.410 ;
        RECT 167.990 122.130 168.270 122.410 ;
        RECT 168.610 122.130 168.890 122.410 ;
        RECT 169.230 122.130 169.510 122.410 ;
        RECT 169.850 122.130 170.130 122.410 ;
        RECT 170.470 122.130 170.750 122.410 ;
        RECT 164.890 121.510 165.170 121.790 ;
        RECT 165.510 121.510 165.790 121.790 ;
        RECT 166.130 121.510 166.410 121.790 ;
        RECT 166.750 121.510 167.030 121.790 ;
        RECT 167.370 121.510 167.650 121.790 ;
        RECT 167.990 121.510 168.270 121.790 ;
        RECT 168.610 121.510 168.890 121.790 ;
        RECT 169.230 121.510 169.510 121.790 ;
        RECT 169.850 121.510 170.130 121.790 ;
        RECT 170.470 121.510 170.750 121.790 ;
        RECT 164.890 120.890 165.170 121.170 ;
        RECT 165.510 120.890 165.790 121.170 ;
        RECT 166.130 120.890 166.410 121.170 ;
        RECT 166.750 120.890 167.030 121.170 ;
        RECT 167.370 120.890 167.650 121.170 ;
        RECT 167.990 120.890 168.270 121.170 ;
        RECT 168.610 120.890 168.890 121.170 ;
        RECT 169.230 120.890 169.510 121.170 ;
        RECT 169.850 120.890 170.130 121.170 ;
        RECT 170.470 120.890 170.750 121.170 ;
        RECT 164.890 120.270 165.170 120.550 ;
        RECT 165.510 120.270 165.790 120.550 ;
        RECT 166.130 120.270 166.410 120.550 ;
        RECT 166.750 120.270 167.030 120.550 ;
        RECT 167.370 120.270 167.650 120.550 ;
        RECT 167.990 120.270 168.270 120.550 ;
        RECT 168.610 120.270 168.890 120.550 ;
        RECT 169.230 120.270 169.510 120.550 ;
        RECT 169.850 120.270 170.130 120.550 ;
        RECT 170.470 120.270 170.750 120.550 ;
        RECT 164.890 119.650 165.170 119.930 ;
        RECT 165.510 119.650 165.790 119.930 ;
        RECT 166.130 119.650 166.410 119.930 ;
        RECT 166.750 119.650 167.030 119.930 ;
        RECT 167.370 119.650 167.650 119.930 ;
        RECT 167.990 119.650 168.270 119.930 ;
        RECT 168.610 119.650 168.890 119.930 ;
        RECT 169.230 119.650 169.510 119.930 ;
        RECT 169.850 119.650 170.130 119.930 ;
        RECT 170.470 119.650 170.750 119.930 ;
        RECT 164.890 119.030 165.170 119.310 ;
        RECT 165.510 119.030 165.790 119.310 ;
        RECT 166.130 119.030 166.410 119.310 ;
        RECT 166.750 119.030 167.030 119.310 ;
        RECT 167.370 119.030 167.650 119.310 ;
        RECT 167.990 119.030 168.270 119.310 ;
        RECT 168.610 119.030 168.890 119.310 ;
        RECT 169.230 119.030 169.510 119.310 ;
        RECT 169.850 119.030 170.130 119.310 ;
        RECT 170.470 119.030 170.750 119.310 ;
        RECT 164.890 118.410 165.170 118.690 ;
        RECT 165.510 118.410 165.790 118.690 ;
        RECT 166.130 118.410 166.410 118.690 ;
        RECT 166.750 118.410 167.030 118.690 ;
        RECT 167.370 118.410 167.650 118.690 ;
        RECT 167.990 118.410 168.270 118.690 ;
        RECT 168.610 118.410 168.890 118.690 ;
        RECT 169.230 118.410 169.510 118.690 ;
        RECT 169.850 118.410 170.130 118.690 ;
        RECT 170.470 118.410 170.750 118.690 ;
        RECT 164.890 117.790 165.170 118.070 ;
        RECT 165.510 117.790 165.790 118.070 ;
        RECT 166.130 117.790 166.410 118.070 ;
        RECT 166.750 117.790 167.030 118.070 ;
        RECT 167.370 117.790 167.650 118.070 ;
        RECT 167.990 117.790 168.270 118.070 ;
        RECT 168.610 117.790 168.890 118.070 ;
        RECT 169.230 117.790 169.510 118.070 ;
        RECT 169.850 117.790 170.130 118.070 ;
        RECT 170.470 117.790 170.750 118.070 ;
        RECT 316.050 117.940 317.370 120.300 ;
        RECT -485.930 -118.070 -485.650 -117.790 ;
        RECT -485.310 -118.070 -485.030 -117.790 ;
        RECT -484.690 -118.070 -484.410 -117.790 ;
        RECT -484.070 -118.070 -483.790 -117.790 ;
        RECT -483.450 -118.070 -483.170 -117.790 ;
        RECT -482.830 -118.070 -482.550 -117.790 ;
        RECT -482.210 -118.070 -481.930 -117.790 ;
        RECT -481.590 -118.070 -481.310 -117.790 ;
        RECT -480.970 -118.070 -480.690 -117.790 ;
        RECT -480.350 -118.070 -480.070 -117.790 ;
        RECT -485.930 -118.690 -485.650 -118.410 ;
        RECT -485.310 -118.690 -485.030 -118.410 ;
        RECT -484.690 -118.690 -484.410 -118.410 ;
        RECT -484.070 -118.690 -483.790 -118.410 ;
        RECT -483.450 -118.690 -483.170 -118.410 ;
        RECT -482.830 -118.690 -482.550 -118.410 ;
        RECT -482.210 -118.690 -481.930 -118.410 ;
        RECT -481.590 -118.690 -481.310 -118.410 ;
        RECT -480.970 -118.690 -480.690 -118.410 ;
        RECT -480.350 -118.690 -480.070 -118.410 ;
        RECT -485.930 -119.310 -485.650 -119.030 ;
        RECT -485.310 -119.310 -485.030 -119.030 ;
        RECT -484.690 -119.310 -484.410 -119.030 ;
        RECT -484.070 -119.310 -483.790 -119.030 ;
        RECT -483.450 -119.310 -483.170 -119.030 ;
        RECT -482.830 -119.310 -482.550 -119.030 ;
        RECT -482.210 -119.310 -481.930 -119.030 ;
        RECT -481.590 -119.310 -481.310 -119.030 ;
        RECT -480.970 -119.310 -480.690 -119.030 ;
        RECT -480.350 -119.310 -480.070 -119.030 ;
        RECT -485.930 -119.930 -485.650 -119.650 ;
        RECT -485.310 -119.930 -485.030 -119.650 ;
        RECT -484.690 -119.930 -484.410 -119.650 ;
        RECT -484.070 -119.930 -483.790 -119.650 ;
        RECT -483.450 -119.930 -483.170 -119.650 ;
        RECT -482.830 -119.930 -482.550 -119.650 ;
        RECT -482.210 -119.930 -481.930 -119.650 ;
        RECT -481.590 -119.930 -481.310 -119.650 ;
        RECT -480.970 -119.930 -480.690 -119.650 ;
        RECT -480.350 -119.930 -480.070 -119.650 ;
        RECT -485.930 -120.550 -485.650 -120.270 ;
        RECT -485.310 -120.550 -485.030 -120.270 ;
        RECT -484.690 -120.550 -484.410 -120.270 ;
        RECT -484.070 -120.550 -483.790 -120.270 ;
        RECT -483.450 -120.550 -483.170 -120.270 ;
        RECT -482.830 -120.550 -482.550 -120.270 ;
        RECT -482.210 -120.550 -481.930 -120.270 ;
        RECT -481.590 -120.550 -481.310 -120.270 ;
        RECT -480.970 -120.550 -480.690 -120.270 ;
        RECT -480.350 -120.550 -480.070 -120.270 ;
        RECT -485.930 -121.170 -485.650 -120.890 ;
        RECT -485.310 -121.170 -485.030 -120.890 ;
        RECT -484.690 -121.170 -484.410 -120.890 ;
        RECT -484.070 -121.170 -483.790 -120.890 ;
        RECT -483.450 -121.170 -483.170 -120.890 ;
        RECT -482.830 -121.170 -482.550 -120.890 ;
        RECT -482.210 -121.170 -481.930 -120.890 ;
        RECT -481.590 -121.170 -481.310 -120.890 ;
        RECT -480.970 -121.170 -480.690 -120.890 ;
        RECT -480.350 -121.170 -480.070 -120.890 ;
        RECT -485.930 -121.790 -485.650 -121.510 ;
        RECT -485.310 -121.790 -485.030 -121.510 ;
        RECT -484.690 -121.790 -484.410 -121.510 ;
        RECT -484.070 -121.790 -483.790 -121.510 ;
        RECT -483.450 -121.790 -483.170 -121.510 ;
        RECT -482.830 -121.790 -482.550 -121.510 ;
        RECT -482.210 -121.790 -481.930 -121.510 ;
        RECT -481.590 -121.790 -481.310 -121.510 ;
        RECT -480.970 -121.790 -480.690 -121.510 ;
        RECT -480.350 -121.790 -480.070 -121.510 ;
        RECT -485.930 -122.410 -485.650 -122.130 ;
        RECT -485.310 -122.410 -485.030 -122.130 ;
        RECT -484.690 -122.410 -484.410 -122.130 ;
        RECT -484.070 -122.410 -483.790 -122.130 ;
        RECT -483.450 -122.410 -483.170 -122.130 ;
        RECT -482.830 -122.410 -482.550 -122.130 ;
        RECT -482.210 -122.410 -481.930 -122.130 ;
        RECT -481.590 -122.410 -481.310 -122.130 ;
        RECT -480.970 -122.410 -480.690 -122.130 ;
        RECT -480.350 -122.410 -480.070 -122.130 ;
        RECT 142.315 -118.070 142.595 -117.790 ;
        RECT 142.935 -118.070 143.215 -117.790 ;
        RECT 142.315 -118.690 142.595 -118.410 ;
        RECT 142.935 -118.690 143.215 -118.410 ;
        RECT 142.315 -119.310 142.595 -119.030 ;
        RECT 142.935 -119.310 143.215 -119.030 ;
        RECT 142.315 -119.930 142.595 -119.650 ;
        RECT 142.935 -119.930 143.215 -119.650 ;
        RECT 142.315 -120.550 142.595 -120.270 ;
        RECT 142.935 -120.550 143.215 -120.270 ;
        RECT 142.315 -121.170 142.595 -120.890 ;
        RECT 142.935 -121.170 143.215 -120.890 ;
        RECT 142.315 -121.790 142.595 -121.510 ;
        RECT 142.935 -121.790 143.215 -121.510 ;
        RECT 142.315 -122.410 142.595 -122.130 ;
        RECT 142.935 -122.410 143.215 -122.130 ;
        RECT 164.890 -118.070 165.170 -117.790 ;
        RECT 165.510 -118.070 165.790 -117.790 ;
        RECT 166.130 -118.070 166.410 -117.790 ;
        RECT 166.750 -118.070 167.030 -117.790 ;
        RECT 167.370 -118.070 167.650 -117.790 ;
        RECT 167.990 -118.070 168.270 -117.790 ;
        RECT 168.610 -118.070 168.890 -117.790 ;
        RECT 169.230 -118.070 169.510 -117.790 ;
        RECT 169.850 -118.070 170.130 -117.790 ;
        RECT 170.470 -118.070 170.750 -117.790 ;
        RECT 164.890 -118.690 165.170 -118.410 ;
        RECT 165.510 -118.690 165.790 -118.410 ;
        RECT 166.130 -118.690 166.410 -118.410 ;
        RECT 166.750 -118.690 167.030 -118.410 ;
        RECT 167.370 -118.690 167.650 -118.410 ;
        RECT 167.990 -118.690 168.270 -118.410 ;
        RECT 168.610 -118.690 168.890 -118.410 ;
        RECT 169.230 -118.690 169.510 -118.410 ;
        RECT 169.850 -118.690 170.130 -118.410 ;
        RECT 170.470 -118.690 170.750 -118.410 ;
        RECT 164.890 -119.310 165.170 -119.030 ;
        RECT 165.510 -119.310 165.790 -119.030 ;
        RECT 166.130 -119.310 166.410 -119.030 ;
        RECT 166.750 -119.310 167.030 -119.030 ;
        RECT 167.370 -119.310 167.650 -119.030 ;
        RECT 167.990 -119.310 168.270 -119.030 ;
        RECT 168.610 -119.310 168.890 -119.030 ;
        RECT 169.230 -119.310 169.510 -119.030 ;
        RECT 169.850 -119.310 170.130 -119.030 ;
        RECT 170.470 -119.310 170.750 -119.030 ;
        RECT 164.890 -119.930 165.170 -119.650 ;
        RECT 165.510 -119.930 165.790 -119.650 ;
        RECT 166.130 -119.930 166.410 -119.650 ;
        RECT 166.750 -119.930 167.030 -119.650 ;
        RECT 167.370 -119.930 167.650 -119.650 ;
        RECT 167.990 -119.930 168.270 -119.650 ;
        RECT 168.610 -119.930 168.890 -119.650 ;
        RECT 169.230 -119.930 169.510 -119.650 ;
        RECT 169.850 -119.930 170.130 -119.650 ;
        RECT 170.470 -119.930 170.750 -119.650 ;
        RECT 164.890 -120.550 165.170 -120.270 ;
        RECT 165.510 -120.550 165.790 -120.270 ;
        RECT 166.130 -120.550 166.410 -120.270 ;
        RECT 166.750 -120.550 167.030 -120.270 ;
        RECT 167.370 -120.550 167.650 -120.270 ;
        RECT 167.990 -120.550 168.270 -120.270 ;
        RECT 168.610 -120.550 168.890 -120.270 ;
        RECT 169.230 -120.550 169.510 -120.270 ;
        RECT 169.850 -120.550 170.130 -120.270 ;
        RECT 170.470 -120.550 170.750 -120.270 ;
        RECT 164.890 -121.170 165.170 -120.890 ;
        RECT 165.510 -121.170 165.790 -120.890 ;
        RECT 166.130 -121.170 166.410 -120.890 ;
        RECT 166.750 -121.170 167.030 -120.890 ;
        RECT 167.370 -121.170 167.650 -120.890 ;
        RECT 167.990 -121.170 168.270 -120.890 ;
        RECT 168.610 -121.170 168.890 -120.890 ;
        RECT 169.230 -121.170 169.510 -120.890 ;
        RECT 169.850 -121.170 170.130 -120.890 ;
        RECT 170.470 -121.170 170.750 -120.890 ;
        RECT 316.050 -120.300 317.370 -117.940 ;
        RECT 357.630 117.940 358.950 120.300 ;
        RECT 357.630 -120.300 358.950 -117.940 ;
        RECT 399.210 117.940 400.530 120.300 ;
        RECT 399.210 -120.300 400.530 -117.940 ;
        RECT 440.790 117.940 442.110 120.300 ;
        RECT 440.790 -120.300 442.110 -117.940 ;
        RECT 164.890 -121.790 165.170 -121.510 ;
        RECT 165.510 -121.790 165.790 -121.510 ;
        RECT 166.130 -121.790 166.410 -121.510 ;
        RECT 166.750 -121.790 167.030 -121.510 ;
        RECT 167.370 -121.790 167.650 -121.510 ;
        RECT 167.990 -121.790 168.270 -121.510 ;
        RECT 168.610 -121.790 168.890 -121.510 ;
        RECT 169.230 -121.790 169.510 -121.510 ;
        RECT 169.850 -121.790 170.130 -121.510 ;
        RECT 170.470 -121.790 170.750 -121.510 ;
        RECT 164.890 -122.410 165.170 -122.130 ;
        RECT 165.510 -122.410 165.790 -122.130 ;
        RECT 166.130 -122.410 166.410 -122.130 ;
        RECT 166.750 -122.410 167.030 -122.130 ;
        RECT 167.370 -122.410 167.650 -122.130 ;
        RECT 167.990 -122.410 168.270 -122.130 ;
        RECT 168.610 -122.410 168.890 -122.130 ;
        RECT 169.230 -122.410 169.510 -122.130 ;
        RECT 169.850 -122.410 170.130 -122.130 ;
        RECT 170.470 -122.410 170.750 -122.130 ;
        RECT -725.780 -435.280 -724.980 -414.720 ;
        RECT -724.580 -435.280 -723.780 -414.720 ;
        RECT -723.380 -435.280 -722.580 -414.720 ;
        RECT -722.180 -435.280 -721.380 -414.720 ;
        RECT -720.980 -435.280 -720.180 -414.720 ;
        RECT -719.780 -435.280 -718.980 -414.720 ;
        RECT -718.580 -435.280 -717.780 -414.720 ;
        RECT -717.380 -435.280 -716.580 -414.720 ;
        RECT -716.180 -435.280 -715.380 -414.720 ;
        RECT -714.980 -435.280 -714.180 -414.720 ;
        RECT -713.780 -435.280 -712.980 -414.720 ;
        RECT -712.580 -435.280 -711.780 -414.720 ;
        RECT -711.380 -435.280 -710.580 -414.720 ;
        RECT -710.180 -435.280 -709.380 -414.720 ;
        RECT -708.980 -435.280 -708.180 -414.720 ;
        RECT -707.780 -435.280 -706.980 -414.720 ;
        RECT -706.580 -435.280 -705.780 -414.720 ;
        RECT -705.380 -435.280 -704.580 -414.720 ;
        RECT -704.180 -435.280 -703.380 -414.720 ;
        RECT -702.980 -435.280 -702.180 -414.720 ;
        RECT -701.780 -435.280 -700.980 -414.720 ;
        RECT -700.580 -435.280 -699.780 -414.720 ;
        RECT -699.380 -435.280 -698.580 -414.720 ;
        RECT -698.180 -435.280 -697.380 -414.720 ;
        RECT -696.980 -435.280 -696.180 -414.720 ;
        RECT -695.780 -435.280 -694.980 -414.720 ;
        RECT -694.580 -435.280 -693.780 -414.720 ;
        RECT -693.380 -435.280 -692.580 -414.720 ;
        RECT -692.180 -435.280 -691.380 -414.720 ;
        RECT -690.980 -435.280 -690.180 -414.720 ;
        RECT -689.780 -435.280 -688.980 -414.720 ;
        RECT -688.580 -435.280 -687.780 -414.720 ;
        RECT -687.380 -435.280 -686.580 -414.720 ;
        RECT -686.180 -435.280 -685.380 -414.720 ;
        RECT -684.980 -435.280 -684.180 -414.720 ;
        RECT -683.780 -435.280 -682.980 -414.720 ;
        RECT -682.580 -435.280 -681.780 -414.720 ;
        RECT -681.380 -435.280 -680.580 -414.720 ;
        RECT -680.180 -435.280 -679.380 -414.720 ;
        RECT -678.980 -435.280 -678.180 -414.720 ;
        RECT -677.780 -435.280 -676.980 -414.720 ;
        RECT -676.580 -435.280 -675.780 -414.720 ;
        RECT -675.380 -435.280 -674.580 -414.720 ;
        RECT -674.180 -435.280 -673.380 -414.720 ;
        RECT -672.980 -435.280 -672.180 -414.720 ;
        RECT -671.780 -435.280 -670.980 -414.720 ;
        RECT -670.580 -435.280 -669.780 -414.720 ;
        RECT -669.380 -435.280 -668.580 -414.720 ;
        RECT -668.180 -435.280 -667.380 -414.720 ;
        RECT -666.980 -435.280 -666.180 -414.720 ;
        RECT -665.780 -435.280 -664.980 -414.720 ;
        RECT -664.580 -435.280 -663.780 -414.720 ;
        RECT -663.380 -435.280 -662.580 -414.720 ;
        RECT -662.180 -435.280 -661.380 -414.720 ;
        RECT -660.980 -435.280 -660.180 -414.720 ;
        RECT -659.780 -435.280 -658.980 -414.720 ;
        RECT -658.580 -435.280 -657.780 -414.720 ;
        RECT -657.380 -435.280 -656.580 -414.720 ;
        RECT -656.180 -435.280 -655.380 -414.720 ;
        RECT -654.980 -435.280 -654.180 -414.720 ;
        RECT -653.780 -435.280 -652.980 -414.720 ;
        RECT -652.580 -435.280 -651.780 -414.720 ;
        RECT 654.820 -435.280 655.620 -414.720 ;
        RECT 656.020 -435.280 656.820 -414.720 ;
        RECT 657.220 -435.280 658.020 -414.720 ;
        RECT 658.420 -435.280 659.220 -414.720 ;
        RECT 659.620 -435.280 660.420 -414.720 ;
        RECT 660.820 -435.280 661.620 -414.720 ;
        RECT 662.020 -435.280 662.820 -414.720 ;
        RECT 663.220 -435.280 664.020 -414.720 ;
        RECT 664.420 -435.280 665.220 -414.720 ;
        RECT 665.620 -435.280 666.420 -414.720 ;
        RECT 666.820 -435.280 667.620 -414.720 ;
        RECT 668.020 -435.280 668.820 -414.720 ;
        RECT 669.220 -435.280 670.020 -414.720 ;
        RECT 670.420 -435.280 671.220 -414.720 ;
        RECT 671.620 -435.280 672.420 -414.720 ;
        RECT 672.820 -435.280 673.620 -414.720 ;
        RECT 674.020 -435.280 674.820 -414.720 ;
        RECT 675.220 -435.280 676.020 -414.720 ;
        RECT 676.420 -435.280 677.220 -414.720 ;
        RECT 677.620 -435.280 678.420 -414.720 ;
        RECT 678.820 -435.280 679.620 -414.720 ;
        RECT 680.020 -435.280 680.820 -414.720 ;
        RECT 681.220 -435.280 682.020 -414.720 ;
        RECT 682.420 -435.280 683.220 -414.720 ;
        RECT 683.620 -435.280 684.420 -414.720 ;
        RECT 684.820 -435.280 685.620 -414.720 ;
        RECT 686.020 -435.280 686.820 -414.720 ;
        RECT 687.220 -435.280 688.020 -414.720 ;
        RECT 688.420 -435.280 689.220 -414.720 ;
        RECT 689.620 -435.280 690.420 -414.720 ;
        RECT 690.820 -435.280 691.620 -414.720 ;
        RECT 692.020 -435.280 692.820 -414.720 ;
        RECT 693.220 -435.280 694.020 -414.720 ;
        RECT 694.420 -435.280 695.220 -414.720 ;
        RECT 695.620 -435.280 696.420 -414.720 ;
        RECT 696.820 -435.280 697.620 -414.720 ;
        RECT 698.020 -435.280 698.820 -414.720 ;
        RECT 699.220 -435.280 700.020 -414.720 ;
        RECT 700.420 -435.280 701.220 -414.720 ;
        RECT 701.620 -435.280 702.420 -414.720 ;
        RECT 702.820 -435.280 703.620 -414.720 ;
        RECT 704.020 -435.280 704.820 -414.720 ;
        RECT 705.220 -435.280 706.020 -414.720 ;
        RECT 706.420 -435.280 707.220 -414.720 ;
        RECT 707.620 -435.280 708.420 -414.720 ;
        RECT 708.820 -435.280 709.620 -414.720 ;
        RECT 710.020 -435.280 710.820 -414.720 ;
        RECT 711.220 -435.280 712.020 -414.720 ;
        RECT 712.420 -435.280 713.220 -414.720 ;
        RECT 713.620 -435.280 714.420 -414.720 ;
        RECT 714.820 -435.280 715.620 -414.720 ;
        RECT 716.020 -435.280 716.820 -414.720 ;
        RECT 717.220 -435.280 718.020 -414.720 ;
        RECT 718.420 -435.280 719.220 -414.720 ;
        RECT 719.620 -435.280 720.420 -414.720 ;
        RECT 720.820 -435.280 721.620 -414.720 ;
        RECT 722.020 -435.280 722.820 -414.720 ;
        RECT 723.220 -435.280 724.020 -414.720 ;
        RECT 724.420 -435.280 725.220 -414.720 ;
        RECT 725.620 -435.280 726.420 -414.720 ;
        RECT 726.820 -435.280 727.620 -414.720 ;
        RECT 728.020 -435.280 728.820 -414.720 ;
        RECT -542.230 -970.775 -541.950 -970.495 ;
        RECT -541.470 -970.775 -541.190 -970.495 ;
        RECT -540.710 -970.775 -540.430 -970.495 ;
        RECT -542.230 -971.535 -541.950 -971.255 ;
        RECT -541.470 -971.535 -541.190 -971.255 ;
        RECT -540.710 -971.535 -540.430 -971.255 ;
        RECT -542.230 -972.295 -541.950 -972.015 ;
        RECT -541.470 -972.295 -541.190 -972.015 ;
        RECT -540.710 -972.295 -540.430 -972.015 ;
        RECT -542.230 -973.055 -541.950 -972.775 ;
        RECT -541.470 -973.055 -541.190 -972.775 ;
        RECT -540.710 -973.055 -540.430 -972.775 ;
        RECT -542.230 -973.815 -541.950 -973.535 ;
        RECT -541.470 -973.815 -541.190 -973.535 ;
        RECT -540.710 -973.815 -540.430 -973.535 ;
        RECT -542.230 -974.575 -541.950 -974.295 ;
        RECT -541.470 -974.575 -541.190 -974.295 ;
        RECT -540.710 -974.575 -540.430 -974.295 ;
        RECT -506.530 -970.775 -506.250 -970.495 ;
        RECT -505.770 -970.775 -505.490 -970.495 ;
        RECT -505.010 -970.775 -504.730 -970.495 ;
        RECT -506.530 -971.535 -506.250 -971.255 ;
        RECT -505.770 -971.535 -505.490 -971.255 ;
        RECT -505.010 -971.535 -504.730 -971.255 ;
        RECT -506.530 -972.295 -506.250 -972.015 ;
        RECT -505.770 -972.295 -505.490 -972.015 ;
        RECT -505.010 -972.295 -504.730 -972.015 ;
        RECT -506.530 -973.055 -506.250 -972.775 ;
        RECT -505.770 -973.055 -505.490 -972.775 ;
        RECT -505.010 -973.055 -504.730 -972.775 ;
        RECT -506.530 -973.815 -506.250 -973.535 ;
        RECT -505.770 -973.815 -505.490 -973.535 ;
        RECT -505.010 -973.815 -504.730 -973.535 ;
        RECT -506.530 -974.575 -506.250 -974.295 ;
        RECT -505.770 -974.575 -505.490 -974.295 ;
        RECT -505.010 -974.575 -504.730 -974.295 ;
        RECT -467.230 -970.775 -466.950 -970.495 ;
        RECT -466.470 -970.775 -466.190 -970.495 ;
        RECT -465.710 -970.775 -465.430 -970.495 ;
        RECT -467.230 -971.535 -466.950 -971.255 ;
        RECT -466.470 -971.535 -466.190 -971.255 ;
        RECT -465.710 -971.535 -465.430 -971.255 ;
        RECT -467.230 -972.295 -466.950 -972.015 ;
        RECT -466.470 -972.295 -466.190 -972.015 ;
        RECT -465.710 -972.295 -465.430 -972.015 ;
        RECT -467.230 -973.055 -466.950 -972.775 ;
        RECT -466.470 -973.055 -466.190 -972.775 ;
        RECT -465.710 -973.055 -465.430 -972.775 ;
        RECT -467.230 -973.815 -466.950 -973.535 ;
        RECT -466.470 -973.815 -466.190 -973.535 ;
        RECT -465.710 -973.815 -465.430 -973.535 ;
        RECT -467.230 -974.575 -466.950 -974.295 ;
        RECT -466.470 -974.575 -466.190 -974.295 ;
        RECT -465.710 -974.575 -465.430 -974.295 ;
        RECT -431.530 -970.775 -431.250 -970.495 ;
        RECT -430.770 -970.775 -430.490 -970.495 ;
        RECT -430.010 -970.775 -429.730 -970.495 ;
        RECT -431.530 -971.535 -431.250 -971.255 ;
        RECT -430.770 -971.535 -430.490 -971.255 ;
        RECT -430.010 -971.535 -429.730 -971.255 ;
        RECT -431.530 -972.295 -431.250 -972.015 ;
        RECT -430.770 -972.295 -430.490 -972.015 ;
        RECT -430.010 -972.295 -429.730 -972.015 ;
        RECT -431.530 -973.055 -431.250 -972.775 ;
        RECT -430.770 -973.055 -430.490 -972.775 ;
        RECT -430.010 -973.055 -429.730 -972.775 ;
        RECT -431.530 -973.815 -431.250 -973.535 ;
        RECT -430.770 -973.815 -430.490 -973.535 ;
        RECT -430.010 -973.815 -429.730 -973.535 ;
        RECT -431.530 -974.575 -431.250 -974.295 ;
        RECT -430.770 -974.575 -430.490 -974.295 ;
        RECT -430.010 -974.575 -429.730 -974.295 ;
        RECT -392.230 -970.775 -391.950 -970.495 ;
        RECT -391.470 -970.775 -391.190 -970.495 ;
        RECT -390.710 -970.775 -390.430 -970.495 ;
        RECT -392.230 -971.535 -391.950 -971.255 ;
        RECT -391.470 -971.535 -391.190 -971.255 ;
        RECT -390.710 -971.535 -390.430 -971.255 ;
        RECT -392.230 -972.295 -391.950 -972.015 ;
        RECT -391.470 -972.295 -391.190 -972.015 ;
        RECT -390.710 -972.295 -390.430 -972.015 ;
        RECT -392.230 -973.055 -391.950 -972.775 ;
        RECT -391.470 -973.055 -391.190 -972.775 ;
        RECT -390.710 -973.055 -390.430 -972.775 ;
        RECT -392.230 -973.815 -391.950 -973.535 ;
        RECT -391.470 -973.815 -391.190 -973.535 ;
        RECT -390.710 -973.815 -390.430 -973.535 ;
        RECT -392.230 -974.575 -391.950 -974.295 ;
        RECT -391.470 -974.575 -391.190 -974.295 ;
        RECT -390.710 -974.575 -390.430 -974.295 ;
        RECT -356.530 -970.775 -356.250 -970.495 ;
        RECT -355.770 -970.775 -355.490 -970.495 ;
        RECT -355.010 -970.775 -354.730 -970.495 ;
        RECT -356.530 -971.535 -356.250 -971.255 ;
        RECT -355.770 -971.535 -355.490 -971.255 ;
        RECT -355.010 -971.535 -354.730 -971.255 ;
        RECT -356.530 -972.295 -356.250 -972.015 ;
        RECT -355.770 -972.295 -355.490 -972.015 ;
        RECT -355.010 -972.295 -354.730 -972.015 ;
        RECT -356.530 -973.055 -356.250 -972.775 ;
        RECT -355.770 -973.055 -355.490 -972.775 ;
        RECT -355.010 -973.055 -354.730 -972.775 ;
        RECT -356.530 -973.815 -356.250 -973.535 ;
        RECT -355.770 -973.815 -355.490 -973.535 ;
        RECT -355.010 -973.815 -354.730 -973.535 ;
        RECT -356.530 -974.575 -356.250 -974.295 ;
        RECT -355.770 -974.575 -355.490 -974.295 ;
        RECT -355.010 -974.575 -354.730 -974.295 ;
        RECT -317.230 -970.775 -316.950 -970.495 ;
        RECT -316.470 -970.775 -316.190 -970.495 ;
        RECT -315.710 -970.775 -315.430 -970.495 ;
        RECT -317.230 -971.535 -316.950 -971.255 ;
        RECT -316.470 -971.535 -316.190 -971.255 ;
        RECT -315.710 -971.535 -315.430 -971.255 ;
        RECT -317.230 -972.295 -316.950 -972.015 ;
        RECT -316.470 -972.295 -316.190 -972.015 ;
        RECT -315.710 -972.295 -315.430 -972.015 ;
        RECT -317.230 -973.055 -316.950 -972.775 ;
        RECT -316.470 -973.055 -316.190 -972.775 ;
        RECT -315.710 -973.055 -315.430 -972.775 ;
        RECT -317.230 -973.815 -316.950 -973.535 ;
        RECT -316.470 -973.815 -316.190 -973.535 ;
        RECT -315.710 -973.815 -315.430 -973.535 ;
        RECT -317.230 -974.575 -316.950 -974.295 ;
        RECT -316.470 -974.575 -316.190 -974.295 ;
        RECT -315.710 -974.575 -315.430 -974.295 ;
        RECT -281.530 -970.775 -281.250 -970.495 ;
        RECT -280.770 -970.775 -280.490 -970.495 ;
        RECT -280.010 -970.775 -279.730 -970.495 ;
        RECT -281.530 -971.535 -281.250 -971.255 ;
        RECT -280.770 -971.535 -280.490 -971.255 ;
        RECT -280.010 -971.535 -279.730 -971.255 ;
        RECT -281.530 -972.295 -281.250 -972.015 ;
        RECT -280.770 -972.295 -280.490 -972.015 ;
        RECT -280.010 -972.295 -279.730 -972.015 ;
        RECT -281.530 -973.055 -281.250 -972.775 ;
        RECT -280.770 -973.055 -280.490 -972.775 ;
        RECT -280.010 -973.055 -279.730 -972.775 ;
        RECT -281.530 -973.815 -281.250 -973.535 ;
        RECT -280.770 -973.815 -280.490 -973.535 ;
        RECT -280.010 -973.815 -279.730 -973.535 ;
        RECT -281.530 -974.575 -281.250 -974.295 ;
        RECT -280.770 -974.575 -280.490 -974.295 ;
        RECT -280.010 -974.575 -279.730 -974.295 ;
        RECT -242.230 -970.775 -241.950 -970.495 ;
        RECT -241.470 -970.775 -241.190 -970.495 ;
        RECT -240.710 -970.775 -240.430 -970.495 ;
        RECT -242.230 -971.535 -241.950 -971.255 ;
        RECT -241.470 -971.535 -241.190 -971.255 ;
        RECT -240.710 -971.535 -240.430 -971.255 ;
        RECT -242.230 -972.295 -241.950 -972.015 ;
        RECT -241.470 -972.295 -241.190 -972.015 ;
        RECT -240.710 -972.295 -240.430 -972.015 ;
        RECT -242.230 -973.055 -241.950 -972.775 ;
        RECT -241.470 -973.055 -241.190 -972.775 ;
        RECT -240.710 -973.055 -240.430 -972.775 ;
        RECT -242.230 -973.815 -241.950 -973.535 ;
        RECT -241.470 -973.815 -241.190 -973.535 ;
        RECT -240.710 -973.815 -240.430 -973.535 ;
        RECT -242.230 -974.575 -241.950 -974.295 ;
        RECT -241.470 -974.575 -241.190 -974.295 ;
        RECT -240.710 -974.575 -240.430 -974.295 ;
        RECT -206.530 -970.775 -206.250 -970.495 ;
        RECT -205.770 -970.775 -205.490 -970.495 ;
        RECT -205.010 -970.775 -204.730 -970.495 ;
        RECT -206.530 -971.535 -206.250 -971.255 ;
        RECT -205.770 -971.535 -205.490 -971.255 ;
        RECT -205.010 -971.535 -204.730 -971.255 ;
        RECT -206.530 -972.295 -206.250 -972.015 ;
        RECT -205.770 -972.295 -205.490 -972.015 ;
        RECT -205.010 -972.295 -204.730 -972.015 ;
        RECT -206.530 -973.055 -206.250 -972.775 ;
        RECT -205.770 -973.055 -205.490 -972.775 ;
        RECT -205.010 -973.055 -204.730 -972.775 ;
        RECT -206.530 -973.815 -206.250 -973.535 ;
        RECT -205.770 -973.815 -205.490 -973.535 ;
        RECT -205.010 -973.815 -204.730 -973.535 ;
        RECT -206.530 -974.575 -206.250 -974.295 ;
        RECT -205.770 -974.575 -205.490 -974.295 ;
        RECT -205.010 -974.575 -204.730 -974.295 ;
        RECT -167.230 -970.775 -166.950 -970.495 ;
        RECT -166.470 -970.775 -166.190 -970.495 ;
        RECT -165.710 -970.775 -165.430 -970.495 ;
        RECT -167.230 -971.535 -166.950 -971.255 ;
        RECT -166.470 -971.535 -166.190 -971.255 ;
        RECT -165.710 -971.535 -165.430 -971.255 ;
        RECT -167.230 -972.295 -166.950 -972.015 ;
        RECT -166.470 -972.295 -166.190 -972.015 ;
        RECT -165.710 -972.295 -165.430 -972.015 ;
        RECT -167.230 -973.055 -166.950 -972.775 ;
        RECT -166.470 -973.055 -166.190 -972.775 ;
        RECT -165.710 -973.055 -165.430 -972.775 ;
        RECT -167.230 -973.815 -166.950 -973.535 ;
        RECT -166.470 -973.815 -166.190 -973.535 ;
        RECT -165.710 -973.815 -165.430 -973.535 ;
        RECT -167.230 -974.575 -166.950 -974.295 ;
        RECT -166.470 -974.575 -166.190 -974.295 ;
        RECT -165.710 -974.575 -165.430 -974.295 ;
        RECT -131.530 -970.775 -131.250 -970.495 ;
        RECT -130.770 -970.775 -130.490 -970.495 ;
        RECT -130.010 -970.775 -129.730 -970.495 ;
        RECT -131.530 -971.535 -131.250 -971.255 ;
        RECT -130.770 -971.535 -130.490 -971.255 ;
        RECT -130.010 -971.535 -129.730 -971.255 ;
        RECT -131.530 -972.295 -131.250 -972.015 ;
        RECT -130.770 -972.295 -130.490 -972.015 ;
        RECT -130.010 -972.295 -129.730 -972.015 ;
        RECT -131.530 -973.055 -131.250 -972.775 ;
        RECT -130.770 -973.055 -130.490 -972.775 ;
        RECT -130.010 -973.055 -129.730 -972.775 ;
        RECT -131.530 -973.815 -131.250 -973.535 ;
        RECT -130.770 -973.815 -130.490 -973.535 ;
        RECT -130.010 -973.815 -129.730 -973.535 ;
        RECT -131.530 -974.575 -131.250 -974.295 ;
        RECT -130.770 -974.575 -130.490 -974.295 ;
        RECT -130.010 -974.575 -129.730 -974.295 ;
        RECT -92.230 -970.775 -91.950 -970.495 ;
        RECT -91.470 -970.775 -91.190 -970.495 ;
        RECT -90.710 -970.775 -90.430 -970.495 ;
        RECT -92.230 -971.535 -91.950 -971.255 ;
        RECT -91.470 -971.535 -91.190 -971.255 ;
        RECT -90.710 -971.535 -90.430 -971.255 ;
        RECT -92.230 -972.295 -91.950 -972.015 ;
        RECT -91.470 -972.295 -91.190 -972.015 ;
        RECT -90.710 -972.295 -90.430 -972.015 ;
        RECT -92.230 -973.055 -91.950 -972.775 ;
        RECT -91.470 -973.055 -91.190 -972.775 ;
        RECT -90.710 -973.055 -90.430 -972.775 ;
        RECT -92.230 -973.815 -91.950 -973.535 ;
        RECT -91.470 -973.815 -91.190 -973.535 ;
        RECT -90.710 -973.815 -90.430 -973.535 ;
        RECT -92.230 -974.575 -91.950 -974.295 ;
        RECT -91.470 -974.575 -91.190 -974.295 ;
        RECT -90.710 -974.575 -90.430 -974.295 ;
        RECT -56.530 -970.775 -56.250 -970.495 ;
        RECT -55.770 -970.775 -55.490 -970.495 ;
        RECT -55.010 -970.775 -54.730 -970.495 ;
        RECT -56.530 -971.535 -56.250 -971.255 ;
        RECT -55.770 -971.535 -55.490 -971.255 ;
        RECT -55.010 -971.535 -54.730 -971.255 ;
        RECT -56.530 -972.295 -56.250 -972.015 ;
        RECT -55.770 -972.295 -55.490 -972.015 ;
        RECT -55.010 -972.295 -54.730 -972.015 ;
        RECT -56.530 -973.055 -56.250 -972.775 ;
        RECT -55.770 -973.055 -55.490 -972.775 ;
        RECT -55.010 -973.055 -54.730 -972.775 ;
        RECT -56.530 -973.815 -56.250 -973.535 ;
        RECT -55.770 -973.815 -55.490 -973.535 ;
        RECT -55.010 -973.815 -54.730 -973.535 ;
        RECT -56.530 -974.575 -56.250 -974.295 ;
        RECT -55.770 -974.575 -55.490 -974.295 ;
        RECT -55.010 -974.575 -54.730 -974.295 ;
        RECT -17.230 -970.775 -16.950 -970.495 ;
        RECT -16.470 -970.775 -16.190 -970.495 ;
        RECT -15.710 -970.775 -15.430 -970.495 ;
        RECT -17.230 -971.535 -16.950 -971.255 ;
        RECT -16.470 -971.535 -16.190 -971.255 ;
        RECT -15.710 -971.535 -15.430 -971.255 ;
        RECT -17.230 -972.295 -16.950 -972.015 ;
        RECT -16.470 -972.295 -16.190 -972.015 ;
        RECT -15.710 -972.295 -15.430 -972.015 ;
        RECT -17.230 -973.055 -16.950 -972.775 ;
        RECT -16.470 -973.055 -16.190 -972.775 ;
        RECT -15.710 -973.055 -15.430 -972.775 ;
        RECT -17.230 -973.815 -16.950 -973.535 ;
        RECT -16.470 -973.815 -16.190 -973.535 ;
        RECT -15.710 -973.815 -15.430 -973.535 ;
        RECT -17.230 -974.575 -16.950 -974.295 ;
        RECT -16.470 -974.575 -16.190 -974.295 ;
        RECT -15.710 -974.575 -15.430 -974.295 ;
        RECT 18.470 -970.775 18.750 -970.495 ;
        RECT 19.230 -970.775 19.510 -970.495 ;
        RECT 19.990 -970.775 20.270 -970.495 ;
        RECT 18.470 -971.535 18.750 -971.255 ;
        RECT 19.230 -971.535 19.510 -971.255 ;
        RECT 19.990 -971.535 20.270 -971.255 ;
        RECT 18.470 -972.295 18.750 -972.015 ;
        RECT 19.230 -972.295 19.510 -972.015 ;
        RECT 19.990 -972.295 20.270 -972.015 ;
        RECT 18.470 -973.055 18.750 -972.775 ;
        RECT 19.230 -973.055 19.510 -972.775 ;
        RECT 19.990 -973.055 20.270 -972.775 ;
        RECT 18.470 -973.815 18.750 -973.535 ;
        RECT 19.230 -973.815 19.510 -973.535 ;
        RECT 19.990 -973.815 20.270 -973.535 ;
        RECT 18.470 -974.575 18.750 -974.295 ;
        RECT 19.230 -974.575 19.510 -974.295 ;
        RECT 19.990 -974.575 20.270 -974.295 ;
        RECT 57.770 -970.775 58.050 -970.495 ;
        RECT 58.530 -970.775 58.810 -970.495 ;
        RECT 59.290 -970.775 59.570 -970.495 ;
        RECT 57.770 -971.535 58.050 -971.255 ;
        RECT 58.530 -971.535 58.810 -971.255 ;
        RECT 59.290 -971.535 59.570 -971.255 ;
        RECT 57.770 -972.295 58.050 -972.015 ;
        RECT 58.530 -972.295 58.810 -972.015 ;
        RECT 59.290 -972.295 59.570 -972.015 ;
        RECT 57.770 -973.055 58.050 -972.775 ;
        RECT 58.530 -973.055 58.810 -972.775 ;
        RECT 59.290 -973.055 59.570 -972.775 ;
        RECT 57.770 -973.815 58.050 -973.535 ;
        RECT 58.530 -973.815 58.810 -973.535 ;
        RECT 59.290 -973.815 59.570 -973.535 ;
        RECT 57.770 -974.575 58.050 -974.295 ;
        RECT 58.530 -974.575 58.810 -974.295 ;
        RECT 59.290 -974.575 59.570 -974.295 ;
        RECT 93.470 -970.775 93.750 -970.495 ;
        RECT 94.230 -970.775 94.510 -970.495 ;
        RECT 94.990 -970.775 95.270 -970.495 ;
        RECT 93.470 -971.535 93.750 -971.255 ;
        RECT 94.230 -971.535 94.510 -971.255 ;
        RECT 94.990 -971.535 95.270 -971.255 ;
        RECT 93.470 -972.295 93.750 -972.015 ;
        RECT 94.230 -972.295 94.510 -972.015 ;
        RECT 94.990 -972.295 95.270 -972.015 ;
        RECT 93.470 -973.055 93.750 -972.775 ;
        RECT 94.230 -973.055 94.510 -972.775 ;
        RECT 94.990 -973.055 95.270 -972.775 ;
        RECT 93.470 -973.815 93.750 -973.535 ;
        RECT 94.230 -973.815 94.510 -973.535 ;
        RECT 94.990 -973.815 95.270 -973.535 ;
        RECT 93.470 -974.575 93.750 -974.295 ;
        RECT 94.230 -974.575 94.510 -974.295 ;
        RECT 94.990 -974.575 95.270 -974.295 ;
        RECT 132.770 -970.775 133.050 -970.495 ;
        RECT 133.530 -970.775 133.810 -970.495 ;
        RECT 134.290 -970.775 134.570 -970.495 ;
        RECT 132.770 -971.535 133.050 -971.255 ;
        RECT 133.530 -971.535 133.810 -971.255 ;
        RECT 134.290 -971.535 134.570 -971.255 ;
        RECT 132.770 -972.295 133.050 -972.015 ;
        RECT 133.530 -972.295 133.810 -972.015 ;
        RECT 134.290 -972.295 134.570 -972.015 ;
        RECT 132.770 -973.055 133.050 -972.775 ;
        RECT 133.530 -973.055 133.810 -972.775 ;
        RECT 134.290 -973.055 134.570 -972.775 ;
        RECT 132.770 -973.815 133.050 -973.535 ;
        RECT 133.530 -973.815 133.810 -973.535 ;
        RECT 134.290 -973.815 134.570 -973.535 ;
        RECT 132.770 -974.575 133.050 -974.295 ;
        RECT 133.530 -974.575 133.810 -974.295 ;
        RECT 134.290 -974.575 134.570 -974.295 ;
        RECT 168.470 -970.775 168.750 -970.495 ;
        RECT 169.230 -970.775 169.510 -970.495 ;
        RECT 169.990 -970.775 170.270 -970.495 ;
        RECT 168.470 -971.535 168.750 -971.255 ;
        RECT 169.230 -971.535 169.510 -971.255 ;
        RECT 169.990 -971.535 170.270 -971.255 ;
        RECT 168.470 -972.295 168.750 -972.015 ;
        RECT 169.230 -972.295 169.510 -972.015 ;
        RECT 169.990 -972.295 170.270 -972.015 ;
        RECT 168.470 -973.055 168.750 -972.775 ;
        RECT 169.230 -973.055 169.510 -972.775 ;
        RECT 169.990 -973.055 170.270 -972.775 ;
        RECT 168.470 -973.815 168.750 -973.535 ;
        RECT 169.230 -973.815 169.510 -973.535 ;
        RECT 169.990 -973.815 170.270 -973.535 ;
        RECT 168.470 -974.575 168.750 -974.295 ;
        RECT 169.230 -974.575 169.510 -974.295 ;
        RECT 169.990 -974.575 170.270 -974.295 ;
        RECT 207.770 -970.775 208.050 -970.495 ;
        RECT 208.530 -970.775 208.810 -970.495 ;
        RECT 209.290 -970.775 209.570 -970.495 ;
        RECT 207.770 -971.535 208.050 -971.255 ;
        RECT 208.530 -971.535 208.810 -971.255 ;
        RECT 209.290 -971.535 209.570 -971.255 ;
        RECT 207.770 -972.295 208.050 -972.015 ;
        RECT 208.530 -972.295 208.810 -972.015 ;
        RECT 209.290 -972.295 209.570 -972.015 ;
        RECT 207.770 -973.055 208.050 -972.775 ;
        RECT 208.530 -973.055 208.810 -972.775 ;
        RECT 209.290 -973.055 209.570 -972.775 ;
        RECT 207.770 -973.815 208.050 -973.535 ;
        RECT 208.530 -973.815 208.810 -973.535 ;
        RECT 209.290 -973.815 209.570 -973.535 ;
        RECT 207.770 -974.575 208.050 -974.295 ;
        RECT 208.530 -974.575 208.810 -974.295 ;
        RECT 209.290 -974.575 209.570 -974.295 ;
        RECT 243.470 -970.775 243.750 -970.495 ;
        RECT 244.230 -970.775 244.510 -970.495 ;
        RECT 244.990 -970.775 245.270 -970.495 ;
        RECT 243.470 -971.535 243.750 -971.255 ;
        RECT 244.230 -971.535 244.510 -971.255 ;
        RECT 244.990 -971.535 245.270 -971.255 ;
        RECT 243.470 -972.295 243.750 -972.015 ;
        RECT 244.230 -972.295 244.510 -972.015 ;
        RECT 244.990 -972.295 245.270 -972.015 ;
        RECT 243.470 -973.055 243.750 -972.775 ;
        RECT 244.230 -973.055 244.510 -972.775 ;
        RECT 244.990 -973.055 245.270 -972.775 ;
        RECT 243.470 -973.815 243.750 -973.535 ;
        RECT 244.230 -973.815 244.510 -973.535 ;
        RECT 244.990 -973.815 245.270 -973.535 ;
        RECT 243.470 -974.575 243.750 -974.295 ;
        RECT 244.230 -974.575 244.510 -974.295 ;
        RECT 244.990 -974.575 245.270 -974.295 ;
        RECT 282.770 -970.775 283.050 -970.495 ;
        RECT 283.530 -970.775 283.810 -970.495 ;
        RECT 284.290 -970.775 284.570 -970.495 ;
        RECT 282.770 -971.535 283.050 -971.255 ;
        RECT 283.530 -971.535 283.810 -971.255 ;
        RECT 284.290 -971.535 284.570 -971.255 ;
        RECT 282.770 -972.295 283.050 -972.015 ;
        RECT 283.530 -972.295 283.810 -972.015 ;
        RECT 284.290 -972.295 284.570 -972.015 ;
        RECT 282.770 -973.055 283.050 -972.775 ;
        RECT 283.530 -973.055 283.810 -972.775 ;
        RECT 284.290 -973.055 284.570 -972.775 ;
        RECT 282.770 -973.815 283.050 -973.535 ;
        RECT 283.530 -973.815 283.810 -973.535 ;
        RECT 284.290 -973.815 284.570 -973.535 ;
        RECT 282.770 -974.575 283.050 -974.295 ;
        RECT 283.530 -974.575 283.810 -974.295 ;
        RECT 284.290 -974.575 284.570 -974.295 ;
        RECT 318.470 -970.775 318.750 -970.495 ;
        RECT 319.230 -970.775 319.510 -970.495 ;
        RECT 319.990 -970.775 320.270 -970.495 ;
        RECT 318.470 -971.535 318.750 -971.255 ;
        RECT 319.230 -971.535 319.510 -971.255 ;
        RECT 319.990 -971.535 320.270 -971.255 ;
        RECT 318.470 -972.295 318.750 -972.015 ;
        RECT 319.230 -972.295 319.510 -972.015 ;
        RECT 319.990 -972.295 320.270 -972.015 ;
        RECT 318.470 -973.055 318.750 -972.775 ;
        RECT 319.230 -973.055 319.510 -972.775 ;
        RECT 319.990 -973.055 320.270 -972.775 ;
        RECT 318.470 -973.815 318.750 -973.535 ;
        RECT 319.230 -973.815 319.510 -973.535 ;
        RECT 319.990 -973.815 320.270 -973.535 ;
        RECT 318.470 -974.575 318.750 -974.295 ;
        RECT 319.230 -974.575 319.510 -974.295 ;
        RECT 319.990 -974.575 320.270 -974.295 ;
        RECT 357.770 -970.775 358.050 -970.495 ;
        RECT 358.530 -970.775 358.810 -970.495 ;
        RECT 359.290 -970.775 359.570 -970.495 ;
        RECT 357.770 -971.535 358.050 -971.255 ;
        RECT 358.530 -971.535 358.810 -971.255 ;
        RECT 359.290 -971.535 359.570 -971.255 ;
        RECT 357.770 -972.295 358.050 -972.015 ;
        RECT 358.530 -972.295 358.810 -972.015 ;
        RECT 359.290 -972.295 359.570 -972.015 ;
        RECT 357.770 -973.055 358.050 -972.775 ;
        RECT 358.530 -973.055 358.810 -972.775 ;
        RECT 359.290 -973.055 359.570 -972.775 ;
        RECT 357.770 -973.815 358.050 -973.535 ;
        RECT 358.530 -973.815 358.810 -973.535 ;
        RECT 359.290 -973.815 359.570 -973.535 ;
        RECT 357.770 -974.575 358.050 -974.295 ;
        RECT 358.530 -974.575 358.810 -974.295 ;
        RECT 359.290 -974.575 359.570 -974.295 ;
        RECT 393.470 -970.775 393.750 -970.495 ;
        RECT 394.230 -970.775 394.510 -970.495 ;
        RECT 394.990 -970.775 395.270 -970.495 ;
        RECT 393.470 -971.535 393.750 -971.255 ;
        RECT 394.230 -971.535 394.510 -971.255 ;
        RECT 394.990 -971.535 395.270 -971.255 ;
        RECT 393.470 -972.295 393.750 -972.015 ;
        RECT 394.230 -972.295 394.510 -972.015 ;
        RECT 394.990 -972.295 395.270 -972.015 ;
        RECT 393.470 -973.055 393.750 -972.775 ;
        RECT 394.230 -973.055 394.510 -972.775 ;
        RECT 394.990 -973.055 395.270 -972.775 ;
        RECT 393.470 -973.815 393.750 -973.535 ;
        RECT 394.230 -973.815 394.510 -973.535 ;
        RECT 394.990 -973.815 395.270 -973.535 ;
        RECT 393.470 -974.575 393.750 -974.295 ;
        RECT 394.230 -974.575 394.510 -974.295 ;
        RECT 394.990 -974.575 395.270 -974.295 ;
        RECT 432.770 -970.775 433.050 -970.495 ;
        RECT 433.530 -970.775 433.810 -970.495 ;
        RECT 434.290 -970.775 434.570 -970.495 ;
        RECT 432.770 -971.535 433.050 -971.255 ;
        RECT 433.530 -971.535 433.810 -971.255 ;
        RECT 434.290 -971.535 434.570 -971.255 ;
        RECT 432.770 -972.295 433.050 -972.015 ;
        RECT 433.530 -972.295 433.810 -972.015 ;
        RECT 434.290 -972.295 434.570 -972.015 ;
        RECT 432.770 -973.055 433.050 -972.775 ;
        RECT 433.530 -973.055 433.810 -972.775 ;
        RECT 434.290 -973.055 434.570 -972.775 ;
        RECT 432.770 -973.815 433.050 -973.535 ;
        RECT 433.530 -973.815 433.810 -973.535 ;
        RECT 434.290 -973.815 434.570 -973.535 ;
        RECT 432.770 -974.575 433.050 -974.295 ;
        RECT 433.530 -974.575 433.810 -974.295 ;
        RECT 434.290 -974.575 434.570 -974.295 ;
        RECT 468.470 -970.775 468.750 -970.495 ;
        RECT 469.230 -970.775 469.510 -970.495 ;
        RECT 469.990 -970.775 470.270 -970.495 ;
        RECT 468.470 -971.535 468.750 -971.255 ;
        RECT 469.230 -971.535 469.510 -971.255 ;
        RECT 469.990 -971.535 470.270 -971.255 ;
        RECT 468.470 -972.295 468.750 -972.015 ;
        RECT 469.230 -972.295 469.510 -972.015 ;
        RECT 469.990 -972.295 470.270 -972.015 ;
        RECT 468.470 -973.055 468.750 -972.775 ;
        RECT 469.230 -973.055 469.510 -972.775 ;
        RECT 469.990 -973.055 470.270 -972.775 ;
        RECT 468.470 -973.815 468.750 -973.535 ;
        RECT 469.230 -973.815 469.510 -973.535 ;
        RECT 469.990 -973.815 470.270 -973.535 ;
        RECT 468.470 -974.575 468.750 -974.295 ;
        RECT 469.230 -974.575 469.510 -974.295 ;
        RECT 469.990 -974.575 470.270 -974.295 ;
        RECT 507.770 -970.775 508.050 -970.495 ;
        RECT 508.530 -970.775 508.810 -970.495 ;
        RECT 509.290 -970.775 509.570 -970.495 ;
        RECT 507.770 -971.535 508.050 -971.255 ;
        RECT 508.530 -971.535 508.810 -971.255 ;
        RECT 509.290 -971.535 509.570 -971.255 ;
        RECT 507.770 -972.295 508.050 -972.015 ;
        RECT 508.530 -972.295 508.810 -972.015 ;
        RECT 509.290 -972.295 509.570 -972.015 ;
        RECT 507.770 -973.055 508.050 -972.775 ;
        RECT 508.530 -973.055 508.810 -972.775 ;
        RECT 509.290 -973.055 509.570 -972.775 ;
        RECT 507.770 -973.815 508.050 -973.535 ;
        RECT 508.530 -973.815 508.810 -973.535 ;
        RECT 509.290 -973.815 509.570 -973.535 ;
        RECT 507.770 -974.575 508.050 -974.295 ;
        RECT 508.530 -974.575 508.810 -974.295 ;
        RECT 509.290 -974.575 509.570 -974.295 ;
        RECT 543.470 -970.775 543.750 -970.495 ;
        RECT 544.230 -970.775 544.510 -970.495 ;
        RECT 544.990 -970.775 545.270 -970.495 ;
        RECT 543.470 -971.535 543.750 -971.255 ;
        RECT 544.230 -971.535 544.510 -971.255 ;
        RECT 544.990 -971.535 545.270 -971.255 ;
        RECT 543.470 -972.295 543.750 -972.015 ;
        RECT 544.230 -972.295 544.510 -972.015 ;
        RECT 544.990 -972.295 545.270 -972.015 ;
        RECT 543.470 -973.055 543.750 -972.775 ;
        RECT 544.230 -973.055 544.510 -972.775 ;
        RECT 544.990 -973.055 545.270 -972.775 ;
        RECT 543.470 -973.815 543.750 -973.535 ;
        RECT 544.230 -973.815 544.510 -973.535 ;
        RECT 544.990 -973.815 545.270 -973.535 ;
        RECT 543.470 -974.575 543.750 -974.295 ;
        RECT 544.230 -974.575 544.510 -974.295 ;
        RECT 544.990 -974.575 545.270 -974.295 ;
    END
  END vdd
  PIN result[9]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 12.360 444.265 12.725 ;
        RECT 446.245 12.360 446.475 12.725 ;
        RECT 448.485 12.360 448.715 12.725 ;
        RECT 450.725 12.360 450.955 12.725 ;
        RECT 444.005 11.980 450.955 12.360 ;
        RECT 447.000 11.070 447.800 11.980 ;
        RECT 444.005 10.690 450.855 11.070 ;
        RECT 444.005 10.020 444.235 10.690 ;
        RECT 446.145 10.020 446.375 10.690 ;
        RECT 448.385 10.020 448.615 10.690 ;
        RECT 450.625 10.020 450.855 10.690 ;
      LAYER Via1 ;
        RECT 444.470 10.750 444.730 11.010 ;
      LAYER Metal2 ;
        RECT 444.460 10.690 444.740 40.750 ;
        RECT 447.260 40.370 447.540 58.670 ;
      LAYER Via2 ;
        RECT 447.260 58.340 447.540 58.620 ;
        RECT 444.460 40.420 444.740 40.700 ;
        RECT 447.260 40.420 447.540 40.700 ;
      LAYER Metal3 ;
        RECT 465.200 58.620 654.000 58.760 ;
        RECT 447.210 58.340 654.000 58.620 ;
        RECT 465.200 58.200 654.000 58.340 ;
        RECT 444.410 40.420 447.590 40.700 ;
    END
  END result[9]
  PIN result[8]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 409.845 39.630 410.075 40.300 ;
        RECT 411.985 39.630 412.215 40.300 ;
        RECT 414.225 39.630 414.455 40.300 ;
        RECT 416.465 39.630 416.695 40.300 ;
        RECT 409.845 39.250 416.695 39.630 ;
        RECT 412.840 38.340 413.640 39.250 ;
        RECT 409.845 37.960 416.795 38.340 ;
        RECT 409.845 37.595 410.105 37.960 ;
        RECT 412.085 37.595 412.315 37.960 ;
        RECT 414.325 37.595 414.555 37.960 ;
        RECT 416.565 37.595 416.795 37.960 ;
      LAYER Via1 ;
        RECT 414.790 39.310 415.050 39.570 ;
      LAYER Metal2 ;
        RECT 414.780 39.250 415.060 50.830 ;
      LAYER Via2 ;
        RECT 414.780 50.500 415.060 50.780 ;
      LAYER Metal3 ;
        RECT 465.200 50.780 654.000 50.920 ;
        RECT 414.730 50.500 654.000 50.780 ;
        RECT 465.200 50.360 654.000 50.500 ;
    END
  END result[8]
  PIN result[7]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 429.445 28.040 429.705 28.405 ;
        RECT 431.685 28.040 431.915 28.405 ;
        RECT 433.925 28.040 434.155 28.405 ;
        RECT 436.165 28.040 436.395 28.405 ;
        RECT 429.445 27.660 436.395 28.040 ;
        RECT 432.440 26.750 433.240 27.660 ;
        RECT 429.445 26.370 436.330 26.750 ;
        RECT 429.445 25.700 429.675 26.370 ;
        RECT 431.585 25.700 431.815 26.370 ;
        RECT 433.825 25.700 434.055 26.370 ;
        RECT 436.065 25.700 436.295 26.370 ;
      LAYER Via1 ;
        RECT 436.070 26.430 436.330 26.690 ;
      LAYER Metal2 ;
        RECT 436.060 26.370 436.340 28.430 ;
        RECT 445.020 28.050 445.300 42.990 ;
      LAYER Via2 ;
        RECT 445.020 42.660 445.300 42.940 ;
        RECT 436.060 28.100 436.340 28.380 ;
        RECT 445.020 28.100 445.300 28.380 ;
      LAYER Metal3 ;
        RECT 465.200 42.940 654.000 43.080 ;
        RECT 444.970 42.660 654.000 42.940 ;
        RECT 465.200 42.520 654.000 42.660 ;
        RECT 436.010 28.100 445.350 28.380 ;
    END
  END result[7]
  PIN result[6]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 424.965 35.880 425.225 36.245 ;
        RECT 427.205 35.880 427.435 36.245 ;
        RECT 429.445 35.880 429.675 36.245 ;
        RECT 431.685 35.880 431.915 36.245 ;
        RECT 424.965 35.500 431.915 35.880 ;
        RECT 427.960 34.590 428.760 35.500 ;
        RECT 424.965 34.210 431.850 34.590 ;
        RECT 424.965 33.540 425.195 34.210 ;
        RECT 427.105 33.540 427.335 34.210 ;
        RECT 429.345 33.540 429.575 34.210 ;
        RECT 431.585 33.540 431.815 34.210 ;
      LAYER Via1 ;
        RECT 431.590 34.270 431.850 34.530 ;
      LAYER Metal2 ;
        RECT 431.580 34.210 431.860 35.150 ;
      LAYER Via2 ;
        RECT 431.580 34.820 431.860 35.100 ;
      LAYER Metal3 ;
        RECT 465.200 35.100 654.000 35.240 ;
        RECT 431.530 34.820 654.000 35.100 ;
        RECT 465.200 34.680 654.000 34.820 ;
    END
  END result[6]
  PIN result[5]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 28.040 444.265 28.405 ;
        RECT 446.245 28.040 446.475 28.405 ;
        RECT 448.485 28.040 448.715 28.405 ;
        RECT 450.725 28.040 450.955 28.405 ;
        RECT 444.005 27.660 450.955 28.040 ;
        RECT 447.000 26.750 447.800 27.660 ;
        RECT 444.005 26.370 450.855 26.750 ;
        RECT 444.005 25.700 444.235 26.370 ;
        RECT 446.145 25.700 446.375 26.370 ;
        RECT 448.385 25.700 448.615 26.370 ;
        RECT 450.625 25.700 450.855 26.370 ;
      LAYER Via1 ;
        RECT 448.390 26.430 448.650 26.690 ;
      LAYER Metal2 ;
        RECT 448.380 26.370 448.660 27.310 ;
      LAYER Via2 ;
        RECT 448.380 26.980 448.660 27.260 ;
      LAYER Metal3 ;
        RECT 465.200 27.260 654.000 27.400 ;
        RECT 448.330 26.980 654.000 27.260 ;
        RECT 465.200 26.840 654.000 26.980 ;
    END
  END result[5]
  PIN result[4]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 20.200 444.265 20.565 ;
        RECT 446.245 20.200 446.475 20.565 ;
        RECT 448.485 20.200 448.715 20.565 ;
        RECT 450.725 20.200 450.955 20.565 ;
        RECT 444.005 19.820 450.955 20.200 ;
        RECT 447.000 18.910 447.800 19.820 ;
        RECT 444.005 18.530 450.855 18.910 ;
        RECT 444.005 17.860 444.235 18.530 ;
        RECT 446.145 17.860 446.375 18.530 ;
        RECT 448.385 17.860 448.615 18.530 ;
        RECT 450.625 17.860 450.855 18.530 ;
      LAYER Via1 ;
        RECT 447.270 19.150 447.530 19.410 ;
      LAYER Metal2 ;
        RECT 447.260 18.950 447.540 19.470 ;
      LAYER Via2 ;
        RECT 447.260 19.140 447.540 19.420 ;
      LAYER Metal3 ;
        RECT 465.200 19.420 654.000 19.560 ;
        RECT 447.210 19.140 654.000 19.420 ;
        RECT 465.200 19.000 654.000 19.140 ;
    END
  END result[4]
  PIN result[3]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 452.405 8.270 452.635 8.940 ;
        RECT 454.545 8.270 454.775 8.940 ;
        RECT 456.785 8.770 457.015 8.940 ;
        RECT 456.730 8.510 457.110 8.770 ;
        RECT 456.785 8.270 457.015 8.510 ;
        RECT 459.025 8.270 459.255 8.940 ;
        RECT 452.405 7.890 459.255 8.270 ;
        RECT 455.400 6.980 456.200 7.890 ;
        RECT 452.405 6.600 459.355 6.980 ;
        RECT 452.405 6.235 452.665 6.600 ;
        RECT 454.645 6.235 454.875 6.600 ;
        RECT 456.885 6.235 457.115 6.600 ;
        RECT 459.125 6.235 459.355 6.600 ;
      LAYER Via1 ;
        RECT 456.790 8.510 457.050 8.770 ;
      LAYER Metal2 ;
        RECT 456.780 8.450 457.060 11.630 ;
      LAYER Via2 ;
        RECT 456.780 11.300 457.060 11.580 ;
      LAYER Metal3 ;
        RECT 465.200 11.580 654.000 11.720 ;
        RECT 456.730 11.300 654.000 11.580 ;
        RECT 465.200 11.160 654.000 11.300 ;
    END
  END result[3]
  PIN result[2]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 4.520 444.265 4.885 ;
        RECT 446.245 4.520 446.475 4.885 ;
        RECT 448.485 4.520 448.715 4.885 ;
        RECT 450.725 4.520 450.955 4.885 ;
        RECT 444.005 4.140 450.955 4.520 ;
        RECT 447.000 3.230 447.800 4.140 ;
        RECT 444.005 2.850 450.855 3.230 ;
        RECT 444.005 2.180 444.235 2.850 ;
        RECT 446.145 2.180 446.375 2.850 ;
        RECT 448.385 2.180 448.615 2.850 ;
        RECT 450.625 2.180 450.855 2.850 ;
      LAYER Via1 ;
        RECT 448.390 2.910 448.650 3.170 ;
      LAYER Metal2 ;
        RECT 448.380 2.710 448.660 3.230 ;
      LAYER Via2 ;
        RECT 448.380 2.900 448.660 3.180 ;
      LAYER Metal3 ;
        RECT 448.660 4.020 457.620 4.300 ;
        RECT 448.660 3.180 448.940 4.020 ;
        RECT 457.340 3.740 457.620 4.020 ;
        RECT 465.200 3.740 654.000 3.880 ;
        RECT 457.340 3.460 654.000 3.740 ;
        RECT 465.200 3.320 654.000 3.460 ;
        RECT 448.330 2.900 448.940 3.180 ;
    END
  END result[2]
  PIN result[1]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 -3.320 444.265 -2.955 ;
        RECT 446.245 -3.320 446.475 -2.955 ;
        RECT 448.485 -3.320 448.715 -2.955 ;
        RECT 450.725 -3.320 450.955 -2.955 ;
        RECT 444.005 -3.700 450.955 -3.320 ;
        RECT 447.000 -4.610 447.800 -3.700 ;
        RECT 444.005 -4.990 450.855 -4.610 ;
        RECT 444.005 -5.660 444.235 -4.990 ;
        RECT 446.145 -5.660 446.375 -4.990 ;
        RECT 448.385 -5.660 448.615 -4.990 ;
        RECT 450.625 -5.660 450.855 -4.990 ;
      LAYER Via1 ;
        RECT 448.390 -4.930 448.650 -4.670 ;
      LAYER Metal2 ;
        RECT 448.380 -5.130 448.660 -4.610 ;
      LAYER Via2 ;
        RECT 448.380 -4.940 448.660 -4.660 ;
      LAYER Metal3 ;
        RECT 465.200 -4.100 654.000 -3.960 ;
        RECT 448.660 -4.380 654.000 -4.100 ;
        RECT 448.660 -4.660 448.940 -4.380 ;
        RECT 465.200 -4.520 654.000 -4.380 ;
        RECT 448.330 -4.940 448.940 -4.660 ;
    END
  END result[1]
  PIN result[0]
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 452.405 -15.250 452.635 -14.580 ;
        RECT 454.545 -15.250 454.775 -14.580 ;
        RECT 456.785 -14.750 457.015 -14.580 ;
        RECT 456.730 -15.010 457.110 -14.750 ;
        RECT 456.785 -15.250 457.015 -15.010 ;
        RECT 459.025 -15.250 459.255 -14.580 ;
        RECT 452.405 -15.630 459.255 -15.250 ;
        RECT 455.400 -16.540 456.200 -15.630 ;
        RECT 452.405 -16.920 459.355 -16.540 ;
        RECT 452.405 -17.285 452.665 -16.920 ;
        RECT 454.645 -17.285 454.875 -16.920 ;
        RECT 456.885 -17.285 457.115 -16.920 ;
        RECT 459.125 -17.285 459.355 -16.920 ;
      LAYER Via1 ;
        RECT 456.790 -15.010 457.050 -14.750 ;
      LAYER Metal2 ;
        RECT 456.780 -15.070 457.060 -11.890 ;
      LAYER Via2 ;
        RECT 456.780 -12.220 457.060 -11.940 ;
      LAYER Metal3 ;
        RECT 465.200 -11.940 654.000 -11.800 ;
        RECT 456.730 -12.220 654.000 -11.940 ;
        RECT 465.200 -12.360 654.000 -12.220 ;
    END
  END result[0]
  PIN valid
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 444.005 -26.840 444.265 -26.475 ;
        RECT 446.245 -26.840 446.475 -26.475 ;
        RECT 448.485 -26.840 448.715 -26.475 ;
        RECT 450.725 -26.840 450.955 -26.475 ;
        RECT 444.005 -27.220 450.955 -26.840 ;
        RECT 447.000 -28.130 447.800 -27.220 ;
        RECT 444.005 -28.510 450.855 -28.130 ;
        RECT 444.005 -29.180 444.235 -28.510 ;
        RECT 446.145 -29.180 446.375 -28.510 ;
        RECT 448.385 -29.180 448.615 -28.510 ;
        RECT 450.625 -29.180 450.855 -28.510 ;
      LAYER Via1 ;
        RECT 448.390 -28.450 448.650 -28.190 ;
      LAYER Metal2 ;
        RECT 448.380 -28.510 448.660 -27.570 ;
      LAYER Via2 ;
        RECT 448.380 -27.900 448.660 -27.620 ;
      LAYER Metal3 ;
        RECT 465.200 -27.620 654.000 -27.480 ;
        RECT 448.330 -27.900 654.000 -27.620 ;
        RECT 465.200 -28.040 654.000 -27.900 ;
    END
  END valid
  PIN cal
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal1 ;
        RECT 452.245 -44.190 452.580 -42.290 ;
        RECT 460.040 -43.220 460.415 -42.515 ;
        RECT 459.530 -43.630 460.415 -43.220 ;
      LAYER Via1 ;
        RECT 452.310 -43.570 452.570 -43.310 ;
        RECT 459.590 -43.570 459.850 -43.310 ;
      LAYER Metal2 ;
        RECT 452.300 -43.770 452.580 -43.250 ;
        RECT 459.580 -43.770 459.860 -35.410 ;
      LAYER Via2 ;
        RECT 459.580 -35.740 459.860 -35.460 ;
        RECT 452.300 -43.580 452.580 -43.300 ;
        RECT 459.580 -43.580 459.860 -43.300 ;
      LAYER Metal3 ;
        RECT 465.200 -35.460 654.000 -35.320 ;
        RECT 459.530 -35.740 654.000 -35.460 ;
        RECT 465.200 -35.880 654.000 -35.740 ;
        RECT 452.250 -43.580 459.910 -43.300 ;
    END
  END cal
  PIN en
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal1 ;
        RECT 456.165 -28.510 456.500 -26.610 ;
        RECT 459.470 -39.855 460.415 -39.330 ;
        RECT 460.105 -40.870 460.415 -39.855 ;
      LAYER Via1 ;
        RECT 456.230 -28.450 456.490 -28.190 ;
        RECT 460.150 -39.650 460.410 -39.390 ;
      LAYER Metal2 ;
        RECT 456.220 -28.180 456.500 -28.130 ;
        RECT 455.660 -28.460 456.500 -28.180 ;
        RECT 455.660 -39.710 455.940 -28.460 ;
        RECT 456.220 -28.510 456.500 -28.460 ;
        RECT 460.140 -39.380 460.420 -39.330 ;
        RECT 460.140 -39.660 460.980 -39.380 ;
        RECT 460.140 -39.850 460.420 -39.660 ;
        RECT 460.700 -43.630 460.980 -39.660 ;
      LAYER Via2 ;
        RECT 455.660 -39.660 455.940 -39.380 ;
        RECT 460.700 -43.580 460.980 -43.300 ;
      LAYER Metal3 ;
        RECT 455.610 -39.660 460.470 -39.380 ;
        RECT 465.200 -43.300 654.000 -43.160 ;
        RECT 460.650 -43.580 654.000 -43.300 ;
        RECT 465.200 -43.720 654.000 -43.580 ;
    END
  END en
  PIN clk
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal1 ;
        RECT 451.685 -48.510 452.020 -46.610 ;
        RECT 459.530 -47.580 460.415 -47.170 ;
        RECT 460.040 -48.285 460.415 -47.580 ;
      LAYER Via1 ;
        RECT 451.750 -48.050 452.010 -47.790 ;
        RECT 460.150 -48.050 460.410 -47.790 ;
      LAYER Metal2 ;
        RECT 451.740 -48.250 452.020 -47.730 ;
        RECT 460.140 -51.470 460.420 -47.730 ;
      LAYER Via2 ;
        RECT 451.740 -48.060 452.020 -47.780 ;
        RECT 460.140 -48.060 460.420 -47.780 ;
        RECT 460.140 -51.420 460.420 -51.140 ;
      LAYER Metal3 ;
        RECT 451.690 -48.060 460.470 -47.780 ;
        RECT 465.200 -51.140 654.000 -51.000 ;
        RECT 460.090 -51.420 654.000 -51.140 ;
        RECT 465.200 -51.560 654.000 -51.420 ;
    END
  END clk
  PIN rstn
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal1 ;
        RECT 447.765 -48.510 448.100 -46.610 ;
        RECT 455.105 -47.580 455.990 -47.170 ;
        RECT 455.105 -48.285 455.480 -47.580 ;
      LAYER Via1 ;
        RECT 447.830 -47.490 448.090 -47.230 ;
        RECT 455.670 -47.490 455.930 -47.230 ;
      LAYER Metal2 ;
        RECT 447.820 -47.690 448.100 -47.170 ;
        RECT 455.660 -59.310 455.940 -47.170 ;
      LAYER Via2 ;
        RECT 447.820 -47.500 448.100 -47.220 ;
        RECT 455.660 -47.500 455.940 -47.220 ;
        RECT 455.660 -59.260 455.940 -58.980 ;
      LAYER Metal3 ;
        RECT 447.770 -47.500 455.990 -47.220 ;
        RECT 465.200 -58.980 654.000 -58.840 ;
        RECT 455.610 -59.260 654.000 -58.980 ;
        RECT 465.200 -59.400 654.000 -59.260 ;
    END
  END rstn
  PIN vinp
    ANTENNADIFFAREA 1.040000 ;
    PORT
      LAYER Metal1 ;
        RECT -497.005 82.660 -496.105 82.735 ;
        RECT -497.005 82.430 -492.560 82.660 ;
        RECT -497.005 82.355 -496.105 82.430 ;
      LAYER Via1 ;
        RECT -496.945 82.415 -496.165 82.675 ;
      LAYER Metal2 ;
        RECT -507.300 82.735 -504.300 83.340 ;
        RECT -507.300 82.355 -496.105 82.735 ;
        RECT -507.300 81.740 -504.300 82.355 ;
      LAYER Via2 ;
        RECT -506.980 81.880 -504.620 83.200 ;
      LAYER Metal3 ;
        RECT -877.500 81.740 -504.300 83.340 ;
    END
  END vinp
  PIN vinn
    ANTENNADIFFAREA 1.040000 ;
    PORT
      LAYER Metal1 ;
        RECT -497.005 -82.430 -496.105 -82.355 ;
        RECT -497.005 -82.660 -492.560 -82.430 ;
        RECT -497.005 -82.735 -496.105 -82.660 ;
      LAYER Via1 ;
        RECT -496.945 -82.675 -496.165 -82.415 ;
      LAYER Metal2 ;
        RECT -507.300 -82.345 -504.300 -81.740 ;
        RECT -507.300 -82.725 -496.105 -82.345 ;
        RECT -507.300 -83.340 -504.300 -82.725 ;
        RECT -498.105 -82.735 -496.105 -82.725 ;
      LAYER Via2 ;
        RECT -506.980 -83.200 -504.620 -81.880 ;
      LAYER Metal3 ;
        RECT -877.500 -83.340 -504.300 -81.740 ;
    END
  END vinn
  OBS
      LAYER Nwell ;
        RECT -490.535 83.595 -486.455 87.615 ;
        RECT 233.175 -2.120 236.275 11.560 ;
        RECT 229.550 -8.550 232.330 -5.450 ;
        RECT 233.065 -8.550 235.845 -5.450 ;
        RECT -490.535 -87.615 -486.455 -83.595 ;
      LAYER Metal1 ;
        RECT 144.285 98.450 145.745 98.750 ;
        RECT -491.830 96.285 -491.430 98.115 ;
        RECT 144.285 97.740 144.605 98.450 ;
        RECT 143.575 97.290 144.605 97.740 ;
        RECT 145.490 97.695 145.745 98.450 ;
        RECT 145.490 97.465 146.435 97.695 ;
        RECT -492.345 95.945 -489.675 96.285 ;
        RECT -491.830 95.830 -491.430 95.945 ;
        RECT -493.475 95.450 -492.575 95.830 ;
        RECT -489.445 95.450 -488.545 95.830 ;
        RECT 144.285 95.090 145.745 95.390 ;
        RECT 144.285 94.380 144.605 95.090 ;
        RECT 143.575 93.930 144.605 94.380 ;
        RECT 144.845 93.340 145.260 94.860 ;
        RECT 145.490 94.335 145.745 95.090 ;
        RECT 145.490 94.105 146.435 94.335 ;
        RECT 144.285 91.730 145.745 92.030 ;
        RECT 144.285 91.020 144.605 91.730 ;
        RECT 143.575 90.570 144.605 91.020 ;
        RECT 144.845 89.980 145.260 91.500 ;
        RECT 145.490 90.975 145.745 91.730 ;
        RECT 145.490 90.745 146.435 90.975 ;
        RECT 144.285 88.370 145.745 88.670 ;
        RECT 144.285 87.660 144.605 88.370 ;
        RECT -494.430 86.965 -487.560 87.265 ;
        RECT 143.575 87.210 144.605 87.660 ;
        RECT -494.430 86.510 -492.560 86.965 ;
        RECT -494.430 85.490 -492.560 85.720 ;
        RECT -492.330 84.775 -492.100 85.335 ;
        RECT -492.330 84.395 -491.430 84.775 ;
        RECT -492.330 83.835 -492.100 84.395 ;
        RECT -497.595 83.680 -495.515 83.765 ;
        RECT -497.595 83.450 -492.560 83.680 ;
        RECT -497.595 83.365 -495.515 83.450 ;
        RECT -492.330 82.660 -492.100 83.295 ;
        RECT -491.110 82.660 -490.880 86.965 ;
        RECT -490.615 86.355 -490.235 86.565 ;
        RECT -489.430 86.510 -487.560 86.965 ;
        RECT -490.615 85.875 -489.660 86.355 ;
        RECT -490.615 85.665 -490.235 85.875 ;
        RECT -486.870 85.720 -486.640 87.105 ;
        RECT 144.845 86.620 145.260 88.140 ;
        RECT 145.490 87.615 145.745 88.370 ;
        RECT 145.490 87.385 146.435 87.615 ;
        RECT -489.430 85.490 -486.640 85.720 ;
        RECT -489.890 82.660 -489.660 85.335 ;
        RECT -486.870 83.235 -486.640 85.490 ;
        RECT 144.285 85.010 145.745 85.310 ;
        RECT 144.285 84.300 144.605 85.010 ;
        RECT 143.575 83.850 144.605 84.300 ;
        RECT 144.845 83.260 145.260 84.780 ;
        RECT 145.490 84.255 145.745 85.010 ;
        RECT 145.490 84.025 146.435 84.255 ;
        RECT -492.330 82.430 -489.660 82.660 ;
        RECT -492.330 81.795 -492.100 82.430 ;
        RECT -494.430 79.615 -492.560 81.640 ;
        RECT -486.955 81.155 -486.555 83.235 ;
        RECT 144.285 81.650 145.745 81.950 ;
        RECT 144.285 80.940 144.605 81.650 ;
        RECT 143.575 80.490 144.605 80.940 ;
        RECT 144.845 79.900 145.260 81.420 ;
        RECT 145.490 80.895 145.745 81.650 ;
        RECT 145.490 80.665 146.435 80.895 ;
        RECT -484.745 79.615 -483.845 79.655 ;
        RECT -494.430 79.315 -483.845 79.615 ;
        RECT -484.745 79.275 -483.845 79.315 ;
        RECT 144.285 78.290 145.745 78.590 ;
        RECT 144.285 77.580 144.605 78.290 ;
        RECT 143.575 77.130 144.605 77.580 ;
        RECT 144.845 76.540 145.260 78.060 ;
        RECT 145.490 77.535 145.745 78.290 ;
        RECT 145.490 77.305 146.435 77.535 ;
        RECT 144.285 74.930 145.745 75.230 ;
        RECT 144.285 74.220 144.605 74.930 ;
        RECT 143.575 73.770 144.605 74.220 ;
        RECT 144.845 73.180 145.260 74.700 ;
        RECT 145.490 74.175 145.745 74.930 ;
        RECT 145.490 73.945 146.435 74.175 ;
        RECT 144.285 71.570 145.745 71.870 ;
        RECT 144.285 70.860 144.605 71.570 ;
        RECT 143.575 70.410 144.605 70.860 ;
        RECT 144.845 69.820 145.260 71.340 ;
        RECT 145.490 70.815 145.745 71.570 ;
        RECT 145.490 70.585 146.435 70.815 ;
        RECT 144.285 68.210 145.745 68.510 ;
        RECT 144.285 67.500 144.605 68.210 ;
        RECT 143.575 67.050 144.605 67.500 ;
        RECT 144.845 66.460 145.260 67.980 ;
        RECT 145.490 67.455 145.745 68.210 ;
        RECT 145.490 67.225 146.435 67.455 ;
        RECT 144.285 64.850 145.745 65.150 ;
        RECT 144.285 64.140 144.605 64.850 ;
        RECT 143.575 63.690 144.605 64.140 ;
        RECT 144.845 63.100 145.260 64.620 ;
        RECT 145.490 64.095 145.745 64.850 ;
        RECT 145.490 63.865 146.435 64.095 ;
        RECT 300.585 48.030 300.815 48.140 ;
        RECT 300.550 47.650 300.815 48.030 ;
        RECT 300.585 47.470 300.815 47.650 ;
        RECT 302.825 47.470 303.055 48.140 ;
        RECT 305.065 47.470 305.295 48.140 ;
        RECT 307.205 47.470 307.435 48.140 ;
        RECT 309.545 47.520 309.775 48.140 ;
        RECT 311.785 47.520 312.015 48.140 ;
        RECT 300.585 47.090 307.435 47.470 ;
        RECT 308.965 47.290 312.015 47.520 ;
        RECT 317.905 47.520 318.135 48.140 ;
        RECT 320.145 47.520 320.375 48.140 ;
        RECT 322.485 48.030 322.715 48.140 ;
        RECT 322.390 47.650 322.715 48.030 ;
        RECT 317.905 47.290 320.955 47.520 ;
        RECT 299.740 46.445 302.940 46.790 ;
        RECT 303.640 46.180 304.440 47.090 ;
        RECT 308.965 46.785 309.300 47.290 ;
        RECT 305.010 46.445 309.300 46.785 ;
        RECT 309.770 46.475 312.630 46.910 ;
        RECT 317.290 46.475 320.150 46.910 ;
        RECT 320.620 46.785 320.955 47.290 ;
        RECT 322.485 47.470 322.715 47.650 ;
        RECT 324.625 47.470 324.855 48.140 ;
        RECT 326.865 47.470 327.095 48.140 ;
        RECT 329.105 47.470 329.335 48.140 ;
        RECT 322.485 47.090 329.335 47.470 ;
        RECT 300.485 45.800 307.435 46.180 ;
        RECT 300.485 45.435 300.715 45.800 ;
        RECT 302.725 45.435 302.955 45.800 ;
        RECT 304.965 45.435 305.195 45.800 ;
        RECT 307.175 45.435 307.435 45.800 ;
        RECT 308.965 46.010 309.300 46.445 ;
        RECT 320.620 46.445 324.910 46.785 ;
        RECT 320.620 46.010 320.955 46.445 ;
        RECT 325.480 46.180 326.280 47.090 ;
        RECT 326.980 46.445 330.180 46.790 ;
        RECT 331.445 46.315 331.675 48.150 ;
        RECT 336.985 48.030 337.215 48.140 ;
        RECT 336.950 47.650 337.215 48.030 ;
        RECT 336.985 47.470 337.215 47.650 ;
        RECT 339.225 47.470 339.455 48.140 ;
        RECT 341.465 47.470 341.695 48.140 ;
        RECT 343.605 47.470 343.835 48.140 ;
        RECT 345.945 47.520 346.175 48.140 ;
        RECT 348.185 47.520 348.415 48.140 ;
        RECT 336.985 47.090 343.835 47.470 ;
        RECT 345.365 47.290 348.415 47.520 ;
        RECT 331.930 46.720 333.195 46.950 ;
        RECT 308.965 45.775 311.915 46.010 ;
        RECT 309.445 45.435 309.675 45.775 ;
        RECT 311.685 45.435 311.915 45.775 ;
        RECT 318.005 45.775 320.955 46.010 ;
        RECT 322.485 45.800 329.435 46.180 ;
        RECT 331.445 46.085 332.720 46.315 ;
        RECT 318.005 45.435 318.235 45.775 ;
        RECT 320.245 45.435 320.475 45.775 ;
        RECT 322.485 45.435 322.745 45.800 ;
        RECT 324.725 45.435 324.955 45.800 ;
        RECT 326.965 45.435 327.195 45.800 ;
        RECT 329.205 45.435 329.435 45.800 ;
        RECT 332.965 45.290 333.195 46.720 ;
        RECT 336.140 46.445 339.340 46.790 ;
        RECT 340.040 46.180 340.840 47.090 ;
        RECT 345.365 46.785 345.700 47.290 ;
        RECT 341.410 46.445 345.700 46.785 ;
        RECT 346.170 46.475 349.030 46.910 ;
        RECT 336.885 45.800 343.835 46.180 ;
        RECT 336.885 45.435 337.115 45.800 ;
        RECT 339.125 45.435 339.355 45.800 ;
        RECT 341.365 45.435 341.595 45.800 ;
        RECT 343.575 45.435 343.835 45.800 ;
        RECT 345.365 46.010 345.700 46.445 ;
        RECT 349.925 46.315 350.155 48.150 ;
        RECT 355.425 47.520 355.655 48.140 ;
        RECT 357.665 47.520 357.895 48.140 ;
        RECT 360.005 48.030 360.235 48.140 ;
        RECT 359.910 47.650 360.235 48.030 ;
        RECT 355.425 47.290 358.475 47.520 ;
        RECT 350.410 46.720 351.675 46.950 ;
        RECT 349.925 46.085 351.200 46.315 ;
        RECT 345.365 45.775 348.315 46.010 ;
        RECT 345.845 45.435 346.075 45.775 ;
        RECT 348.085 45.435 348.315 45.775 ;
        RECT 351.445 45.290 351.675 46.720 ;
        RECT 354.810 46.475 357.670 46.910 ;
        RECT 358.140 46.785 358.475 47.290 ;
        RECT 360.005 47.470 360.235 47.650 ;
        RECT 362.145 47.470 362.375 48.140 ;
        RECT 364.385 47.470 364.615 48.140 ;
        RECT 366.625 47.470 366.855 48.140 ;
        RECT 360.005 47.090 366.855 47.470 ;
        RECT 358.140 46.445 362.430 46.785 ;
        RECT 358.140 46.010 358.475 46.445 ;
        RECT 363.000 46.180 363.800 47.090 ;
        RECT 364.500 46.445 367.700 46.790 ;
        RECT 368.965 46.315 369.195 48.150 ;
        RECT 375.065 48.030 375.295 48.140 ;
        RECT 375.030 47.650 375.295 48.030 ;
        RECT 375.065 47.470 375.295 47.650 ;
        RECT 377.305 47.470 377.535 48.140 ;
        RECT 379.545 47.470 379.775 48.140 ;
        RECT 381.685 47.470 381.915 48.140 ;
        RECT 384.025 47.520 384.255 48.140 ;
        RECT 386.265 47.520 386.495 48.140 ;
        RECT 394.105 48.030 394.335 48.140 ;
        RECT 394.070 47.650 394.335 48.030 ;
        RECT 375.065 47.090 381.915 47.470 ;
        RECT 383.445 47.290 386.495 47.520 ;
        RECT 394.105 47.470 394.335 47.650 ;
        RECT 396.345 47.470 396.575 48.140 ;
        RECT 398.585 47.470 398.815 48.140 ;
        RECT 400.725 47.470 400.955 48.140 ;
        RECT 403.065 47.520 403.295 48.140 ;
        RECT 405.305 47.520 405.535 48.140 ;
        RECT 369.450 46.720 370.715 46.950 ;
        RECT 355.525 45.775 358.475 46.010 ;
        RECT 360.005 45.800 366.955 46.180 ;
        RECT 368.965 46.085 370.240 46.315 ;
        RECT 355.525 45.435 355.755 45.775 ;
        RECT 357.765 45.435 357.995 45.775 ;
        RECT 360.005 45.435 360.265 45.800 ;
        RECT 362.245 45.435 362.475 45.800 ;
        RECT 364.485 45.435 364.715 45.800 ;
        RECT 366.725 45.435 366.955 45.800 ;
        RECT 370.485 45.290 370.715 46.720 ;
        RECT 374.220 46.445 377.420 46.790 ;
        RECT 378.120 46.180 378.920 47.090 ;
        RECT 383.445 46.785 383.780 47.290 ;
        RECT 379.490 46.445 383.780 46.785 ;
        RECT 384.250 46.475 387.110 46.910 ;
        RECT 374.965 45.800 381.915 46.180 ;
        RECT 374.965 45.435 375.195 45.800 ;
        RECT 377.205 45.435 377.435 45.800 ;
        RECT 379.445 45.435 379.675 45.800 ;
        RECT 381.655 45.435 381.915 45.800 ;
        RECT 383.445 46.010 383.780 46.445 ;
        RECT 383.445 45.775 386.395 46.010 ;
        RECT 383.925 45.435 384.155 45.775 ;
        RECT 386.165 45.435 386.395 45.775 ;
        RECT 389.020 45.570 389.355 47.470 ;
        RECT 394.105 47.090 400.955 47.470 ;
        RECT 402.485 47.290 405.535 47.520 ;
        RECT 412.545 47.520 412.775 48.140 ;
        RECT 414.785 47.520 415.015 48.140 ;
        RECT 417.125 48.030 417.355 48.140 ;
        RECT 417.030 47.650 417.355 48.030 ;
        RECT 393.260 46.445 396.460 46.790 ;
        RECT 397.160 46.180 397.960 47.090 ;
        RECT 402.485 46.785 402.820 47.290 ;
        RECT 398.530 46.445 402.820 46.785 ;
        RECT 403.290 46.475 406.150 46.910 ;
        RECT 394.005 45.800 400.955 46.180 ;
        RECT 389.030 45.410 389.290 45.570 ;
        RECT 394.005 45.435 394.235 45.800 ;
        RECT 396.245 45.435 396.475 45.800 ;
        RECT 398.485 45.435 398.715 45.800 ;
        RECT 400.695 45.435 400.955 45.800 ;
        RECT 402.485 46.010 402.820 46.445 ;
        RECT 402.485 45.775 405.435 46.010 ;
        RECT 402.965 45.435 403.195 45.775 ;
        RECT 405.205 45.435 405.435 45.775 ;
        RECT 408.060 45.570 408.395 47.470 ;
        RECT 412.545 47.290 415.595 47.520 ;
        RECT 411.930 46.475 414.790 46.910 ;
        RECT 415.260 46.785 415.595 47.290 ;
        RECT 417.125 47.470 417.355 47.650 ;
        RECT 419.265 47.470 419.495 48.140 ;
        RECT 421.505 47.470 421.735 48.140 ;
        RECT 423.745 47.470 423.975 48.140 ;
        RECT 417.125 47.090 423.975 47.470 ;
        RECT 415.260 46.445 419.550 46.785 ;
        RECT 415.260 46.010 415.595 46.445 ;
        RECT 420.120 46.180 420.920 47.090 ;
        RECT 421.620 46.445 424.820 46.790 ;
        RECT 412.645 45.775 415.595 46.010 ;
        RECT 417.125 45.800 424.075 46.180 ;
        RECT 426.545 45.940 426.850 48.080 ;
        RECT 428.225 47.440 428.505 48.140 ;
        RECT 432.185 48.030 432.415 48.140 ;
        RECT 432.150 47.650 432.415 48.030 ;
        RECT 427.080 47.120 428.505 47.440 ;
        RECT 432.185 47.470 432.415 47.650 ;
        RECT 434.425 47.470 434.655 48.140 ;
        RECT 436.665 47.470 436.895 48.140 ;
        RECT 438.805 47.470 439.035 48.140 ;
        RECT 441.145 47.520 441.375 48.140 ;
        RECT 443.385 47.520 443.615 48.140 ;
        RECT 408.070 45.410 408.330 45.570 ;
        RECT 412.645 45.435 412.875 45.775 ;
        RECT 414.885 45.435 415.115 45.775 ;
        RECT 417.125 45.435 417.385 45.800 ;
        RECT 419.365 45.435 419.595 45.800 ;
        RECT 421.605 45.435 421.835 45.800 ;
        RECT 423.845 45.435 424.075 45.800 ;
        RECT 427.080 45.360 427.435 47.120 ;
        RECT 432.185 47.090 439.035 47.470 ;
        RECT 440.565 47.290 443.615 47.520 ;
        RECT 427.665 46.550 428.695 46.890 ;
        RECT 427.665 45.360 427.970 46.550 ;
        RECT 431.340 46.445 434.540 46.790 ;
        RECT 435.240 46.180 436.040 47.090 ;
        RECT 440.565 46.785 440.900 47.290 ;
        RECT 436.610 46.445 440.900 46.785 ;
        RECT 441.370 46.475 444.230 46.910 ;
        RECT 432.085 45.800 439.035 46.180 ;
        RECT 432.085 45.435 432.315 45.800 ;
        RECT 434.325 45.435 434.555 45.800 ;
        RECT 436.565 45.435 436.795 45.800 ;
        RECT 438.775 45.435 439.035 45.800 ;
        RECT 440.565 46.010 440.900 46.445 ;
        RECT 440.565 45.775 443.515 46.010 ;
        RECT 441.045 45.435 441.275 45.775 ;
        RECT 443.285 45.435 443.515 45.775 ;
        RECT 446.140 45.570 446.475 47.470 ;
        RECT 449.605 46.315 449.835 48.150 ;
        RECT 450.090 46.720 451.355 46.950 ;
        RECT 449.605 46.085 450.880 46.315 ;
        RECT 446.150 45.410 446.410 45.570 ;
        RECT 451.125 45.290 451.355 46.720 ;
        RECT 451.845 46.315 452.075 48.150 ;
        RECT 452.330 46.720 453.595 46.950 ;
        RECT 451.845 46.085 453.120 46.315 ;
        RECT 453.365 45.290 453.595 46.720 ;
        RECT 454.085 46.315 454.315 48.150 ;
        RECT 454.570 46.720 455.835 46.950 ;
        RECT 454.085 46.085 455.360 46.315 ;
        RECT 455.605 45.290 455.835 46.720 ;
        RECT 456.325 46.315 456.555 48.150 ;
        RECT 456.810 46.720 458.075 46.950 ;
        RECT 456.325 46.085 457.600 46.315 ;
        RECT 457.845 45.290 458.075 46.720 ;
        RECT 458.565 46.315 458.795 48.150 ;
        RECT 459.050 46.720 460.315 46.950 ;
        RECT 458.565 46.085 459.840 46.315 ;
        RECT 460.085 45.290 460.315 46.720 ;
        RECT 298.805 43.720 299.035 44.085 ;
        RECT 301.045 43.720 301.275 44.085 ;
        RECT 303.285 43.720 303.515 44.085 ;
        RECT 305.495 43.720 305.755 44.085 ;
        RECT 307.765 43.745 307.995 44.085 ;
        RECT 310.005 43.745 310.235 44.085 ;
        RECT 298.805 43.340 305.755 43.720 ;
        RECT 307.285 43.510 310.235 43.745 ;
        RECT 298.060 42.730 301.260 43.075 ;
        RECT 301.960 42.430 302.760 43.340 ;
        RECT 307.285 43.075 307.620 43.510 ;
        RECT 303.330 42.735 307.620 43.075 ;
        RECT 298.870 42.050 305.755 42.430 ;
        RECT 298.905 41.380 299.135 42.050 ;
        RECT 301.145 41.380 301.375 42.050 ;
        RECT 303.385 41.380 303.615 42.050 ;
        RECT 305.525 41.380 305.755 42.050 ;
        RECT 307.285 42.230 307.620 42.735 ;
        RECT 308.090 42.610 310.950 43.045 ;
        RECT 307.285 42.000 310.335 42.230 ;
        RECT 307.865 41.380 308.095 42.000 ;
        RECT 310.105 41.380 310.335 42.000 ;
        RECT 312.245 41.390 312.580 44.160 ;
        RECT 312.810 41.810 313.135 43.790 ;
        RECT 314.485 41.390 314.820 44.160 ;
        RECT 315.050 41.810 315.375 43.790 ;
        RECT 317.340 42.050 317.675 43.950 ;
        RECT 319.580 42.050 319.915 43.950 ;
        RECT 320.805 43.205 322.080 43.435 ;
        RECT 320.805 41.370 321.035 43.205 ;
        RECT 322.325 42.800 322.555 44.230 ;
        RECT 321.290 42.570 322.555 42.800 ;
        RECT 323.045 43.205 324.320 43.435 ;
        RECT 323.045 41.370 323.275 43.205 ;
        RECT 324.565 42.800 324.795 44.230 ;
        RECT 323.530 42.570 324.795 42.800 ;
        RECT 325.285 43.205 326.560 43.435 ;
        RECT 325.285 41.370 325.515 43.205 ;
        RECT 326.805 42.800 327.035 44.230 ;
        RECT 325.770 42.570 327.035 42.800 ;
        RECT 327.525 43.205 328.800 43.435 ;
        RECT 327.525 41.370 327.755 43.205 ;
        RECT 329.045 42.800 329.275 44.230 ;
        RECT 328.010 42.570 329.275 42.800 ;
        RECT 329.765 43.205 331.040 43.435 ;
        RECT 329.765 41.370 329.995 43.205 ;
        RECT 331.285 42.800 331.515 44.230 ;
        RECT 330.250 42.570 331.515 42.800 ;
        RECT 333.525 41.370 333.855 44.230 ;
        RECT 334.085 42.560 334.410 43.560 ;
        RECT 338.020 41.880 338.440 43.685 ;
        RECT 338.670 43.480 339.065 44.230 ;
        RECT 340.725 43.720 341.490 44.150 ;
        RECT 338.670 43.250 340.895 43.480 ;
        RECT 338.670 41.630 338.900 43.250 ;
        RECT 340.040 43.120 340.895 43.250 ;
        RECT 337.695 41.400 338.900 41.630 ;
        RECT 339.140 41.415 339.500 43.020 ;
        RECT 341.160 42.470 341.490 43.720 ;
        RECT 340.860 41.415 341.490 42.470 ;
        RECT 342.085 42.180 342.315 43.960 ;
        RECT 342.545 43.130 343.060 44.110 ;
        RECT 344.170 43.160 344.795 44.185 ;
        RECT 342.545 42.570 343.430 43.130 ;
        RECT 343.810 42.180 344.095 42.930 ;
        RECT 342.085 41.945 344.095 42.180 ;
        RECT 342.085 41.370 342.470 41.945 ;
        RECT 344.325 41.380 344.795 43.160 ;
        RECT 345.445 43.205 346.720 43.435 ;
        RECT 345.445 41.370 345.675 43.205 ;
        RECT 346.965 42.800 347.195 44.230 ;
        RECT 345.930 42.570 347.195 42.800 ;
        RECT 349.830 42.560 350.155 43.560 ;
        RECT 350.385 41.370 350.715 44.230 ;
        RECT 351.765 43.160 352.390 44.185 ;
        RECT 351.765 41.380 352.235 43.160 ;
        RECT 353.500 43.130 354.015 44.110 ;
        RECT 364.280 44.000 367.630 44.230 ;
        RECT 352.465 42.180 352.750 42.930 ;
        RECT 353.130 42.570 354.015 43.130 ;
        RECT 354.245 42.180 354.475 43.960 ;
        RECT 355.525 43.480 355.755 43.950 ;
        RECT 357.545 43.665 358.050 43.895 ;
        RECT 359.505 43.685 359.910 43.915 ;
        RECT 355.525 43.250 357.315 43.480 ;
        RECT 355.430 42.610 356.850 42.990 ;
        RECT 357.085 42.355 357.315 43.250 ;
        RECT 352.465 41.945 354.475 42.180 ;
        RECT 354.090 41.370 354.475 41.945 ;
        RECT 355.625 42.125 357.315 42.355 ;
        RECT 357.545 42.375 357.775 43.665 ;
        RECT 358.170 42.610 359.200 42.990 ;
        RECT 357.545 42.145 359.175 42.375 ;
        RECT 359.505 42.340 359.735 43.685 ;
        RECT 355.625 41.535 355.855 42.125 ;
        RECT 357.545 41.545 357.895 42.145 ;
        RECT 358.945 41.770 359.175 42.145 ;
        RECT 359.405 42.000 359.735 42.340 ;
        RECT 359.965 41.770 360.195 42.850 ;
        RECT 360.745 42.690 360.975 43.970 ;
        RECT 364.280 43.610 364.510 44.000 ;
        RECT 361.325 43.380 364.510 43.610 ;
        RECT 361.325 43.170 361.555 43.380 ;
        RECT 365.270 43.150 365.610 43.760 ;
        RECT 366.205 43.170 366.435 44.000 ;
        RECT 361.970 42.920 365.950 43.150 ;
        RECT 360.425 42.460 365.435 42.690 ;
        RECT 360.425 42.000 360.655 42.460 ;
        RECT 365.135 42.235 365.435 42.460 ;
        RECT 361.445 42.000 364.275 42.230 ;
        RECT 361.445 41.805 361.675 42.000 ;
        RECT 358.945 41.540 360.195 41.770 ;
        RECT 364.045 41.630 364.275 42.000 ;
        RECT 365.720 41.915 365.950 42.920 ;
        RECT 366.830 42.940 367.170 43.760 ;
        RECT 367.400 43.400 367.630 44.000 ;
        RECT 368.230 43.630 369.035 43.970 ;
        RECT 367.400 43.170 368.400 43.400 ;
        RECT 366.830 42.710 367.720 42.940 ;
        RECT 365.720 41.685 366.360 41.915 ;
        RECT 367.490 41.600 367.720 42.710 ;
        RECT 368.170 42.235 368.400 43.170 ;
        RECT 368.695 41.830 369.035 43.630 ;
        RECT 369.940 43.740 371.575 44.100 ;
        RECT 369.940 42.930 370.485 43.740 ;
        RECT 371.930 43.310 372.160 43.970 ;
        RECT 371.010 43.080 373.510 43.310 ;
        RECT 371.010 42.585 371.240 43.080 ;
        RECT 369.275 42.355 371.240 42.585 ;
        RECT 369.475 41.710 370.745 41.940 ;
        RECT 371.010 41.830 371.240 42.355 ;
        RECT 369.475 41.600 369.705 41.710 ;
        RECT 367.490 41.370 369.705 41.600 ;
        RECT 370.515 41.600 370.745 41.710 ;
        RECT 371.470 41.600 371.700 42.850 ;
        RECT 370.515 41.370 371.700 41.600 ;
        RECT 373.755 41.380 374.190 44.210 ;
        RECT 375.790 43.720 376.555 44.150 ;
        RECT 375.790 42.470 376.120 43.720 ;
        RECT 378.215 43.480 378.610 44.230 ;
        RECT 376.385 43.250 378.610 43.480 ;
        RECT 376.385 43.120 377.240 43.250 ;
        RECT 375.790 41.415 376.420 42.470 ;
        RECT 377.780 41.415 378.140 43.020 ;
        RECT 378.380 41.630 378.610 43.250 ;
        RECT 378.840 41.880 379.260 43.685 ;
        RECT 382.065 43.480 382.295 43.960 ;
        RECT 381.150 43.250 382.295 43.480 ;
        RECT 381.150 42.400 381.490 43.250 ;
        RECT 383.880 43.020 384.255 44.210 ;
        RECT 381.750 42.720 383.070 43.020 ;
        RECT 381.150 42.050 382.295 42.400 ;
        RECT 378.380 41.400 379.585 41.630 ;
        RECT 382.065 41.370 382.295 42.050 ;
        RECT 382.745 42.170 383.070 42.720 ;
        RECT 383.310 42.610 384.255 43.020 ;
        RECT 384.485 42.170 384.715 43.955 ;
        RECT 385.570 42.990 385.965 43.675 ;
        RECT 385.570 42.610 386.530 42.990 ;
        RECT 386.760 42.610 387.080 44.210 ;
        RECT 387.310 42.380 387.640 44.175 ;
        RECT 387.880 42.610 388.200 44.210 ;
        RECT 388.440 42.960 388.760 44.210 ;
        RECT 388.440 42.610 389.505 42.960 ;
        RECT 382.745 41.940 384.715 42.170 ;
        RECT 384.485 41.370 384.715 41.940 ;
        RECT 385.215 42.000 387.010 42.230 ;
        RECT 387.310 42.050 388.850 42.380 ;
        RECT 385.215 41.380 385.555 42.000 ;
        RECT 386.780 41.615 387.010 42.000 ;
        RECT 389.295 41.615 389.635 42.230 ;
        RECT 391.825 41.810 392.150 43.790 ;
        RECT 386.780 41.380 389.635 41.615 ;
        RECT 392.380 41.390 392.715 44.160 ;
        RECT 402.920 44.000 406.270 44.230 ;
        RECT 394.165 43.480 394.395 43.950 ;
        RECT 396.185 43.665 396.690 43.895 ;
        RECT 398.145 43.685 398.550 43.915 ;
        RECT 394.165 43.250 395.955 43.480 ;
        RECT 394.070 42.610 395.490 42.990 ;
        RECT 395.725 42.355 395.955 43.250 ;
        RECT 394.265 42.125 395.955 42.355 ;
        RECT 396.185 42.375 396.415 43.665 ;
        RECT 396.810 42.610 397.840 42.990 ;
        RECT 396.185 42.145 397.815 42.375 ;
        RECT 398.145 42.340 398.375 43.685 ;
        RECT 394.265 41.535 394.495 42.125 ;
        RECT 396.185 41.545 396.535 42.145 ;
        RECT 397.585 41.770 397.815 42.145 ;
        RECT 398.045 42.000 398.375 42.340 ;
        RECT 398.605 41.770 398.835 42.850 ;
        RECT 399.385 42.690 399.615 43.970 ;
        RECT 402.920 43.610 403.150 44.000 ;
        RECT 399.965 43.380 403.150 43.610 ;
        RECT 399.965 43.170 400.195 43.380 ;
        RECT 403.910 43.150 404.250 43.760 ;
        RECT 404.845 43.170 405.075 44.000 ;
        RECT 400.610 42.920 404.590 43.150 ;
        RECT 399.065 42.460 404.075 42.690 ;
        RECT 399.065 42.000 399.295 42.460 ;
        RECT 403.775 42.235 404.075 42.460 ;
        RECT 400.085 42.000 402.915 42.230 ;
        RECT 400.085 41.805 400.315 42.000 ;
        RECT 397.585 41.540 398.835 41.770 ;
        RECT 402.685 41.630 402.915 42.000 ;
        RECT 404.360 41.915 404.590 42.920 ;
        RECT 405.470 42.940 405.810 43.760 ;
        RECT 406.040 43.400 406.270 44.000 ;
        RECT 406.870 43.630 407.675 43.970 ;
        RECT 406.040 43.170 407.040 43.400 ;
        RECT 405.470 42.710 406.360 42.940 ;
        RECT 404.360 41.685 405.000 41.915 ;
        RECT 406.130 41.600 406.360 42.710 ;
        RECT 406.810 42.235 407.040 43.170 ;
        RECT 407.335 41.830 407.675 43.630 ;
        RECT 408.580 43.740 410.215 44.100 ;
        RECT 408.580 42.930 409.125 43.740 ;
        RECT 410.570 43.310 410.800 43.970 ;
        RECT 409.650 43.080 412.150 43.310 ;
        RECT 409.650 42.585 409.880 43.080 ;
        RECT 407.915 42.355 409.880 42.585 ;
        RECT 408.115 41.710 409.385 41.940 ;
        RECT 409.650 41.830 409.880 42.355 ;
        RECT 408.115 41.600 408.345 41.710 ;
        RECT 406.130 41.370 408.345 41.600 ;
        RECT 409.155 41.600 409.385 41.710 ;
        RECT 410.110 41.600 410.340 42.850 ;
        RECT 409.155 41.370 410.340 41.600 ;
        RECT 412.395 41.380 412.830 44.210 ;
        RECT 416.540 43.890 417.880 44.210 ;
        RECT 421.020 43.890 422.360 44.210 ;
        RECT 415.305 42.990 415.645 43.600 ;
        RECT 416.440 42.990 416.780 43.600 ;
        RECT 415.305 42.610 416.210 42.990 ;
        RECT 416.440 42.610 417.345 42.990 ;
        RECT 416.550 41.600 416.890 42.265 ;
        RECT 417.575 42.035 417.880 43.890 ;
        RECT 418.110 42.990 418.460 43.600 ;
        RECT 419.785 42.990 420.125 43.600 ;
        RECT 420.920 42.990 421.260 43.600 ;
        RECT 418.110 42.610 419.005 42.990 ;
        RECT 419.785 42.610 420.690 42.990 ;
        RECT 420.920 42.610 421.825 42.990 ;
        RECT 418.590 41.600 418.930 42.265 ;
        RECT 416.550 41.370 418.930 41.600 ;
        RECT 421.030 41.600 421.370 42.265 ;
        RECT 422.055 42.035 422.360 43.890 ;
        RECT 422.590 42.990 422.940 43.600 ;
        RECT 422.590 42.610 423.485 42.990 ;
        RECT 423.070 41.600 423.410 42.265 ;
        RECT 421.030 41.370 423.410 41.600 ;
        RECT 424.850 41.380 425.285 44.210 ;
        RECT 426.880 43.310 427.110 43.970 ;
        RECT 427.465 43.740 429.100 44.100 ;
        RECT 431.410 44.000 434.760 44.230 ;
        RECT 425.530 43.080 428.030 43.310 ;
        RECT 427.340 41.600 427.570 42.850 ;
        RECT 427.800 42.585 428.030 43.080 ;
        RECT 428.555 42.930 429.100 43.740 ;
        RECT 430.005 43.630 430.810 43.970 ;
        RECT 427.800 42.355 429.765 42.585 ;
        RECT 427.800 41.830 428.030 42.355 ;
        RECT 428.295 41.710 429.565 41.940 ;
        RECT 430.005 41.830 430.345 43.630 ;
        RECT 431.410 43.400 431.640 44.000 ;
        RECT 430.640 43.170 431.640 43.400 ;
        RECT 430.640 42.235 430.870 43.170 ;
        RECT 431.870 42.940 432.210 43.760 ;
        RECT 432.605 43.170 432.835 44.000 ;
        RECT 433.430 43.150 433.770 43.760 ;
        RECT 434.530 43.610 434.760 44.000 ;
        RECT 434.530 43.380 437.715 43.610 ;
        RECT 437.485 43.170 437.715 43.380 ;
        RECT 431.320 42.710 432.210 42.940 ;
        RECT 433.090 42.920 437.070 43.150 ;
        RECT 428.295 41.600 428.525 41.710 ;
        RECT 427.340 41.370 428.525 41.600 ;
        RECT 429.335 41.600 429.565 41.710 ;
        RECT 431.320 41.600 431.550 42.710 ;
        RECT 433.090 41.915 433.320 42.920 ;
        RECT 438.065 42.690 438.295 43.970 ;
        RECT 439.130 43.685 439.535 43.915 ;
        RECT 433.605 42.460 438.615 42.690 ;
        RECT 433.605 42.235 433.905 42.460 ;
        RECT 432.680 41.685 433.320 41.915 ;
        RECT 434.765 42.000 437.595 42.230 ;
        RECT 438.385 42.000 438.615 42.460 ;
        RECT 434.765 41.630 434.995 42.000 ;
        RECT 437.365 41.805 437.595 42.000 ;
        RECT 438.845 41.770 439.075 42.850 ;
        RECT 439.305 42.340 439.535 43.685 ;
        RECT 440.990 43.665 441.495 43.895 ;
        RECT 439.840 42.610 440.870 42.990 ;
        RECT 441.265 42.375 441.495 43.665 ;
        RECT 443.285 43.480 443.515 43.950 ;
        RECT 439.305 42.000 439.635 42.340 ;
        RECT 439.865 42.145 441.495 42.375 ;
        RECT 439.865 41.770 440.095 42.145 ;
        RECT 429.335 41.370 431.550 41.600 ;
        RECT 438.845 41.540 440.095 41.770 ;
        RECT 441.145 41.545 441.495 42.145 ;
        RECT 441.725 43.250 443.515 43.480 ;
        RECT 441.725 42.355 441.955 43.250 ;
        RECT 442.190 42.610 443.610 42.990 ;
        RECT 441.725 42.125 443.415 42.355 ;
        RECT 443.185 41.535 443.415 42.125 ;
        RECT 444.465 41.440 444.770 43.580 ;
        RECT 445.000 42.400 445.355 44.160 ;
        RECT 445.585 42.970 445.890 44.160 ;
        RECT 445.585 42.630 446.615 42.970 ;
        RECT 445.000 42.080 446.425 42.400 ;
        RECT 446.145 41.380 446.425 42.080 ;
        RECT 448.380 42.050 448.715 43.950 ;
        RECT 449.605 43.205 450.880 43.435 ;
        RECT 449.605 41.370 449.835 43.205 ;
        RECT 451.125 42.800 451.355 44.230 ;
        RECT 450.090 42.570 451.355 42.800 ;
        RECT 454.085 43.205 455.360 43.435 ;
        RECT 454.085 41.370 454.315 43.205 ;
        RECT 455.605 42.800 455.835 44.230 ;
        RECT 454.570 42.570 455.835 42.800 ;
        RECT 456.325 43.205 457.600 43.435 ;
        RECT 456.325 41.370 456.555 43.205 ;
        RECT 457.845 42.800 458.075 44.230 ;
        RECT 456.810 42.570 458.075 42.800 ;
        RECT 458.565 43.205 459.840 43.435 ;
        RECT 458.565 41.370 458.795 43.205 ;
        RECT 460.085 42.800 460.315 44.230 ;
        RECT 459.050 42.570 460.315 42.800 ;
        RECT 298.905 39.630 299.135 40.300 ;
        RECT 301.145 39.630 301.375 40.300 ;
        RECT 303.385 39.630 303.615 40.300 ;
        RECT 305.525 39.630 305.755 40.300 ;
        RECT 307.865 39.680 308.095 40.300 ;
        RECT 310.105 39.680 310.335 40.300 ;
        RECT 298.870 39.250 305.755 39.630 ;
        RECT 307.285 39.450 310.335 39.680 ;
        RECT 298.060 38.605 301.260 38.950 ;
        RECT 301.960 38.340 302.760 39.250 ;
        RECT 307.285 38.945 307.620 39.450 ;
        RECT 303.330 38.605 307.620 38.945 ;
        RECT 308.090 38.635 310.950 39.070 ;
        RECT 298.805 37.960 305.755 38.340 ;
        RECT 298.805 37.595 299.035 37.960 ;
        RECT 301.045 37.595 301.275 37.960 ;
        RECT 303.285 37.595 303.515 37.960 ;
        RECT 305.495 37.595 305.755 37.960 ;
        RECT 307.285 38.170 307.620 38.605 ;
        RECT 307.285 37.935 310.235 38.170 ;
        RECT 307.765 37.595 307.995 37.935 ;
        RECT 310.005 37.595 310.235 37.935 ;
        RECT 312.860 37.730 313.195 39.630 ;
        RECT 318.665 39.555 318.895 40.145 ;
        RECT 318.665 39.325 320.355 39.555 ;
        RECT 318.470 38.690 319.890 39.070 ;
        RECT 320.125 38.430 320.355 39.325 ;
        RECT 318.565 38.200 320.355 38.430 ;
        RECT 320.585 39.535 320.935 40.135 ;
        RECT 321.985 39.910 323.235 40.140 ;
        RECT 330.530 40.080 332.745 40.310 ;
        RECT 321.985 39.535 322.215 39.910 ;
        RECT 320.585 39.305 322.215 39.535 ;
        RECT 322.445 39.340 322.775 39.680 ;
        RECT 318.565 37.730 318.795 38.200 ;
        RECT 320.585 38.015 320.815 39.305 ;
        RECT 321.210 38.690 322.240 39.070 ;
        RECT 320.585 37.785 321.090 38.015 ;
        RECT 322.545 37.995 322.775 39.340 ;
        RECT 323.005 38.830 323.235 39.910 ;
        RECT 324.485 39.680 324.715 39.875 ;
        RECT 327.085 39.680 327.315 40.050 ;
        RECT 323.465 39.220 323.695 39.680 ;
        RECT 324.485 39.450 327.315 39.680 ;
        RECT 328.760 39.765 329.400 39.995 ;
        RECT 328.175 39.220 328.475 39.445 ;
        RECT 323.465 38.990 328.475 39.220 ;
        RECT 322.545 37.765 322.950 37.995 ;
        RECT 323.785 37.710 324.015 38.990 ;
        RECT 328.760 38.760 328.990 39.765 ;
        RECT 330.530 38.970 330.760 40.080 ;
        RECT 332.515 39.970 332.745 40.080 ;
        RECT 333.555 40.080 334.740 40.310 ;
        RECT 333.555 39.970 333.785 40.080 ;
        RECT 325.010 38.530 328.990 38.760 ;
        RECT 329.870 38.740 330.760 38.970 ;
        RECT 324.365 38.300 324.595 38.510 ;
        RECT 324.365 38.070 327.550 38.300 ;
        RECT 327.320 37.680 327.550 38.070 ;
        RECT 328.310 37.920 328.650 38.530 ;
        RECT 329.245 37.680 329.475 38.510 ;
        RECT 329.870 37.920 330.210 38.740 ;
        RECT 331.210 38.510 331.440 39.445 ;
        RECT 330.440 38.280 331.440 38.510 ;
        RECT 330.440 37.680 330.670 38.280 ;
        RECT 331.735 38.050 332.075 39.850 ;
        RECT 332.515 39.740 333.785 39.970 ;
        RECT 334.050 39.325 334.280 39.850 ;
        RECT 332.315 39.095 334.280 39.325 ;
        RECT 331.270 37.710 332.075 38.050 ;
        RECT 332.980 37.940 333.525 38.750 ;
        RECT 334.050 38.600 334.280 39.095 ;
        RECT 334.510 38.830 334.740 40.080 ;
        RECT 334.050 38.370 336.550 38.600 ;
        RECT 332.980 37.890 334.615 37.940 ;
        RECT 327.320 37.450 330.670 37.680 ;
        RECT 332.970 37.630 334.615 37.890 ;
        RECT 334.970 37.710 335.200 38.370 ;
        RECT 332.980 37.580 334.615 37.630 ;
        RECT 336.795 37.470 337.230 40.300 ;
        RECT 339.270 40.080 341.650 40.310 ;
        RECT 339.270 39.415 339.610 40.080 ;
        RECT 338.025 38.690 338.930 39.070 ;
        RECT 339.160 38.690 340.065 39.070 ;
        RECT 338.025 38.080 338.365 38.690 ;
        RECT 339.160 38.080 339.500 38.690 ;
        RECT 339.750 37.790 340.010 37.950 ;
        RECT 340.295 37.790 340.600 39.645 ;
        RECT 341.310 39.415 341.650 40.080 ;
        RECT 340.830 38.690 341.725 39.070 ;
        RECT 340.830 38.080 341.180 38.690 ;
        RECT 339.260 37.470 340.600 37.790 ;
        RECT 343.605 37.730 343.940 39.630 ;
        RECT 344.325 38.475 344.555 40.310 ;
        RECT 344.810 38.880 346.075 39.110 ;
        RECT 344.325 38.245 345.600 38.475 ;
        RECT 343.670 37.570 343.930 37.730 ;
        RECT 345.845 37.450 346.075 38.880 ;
        RECT 346.565 38.475 346.795 40.310 ;
        RECT 347.050 38.880 348.315 39.110 ;
        RECT 346.565 38.245 347.840 38.475 ;
        RECT 348.085 37.450 348.315 38.880 ;
        RECT 348.805 38.475 349.035 40.310 ;
        RECT 349.290 38.880 350.555 39.110 ;
        RECT 348.805 38.245 350.080 38.475 ;
        RECT 350.325 37.450 350.555 38.880 ;
        RECT 351.045 38.475 351.275 40.310 ;
        RECT 351.530 38.880 352.795 39.110 ;
        RECT 351.045 38.245 352.320 38.475 ;
        RECT 352.565 37.450 352.795 38.880 ;
        RECT 356.085 38.475 356.315 40.310 ;
        RECT 356.570 38.880 357.835 39.110 ;
        RECT 356.085 38.245 357.360 38.475 ;
        RECT 357.605 37.450 357.835 38.880 ;
        RECT 358.325 38.475 358.555 40.310 ;
        RECT 358.810 38.880 360.075 39.110 ;
        RECT 358.325 38.245 359.600 38.475 ;
        RECT 359.845 37.450 360.075 38.880 ;
        RECT 360.965 37.520 361.300 40.290 ;
        RECT 361.530 37.890 361.855 39.870 ;
        RECT 362.815 39.680 363.155 40.300 ;
        RECT 364.380 40.065 367.235 40.300 ;
        RECT 364.380 39.680 364.610 40.065 ;
        RECT 362.815 39.450 364.610 39.680 ;
        RECT 364.910 39.300 366.450 39.630 ;
        RECT 366.895 39.450 367.235 40.065 ;
        RECT 363.170 38.690 364.130 39.070 ;
        RECT 363.170 38.005 363.565 38.690 ;
        RECT 364.360 37.470 364.680 39.070 ;
        RECT 364.910 37.505 365.240 39.300 ;
        RECT 365.480 37.470 365.800 39.070 ;
        RECT 366.040 38.720 367.105 39.070 ;
        RECT 366.040 37.470 366.360 38.720 ;
        RECT 367.845 38.475 368.075 40.310 ;
        RECT 368.330 38.880 369.595 39.110 ;
        RECT 367.845 38.245 369.120 38.475 ;
        RECT 369.365 37.450 369.595 38.880 ;
        RECT 370.085 38.475 370.315 40.310 ;
        RECT 370.570 38.880 371.835 39.110 ;
        RECT 370.085 38.245 371.360 38.475 ;
        RECT 371.605 37.450 371.835 38.880 ;
        RECT 372.325 38.475 372.555 40.310 ;
        RECT 372.810 38.880 374.075 39.110 ;
        RECT 372.325 38.245 373.600 38.475 ;
        RECT 373.845 37.450 374.075 38.880 ;
        RECT 374.565 38.475 374.795 40.310 ;
        RECT 375.050 38.880 376.315 39.110 ;
        RECT 374.565 38.245 375.840 38.475 ;
        RECT 376.085 37.450 376.315 38.880 ;
        RECT 376.805 38.475 377.035 40.310 ;
        RECT 377.290 38.880 378.555 39.110 ;
        RECT 376.805 38.245 378.080 38.475 ;
        RECT 378.325 37.450 378.555 38.880 ;
        RECT 379.045 38.475 379.275 40.310 ;
        RECT 379.530 38.880 380.795 39.110 ;
        RECT 379.045 38.245 380.320 38.475 ;
        RECT 380.565 37.450 380.795 38.880 ;
        RECT 381.285 38.475 381.515 40.310 ;
        RECT 381.770 38.880 383.035 39.110 ;
        RECT 381.285 38.245 382.560 38.475 ;
        RECT 382.805 37.450 383.035 38.880 ;
        RECT 383.525 38.475 383.755 40.310 ;
        RECT 385.870 39.210 386.500 40.265 ;
        RECT 384.010 38.880 385.275 39.110 ;
        RECT 383.525 38.245 384.800 38.475 ;
        RECT 385.045 37.450 385.275 38.880 ;
        RECT 385.870 37.960 386.200 39.210 ;
        RECT 387.860 38.660 388.220 40.265 ;
        RECT 388.460 40.050 389.665 40.280 ;
        RECT 386.465 38.430 387.320 38.560 ;
        RECT 388.460 38.430 388.690 40.050 ;
        RECT 386.465 38.200 388.690 38.430 ;
        RECT 385.870 37.530 386.635 37.960 ;
        RECT 388.295 37.450 388.690 38.200 ;
        RECT 388.920 37.995 389.340 39.800 ;
        RECT 390.705 37.890 391.030 39.870 ;
        RECT 391.260 37.520 391.595 40.290 ;
        RECT 395.285 38.475 395.515 40.310 ;
        RECT 395.770 38.880 397.035 39.110 ;
        RECT 395.285 38.245 396.560 38.475 ;
        RECT 396.805 37.450 397.035 38.880 ;
        RECT 397.525 38.475 397.755 40.310 ;
        RECT 398.010 38.880 399.275 39.110 ;
        RECT 397.525 38.245 398.800 38.475 ;
        RECT 399.045 37.450 399.275 38.880 ;
        RECT 399.765 38.475 399.995 40.310 ;
        RECT 400.250 38.880 401.515 39.110 ;
        RECT 399.765 38.245 401.040 38.475 ;
        RECT 401.285 37.450 401.515 38.880 ;
        RECT 402.005 38.475 402.235 40.310 ;
        RECT 405.265 39.680 405.495 40.300 ;
        RECT 407.505 39.680 407.735 40.300 ;
        RECT 405.265 39.450 408.315 39.680 ;
        RECT 402.490 38.880 403.755 39.110 ;
        RECT 402.005 38.245 403.280 38.475 ;
        RECT 403.525 37.450 403.755 38.880 ;
        RECT 404.650 38.635 407.510 39.070 ;
        RECT 407.980 38.945 408.315 39.450 ;
        RECT 420.425 39.630 420.655 40.300 ;
        RECT 422.665 39.630 422.895 40.300 ;
        RECT 424.905 39.630 425.135 40.300 ;
        RECT 427.045 39.630 427.275 40.300 ;
        RECT 429.385 39.680 429.615 40.300 ;
        RECT 431.625 39.680 431.855 40.300 ;
        RECT 420.425 39.250 427.370 39.630 ;
        RECT 428.805 39.450 431.855 39.680 ;
        RECT 436.150 40.080 438.530 40.310 ;
        RECT 407.980 38.605 412.270 38.945 ;
        RECT 414.340 38.605 417.540 38.950 ;
        RECT 419.580 38.605 422.780 38.950 ;
        RECT 407.980 38.170 408.315 38.605 ;
        RECT 423.480 38.340 424.280 39.250 ;
        RECT 428.805 38.945 429.140 39.450 ;
        RECT 436.150 39.415 436.490 40.080 ;
        RECT 424.850 38.605 429.140 38.945 ;
        RECT 429.610 38.635 432.470 39.070 ;
        RECT 434.905 38.690 435.810 39.070 ;
        RECT 436.040 38.690 436.945 39.070 ;
        RECT 405.365 37.935 408.315 38.170 ;
        RECT 420.325 37.960 427.275 38.340 ;
        RECT 405.365 37.595 405.595 37.935 ;
        RECT 407.605 37.595 407.835 37.935 ;
        RECT 420.325 37.595 420.555 37.960 ;
        RECT 422.565 37.595 422.795 37.960 ;
        RECT 424.805 37.595 425.035 37.960 ;
        RECT 427.015 37.595 427.275 37.960 ;
        RECT 428.805 38.170 429.140 38.605 ;
        RECT 428.805 37.935 431.755 38.170 ;
        RECT 434.905 38.080 435.245 38.690 ;
        RECT 436.040 38.080 436.380 38.690 ;
        RECT 429.285 37.595 429.515 37.935 ;
        RECT 431.525 37.595 431.755 37.935 ;
        RECT 437.175 37.790 437.480 39.645 ;
        RECT 438.190 39.415 438.530 40.080 ;
        RECT 437.710 38.690 438.605 39.070 ;
        RECT 437.710 38.080 438.060 38.690 ;
        RECT 439.425 38.100 439.730 40.240 ;
        RECT 439.990 39.600 440.250 39.630 ;
        RECT 441.105 39.600 441.385 40.300 ;
        RECT 439.960 39.280 441.385 39.600 ;
        RECT 436.140 37.470 437.480 37.790 ;
        RECT 439.960 37.520 440.315 39.280 ;
        RECT 440.545 38.710 441.575 39.050 ;
        RECT 440.545 37.520 440.850 38.710 ;
        RECT 442.210 37.470 442.645 40.300 ;
        RECT 444.700 40.080 445.885 40.310 ;
        RECT 444.700 38.830 444.930 40.080 ;
        RECT 445.655 39.970 445.885 40.080 ;
        RECT 446.695 40.080 448.910 40.310 ;
        RECT 446.695 39.970 446.925 40.080 ;
        RECT 445.160 39.325 445.390 39.850 ;
        RECT 445.655 39.740 446.925 39.970 ;
        RECT 445.160 39.095 447.125 39.325 ;
        RECT 445.160 38.600 445.390 39.095 ;
        RECT 442.890 38.370 445.390 38.600 ;
        RECT 444.240 37.710 444.470 38.370 ;
        RECT 445.915 37.940 446.460 38.750 ;
        RECT 444.825 37.890 446.460 37.940 ;
        RECT 447.365 38.050 447.705 39.850 ;
        RECT 448.000 38.510 448.230 39.445 ;
        RECT 448.680 38.970 448.910 40.080 ;
        RECT 450.040 39.765 450.680 39.995 ;
        RECT 448.680 38.740 449.570 38.970 ;
        RECT 448.000 38.280 449.000 38.510 ;
        RECT 444.825 37.630 446.470 37.890 ;
        RECT 447.365 37.710 448.170 38.050 ;
        RECT 448.770 37.680 449.000 38.280 ;
        RECT 449.230 37.920 449.570 38.740 ;
        RECT 450.450 38.760 450.680 39.765 ;
        RECT 452.125 39.680 452.355 40.050 ;
        RECT 456.205 39.910 457.455 40.140 ;
        RECT 454.725 39.680 454.955 39.875 ;
        RECT 452.125 39.450 454.955 39.680 ;
        RECT 450.965 39.220 451.265 39.445 ;
        RECT 455.745 39.220 455.975 39.680 ;
        RECT 450.965 38.990 455.975 39.220 ;
        RECT 450.450 38.530 454.430 38.760 ;
        RECT 449.965 37.680 450.195 38.510 ;
        RECT 450.790 37.920 451.130 38.530 ;
        RECT 454.845 38.300 455.075 38.510 ;
        RECT 451.890 38.070 455.075 38.300 ;
        RECT 451.890 37.680 452.120 38.070 ;
        RECT 455.425 37.710 455.655 38.990 ;
        RECT 456.205 38.830 456.435 39.910 ;
        RECT 456.665 39.340 456.995 39.680 ;
        RECT 457.225 39.535 457.455 39.910 ;
        RECT 458.505 39.535 458.855 40.135 ;
        RECT 460.545 39.555 460.775 40.145 ;
        RECT 456.665 37.995 456.895 39.340 ;
        RECT 457.225 39.305 458.855 39.535 ;
        RECT 457.200 38.690 458.230 39.070 ;
        RECT 458.625 38.015 458.855 39.305 ;
        RECT 459.085 39.325 460.775 39.555 ;
        RECT 459.085 38.430 459.315 39.325 ;
        RECT 459.550 38.690 460.840 39.070 ;
        RECT 459.085 38.200 460.875 38.430 ;
        RECT 456.490 37.765 456.895 37.995 ;
        RECT 458.350 37.785 458.855 38.015 ;
        RECT 460.645 37.730 460.875 38.200 ;
        RECT 444.825 37.580 446.460 37.630 ;
        RECT 448.770 37.450 452.120 37.680 ;
        RECT 298.805 35.880 299.035 36.245 ;
        RECT 301.045 35.880 301.275 36.245 ;
        RECT 303.285 35.880 303.515 36.245 ;
        RECT 305.495 35.880 305.755 36.245 ;
        RECT 307.765 35.905 307.995 36.245 ;
        RECT 310.005 35.905 310.235 36.245 ;
        RECT 298.805 35.500 305.755 35.880 ;
        RECT 307.285 35.670 310.235 35.905 ;
        RECT 168.115 34.250 168.495 35.150 ;
        RECT 174.115 34.250 174.495 35.150 ;
        RECT 178.045 34.355 178.425 35.215 ;
        RECT 180.185 34.355 180.565 35.215 ;
        RECT 166.935 34.020 169.675 34.250 ;
        RECT 173.735 34.020 174.875 34.250 ;
        RECT 178.045 34.020 179.075 34.355 ;
        RECT 179.535 34.020 180.565 34.355 ;
        RECT 186.615 34.250 186.995 35.150 ;
        RECT 298.060 34.890 301.260 35.235 ;
        RECT 301.960 34.590 302.760 35.500 ;
        RECT 307.285 35.235 307.620 35.670 ;
        RECT 303.330 34.895 307.620 35.235 ;
        RECT 311.845 35.365 313.120 35.595 ;
        RECT 183.835 34.020 189.775 34.250 ;
        RECT 298.905 34.210 305.755 34.590 ;
        RECT 166.590 30.810 166.820 33.790 ;
        RECT 168.190 30.810 168.420 33.790 ;
        RECT 169.790 30.810 170.020 33.790 ;
        RECT 166.590 30.510 170.020 30.810 ;
        RECT 173.390 30.810 173.620 33.790 ;
        RECT 174.990 30.810 175.220 33.790 ;
        RECT 173.390 30.510 175.220 30.810 ;
        RECT 166.590 25.250 166.890 30.510 ;
        RECT 173.390 27.250 173.690 30.510 ;
        RECT 178.355 29.640 178.655 33.790 ;
        RECT 179.955 29.640 180.255 33.790 ;
        RECT 184.290 30.810 184.520 33.790 ;
        RECT 185.890 30.810 186.120 33.790 ;
        RECT 187.490 30.810 187.720 33.790 ;
        RECT 189.090 30.810 189.320 33.790 ;
        RECT 298.905 33.540 299.135 34.210 ;
        RECT 301.145 33.540 301.375 34.210 ;
        RECT 303.385 33.540 303.615 34.210 ;
        RECT 305.525 33.540 305.755 34.210 ;
        RECT 307.285 34.390 307.620 34.895 ;
        RECT 308.090 34.770 310.950 35.205 ;
        RECT 307.285 34.160 310.335 34.390 ;
        RECT 307.865 33.540 308.095 34.160 ;
        RECT 310.105 33.540 310.335 34.160 ;
        RECT 311.845 33.530 312.075 35.365 ;
        RECT 313.365 34.960 313.595 36.390 ;
        RECT 312.330 34.730 313.595 34.960 ;
        RECT 314.085 35.365 315.360 35.595 ;
        RECT 314.085 33.530 314.315 35.365 ;
        RECT 315.605 34.960 315.835 36.390 ;
        RECT 314.570 34.730 315.835 34.960 ;
        RECT 316.325 35.365 317.600 35.595 ;
        RECT 316.325 33.530 316.555 35.365 ;
        RECT 317.845 34.960 318.075 36.390 ;
        RECT 316.810 34.730 318.075 34.960 ;
        RECT 318.565 35.365 319.840 35.595 ;
        RECT 318.565 33.530 318.795 35.365 ;
        RECT 320.085 34.960 320.315 36.390 ;
        RECT 319.050 34.730 320.315 34.960 ;
        RECT 320.805 35.365 322.080 35.595 ;
        RECT 320.805 33.530 321.035 35.365 ;
        RECT 322.325 34.960 322.555 36.390 ;
        RECT 321.290 34.730 322.555 34.960 ;
        RECT 323.045 35.365 324.320 35.595 ;
        RECT 323.045 33.530 323.275 35.365 ;
        RECT 324.565 34.960 324.795 36.390 ;
        RECT 323.530 34.730 324.795 34.960 ;
        RECT 325.285 35.365 326.560 35.595 ;
        RECT 325.285 33.530 325.515 35.365 ;
        RECT 326.805 34.960 327.035 36.390 ;
        RECT 325.770 34.730 327.035 34.960 ;
        RECT 327.525 35.365 328.800 35.595 ;
        RECT 327.525 33.530 327.755 35.365 ;
        RECT 329.045 34.960 329.275 36.390 ;
        RECT 328.010 34.730 329.275 34.960 ;
        RECT 329.765 35.365 331.040 35.595 ;
        RECT 329.765 33.530 329.995 35.365 ;
        RECT 331.285 34.960 331.515 36.390 ;
        RECT 330.250 34.730 331.515 34.960 ;
        RECT 332.005 35.365 333.280 35.595 ;
        RECT 332.005 33.530 332.235 35.365 ;
        RECT 333.525 34.960 333.755 36.390 ;
        RECT 337.470 35.130 337.775 36.320 ;
        RECT 332.490 34.730 333.755 34.960 ;
        RECT 336.745 34.790 337.775 35.130 ;
        RECT 338.005 34.560 338.360 36.320 ;
        RECT 350.840 36.160 354.190 36.390 ;
        RECT 336.935 34.240 338.360 34.560 ;
        RECT 336.935 33.540 337.215 34.240 ;
        RECT 338.590 33.600 338.895 35.740 ;
        RECT 340.860 34.210 341.195 36.110 ;
        RECT 342.085 35.640 342.315 36.110 ;
        RECT 344.105 35.825 344.610 36.055 ;
        RECT 346.065 35.845 346.470 36.075 ;
        RECT 342.085 35.410 343.875 35.640 ;
        RECT 341.990 34.770 343.410 35.150 ;
        RECT 343.645 34.515 343.875 35.410 ;
        RECT 342.185 34.285 343.875 34.515 ;
        RECT 344.105 34.535 344.335 35.825 ;
        RECT 344.730 34.770 345.760 35.150 ;
        RECT 344.105 34.305 345.735 34.535 ;
        RECT 346.065 34.500 346.295 35.845 ;
        RECT 342.185 33.695 342.415 34.285 ;
        RECT 344.105 33.705 344.455 34.305 ;
        RECT 345.505 33.930 345.735 34.305 ;
        RECT 345.965 34.160 346.295 34.500 ;
        RECT 346.525 33.930 346.755 35.010 ;
        RECT 347.305 34.850 347.535 36.130 ;
        RECT 350.840 35.770 351.070 36.160 ;
        RECT 347.885 35.540 351.070 35.770 ;
        RECT 347.885 35.330 348.115 35.540 ;
        RECT 351.830 35.310 352.170 35.920 ;
        RECT 352.765 35.330 352.995 36.160 ;
        RECT 348.530 35.080 352.510 35.310 ;
        RECT 346.985 34.620 351.995 34.850 ;
        RECT 346.985 34.160 347.215 34.620 ;
        RECT 351.695 34.395 351.995 34.620 ;
        RECT 348.005 34.160 350.835 34.390 ;
        RECT 348.005 33.965 348.235 34.160 ;
        RECT 345.505 33.700 346.755 33.930 ;
        RECT 350.605 33.790 350.835 34.160 ;
        RECT 352.280 34.075 352.510 35.080 ;
        RECT 353.390 35.100 353.730 35.920 ;
        RECT 353.960 35.560 354.190 36.160 ;
        RECT 354.790 35.790 355.595 36.130 ;
        RECT 353.960 35.330 354.960 35.560 ;
        RECT 353.390 34.870 354.280 35.100 ;
        RECT 352.280 33.845 352.920 34.075 ;
        RECT 354.050 33.760 354.280 34.870 ;
        RECT 354.730 34.395 354.960 35.330 ;
        RECT 355.255 33.990 355.595 35.790 ;
        RECT 356.500 35.900 358.135 36.260 ;
        RECT 356.500 35.090 357.045 35.900 ;
        RECT 358.490 35.470 358.720 36.130 ;
        RECT 357.570 35.240 360.070 35.470 ;
        RECT 357.570 34.745 357.800 35.240 ;
        RECT 355.835 34.515 357.800 34.745 ;
        RECT 356.035 33.870 357.305 34.100 ;
        RECT 357.570 33.990 357.800 34.515 ;
        RECT 356.035 33.760 356.265 33.870 ;
        RECT 354.050 33.530 356.265 33.760 ;
        RECT 357.075 33.760 357.305 33.870 ;
        RECT 358.030 33.760 358.260 35.010 ;
        RECT 357.075 33.530 358.260 33.760 ;
        RECT 360.315 33.540 360.750 36.370 ;
        RECT 361.490 35.150 361.885 35.835 ;
        RECT 361.490 34.770 362.450 35.150 ;
        RECT 362.680 34.770 363.000 36.370 ;
        RECT 363.230 34.540 363.560 36.335 ;
        RECT 363.800 34.770 364.120 36.370 ;
        RECT 364.360 35.120 364.680 36.370 ;
        RECT 366.165 35.365 367.440 35.595 ;
        RECT 364.360 34.770 365.425 35.120 ;
        RECT 361.135 34.160 362.930 34.390 ;
        RECT 363.230 34.210 364.770 34.540 ;
        RECT 361.135 33.540 361.475 34.160 ;
        RECT 362.700 33.775 362.930 34.160 ;
        RECT 365.215 33.775 365.555 34.390 ;
        RECT 362.700 33.540 365.555 33.775 ;
        RECT 366.165 33.530 366.395 35.365 ;
        RECT 367.685 34.960 367.915 36.390 ;
        RECT 366.650 34.730 367.915 34.960 ;
        RECT 368.405 35.365 369.680 35.595 ;
        RECT 368.405 33.530 368.635 35.365 ;
        RECT 369.925 34.960 370.155 36.390 ;
        RECT 368.890 34.730 370.155 34.960 ;
        RECT 370.645 35.365 371.920 35.595 ;
        RECT 370.645 33.530 370.875 35.365 ;
        RECT 372.165 34.960 372.395 36.390 ;
        RECT 371.130 34.730 372.395 34.960 ;
        RECT 375.685 35.365 376.960 35.595 ;
        RECT 375.685 33.530 375.915 35.365 ;
        RECT 377.205 34.960 377.435 36.390 ;
        RECT 376.170 34.730 377.435 34.960 ;
        RECT 377.925 35.365 379.200 35.595 ;
        RECT 377.925 33.530 378.155 35.365 ;
        RECT 379.445 34.960 379.675 36.390 ;
        RECT 378.410 34.730 379.675 34.960 ;
        RECT 380.165 35.365 381.440 35.595 ;
        RECT 380.165 33.530 380.395 35.365 ;
        RECT 381.685 34.960 381.915 36.390 ;
        RECT 385.080 35.120 385.400 36.370 ;
        RECT 380.650 34.730 381.915 34.960 ;
        RECT 384.335 34.770 385.400 35.120 ;
        RECT 385.640 34.770 385.960 36.370 ;
        RECT 386.200 34.540 386.530 36.335 ;
        RECT 386.760 34.770 387.080 36.370 ;
        RECT 399.000 36.160 402.350 36.390 ;
        RECT 404.660 36.210 406.295 36.260 ;
        RECT 387.875 35.150 388.270 35.835 ;
        RECT 390.245 35.640 390.475 36.110 ;
        RECT 392.265 35.825 392.770 36.055 ;
        RECT 394.225 35.845 394.630 36.075 ;
        RECT 390.245 35.410 392.035 35.640 ;
        RECT 387.310 34.770 388.270 35.150 ;
        RECT 390.280 34.770 391.570 35.150 ;
        RECT 384.205 33.775 384.545 34.390 ;
        RECT 384.990 34.210 386.530 34.540 ;
        RECT 391.805 34.515 392.035 35.410 ;
        RECT 386.830 34.160 388.625 34.390 ;
        RECT 386.830 33.775 387.060 34.160 ;
        RECT 384.205 33.540 387.060 33.775 ;
        RECT 388.285 33.540 388.625 34.160 ;
        RECT 390.345 34.285 392.035 34.515 ;
        RECT 392.265 34.535 392.495 35.825 ;
        RECT 392.890 34.770 393.920 35.150 ;
        RECT 392.265 34.305 393.895 34.535 ;
        RECT 394.225 34.500 394.455 35.845 ;
        RECT 390.345 33.695 390.575 34.285 ;
        RECT 392.265 33.705 392.615 34.305 ;
        RECT 393.665 33.930 393.895 34.305 ;
        RECT 394.125 34.160 394.455 34.500 ;
        RECT 394.685 33.930 394.915 35.010 ;
        RECT 395.465 34.850 395.695 36.130 ;
        RECT 399.000 35.770 399.230 36.160 ;
        RECT 396.045 35.540 399.230 35.770 ;
        RECT 396.045 35.330 396.275 35.540 ;
        RECT 399.990 35.310 400.330 35.920 ;
        RECT 400.925 35.330 401.155 36.160 ;
        RECT 396.690 35.080 400.670 35.310 ;
        RECT 395.145 34.620 400.155 34.850 ;
        RECT 395.145 34.160 395.375 34.620 ;
        RECT 399.855 34.395 400.155 34.620 ;
        RECT 396.165 34.160 398.995 34.390 ;
        RECT 396.165 33.965 396.395 34.160 ;
        RECT 393.665 33.700 394.915 33.930 ;
        RECT 398.765 33.790 398.995 34.160 ;
        RECT 400.440 34.075 400.670 35.080 ;
        RECT 401.550 35.100 401.890 35.920 ;
        RECT 402.120 35.560 402.350 36.160 ;
        RECT 402.950 35.790 403.755 36.130 ;
        RECT 404.650 35.950 406.295 36.210 ;
        RECT 402.120 35.330 403.120 35.560 ;
        RECT 401.550 34.870 402.440 35.100 ;
        RECT 400.440 33.845 401.080 34.075 ;
        RECT 402.210 33.760 402.440 34.870 ;
        RECT 402.890 34.395 403.120 35.330 ;
        RECT 403.415 33.990 403.755 35.790 ;
        RECT 404.660 35.900 406.295 35.950 ;
        RECT 404.660 35.090 405.205 35.900 ;
        RECT 406.650 35.470 406.880 36.130 ;
        RECT 405.730 35.240 408.230 35.470 ;
        RECT 405.730 34.745 405.960 35.240 ;
        RECT 403.995 34.515 405.960 34.745 ;
        RECT 404.195 33.870 405.465 34.100 ;
        RECT 405.730 33.990 405.960 34.515 ;
        RECT 404.195 33.760 404.425 33.870 ;
        RECT 402.210 33.530 404.425 33.760 ;
        RECT 405.235 33.760 405.465 33.870 ;
        RECT 406.190 33.760 406.420 35.010 ;
        RECT 405.235 33.530 406.420 33.760 ;
        RECT 408.475 33.540 408.910 36.370 ;
        RECT 410.300 34.210 410.635 36.110 ;
        RECT 411.525 35.365 412.800 35.595 ;
        RECT 411.525 33.530 411.755 35.365 ;
        RECT 413.045 34.960 413.275 36.390 ;
        RECT 412.010 34.730 413.275 34.960 ;
        RECT 414.990 35.880 415.755 36.310 ;
        RECT 414.990 34.630 415.320 35.880 ;
        RECT 417.415 35.640 417.810 36.390 ;
        RECT 420.485 35.905 420.715 36.245 ;
        RECT 422.725 35.905 422.955 36.245 ;
        RECT 415.585 35.410 417.810 35.640 ;
        RECT 415.585 35.280 416.440 35.410 ;
        RECT 414.990 33.575 415.620 34.630 ;
        RECT 416.980 33.575 417.340 35.180 ;
        RECT 417.580 33.790 417.810 35.410 ;
        RECT 418.040 34.040 418.460 35.845 ;
        RECT 420.485 35.670 423.435 35.905 ;
        RECT 423.100 35.235 423.435 35.670 ;
        RECT 419.770 34.770 422.630 35.205 ;
        RECT 423.100 34.895 427.390 35.235 ;
        RECT 423.100 34.390 423.435 34.895 ;
        RECT 429.460 34.890 432.660 35.235 ;
        RECT 420.385 34.160 423.435 34.390 ;
        RECT 417.580 33.560 418.785 33.790 ;
        RECT 420.385 33.540 420.615 34.160 ;
        RECT 422.625 33.540 422.855 34.160 ;
        RECT 433.810 33.540 434.245 36.370 ;
        RECT 435.840 35.470 436.070 36.130 ;
        RECT 436.425 35.900 438.060 36.260 ;
        RECT 440.370 36.160 443.720 36.390 ;
        RECT 434.490 35.240 436.990 35.470 ;
        RECT 436.300 33.760 436.530 35.010 ;
        RECT 436.760 34.745 436.990 35.240 ;
        RECT 437.515 35.090 438.060 35.900 ;
        RECT 438.965 35.790 439.770 36.130 ;
        RECT 436.760 34.515 438.725 34.745 ;
        RECT 436.760 33.990 436.990 34.515 ;
        RECT 437.255 33.870 438.525 34.100 ;
        RECT 438.965 33.990 439.305 35.790 ;
        RECT 440.370 35.560 440.600 36.160 ;
        RECT 439.600 35.330 440.600 35.560 ;
        RECT 439.600 34.395 439.830 35.330 ;
        RECT 440.830 35.100 441.170 35.920 ;
        RECT 441.565 35.330 441.795 36.160 ;
        RECT 442.390 35.310 442.730 35.920 ;
        RECT 443.490 35.770 443.720 36.160 ;
        RECT 443.490 35.540 446.675 35.770 ;
        RECT 446.445 35.330 446.675 35.540 ;
        RECT 440.280 34.870 441.170 35.100 ;
        RECT 442.050 35.080 446.030 35.310 ;
        RECT 437.255 33.760 437.485 33.870 ;
        RECT 436.300 33.530 437.485 33.760 ;
        RECT 438.295 33.760 438.525 33.870 ;
        RECT 440.280 33.760 440.510 34.870 ;
        RECT 442.050 34.075 442.280 35.080 ;
        RECT 447.025 34.850 447.255 36.130 ;
        RECT 448.090 35.845 448.495 36.075 ;
        RECT 442.565 34.620 447.575 34.850 ;
        RECT 442.565 34.395 442.865 34.620 ;
        RECT 441.640 33.845 442.280 34.075 ;
        RECT 443.725 34.160 446.555 34.390 ;
        RECT 447.345 34.160 447.575 34.620 ;
        RECT 443.725 33.790 443.955 34.160 ;
        RECT 446.325 33.965 446.555 34.160 ;
        RECT 447.805 33.930 448.035 35.010 ;
        RECT 448.265 34.500 448.495 35.845 ;
        RECT 449.950 35.825 450.455 36.055 ;
        RECT 448.800 34.770 449.830 35.150 ;
        RECT 450.225 34.535 450.455 35.825 ;
        RECT 452.245 35.640 452.475 36.110 ;
        RECT 448.265 34.160 448.595 34.500 ;
        RECT 448.825 34.305 450.455 34.535 ;
        RECT 448.825 33.930 449.055 34.305 ;
        RECT 438.295 33.530 440.510 33.760 ;
        RECT 447.805 33.700 449.055 33.930 ;
        RECT 450.105 33.705 450.455 34.305 ;
        RECT 450.685 35.410 452.475 35.640 ;
        RECT 450.685 34.515 450.915 35.410 ;
        RECT 451.150 34.770 452.570 35.150 ;
        RECT 450.685 34.285 452.375 34.515 ;
        RECT 452.145 33.695 452.375 34.285 ;
        RECT 455.605 34.210 455.940 36.110 ;
        RECT 456.325 35.365 457.600 35.595 ;
        RECT 456.325 33.530 456.555 35.365 ;
        RECT 457.845 34.960 458.075 36.390 ;
        RECT 456.810 34.730 458.075 34.960 ;
        RECT 458.565 35.365 459.840 35.595 ;
        RECT 458.565 33.530 458.795 35.365 ;
        RECT 460.085 34.960 460.315 36.390 ;
        RECT 459.050 34.730 460.315 34.960 ;
        RECT 184.290 30.510 189.320 30.810 ;
        RECT 178.355 28.740 178.970 29.640 ;
        RECT 179.710 28.740 180.255 29.640 ;
        RECT 173.390 26.950 184.570 27.250 ;
        RECT 174.110 26.350 174.490 26.950 ;
        RECT 184.190 26.350 184.570 26.950 ;
        RECT 166.590 24.950 186.810 25.250 ;
        RECT 171.870 24.350 172.250 24.950 ;
        RECT 176.350 24.350 176.730 24.950 ;
        RECT 181.950 24.350 182.330 24.950 ;
        RECT 186.430 24.350 186.810 24.950 ;
        RECT 189.020 23.250 189.320 30.510 ;
        RECT 297.285 30.635 297.515 32.470 ;
        RECT 297.770 31.040 299.035 31.270 ;
        RECT 297.285 30.405 298.560 30.635 ;
        RECT 298.805 29.610 299.035 31.040 ;
        RECT 299.525 30.635 299.755 32.470 ;
        RECT 300.010 31.040 301.275 31.270 ;
        RECT 299.525 30.405 300.800 30.635 ;
        RECT 301.045 29.610 301.275 31.040 ;
        RECT 302.725 29.680 303.060 32.450 ;
        RECT 303.290 30.050 303.615 32.030 ;
        RECT 304.565 30.635 304.795 32.470 ;
        RECT 305.050 31.040 306.315 31.270 ;
        RECT 304.565 30.405 305.840 30.635 ;
        RECT 306.085 29.610 306.315 31.040 ;
        RECT 306.805 30.635 307.035 32.470 ;
        RECT 307.290 31.040 308.555 31.270 ;
        RECT 306.805 30.405 308.080 30.635 ;
        RECT 308.325 29.610 308.555 31.040 ;
        RECT 309.045 30.635 309.275 32.470 ;
        RECT 309.530 31.040 310.795 31.270 ;
        RECT 309.045 30.405 310.320 30.635 ;
        RECT 310.565 29.610 310.795 31.040 ;
        RECT 311.285 30.635 311.515 32.470 ;
        RECT 311.770 31.040 313.035 31.270 ;
        RECT 311.285 30.405 312.560 30.635 ;
        RECT 312.805 29.610 313.035 31.040 ;
        RECT 313.525 30.635 313.755 32.470 ;
        RECT 316.985 31.715 317.215 32.305 ;
        RECT 316.985 31.485 318.675 31.715 ;
        RECT 314.010 31.040 315.275 31.270 ;
        RECT 313.525 30.405 314.800 30.635 ;
        RECT 315.045 29.610 315.275 31.040 ;
        RECT 316.920 30.850 318.210 31.230 ;
        RECT 318.445 30.590 318.675 31.485 ;
        RECT 316.885 30.360 318.675 30.590 ;
        RECT 318.905 31.695 319.255 32.295 ;
        RECT 320.305 32.070 321.555 32.300 ;
        RECT 328.850 32.240 331.065 32.470 ;
        RECT 320.305 31.695 320.535 32.070 ;
        RECT 318.905 31.465 320.535 31.695 ;
        RECT 320.765 31.500 321.095 31.840 ;
        RECT 316.885 29.890 317.115 30.360 ;
        RECT 318.905 30.175 319.135 31.465 ;
        RECT 319.530 30.850 320.560 31.230 ;
        RECT 318.905 29.945 319.410 30.175 ;
        RECT 320.865 30.155 321.095 31.500 ;
        RECT 321.325 30.990 321.555 32.070 ;
        RECT 322.805 31.840 323.035 32.035 ;
        RECT 325.405 31.840 325.635 32.210 ;
        RECT 321.785 31.380 322.015 31.840 ;
        RECT 322.805 31.610 325.635 31.840 ;
        RECT 327.080 31.925 327.720 32.155 ;
        RECT 326.495 31.380 326.795 31.605 ;
        RECT 321.785 31.150 326.795 31.380 ;
        RECT 320.865 29.925 321.270 30.155 ;
        RECT 322.105 29.870 322.335 31.150 ;
        RECT 327.080 30.920 327.310 31.925 ;
        RECT 328.850 31.130 329.080 32.240 ;
        RECT 330.835 32.130 331.065 32.240 ;
        RECT 331.875 32.240 333.060 32.470 ;
        RECT 331.875 32.130 332.105 32.240 ;
        RECT 323.330 30.690 327.310 30.920 ;
        RECT 328.190 30.900 329.080 31.130 ;
        RECT 322.685 30.460 322.915 30.670 ;
        RECT 322.685 30.230 325.870 30.460 ;
        RECT 325.640 29.840 325.870 30.230 ;
        RECT 326.630 30.080 326.970 30.690 ;
        RECT 327.565 29.840 327.795 30.670 ;
        RECT 328.190 30.080 328.530 30.900 ;
        RECT 329.530 30.670 329.760 31.605 ;
        RECT 328.760 30.440 329.760 30.670 ;
        RECT 328.760 29.840 328.990 30.440 ;
        RECT 330.055 30.210 330.395 32.010 ;
        RECT 330.835 31.900 332.105 32.130 ;
        RECT 332.370 31.485 332.600 32.010 ;
        RECT 330.635 31.255 332.600 31.485 ;
        RECT 329.590 29.870 330.395 30.210 ;
        RECT 331.300 30.100 331.845 30.910 ;
        RECT 332.370 30.760 332.600 31.255 ;
        RECT 332.830 30.990 333.060 32.240 ;
        RECT 332.370 30.530 334.870 30.760 ;
        RECT 325.640 29.610 328.990 29.840 ;
        RECT 331.300 29.740 332.935 30.100 ;
        RECT 333.290 29.870 333.520 30.530 ;
        RECT 335.115 29.630 335.550 32.460 ;
        RECT 337.590 32.240 339.970 32.470 ;
        RECT 337.590 31.575 337.930 32.240 ;
        RECT 336.345 30.850 337.250 31.230 ;
        RECT 337.480 30.850 338.385 31.230 ;
        RECT 336.345 30.240 336.685 30.850 ;
        RECT 337.480 30.240 337.820 30.850 ;
        RECT 338.615 29.950 338.920 31.805 ;
        RECT 339.630 31.575 339.970 32.240 ;
        RECT 339.150 30.850 340.045 31.230 ;
        RECT 339.150 30.240 339.500 30.850 ;
        RECT 337.580 29.630 338.920 29.950 ;
        RECT 341.420 29.890 341.755 31.790 ;
        RECT 343.660 29.890 343.995 31.790 ;
        RECT 344.885 30.635 345.115 32.470 ;
        RECT 345.370 31.040 346.635 31.270 ;
        RECT 344.885 30.405 346.160 30.635 ;
        RECT 343.670 29.730 343.930 29.890 ;
        RECT 346.405 29.610 346.635 31.040 ;
        RECT 349.205 29.680 349.540 32.450 ;
        RECT 349.770 30.050 350.095 32.030 ;
        RECT 351.045 30.635 351.275 32.470 ;
        RECT 351.530 31.040 352.795 31.270 ;
        RECT 351.045 30.405 352.320 30.635 ;
        RECT 352.565 29.610 352.795 31.040 ;
        RECT 356.085 30.635 356.315 32.470 ;
        RECT 356.570 31.040 357.835 31.270 ;
        RECT 356.085 30.405 357.360 30.635 ;
        RECT 357.605 29.610 357.835 31.040 ;
        RECT 360.190 30.685 360.555 32.400 ;
        RECT 362.545 31.835 362.875 32.460 ;
        RECT 360.850 31.600 362.875 31.835 ;
        RECT 360.850 30.960 361.190 31.600 ;
        RECT 361.530 30.820 362.415 31.230 ;
        RECT 360.190 29.645 360.780 30.685 ;
        RECT 362.040 30.115 362.415 30.820 ;
        RECT 362.645 29.645 362.875 31.600 ;
        RECT 363.465 31.715 363.695 32.305 ;
        RECT 363.465 31.485 365.155 31.715 ;
        RECT 363.270 30.850 364.690 31.230 ;
        RECT 364.925 30.590 365.155 31.485 ;
        RECT 363.365 30.360 365.155 30.590 ;
        RECT 365.385 31.695 365.735 32.295 ;
        RECT 366.785 32.070 368.035 32.300 ;
        RECT 375.330 32.240 377.545 32.470 ;
        RECT 366.785 31.695 367.015 32.070 ;
        RECT 365.385 31.465 367.015 31.695 ;
        RECT 367.245 31.500 367.575 31.840 ;
        RECT 363.365 29.890 363.595 30.360 ;
        RECT 365.385 30.175 365.615 31.465 ;
        RECT 366.010 30.850 367.040 31.230 ;
        RECT 365.385 29.945 365.890 30.175 ;
        RECT 367.345 30.155 367.575 31.500 ;
        RECT 367.805 30.990 368.035 32.070 ;
        RECT 369.285 31.840 369.515 32.035 ;
        RECT 371.885 31.840 372.115 32.210 ;
        RECT 368.265 31.380 368.495 31.840 ;
        RECT 369.285 31.610 372.115 31.840 ;
        RECT 373.560 31.925 374.200 32.155 ;
        RECT 372.975 31.380 373.275 31.605 ;
        RECT 368.265 31.150 373.275 31.380 ;
        RECT 367.345 29.925 367.750 30.155 ;
        RECT 368.585 29.870 368.815 31.150 ;
        RECT 373.560 30.920 373.790 31.925 ;
        RECT 375.330 31.130 375.560 32.240 ;
        RECT 377.315 32.130 377.545 32.240 ;
        RECT 378.355 32.240 379.540 32.470 ;
        RECT 378.355 32.130 378.585 32.240 ;
        RECT 369.810 30.690 373.790 30.920 ;
        RECT 374.670 30.900 375.560 31.130 ;
        RECT 369.165 30.460 369.395 30.670 ;
        RECT 369.165 30.230 372.350 30.460 ;
        RECT 372.120 29.840 372.350 30.230 ;
        RECT 373.110 30.080 373.450 30.690 ;
        RECT 374.045 29.840 374.275 30.670 ;
        RECT 374.670 30.080 375.010 30.900 ;
        RECT 376.010 30.670 376.240 31.605 ;
        RECT 375.240 30.440 376.240 30.670 ;
        RECT 375.240 29.840 375.470 30.440 ;
        RECT 376.535 30.210 376.875 32.010 ;
        RECT 377.315 31.900 378.585 32.130 ;
        RECT 378.850 31.485 379.080 32.010 ;
        RECT 377.115 31.255 379.080 31.485 ;
        RECT 376.070 29.870 376.875 30.210 ;
        RECT 377.780 30.100 378.325 30.910 ;
        RECT 378.850 30.760 379.080 31.255 ;
        RECT 379.310 30.990 379.540 32.240 ;
        RECT 378.850 30.530 381.350 30.760 ;
        RECT 372.120 29.610 375.470 29.840 ;
        RECT 377.780 29.740 379.415 30.100 ;
        RECT 379.770 29.870 380.000 30.530 ;
        RECT 381.595 29.630 382.030 32.460 ;
        RECT 382.525 32.225 385.380 32.460 ;
        RECT 382.525 31.610 382.865 32.225 ;
        RECT 385.150 31.840 385.380 32.225 ;
        RECT 386.605 31.840 386.945 32.460 ;
        RECT 383.310 31.460 384.850 31.790 ;
        RECT 385.150 31.610 386.945 31.840 ;
        RECT 382.655 30.880 383.720 31.230 ;
        RECT 383.400 29.630 383.720 30.880 ;
        RECT 383.960 29.630 384.280 31.230 ;
        RECT 384.520 29.665 384.850 31.460 ;
        RECT 385.080 29.630 385.400 31.230 ;
        RECT 385.630 30.850 386.590 31.230 ;
        RECT 386.195 30.165 386.590 30.850 ;
        RECT 387.605 30.680 388.075 32.460 ;
        RECT 389.930 31.895 390.315 32.470 ;
        RECT 388.305 31.660 390.315 31.895 ;
        RECT 388.305 30.910 388.590 31.660 ;
        RECT 388.970 30.710 389.855 31.270 ;
        RECT 387.605 29.655 388.230 30.680 ;
        RECT 389.340 29.730 389.855 30.710 ;
        RECT 390.085 29.880 390.315 31.660 ;
        RECT 390.805 30.635 391.035 32.470 ;
        RECT 391.290 31.040 392.555 31.270 ;
        RECT 390.805 30.405 392.080 30.635 ;
        RECT 392.325 29.610 392.555 31.040 ;
        RECT 395.285 30.635 395.515 32.470 ;
        RECT 395.770 31.040 397.035 31.270 ;
        RECT 395.285 30.405 396.560 30.635 ;
        RECT 396.805 29.610 397.035 31.040 ;
        RECT 397.525 30.635 397.755 32.470 ;
        RECT 398.010 31.040 399.275 31.270 ;
        RECT 397.525 30.405 398.800 30.635 ;
        RECT 399.045 29.610 399.275 31.040 ;
        RECT 399.765 30.635 399.995 32.470 ;
        RECT 400.250 31.040 401.515 31.270 ;
        RECT 399.765 30.405 401.040 30.635 ;
        RECT 401.285 29.610 401.515 31.040 ;
        RECT 402.005 30.635 402.235 32.470 ;
        RECT 402.490 31.040 403.755 31.270 ;
        RECT 402.005 30.405 403.280 30.635 ;
        RECT 403.525 29.610 403.755 31.040 ;
        RECT 404.245 30.635 404.475 32.470 ;
        RECT 404.730 31.040 405.995 31.270 ;
        RECT 404.245 30.405 405.520 30.635 ;
        RECT 405.765 29.610 405.995 31.040 ;
        RECT 406.485 30.635 406.715 32.470 ;
        RECT 411.745 31.790 411.975 32.470 ;
        RECT 414.165 31.900 414.395 32.470 ;
        RECT 406.970 31.040 408.235 31.270 ;
        RECT 406.485 30.405 407.760 30.635 ;
        RECT 408.005 29.610 408.235 31.040 ;
        RECT 409.180 29.890 409.515 31.790 ;
        RECT 410.830 31.440 411.975 31.790 ;
        RECT 412.425 31.670 414.395 31.900 ;
        RECT 410.830 30.590 411.170 31.440 ;
        RECT 412.425 31.120 412.750 31.670 ;
        RECT 411.430 30.820 412.750 31.120 ;
        RECT 412.990 30.820 413.935 31.230 ;
        RECT 410.830 30.360 411.975 30.590 ;
        RECT 411.745 29.880 411.975 30.360 ;
        RECT 413.560 29.630 413.935 30.820 ;
        RECT 414.165 29.885 414.395 31.670 ;
        RECT 415.445 31.895 415.830 32.470 ;
        RECT 415.445 31.660 417.455 31.895 ;
        RECT 415.445 29.880 415.675 31.660 ;
        RECT 415.905 30.710 416.790 31.270 ;
        RECT 417.170 30.910 417.455 31.660 ;
        RECT 415.905 29.730 416.420 30.710 ;
        RECT 417.685 30.680 418.155 32.460 ;
        RECT 420.425 31.790 420.655 32.460 ;
        RECT 422.665 31.790 422.895 32.460 ;
        RECT 424.905 31.790 425.135 32.460 ;
        RECT 427.045 32.350 427.275 32.460 ;
        RECT 427.045 31.970 427.370 32.350 ;
        RECT 427.045 31.790 427.275 31.970 ;
        RECT 429.385 31.840 429.615 32.460 ;
        RECT 431.625 31.840 431.855 32.460 ;
        RECT 420.425 31.410 427.275 31.790 ;
        RECT 428.805 31.610 431.855 31.840 ;
        RECT 419.580 30.765 422.780 31.110 ;
        RECT 417.530 29.655 418.155 30.680 ;
        RECT 423.480 30.500 424.280 31.410 ;
        RECT 428.805 31.105 429.140 31.610 ;
        RECT 424.850 30.765 429.140 31.105 ;
        RECT 429.610 30.795 432.470 31.230 ;
        RECT 420.325 30.120 427.275 30.500 ;
        RECT 420.325 29.755 420.555 30.120 ;
        RECT 422.565 29.755 422.795 30.120 ;
        RECT 424.805 29.755 425.035 30.120 ;
        RECT 427.015 29.755 427.275 30.120 ;
        RECT 428.805 30.330 429.140 30.765 ;
        RECT 428.805 30.095 431.755 30.330 ;
        RECT 429.285 29.755 429.515 30.095 ;
        RECT 431.525 29.755 431.755 30.095 ;
        RECT 434.370 29.630 434.805 32.460 ;
        RECT 436.860 32.240 438.045 32.470 ;
        RECT 436.860 30.990 437.090 32.240 ;
        RECT 437.815 32.130 438.045 32.240 ;
        RECT 438.855 32.240 441.070 32.470 ;
        RECT 438.855 32.130 439.085 32.240 ;
        RECT 437.320 31.485 437.550 32.010 ;
        RECT 437.815 31.900 439.085 32.130 ;
        RECT 437.320 31.255 439.285 31.485 ;
        RECT 437.320 30.760 437.550 31.255 ;
        RECT 435.050 30.530 437.550 30.760 ;
        RECT 436.400 29.870 436.630 30.530 ;
        RECT 438.075 30.100 438.620 30.910 ;
        RECT 436.985 30.050 438.620 30.100 ;
        RECT 439.525 30.210 439.865 32.010 ;
        RECT 440.160 30.670 440.390 31.605 ;
        RECT 440.840 31.130 441.070 32.240 ;
        RECT 442.200 31.925 442.840 32.155 ;
        RECT 440.840 30.900 441.730 31.130 ;
        RECT 440.160 30.440 441.160 30.670 ;
        RECT 436.985 29.790 438.630 30.050 ;
        RECT 439.525 29.870 440.330 30.210 ;
        RECT 440.930 29.840 441.160 30.440 ;
        RECT 441.390 30.080 441.730 30.900 ;
        RECT 442.610 30.920 442.840 31.925 ;
        RECT 444.285 31.840 444.515 32.210 ;
        RECT 448.365 32.070 449.615 32.300 ;
        RECT 446.885 31.840 447.115 32.035 ;
        RECT 444.285 31.610 447.115 31.840 ;
        RECT 443.125 31.380 443.425 31.605 ;
        RECT 447.905 31.380 448.135 31.840 ;
        RECT 443.125 31.150 448.135 31.380 ;
        RECT 442.610 30.690 446.590 30.920 ;
        RECT 442.125 29.840 442.355 30.670 ;
        RECT 442.950 30.080 443.290 30.690 ;
        RECT 447.005 30.460 447.235 30.670 ;
        RECT 444.050 30.230 447.235 30.460 ;
        RECT 444.050 29.840 444.280 30.230 ;
        RECT 447.585 29.870 447.815 31.150 ;
        RECT 448.365 30.990 448.595 32.070 ;
        RECT 448.825 31.500 449.155 31.840 ;
        RECT 449.385 31.695 449.615 32.070 ;
        RECT 450.665 31.695 451.015 32.295 ;
        RECT 452.705 31.715 452.935 32.305 ;
        RECT 448.825 30.155 449.055 31.500 ;
        RECT 449.385 31.465 451.015 31.695 ;
        RECT 449.360 30.850 450.390 31.230 ;
        RECT 450.785 30.175 451.015 31.465 ;
        RECT 451.245 31.485 452.935 31.715 ;
        RECT 451.245 30.590 451.475 31.485 ;
        RECT 451.710 30.850 453.130 31.230 ;
        RECT 453.710 30.685 454.075 32.400 ;
        RECT 456.065 31.835 456.395 32.460 ;
        RECT 454.370 31.600 456.395 31.835 ;
        RECT 454.370 30.960 454.710 31.600 ;
        RECT 455.050 30.820 455.935 31.230 ;
        RECT 451.245 30.360 453.035 30.590 ;
        RECT 448.650 29.925 449.055 30.155 ;
        RECT 450.510 29.945 451.015 30.175 ;
        RECT 452.805 29.890 453.035 30.360 ;
        RECT 436.985 29.740 438.620 29.790 ;
        RECT 440.930 29.610 444.280 29.840 ;
        RECT 453.710 29.645 454.300 30.685 ;
        RECT 455.560 30.115 455.935 30.820 ;
        RECT 456.165 29.645 456.395 31.600 ;
        RECT 458.190 30.685 458.555 32.400 ;
        RECT 460.545 31.835 460.875 32.460 ;
        RECT 458.850 31.600 460.875 31.835 ;
        RECT 458.850 30.960 459.190 31.600 ;
        RECT 459.530 30.820 460.415 31.230 ;
        RECT 458.190 29.645 458.780 30.685 ;
        RECT 460.040 30.115 460.415 30.820 ;
        RECT 460.645 29.645 460.875 31.600 ;
        RECT 298.405 28.065 298.635 28.405 ;
        RECT 300.645 28.065 300.875 28.405 ;
        RECT 298.405 27.830 301.355 28.065 ;
        RECT 301.020 27.395 301.355 27.830 ;
        RECT 302.885 28.040 303.145 28.405 ;
        RECT 305.125 28.040 305.355 28.405 ;
        RECT 307.365 28.040 307.595 28.405 ;
        RECT 309.605 28.040 309.835 28.405 ;
        RECT 302.885 27.660 309.835 28.040 ;
        RECT 297.690 26.930 300.550 27.365 ;
        RECT 301.020 27.055 305.310 27.395 ;
        RECT 301.020 26.550 301.355 27.055 ;
        RECT 305.880 26.750 306.680 27.660 ;
        RECT 311.845 27.525 313.120 27.755 ;
        RECT 307.380 27.050 310.580 27.395 ;
        RECT 298.305 26.320 301.355 26.550 ;
        RECT 302.885 26.370 309.735 26.750 ;
        RECT 298.305 25.700 298.535 26.320 ;
        RECT 300.545 25.700 300.775 26.320 ;
        RECT 302.885 26.190 303.115 26.370 ;
        RECT 302.790 25.810 303.115 26.190 ;
        RECT 302.885 25.700 303.115 25.810 ;
        RECT 305.025 25.700 305.255 26.370 ;
        RECT 307.265 25.700 307.495 26.370 ;
        RECT 309.505 25.700 309.735 26.370 ;
        RECT 311.845 25.690 312.075 27.525 ;
        RECT 313.365 27.120 313.595 28.550 ;
        RECT 312.330 26.890 313.595 27.120 ;
        RECT 314.085 27.525 315.360 27.755 ;
        RECT 314.085 25.690 314.315 27.525 ;
        RECT 315.605 27.120 315.835 28.550 ;
        RECT 314.570 26.890 315.835 27.120 ;
        RECT 316.885 26.500 317.115 28.280 ;
        RECT 317.345 27.450 317.860 28.430 ;
        RECT 318.970 27.480 319.595 28.505 ;
        RECT 317.345 26.890 318.230 27.450 ;
        RECT 318.610 26.500 318.895 27.250 ;
        RECT 316.885 26.265 318.895 26.500 ;
        RECT 316.885 25.690 317.270 26.265 ;
        RECT 319.125 25.700 319.595 27.480 ;
        RECT 320.645 25.690 320.975 28.550 ;
        RECT 321.205 26.880 321.530 27.880 ;
        RECT 322.485 27.525 323.760 27.755 ;
        RECT 322.485 25.690 322.715 27.525 ;
        RECT 324.005 27.120 324.235 28.550 ;
        RECT 322.970 26.890 324.235 27.120 ;
        RECT 324.725 27.525 326.000 27.755 ;
        RECT 324.725 25.690 324.955 27.525 ;
        RECT 326.245 27.120 326.475 28.550 ;
        RECT 325.210 26.890 326.475 27.120 ;
        RECT 326.965 27.525 328.240 27.755 ;
        RECT 326.965 25.690 327.195 27.525 ;
        RECT 328.485 27.120 328.715 28.550 ;
        RECT 327.450 26.890 328.715 27.120 ;
        RECT 330.990 28.040 331.755 28.470 ;
        RECT 330.990 26.790 331.320 28.040 ;
        RECT 333.415 27.800 333.810 28.550 ;
        RECT 337.510 28.270 337.770 28.430 ;
        RECT 348.040 28.320 351.390 28.550 ;
        RECT 331.585 27.570 333.810 27.800 ;
        RECT 331.585 27.440 332.440 27.570 ;
        RECT 330.990 25.735 331.620 26.790 ;
        RECT 332.980 25.735 333.340 27.340 ;
        RECT 333.580 25.950 333.810 27.570 ;
        RECT 334.040 26.200 334.460 28.005 ;
        RECT 337.500 26.370 337.835 28.270 ;
        RECT 339.285 27.800 339.515 28.270 ;
        RECT 341.305 27.985 341.810 28.215 ;
        RECT 343.265 28.005 343.670 28.235 ;
        RECT 339.285 27.570 341.075 27.800 ;
        RECT 339.320 26.930 340.610 27.310 ;
        RECT 340.845 26.675 341.075 27.570 ;
        RECT 339.385 26.445 341.075 26.675 ;
        RECT 341.305 26.695 341.535 27.985 ;
        RECT 341.930 26.930 342.960 27.310 ;
        RECT 341.305 26.465 342.935 26.695 ;
        RECT 343.265 26.660 343.495 28.005 ;
        RECT 333.580 25.720 334.785 25.950 ;
        RECT 339.385 25.855 339.615 26.445 ;
        RECT 341.305 25.865 341.655 26.465 ;
        RECT 342.705 26.090 342.935 26.465 ;
        RECT 343.165 26.320 343.495 26.660 ;
        RECT 343.725 26.090 343.955 27.170 ;
        RECT 344.505 27.010 344.735 28.290 ;
        RECT 348.040 27.930 348.270 28.320 ;
        RECT 345.085 27.700 348.270 27.930 ;
        RECT 345.085 27.490 345.315 27.700 ;
        RECT 349.030 27.470 349.370 28.080 ;
        RECT 349.965 27.490 350.195 28.320 ;
        RECT 345.730 27.240 349.710 27.470 ;
        RECT 344.185 26.780 349.195 27.010 ;
        RECT 344.185 26.320 344.415 26.780 ;
        RECT 348.895 26.555 349.195 26.780 ;
        RECT 345.205 26.320 348.035 26.550 ;
        RECT 345.205 26.125 345.435 26.320 ;
        RECT 342.705 25.860 343.955 26.090 ;
        RECT 347.805 25.950 348.035 26.320 ;
        RECT 349.480 26.235 349.710 27.240 ;
        RECT 350.590 27.260 350.930 28.080 ;
        RECT 351.160 27.720 351.390 28.320 ;
        RECT 351.990 27.950 352.795 28.290 ;
        RECT 351.160 27.490 352.160 27.720 ;
        RECT 350.590 27.030 351.480 27.260 ;
        RECT 349.480 26.005 350.120 26.235 ;
        RECT 351.250 25.920 351.480 27.030 ;
        RECT 351.930 26.555 352.160 27.490 ;
        RECT 352.455 26.150 352.795 27.950 ;
        RECT 353.700 28.060 355.335 28.420 ;
        RECT 353.700 27.250 354.245 28.060 ;
        RECT 355.690 27.630 355.920 28.290 ;
        RECT 354.770 27.400 357.270 27.630 ;
        RECT 354.770 26.905 355.000 27.400 ;
        RECT 353.035 26.675 355.000 26.905 ;
        RECT 353.235 26.030 354.505 26.260 ;
        RECT 354.770 26.150 355.000 26.675 ;
        RECT 353.235 25.920 353.465 26.030 ;
        RECT 351.250 25.690 353.465 25.920 ;
        RECT 354.275 25.920 354.505 26.030 ;
        RECT 355.230 25.920 355.460 27.170 ;
        RECT 354.275 25.690 355.460 25.920 ;
        RECT 357.515 25.700 357.950 28.530 ;
        RECT 358.325 27.525 359.600 27.755 ;
        RECT 358.325 25.690 358.555 27.525 ;
        RECT 359.845 27.120 360.075 28.550 ;
        RECT 358.810 26.890 360.075 27.120 ;
        RECT 360.565 27.525 361.840 27.755 ;
        RECT 360.565 25.690 360.795 27.525 ;
        RECT 362.085 27.120 362.315 28.550 ;
        RECT 361.050 26.890 362.315 27.120 ;
        RECT 362.805 26.500 363.035 28.280 ;
        RECT 363.265 27.450 363.780 28.430 ;
        RECT 364.890 27.480 365.515 28.505 ;
        RECT 363.265 26.890 364.150 27.450 ;
        RECT 364.530 26.500 364.815 27.250 ;
        RECT 362.805 26.265 364.815 26.500 ;
        RECT 362.805 25.690 363.190 26.265 ;
        RECT 365.045 25.700 365.515 27.480 ;
        RECT 366.165 27.525 367.440 27.755 ;
        RECT 366.165 25.690 366.395 27.525 ;
        RECT 367.685 27.120 367.915 28.550 ;
        RECT 366.650 26.890 367.915 27.120 ;
        RECT 369.365 25.710 369.700 28.480 ;
        RECT 369.930 26.130 370.255 28.110 ;
        RECT 371.205 27.525 372.480 27.755 ;
        RECT 371.205 25.690 371.435 27.525 ;
        RECT 372.725 27.120 372.955 28.550 ;
        RECT 371.690 26.890 372.955 27.120 ;
        RECT 375.685 27.525 376.960 27.755 ;
        RECT 375.685 25.690 375.915 27.525 ;
        RECT 377.205 27.120 377.435 28.550 ;
        RECT 379.825 27.800 380.055 28.280 ;
        RECT 376.170 26.890 377.435 27.120 ;
        RECT 378.910 27.570 380.055 27.800 ;
        RECT 378.910 26.720 379.250 27.570 ;
        RECT 381.640 27.340 382.015 28.530 ;
        RECT 379.510 27.040 380.830 27.340 ;
        RECT 378.910 26.370 380.055 26.720 ;
        RECT 379.825 25.690 380.055 26.370 ;
        RECT 380.505 26.490 380.830 27.040 ;
        RECT 381.070 26.930 382.015 27.340 ;
        RECT 382.245 26.490 382.475 28.275 ;
        RECT 380.505 26.260 382.475 26.490 ;
        RECT 382.245 25.690 382.475 26.260 ;
        RECT 382.965 27.525 384.240 27.755 ;
        RECT 382.965 25.690 383.195 27.525 ;
        RECT 384.485 27.120 384.715 28.550 ;
        RECT 383.450 26.890 384.715 27.120 ;
        RECT 385.205 27.525 386.480 27.755 ;
        RECT 385.205 25.690 385.435 27.525 ;
        RECT 386.725 27.120 386.955 28.550 ;
        RECT 385.690 26.890 386.955 27.120 ;
        RECT 388.725 27.480 389.350 28.505 ;
        RECT 388.725 25.700 389.195 27.480 ;
        RECT 390.460 27.450 390.975 28.430 ;
        RECT 389.425 26.500 389.710 27.250 ;
        RECT 390.090 26.890 390.975 27.450 ;
        RECT 391.205 26.500 391.435 28.280 ;
        RECT 389.425 26.265 391.435 26.500 ;
        RECT 391.050 25.690 391.435 26.265 ;
        RECT 391.925 27.525 393.200 27.755 ;
        RECT 391.925 25.690 392.155 27.525 ;
        RECT 393.445 27.120 393.675 28.550 ;
        RECT 392.410 26.890 393.675 27.120 ;
        RECT 394.165 27.525 395.440 27.755 ;
        RECT 394.165 25.690 394.395 27.525 ;
        RECT 395.685 27.120 395.915 28.550 ;
        RECT 394.650 26.890 395.915 27.120 ;
        RECT 396.405 27.525 397.680 27.755 ;
        RECT 396.405 25.690 396.635 27.525 ;
        RECT 397.925 27.120 398.155 28.550 ;
        RECT 396.890 26.890 398.155 27.120 ;
        RECT 398.645 27.525 399.920 27.755 ;
        RECT 398.645 25.690 398.875 27.525 ;
        RECT 400.165 27.120 400.395 28.550 ;
        RECT 399.130 26.890 400.395 27.120 ;
        RECT 400.885 27.525 402.160 27.755 ;
        RECT 400.885 25.690 401.115 27.525 ;
        RECT 402.405 27.120 402.635 28.550 ;
        RECT 401.370 26.890 402.635 27.120 ;
        RECT 403.125 27.525 404.400 27.755 ;
        RECT 403.125 25.690 403.355 27.525 ;
        RECT 404.645 27.120 404.875 28.550 ;
        RECT 403.610 26.890 404.875 27.120 ;
        RECT 405.365 27.525 406.640 27.755 ;
        RECT 405.365 25.690 405.595 27.525 ;
        RECT 406.885 27.120 407.115 28.550 ;
        RECT 409.505 27.800 409.735 28.280 ;
        RECT 405.850 26.890 407.115 27.120 ;
        RECT 408.590 27.570 409.735 27.800 ;
        RECT 408.590 26.720 408.930 27.570 ;
        RECT 411.320 27.340 411.695 28.530 ;
        RECT 409.190 27.040 410.510 27.340 ;
        RECT 408.590 26.370 409.735 26.720 ;
        RECT 409.505 25.690 409.735 26.370 ;
        RECT 410.185 26.490 410.510 27.040 ;
        RECT 410.750 26.930 411.695 27.340 ;
        RECT 411.925 26.490 412.155 28.275 ;
        RECT 410.185 26.260 412.155 26.490 ;
        RECT 411.925 25.690 412.155 26.260 ;
        RECT 414.990 28.040 415.755 28.470 ;
        RECT 414.990 26.790 415.320 28.040 ;
        RECT 417.415 27.800 417.810 28.550 ;
        RECT 421.020 28.210 422.360 28.530 ;
        RECT 415.585 27.570 417.810 27.800 ;
        RECT 415.585 27.440 416.440 27.570 ;
        RECT 414.990 25.735 415.620 26.790 ;
        RECT 416.980 25.735 417.340 27.340 ;
        RECT 417.580 25.950 417.810 27.570 ;
        RECT 418.040 26.200 418.460 28.005 ;
        RECT 419.785 27.310 420.125 27.920 ;
        RECT 420.920 27.310 421.260 27.920 ;
        RECT 419.785 26.930 420.690 27.310 ;
        RECT 420.920 26.930 421.825 27.310 ;
        RECT 417.580 25.720 418.785 25.950 ;
        RECT 421.030 25.920 421.370 26.585 ;
        RECT 422.055 26.355 422.360 28.210 ;
        RECT 424.965 28.065 425.195 28.405 ;
        RECT 427.205 28.065 427.435 28.405 ;
        RECT 439.525 28.065 439.755 28.405 ;
        RECT 441.765 28.065 441.995 28.405 ;
        RECT 422.590 27.310 422.940 27.920 ;
        RECT 424.965 27.830 427.915 28.065 ;
        RECT 439.525 27.830 442.475 28.065 ;
        RECT 427.580 27.395 427.915 27.830 ;
        RECT 442.140 27.395 442.475 27.830 ;
        RECT 422.590 26.930 423.485 27.310 ;
        RECT 424.250 26.930 427.110 27.365 ;
        RECT 427.580 27.055 431.870 27.395 ;
        RECT 423.070 25.920 423.410 26.585 ;
        RECT 427.580 26.550 427.915 27.055 ;
        RECT 433.940 27.050 437.140 27.395 ;
        RECT 438.810 26.930 441.670 27.365 ;
        RECT 442.140 27.055 446.430 27.395 ;
        RECT 442.140 26.550 442.475 27.055 ;
        RECT 448.500 27.050 451.700 27.395 ;
        RECT 421.030 25.690 423.410 25.920 ;
        RECT 424.865 26.320 427.915 26.550 ;
        RECT 439.425 26.320 442.475 26.550 ;
        RECT 424.865 25.700 425.095 26.320 ;
        RECT 427.105 25.700 427.335 26.320 ;
        RECT 439.425 25.700 439.655 26.320 ;
        RECT 441.665 25.700 441.895 26.320 ;
        RECT 454.545 25.760 454.850 27.900 ;
        RECT 455.080 26.720 455.435 28.480 ;
        RECT 455.665 27.290 455.970 28.480 ;
        RECT 457.630 27.475 458.220 28.515 ;
        RECT 455.665 26.950 456.695 27.290 ;
        RECT 455.080 26.400 456.505 26.720 ;
        RECT 456.225 25.700 456.505 26.400 ;
        RECT 457.630 25.760 457.995 27.475 ;
        RECT 459.480 27.340 459.855 28.045 ;
        RECT 458.290 26.560 458.630 27.200 ;
        RECT 458.970 26.930 459.855 27.340 ;
        RECT 460.085 26.560 460.315 28.515 ;
        RECT 458.290 26.325 460.315 26.560 ;
        RECT 459.985 25.700 460.315 26.325 ;
        RECT 170.750 22.950 189.320 23.250 ;
        RECT 170.750 22.350 171.130 22.950 ;
        RECT 172.990 22.350 173.370 22.950 ;
        RECT 175.230 22.350 175.610 22.950 ;
        RECT 177.470 22.350 177.850 22.950 ;
        RECT 180.830 22.350 181.210 22.950 ;
        RECT 183.070 22.350 183.450 22.950 ;
        RECT 185.310 22.350 185.690 22.950 ;
        RECT 187.550 22.350 187.930 22.950 ;
        RECT 297.285 22.795 297.515 24.630 ;
        RECT 297.770 23.200 299.035 23.430 ;
        RECT 297.285 22.565 298.560 22.795 ;
        RECT 298.805 21.770 299.035 23.200 ;
        RECT 299.525 22.795 299.755 24.630 ;
        RECT 300.010 23.200 301.275 23.430 ;
        RECT 299.525 22.565 300.800 22.795 ;
        RECT 301.045 21.770 301.275 23.200 ;
        RECT 301.765 22.795 301.995 24.630 ;
        RECT 302.250 23.200 303.515 23.430 ;
        RECT 301.765 22.565 303.040 22.795 ;
        RECT 303.285 21.770 303.515 23.200 ;
        RECT 304.005 22.795 304.235 24.630 ;
        RECT 304.490 23.200 305.755 23.430 ;
        RECT 304.005 22.565 305.280 22.795 ;
        RECT 305.525 21.770 305.755 23.200 ;
        RECT 306.245 22.795 306.475 24.630 ;
        RECT 306.730 23.200 307.995 23.430 ;
        RECT 306.245 22.565 307.520 22.795 ;
        RECT 307.765 21.770 307.995 23.200 ;
        RECT 308.485 22.795 308.715 24.630 ;
        RECT 308.970 23.200 310.235 23.430 ;
        RECT 308.485 22.565 309.760 22.795 ;
        RECT 310.005 21.770 310.235 23.200 ;
        RECT 310.725 22.795 310.955 24.630 ;
        RECT 311.210 23.200 312.475 23.430 ;
        RECT 310.725 22.565 312.000 22.795 ;
        RECT 312.245 21.770 312.475 23.200 ;
        RECT 312.965 22.795 313.195 24.630 ;
        RECT 313.450 23.200 314.715 23.430 ;
        RECT 312.965 22.565 314.240 22.795 ;
        RECT 314.485 21.770 314.715 23.200 ;
        RECT 316.885 22.795 317.115 24.630 ;
        RECT 317.370 23.200 318.635 23.430 ;
        RECT 316.885 22.565 318.160 22.795 ;
        RECT 318.405 21.770 318.635 23.200 ;
        RECT 319.125 22.795 319.355 24.630 ;
        RECT 319.610 23.200 320.875 23.430 ;
        RECT 319.125 22.565 320.400 22.795 ;
        RECT 320.645 21.770 320.875 23.200 ;
        RECT 321.365 22.795 321.595 24.630 ;
        RECT 321.850 23.200 323.115 23.430 ;
        RECT 321.365 22.565 322.640 22.795 ;
        RECT 322.885 21.770 323.115 23.200 ;
        RECT 323.605 22.795 323.835 24.630 ;
        RECT 324.090 23.200 325.355 23.430 ;
        RECT 323.605 22.565 324.880 22.795 ;
        RECT 325.125 21.770 325.355 23.200 ;
        RECT 325.845 22.795 326.075 24.630 ;
        RECT 326.330 23.200 327.595 23.430 ;
        RECT 325.845 22.565 327.120 22.795 ;
        RECT 327.365 21.770 327.595 23.200 ;
        RECT 328.085 22.795 328.315 24.630 ;
        RECT 328.570 23.200 329.835 23.430 ;
        RECT 328.085 22.565 329.360 22.795 ;
        RECT 329.605 21.770 329.835 23.200 ;
        RECT 330.325 22.795 330.555 24.630 ;
        RECT 333.575 23.920 333.855 24.620 ;
        RECT 333.575 23.600 335.000 23.920 ;
        RECT 330.810 23.200 332.075 23.430 ;
        RECT 330.325 22.565 331.600 22.795 ;
        RECT 331.845 21.770 332.075 23.200 ;
        RECT 333.385 23.030 334.415 23.370 ;
        RECT 334.110 21.840 334.415 23.030 ;
        RECT 334.645 21.840 335.000 23.600 ;
        RECT 335.230 22.420 335.535 24.560 ;
        RECT 337.500 22.050 337.835 23.950 ;
        RECT 338.725 22.795 338.955 24.630 ;
        RECT 339.210 23.200 340.475 23.430 ;
        RECT 338.725 22.565 340.000 22.795 ;
        RECT 340.245 21.770 340.475 23.200 ;
        RECT 340.965 22.795 341.195 24.630 ;
        RECT 341.450 23.200 342.715 23.430 ;
        RECT 340.965 22.565 342.240 22.795 ;
        RECT 342.485 21.770 342.715 23.200 ;
        RECT 343.605 21.840 343.940 24.610 ;
        RECT 347.110 24.400 349.490 24.630 ;
        RECT 344.170 22.210 344.495 24.190 ;
        RECT 347.110 23.735 347.450 24.400 ;
        RECT 345.865 23.010 346.770 23.390 ;
        RECT 347.000 23.010 347.905 23.390 ;
        RECT 345.865 22.400 346.205 23.010 ;
        RECT 347.000 22.400 347.340 23.010 ;
        RECT 348.135 22.110 348.440 23.965 ;
        RECT 349.150 23.735 349.490 24.400 ;
        RECT 348.670 23.010 349.565 23.390 ;
        RECT 348.670 22.400 349.020 23.010 ;
        RECT 347.100 21.790 348.440 22.110 ;
        RECT 350.940 22.050 351.275 23.950 ;
        RECT 352.165 22.795 352.395 24.630 ;
        RECT 352.650 23.200 353.915 23.430 ;
        RECT 352.165 22.565 353.440 22.795 ;
        RECT 350.950 21.890 351.210 22.050 ;
        RECT 353.685 21.770 353.915 23.200 ;
        RECT 356.085 22.795 356.315 24.630 ;
        RECT 356.570 23.200 357.835 23.430 ;
        RECT 356.085 22.565 357.360 22.795 ;
        RECT 357.605 21.770 357.835 23.200 ;
        RECT 358.325 22.795 358.555 24.630 ;
        RECT 358.810 23.200 360.075 23.430 ;
        RECT 358.325 22.565 359.600 22.795 ;
        RECT 359.845 21.770 360.075 23.200 ;
        RECT 360.565 22.795 360.795 24.630 ;
        RECT 361.050 23.200 362.315 23.430 ;
        RECT 360.565 22.565 361.840 22.795 ;
        RECT 362.085 21.770 362.315 23.200 ;
        RECT 362.805 22.795 363.035 24.630 ;
        RECT 363.290 23.200 364.555 23.430 ;
        RECT 362.805 22.565 364.080 22.795 ;
        RECT 364.325 21.770 364.555 23.200 ;
        RECT 365.045 22.795 365.275 24.630 ;
        RECT 365.530 23.200 366.795 23.430 ;
        RECT 365.045 22.565 366.320 22.795 ;
        RECT 366.565 21.770 366.795 23.200 ;
        RECT 367.285 22.795 367.515 24.630 ;
        RECT 367.770 23.200 369.035 23.430 ;
        RECT 367.285 22.565 368.560 22.795 ;
        RECT 368.805 21.770 369.035 23.200 ;
        RECT 369.525 22.795 369.755 24.630 ;
        RECT 370.010 23.200 371.275 23.430 ;
        RECT 369.525 22.565 370.800 22.795 ;
        RECT 371.045 21.770 371.275 23.200 ;
        RECT 371.765 22.795 371.995 24.630 ;
        RECT 372.250 23.200 373.515 23.430 ;
        RECT 371.765 22.565 373.040 22.795 ;
        RECT 373.285 21.770 373.515 23.200 ;
        RECT 374.005 22.795 374.235 24.630 ;
        RECT 374.490 23.200 375.755 23.430 ;
        RECT 374.005 22.565 375.280 22.795 ;
        RECT 375.525 21.770 375.755 23.200 ;
        RECT 376.245 22.795 376.475 24.630 ;
        RECT 376.730 23.200 377.995 23.430 ;
        RECT 376.245 22.565 377.520 22.795 ;
        RECT 377.765 21.770 377.995 23.200 ;
        RECT 378.485 22.795 378.715 24.630 ;
        RECT 378.970 23.200 380.235 23.430 ;
        RECT 378.485 22.565 379.760 22.795 ;
        RECT 380.005 21.770 380.235 23.200 ;
        RECT 380.725 22.795 380.955 24.630 ;
        RECT 384.655 24.000 384.995 24.620 ;
        RECT 386.220 24.385 389.075 24.620 ;
        RECT 386.220 24.000 386.450 24.385 ;
        RECT 384.655 23.770 386.450 24.000 ;
        RECT 386.750 23.620 388.290 23.950 ;
        RECT 388.735 23.770 389.075 24.385 ;
        RECT 381.210 23.200 382.475 23.430 ;
        RECT 380.725 22.565 382.000 22.795 ;
        RECT 382.245 21.770 382.475 23.200 ;
        RECT 385.010 23.010 385.970 23.390 ;
        RECT 385.010 22.325 385.405 23.010 ;
        RECT 386.200 21.790 386.520 23.390 ;
        RECT 386.750 21.825 387.080 23.620 ;
        RECT 387.320 21.790 387.640 23.390 ;
        RECT 387.880 23.040 388.945 23.390 ;
        RECT 387.880 21.790 388.200 23.040 ;
        RECT 390.145 22.210 390.470 24.190 ;
        RECT 390.700 21.840 391.035 24.610 ;
        RECT 391.925 22.795 392.155 24.630 ;
        RECT 392.410 23.200 393.675 23.430 ;
        RECT 391.925 22.565 393.200 22.795 ;
        RECT 393.445 21.770 393.675 23.200 ;
        RECT 395.285 22.795 395.515 24.630 ;
        RECT 395.770 23.200 397.035 23.430 ;
        RECT 395.285 22.565 396.560 22.795 ;
        RECT 396.805 21.770 397.035 23.200 ;
        RECT 397.525 22.795 397.755 24.630 ;
        RECT 398.010 23.200 399.275 23.430 ;
        RECT 397.525 22.565 398.800 22.795 ;
        RECT 399.045 21.770 399.275 23.200 ;
        RECT 399.765 22.795 399.995 24.630 ;
        RECT 400.250 23.200 401.515 23.430 ;
        RECT 399.765 22.565 401.040 22.795 ;
        RECT 401.285 21.770 401.515 23.200 ;
        RECT 402.005 22.795 402.235 24.630 ;
        RECT 402.490 23.200 403.755 23.430 ;
        RECT 402.005 22.565 403.280 22.795 ;
        RECT 403.525 21.770 403.755 23.200 ;
        RECT 404.245 22.795 404.475 24.630 ;
        RECT 404.730 23.200 405.995 23.430 ;
        RECT 404.245 22.565 405.520 22.795 ;
        RECT 405.765 21.770 405.995 23.200 ;
        RECT 406.485 22.795 406.715 24.630 ;
        RECT 406.970 23.200 408.235 23.430 ;
        RECT 406.485 22.565 407.760 22.795 ;
        RECT 408.005 21.770 408.235 23.200 ;
        RECT 408.725 22.795 408.955 24.630 ;
        RECT 409.210 23.200 410.475 23.430 ;
        RECT 408.725 22.565 410.000 22.795 ;
        RECT 410.245 21.770 410.475 23.200 ;
        RECT 410.965 22.795 411.195 24.630 ;
        RECT 411.450 23.200 412.715 23.430 ;
        RECT 410.965 22.565 412.240 22.795 ;
        RECT 412.485 21.770 412.715 23.200 ;
        RECT 413.205 22.795 413.435 24.630 ;
        RECT 413.690 23.200 414.955 23.430 ;
        RECT 413.205 22.565 414.480 22.795 ;
        RECT 414.725 21.770 414.955 23.200 ;
        RECT 415.445 22.795 415.675 24.630 ;
        RECT 415.930 23.200 417.195 23.430 ;
        RECT 415.445 22.565 416.720 22.795 ;
        RECT 416.965 21.770 417.195 23.200 ;
        RECT 418.405 22.840 418.875 24.620 ;
        RECT 420.730 24.055 421.115 24.630 ;
        RECT 419.105 23.820 421.115 24.055 ;
        RECT 419.105 23.070 419.390 23.820 ;
        RECT 419.770 22.870 420.655 23.430 ;
        RECT 418.405 21.815 419.030 22.840 ;
        RECT 420.140 21.890 420.655 22.870 ;
        RECT 420.885 22.040 421.115 23.820 ;
        RECT 421.605 24.055 421.990 24.630 ;
        RECT 421.605 23.820 423.615 24.055 ;
        RECT 421.605 22.040 421.835 23.820 ;
        RECT 422.065 22.870 422.950 23.430 ;
        RECT 423.330 23.070 423.615 23.820 ;
        RECT 422.065 21.890 422.580 22.870 ;
        RECT 423.845 22.840 424.315 24.620 ;
        RECT 427.425 23.950 427.655 24.630 ;
        RECT 429.845 24.060 430.075 24.630 ;
        RECT 423.690 21.815 424.315 22.840 ;
        RECT 426.510 23.600 427.655 23.950 ;
        RECT 428.105 23.830 430.075 24.060 ;
        RECT 434.485 24.055 434.870 24.630 ;
        RECT 426.510 22.750 426.850 23.600 ;
        RECT 428.105 23.280 428.430 23.830 ;
        RECT 427.110 22.980 428.430 23.280 ;
        RECT 428.670 22.980 429.615 23.390 ;
        RECT 426.510 22.520 427.655 22.750 ;
        RECT 427.425 22.040 427.655 22.520 ;
        RECT 429.240 21.790 429.615 22.980 ;
        RECT 429.845 22.045 430.075 23.830 ;
        RECT 432.140 22.050 432.475 23.950 ;
        RECT 434.485 23.820 436.495 24.055 ;
        RECT 432.150 21.890 432.410 22.050 ;
        RECT 434.485 22.040 434.715 23.820 ;
        RECT 434.945 22.870 435.830 23.430 ;
        RECT 436.210 23.070 436.495 23.820 ;
        RECT 434.945 21.890 435.460 22.870 ;
        RECT 436.725 22.840 437.195 24.620 ;
        RECT 436.570 21.815 437.195 22.840 ;
        RECT 438.865 22.420 439.170 24.560 ;
        RECT 440.545 23.920 440.825 24.620 ;
        RECT 439.400 23.600 440.825 23.920 ;
        RECT 439.400 21.840 439.755 23.600 ;
        RECT 439.985 23.030 441.015 23.370 ;
        RECT 439.985 21.840 440.290 23.030 ;
        RECT 442.210 21.790 442.645 24.620 ;
        RECT 444.700 24.400 445.885 24.630 ;
        RECT 444.700 23.150 444.930 24.400 ;
        RECT 445.655 24.290 445.885 24.400 ;
        RECT 446.695 24.400 448.910 24.630 ;
        RECT 446.695 24.290 446.925 24.400 ;
        RECT 445.160 23.645 445.390 24.170 ;
        RECT 445.655 24.060 446.925 24.290 ;
        RECT 445.160 23.415 447.125 23.645 ;
        RECT 445.160 22.920 445.390 23.415 ;
        RECT 442.890 22.690 445.390 22.920 ;
        RECT 444.240 22.030 444.470 22.690 ;
        RECT 445.915 22.260 446.460 23.070 ;
        RECT 444.825 22.210 446.460 22.260 ;
        RECT 447.365 22.370 447.705 24.170 ;
        RECT 448.000 22.830 448.230 23.765 ;
        RECT 448.680 23.290 448.910 24.400 ;
        RECT 450.040 24.085 450.680 24.315 ;
        RECT 448.680 23.060 449.570 23.290 ;
        RECT 448.000 22.600 449.000 22.830 ;
        RECT 444.825 21.950 446.470 22.210 ;
        RECT 447.365 22.030 448.170 22.370 ;
        RECT 448.770 22.000 449.000 22.600 ;
        RECT 449.230 22.240 449.570 23.060 ;
        RECT 450.450 23.080 450.680 24.085 ;
        RECT 452.125 24.000 452.355 24.370 ;
        RECT 456.205 24.230 457.455 24.460 ;
        RECT 454.725 24.000 454.955 24.195 ;
        RECT 452.125 23.770 454.955 24.000 ;
        RECT 450.965 23.540 451.265 23.765 ;
        RECT 455.745 23.540 455.975 24.000 ;
        RECT 450.965 23.310 455.975 23.540 ;
        RECT 450.450 22.850 454.430 23.080 ;
        RECT 449.965 22.000 450.195 22.830 ;
        RECT 450.790 22.240 451.130 22.850 ;
        RECT 454.845 22.620 455.075 22.830 ;
        RECT 451.890 22.390 455.075 22.620 ;
        RECT 451.890 22.000 452.120 22.390 ;
        RECT 455.425 22.030 455.655 23.310 ;
        RECT 456.205 23.150 456.435 24.230 ;
        RECT 456.665 23.660 456.995 24.000 ;
        RECT 457.225 23.855 457.455 24.230 ;
        RECT 458.505 23.855 458.855 24.455 ;
        RECT 460.545 23.875 460.775 24.465 ;
        RECT 456.665 22.315 456.895 23.660 ;
        RECT 457.225 23.625 458.855 23.855 ;
        RECT 457.200 23.010 458.230 23.390 ;
        RECT 458.625 22.335 458.855 23.625 ;
        RECT 459.085 23.645 460.775 23.875 ;
        RECT 459.085 22.750 459.315 23.645 ;
        RECT 459.550 23.010 460.840 23.390 ;
        RECT 459.085 22.520 460.875 22.750 ;
        RECT 456.490 22.085 456.895 22.315 ;
        RECT 458.350 22.105 458.855 22.335 ;
        RECT 460.645 22.050 460.875 22.520 ;
        RECT 444.825 21.900 446.460 21.950 ;
        RECT 448.770 21.770 452.120 22.000 ;
        RECT 297.385 20.080 297.900 20.690 ;
        RECT 301.090 20.480 305.270 20.710 ;
        RECT 297.385 19.050 297.775 20.080 ;
        RECT 299.240 19.740 299.470 20.435 ;
        RECT 301.090 19.845 301.320 20.480 ;
        RECT 305.040 20.450 305.270 20.480 ;
        RECT 306.160 20.480 309.090 20.710 ;
        RECT 302.705 20.020 304.645 20.250 ;
        RECT 305.040 20.110 305.930 20.450 ;
        RECT 298.080 19.400 299.470 19.740 ;
        RECT 299.865 19.610 301.320 19.845 ;
        RECT 299.240 19.380 299.470 19.400 ;
        RECT 299.240 19.135 301.445 19.380 ;
        RECT 297.385 17.860 298.155 19.050 ;
        RECT 299.240 17.860 299.470 19.135 ;
        RECT 301.915 19.090 303.110 19.470 ;
        RECT 303.340 18.700 303.570 20.020 ;
        RECT 301.600 18.465 303.570 18.700 ;
        RECT 305.040 18.690 305.270 20.110 ;
        RECT 306.160 19.625 306.390 20.480 ;
        RECT 306.985 19.160 307.325 20.250 ;
        RECT 308.860 19.935 309.090 20.480 ;
        RECT 308.860 19.705 311.200 19.935 ;
        RECT 311.525 19.475 311.855 20.450 ;
        RECT 308.965 19.245 311.855 19.475 ;
        RECT 301.600 18.355 301.830 18.465 ;
        RECT 303.340 18.395 303.570 18.465 ;
        RECT 304.305 18.460 305.270 18.690 ;
        RECT 305.555 19.015 308.165 19.160 ;
        RECT 305.555 18.930 310.185 19.015 ;
        RECT 305.555 18.460 305.895 18.930 ;
        RECT 307.825 18.785 310.185 18.930 ;
        RECT 306.125 18.465 307.515 18.700 ;
        RECT 306.125 18.175 306.355 18.465 ;
        RECT 304.885 17.945 306.355 18.175 ;
        RECT 307.285 18.080 307.515 18.465 ;
        RECT 307.825 18.310 308.165 18.785 ;
        RECT 310.745 18.255 311.085 19.000 ;
        RECT 311.625 18.255 311.855 19.245 ;
        RECT 308.700 18.080 311.085 18.255 ;
        RECT 307.285 18.025 311.085 18.080 ;
        RECT 312.085 18.080 312.315 19.310 ;
        RECT 312.590 18.310 312.930 20.450 ;
        RECT 314.485 20.090 314.815 20.430 ;
        RECT 313.170 19.090 314.310 19.470 ;
        RECT 314.580 18.860 314.815 20.090 ;
        RECT 316.725 19.960 316.955 20.430 ;
        RECT 313.160 18.625 314.815 18.860 ;
        RECT 315.110 19.730 316.955 19.960 ;
        RECT 315.110 18.880 315.340 19.730 ;
        RECT 317.445 19.685 318.720 19.915 ;
        RECT 315.610 19.410 316.920 19.475 ;
        RECT 315.610 19.150 317.110 19.410 ;
        RECT 315.610 19.110 316.920 19.150 ;
        RECT 315.110 18.645 316.855 18.880 ;
        RECT 313.160 18.080 313.390 18.625 ;
        RECT 307.285 17.850 308.930 18.025 ;
        RECT 312.085 17.850 313.390 18.080 ;
        RECT 314.585 18.015 314.815 18.625 ;
        RECT 316.625 18.015 316.855 18.645 ;
        RECT 317.445 17.850 317.675 19.685 ;
        RECT 318.965 19.280 319.195 20.710 ;
        RECT 317.930 19.050 319.195 19.280 ;
        RECT 319.685 19.685 320.960 19.915 ;
        RECT 319.685 17.850 319.915 19.685 ;
        RECT 321.205 19.280 321.435 20.710 ;
        RECT 324.040 20.370 325.380 20.690 ;
        RECT 323.460 19.470 323.810 20.080 ;
        RECT 320.170 19.050 321.435 19.280 ;
        RECT 322.915 19.090 323.810 19.470 ;
        RECT 322.990 18.080 323.330 18.745 ;
        RECT 324.040 18.515 324.345 20.370 ;
        RECT 325.140 19.470 325.480 20.080 ;
        RECT 326.275 19.470 326.615 20.080 ;
        RECT 324.575 19.090 325.480 19.470 ;
        RECT 325.710 19.090 326.615 19.470 ;
        RECT 327.525 19.685 328.800 19.915 ;
        RECT 325.030 18.080 325.370 18.745 ;
        RECT 322.990 17.850 325.370 18.080 ;
        RECT 327.525 17.850 327.755 19.685 ;
        RECT 329.045 19.280 329.275 20.710 ;
        RECT 328.010 19.050 329.275 19.280 ;
        RECT 329.765 19.685 331.040 19.915 ;
        RECT 329.765 17.850 329.995 19.685 ;
        RECT 331.285 19.280 331.515 20.710 ;
        RECT 330.250 19.050 331.515 19.280 ;
        RECT 332.005 19.685 333.280 19.915 ;
        RECT 332.005 17.850 332.235 19.685 ;
        RECT 333.525 19.280 333.755 20.710 ;
        RECT 332.490 19.050 333.755 19.280 ;
        RECT 336.485 19.685 337.760 19.915 ;
        RECT 336.485 17.850 336.715 19.685 ;
        RECT 338.005 19.280 338.235 20.710 ;
        RECT 336.970 19.050 338.235 19.280 ;
        RECT 338.725 19.685 340.000 19.915 ;
        RECT 338.725 17.850 338.955 19.685 ;
        RECT 340.245 19.280 340.475 20.710 ;
        RECT 339.210 19.050 340.475 19.280 ;
        RECT 340.965 19.685 342.240 19.915 ;
        RECT 340.965 17.850 341.195 19.685 ;
        RECT 342.485 19.280 342.715 20.710 ;
        RECT 341.450 19.050 342.715 19.280 ;
        RECT 343.205 19.685 344.480 19.915 ;
        RECT 343.205 17.850 343.435 19.685 ;
        RECT 344.725 19.280 344.955 20.710 ;
        RECT 343.690 19.050 344.955 19.280 ;
        RECT 345.445 19.685 346.720 19.915 ;
        RECT 345.445 17.850 345.675 19.685 ;
        RECT 346.965 19.280 347.195 20.710 ;
        RECT 345.930 19.050 347.195 19.280 ;
        RECT 347.685 19.685 348.960 19.915 ;
        RECT 347.685 17.850 347.915 19.685 ;
        RECT 349.205 19.280 349.435 20.710 ;
        RECT 348.170 19.050 349.435 19.280 ;
        RECT 349.925 19.685 351.200 19.915 ;
        RECT 349.925 17.850 350.155 19.685 ;
        RECT 351.445 19.280 351.675 20.710 ;
        RECT 350.410 19.050 351.675 19.280 ;
        RECT 352.165 19.685 353.440 19.915 ;
        RECT 352.165 17.850 352.395 19.685 ;
        RECT 353.685 19.280 353.915 20.710 ;
        RECT 352.650 19.050 353.915 19.280 ;
        RECT 354.405 19.685 355.680 19.915 ;
        RECT 354.405 17.850 354.635 19.685 ;
        RECT 355.925 19.280 356.155 20.710 ;
        RECT 354.890 19.050 356.155 19.280 ;
        RECT 356.645 19.685 357.920 19.915 ;
        RECT 356.645 17.850 356.875 19.685 ;
        RECT 358.165 19.280 358.395 20.710 ;
        RECT 357.130 19.050 358.395 19.280 ;
        RECT 358.885 19.685 360.160 19.915 ;
        RECT 358.885 17.850 359.115 19.685 ;
        RECT 360.405 19.280 360.635 20.710 ;
        RECT 359.370 19.050 360.635 19.280 ;
        RECT 361.125 19.685 362.400 19.915 ;
        RECT 361.125 17.850 361.355 19.685 ;
        RECT 362.645 19.280 362.875 20.710 ;
        RECT 361.610 19.050 362.875 19.280 ;
        RECT 365.045 18.660 365.275 20.440 ;
        RECT 365.505 19.610 366.020 20.590 ;
        RECT 367.130 19.640 367.755 20.665 ;
        RECT 365.505 19.050 366.390 19.610 ;
        RECT 366.770 18.660 367.055 19.410 ;
        RECT 365.045 18.425 367.055 18.660 ;
        RECT 365.045 17.850 365.430 18.425 ;
        RECT 367.285 17.860 367.755 19.640 ;
        RECT 368.805 17.870 369.140 20.640 ;
        RECT 369.370 18.290 369.695 20.270 ;
        RECT 370.645 19.685 371.920 19.915 ;
        RECT 370.645 17.850 370.875 19.685 ;
        RECT 372.165 19.280 372.395 20.710 ;
        RECT 371.130 19.050 372.395 19.280 ;
        RECT 375.685 19.685 376.960 19.915 ;
        RECT 375.685 17.850 375.915 19.685 ;
        RECT 377.205 19.280 377.435 20.710 ;
        RECT 376.170 19.050 377.435 19.280 ;
        RECT 377.925 19.685 379.200 19.915 ;
        RECT 377.925 17.850 378.155 19.685 ;
        RECT 379.445 19.280 379.675 20.710 ;
        RECT 382.280 19.440 382.600 20.690 ;
        RECT 378.410 19.050 379.675 19.280 ;
        RECT 381.535 19.090 382.600 19.440 ;
        RECT 382.840 19.090 383.160 20.690 ;
        RECT 383.400 18.860 383.730 20.655 ;
        RECT 383.960 19.090 384.280 20.690 ;
        RECT 385.075 19.470 385.470 20.155 ;
        RECT 384.510 19.090 385.470 19.470 ;
        RECT 386.325 19.685 387.600 19.915 ;
        RECT 381.405 18.095 381.745 18.710 ;
        RECT 382.190 18.530 383.730 18.860 ;
        RECT 384.030 18.480 385.825 18.710 ;
        RECT 384.030 18.095 384.260 18.480 ;
        RECT 381.405 17.860 384.260 18.095 ;
        RECT 385.485 17.860 385.825 18.480 ;
        RECT 386.325 17.850 386.555 19.685 ;
        RECT 387.845 19.280 388.075 20.710 ;
        RECT 397.880 20.480 401.230 20.710 ;
        RECT 389.125 19.960 389.355 20.430 ;
        RECT 391.145 20.145 391.650 20.375 ;
        RECT 393.105 20.165 393.510 20.395 ;
        RECT 389.125 19.730 390.915 19.960 ;
        RECT 386.810 19.050 388.075 19.280 ;
        RECT 389.160 19.090 390.450 19.470 ;
        RECT 390.685 18.835 390.915 19.730 ;
        RECT 389.225 18.605 390.915 18.835 ;
        RECT 391.145 18.855 391.375 20.145 ;
        RECT 391.770 19.090 392.800 19.470 ;
        RECT 391.145 18.625 392.775 18.855 ;
        RECT 393.105 18.820 393.335 20.165 ;
        RECT 389.225 18.015 389.455 18.605 ;
        RECT 391.145 18.025 391.495 18.625 ;
        RECT 392.545 18.250 392.775 18.625 ;
        RECT 393.005 18.480 393.335 18.820 ;
        RECT 393.565 18.250 393.795 19.330 ;
        RECT 394.345 19.170 394.575 20.450 ;
        RECT 397.880 20.090 398.110 20.480 ;
        RECT 394.925 19.860 398.110 20.090 ;
        RECT 394.925 19.650 395.155 19.860 ;
        RECT 398.870 19.630 399.210 20.240 ;
        RECT 399.805 19.650 400.035 20.480 ;
        RECT 395.570 19.400 399.550 19.630 ;
        RECT 394.025 18.940 399.035 19.170 ;
        RECT 394.025 18.480 394.255 18.940 ;
        RECT 398.735 18.715 399.035 18.940 ;
        RECT 395.045 18.480 397.875 18.710 ;
        RECT 395.045 18.285 395.275 18.480 ;
        RECT 392.545 18.020 393.795 18.250 ;
        RECT 397.645 18.110 397.875 18.480 ;
        RECT 399.320 18.395 399.550 19.400 ;
        RECT 400.430 19.420 400.770 20.240 ;
        RECT 401.000 19.880 401.230 20.480 ;
        RECT 401.830 20.110 402.635 20.450 ;
        RECT 401.000 19.650 402.000 19.880 ;
        RECT 400.430 19.190 401.320 19.420 ;
        RECT 399.320 18.165 399.960 18.395 ;
        RECT 401.090 18.080 401.320 19.190 ;
        RECT 401.770 18.715 402.000 19.650 ;
        RECT 402.295 18.310 402.635 20.110 ;
        RECT 403.540 20.220 405.175 20.580 ;
        RECT 403.540 19.410 404.085 20.220 ;
        RECT 405.530 19.790 405.760 20.450 ;
        RECT 404.610 19.560 407.110 19.790 ;
        RECT 404.610 19.065 404.840 19.560 ;
        RECT 402.875 18.835 404.840 19.065 ;
        RECT 403.075 18.190 404.345 18.420 ;
        RECT 404.610 18.310 404.840 18.835 ;
        RECT 403.075 18.080 403.305 18.190 ;
        RECT 401.090 17.850 403.305 18.080 ;
        RECT 404.115 18.080 404.345 18.190 ;
        RECT 405.070 18.080 405.300 19.330 ;
        RECT 404.115 17.850 405.300 18.080 ;
        RECT 407.355 17.860 407.790 20.690 ;
        RECT 408.165 19.685 409.440 19.915 ;
        RECT 408.165 17.850 408.395 19.685 ;
        RECT 409.685 19.280 409.915 20.710 ;
        RECT 408.650 19.050 409.915 19.280 ;
        RECT 410.405 19.685 411.680 19.915 ;
        RECT 410.405 17.850 410.635 19.685 ;
        RECT 411.925 19.280 412.155 20.710 ;
        RECT 415.870 19.450 416.175 20.640 ;
        RECT 410.890 19.050 412.155 19.280 ;
        RECT 415.145 19.110 416.175 19.450 ;
        RECT 416.405 18.880 416.760 20.640 ;
        RECT 415.335 18.560 416.760 18.880 ;
        RECT 415.335 17.860 415.615 18.560 ;
        RECT 416.990 17.920 417.295 20.060 ;
        RECT 418.245 19.685 419.520 19.915 ;
        RECT 418.245 17.850 418.475 19.685 ;
        RECT 419.765 19.280 419.995 20.710 ;
        RECT 418.730 19.050 419.995 19.280 ;
        RECT 420.485 19.685 421.760 19.915 ;
        RECT 420.485 17.850 420.715 19.685 ;
        RECT 422.005 19.280 422.235 20.710 ;
        RECT 420.970 19.050 422.235 19.280 ;
        RECT 422.725 19.685 424.000 19.915 ;
        RECT 422.725 17.850 422.955 19.685 ;
        RECT 424.245 19.280 424.475 20.710 ;
        RECT 423.210 19.050 424.475 19.280 ;
        RECT 425.985 17.920 426.290 20.060 ;
        RECT 426.520 18.880 426.875 20.640 ;
        RECT 427.105 19.450 427.410 20.640 ;
        RECT 429.550 20.200 430.315 20.630 ;
        RECT 427.105 19.110 428.135 19.450 ;
        RECT 429.550 18.950 429.880 20.200 ;
        RECT 431.975 19.960 432.370 20.710 ;
        RECT 434.920 20.370 436.260 20.690 ;
        RECT 430.145 19.730 432.370 19.960 ;
        RECT 430.145 19.600 431.000 19.730 ;
        RECT 426.520 18.850 427.945 18.880 ;
        RECT 426.520 18.590 427.990 18.850 ;
        RECT 426.520 18.560 427.945 18.590 ;
        RECT 427.665 17.860 427.945 18.560 ;
        RECT 429.550 17.895 430.180 18.950 ;
        RECT 431.540 17.895 431.900 19.500 ;
        RECT 432.140 18.110 432.370 19.730 ;
        RECT 432.600 18.360 433.020 20.165 ;
        RECT 434.340 19.470 434.690 20.080 ;
        RECT 433.795 19.090 434.690 19.470 ;
        RECT 432.140 17.880 433.345 18.110 ;
        RECT 433.870 18.080 434.210 18.745 ;
        RECT 434.920 18.515 435.225 20.370 ;
        RECT 439.525 20.225 439.755 20.565 ;
        RECT 441.765 20.225 441.995 20.565 ;
        RECT 436.020 19.470 436.360 20.080 ;
        RECT 437.155 19.470 437.495 20.080 ;
        RECT 439.525 19.990 442.475 20.225 ;
        RECT 442.140 19.555 442.475 19.990 ;
        RECT 454.085 19.685 455.360 19.915 ;
        RECT 435.455 19.090 436.360 19.470 ;
        RECT 436.590 19.090 437.495 19.470 ;
        RECT 438.810 19.090 441.670 19.525 ;
        RECT 442.140 19.215 446.430 19.555 ;
        RECT 435.910 18.080 436.250 18.745 ;
        RECT 442.140 18.710 442.475 19.215 ;
        RECT 448.500 19.210 451.700 19.555 ;
        RECT 433.870 17.850 436.250 18.080 ;
        RECT 439.425 18.480 442.475 18.710 ;
        RECT 439.425 17.860 439.655 18.480 ;
        RECT 441.665 17.860 441.895 18.480 ;
        RECT 454.085 17.850 454.315 19.685 ;
        RECT 455.605 19.280 455.835 20.710 ;
        RECT 458.225 19.960 458.455 20.440 ;
        RECT 454.570 19.050 455.835 19.280 ;
        RECT 457.310 19.730 458.455 19.960 ;
        RECT 457.310 18.880 457.650 19.730 ;
        RECT 460.040 19.500 460.415 20.690 ;
        RECT 457.910 19.200 459.230 19.500 ;
        RECT 457.310 18.530 458.455 18.880 ;
        RECT 458.225 17.850 458.455 18.530 ;
        RECT 458.905 18.650 459.230 19.200 ;
        RECT 459.470 19.090 460.415 19.500 ;
        RECT 460.645 18.650 460.875 20.435 ;
        RECT 458.905 18.420 460.875 18.650 ;
        RECT 460.645 17.850 460.875 18.420 ;
        RECT 298.905 16.110 299.135 16.780 ;
        RECT 301.145 16.110 301.375 16.780 ;
        RECT 303.385 16.110 303.615 16.780 ;
        RECT 305.525 16.110 305.755 16.780 ;
        RECT 307.865 16.160 308.095 16.780 ;
        RECT 310.105 16.160 310.335 16.780 ;
        RECT 298.870 15.730 305.755 16.110 ;
        RECT 307.285 15.930 310.335 16.160 ;
        RECT 298.060 15.085 301.260 15.430 ;
        RECT 301.960 14.820 302.760 15.730 ;
        RECT 307.285 15.425 307.620 15.930 ;
        RECT 303.330 15.085 307.620 15.425 ;
        RECT 308.090 15.115 310.950 15.550 ;
        RECT 298.805 14.440 305.755 14.820 ;
        RECT 298.805 14.075 299.035 14.440 ;
        RECT 301.045 14.075 301.275 14.440 ;
        RECT 303.285 14.075 303.515 14.440 ;
        RECT 305.495 14.075 305.755 14.440 ;
        RECT 307.285 14.650 307.620 15.085 ;
        RECT 307.285 14.415 310.235 14.650 ;
        RECT 307.765 14.075 307.995 14.415 ;
        RECT 310.005 14.075 310.235 14.415 ;
        RECT 312.860 14.210 313.195 16.110 ;
        RECT 316.885 14.955 317.115 16.790 ;
        RECT 317.370 15.360 318.635 15.590 ;
        RECT 316.885 14.725 318.160 14.955 ;
        RECT 318.405 13.930 318.635 15.360 ;
        RECT 320.145 14.580 320.450 16.720 ;
        RECT 321.825 16.080 322.105 16.780 ;
        RECT 320.680 15.760 322.105 16.080 ;
        RECT 325.175 16.080 325.455 16.780 ;
        RECT 326.310 16.080 326.570 16.110 ;
        RECT 325.175 15.760 326.600 16.080 ;
        RECT 320.680 14.000 321.035 15.760 ;
        RECT 321.265 15.190 322.295 15.530 ;
        RECT 324.985 15.190 326.015 15.530 ;
        RECT 321.265 14.000 321.570 15.190 ;
        RECT 325.710 14.000 326.015 15.190 ;
        RECT 326.245 14.000 326.600 15.760 ;
        RECT 326.830 14.580 327.135 16.720 ;
        RECT 328.085 14.955 328.315 16.790 ;
        RECT 328.570 15.360 329.835 15.590 ;
        RECT 328.085 14.725 329.360 14.955 ;
        RECT 329.605 13.930 329.835 15.360 ;
        RECT 330.325 14.955 330.555 16.790 ;
        RECT 330.810 15.360 332.075 15.590 ;
        RECT 330.325 14.725 331.600 14.955 ;
        RECT 331.845 13.930 332.075 15.360 ;
        RECT 332.565 14.955 332.795 16.790 ;
        RECT 333.050 15.360 334.315 15.590 ;
        RECT 332.565 14.725 333.840 14.955 ;
        RECT 334.085 13.930 334.315 15.360 ;
        RECT 334.805 14.955 335.035 16.790 ;
        RECT 335.290 15.360 336.555 15.590 ;
        RECT 334.805 14.725 336.080 14.955 ;
        RECT 336.325 13.930 336.555 15.360 ;
        RECT 337.045 14.955 337.275 16.790 ;
        RECT 337.530 15.360 338.795 15.590 ;
        RECT 337.045 14.725 338.320 14.955 ;
        RECT 338.565 13.930 338.795 15.360 ;
        RECT 339.285 14.955 339.515 16.790 ;
        RECT 341.470 16.560 343.850 16.790 ;
        RECT 341.470 15.895 341.810 16.560 ;
        RECT 339.770 15.360 341.035 15.590 ;
        RECT 339.285 14.725 340.560 14.955 ;
        RECT 340.805 13.930 341.035 15.360 ;
        RECT 341.395 15.170 342.290 15.550 ;
        RECT 341.940 14.560 342.290 15.170 ;
        RECT 342.520 14.270 342.825 16.125 ;
        RECT 343.510 15.895 343.850 16.560 ;
        RECT 343.055 15.170 343.960 15.550 ;
        RECT 344.190 15.170 345.095 15.550 ;
        RECT 343.620 14.560 343.960 15.170 ;
        RECT 344.755 14.560 345.095 15.170 ;
        RECT 346.005 14.955 346.235 16.790 ;
        RECT 346.490 15.360 347.755 15.590 ;
        RECT 346.005 14.725 347.280 14.955 ;
        RECT 343.110 14.270 343.370 14.430 ;
        RECT 342.520 13.950 343.860 14.270 ;
        RECT 347.525 13.930 347.755 15.360 ;
        RECT 348.245 14.955 348.475 16.790 ;
        RECT 348.730 15.360 349.995 15.590 ;
        RECT 348.245 14.725 349.520 14.955 ;
        RECT 349.765 13.930 349.995 15.360 ;
        RECT 350.485 14.955 350.715 16.790 ;
        RECT 350.970 15.360 352.235 15.590 ;
        RECT 350.485 14.725 351.760 14.955 ;
        RECT 352.005 13.930 352.235 15.360 ;
        RECT 352.725 14.955 352.955 16.790 ;
        RECT 353.210 15.360 354.475 15.590 ;
        RECT 352.725 14.725 354.000 14.955 ;
        RECT 354.245 13.930 354.475 15.360 ;
        RECT 356.085 14.955 356.315 16.790 ;
        RECT 356.570 15.360 357.835 15.590 ;
        RECT 356.085 14.725 357.360 14.955 ;
        RECT 357.605 13.930 357.835 15.360 ;
        RECT 358.325 14.955 358.555 16.790 ;
        RECT 358.810 15.360 360.075 15.590 ;
        RECT 358.325 14.725 359.600 14.955 ;
        RECT 359.845 13.930 360.075 15.360 ;
        RECT 360.565 14.955 360.795 16.790 ;
        RECT 363.465 16.035 363.695 16.625 ;
        RECT 363.465 15.805 365.155 16.035 ;
        RECT 361.050 15.360 362.315 15.590 ;
        RECT 360.565 14.725 361.840 14.955 ;
        RECT 362.085 13.930 362.315 15.360 ;
        RECT 363.270 15.170 364.690 15.550 ;
        RECT 364.925 14.910 365.155 15.805 ;
        RECT 363.365 14.680 365.155 14.910 ;
        RECT 365.385 16.015 365.735 16.615 ;
        RECT 366.785 16.390 368.035 16.620 ;
        RECT 375.330 16.560 377.545 16.790 ;
        RECT 366.785 16.015 367.015 16.390 ;
        RECT 365.385 15.785 367.015 16.015 ;
        RECT 367.245 15.820 367.575 16.160 ;
        RECT 363.365 14.210 363.595 14.680 ;
        RECT 365.385 14.495 365.615 15.785 ;
        RECT 366.010 15.170 367.040 15.550 ;
        RECT 365.385 14.265 365.890 14.495 ;
        RECT 367.345 14.475 367.575 15.820 ;
        RECT 367.805 15.310 368.035 16.390 ;
        RECT 369.285 16.160 369.515 16.355 ;
        RECT 371.885 16.160 372.115 16.530 ;
        RECT 368.265 15.700 368.495 16.160 ;
        RECT 369.285 15.930 372.115 16.160 ;
        RECT 373.560 16.245 374.200 16.475 ;
        RECT 372.975 15.700 373.275 15.925 ;
        RECT 368.265 15.470 373.275 15.700 ;
        RECT 367.345 14.245 367.750 14.475 ;
        RECT 368.585 14.190 368.815 15.470 ;
        RECT 373.560 15.240 373.790 16.245 ;
        RECT 375.330 15.450 375.560 16.560 ;
        RECT 377.315 16.450 377.545 16.560 ;
        RECT 378.355 16.560 379.540 16.790 ;
        RECT 378.355 16.450 378.585 16.560 ;
        RECT 369.810 15.010 373.790 15.240 ;
        RECT 374.670 15.220 375.560 15.450 ;
        RECT 369.165 14.780 369.395 14.990 ;
        RECT 369.165 14.550 372.350 14.780 ;
        RECT 372.120 14.160 372.350 14.550 ;
        RECT 373.110 14.400 373.450 15.010 ;
        RECT 374.045 14.160 374.275 14.990 ;
        RECT 374.670 14.400 375.010 15.220 ;
        RECT 376.010 14.990 376.240 15.925 ;
        RECT 375.240 14.760 376.240 14.990 ;
        RECT 375.240 14.160 375.470 14.760 ;
        RECT 376.535 14.530 376.875 16.330 ;
        RECT 377.315 16.220 378.585 16.450 ;
        RECT 378.850 15.805 379.080 16.330 ;
        RECT 377.115 15.575 379.080 15.805 ;
        RECT 376.070 14.190 376.875 14.530 ;
        RECT 377.780 14.420 378.325 15.230 ;
        RECT 378.850 15.080 379.080 15.575 ;
        RECT 379.310 15.310 379.540 16.560 ;
        RECT 378.850 14.850 381.350 15.080 ;
        RECT 377.780 14.370 379.415 14.420 ;
        RECT 372.120 13.930 375.470 14.160 ;
        RECT 377.770 14.110 379.415 14.370 ;
        RECT 379.770 14.190 380.000 14.850 ;
        RECT 377.780 14.060 379.415 14.110 ;
        RECT 381.595 13.950 382.030 16.780 ;
        RECT 382.405 14.955 382.635 16.790 ;
        RECT 382.890 15.360 384.155 15.590 ;
        RECT 382.405 14.725 383.680 14.955 ;
        RECT 383.925 13.930 384.155 15.360 ;
        RECT 384.645 14.955 384.875 16.790 ;
        RECT 385.130 15.360 386.395 15.590 ;
        RECT 384.645 14.725 385.920 14.955 ;
        RECT 386.165 13.930 386.395 15.360 ;
        RECT 386.885 14.955 387.115 16.790 ;
        RECT 387.370 15.360 388.635 15.590 ;
        RECT 386.885 14.725 388.160 14.955 ;
        RECT 388.405 13.930 388.635 15.360 ;
        RECT 389.125 14.955 389.355 16.790 ;
        RECT 395.285 16.215 395.670 16.790 ;
        RECT 389.610 15.360 390.875 15.590 ;
        RECT 389.125 14.725 390.400 14.955 ;
        RECT 390.645 13.930 390.875 15.360 ;
        RECT 391.260 14.210 391.595 16.110 ;
        RECT 395.285 15.980 397.295 16.215 ;
        RECT 391.270 14.050 391.530 14.210 ;
        RECT 395.285 14.200 395.515 15.980 ;
        RECT 395.745 15.030 396.630 15.590 ;
        RECT 397.010 15.230 397.295 15.980 ;
        RECT 395.745 14.050 396.260 15.030 ;
        RECT 397.525 15.000 397.995 16.780 ;
        RECT 398.655 16.160 398.995 16.780 ;
        RECT 400.220 16.545 403.075 16.780 ;
        RECT 400.220 16.160 400.450 16.545 ;
        RECT 398.655 15.930 400.450 16.160 ;
        RECT 400.750 15.780 402.290 16.110 ;
        RECT 402.735 15.930 403.075 16.545 ;
        RECT 404.345 16.035 404.575 16.625 ;
        RECT 404.345 15.805 406.035 16.035 ;
        RECT 397.370 13.975 397.995 15.000 ;
        RECT 399.010 15.170 399.970 15.550 ;
        RECT 399.010 14.485 399.405 15.170 ;
        RECT 400.200 13.950 400.520 15.550 ;
        RECT 400.750 13.985 401.080 15.780 ;
        RECT 401.320 13.950 401.640 15.550 ;
        RECT 401.880 15.200 402.945 15.550 ;
        RECT 401.880 13.950 402.200 15.200 ;
        RECT 404.150 15.170 405.570 15.550 ;
        RECT 405.805 14.910 406.035 15.805 ;
        RECT 404.245 14.680 406.035 14.910 ;
        RECT 406.265 16.015 406.615 16.615 ;
        RECT 407.665 16.390 408.915 16.620 ;
        RECT 416.210 16.560 418.425 16.790 ;
        RECT 407.665 16.015 407.895 16.390 ;
        RECT 406.265 15.785 407.895 16.015 ;
        RECT 408.125 15.820 408.455 16.160 ;
        RECT 404.245 14.210 404.475 14.680 ;
        RECT 406.265 14.495 406.495 15.785 ;
        RECT 406.890 15.170 407.920 15.550 ;
        RECT 406.265 14.265 406.770 14.495 ;
        RECT 408.225 14.475 408.455 15.820 ;
        RECT 408.685 15.310 408.915 16.390 ;
        RECT 410.165 16.160 410.395 16.355 ;
        RECT 412.765 16.160 412.995 16.530 ;
        RECT 409.145 15.700 409.375 16.160 ;
        RECT 410.165 15.930 412.995 16.160 ;
        RECT 414.440 16.245 415.080 16.475 ;
        RECT 413.855 15.700 414.155 15.925 ;
        RECT 409.145 15.470 414.155 15.700 ;
        RECT 408.225 14.245 408.630 14.475 ;
        RECT 409.465 14.190 409.695 15.470 ;
        RECT 414.440 15.240 414.670 16.245 ;
        RECT 416.210 15.450 416.440 16.560 ;
        RECT 418.195 16.450 418.425 16.560 ;
        RECT 419.235 16.560 420.420 16.790 ;
        RECT 419.235 16.450 419.465 16.560 ;
        RECT 410.690 15.010 414.670 15.240 ;
        RECT 415.550 15.220 416.440 15.450 ;
        RECT 410.045 14.780 410.275 14.990 ;
        RECT 410.045 14.550 413.230 14.780 ;
        RECT 413.000 14.160 413.230 14.550 ;
        RECT 413.990 14.400 414.330 15.010 ;
        RECT 414.925 14.160 415.155 14.990 ;
        RECT 415.550 14.400 415.890 15.220 ;
        RECT 416.890 14.990 417.120 15.925 ;
        RECT 416.120 14.760 417.120 14.990 ;
        RECT 416.120 14.160 416.350 14.760 ;
        RECT 417.415 14.530 417.755 16.330 ;
        RECT 418.195 16.220 419.465 16.450 ;
        RECT 419.730 15.805 419.960 16.330 ;
        RECT 417.995 15.575 419.960 15.805 ;
        RECT 416.950 14.190 417.755 14.530 ;
        RECT 418.660 14.420 419.205 15.230 ;
        RECT 419.730 15.080 419.960 15.575 ;
        RECT 420.190 15.310 420.420 16.560 ;
        RECT 419.730 14.850 422.230 15.080 ;
        RECT 413.000 13.930 416.350 14.160 ;
        RECT 418.660 14.060 420.295 14.420 ;
        RECT 420.650 14.190 420.880 14.850 ;
        RECT 422.475 13.950 422.910 16.780 ;
        RECT 424.625 16.110 424.855 16.790 ;
        RECT 427.045 16.220 427.275 16.790 ;
        RECT 423.710 15.760 424.855 16.110 ;
        RECT 425.305 15.990 427.275 16.220 ;
        RECT 423.710 14.910 424.050 15.760 ;
        RECT 425.305 15.440 425.630 15.990 ;
        RECT 424.310 15.140 425.630 15.440 ;
        RECT 425.870 15.140 426.815 15.550 ;
        RECT 423.710 14.680 424.855 14.910 ;
        RECT 424.625 14.200 424.855 14.680 ;
        RECT 426.440 13.950 426.815 15.140 ;
        RECT 427.045 14.205 427.275 15.990 ;
        RECT 427.765 16.215 428.150 16.790 ;
        RECT 427.765 15.980 429.775 16.215 ;
        RECT 427.765 14.200 427.995 15.980 ;
        RECT 428.225 15.030 429.110 15.590 ;
        RECT 429.490 15.230 429.775 15.980 ;
        RECT 428.225 14.050 428.740 15.030 ;
        RECT 430.005 15.000 430.475 16.780 ;
        RECT 429.850 13.975 430.475 15.000 ;
        RECT 431.125 14.955 431.355 16.790 ;
        RECT 434.430 16.560 436.810 16.790 ;
        RECT 434.430 15.895 434.770 16.560 ;
        RECT 431.610 15.360 432.875 15.590 ;
        RECT 431.125 14.725 432.400 14.955 ;
        RECT 432.645 13.930 432.875 15.360 ;
        RECT 434.355 15.170 435.250 15.550 ;
        RECT 434.900 14.560 435.250 15.170 ;
        RECT 435.480 14.270 435.785 16.125 ;
        RECT 436.470 15.895 436.810 16.560 ;
        RECT 436.015 15.170 436.920 15.550 ;
        RECT 437.150 15.170 438.055 15.550 ;
        RECT 436.580 14.560 436.920 15.170 ;
        RECT 437.715 14.560 438.055 15.170 ;
        RECT 438.965 14.955 439.195 16.790 ;
        RECT 439.450 15.360 440.715 15.590 ;
        RECT 438.965 14.725 440.240 14.955 ;
        RECT 435.480 13.950 436.820 14.270 ;
        RECT 440.485 13.930 440.715 15.360 ;
        RECT 442.210 13.950 442.645 16.780 ;
        RECT 444.700 16.560 445.885 16.790 ;
        RECT 444.700 15.310 444.930 16.560 ;
        RECT 445.655 16.450 445.885 16.560 ;
        RECT 446.695 16.560 448.910 16.790 ;
        RECT 446.695 16.450 446.925 16.560 ;
        RECT 445.160 15.805 445.390 16.330 ;
        RECT 445.655 16.220 446.925 16.450 ;
        RECT 445.160 15.575 447.125 15.805 ;
        RECT 445.160 15.080 445.390 15.575 ;
        RECT 442.890 14.850 445.390 15.080 ;
        RECT 444.240 14.190 444.470 14.850 ;
        RECT 445.915 14.420 446.460 15.230 ;
        RECT 444.825 14.370 446.460 14.420 ;
        RECT 447.365 14.530 447.705 16.330 ;
        RECT 448.000 14.990 448.230 15.925 ;
        RECT 448.680 15.450 448.910 16.560 ;
        RECT 450.040 16.245 450.680 16.475 ;
        RECT 448.680 15.220 449.570 15.450 ;
        RECT 448.000 14.760 449.000 14.990 ;
        RECT 444.825 14.110 446.470 14.370 ;
        RECT 447.365 14.190 448.170 14.530 ;
        RECT 448.770 14.160 449.000 14.760 ;
        RECT 449.230 14.400 449.570 15.220 ;
        RECT 450.450 15.240 450.680 16.245 ;
        RECT 452.125 16.160 452.355 16.530 ;
        RECT 456.205 16.390 457.455 16.620 ;
        RECT 454.725 16.160 454.955 16.355 ;
        RECT 452.125 15.930 454.955 16.160 ;
        RECT 450.965 15.700 451.265 15.925 ;
        RECT 455.745 15.700 455.975 16.160 ;
        RECT 450.965 15.470 455.975 15.700 ;
        RECT 450.450 15.010 454.430 15.240 ;
        RECT 449.965 14.160 450.195 14.990 ;
        RECT 450.790 14.400 451.130 15.010 ;
        RECT 454.845 14.780 455.075 14.990 ;
        RECT 451.890 14.550 455.075 14.780 ;
        RECT 451.890 14.160 452.120 14.550 ;
        RECT 455.425 14.190 455.655 15.470 ;
        RECT 456.205 15.310 456.435 16.390 ;
        RECT 456.665 15.820 456.995 16.160 ;
        RECT 457.225 16.015 457.455 16.390 ;
        RECT 458.505 16.015 458.855 16.615 ;
        RECT 460.545 16.035 460.775 16.625 ;
        RECT 456.665 14.475 456.895 15.820 ;
        RECT 457.225 15.785 458.855 16.015 ;
        RECT 457.200 15.170 458.230 15.550 ;
        RECT 458.625 14.495 458.855 15.785 ;
        RECT 459.085 15.805 460.775 16.035 ;
        RECT 459.085 14.910 459.315 15.805 ;
        RECT 459.550 15.170 460.840 15.550 ;
        RECT 459.085 14.680 460.875 14.910 ;
        RECT 456.490 14.245 456.895 14.475 ;
        RECT 458.350 14.265 458.855 14.495 ;
        RECT 460.645 14.210 460.875 14.680 ;
        RECT 444.825 14.060 446.460 14.110 ;
        RECT 448.770 13.930 452.120 14.160 ;
        RECT 223.900 11.955 232.945 12.355 ;
        RECT 183.905 10.305 184.805 10.685 ;
        RECT 184.205 8.150 184.505 10.305 ;
        RECT 171.420 7.850 184.505 8.150 ;
        RECT 171.420 6.785 172.290 7.850 ;
        RECT 172.520 6.300 172.750 6.670 ;
        RECT 172.520 6.290 181.855 6.300 ;
        RECT 172.520 5.910 182.305 6.290 ;
        RECT 172.520 5.900 181.855 5.910 ;
        RECT 172.520 5.530 172.750 5.900 ;
        RECT 171.420 5.185 172.290 5.415 ;
        RECT 171.655 3.190 172.055 5.185 ;
        RECT 179.705 4.950 180.005 5.000 ;
        RECT 179.665 4.050 180.045 4.950 ;
        RECT 171.405 2.810 172.305 3.190 ;
        RECT 175.905 2.810 177.855 3.190 ;
        RECT 171.655 0.915 172.055 2.810 ;
        RECT 173.200 1.350 174.100 1.390 ;
        RECT 172.520 1.050 174.100 1.350 ;
        RECT 171.420 0.685 172.290 0.915 ;
        RECT 172.520 0.230 172.750 1.050 ;
        RECT 173.200 1.010 174.100 1.050 ;
        RECT 174.855 1.010 176.805 1.390 ;
        RECT 171.420 -0.915 172.290 -0.685 ;
        RECT 171.655 -2.810 172.055 -0.915 ;
        RECT 172.520 -1.050 172.750 -0.230 ;
        RECT 173.200 -1.050 174.100 -1.010 ;
        RECT 172.520 -1.350 174.100 -1.050 ;
        RECT 173.200 -1.390 174.100 -1.350 ;
        RECT 174.855 -2.810 175.155 1.010 ;
        RECT 177.555 -1.010 177.855 2.810 ;
        RECT 179.705 0.515 180.005 4.050 ;
        RECT 181.905 2.810 182.805 3.190 ;
        RECT 181.920 1.485 182.790 2.810 ;
        RECT 180.625 1.370 181.525 1.390 ;
        RECT 180.625 1.030 181.690 1.370 ;
        RECT 180.625 1.010 181.525 1.030 ;
        RECT 184.205 0.915 184.505 7.850 ;
        RECT 185.405 6.255 186.305 6.295 ;
        RECT 185.405 5.955 187.620 6.255 ;
        RECT 185.405 5.915 186.305 5.955 ;
        RECT 181.920 0.685 184.505 0.915 ;
        RECT 187.320 0.570 187.620 5.955 ;
        RECT 223.900 3.300 224.270 11.955 ;
        RECT 232.545 10.340 232.945 11.955 ;
        RECT 297.285 11.845 298.560 12.075 ;
        RECT 235.860 10.685 236.090 11.170 ;
        RECT 234.290 10.620 236.090 10.685 ;
        RECT 234.290 10.455 236.240 10.620 ;
        RECT 231.390 10.000 234.060 10.340 ;
        RECT 230.260 9.505 231.160 9.885 ;
        RECT 234.290 9.505 235.190 9.885 ;
        RECT 235.860 9.720 236.240 10.455 ;
        RECT 297.285 10.010 297.515 11.845 ;
        RECT 298.805 11.440 299.035 12.870 ;
        RECT 297.770 11.210 299.035 11.440 ;
        RECT 299.525 11.845 300.800 12.075 ;
        RECT 299.525 10.010 299.755 11.845 ;
        RECT 301.045 11.440 301.275 12.870 ;
        RECT 300.010 11.210 301.275 11.440 ;
        RECT 301.765 11.845 303.040 12.075 ;
        RECT 301.765 10.010 301.995 11.845 ;
        RECT 303.285 11.440 303.515 12.870 ;
        RECT 302.250 11.210 303.515 11.440 ;
        RECT 306.085 10.690 306.420 12.590 ;
        RECT 306.805 12.345 307.035 12.595 ;
        RECT 306.805 12.110 309.735 12.345 ;
        RECT 307.220 10.590 307.580 11.860 ;
        RECT 307.825 10.075 308.055 12.110 ;
        RECT 308.340 10.030 308.700 11.860 ;
        RECT 309.505 11.415 309.735 12.110 ;
        RECT 310.010 10.020 310.430 12.845 ;
        RECT 312.345 12.410 312.690 12.870 ;
        RECT 314.770 12.410 315.110 12.870 ;
        RECT 317.530 12.410 317.870 12.870 ;
        RECT 320.780 12.640 323.900 12.870 ;
        RECT 311.385 12.180 314.535 12.410 ;
        RECT 311.385 10.205 311.615 12.180 ;
        RECT 314.770 12.175 317.150 12.410 ;
        RECT 317.530 12.175 320.580 12.410 ;
        RECT 312.810 11.575 313.265 11.945 ;
        RECT 314.710 11.710 315.810 11.945 ;
        RECT 314.710 11.575 314.940 11.710 ;
        RECT 312.810 11.305 314.940 11.575 ;
        RECT 316.215 11.480 316.660 11.805 ;
        RECT 315.170 11.250 316.660 11.480 ;
        RECT 315.170 11.015 315.400 11.250 ;
        RECT 316.920 11.020 317.150 12.175 ;
        RECT 318.070 11.020 318.300 11.865 ;
        RECT 311.910 10.745 315.400 11.015 ;
        RECT 315.780 10.790 318.300 11.020 ;
        RECT 314.760 10.240 315.120 10.500 ;
        RECT 315.780 10.470 316.140 10.790 ;
        RECT 316.800 10.240 317.160 10.500 ;
        RECT 314.760 10.010 317.160 10.240 ;
        RECT 318.070 10.240 318.300 10.790 ;
        RECT 318.550 10.470 318.890 12.175 ;
        RECT 320.240 11.835 320.580 12.175 ;
        RECT 322.210 11.820 323.800 12.410 ;
        RECT 319.125 11.305 321.805 11.575 ;
        RECT 322.260 11.305 323.210 11.540 ;
        RECT 322.260 11.070 322.490 11.305 ;
        RECT 319.310 10.835 322.490 11.070 ;
        RECT 323.480 11.040 323.800 11.820 ;
        RECT 319.310 10.240 319.540 10.835 ;
        RECT 322.920 10.720 323.800 11.040 ;
        RECT 324.725 10.940 324.955 12.850 ;
        RECT 325.185 11.170 325.480 12.850 ;
        RECT 322.920 10.480 323.255 10.720 ;
        RECT 324.725 10.710 325.465 10.940 ;
        RECT 318.070 10.010 319.540 10.240 ;
        RECT 320.610 10.160 323.255 10.480 ;
        RECT 325.235 10.240 325.465 10.710 ;
        RECT 325.710 10.810 326.075 12.850 ;
        RECT 326.305 11.080 326.640 12.850 ;
        RECT 326.965 11.270 327.195 12.850 ;
        RECT 327.425 11.800 327.760 12.850 ;
        RECT 329.205 11.845 330.480 12.075 ;
        RECT 327.425 11.500 328.830 11.800 ;
        RECT 326.965 11.040 327.555 11.270 ;
        RECT 327.855 11.250 328.830 11.500 ;
        RECT 325.710 10.470 327.095 10.810 ;
        RECT 327.325 10.240 327.555 11.040 ;
        RECT 325.235 10.010 327.555 10.240 ;
        RECT 329.205 10.010 329.435 11.845 ;
        RECT 330.725 11.440 330.955 12.870 ;
        RECT 329.690 11.210 330.955 11.440 ;
        RECT 331.445 11.845 332.720 12.075 ;
        RECT 331.445 10.010 331.675 11.845 ;
        RECT 332.965 11.440 333.195 12.870 ;
        RECT 331.930 11.210 333.195 11.440 ;
        RECT 336.485 11.845 337.760 12.075 ;
        RECT 336.485 10.010 336.715 11.845 ;
        RECT 338.005 11.440 338.235 12.870 ;
        RECT 336.970 11.210 338.235 11.440 ;
        RECT 338.725 11.845 340.000 12.075 ;
        RECT 338.725 10.010 338.955 11.845 ;
        RECT 340.245 11.440 340.475 12.870 ;
        RECT 339.210 11.210 340.475 11.440 ;
        RECT 341.065 12.240 341.580 12.850 ;
        RECT 344.770 12.640 348.950 12.870 ;
        RECT 341.065 11.210 341.455 12.240 ;
        RECT 342.920 11.900 343.150 12.595 ;
        RECT 344.770 12.005 345.000 12.640 ;
        RECT 348.720 12.610 348.950 12.640 ;
        RECT 349.840 12.640 352.770 12.870 ;
        RECT 346.385 12.180 348.325 12.410 ;
        RECT 348.720 12.270 349.610 12.610 ;
        RECT 341.760 11.560 343.150 11.900 ;
        RECT 343.545 11.770 345.000 12.005 ;
        RECT 342.920 11.540 343.150 11.560 ;
        RECT 342.920 11.295 345.125 11.540 ;
        RECT 341.065 10.020 341.835 11.210 ;
        RECT 342.920 10.020 343.150 11.295 ;
        RECT 345.595 11.250 346.790 11.630 ;
        RECT 347.020 10.860 347.250 12.180 ;
        RECT 345.280 10.625 347.250 10.860 ;
        RECT 348.720 10.850 348.950 12.270 ;
        RECT 349.840 11.785 350.070 12.640 ;
        RECT 350.665 11.320 351.005 12.410 ;
        RECT 352.540 12.095 352.770 12.640 ;
        RECT 352.540 11.865 354.880 12.095 ;
        RECT 355.205 11.635 355.535 12.610 ;
        RECT 352.645 11.405 355.535 11.635 ;
        RECT 345.280 10.515 345.510 10.625 ;
        RECT 347.020 10.555 347.250 10.625 ;
        RECT 347.985 10.620 348.950 10.850 ;
        RECT 349.235 11.175 351.845 11.320 ;
        RECT 349.235 11.090 353.865 11.175 ;
        RECT 349.235 10.620 349.575 11.090 ;
        RECT 351.505 10.945 353.865 11.090 ;
        RECT 349.805 10.625 351.195 10.860 ;
        RECT 349.805 10.335 350.035 10.625 ;
        RECT 348.565 10.105 350.035 10.335 ;
        RECT 350.965 10.240 351.195 10.625 ;
        RECT 351.505 10.470 351.845 10.945 ;
        RECT 354.425 10.415 354.765 11.160 ;
        RECT 355.305 10.415 355.535 11.405 ;
        RECT 352.380 10.240 354.765 10.415 ;
        RECT 350.965 10.185 354.765 10.240 ;
        RECT 355.765 10.240 355.995 11.470 ;
        RECT 356.270 10.470 356.610 12.610 ;
        RECT 358.165 12.250 358.495 12.590 ;
        RECT 356.850 11.250 357.990 11.630 ;
        RECT 358.260 11.020 358.495 12.250 ;
        RECT 360.405 12.120 360.635 12.590 ;
        RECT 356.840 10.785 358.495 11.020 ;
        RECT 358.790 11.890 360.635 12.120 ;
        RECT 358.790 11.040 359.020 11.890 ;
        RECT 361.125 11.845 362.400 12.075 ;
        RECT 359.290 11.270 360.600 11.635 ;
        RECT 358.790 10.805 360.535 11.040 ;
        RECT 356.840 10.240 357.070 10.785 ;
        RECT 350.965 10.010 352.610 10.185 ;
        RECT 355.765 10.010 357.070 10.240 ;
        RECT 358.265 10.175 358.495 10.785 ;
        RECT 360.305 10.175 360.535 10.805 ;
        RECT 361.125 10.010 361.355 11.845 ;
        RECT 362.645 11.440 362.875 12.870 ;
        RECT 361.610 11.210 362.875 11.440 ;
        RECT 363.365 11.845 364.640 12.075 ;
        RECT 363.365 10.010 363.595 11.845 ;
        RECT 364.885 11.440 365.115 12.870 ;
        RECT 363.850 11.210 365.115 11.440 ;
        RECT 366.910 11.795 367.500 12.835 ;
        RECT 366.910 10.080 367.275 11.795 ;
        RECT 368.760 11.660 369.135 12.365 ;
        RECT 367.570 10.880 367.910 11.520 ;
        RECT 368.250 11.250 369.135 11.660 ;
        RECT 369.365 10.880 369.595 12.835 ;
        RECT 367.570 10.645 369.595 10.880 ;
        RECT 369.265 10.020 369.595 10.645 ;
        RECT 370.270 11.795 370.860 12.835 ;
        RECT 370.270 10.080 370.635 11.795 ;
        RECT 372.120 11.660 372.495 12.365 ;
        RECT 370.930 10.880 371.270 11.520 ;
        RECT 371.610 11.250 372.495 11.660 ;
        RECT 372.725 10.880 372.955 12.835 ;
        RECT 370.930 10.645 372.955 10.880 ;
        RECT 372.625 10.020 372.955 10.645 ;
        RECT 375.685 11.845 376.960 12.075 ;
        RECT 375.685 10.010 375.915 11.845 ;
        RECT 377.205 11.440 377.435 12.870 ;
        RECT 376.170 11.210 377.435 11.440 ;
        RECT 377.925 11.845 379.200 12.075 ;
        RECT 377.925 10.010 378.155 11.845 ;
        RECT 379.445 11.440 379.675 12.870 ;
        RECT 378.410 11.210 379.675 11.440 ;
        RECT 380.165 11.845 381.440 12.075 ;
        RECT 380.165 10.010 380.395 11.845 ;
        RECT 381.685 11.440 381.915 12.870 ;
        RECT 384.865 12.120 385.095 12.600 ;
        RECT 380.650 11.210 381.915 11.440 ;
        RECT 383.950 11.890 385.095 12.120 ;
        RECT 383.950 11.040 384.290 11.890 ;
        RECT 386.680 11.660 387.055 12.850 ;
        RECT 384.550 11.360 385.870 11.660 ;
        RECT 383.950 10.690 385.095 11.040 ;
        RECT 384.865 10.010 385.095 10.690 ;
        RECT 385.545 10.810 385.870 11.360 ;
        RECT 386.110 11.250 387.055 11.660 ;
        RECT 387.285 10.810 387.515 12.595 ;
        RECT 385.545 10.580 387.515 10.810 ;
        RECT 387.285 10.010 387.515 10.580 ;
        RECT 388.190 11.795 388.780 12.835 ;
        RECT 388.190 10.080 388.555 11.795 ;
        RECT 390.040 11.660 390.415 12.365 ;
        RECT 388.850 10.880 389.190 11.520 ;
        RECT 389.530 11.250 390.415 11.660 ;
        RECT 390.645 10.880 390.875 12.835 ;
        RECT 392.485 12.750 392.715 12.870 ;
        RECT 392.390 12.370 392.715 12.750 ;
        RECT 392.485 12.350 392.715 12.370 ;
        RECT 394.725 12.350 394.955 12.870 ;
        RECT 392.485 12.080 396.015 12.350 ;
        RECT 391.930 11.630 392.180 11.820 ;
        RECT 391.830 11.250 392.180 11.630 ;
        RECT 392.600 11.250 394.340 11.630 ;
        RECT 394.600 11.250 395.510 11.630 ;
        RECT 388.850 10.645 390.875 10.880 ;
        RECT 391.930 11.020 392.180 11.250 ;
        RECT 394.600 11.020 394.900 11.250 ;
        RECT 391.930 10.700 394.900 11.020 ;
        RECT 390.545 10.020 390.875 10.645 ;
        RECT 395.745 10.600 396.015 12.080 ;
        RECT 395.215 10.365 396.015 10.600 ;
        RECT 396.965 11.845 398.240 12.075 ;
        RECT 395.215 10.260 395.445 10.365 ;
        RECT 393.510 10.030 395.445 10.260 ;
        RECT 396.965 10.010 397.195 11.845 ;
        RECT 398.485 11.440 398.715 12.870 ;
        RECT 397.450 11.210 398.715 11.440 ;
        RECT 399.205 11.845 400.480 12.075 ;
        RECT 399.205 10.010 399.435 11.845 ;
        RECT 400.725 11.440 400.955 12.870 ;
        RECT 399.690 11.210 400.955 11.440 ;
        RECT 403.585 10.450 403.910 12.430 ;
        RECT 404.140 10.030 404.475 12.800 ;
        RECT 405.550 11.795 406.140 12.835 ;
        RECT 405.550 10.080 405.915 11.795 ;
        RECT 407.400 11.660 407.775 12.365 ;
        RECT 406.210 10.880 406.550 11.520 ;
        RECT 406.890 11.250 407.775 11.660 ;
        RECT 408.005 10.880 408.235 12.835 ;
        RECT 406.210 10.645 408.235 10.880 ;
        RECT 409.740 10.690 410.075 12.590 ;
        RECT 410.965 11.845 412.240 12.075 ;
        RECT 407.905 10.020 408.235 10.645 ;
        RECT 410.965 10.010 411.195 11.845 ;
        RECT 412.485 11.440 412.715 12.870 ;
        RECT 411.450 11.210 412.715 11.440 ;
        RECT 414.885 11.845 416.160 12.075 ;
        RECT 414.885 10.010 415.115 11.845 ;
        RECT 416.405 11.440 416.635 12.870 ;
        RECT 415.370 11.210 416.635 11.440 ;
        RECT 417.125 11.845 418.400 12.075 ;
        RECT 417.125 10.010 417.355 11.845 ;
        RECT 418.645 11.440 418.875 12.870 ;
        RECT 417.610 11.210 418.875 11.440 ;
        RECT 419.365 11.845 420.640 12.075 ;
        RECT 419.365 10.010 419.595 11.845 ;
        RECT 420.885 11.440 421.115 12.870 ;
        RECT 419.850 11.210 421.115 11.440 ;
        RECT 421.605 11.845 422.880 12.075 ;
        RECT 421.605 10.010 421.835 11.845 ;
        RECT 423.125 11.440 423.355 12.870 ;
        RECT 422.090 11.210 423.355 11.440 ;
        RECT 423.845 11.845 425.120 12.075 ;
        RECT 423.845 10.010 424.075 11.845 ;
        RECT 425.365 11.440 425.595 12.870 ;
        RECT 426.550 12.590 426.810 12.750 ;
        RECT 424.330 11.210 425.595 11.440 ;
        RECT 426.540 10.690 426.875 12.590 ;
        RECT 427.765 11.845 429.040 12.075 ;
        RECT 427.765 10.010 427.995 11.845 ;
        RECT 429.285 11.440 429.515 12.870 ;
        RECT 428.250 11.210 429.515 11.440 ;
        RECT 430.005 11.845 431.280 12.075 ;
        RECT 430.005 10.010 430.235 11.845 ;
        RECT 431.525 11.440 431.755 12.870 ;
        RECT 432.710 12.590 432.970 12.750 ;
        RECT 430.490 11.210 431.755 11.440 ;
        RECT 432.700 10.690 433.035 12.590 ;
        RECT 434.340 10.520 434.760 12.325 ;
        RECT 434.990 12.120 435.385 12.870 ;
        RECT 437.045 12.360 437.810 12.790 ;
        RECT 434.990 11.890 437.215 12.120 ;
        RECT 434.990 10.270 435.220 11.890 ;
        RECT 436.360 11.760 437.215 11.890 ;
        RECT 434.015 10.040 435.220 10.270 ;
        RECT 435.460 10.055 435.820 11.660 ;
        RECT 437.480 11.110 437.810 12.360 ;
        RECT 439.525 12.385 439.755 12.725 ;
        RECT 441.765 12.385 441.995 12.725 ;
        RECT 439.525 12.150 442.475 12.385 ;
        RECT 442.140 11.715 442.475 12.150 ;
        RECT 454.085 11.845 455.360 12.075 ;
        RECT 438.810 11.250 441.670 11.685 ;
        RECT 442.140 11.375 446.430 11.715 ;
        RECT 437.180 10.055 437.810 11.110 ;
        RECT 442.140 10.870 442.475 11.375 ;
        RECT 448.500 11.370 451.700 11.715 ;
        RECT 439.425 10.640 442.475 10.870 ;
        RECT 439.425 10.020 439.655 10.640 ;
        RECT 441.665 10.020 441.895 10.640 ;
        RECT 454.085 10.010 454.315 11.845 ;
        RECT 455.605 11.440 455.835 12.870 ;
        RECT 454.570 11.210 455.835 11.440 ;
        RECT 456.325 11.845 457.600 12.075 ;
        RECT 456.325 10.010 456.555 11.845 ;
        RECT 457.845 11.440 458.075 12.870 ;
        RECT 456.810 11.210 458.075 11.440 ;
        RECT 458.565 11.845 459.840 12.075 ;
        RECT 458.565 10.010 458.795 11.845 ;
        RECT 460.085 11.440 460.315 12.870 ;
        RECT 459.050 11.210 460.315 11.440 ;
        RECT 232.295 9.105 233.195 9.505 ;
        RECT 235.860 9.170 236.090 9.720 ;
        RECT 230.290 8.275 231.160 8.505 ;
        RECT 232.545 8.160 232.945 9.105 ;
        RECT 231.390 7.820 232.945 8.160 ;
        RECT 297.285 8.315 297.615 8.940 ;
        RECT 297.285 8.080 299.310 8.315 ;
        RECT 230.290 7.475 231.160 7.705 ;
        RECT 230.525 7.050 230.925 7.475 ;
        RECT 230.525 6.730 232.945 7.050 ;
        RECT 232.545 5.980 232.945 6.730 ;
        RECT 235.860 6.325 236.090 6.810 ;
        RECT 234.290 6.260 236.090 6.325 ;
        RECT 234.290 6.095 236.240 6.260 ;
        RECT 297.285 6.125 297.515 8.080 ;
        RECT 297.745 7.300 298.630 7.710 ;
        RECT 298.970 7.440 299.310 8.080 ;
        RECT 297.745 6.595 298.120 7.300 ;
        RECT 299.605 7.165 299.970 8.880 ;
        RECT 299.380 6.125 299.970 7.165 ;
        RECT 301.765 8.315 302.095 8.940 ;
        RECT 301.765 8.080 303.790 8.315 ;
        RECT 301.765 6.125 301.995 8.080 ;
        RECT 302.225 7.300 303.110 7.710 ;
        RECT 303.450 7.440 303.790 8.080 ;
        RECT 302.225 6.595 302.600 7.300 ;
        RECT 304.085 7.165 304.450 8.880 ;
        RECT 303.860 6.125 304.450 7.165 ;
        RECT 305.125 8.380 305.355 8.950 ;
        RECT 305.125 8.150 307.095 8.380 ;
        RECT 305.125 6.365 305.355 8.150 ;
        RECT 305.585 7.300 306.530 7.710 ;
        RECT 306.770 7.600 307.095 8.150 ;
        RECT 307.545 8.270 307.775 8.950 ;
        RECT 309.695 8.690 310.900 8.920 ;
        RECT 307.545 7.920 308.690 8.270 ;
        RECT 306.770 7.300 308.090 7.600 ;
        RECT 305.585 6.110 305.960 7.300 ;
        RECT 308.350 7.070 308.690 7.920 ;
        RECT 307.545 6.840 308.690 7.070 ;
        RECT 307.545 6.360 307.775 6.840 ;
        RECT 310.020 6.635 310.440 8.440 ;
        RECT 310.670 7.070 310.900 8.690 ;
        RECT 311.140 7.300 311.500 8.905 ;
        RECT 312.860 7.850 313.490 8.905 ;
        RECT 316.830 8.720 319.210 8.950 ;
        RECT 316.830 8.055 317.170 8.720 ;
        RECT 312.040 7.070 312.895 7.200 ;
        RECT 310.670 6.840 312.895 7.070 ;
        RECT 231.390 5.640 234.060 5.980 ;
        RECT 230.260 5.145 231.160 5.525 ;
        RECT 231.390 4.500 231.620 5.640 ;
        RECT 232.255 4.940 234.060 5.340 ;
        RECT 234.290 5.145 235.190 5.525 ;
        RECT 235.860 5.360 236.240 6.095 ;
        RECT 310.670 6.090 311.065 6.840 ;
        RECT 313.160 6.600 313.490 7.850 ;
        RECT 316.755 7.330 317.650 7.710 ;
        RECT 317.300 6.720 317.650 7.330 ;
        RECT 312.725 6.170 313.490 6.600 ;
        RECT 317.880 6.430 318.185 8.285 ;
        RECT 318.870 8.055 319.210 8.720 ;
        RECT 322.390 7.860 322.620 8.940 ;
        RECT 318.415 7.330 319.320 7.710 ;
        RECT 319.550 7.330 320.455 7.710 ;
        RECT 318.980 6.720 319.320 7.330 ;
        RECT 320.115 6.720 320.455 7.330 ;
        RECT 321.755 6.620 322.120 7.750 ;
        RECT 322.390 7.630 323.800 7.860 ;
        RECT 322.360 7.000 323.175 7.380 ;
        RECT 317.880 6.110 319.220 6.430 ;
        RECT 322.360 6.115 322.725 7.000 ;
        RECT 323.410 6.090 323.800 7.630 ;
        RECT 324.165 7.115 324.395 8.950 ;
        RECT 332.130 8.720 334.455 8.950 ;
        RECT 324.650 7.520 325.915 7.750 ;
        RECT 324.165 6.885 325.440 7.115 ;
        RECT 325.685 6.090 325.915 7.520 ;
        RECT 327.420 6.370 327.755 8.270 ;
        RECT 328.745 6.865 328.975 8.540 ;
        RECT 332.130 8.315 332.470 8.720 ;
        RECT 329.265 8.015 330.500 8.270 ;
        RECT 333.150 8.115 333.490 8.475 ;
        RECT 334.225 8.375 334.455 8.720 ;
        RECT 334.685 8.720 336.325 8.950 ;
        RECT 338.040 8.720 340.560 8.950 ;
        RECT 334.685 8.115 334.915 8.720 ;
        RECT 329.265 7.785 332.595 8.015 ;
        RECT 333.150 7.885 334.915 8.115 ;
        RECT 329.265 7.130 329.495 7.785 ;
        RECT 332.315 7.655 332.595 7.785 ;
        RECT 329.785 7.325 331.910 7.555 ;
        RECT 332.315 7.380 334.000 7.655 ;
        RECT 329.785 6.865 330.050 7.325 ;
        RECT 328.745 6.630 330.050 6.865 ;
        RECT 330.290 6.825 333.000 7.095 ;
        RECT 334.280 6.865 334.510 7.885 ;
        RECT 335.145 7.325 335.375 8.485 ;
        RECT 336.095 8.120 336.325 8.720 ;
        RECT 339.170 8.260 340.600 8.490 ;
        RECT 336.095 8.030 338.985 8.120 ;
        RECT 336.095 7.890 339.985 8.030 ;
        RECT 338.795 7.800 339.985 7.890 ;
        RECT 336.605 7.385 338.605 7.660 ;
        RECT 335.145 7.095 336.330 7.325 ;
        RECT 327.430 6.210 327.690 6.370 ;
        RECT 329.710 6.090 330.050 6.630 ;
        RECT 333.595 6.630 335.790 6.865 ;
        RECT 336.025 6.780 336.330 7.095 ;
        RECT 336.605 7.015 336.945 7.385 ;
        RECT 338.375 7.120 338.605 7.385 ;
        RECT 339.750 7.320 339.985 7.800 ;
        RECT 337.795 6.780 338.145 7.115 ;
        RECT 338.375 6.825 339.510 7.120 ;
        RECT 340.280 6.855 340.600 8.260 ;
        RECT 341.525 7.115 341.755 8.950 ;
        RECT 344.215 8.240 344.495 8.940 ;
        RECT 344.215 7.920 345.640 8.240 ;
        RECT 342.010 7.520 343.275 7.750 ;
        RECT 341.525 6.885 342.800 7.115 ;
        RECT 333.595 6.320 333.825 6.630 ;
        RECT 332.100 6.090 333.825 6.320 ;
        RECT 336.025 6.550 338.145 6.780 ;
        RECT 339.960 6.575 340.600 6.855 ;
        RECT 339.960 6.560 340.230 6.575 ;
        RECT 336.025 6.090 336.365 6.550 ;
        RECT 338.445 6.230 340.230 6.560 ;
        RECT 343.045 6.090 343.275 7.520 ;
        RECT 344.025 7.350 345.055 7.690 ;
        RECT 344.750 6.160 345.055 7.350 ;
        RECT 345.285 6.160 345.640 7.920 ;
        RECT 345.870 6.740 346.175 8.880 ;
        RECT 347.125 7.115 347.355 8.950 ;
        RECT 347.610 7.520 348.875 7.750 ;
        RECT 347.125 6.885 348.400 7.115 ;
        RECT 348.645 6.090 348.875 7.520 ;
        RECT 349.365 7.115 349.595 8.950 ;
        RECT 349.850 7.520 351.115 7.750 ;
        RECT 349.365 6.885 350.640 7.115 ;
        RECT 350.885 6.090 351.115 7.520 ;
        RECT 351.605 7.115 351.835 8.950 ;
        RECT 352.090 7.520 353.355 7.750 ;
        RECT 351.605 6.885 352.880 7.115 ;
        RECT 353.125 6.090 353.355 7.520 ;
        RECT 356.085 7.115 356.315 8.950 ;
        RECT 356.570 7.520 357.835 7.750 ;
        RECT 356.085 6.885 357.360 7.115 ;
        RECT 357.605 6.090 357.835 7.520 ;
        RECT 358.325 7.115 358.555 8.950 ;
        RECT 358.810 7.520 360.075 7.750 ;
        RECT 358.325 6.885 359.600 7.115 ;
        RECT 359.845 6.090 360.075 7.520 ;
        RECT 360.565 7.115 360.795 8.950 ;
        RECT 361.050 7.520 362.315 7.750 ;
        RECT 360.565 6.885 361.840 7.115 ;
        RECT 362.085 6.090 362.315 7.520 ;
        RECT 362.805 7.115 363.035 8.950 ;
        RECT 363.290 7.520 364.555 7.750 ;
        RECT 362.805 6.885 364.080 7.115 ;
        RECT 364.325 6.090 364.555 7.520 ;
        RECT 365.045 7.115 365.275 8.950 ;
        RECT 368.505 8.195 368.735 8.785 ;
        RECT 368.505 7.965 370.195 8.195 ;
        RECT 365.530 7.520 366.795 7.750 ;
        RECT 365.045 6.885 366.320 7.115 ;
        RECT 366.565 6.090 366.795 7.520 ;
        RECT 368.310 7.330 369.730 7.710 ;
        RECT 369.965 7.070 370.195 7.965 ;
        RECT 368.405 6.840 370.195 7.070 ;
        RECT 370.425 8.175 370.775 8.775 ;
        RECT 371.825 8.550 373.075 8.780 ;
        RECT 380.370 8.720 382.585 8.950 ;
        RECT 371.825 8.175 372.055 8.550 ;
        RECT 370.425 7.945 372.055 8.175 ;
        RECT 372.285 7.980 372.615 8.320 ;
        RECT 368.405 6.370 368.635 6.840 ;
        RECT 370.425 6.655 370.655 7.945 ;
        RECT 371.050 7.330 372.080 7.710 ;
        RECT 370.425 6.425 370.930 6.655 ;
        RECT 372.385 6.635 372.615 7.980 ;
        RECT 372.845 7.470 373.075 8.550 ;
        RECT 374.325 8.320 374.555 8.515 ;
        RECT 376.925 8.320 377.155 8.690 ;
        RECT 373.305 7.860 373.535 8.320 ;
        RECT 374.325 8.090 377.155 8.320 ;
        RECT 378.600 8.405 379.240 8.635 ;
        RECT 378.015 7.860 378.315 8.085 ;
        RECT 373.305 7.630 378.315 7.860 ;
        RECT 372.385 6.405 372.790 6.635 ;
        RECT 373.625 6.350 373.855 7.630 ;
        RECT 378.600 7.400 378.830 8.405 ;
        RECT 380.370 7.610 380.600 8.720 ;
        RECT 382.355 8.610 382.585 8.720 ;
        RECT 383.395 8.720 384.580 8.950 ;
        RECT 383.395 8.610 383.625 8.720 ;
        RECT 374.850 7.170 378.830 7.400 ;
        RECT 379.710 7.380 380.600 7.610 ;
        RECT 374.205 6.940 374.435 7.150 ;
        RECT 374.205 6.710 377.390 6.940 ;
        RECT 377.160 6.320 377.390 6.710 ;
        RECT 378.150 6.560 378.490 7.170 ;
        RECT 379.085 6.320 379.315 7.150 ;
        RECT 379.710 6.560 380.050 7.380 ;
        RECT 381.050 7.150 381.280 8.085 ;
        RECT 380.280 6.920 381.280 7.150 ;
        RECT 380.280 6.320 380.510 6.920 ;
        RECT 381.575 6.690 381.915 8.490 ;
        RECT 382.355 8.380 383.625 8.610 ;
        RECT 383.890 7.965 384.120 8.490 ;
        RECT 382.155 7.735 384.120 7.965 ;
        RECT 381.110 6.350 381.915 6.690 ;
        RECT 382.820 6.580 383.365 7.390 ;
        RECT 383.890 7.240 384.120 7.735 ;
        RECT 384.350 7.470 384.580 8.720 ;
        RECT 386.635 7.840 387.100 8.940 ;
        RECT 390.695 8.240 390.975 8.940 ;
        RECT 391.830 8.240 392.090 8.270 ;
        RECT 390.695 7.920 392.120 8.240 ;
        RECT 386.635 7.610 387.660 7.840 ;
        RECT 384.810 7.240 386.850 7.315 ;
        RECT 383.890 7.085 386.850 7.240 ;
        RECT 383.890 7.010 385.040 7.085 ;
        RECT 377.160 6.090 380.510 6.320 ;
        RECT 382.820 6.220 384.415 6.580 ;
        RECT 384.810 6.370 385.040 7.010 ;
        RECT 387.300 6.830 387.660 7.610 ;
        RECT 390.505 7.350 391.535 7.690 ;
        RECT 386.635 6.600 387.660 6.830 ;
        RECT 386.635 6.110 387.100 6.600 ;
        RECT 391.230 6.160 391.535 7.350 ;
        RECT 391.765 6.160 392.120 7.920 ;
        RECT 392.350 6.740 392.655 8.880 ;
        RECT 396.300 6.370 396.635 8.270 ;
        RECT 397.525 7.115 397.755 8.950 ;
        RECT 400.335 8.320 400.675 8.940 ;
        RECT 401.900 8.705 404.755 8.940 ;
        RECT 401.900 8.320 402.130 8.705 ;
        RECT 400.335 8.090 402.130 8.320 ;
        RECT 402.430 7.940 403.970 8.270 ;
        RECT 404.415 8.090 404.755 8.705 ;
        RECT 398.010 7.520 399.275 7.750 ;
        RECT 397.525 6.885 398.800 7.115 ;
        RECT 396.310 6.210 396.570 6.370 ;
        RECT 399.045 6.090 399.275 7.520 ;
        RECT 400.690 7.330 401.650 7.710 ;
        RECT 400.690 6.645 401.085 7.330 ;
        RECT 401.880 6.110 402.200 7.710 ;
        RECT 402.430 6.145 402.760 7.940 ;
        RECT 403.000 6.110 403.320 7.710 ;
        RECT 403.560 7.360 404.625 7.710 ;
        RECT 403.560 6.110 403.880 7.360 ;
        RECT 406.945 6.530 407.270 8.510 ;
        RECT 407.500 6.160 407.835 8.930 ;
        RECT 408.825 8.195 409.055 8.785 ;
        RECT 408.825 7.965 410.515 8.195 ;
        RECT 408.760 7.330 410.050 7.710 ;
        RECT 410.285 7.070 410.515 7.965 ;
        RECT 408.725 6.840 410.515 7.070 ;
        RECT 410.745 8.175 411.095 8.775 ;
        RECT 412.145 8.550 413.395 8.780 ;
        RECT 420.690 8.720 422.905 8.950 ;
        RECT 412.145 8.175 412.375 8.550 ;
        RECT 410.745 7.945 412.375 8.175 ;
        RECT 412.605 7.980 412.935 8.320 ;
        RECT 408.725 6.370 408.955 6.840 ;
        RECT 410.745 6.655 410.975 7.945 ;
        RECT 411.370 7.330 412.400 7.710 ;
        RECT 410.745 6.425 411.250 6.655 ;
        RECT 412.705 6.635 412.935 7.980 ;
        RECT 413.165 7.470 413.395 8.550 ;
        RECT 414.645 8.320 414.875 8.515 ;
        RECT 417.245 8.320 417.475 8.690 ;
        RECT 413.625 7.860 413.855 8.320 ;
        RECT 414.645 8.090 417.475 8.320 ;
        RECT 418.920 8.405 419.560 8.635 ;
        RECT 418.335 7.860 418.635 8.085 ;
        RECT 413.625 7.630 418.635 7.860 ;
        RECT 412.705 6.405 413.110 6.635 ;
        RECT 413.945 6.350 414.175 7.630 ;
        RECT 418.920 7.400 419.150 8.405 ;
        RECT 420.690 7.610 420.920 8.720 ;
        RECT 422.675 8.610 422.905 8.720 ;
        RECT 423.715 8.720 424.900 8.950 ;
        RECT 423.715 8.610 423.945 8.720 ;
        RECT 415.170 7.170 419.150 7.400 ;
        RECT 420.030 7.380 420.920 7.610 ;
        RECT 414.525 6.940 414.755 7.150 ;
        RECT 414.525 6.710 417.710 6.940 ;
        RECT 417.480 6.320 417.710 6.710 ;
        RECT 418.470 6.560 418.810 7.170 ;
        RECT 419.405 6.320 419.635 7.150 ;
        RECT 420.030 6.560 420.370 7.380 ;
        RECT 421.370 7.150 421.600 8.085 ;
        RECT 420.600 6.920 421.600 7.150 ;
        RECT 420.600 6.320 420.830 6.920 ;
        RECT 421.895 6.690 422.235 8.490 ;
        RECT 422.675 8.380 423.945 8.610 ;
        RECT 424.210 7.965 424.440 8.490 ;
        RECT 422.475 7.735 424.440 7.965 ;
        RECT 421.430 6.350 422.235 6.690 ;
        RECT 423.140 6.580 423.685 7.390 ;
        RECT 424.210 7.240 424.440 7.735 ;
        RECT 424.670 7.470 424.900 8.720 ;
        RECT 424.210 7.010 426.710 7.240 ;
        RECT 417.480 6.090 420.830 6.320 ;
        RECT 423.140 6.220 424.775 6.580 ;
        RECT 425.130 6.350 425.360 7.010 ;
        RECT 426.955 6.110 427.390 8.940 ;
        RECT 427.765 7.115 427.995 8.950 ;
        RECT 428.250 7.520 429.515 7.750 ;
        RECT 427.765 6.885 429.040 7.115 ;
        RECT 429.285 6.090 429.515 7.520 ;
        RECT 430.005 7.115 430.235 8.950 ;
        RECT 434.430 8.720 436.810 8.950 ;
        RECT 434.430 8.055 434.770 8.720 ;
        RECT 430.490 7.520 431.755 7.750 ;
        RECT 430.005 6.885 431.280 7.115 ;
        RECT 431.525 6.090 431.755 7.520 ;
        RECT 434.355 7.330 435.250 7.710 ;
        RECT 434.900 6.720 435.250 7.330 ;
        RECT 435.480 6.430 435.785 8.285 ;
        RECT 436.470 8.055 436.810 8.720 ;
        RECT 438.965 8.380 439.195 8.950 ;
        RECT 438.965 8.150 440.935 8.380 ;
        RECT 436.015 7.330 436.920 7.710 ;
        RECT 437.150 7.330 438.055 7.710 ;
        RECT 436.580 6.720 436.920 7.330 ;
        RECT 437.715 6.720 438.055 7.330 ;
        RECT 435.480 6.110 436.820 6.430 ;
        RECT 438.965 6.365 439.195 8.150 ;
        RECT 439.425 7.300 440.370 7.710 ;
        RECT 440.610 7.600 440.935 8.150 ;
        RECT 441.385 8.270 441.615 8.950 ;
        RECT 441.385 7.920 442.530 8.270 ;
        RECT 440.610 7.300 441.930 7.600 ;
        RECT 439.425 6.110 439.800 7.300 ;
        RECT 442.190 7.070 442.530 7.920 ;
        RECT 441.385 6.840 442.530 7.070 ;
        RECT 443.445 7.115 443.675 8.950 ;
        RECT 447.825 8.320 448.055 8.940 ;
        RECT 450.065 8.320 450.295 8.940 ;
        RECT 447.825 8.090 450.875 8.320 ;
        RECT 443.930 7.520 445.195 7.750 ;
        RECT 443.445 6.885 444.720 7.115 ;
        RECT 441.385 6.360 441.615 6.840 ;
        RECT 444.965 6.090 445.195 7.520 ;
        RECT 447.210 7.275 450.070 7.710 ;
        RECT 450.540 7.585 450.875 8.090 ;
        RECT 450.540 7.245 454.830 7.585 ;
        RECT 456.900 7.245 460.100 7.590 ;
        RECT 450.540 6.810 450.875 7.245 ;
        RECT 447.925 6.575 450.875 6.810 ;
        RECT 447.925 6.235 448.155 6.575 ;
        RECT 450.165 6.235 450.395 6.575 ;
        RECT 233.830 4.910 234.060 4.940 ;
        RECT 235.860 4.920 236.090 5.360 ;
        RECT 286.700 4.920 289.200 5.220 ;
        RECT 235.860 4.910 289.200 4.920 ;
        RECT 233.830 4.530 289.200 4.910 ;
        RECT 298.310 4.750 298.570 4.910 ;
        RECT 230.260 3.915 231.160 4.295 ;
        RECT 231.390 4.100 233.195 4.500 ;
        RECT 233.830 3.800 234.060 4.530 ;
        RECT 235.860 4.520 289.200 4.530 ;
        RECT 234.290 3.915 235.190 4.295 ;
        RECT 235.860 4.080 236.090 4.520 ;
        RECT 286.700 4.220 289.200 4.520 ;
        RECT 231.390 3.460 234.060 3.800 ;
        RECT 223.200 2.700 224.400 3.300 ;
        RECT 232.545 2.710 232.945 3.460 ;
        RECT 235.860 3.345 236.240 4.080 ;
        RECT 234.290 3.180 236.240 3.345 ;
        RECT 234.290 3.115 236.090 3.180 ;
        RECT 230.525 2.390 232.945 2.710 ;
        RECT 235.860 2.630 236.090 3.115 ;
        RECT 298.300 2.850 298.635 4.750 ;
        RECT 301.985 4.280 302.215 4.760 ;
        RECT 301.070 4.050 302.215 4.280 ;
        RECT 301.070 3.200 301.410 4.050 ;
        RECT 303.800 3.820 304.175 5.010 ;
        RECT 301.670 3.520 302.990 3.820 ;
        RECT 301.070 2.850 302.215 3.200 ;
        RECT 230.525 1.965 230.925 2.390 ;
        RECT 301.985 2.170 302.215 2.850 ;
        RECT 302.665 2.970 302.990 3.520 ;
        RECT 303.230 3.410 304.175 3.820 ;
        RECT 304.405 2.970 304.635 4.755 ;
        RECT 302.665 2.740 304.635 2.970 ;
        RECT 306.140 2.850 306.475 4.750 ;
        RECT 308.430 4.490 308.770 5.030 ;
        RECT 310.820 4.800 312.545 5.030 ;
        RECT 307.465 4.255 308.770 4.490 ;
        RECT 312.315 4.490 312.545 4.800 ;
        RECT 314.745 4.570 315.085 5.030 ;
        RECT 304.405 2.170 304.635 2.740 ;
        RECT 307.465 2.580 307.695 4.255 ;
        RECT 307.985 3.335 308.215 3.990 ;
        RECT 308.505 3.795 308.770 4.255 ;
        RECT 309.010 4.025 311.720 4.295 ;
        RECT 312.315 4.255 314.510 4.490 ;
        RECT 314.745 4.340 316.865 4.570 ;
        RECT 317.165 4.560 318.950 4.890 ;
        RECT 308.505 3.565 310.630 3.795 ;
        RECT 311.035 3.465 312.720 3.740 ;
        RECT 311.035 3.335 311.315 3.465 ;
        RECT 307.985 3.105 311.315 3.335 ;
        RECT 313.000 3.235 313.230 4.255 ;
        RECT 314.745 4.025 315.050 4.340 ;
        RECT 313.865 3.795 315.050 4.025 ;
        RECT 307.985 2.850 309.220 3.105 ;
        RECT 311.870 3.005 313.635 3.235 ;
        RECT 310.850 2.400 311.190 2.805 ;
        RECT 311.870 2.645 312.210 3.005 ;
        RECT 312.945 2.400 313.175 2.745 ;
        RECT 310.850 2.170 313.175 2.400 ;
        RECT 313.405 2.400 313.635 3.005 ;
        RECT 313.865 2.635 314.095 3.795 ;
        RECT 315.325 3.735 315.665 4.105 ;
        RECT 316.515 4.005 316.865 4.340 ;
        RECT 318.680 4.545 318.950 4.560 ;
        RECT 317.095 4.000 318.230 4.295 ;
        RECT 318.680 4.265 319.320 4.545 ;
        RECT 317.095 3.735 317.325 4.000 ;
        RECT 315.325 3.460 317.325 3.735 ;
        RECT 318.470 3.320 318.705 3.800 ;
        RECT 317.515 3.230 318.705 3.320 ;
        RECT 314.815 3.090 318.705 3.230 ;
        RECT 314.815 3.000 317.705 3.090 ;
        RECT 314.815 2.400 315.045 3.000 ;
        RECT 319.000 2.860 319.320 4.265 ;
        RECT 317.890 2.630 319.320 2.860 ;
        RECT 321.265 2.610 321.590 4.590 ;
        RECT 313.405 2.170 315.045 2.400 ;
        RECT 316.760 2.170 319.280 2.400 ;
        RECT 321.820 2.190 322.155 4.960 ;
        RECT 326.870 4.750 327.130 4.910 ;
        RECT 324.565 2.850 324.900 4.750 ;
        RECT 326.805 2.850 327.140 4.750 ;
        RECT 329.390 3.955 329.980 4.995 ;
        RECT 329.390 2.240 329.755 3.955 ;
        RECT 331.240 3.820 331.615 4.525 ;
        RECT 330.050 3.040 330.390 3.680 ;
        RECT 330.730 3.410 331.615 3.820 ;
        RECT 331.845 3.040 332.075 4.995 ;
        RECT 330.050 2.805 332.075 3.040 ;
        RECT 331.745 2.180 332.075 2.805 ;
        RECT 332.565 4.005 333.840 4.235 ;
        RECT 332.565 2.170 332.795 4.005 ;
        RECT 334.085 3.600 334.315 5.030 ;
        RECT 333.050 3.370 334.315 3.600 ;
        RECT 336.485 4.005 337.760 4.235 ;
        RECT 336.485 2.170 336.715 4.005 ;
        RECT 338.005 3.600 338.235 5.030 ;
        RECT 336.970 3.370 338.235 3.600 ;
        RECT 338.725 4.005 340.000 4.235 ;
        RECT 338.725 2.170 338.955 4.005 ;
        RECT 340.245 3.600 340.475 5.030 ;
        RECT 339.210 3.370 340.475 3.600 ;
        RECT 340.965 4.005 342.240 4.235 ;
        RECT 340.965 2.170 341.195 4.005 ;
        RECT 342.485 3.600 342.715 5.030 ;
        RECT 344.545 4.280 344.775 4.760 ;
        RECT 341.450 3.370 342.715 3.600 ;
        RECT 343.630 4.050 344.775 4.280 ;
        RECT 343.630 3.200 343.970 4.050 ;
        RECT 346.360 3.820 346.735 5.010 ;
        RECT 344.230 3.520 345.550 3.820 ;
        RECT 343.630 2.850 344.775 3.200 ;
        RECT 344.545 2.170 344.775 2.850 ;
        RECT 345.225 2.970 345.550 3.520 ;
        RECT 345.790 3.410 346.735 3.820 ;
        RECT 346.965 2.970 347.195 4.755 ;
        RECT 345.225 2.740 347.195 2.970 ;
        RECT 346.965 2.170 347.195 2.740 ;
        RECT 348.085 2.190 348.420 4.960 ;
        RECT 348.650 2.610 348.975 4.590 ;
        RECT 350.940 2.850 351.275 4.750 ;
        RECT 352.165 4.005 353.440 4.235 ;
        RECT 352.165 2.170 352.395 4.005 ;
        RECT 353.685 3.600 353.915 5.030 ;
        RECT 364.280 4.800 367.630 5.030 ;
        RECT 369.940 4.850 371.575 4.900 ;
        RECT 355.525 4.280 355.755 4.750 ;
        RECT 357.545 4.465 358.050 4.695 ;
        RECT 359.505 4.485 359.910 4.715 ;
        RECT 355.525 4.050 357.315 4.280 ;
        RECT 352.650 3.370 353.915 3.600 ;
        RECT 355.560 3.410 356.850 3.790 ;
        RECT 357.085 3.155 357.315 4.050 ;
        RECT 355.625 2.925 357.315 3.155 ;
        RECT 357.545 3.175 357.775 4.465 ;
        RECT 358.170 3.410 359.200 3.790 ;
        RECT 357.545 2.945 359.175 3.175 ;
        RECT 359.505 3.140 359.735 4.485 ;
        RECT 355.625 2.335 355.855 2.925 ;
        RECT 357.545 2.345 357.895 2.945 ;
        RECT 358.945 2.570 359.175 2.945 ;
        RECT 359.405 2.800 359.735 3.140 ;
        RECT 359.965 2.570 360.195 3.650 ;
        RECT 360.745 3.490 360.975 4.770 ;
        RECT 364.280 4.410 364.510 4.800 ;
        RECT 361.325 4.180 364.510 4.410 ;
        RECT 361.325 3.970 361.555 4.180 ;
        RECT 365.270 3.950 365.610 4.560 ;
        RECT 366.205 3.970 366.435 4.800 ;
        RECT 361.970 3.720 365.950 3.950 ;
        RECT 360.425 3.260 365.435 3.490 ;
        RECT 360.425 2.800 360.655 3.260 ;
        RECT 365.135 3.035 365.435 3.260 ;
        RECT 361.445 2.800 364.275 3.030 ;
        RECT 361.445 2.605 361.675 2.800 ;
        RECT 358.945 2.340 360.195 2.570 ;
        RECT 364.045 2.430 364.275 2.800 ;
        RECT 365.720 2.715 365.950 3.720 ;
        RECT 366.830 3.740 367.170 4.560 ;
        RECT 367.400 4.200 367.630 4.800 ;
        RECT 368.230 4.430 369.035 4.770 ;
        RECT 369.930 4.590 371.575 4.850 ;
        RECT 367.400 3.970 368.400 4.200 ;
        RECT 366.830 3.510 367.720 3.740 ;
        RECT 365.720 2.485 366.360 2.715 ;
        RECT 367.490 2.400 367.720 3.510 ;
        RECT 368.170 3.035 368.400 3.970 ;
        RECT 368.695 2.630 369.035 4.430 ;
        RECT 369.940 4.540 371.575 4.590 ;
        RECT 369.940 3.730 370.485 4.540 ;
        RECT 371.930 4.110 372.160 4.770 ;
        RECT 371.010 3.880 373.510 4.110 ;
        RECT 371.010 3.385 371.240 3.880 ;
        RECT 369.275 3.155 371.240 3.385 ;
        RECT 369.475 2.510 370.745 2.740 ;
        RECT 371.010 2.630 371.240 3.155 ;
        RECT 369.475 2.400 369.705 2.510 ;
        RECT 367.490 2.170 369.705 2.400 ;
        RECT 370.515 2.400 370.745 2.510 ;
        RECT 371.470 2.400 371.700 3.650 ;
        RECT 370.515 2.170 371.700 2.400 ;
        RECT 373.755 2.180 374.190 5.010 ;
        RECT 375.685 4.005 376.960 4.235 ;
        RECT 375.685 2.170 375.915 4.005 ;
        RECT 377.205 3.600 377.435 5.030 ;
        RECT 376.170 3.370 377.435 3.600 ;
        RECT 377.925 4.005 379.200 4.235 ;
        RECT 377.925 2.170 378.155 4.005 ;
        RECT 379.445 3.600 379.675 5.030 ;
        RECT 378.410 3.370 379.675 3.600 ;
        RECT 380.165 4.005 381.440 4.235 ;
        RECT 380.165 2.170 380.395 4.005 ;
        RECT 381.685 3.600 381.915 5.030 ;
        RECT 380.650 3.370 381.915 3.600 ;
        RECT 382.405 4.005 383.680 4.235 ;
        RECT 382.405 2.170 382.635 4.005 ;
        RECT 383.925 3.600 384.155 5.030 ;
        RECT 382.890 3.370 384.155 3.600 ;
        RECT 386.325 2.980 386.555 4.760 ;
        RECT 386.785 3.930 387.300 4.910 ;
        RECT 388.410 3.960 389.035 4.985 ;
        RECT 392.885 4.510 393.115 5.030 ;
        RECT 395.125 4.510 395.355 5.030 ;
        RECT 386.785 3.370 387.670 3.930 ;
        RECT 388.050 2.980 388.335 3.730 ;
        RECT 386.325 2.745 388.335 2.980 ;
        RECT 386.325 2.170 386.710 2.745 ;
        RECT 388.565 2.180 389.035 3.960 ;
        RECT 391.825 4.240 395.355 4.510 ;
        RECT 397.975 4.615 398.370 5.030 ;
        RECT 399.720 4.800 401.160 5.030 ;
        RECT 399.720 4.615 399.950 4.800 ;
        RECT 397.975 4.380 399.950 4.615 ;
        RECT 400.930 4.615 401.160 4.800 ;
        RECT 401.960 4.800 403.400 5.030 ;
        RECT 401.960 4.615 402.190 4.800 ;
        RECT 391.825 2.760 392.095 4.240 ;
        RECT 400.190 4.150 400.630 4.550 ;
        RECT 400.930 4.380 402.190 4.615 ;
        RECT 403.170 4.615 403.400 4.800 ;
        RECT 404.670 4.615 405.540 5.030 ;
        RECT 406.440 4.615 407.880 5.030 ;
        RECT 409.180 4.615 409.570 5.030 ;
        RECT 402.420 4.150 402.870 4.550 ;
        RECT 403.170 4.380 409.570 4.615 ;
        RECT 392.330 3.410 393.240 3.790 ;
        RECT 393.500 3.410 395.240 3.790 ;
        RECT 392.940 3.180 393.240 3.410 ;
        RECT 395.660 3.180 395.910 3.980 ;
        RECT 398.510 3.920 404.455 4.150 ;
        RECT 406.270 3.920 408.900 4.150 ;
        RECT 397.125 3.690 398.290 3.810 ;
        RECT 404.690 3.690 405.750 3.810 ;
        RECT 397.125 3.410 405.750 3.690 ;
        RECT 392.940 2.860 395.910 3.180 ;
        RECT 396.965 2.760 404.940 2.990 ;
        RECT 391.825 2.525 392.625 2.760 ;
        RECT 392.395 2.420 392.625 2.525 ;
        RECT 392.395 2.190 394.330 2.420 ;
        RECT 396.965 2.180 397.195 2.760 ;
        RECT 401.345 2.180 401.575 2.760 ;
        RECT 404.710 2.400 404.940 2.760 ;
        RECT 406.270 2.710 406.680 3.920 ;
        RECT 409.140 3.685 409.570 4.380 ;
        RECT 406.910 3.450 409.570 3.685 ;
        RECT 406.910 2.650 407.275 3.450 ;
        RECT 408.065 2.400 408.295 3.030 ;
        RECT 409.180 2.650 409.570 3.450 ;
        RECT 411.525 4.005 412.800 4.235 ;
        RECT 410.305 2.400 410.535 3.030 ;
        RECT 404.710 2.170 410.535 2.400 ;
        RECT 411.525 2.170 411.755 4.005 ;
        RECT 413.045 3.600 413.275 5.030 ;
        RECT 412.010 3.370 413.275 3.600 ;
        RECT 414.885 4.005 416.160 4.235 ;
        RECT 414.885 2.170 415.115 4.005 ;
        RECT 416.405 3.600 416.635 5.030 ;
        RECT 415.370 3.370 416.635 3.600 ;
        RECT 417.125 4.005 418.400 4.235 ;
        RECT 417.125 2.170 417.355 4.005 ;
        RECT 418.645 3.600 418.875 5.030 ;
        RECT 417.610 3.370 418.875 3.600 ;
        RECT 419.365 4.005 420.640 4.235 ;
        RECT 419.365 2.170 419.595 4.005 ;
        RECT 420.885 3.600 421.115 5.030 ;
        RECT 419.850 3.370 421.115 3.600 ;
        RECT 421.605 4.005 422.880 4.235 ;
        RECT 421.605 2.170 421.835 4.005 ;
        RECT 423.125 3.600 423.355 5.030 ;
        RECT 422.090 3.370 423.355 3.600 ;
        RECT 423.845 4.005 425.120 4.235 ;
        RECT 423.845 2.170 424.075 4.005 ;
        RECT 425.365 3.600 425.595 5.030 ;
        RECT 424.330 3.370 425.595 3.600 ;
        RECT 426.190 4.520 426.955 4.950 ;
        RECT 426.190 3.270 426.520 4.520 ;
        RECT 428.615 4.280 429.010 5.030 ;
        RECT 432.220 4.690 433.560 5.010 ;
        RECT 426.785 4.050 429.010 4.280 ;
        RECT 426.785 3.920 427.640 4.050 ;
        RECT 426.190 2.215 426.820 3.270 ;
        RECT 428.180 2.215 428.540 3.820 ;
        RECT 428.780 2.430 429.010 4.050 ;
        RECT 429.240 2.680 429.660 4.485 ;
        RECT 430.985 3.790 431.325 4.400 ;
        RECT 432.120 3.790 432.460 4.400 ;
        RECT 430.985 3.410 431.890 3.790 ;
        RECT 432.120 3.410 433.025 3.790 ;
        RECT 428.780 2.200 429.985 2.430 ;
        RECT 432.230 2.400 432.570 3.065 ;
        RECT 433.255 2.835 433.560 4.690 ;
        RECT 433.790 3.790 434.140 4.400 ;
        RECT 433.790 3.410 434.685 3.790 ;
        RECT 434.270 2.400 434.610 3.065 ;
        RECT 432.230 2.170 434.610 2.400 ;
        RECT 435.505 2.240 435.810 4.380 ;
        RECT 436.040 3.200 436.395 4.960 ;
        RECT 436.625 3.770 436.930 4.960 ;
        RECT 439.525 4.545 439.755 4.885 ;
        RECT 441.765 4.545 441.995 4.885 ;
        RECT 439.525 4.310 442.475 4.545 ;
        RECT 442.140 3.875 442.475 4.310 ;
        RECT 436.625 3.430 437.655 3.770 ;
        RECT 438.810 3.410 441.670 3.845 ;
        RECT 442.140 3.535 446.430 3.875 ;
        RECT 436.040 2.880 437.465 3.200 ;
        RECT 442.140 3.030 442.475 3.535 ;
        RECT 448.500 3.530 451.700 3.875 ;
        RECT 437.185 2.180 437.465 2.880 ;
        RECT 439.425 2.800 442.475 3.030 ;
        RECT 454.085 2.970 454.315 4.755 ;
        RECT 454.545 3.820 454.920 5.010 ;
        RECT 456.505 4.280 456.735 4.760 ;
        RECT 456.505 4.050 457.650 4.280 ;
        RECT 454.545 3.410 455.490 3.820 ;
        RECT 455.730 3.520 457.050 3.820 ;
        RECT 455.730 2.970 456.055 3.520 ;
        RECT 457.310 3.200 457.650 4.050 ;
        RECT 439.425 2.180 439.655 2.800 ;
        RECT 441.665 2.180 441.895 2.800 ;
        RECT 454.085 2.740 456.055 2.970 ;
        RECT 456.505 2.850 457.650 3.200 ;
        RECT 458.565 4.005 459.840 4.235 ;
        RECT 454.085 2.170 454.315 2.740 ;
        RECT 456.505 2.170 456.735 2.850 ;
        RECT 458.565 2.170 458.795 4.005 ;
        RECT 460.085 3.600 460.315 5.030 ;
        RECT 459.050 3.370 460.315 3.600 ;
        RECT 230.290 1.735 231.160 1.965 ;
        RECT 231.390 1.280 232.945 1.620 ;
        RECT 230.290 0.935 231.160 1.165 ;
        RECT 181.460 0.515 181.690 0.570 ;
        RECT 179.705 0.285 181.690 0.515 ;
        RECT 181.460 0.230 181.690 0.285 ;
        RECT 187.020 0.250 187.620 0.570 ;
        RECT 232.545 0.335 232.945 1.280 ;
        RECT 181.920 -0.115 186.790 0.115 ;
        RECT 181.460 -0.285 181.690 -0.230 ;
        RECT 175.905 -1.390 177.855 -1.010 ;
        RECT 179.705 -0.515 181.690 -0.285 ;
        RECT 171.405 -3.190 172.305 -2.810 ;
        RECT 174.855 -3.190 176.805 -2.810 ;
        RECT 171.655 -5.185 172.055 -3.190 ;
        RECT 179.705 -4.050 180.005 -0.515 ;
        RECT 181.460 -0.570 181.690 -0.515 ;
        RECT 187.020 -0.250 192.105 0.250 ;
        RECT 232.295 -0.065 233.195 0.335 ;
        RECT 187.020 -0.570 187.620 -0.250 ;
        RECT 181.920 -0.915 184.505 -0.685 ;
        RECT 180.625 -1.030 181.525 -1.010 ;
        RECT 180.625 -1.370 181.690 -1.030 ;
        RECT 180.625 -1.390 181.525 -1.370 ;
        RECT 181.920 -2.810 182.790 -1.485 ;
        RECT 181.905 -3.190 182.805 -2.810 ;
        RECT 179.665 -4.950 180.045 -4.050 ;
        RECT 179.705 -5.000 180.005 -4.950 ;
        RECT 171.420 -5.415 172.290 -5.185 ;
        RECT 172.520 -5.900 172.750 -5.530 ;
        RECT 172.520 -5.910 181.855 -5.900 ;
        RECT 172.520 -6.290 182.305 -5.910 ;
        RECT 172.520 -6.300 181.855 -6.290 ;
        RECT 172.520 -6.670 172.750 -6.300 ;
        RECT 171.420 -7.850 172.290 -6.785 ;
        RECT 184.205 -7.850 184.505 -0.915 ;
        RECT 185.405 -5.950 186.305 -5.910 ;
        RECT 187.320 -5.950 187.620 -0.570 ;
        RECT 185.405 -6.250 187.620 -5.950 ;
        RECT 185.405 -6.290 186.305 -6.250 ;
        RECT 171.420 -8.150 184.505 -7.850 ;
        RECT 184.205 -10.305 184.505 -8.150 ;
        RECT 191.600 -8.830 192.100 -0.250 ;
        RECT 230.260 -0.445 231.160 -0.065 ;
        RECT 234.290 -0.445 235.190 -0.065 ;
        RECT 235.860 -0.280 236.090 0.270 ;
        RECT 231.390 -0.900 234.060 -0.560 ;
        RECT 223.320 -2.810 224.520 -2.700 ;
        RECT 232.545 -2.810 232.945 -0.900 ;
        RECT 235.860 -1.015 236.240 -0.280 ;
        RECT 297.285 -0.725 297.515 1.110 ;
        RECT 297.770 -0.320 299.035 -0.090 ;
        RECT 297.285 -0.955 298.560 -0.725 ;
        RECT 234.290 -1.180 236.240 -1.015 ;
        RECT 234.290 -1.245 236.090 -1.180 ;
        RECT 235.860 -1.730 236.090 -1.245 ;
        RECT 298.805 -1.750 299.035 -0.320 ;
        RECT 299.525 -0.725 299.755 1.110 ;
        RECT 302.795 0.860 304.730 1.090 ;
        RECT 302.795 0.755 303.025 0.860 ;
        RECT 302.225 0.520 303.025 0.755 ;
        RECT 300.010 -0.320 301.275 -0.090 ;
        RECT 299.525 -0.955 300.800 -0.725 ;
        RECT 301.045 -1.750 301.275 -0.320 ;
        RECT 302.225 -0.960 302.495 0.520 ;
        RECT 303.340 0.100 306.310 0.420 ;
        RECT 303.340 -0.130 303.640 0.100 ;
        RECT 302.730 -0.510 303.640 -0.130 ;
        RECT 303.900 -0.510 305.640 -0.130 ;
        RECT 306.060 -0.700 306.310 0.100 ;
        RECT 307.365 -0.725 307.595 1.110 ;
        RECT 307.850 -0.320 309.115 -0.090 ;
        RECT 307.365 -0.955 308.640 -0.725 ;
        RECT 302.225 -1.230 305.755 -0.960 ;
        RECT 303.285 -1.750 303.515 -1.230 ;
        RECT 305.525 -1.250 305.755 -1.230 ;
        RECT 305.525 -1.630 305.850 -1.250 ;
        RECT 305.525 -1.750 305.755 -1.630 ;
        RECT 308.885 -1.750 309.115 -0.320 ;
        RECT 309.605 -0.725 309.835 1.110 ;
        RECT 310.090 -0.320 311.355 -0.090 ;
        RECT 309.605 -0.955 310.880 -0.725 ;
        RECT 311.125 -1.750 311.355 -0.320 ;
        RECT 311.845 -0.725 312.075 1.110 ;
        RECT 318.605 0.880 320.925 1.110 ;
        RECT 318.605 0.080 318.835 0.880 ;
        RECT 319.065 0.310 320.450 0.650 ;
        RECT 312.330 -0.320 313.595 -0.090 ;
        RECT 311.845 -0.955 313.120 -0.725 ;
        RECT 313.365 -1.750 313.595 -0.320 ;
        RECT 317.330 -0.380 318.305 -0.130 ;
        RECT 318.605 -0.150 319.195 0.080 ;
        RECT 317.330 -0.680 318.735 -0.380 ;
        RECT 318.400 -1.730 318.735 -0.680 ;
        RECT 318.965 -1.730 319.195 -0.150 ;
        RECT 319.520 -1.730 319.855 0.040 ;
        RECT 320.085 -1.730 320.450 0.310 ;
        RECT 320.695 0.410 320.925 0.880 ;
        RECT 320.695 0.180 321.435 0.410 ;
        RECT 320.680 -1.730 320.975 -0.050 ;
        RECT 321.205 -1.730 321.435 0.180 ;
        RECT 323.445 -1.470 323.780 0.430 ;
        RECT 324.165 -0.725 324.395 1.110 ;
        RECT 328.185 0.355 328.415 0.945 ;
        RECT 328.185 0.125 329.875 0.355 ;
        RECT 324.650 -0.320 325.915 -0.090 ;
        RECT 324.165 -0.955 325.440 -0.725 ;
        RECT 323.510 -1.630 323.770 -1.470 ;
        RECT 325.685 -1.750 325.915 -0.320 ;
        RECT 328.120 -0.510 329.410 -0.130 ;
        RECT 329.645 -0.770 329.875 0.125 ;
        RECT 328.085 -1.000 329.875 -0.770 ;
        RECT 330.105 0.335 330.455 0.935 ;
        RECT 331.505 0.710 332.755 0.940 ;
        RECT 340.050 0.880 342.265 1.110 ;
        RECT 331.505 0.335 331.735 0.710 ;
        RECT 330.105 0.105 331.735 0.335 ;
        RECT 331.965 0.140 332.295 0.480 ;
        RECT 328.085 -1.470 328.315 -1.000 ;
        RECT 330.105 -1.185 330.335 0.105 ;
        RECT 330.730 -0.510 331.760 -0.130 ;
        RECT 330.105 -1.415 330.610 -1.185 ;
        RECT 332.065 -1.205 332.295 0.140 ;
        RECT 332.525 -0.370 332.755 0.710 ;
        RECT 334.005 0.480 334.235 0.675 ;
        RECT 336.605 0.480 336.835 0.850 ;
        RECT 332.985 0.020 333.215 0.480 ;
        RECT 334.005 0.250 336.835 0.480 ;
        RECT 338.280 0.565 338.920 0.795 ;
        RECT 337.695 0.020 337.995 0.245 ;
        RECT 332.985 -0.210 337.995 0.020 ;
        RECT 332.065 -1.435 332.470 -1.205 ;
        RECT 333.305 -1.490 333.535 -0.210 ;
        RECT 338.280 -0.440 338.510 0.565 ;
        RECT 340.050 -0.230 340.280 0.880 ;
        RECT 342.035 0.770 342.265 0.880 ;
        RECT 343.075 0.880 344.260 1.110 ;
        RECT 343.075 0.770 343.305 0.880 ;
        RECT 334.530 -0.670 338.510 -0.440 ;
        RECT 339.390 -0.460 340.280 -0.230 ;
        RECT 333.885 -0.900 334.115 -0.690 ;
        RECT 333.885 -1.130 337.070 -0.900 ;
        RECT 336.840 -1.520 337.070 -1.130 ;
        RECT 337.830 -1.280 338.170 -0.670 ;
        RECT 338.765 -1.520 338.995 -0.690 ;
        RECT 339.390 -1.280 339.730 -0.460 ;
        RECT 340.730 -0.690 340.960 0.245 ;
        RECT 339.960 -0.920 340.960 -0.690 ;
        RECT 339.960 -1.520 340.190 -0.920 ;
        RECT 341.255 -1.150 341.595 0.650 ;
        RECT 342.035 0.540 343.305 0.770 ;
        RECT 343.570 0.125 343.800 0.650 ;
        RECT 341.835 -0.105 343.800 0.125 ;
        RECT 340.790 -1.490 341.595 -1.150 ;
        RECT 342.500 -1.260 343.045 -0.450 ;
        RECT 343.570 -0.600 343.800 -0.105 ;
        RECT 344.030 -0.370 344.260 0.880 ;
        RECT 343.570 -0.830 346.070 -0.600 ;
        RECT 336.840 -1.750 340.190 -1.520 ;
        RECT 342.500 -1.620 344.135 -1.260 ;
        RECT 344.490 -1.490 344.720 -0.830 ;
        RECT 346.315 -1.730 346.750 1.100 ;
        RECT 347.585 -0.670 347.910 1.040 ;
        RECT 348.200 0.860 351.245 1.090 ;
        RECT 348.200 -1.185 348.430 0.860 ;
        RECT 348.680 -0.090 349.040 0.565 ;
        RECT 349.320 0.400 350.715 0.630 ;
        RECT 348.680 -0.595 349.595 -0.090 ;
        RECT 347.125 -1.415 349.595 -1.185 ;
        RECT 347.125 -1.730 347.355 -1.415 ;
        RECT 349.365 -1.730 349.595 -1.415 ;
        RECT 349.825 -1.730 350.120 -0.060 ;
        RECT 350.360 -1.730 350.715 0.400 ;
        RECT 351.015 0.400 351.245 0.860 ;
        RECT 356.085 0.475 356.415 1.100 ;
        RECT 351.015 0.170 351.835 0.400 ;
        RECT 350.945 -1.730 351.260 -0.060 ;
        RECT 351.605 -1.730 351.835 0.170 ;
        RECT 353.740 -1.470 354.075 0.430 ;
        RECT 356.085 0.240 358.110 0.475 ;
        RECT 353.750 -1.630 354.010 -1.470 ;
        RECT 356.085 -1.715 356.315 0.240 ;
        RECT 356.545 -0.540 357.430 -0.130 ;
        RECT 357.770 -0.400 358.110 0.240 ;
        RECT 356.545 -1.245 356.920 -0.540 ;
        RECT 358.405 -0.675 358.770 1.040 ;
        RECT 361.070 0.880 363.450 1.110 ;
        RECT 361.070 0.215 361.410 0.880 ;
        RECT 360.995 -0.510 361.890 -0.130 ;
        RECT 358.180 -1.715 358.770 -0.675 ;
        RECT 361.540 -1.120 361.890 -0.510 ;
        RECT 362.120 -1.410 362.425 0.445 ;
        RECT 363.110 0.215 363.450 0.880 ;
        RECT 362.655 -0.510 363.560 -0.130 ;
        RECT 363.790 -0.510 364.695 -0.130 ;
        RECT 363.220 -1.120 363.560 -0.510 ;
        RECT 364.355 -1.120 364.695 -0.510 ;
        RECT 365.605 -0.725 365.835 1.110 ;
        RECT 369.510 0.880 371.890 1.110 ;
        RECT 369.510 0.215 369.850 0.880 ;
        RECT 366.090 -0.320 367.355 -0.090 ;
        RECT 365.605 -0.955 366.880 -0.725 ;
        RECT 362.120 -1.730 363.460 -1.410 ;
        RECT 367.125 -1.750 367.355 -0.320 ;
        RECT 368.265 -0.510 369.170 -0.130 ;
        RECT 369.400 -0.510 370.305 -0.130 ;
        RECT 368.265 -1.120 368.605 -0.510 ;
        RECT 369.400 -1.120 369.740 -0.510 ;
        RECT 370.535 -1.410 370.840 0.445 ;
        RECT 371.550 0.215 371.890 0.880 ;
        RECT 371.070 -0.510 371.965 -0.130 ;
        RECT 371.070 -1.120 371.420 -0.510 ;
        RECT 372.325 -0.725 372.555 1.110 ;
        RECT 372.810 -0.320 374.075 -0.090 ;
        RECT 372.325 -0.955 373.600 -0.725 ;
        RECT 369.500 -1.730 370.840 -1.410 ;
        RECT 373.845 -1.750 374.075 -0.320 ;
        RECT 374.565 -0.725 374.795 1.110 ;
        RECT 375.050 -0.320 376.315 -0.090 ;
        RECT 374.565 -0.955 375.840 -0.725 ;
        RECT 376.085 -1.750 376.315 -0.320 ;
        RECT 376.805 -0.725 377.035 1.110 ;
        RECT 377.290 -0.320 378.555 -0.090 ;
        RECT 376.805 -0.955 378.080 -0.725 ;
        RECT 378.325 -1.750 378.555 -0.320 ;
        RECT 379.045 -0.725 379.275 1.110 ;
        RECT 379.530 -0.320 380.795 -0.090 ;
        RECT 379.045 -0.955 380.320 -0.725 ;
        RECT 380.565 -1.750 380.795 -0.320 ;
        RECT 382.310 -1.080 382.635 -0.080 ;
        RECT 382.865 -1.750 383.195 1.110 ;
        RECT 384.085 0.345 384.315 1.110 ;
        RECT 386.515 0.420 386.745 1.110 ;
        RECT 384.085 0.110 385.970 0.345 ;
        RECT 384.085 -1.710 384.315 0.110 ;
        RECT 384.545 -0.655 385.490 -0.130 ;
        RECT 385.740 -0.390 385.970 0.110 ;
        RECT 386.515 -0.070 387.640 0.420 ;
        RECT 384.545 -1.670 384.855 -0.655 ;
        RECT 385.740 -0.730 387.080 -0.390 ;
        RECT 387.320 -0.980 387.640 -0.070 ;
        RECT 386.515 -1.215 387.640 -0.980 ;
        RECT 389.685 0.345 389.915 1.110 ;
        RECT 392.115 0.420 392.345 1.110 ;
        RECT 396.905 0.455 397.135 1.100 ;
        RECT 392.950 0.420 393.210 0.430 ;
        RECT 389.685 0.110 391.570 0.345 ;
        RECT 386.515 -1.710 386.745 -1.215 ;
        RECT 389.685 -1.710 389.915 0.110 ;
        RECT 390.145 -0.655 391.090 -0.130 ;
        RECT 391.340 -0.390 391.570 0.110 ;
        RECT 392.115 -0.070 393.240 0.420 ;
        RECT 390.145 -1.670 390.455 -0.655 ;
        RECT 391.340 -0.730 392.680 -0.390 ;
        RECT 392.920 -0.980 393.240 -0.070 ;
        RECT 392.115 -1.215 393.240 -0.980 ;
        RECT 395.690 0.080 397.135 0.455 ;
        RECT 395.690 -0.775 396.070 0.080 ;
        RECT 397.365 -0.160 397.695 0.595 ;
        RECT 399.905 0.400 400.135 1.100 ;
        RECT 401.860 0.400 402.220 1.100 ;
        RECT 396.430 -0.545 397.695 -0.160 ;
        RECT 395.690 -1.010 397.035 -0.775 ;
        RECT 392.115 -1.710 392.345 -1.215 ;
        RECT 396.805 -1.600 397.035 -1.010 ;
        RECT 397.365 -1.090 397.695 -0.545 ;
        RECT 398.950 0.080 402.220 0.400 ;
        RECT 398.950 -0.745 399.180 0.080 ;
        RECT 399.410 -0.480 402.820 -0.160 ;
        RECT 398.950 -1.015 399.980 -0.745 ;
        RECT 399.620 -1.280 399.980 -1.015 ;
        RECT 400.280 -1.040 402.820 -0.720 ;
        RECT 399.620 -1.600 401.290 -1.280 ;
        RECT 404.700 -1.470 405.035 0.430 ;
        RECT 405.925 -0.725 406.155 1.110 ;
        RECT 409.140 0.400 409.590 1.110 ;
        RECT 409.140 0.080 410.600 0.400 ;
        RECT 406.410 -0.320 407.675 -0.090 ;
        RECT 405.925 -0.955 407.200 -0.725 ;
        RECT 404.710 -1.630 404.970 -1.470 ;
        RECT 407.445 -1.750 407.675 -0.320 ;
        RECT 408.550 -0.575 410.070 -0.160 ;
        RECT 410.300 -0.805 410.600 0.080 ;
        RECT 409.315 -1.060 410.600 -0.805 ;
        RECT 409.315 -1.250 409.545 -1.060 ;
        RECT 409.190 -1.630 409.545 -1.250 ;
        RECT 409.315 -1.750 409.545 -1.630 ;
        RECT 411.925 -1.750 412.255 1.110 ;
        RECT 414.885 0.345 415.115 1.110 ;
        RECT 417.315 0.420 417.545 1.110 ;
        RECT 414.885 0.110 416.770 0.345 ;
        RECT 412.485 -1.080 412.810 -0.080 ;
        RECT 414.885 -1.710 415.115 0.110 ;
        RECT 415.345 -0.655 416.290 -0.130 ;
        RECT 416.540 -0.390 416.770 0.110 ;
        RECT 417.315 -0.070 418.440 0.420 ;
        RECT 415.345 -1.670 415.655 -0.655 ;
        RECT 416.540 -0.730 417.880 -0.390 ;
        RECT 418.120 -0.980 418.440 -0.070 ;
        RECT 419.365 -0.725 419.595 1.110 ;
        RECT 419.850 -0.320 421.115 -0.090 ;
        RECT 419.365 -0.955 420.640 -0.725 ;
        RECT 417.315 -1.215 418.440 -0.980 ;
        RECT 417.315 -1.710 417.545 -1.215 ;
        RECT 420.885 -1.750 421.115 -0.320 ;
        RECT 421.605 -0.725 421.835 1.110 ;
        RECT 422.090 -0.320 423.355 -0.090 ;
        RECT 421.605 -0.955 422.880 -0.725 ;
        RECT 423.125 -1.750 423.355 -0.320 ;
        RECT 423.845 -0.725 424.075 1.110 ;
        RECT 424.330 -0.320 425.595 -0.090 ;
        RECT 423.845 -0.955 425.120 -0.725 ;
        RECT 425.365 -1.750 425.595 -0.320 ;
        RECT 426.085 -0.725 426.315 1.110 ;
        RECT 426.570 -0.320 427.835 -0.090 ;
        RECT 426.085 -0.955 427.360 -0.725 ;
        RECT 427.605 -1.750 427.835 -0.320 ;
        RECT 428.325 -0.725 428.555 1.110 ;
        RECT 428.810 -0.320 430.075 -0.090 ;
        RECT 428.325 -0.955 429.600 -0.725 ;
        RECT 429.845 -1.750 430.075 -0.320 ;
        RECT 430.565 -0.725 430.795 1.110 ;
        RECT 431.050 -0.320 432.315 -0.090 ;
        RECT 430.565 -0.955 431.840 -0.725 ;
        RECT 432.085 -1.750 432.315 -0.320 ;
        RECT 434.945 -1.100 435.250 1.040 ;
        RECT 436.625 0.400 436.905 1.100 ;
        RECT 437.935 0.850 439.140 1.080 ;
        RECT 435.480 0.370 436.905 0.400 ;
        RECT 435.480 0.110 436.950 0.370 ;
        RECT 435.480 0.080 436.905 0.110 ;
        RECT 435.480 -1.680 435.835 0.080 ;
        RECT 436.065 -0.490 437.095 -0.150 ;
        RECT 436.065 -1.680 436.370 -0.490 ;
        RECT 438.260 -1.205 438.680 0.600 ;
        RECT 438.910 -0.770 439.140 0.850 ;
        RECT 439.380 -0.540 439.740 1.065 ;
        RECT 441.100 0.010 441.730 1.065 ;
        RECT 440.280 -0.770 441.135 -0.640 ;
        RECT 438.910 -1.000 441.135 -0.770 ;
        RECT 438.910 -1.750 439.305 -1.000 ;
        RECT 441.400 -1.240 441.730 0.010 ;
        RECT 440.965 -1.670 441.730 -1.240 ;
        RECT 442.210 -1.730 442.645 1.100 ;
        RECT 444.700 0.880 445.885 1.110 ;
        RECT 444.700 -0.370 444.930 0.880 ;
        RECT 445.655 0.770 445.885 0.880 ;
        RECT 446.695 0.880 448.910 1.110 ;
        RECT 446.695 0.770 446.925 0.880 ;
        RECT 445.160 0.125 445.390 0.650 ;
        RECT 445.655 0.540 446.925 0.770 ;
        RECT 445.160 -0.105 447.125 0.125 ;
        RECT 445.160 -0.600 445.390 -0.105 ;
        RECT 442.890 -0.830 445.390 -0.600 ;
        RECT 444.240 -1.490 444.470 -0.830 ;
        RECT 445.915 -1.260 446.460 -0.450 ;
        RECT 444.825 -1.620 446.460 -1.260 ;
        RECT 447.365 -1.150 447.705 0.650 ;
        RECT 448.000 -0.690 448.230 0.245 ;
        RECT 448.680 -0.230 448.910 0.880 ;
        RECT 450.040 0.565 450.680 0.795 ;
        RECT 448.680 -0.460 449.570 -0.230 ;
        RECT 448.000 -0.920 449.000 -0.690 ;
        RECT 447.365 -1.490 448.170 -1.150 ;
        RECT 448.770 -1.520 449.000 -0.920 ;
        RECT 449.230 -1.280 449.570 -0.460 ;
        RECT 450.450 -0.440 450.680 0.565 ;
        RECT 452.125 0.480 452.355 0.850 ;
        RECT 456.205 0.710 457.455 0.940 ;
        RECT 454.725 0.480 454.955 0.675 ;
        RECT 452.125 0.250 454.955 0.480 ;
        RECT 450.965 0.020 451.265 0.245 ;
        RECT 455.745 0.020 455.975 0.480 ;
        RECT 450.965 -0.210 455.975 0.020 ;
        RECT 450.450 -0.670 454.430 -0.440 ;
        RECT 449.965 -1.520 450.195 -0.690 ;
        RECT 450.790 -1.280 451.130 -0.670 ;
        RECT 454.845 -0.900 455.075 -0.690 ;
        RECT 451.890 -1.130 455.075 -0.900 ;
        RECT 451.890 -1.520 452.120 -1.130 ;
        RECT 455.425 -1.490 455.655 -0.210 ;
        RECT 456.205 -0.370 456.435 0.710 ;
        RECT 456.665 0.140 456.995 0.480 ;
        RECT 457.225 0.335 457.455 0.710 ;
        RECT 458.505 0.335 458.855 0.935 ;
        RECT 460.545 0.355 460.775 0.945 ;
        RECT 456.665 -1.205 456.895 0.140 ;
        RECT 457.225 0.105 458.855 0.335 ;
        RECT 457.200 -0.510 458.230 -0.130 ;
        RECT 458.625 -1.185 458.855 0.105 ;
        RECT 459.085 0.125 460.775 0.355 ;
        RECT 459.085 -0.770 459.315 0.125 ;
        RECT 459.550 -0.510 460.840 -0.130 ;
        RECT 459.085 -1.000 460.875 -0.770 ;
        RECT 456.490 -1.435 456.895 -1.205 ;
        RECT 458.350 -1.415 458.855 -1.185 ;
        RECT 460.645 -1.470 460.875 -1.000 ;
        RECT 448.770 -1.750 452.120 -1.520 ;
        RECT 223.320 -3.190 232.945 -2.810 ;
        RECT 305.150 -3.040 308.080 -2.810 ;
        RECT 223.320 -3.300 224.520 -3.190 ;
        RECT 297.285 -3.560 297.515 -3.090 ;
        RECT 299.425 -3.430 299.755 -3.090 ;
        RECT 297.285 -3.790 299.130 -3.560 ;
        RECT 297.320 -4.410 298.630 -4.045 ;
        RECT 298.900 -4.640 299.130 -3.790 ;
        RECT 286.700 -5.160 289.200 -4.860 ;
        RECT 230.490 -5.635 231.390 -5.485 ;
        RECT 234.005 -5.635 234.905 -5.485 ;
        RECT 236.240 -5.560 289.200 -5.160 ;
        RECT 297.385 -4.875 299.130 -4.640 ;
        RECT 299.425 -4.660 299.660 -3.430 ;
        RECT 299.930 -4.430 301.070 -4.050 ;
        RECT 297.385 -5.505 297.615 -4.875 ;
        RECT 299.425 -4.895 301.080 -4.660 ;
        RECT 299.425 -5.505 299.655 -4.895 ;
        RECT 300.850 -5.440 301.080 -4.895 ;
        RECT 301.310 -5.210 301.650 -3.070 ;
        RECT 302.385 -4.045 302.715 -3.070 ;
        RECT 305.150 -3.585 305.380 -3.040 ;
        RECT 303.040 -3.815 305.380 -3.585 ;
        RECT 301.925 -5.440 302.155 -4.210 ;
        RECT 302.385 -4.275 305.275 -4.045 ;
        RECT 302.385 -5.265 302.615 -4.275 ;
        RECT 306.915 -4.360 307.255 -3.270 ;
        RECT 307.850 -3.895 308.080 -3.040 ;
        RECT 308.970 -3.040 313.150 -2.810 ;
        RECT 316.340 -2.930 316.855 -2.830 ;
        RECT 308.970 -3.070 309.200 -3.040 ;
        RECT 308.310 -3.410 309.200 -3.070 ;
        RECT 306.075 -4.505 308.685 -4.360 ;
        RECT 303.155 -5.265 303.495 -4.520 ;
        RECT 304.055 -4.590 308.685 -4.505 ;
        RECT 304.055 -4.735 306.415 -4.590 ;
        RECT 306.075 -5.210 306.415 -4.735 ;
        RECT 306.725 -5.055 308.115 -4.820 ;
        RECT 229.940 -5.865 231.940 -5.635 ;
        RECT 233.455 -5.865 235.455 -5.635 ;
        RECT 230.275 -7.435 230.655 -6.535 ;
        RECT 231.225 -7.435 231.455 -5.865 ;
        RECT 233.790 -7.435 234.170 -6.535 ;
        RECT 234.740 -7.435 234.970 -5.865 ;
        RECT 229.895 -8.830 230.275 -8.550 ;
        RECT 191.600 -9.170 230.275 -8.830 ;
        RECT 229.895 -9.450 230.275 -9.170 ;
        RECT 230.770 -8.830 231.110 -7.665 ;
        RECT 233.410 -8.830 233.790 -8.550 ;
        RECT 230.770 -9.170 233.790 -8.830 ;
        RECT 183.905 -10.685 184.805 -10.305 ;
        RECT 230.770 -10.335 231.110 -9.170 ;
        RECT 233.410 -9.450 233.790 -9.170 ;
        RECT 234.285 -8.830 234.625 -7.665 ;
        RECT 236.240 -8.830 236.540 -5.560 ;
        RECT 286.700 -5.860 289.200 -5.560 ;
        RECT 300.850 -5.670 302.155 -5.440 ;
        RECT 303.155 -5.440 305.540 -5.265 ;
        RECT 306.725 -5.440 306.955 -5.055 ;
        RECT 303.155 -5.495 306.955 -5.440 ;
        RECT 305.310 -5.670 306.955 -5.495 ;
        RECT 307.885 -5.345 308.115 -5.055 ;
        RECT 308.345 -5.060 308.685 -4.590 ;
        RECT 308.970 -4.830 309.200 -3.410 ;
        RECT 309.595 -3.500 311.535 -3.270 ;
        RECT 310.670 -4.820 310.900 -3.500 ;
        RECT 312.920 -3.675 313.150 -3.040 ;
        RECT 312.920 -3.910 314.375 -3.675 ;
        RECT 314.770 -3.780 315.000 -3.085 ;
        RECT 316.230 -3.310 316.855 -2.930 ;
        RECT 316.340 -3.440 316.855 -3.310 ;
        RECT 311.130 -4.430 312.325 -4.050 ;
        RECT 314.770 -4.120 316.160 -3.780 ;
        RECT 314.770 -4.140 315.000 -4.120 ;
        RECT 312.795 -4.385 315.000 -4.140 ;
        RECT 308.970 -5.060 309.935 -4.830 ;
        RECT 310.670 -5.055 312.640 -4.820 ;
        RECT 310.670 -5.125 310.900 -5.055 ;
        RECT 312.410 -5.165 312.640 -5.055 ;
        RECT 307.885 -5.575 309.355 -5.345 ;
        RECT 314.770 -5.660 315.000 -4.385 ;
        RECT 316.465 -4.470 316.855 -3.440 ;
        RECT 316.085 -5.660 316.855 -4.470 ;
        RECT 317.320 -4.350 317.710 -2.810 ;
        RECT 318.395 -3.720 318.760 -2.835 ;
        RECT 317.945 -4.100 318.760 -3.720 ;
        RECT 317.320 -4.580 318.730 -4.350 ;
        RECT 319.000 -4.470 319.365 -3.340 ;
        RECT 318.500 -5.660 318.730 -4.580 ;
        RECT 320.245 -4.740 320.475 -2.830 ;
        RECT 320.705 -4.510 321.000 -2.830 ;
        RECT 320.245 -4.970 320.985 -4.740 ;
        RECT 320.755 -5.440 320.985 -4.970 ;
        RECT 321.230 -4.870 321.595 -2.830 ;
        RECT 321.825 -4.600 322.160 -2.830 ;
        RECT 322.485 -4.410 322.715 -2.830 ;
        RECT 322.945 -3.880 323.280 -2.830 ;
        RECT 322.945 -4.180 324.350 -3.880 ;
        RECT 322.485 -4.640 323.075 -4.410 ;
        RECT 323.375 -4.430 324.350 -4.180 ;
        RECT 324.600 -4.350 324.990 -2.810 ;
        RECT 325.675 -3.720 326.040 -2.835 ;
        RECT 328.550 -3.090 328.810 -2.930 ;
        RECT 325.225 -4.100 326.040 -3.720 ;
        RECT 324.600 -4.580 326.010 -4.350 ;
        RECT 326.280 -4.470 326.645 -3.340 ;
        RECT 321.230 -5.210 322.615 -4.870 ;
        RECT 322.845 -5.440 323.075 -4.640 ;
        RECT 320.755 -5.670 323.075 -5.440 ;
        RECT 325.780 -5.660 326.010 -4.580 ;
        RECT 328.540 -4.990 328.875 -3.090 ;
        RECT 330.780 -4.990 331.115 -3.090 ;
        RECT 332.005 -3.835 333.280 -3.605 ;
        RECT 332.005 -5.670 332.235 -3.835 ;
        RECT 333.525 -4.240 333.755 -2.810 ;
        RECT 332.490 -4.470 333.755 -4.240 ;
        RECT 336.670 -3.885 337.260 -2.845 ;
        RECT 336.670 -5.600 337.035 -3.885 ;
        RECT 338.520 -4.020 338.895 -3.315 ;
        RECT 337.330 -4.800 337.670 -4.160 ;
        RECT 338.010 -4.430 338.895 -4.020 ;
        RECT 339.125 -4.800 339.355 -2.845 ;
        RECT 337.330 -5.035 339.355 -4.800 ;
        RECT 339.025 -5.660 339.355 -5.035 ;
        RECT 339.845 -3.835 341.120 -3.605 ;
        RECT 339.845 -5.670 340.075 -3.835 ;
        RECT 341.365 -4.240 341.595 -2.810 ;
        RECT 340.330 -4.470 341.595 -4.240 ;
        RECT 342.085 -3.835 343.360 -3.605 ;
        RECT 342.085 -5.670 342.315 -3.835 ;
        RECT 343.605 -4.240 343.835 -2.810 ;
        RECT 344.830 -3.085 348.055 -2.855 ;
        RECT 344.830 -3.315 345.170 -3.085 ;
        RECT 345.890 -4.050 346.210 -3.400 ;
        RECT 342.570 -4.470 343.835 -4.240 ;
        RECT 345.180 -4.430 346.210 -4.050 ;
        RECT 346.440 -4.695 346.760 -3.400 ;
        RECT 347.000 -4.695 347.550 -3.400 ;
        RECT 347.825 -3.740 348.055 -3.085 ;
        RECT 347.825 -4.080 348.955 -3.740 ;
        RECT 347.825 -5.105 348.055 -4.080 ;
        RECT 344.830 -5.335 348.055 -5.105 ;
        RECT 344.830 -5.620 345.170 -5.335 ;
        RECT 346.870 -5.620 347.210 -5.335 ;
        RECT 349.210 -5.660 349.650 -2.930 ;
        RECT 350.885 -5.650 351.220 -2.880 ;
        RECT 351.450 -5.230 351.775 -3.250 ;
        RECT 352.725 -3.835 354.000 -3.605 ;
        RECT 352.725 -5.670 352.955 -3.835 ;
        RECT 354.245 -4.240 354.475 -2.810 ;
        RECT 353.210 -4.470 354.475 -4.240 ;
        RECT 354.965 -3.835 356.240 -3.605 ;
        RECT 354.965 -5.670 355.195 -3.835 ;
        RECT 356.485 -4.240 356.715 -2.810 ;
        RECT 355.450 -4.470 356.715 -4.240 ;
        RECT 357.205 -3.835 358.480 -3.605 ;
        RECT 357.205 -5.670 357.435 -3.835 ;
        RECT 358.725 -4.240 358.955 -2.810 ;
        RECT 362.150 -2.975 362.410 -2.930 ;
        RECT 362.150 -3.310 362.530 -2.975 ;
        RECT 362.190 -3.330 362.530 -3.310 ;
        RECT 364.430 -3.330 364.770 -2.975 ;
        RECT 362.190 -3.565 364.770 -3.330 ;
        RECT 357.690 -4.470 358.955 -4.240 ;
        RECT 361.370 -4.470 362.440 -4.040 ;
        RECT 362.100 -5.670 362.440 -4.470 ;
        RECT 362.670 -5.670 363.010 -3.855 ;
        RECT 363.790 -5.670 364.130 -3.855 ;
        RECT 364.370 -5.670 364.770 -3.565 ;
        RECT 365.605 -3.835 366.880 -3.605 ;
        RECT 365.605 -5.670 365.835 -3.835 ;
        RECT 367.125 -4.240 367.355 -2.810 ;
        RECT 369.390 -4.070 369.695 -2.880 ;
        RECT 366.090 -4.470 367.355 -4.240 ;
        RECT 368.665 -4.410 369.695 -4.070 ;
        RECT 369.925 -4.640 370.280 -2.880 ;
        RECT 368.855 -4.960 370.280 -4.640 ;
        RECT 368.855 -5.660 369.135 -4.960 ;
        RECT 370.510 -5.600 370.815 -3.460 ;
        RECT 371.765 -3.835 373.040 -3.605 ;
        RECT 371.765 -5.670 371.995 -3.835 ;
        RECT 373.285 -4.240 373.515 -2.810 ;
        RECT 372.250 -4.470 373.515 -4.240 ;
        RECT 375.685 -3.835 376.960 -3.605 ;
        RECT 375.685 -5.670 375.915 -3.835 ;
        RECT 377.205 -4.240 377.435 -2.810 ;
        RECT 376.170 -4.470 377.435 -4.240 ;
        RECT 377.925 -3.835 379.200 -3.605 ;
        RECT 377.925 -5.670 378.155 -3.835 ;
        RECT 379.445 -4.240 379.675 -2.810 ;
        RECT 378.410 -4.470 379.675 -4.240 ;
        RECT 382.305 -5.600 382.610 -3.460 ;
        RECT 382.840 -4.640 383.195 -2.880 ;
        RECT 383.425 -4.070 383.730 -2.880 ;
        RECT 386.215 -3.225 386.610 -2.810 ;
        RECT 387.960 -3.040 389.400 -2.810 ;
        RECT 387.960 -3.225 388.190 -3.040 ;
        RECT 386.215 -3.460 388.190 -3.225 ;
        RECT 389.170 -3.225 389.400 -3.040 ;
        RECT 390.200 -3.040 391.640 -2.810 ;
        RECT 390.200 -3.225 390.430 -3.040 ;
        RECT 388.430 -3.690 388.870 -3.290 ;
        RECT 389.170 -3.460 390.430 -3.225 ;
        RECT 391.410 -3.225 391.640 -3.040 ;
        RECT 392.910 -3.225 393.780 -2.810 ;
        RECT 394.680 -3.225 396.120 -2.810 ;
        RECT 397.420 -3.225 397.810 -2.810 ;
        RECT 390.660 -3.690 391.110 -3.290 ;
        RECT 391.410 -3.460 397.810 -3.225 ;
        RECT 386.750 -3.920 392.695 -3.690 ;
        RECT 394.510 -3.920 397.140 -3.690 ;
        RECT 383.425 -4.410 384.455 -4.070 ;
        RECT 385.365 -4.150 386.530 -4.030 ;
        RECT 392.930 -4.150 393.990 -4.030 ;
        RECT 385.365 -4.430 393.990 -4.150 ;
        RECT 382.840 -4.960 384.265 -4.640 ;
        RECT 383.985 -5.660 384.265 -4.960 ;
        RECT 385.205 -5.080 393.180 -4.850 ;
        RECT 385.205 -5.660 385.435 -5.080 ;
        RECT 389.585 -5.660 389.815 -5.080 ;
        RECT 392.950 -5.440 393.180 -5.080 ;
        RECT 394.510 -5.130 394.920 -3.920 ;
        RECT 397.380 -4.155 397.810 -3.460 ;
        RECT 400.785 -3.040 404.300 -2.810 ;
        RECT 400.785 -3.545 401.055 -3.040 ;
        RECT 404.350 -3.270 406.725 -3.265 ;
        RECT 395.150 -4.390 397.810 -4.155 ;
        RECT 395.150 -5.190 395.515 -4.390 ;
        RECT 396.305 -5.440 396.535 -4.810 ;
        RECT 397.420 -5.190 397.810 -4.390 ;
        RECT 399.665 -3.815 401.055 -3.545 ;
        RECT 401.290 -3.490 406.725 -3.270 ;
        RECT 401.290 -3.495 407.870 -3.490 ;
        RECT 401.290 -3.500 404.400 -3.495 ;
        RECT 399.665 -4.805 399.985 -3.815 ;
        RECT 401.290 -3.835 401.670 -3.500 ;
        RECT 402.330 -3.975 402.980 -3.745 ;
        RECT 404.450 -3.955 406.130 -3.725 ;
        RECT 406.385 -3.870 407.870 -3.495 ;
        RECT 402.705 -4.030 402.980 -3.975 ;
        RECT 400.290 -4.540 402.100 -4.105 ;
        RECT 402.705 -4.185 404.025 -4.030 ;
        RECT 405.900 -4.100 406.130 -3.955 ;
        RECT 402.705 -4.415 405.670 -4.185 ;
        RECT 405.900 -4.380 407.870 -4.100 ;
        RECT 401.820 -4.645 402.100 -4.540 ;
        RECT 406.635 -4.645 407.790 -4.620 ;
        RECT 398.545 -5.440 398.775 -4.810 ;
        RECT 392.950 -5.670 398.775 -5.440 ;
        RECT 399.665 -5.040 401.570 -4.805 ;
        RECT 401.820 -4.875 407.790 -4.645 ;
        RECT 408.725 -4.670 408.955 -2.850 ;
        RECT 409.185 -3.905 409.495 -2.890 ;
        RECT 411.155 -3.345 411.385 -2.850 ;
        RECT 417.560 -3.040 420.800 -2.810 ;
        RECT 417.560 -3.145 417.790 -3.040 ;
        RECT 411.155 -3.580 412.280 -3.345 ;
        RECT 414.920 -3.375 417.790 -3.145 ;
        RECT 420.570 -3.145 420.800 -3.040 ;
        RECT 422.235 -3.040 432.940 -2.810 ;
        RECT 422.235 -3.145 422.465 -3.040 ;
        RECT 420.570 -3.375 422.465 -3.145 ;
        RECT 423.160 -3.500 431.600 -3.270 ;
        RECT 409.185 -4.430 410.130 -3.905 ;
        RECT 410.380 -4.170 411.720 -3.830 ;
        RECT 410.380 -4.670 410.610 -4.170 ;
        RECT 411.960 -4.490 412.280 -3.580 ;
        RECT 418.040 -3.605 420.190 -3.500 ;
        RECT 415.360 -3.835 422.920 -3.605 ;
        RECT 416.280 -4.400 422.370 -4.080 ;
        RECT 399.665 -5.670 400.075 -5.040 ;
        RECT 401.340 -5.105 401.570 -5.040 ;
        RECT 408.725 -4.905 410.610 -4.670 ;
        RECT 401.340 -5.335 408.300 -5.105 ;
        RECT 401.340 -5.590 402.425 -5.335 ;
        RECT 403.580 -5.590 404.545 -5.335 ;
        RECT 405.460 -5.590 406.670 -5.335 ;
        RECT 407.500 -5.590 408.300 -5.335 ;
        RECT 408.725 -5.670 408.955 -4.905 ;
        RECT 411.155 -4.980 412.280 -4.490 ;
        RECT 422.600 -4.705 422.920 -3.835 ;
        RECT 411.155 -5.670 411.385 -4.980 ;
        RECT 423.160 -5.075 423.480 -3.500 ;
        RECT 426.330 -3.960 431.160 -3.730 ;
        RECT 435.205 -3.880 435.830 -2.855 ;
        RECT 426.330 -4.050 426.580 -3.960 ;
        RECT 423.710 -4.400 424.580 -4.050 ;
        RECT 424.810 -4.400 426.580 -4.050 ;
        RECT 423.750 -4.430 424.010 -4.400 ;
        RECT 424.240 -4.640 424.580 -4.400 ;
        RECT 426.915 -4.420 432.500 -4.190 ;
        RECT 426.915 -4.640 427.165 -4.420 ;
        RECT 424.240 -4.960 427.165 -4.640 ;
        RECT 415.670 -5.200 424.030 -5.075 ;
        RECT 427.395 -5.200 428.730 -5.075 ;
        RECT 430.130 -5.200 430.470 -4.755 ;
        RECT 415.670 -5.305 430.470 -5.200 ;
        RECT 415.670 -5.335 422.945 -5.305 ;
        RECT 415.670 -5.520 416.720 -5.335 ;
        RECT 417.560 -5.520 418.760 -5.335 ;
        RECT 419.600 -5.520 420.800 -5.335 ;
        RECT 421.640 -5.520 422.945 -5.335 ;
        RECT 423.780 -5.520 427.645 -5.305 ;
        RECT 428.480 -5.520 430.470 -5.305 ;
        RECT 417.590 -5.550 417.850 -5.520 ;
        RECT 430.130 -5.605 430.470 -5.520 ;
        RECT 435.205 -5.660 435.675 -3.880 ;
        RECT 436.940 -3.910 437.455 -2.930 ;
        RECT 435.905 -4.860 436.190 -4.110 ;
        RECT 436.570 -4.470 437.455 -3.910 ;
        RECT 437.685 -4.860 437.915 -3.080 ;
        RECT 439.525 -3.295 439.755 -2.955 ;
        RECT 441.765 -3.295 441.995 -2.955 ;
        RECT 439.525 -3.530 442.475 -3.295 ;
        RECT 442.140 -3.965 442.475 -3.530 ;
        RECT 454.085 -3.835 455.360 -3.605 ;
        RECT 438.810 -4.430 441.670 -3.995 ;
        RECT 442.140 -4.305 446.430 -3.965 ;
        RECT 442.140 -4.810 442.475 -4.305 ;
        RECT 448.500 -4.310 451.700 -3.965 ;
        RECT 435.905 -5.095 437.915 -4.860 ;
        RECT 437.530 -5.670 437.915 -5.095 ;
        RECT 439.425 -5.040 442.475 -4.810 ;
        RECT 439.425 -5.660 439.655 -5.040 ;
        RECT 441.665 -5.660 441.895 -5.040 ;
        RECT 454.085 -5.670 454.315 -3.835 ;
        RECT 455.605 -4.240 455.835 -2.810 ;
        RECT 454.570 -4.470 455.835 -4.240 ;
        RECT 456.885 -4.870 457.115 -3.085 ;
        RECT 457.345 -4.020 457.720 -2.830 ;
        RECT 459.305 -3.560 459.535 -3.080 ;
        RECT 459.305 -3.790 460.450 -3.560 ;
        RECT 457.345 -4.430 458.290 -4.020 ;
        RECT 458.530 -4.320 459.850 -4.020 ;
        RECT 458.530 -4.870 458.855 -4.320 ;
        RECT 460.110 -4.640 460.450 -3.790 ;
        RECT 456.885 -5.100 458.855 -4.870 ;
        RECT 459.305 -4.990 460.450 -4.640 ;
        RECT 456.885 -5.670 457.115 -5.100 ;
        RECT 459.305 -5.670 459.535 -4.990 ;
        RECT 298.905 -6.850 299.135 -6.740 ;
        RECT 298.870 -7.230 299.135 -6.850 ;
        RECT 298.905 -7.410 299.135 -7.230 ;
        RECT 301.145 -7.410 301.375 -6.740 ;
        RECT 303.385 -7.410 303.615 -6.740 ;
        RECT 305.525 -7.410 305.755 -6.740 ;
        RECT 307.865 -7.360 308.095 -6.740 ;
        RECT 310.105 -7.360 310.335 -6.740 ;
        RECT 298.905 -7.790 305.755 -7.410 ;
        RECT 307.285 -7.590 310.335 -7.360 ;
        RECT 298.060 -8.435 301.260 -8.090 ;
        RECT 301.960 -8.700 302.760 -7.790 ;
        RECT 307.285 -8.095 307.620 -7.590 ;
        RECT 303.330 -8.435 307.620 -8.095 ;
        RECT 308.090 -8.405 310.950 -7.970 ;
        RECT 234.285 -9.170 236.540 -8.830 ;
        RECT 298.805 -9.080 305.755 -8.700 ;
        RECT 234.285 -10.335 234.625 -9.170 ;
        RECT 298.805 -9.445 299.035 -9.080 ;
        RECT 301.045 -9.445 301.275 -9.080 ;
        RECT 303.285 -9.445 303.515 -9.080 ;
        RECT 305.495 -9.445 305.755 -9.080 ;
        RECT 307.285 -8.870 307.620 -8.435 ;
        RECT 311.845 -8.565 312.075 -6.730 ;
        RECT 312.330 -8.160 313.595 -7.930 ;
        RECT 311.845 -8.795 313.120 -8.565 ;
        RECT 307.285 -9.105 310.235 -8.870 ;
        RECT 307.765 -9.445 307.995 -9.105 ;
        RECT 310.005 -9.445 310.235 -9.105 ;
        RECT 313.365 -9.590 313.595 -8.160 ;
        RECT 316.885 -8.565 317.115 -6.730 ;
        RECT 320.905 -7.485 321.135 -6.895 ;
        RECT 320.905 -7.715 322.595 -7.485 ;
        RECT 317.370 -8.160 318.635 -7.930 ;
        RECT 316.885 -8.795 318.160 -8.565 ;
        RECT 318.405 -9.590 318.635 -8.160 ;
        RECT 320.840 -8.350 322.130 -7.970 ;
        RECT 322.365 -8.610 322.595 -7.715 ;
        RECT 320.805 -8.840 322.595 -8.610 ;
        RECT 322.825 -7.505 323.175 -6.905 ;
        RECT 324.225 -7.130 325.475 -6.900 ;
        RECT 332.770 -6.960 334.985 -6.730 ;
        RECT 324.225 -7.505 324.455 -7.130 ;
        RECT 322.825 -7.735 324.455 -7.505 ;
        RECT 324.685 -7.700 325.015 -7.360 ;
        RECT 320.805 -9.310 321.035 -8.840 ;
        RECT 322.825 -9.025 323.055 -7.735 ;
        RECT 323.450 -8.350 324.480 -7.970 ;
        RECT 322.825 -9.255 323.330 -9.025 ;
        RECT 324.785 -9.045 325.015 -7.700 ;
        RECT 325.245 -8.210 325.475 -7.130 ;
        RECT 326.725 -7.360 326.955 -7.165 ;
        RECT 329.325 -7.360 329.555 -6.990 ;
        RECT 325.705 -7.820 325.935 -7.360 ;
        RECT 326.725 -7.590 329.555 -7.360 ;
        RECT 331.000 -7.275 331.640 -7.045 ;
        RECT 330.415 -7.820 330.715 -7.595 ;
        RECT 325.705 -8.050 330.715 -7.820 ;
        RECT 324.785 -9.275 325.190 -9.045 ;
        RECT 326.025 -9.330 326.255 -8.050 ;
        RECT 331.000 -8.280 331.230 -7.275 ;
        RECT 332.770 -8.070 333.000 -6.960 ;
        RECT 334.755 -7.070 334.985 -6.960 ;
        RECT 335.795 -6.960 336.980 -6.730 ;
        RECT 335.795 -7.070 336.025 -6.960 ;
        RECT 327.250 -8.510 331.230 -8.280 ;
        RECT 332.110 -8.300 333.000 -8.070 ;
        RECT 326.605 -8.740 326.835 -8.530 ;
        RECT 326.605 -8.970 329.790 -8.740 ;
        RECT 329.560 -9.360 329.790 -8.970 ;
        RECT 330.550 -9.120 330.890 -8.510 ;
        RECT 331.485 -9.360 331.715 -8.530 ;
        RECT 332.110 -9.120 332.450 -8.300 ;
        RECT 333.450 -8.530 333.680 -7.595 ;
        RECT 332.680 -8.760 333.680 -8.530 ;
        RECT 332.680 -9.360 332.910 -8.760 ;
        RECT 333.975 -8.990 334.315 -7.190 ;
        RECT 334.755 -7.300 336.025 -7.070 ;
        RECT 336.290 -7.715 336.520 -7.190 ;
        RECT 334.555 -7.945 336.520 -7.715 ;
        RECT 333.510 -9.330 334.315 -8.990 ;
        RECT 335.220 -9.100 335.765 -8.290 ;
        RECT 336.290 -8.440 336.520 -7.945 ;
        RECT 336.750 -8.210 336.980 -6.960 ;
        RECT 336.290 -8.670 338.790 -8.440 ;
        RECT 329.560 -9.590 332.910 -9.360 ;
        RECT 335.220 -9.460 336.855 -9.100 ;
        RECT 337.210 -9.330 337.440 -8.670 ;
        RECT 339.035 -9.570 339.470 -6.740 ;
        RECT 339.845 -8.565 340.075 -6.730 ;
        RECT 340.330 -8.160 341.595 -7.930 ;
        RECT 339.845 -8.795 341.120 -8.565 ;
        RECT 341.365 -9.590 341.595 -8.160 ;
        RECT 342.085 -8.565 342.315 -6.730 ;
        RECT 342.570 -8.160 343.835 -7.930 ;
        RECT 342.085 -8.795 343.360 -8.565 ;
        RECT 343.605 -9.590 343.835 -8.160 ;
        RECT 344.325 -8.565 344.555 -6.730 ;
        RECT 344.810 -8.160 346.075 -7.930 ;
        RECT 344.325 -8.795 345.600 -8.565 ;
        RECT 345.845 -9.590 346.075 -8.160 ;
        RECT 346.565 -8.565 346.795 -6.730 ;
        RECT 347.050 -8.160 348.315 -7.930 ;
        RECT 346.565 -8.795 347.840 -8.565 ;
        RECT 348.085 -9.590 348.315 -8.160 ;
        RECT 348.805 -8.565 349.035 -6.730 ;
        RECT 349.290 -8.160 350.555 -7.930 ;
        RECT 348.805 -8.795 350.080 -8.565 ;
        RECT 350.325 -9.590 350.555 -8.160 ;
        RECT 351.045 -8.565 351.275 -6.730 ;
        RECT 351.530 -8.160 352.795 -7.930 ;
        RECT 351.045 -8.795 352.320 -8.565 ;
        RECT 352.565 -9.590 352.795 -8.160 ;
        RECT 356.085 -8.565 356.315 -6.730 ;
        RECT 356.570 -8.160 357.835 -7.930 ;
        RECT 356.085 -8.795 357.360 -8.565 ;
        RECT 357.605 -9.590 357.835 -8.160 ;
        RECT 358.325 -8.565 358.555 -6.730 ;
        RECT 361.575 -7.440 361.855 -6.740 ;
        RECT 361.575 -7.760 363.000 -7.440 ;
        RECT 358.810 -8.160 360.075 -7.930 ;
        RECT 358.325 -8.795 359.600 -8.565 ;
        RECT 359.845 -9.590 360.075 -8.160 ;
        RECT 361.385 -8.330 362.415 -7.990 ;
        RECT 362.110 -9.520 362.415 -8.330 ;
        RECT 362.645 -9.520 363.000 -7.760 ;
        RECT 363.230 -8.940 363.535 -6.800 ;
        RECT 364.645 -7.065 364.875 -6.740 ;
        RECT 374.990 -6.960 383.540 -6.730 ;
        RECT 374.990 -7.065 375.330 -6.960 ;
        RECT 364.645 -7.295 375.330 -7.065 ;
        RECT 364.645 -7.590 364.875 -7.295 ;
        RECT 365.600 -7.760 374.060 -7.525 ;
        RECT 374.990 -7.590 375.330 -7.295 ;
        RECT 384.965 -7.065 385.195 -6.730 ;
        RECT 387.780 -6.960 393.675 -6.730 ;
        RECT 387.780 -7.065 388.010 -6.960 ;
        RECT 384.965 -7.295 388.010 -7.065 ;
        RECT 376.060 -7.760 383.420 -7.440 ;
        RECT 384.965 -7.620 385.195 -7.295 ;
        RECT 388.255 -7.525 389.320 -7.410 ;
        RECT 365.600 -8.000 365.830 -7.760 ;
        RECT 364.810 -8.320 365.830 -8.000 ;
        RECT 366.150 -8.385 368.320 -7.990 ;
        RECT 368.855 -8.155 369.195 -7.760 ;
        RECT 370.530 -8.155 370.870 -7.760 ;
        RECT 373.830 -8.000 374.060 -7.760 ;
        RECT 373.830 -8.320 374.850 -8.000 ;
        RECT 375.365 -8.320 382.960 -8.000 ;
        RECT 366.150 -8.615 373.560 -8.385 ;
        RECT 376.465 -8.780 382.690 -8.550 ;
        RECT 365.660 -9.020 375.895 -8.845 ;
        RECT 380.570 -8.910 382.690 -8.780 ;
        RECT 383.190 -8.935 383.420 -7.760 ;
        RECT 385.490 -7.760 389.320 -7.525 ;
        RECT 385.490 -8.000 386.035 -7.760 ;
        RECT 384.895 -8.320 386.035 -8.000 ;
        RECT 386.525 -8.320 388.270 -8.000 ;
        RECT 388.700 -8.320 389.320 -7.760 ;
        RECT 389.560 -7.760 392.750 -7.340 ;
        RECT 393.445 -7.620 393.675 -6.960 ;
        RECT 398.150 -7.360 398.380 -6.740 ;
        RECT 399.640 -7.025 404.720 -6.795 ;
        RECT 399.640 -7.360 399.875 -7.025 ;
        RECT 389.560 -8.560 389.880 -7.760 ;
        RECT 390.150 -8.320 393.500 -8.000 ;
        RECT 365.660 -9.075 379.920 -9.020 ;
        RECT 365.660 -9.345 366.000 -9.075 ;
        RECT 368.340 -9.345 368.680 -9.075 ;
        RECT 371.020 -9.345 371.360 -9.075 ;
        RECT 373.700 -9.345 374.040 -9.075 ;
        RECT 375.665 -9.190 379.920 -9.075 ;
        RECT 382.980 -9.165 383.420 -8.935 ;
        RECT 388.775 -8.880 390.265 -8.560 ;
        RECT 390.610 -8.880 392.760 -8.560 ;
        RECT 388.775 -9.020 389.005 -8.880 ;
        RECT 382.980 -9.190 383.210 -9.165 ;
        RECT 375.665 -9.250 383.210 -9.190 ;
        RECT 377.080 -9.410 377.590 -9.250 ;
        RECT 377.080 -9.545 377.420 -9.410 ;
        RECT 379.690 -9.420 383.210 -9.250 ;
        RECT 385.930 -9.250 389.005 -9.020 ;
        RECT 390.005 -9.120 390.265 -8.880 ;
        RECT 381.160 -9.590 381.500 -9.420 ;
        RECT 385.930 -9.560 386.270 -9.250 ;
        RECT 388.170 -9.560 388.510 -9.250 ;
        RECT 390.005 -9.440 391.770 -9.120 ;
        RECT 396.300 -9.310 396.635 -7.410 ;
        RECT 398.150 -7.590 399.875 -7.360 ;
        RECT 400.490 -7.470 403.795 -7.420 ;
        RECT 400.490 -7.730 403.910 -7.470 ;
        RECT 404.490 -7.685 404.720 -7.025 ;
        RECT 406.625 -7.440 406.855 -6.740 ;
        RECT 408.580 -7.440 408.940 -6.740 ;
        RECT 400.490 -7.760 403.795 -7.730 ;
        RECT 405.670 -7.760 408.940 -7.440 ;
        RECT 411.525 -7.300 411.755 -6.730 ;
        RECT 411.525 -7.530 413.495 -7.300 ;
        RECT 398.420 -8.320 400.120 -7.995 ;
        RECT 400.490 -9.020 400.810 -7.760 ;
        RECT 401.130 -8.320 404.565 -8.000 ;
        RECT 401.130 -8.720 401.470 -8.320 ;
        RECT 401.840 -8.880 404.565 -8.560 ;
        RECT 405.670 -8.585 405.900 -7.760 ;
        RECT 406.130 -8.320 409.540 -8.000 ;
        RECT 405.670 -8.855 406.700 -8.585 ;
        RECT 398.810 -9.250 401.165 -9.020 ;
        RECT 406.340 -9.120 406.700 -8.855 ;
        RECT 407.000 -8.880 409.540 -8.560 ;
        RECT 406.340 -9.150 408.010 -9.120 ;
        RECT 396.310 -9.470 396.570 -9.310 ;
        RECT 398.810 -9.560 400.085 -9.250 ;
        RECT 400.935 -9.315 401.165 -9.250 ;
        RECT 400.935 -9.545 402.815 -9.315 ;
        RECT 406.330 -9.410 408.010 -9.150 ;
        RECT 411.525 -9.315 411.755 -7.530 ;
        RECT 411.985 -8.380 412.930 -7.970 ;
        RECT 413.170 -8.080 413.495 -7.530 ;
        RECT 413.945 -7.410 414.175 -6.730 ;
        RECT 413.945 -7.760 415.090 -7.410 ;
        RECT 413.170 -8.380 414.490 -8.080 ;
        RECT 406.340 -9.440 408.010 -9.410 ;
        RECT 411.985 -9.570 412.360 -8.380 ;
        RECT 414.750 -8.610 415.090 -7.760 ;
        RECT 413.945 -8.840 415.090 -8.610 ;
        RECT 416.005 -8.565 416.235 -6.730 ;
        RECT 419.830 -7.420 420.090 -7.410 ;
        RECT 420.695 -7.420 420.925 -6.730 ;
        RECT 419.800 -7.910 420.925 -7.420 ;
        RECT 423.125 -7.495 423.355 -6.730 ;
        RECT 425.185 -7.410 425.415 -6.730 ;
        RECT 427.605 -7.300 427.835 -6.730 ;
        RECT 421.470 -7.730 423.355 -7.495 ;
        RECT 416.490 -8.160 417.755 -7.930 ;
        RECT 416.005 -8.795 417.280 -8.565 ;
        RECT 413.945 -9.320 414.175 -8.840 ;
        RECT 417.525 -9.590 417.755 -8.160 ;
        RECT 419.800 -8.820 420.120 -7.910 ;
        RECT 421.470 -8.230 421.700 -7.730 ;
        RECT 420.360 -8.570 421.700 -8.230 ;
        RECT 421.950 -8.495 422.895 -7.970 ;
        RECT 419.800 -9.055 420.925 -8.820 ;
        RECT 420.695 -9.550 420.925 -9.055 ;
        RECT 422.585 -9.510 422.895 -8.495 ;
        RECT 423.125 -9.550 423.355 -7.730 ;
        RECT 424.270 -7.760 425.415 -7.410 ;
        RECT 425.865 -7.530 427.835 -7.300 ;
        RECT 424.270 -8.610 424.610 -7.760 ;
        RECT 425.865 -8.080 426.190 -7.530 ;
        RECT 424.870 -8.380 426.190 -8.080 ;
        RECT 426.430 -8.380 427.375 -7.970 ;
        RECT 424.270 -8.840 425.415 -8.610 ;
        RECT 425.185 -9.320 425.415 -8.840 ;
        RECT 427.000 -9.570 427.375 -8.380 ;
        RECT 427.605 -9.315 427.835 -7.530 ;
        RECT 428.325 -7.365 428.655 -6.740 ;
        RECT 428.325 -7.600 430.350 -7.365 ;
        RECT 428.325 -9.555 428.555 -7.600 ;
        RECT 428.785 -8.380 429.670 -7.970 ;
        RECT 430.010 -8.240 430.350 -7.600 ;
        RECT 428.785 -9.085 429.160 -8.380 ;
        RECT 430.645 -8.515 431.010 -6.800 ;
        RECT 430.420 -9.555 431.010 -8.515 ;
        RECT 434.485 -8.565 434.715 -6.730 ;
        RECT 434.970 -8.160 436.235 -7.930 ;
        RECT 434.485 -8.795 435.760 -8.565 ;
        RECT 436.005 -9.590 436.235 -8.160 ;
        RECT 438.300 -9.310 438.635 -7.410 ;
        RECT 439.525 -8.565 439.755 -6.730 ;
        RECT 442.425 -7.485 442.655 -6.895 ;
        RECT 442.425 -7.715 444.115 -7.485 ;
        RECT 440.010 -8.160 441.275 -7.930 ;
        RECT 439.525 -8.795 440.800 -8.565 ;
        RECT 441.045 -9.590 441.275 -8.160 ;
        RECT 442.360 -8.350 443.650 -7.970 ;
        RECT 443.885 -8.610 444.115 -7.715 ;
        RECT 442.325 -8.840 444.115 -8.610 ;
        RECT 444.345 -7.505 444.695 -6.905 ;
        RECT 445.745 -7.130 446.995 -6.900 ;
        RECT 454.290 -6.960 456.505 -6.730 ;
        RECT 445.745 -7.505 445.975 -7.130 ;
        RECT 444.345 -7.735 445.975 -7.505 ;
        RECT 446.205 -7.700 446.535 -7.360 ;
        RECT 442.325 -9.310 442.555 -8.840 ;
        RECT 444.345 -9.025 444.575 -7.735 ;
        RECT 444.970 -8.350 446.000 -7.970 ;
        RECT 444.345 -9.255 444.850 -9.025 ;
        RECT 446.305 -9.045 446.535 -7.700 ;
        RECT 446.765 -8.210 446.995 -7.130 ;
        RECT 448.245 -7.360 448.475 -7.165 ;
        RECT 450.845 -7.360 451.075 -6.990 ;
        RECT 447.225 -7.820 447.455 -7.360 ;
        RECT 448.245 -7.590 451.075 -7.360 ;
        RECT 452.520 -7.275 453.160 -7.045 ;
        RECT 451.935 -7.820 452.235 -7.595 ;
        RECT 447.225 -8.050 452.235 -7.820 ;
        RECT 446.305 -9.275 446.710 -9.045 ;
        RECT 447.545 -9.330 447.775 -8.050 ;
        RECT 452.520 -8.280 452.750 -7.275 ;
        RECT 454.290 -8.070 454.520 -6.960 ;
        RECT 456.275 -7.070 456.505 -6.960 ;
        RECT 457.315 -6.960 458.500 -6.730 ;
        RECT 457.315 -7.070 457.545 -6.960 ;
        RECT 448.770 -8.510 452.750 -8.280 ;
        RECT 453.630 -8.300 454.520 -8.070 ;
        RECT 448.125 -8.740 448.355 -8.530 ;
        RECT 448.125 -8.970 451.310 -8.740 ;
        RECT 451.080 -9.360 451.310 -8.970 ;
        RECT 452.070 -9.120 452.410 -8.510 ;
        RECT 453.005 -9.360 453.235 -8.530 ;
        RECT 453.630 -9.120 453.970 -8.300 ;
        RECT 454.970 -8.530 455.200 -7.595 ;
        RECT 454.200 -8.760 455.200 -8.530 ;
        RECT 454.200 -9.360 454.430 -8.760 ;
        RECT 455.495 -8.990 455.835 -7.190 ;
        RECT 456.275 -7.300 457.545 -7.070 ;
        RECT 457.810 -7.715 458.040 -7.190 ;
        RECT 456.075 -7.945 458.040 -7.715 ;
        RECT 455.030 -9.330 455.835 -8.990 ;
        RECT 456.740 -9.100 457.285 -8.290 ;
        RECT 457.810 -8.440 458.040 -7.945 ;
        RECT 458.270 -8.210 458.500 -6.960 ;
        RECT 457.810 -8.670 460.310 -8.440 ;
        RECT 456.740 -9.150 458.375 -9.100 ;
        RECT 451.080 -9.590 454.430 -9.360 ;
        RECT 456.730 -9.410 458.375 -9.150 ;
        RECT 458.730 -9.330 458.960 -8.670 ;
        RECT 456.740 -9.460 458.375 -9.410 ;
        RECT 460.555 -9.570 460.990 -6.740 ;
        RECT 230.275 -11.465 230.655 -10.565 ;
        RECT 233.790 -11.465 234.170 -10.565 ;
        RECT 298.805 -11.160 299.035 -10.795 ;
        RECT 301.045 -11.160 301.275 -10.795 ;
        RECT 303.285 -11.160 303.515 -10.795 ;
        RECT 305.495 -11.160 305.755 -10.795 ;
        RECT 307.765 -11.135 307.995 -10.795 ;
        RECT 310.005 -11.135 310.235 -10.795 ;
        RECT 298.805 -11.540 305.755 -11.160 ;
        RECT 307.285 -11.370 310.235 -11.135 ;
        RECT 298.060 -12.150 301.260 -11.805 ;
        RECT 301.960 -12.450 302.760 -11.540 ;
        RECT 307.285 -11.805 307.620 -11.370 ;
        RECT 303.330 -12.145 307.620 -11.805 ;
        RECT 311.845 -11.675 313.120 -11.445 ;
        RECT 298.905 -12.830 305.755 -12.450 ;
        RECT 298.905 -13.010 299.135 -12.830 ;
        RECT 298.870 -13.390 299.135 -13.010 ;
        RECT 298.905 -13.500 299.135 -13.390 ;
        RECT 301.145 -13.500 301.375 -12.830 ;
        RECT 303.385 -13.500 303.615 -12.830 ;
        RECT 305.525 -13.500 305.755 -12.830 ;
        RECT 307.285 -12.650 307.620 -12.145 ;
        RECT 308.090 -12.270 310.950 -11.835 ;
        RECT 307.285 -12.880 310.335 -12.650 ;
        RECT 307.865 -13.500 308.095 -12.880 ;
        RECT 310.105 -13.500 310.335 -12.880 ;
        RECT 311.845 -13.510 312.075 -11.675 ;
        RECT 313.365 -12.080 313.595 -10.650 ;
        RECT 312.330 -12.310 313.595 -12.080 ;
        RECT 314.085 -11.675 315.360 -11.445 ;
        RECT 314.085 -13.510 314.315 -11.675 ;
        RECT 315.605 -12.080 315.835 -10.650 ;
        RECT 314.570 -12.310 315.835 -12.080 ;
        RECT 316.325 -11.675 317.600 -11.445 ;
        RECT 316.325 -13.510 316.555 -11.675 ;
        RECT 317.845 -12.080 318.075 -10.650 ;
        RECT 316.810 -12.310 318.075 -12.080 ;
        RECT 318.565 -11.675 319.840 -11.445 ;
        RECT 318.565 -13.510 318.795 -11.675 ;
        RECT 320.085 -12.080 320.315 -10.650 ;
        RECT 319.050 -12.310 320.315 -12.080 ;
        RECT 320.805 -11.675 322.080 -11.445 ;
        RECT 320.805 -13.510 321.035 -11.675 ;
        RECT 322.325 -12.080 322.555 -10.650 ;
        RECT 321.290 -12.310 322.555 -12.080 ;
        RECT 323.045 -11.675 324.320 -11.445 ;
        RECT 323.045 -13.510 323.275 -11.675 ;
        RECT 324.565 -12.080 324.795 -10.650 ;
        RECT 323.530 -12.310 324.795 -12.080 ;
        RECT 325.285 -11.675 326.560 -11.445 ;
        RECT 325.285 -13.510 325.515 -11.675 ;
        RECT 326.805 -12.080 327.035 -10.650 ;
        RECT 325.770 -12.310 327.035 -12.080 ;
        RECT 327.525 -11.675 328.800 -11.445 ;
        RECT 327.525 -13.510 327.755 -11.675 ;
        RECT 329.045 -12.080 329.275 -10.650 ;
        RECT 328.010 -12.310 329.275 -12.080 ;
        RECT 329.765 -11.675 331.040 -11.445 ;
        RECT 329.765 -13.510 329.995 -11.675 ;
        RECT 331.285 -12.080 331.515 -10.650 ;
        RECT 330.250 -12.310 331.515 -12.080 ;
        RECT 332.005 -11.675 333.280 -11.445 ;
        RECT 332.005 -13.510 332.235 -11.675 ;
        RECT 333.525 -12.080 333.755 -10.650 ;
        RECT 332.490 -12.310 333.755 -12.080 ;
        RECT 336.485 -11.675 337.760 -11.445 ;
        RECT 336.485 -13.510 336.715 -11.675 ;
        RECT 338.005 -12.080 338.235 -10.650 ;
        RECT 336.970 -12.310 338.235 -12.080 ;
        RECT 338.725 -11.675 340.000 -11.445 ;
        RECT 338.725 -13.510 338.955 -11.675 ;
        RECT 340.245 -12.080 340.475 -10.650 ;
        RECT 339.210 -12.310 340.475 -12.080 ;
        RECT 340.965 -11.675 342.240 -11.445 ;
        RECT 340.965 -13.510 341.195 -11.675 ;
        RECT 342.485 -12.080 342.715 -10.650 ;
        RECT 341.450 -12.310 342.715 -12.080 ;
        RECT 343.205 -11.675 344.480 -11.445 ;
        RECT 343.205 -13.510 343.435 -11.675 ;
        RECT 344.725 -12.080 344.955 -10.650 ;
        RECT 343.690 -12.310 344.955 -12.080 ;
        RECT 347.570 -13.500 347.970 -10.660 ;
        RECT 349.780 -10.900 351.140 -10.670 ;
        RECT 349.780 -11.205 350.010 -10.900 ;
        RECT 348.265 -11.435 350.010 -11.205 ;
        RECT 348.265 -11.900 348.495 -11.435 ;
        RECT 349.200 -13.405 349.550 -11.665 ;
        RECT 349.780 -13.085 350.010 -11.435 ;
        RECT 350.240 -11.770 351.540 -11.370 ;
        RECT 351.895 -11.700 353.545 -11.370 ;
        RECT 351.230 -11.930 351.540 -11.770 ;
        RECT 350.640 -12.610 350.980 -12.080 ;
        RECT 351.230 -12.315 353.690 -11.930 ;
        RECT 354.030 -12.610 354.370 -10.660 ;
        RECT 350.640 -12.845 354.370 -12.610 ;
        RECT 349.780 -13.315 351.580 -13.085 ;
        RECT 353.985 -13.510 354.370 -12.845 ;
        RECT 354.965 -11.675 356.240 -11.445 ;
        RECT 354.965 -13.510 355.195 -11.675 ;
        RECT 356.485 -12.080 356.715 -10.650 ;
        RECT 355.450 -12.310 356.715 -12.080 ;
        RECT 357.205 -11.675 358.480 -11.445 ;
        RECT 357.205 -13.510 357.435 -11.675 ;
        RECT 358.725 -12.080 358.955 -10.650 ;
        RECT 361.345 -11.400 361.575 -10.920 ;
        RECT 357.690 -12.310 358.955 -12.080 ;
        RECT 360.430 -11.630 361.575 -11.400 ;
        RECT 360.430 -12.480 360.770 -11.630 ;
        RECT 363.160 -11.860 363.535 -10.670 ;
        RECT 361.030 -12.160 362.350 -11.860 ;
        RECT 360.430 -12.830 361.575 -12.480 ;
        RECT 361.345 -13.510 361.575 -12.830 ;
        RECT 362.025 -12.710 362.350 -12.160 ;
        RECT 362.590 -12.270 363.535 -11.860 ;
        RECT 363.765 -12.710 363.995 -10.925 ;
        RECT 362.025 -12.940 363.995 -12.710 ;
        RECT 363.765 -13.510 363.995 -12.940 ;
        RECT 366.610 -13.500 367.010 -10.660 ;
        RECT 368.820 -10.900 370.180 -10.670 ;
        RECT 368.820 -11.205 369.050 -10.900 ;
        RECT 367.305 -11.435 369.050 -11.205 ;
        RECT 367.305 -11.900 367.535 -11.435 ;
        RECT 368.240 -13.405 368.590 -11.665 ;
        RECT 368.820 -13.085 369.050 -11.435 ;
        RECT 369.280 -11.770 370.580 -11.370 ;
        RECT 370.935 -11.700 372.585 -11.370 ;
        RECT 370.270 -11.930 370.580 -11.770 ;
        RECT 369.680 -12.610 370.020 -12.080 ;
        RECT 370.270 -12.315 372.730 -11.930 ;
        RECT 373.070 -12.610 373.410 -10.660 ;
        RECT 369.680 -12.845 373.410 -12.610 ;
        RECT 368.820 -13.315 370.620 -13.085 ;
        RECT 373.025 -13.510 373.410 -12.845 ;
        RECT 375.685 -11.675 376.960 -11.445 ;
        RECT 375.685 -13.510 375.915 -11.675 ;
        RECT 377.205 -12.080 377.435 -10.650 ;
        RECT 377.860 -10.880 384.645 -10.650 ;
        RECT 384.415 -10.985 384.645 -10.880 ;
        RECT 385.530 -10.880 387.325 -10.650 ;
        RECT 385.530 -10.985 385.760 -10.880 ;
        RECT 376.170 -12.310 377.435 -12.080 ;
        RECT 378.505 -12.470 378.825 -11.280 ;
        RECT 379.210 -11.340 379.550 -11.110 ;
        RECT 381.450 -11.340 381.790 -11.110 ;
        RECT 384.415 -11.215 385.760 -10.985 ;
        RECT 390.610 -11.095 391.960 -10.650 ;
        RECT 391.730 -11.110 391.960 -11.095 ;
        RECT 392.770 -11.040 394.560 -10.650 ;
        RECT 392.770 -11.110 393.000 -11.040 ;
        RECT 379.210 -11.680 383.160 -11.340 ;
        RECT 379.240 -12.240 381.550 -11.910 ;
        RECT 381.800 -12.240 382.580 -11.910 ;
        RECT 381.800 -12.470 382.060 -12.240 ;
        RECT 378.505 -12.800 382.060 -12.470 ;
        RECT 382.830 -12.490 383.160 -11.680 ;
        RECT 383.400 -11.445 384.165 -11.310 ;
        RECT 386.060 -11.445 387.100 -11.310 ;
        RECT 391.730 -11.340 393.000 -11.110 ;
        RECT 394.330 -11.110 394.560 -11.040 ;
        RECT 395.360 -11.040 397.150 -10.650 ;
        RECT 395.360 -11.110 395.590 -11.040 ;
        RECT 383.400 -11.675 387.100 -11.445 ;
        RECT 390.050 -11.570 391.500 -11.385 ;
        RECT 393.475 -11.570 393.835 -11.290 ;
        RECT 394.330 -11.340 395.590 -11.110 ;
        RECT 396.920 -11.110 397.150 -11.040 ;
        RECT 397.950 -11.110 399.755 -10.650 ;
        RECT 400.650 -11.095 402.270 -10.650 ;
        RECT 400.650 -11.110 401.625 -11.095 ;
        RECT 396.270 -11.570 396.615 -11.290 ;
        RECT 396.920 -11.340 401.625 -11.110 ;
        RECT 402.040 -11.110 402.270 -11.095 ;
        RECT 403.070 -11.040 404.690 -10.650 ;
        RECT 403.070 -11.110 403.300 -11.040 ;
        RECT 402.040 -11.340 403.300 -11.110 ;
        RECT 404.460 -11.110 404.690 -11.040 ;
        RECT 405.490 -11.040 407.110 -10.650 ;
        RECT 405.490 -11.110 405.720 -11.040 ;
        RECT 390.050 -11.655 398.305 -11.570 ;
        RECT 399.090 -11.600 401.625 -11.340 ;
        RECT 403.575 -11.570 403.920 -11.290 ;
        RECT 404.460 -11.340 405.720 -11.110 ;
        RECT 406.880 -11.110 407.110 -11.040 ;
        RECT 407.910 -11.095 408.990 -10.650 ;
        RECT 407.910 -11.110 408.140 -11.095 ;
        RECT 406.310 -11.570 406.650 -11.290 ;
        RECT 406.880 -11.340 408.140 -11.110 ;
        RECT 408.400 -11.570 409.550 -11.385 ;
        RECT 399.090 -11.640 400.500 -11.600 ;
        RECT 383.400 -12.270 383.720 -11.675 ;
        RECT 383.960 -12.260 386.000 -11.920 ;
        RECT 386.545 -12.310 387.100 -11.675 ;
        RECT 391.270 -11.800 398.305 -11.655 ;
        RECT 390.050 -12.030 391.020 -11.890 ;
        RECT 398.535 -12.030 399.650 -11.890 ;
        RECT 390.050 -12.270 399.650 -12.030 ;
        RECT 382.310 -12.500 383.160 -12.490 ;
        RECT 399.920 -12.500 400.500 -11.640 ;
        RECT 401.950 -11.655 409.550 -11.570 ;
        RECT 401.950 -11.800 408.620 -11.655 ;
        RECT 400.765 -12.030 401.700 -11.850 ;
        RECT 408.865 -12.030 409.550 -11.940 ;
        RECT 400.765 -12.270 409.550 -12.030 ;
        RECT 382.310 -12.800 386.240 -12.500 ;
        RECT 382.310 -13.040 382.540 -12.800 ;
        RECT 379.810 -13.400 382.540 -13.040 ;
        RECT 383.970 -13.070 384.200 -12.800 ;
        RECT 383.930 -13.330 384.310 -13.070 ;
        RECT 383.970 -13.395 384.200 -13.330 ;
        RECT 386.010 -13.395 386.240 -12.800 ;
        RECT 389.780 -13.270 390.120 -12.650 ;
        RECT 392.090 -12.775 400.500 -12.500 ;
        RECT 392.090 -12.955 392.945 -12.775 ;
        RECT 397.250 -12.785 400.500 -12.775 ;
        RECT 401.420 -12.770 409.765 -12.535 ;
        RECT 397.250 -12.960 397.590 -12.785 ;
        RECT 394.930 -13.270 395.270 -13.065 ;
        RECT 401.420 -13.270 401.650 -12.770 ;
        RECT 389.780 -13.505 401.650 -13.270 ;
        RECT 405.025 -13.510 405.255 -12.770 ;
        RECT 409.535 -13.500 409.765 -12.770 ;
        RECT 410.865 -13.440 411.170 -11.300 ;
        RECT 411.400 -12.480 411.755 -10.720 ;
        RECT 411.985 -11.910 412.290 -10.720 ;
        RECT 411.985 -12.250 413.015 -11.910 ;
        RECT 411.400 -12.510 412.825 -12.480 ;
        RECT 416.565 -12.510 416.795 -10.690 ;
        RECT 417.025 -11.745 417.335 -10.730 ;
        RECT 418.995 -11.185 419.225 -10.690 ;
        RECT 418.995 -11.420 420.120 -11.185 ;
        RECT 417.025 -12.270 417.970 -11.745 ;
        RECT 418.220 -12.010 419.560 -11.670 ;
        RECT 418.220 -12.510 418.450 -12.010 ;
        RECT 419.800 -12.330 420.120 -11.420 ;
        RECT 411.400 -12.770 412.870 -12.510 ;
        RECT 416.565 -12.745 418.450 -12.510 ;
        RECT 411.400 -12.800 412.825 -12.770 ;
        RECT 412.545 -13.500 412.825 -12.800 ;
        RECT 416.565 -13.510 416.795 -12.745 ;
        RECT 418.995 -12.820 420.120 -12.330 ;
        RECT 421.045 -11.675 422.320 -11.445 ;
        RECT 418.995 -13.510 419.225 -12.820 ;
        RECT 421.045 -13.510 421.275 -11.675 ;
        RECT 422.565 -12.080 422.795 -10.650 ;
        RECT 421.530 -12.310 422.795 -12.080 ;
        RECT 423.285 -11.675 424.560 -11.445 ;
        RECT 423.285 -13.510 423.515 -11.675 ;
        RECT 424.805 -12.080 425.035 -10.650 ;
        RECT 423.770 -12.310 425.035 -12.080 ;
        RECT 425.970 -13.500 426.405 -10.670 ;
        RECT 428.000 -11.570 428.230 -10.910 ;
        RECT 428.585 -11.140 430.220 -10.780 ;
        RECT 432.530 -10.880 435.880 -10.650 ;
        RECT 426.650 -11.800 429.150 -11.570 ;
        RECT 428.460 -13.280 428.690 -12.030 ;
        RECT 428.920 -12.295 429.150 -11.800 ;
        RECT 429.675 -11.950 430.220 -11.140 ;
        RECT 431.125 -11.250 431.930 -10.910 ;
        RECT 428.920 -12.525 430.885 -12.295 ;
        RECT 428.920 -13.050 429.150 -12.525 ;
        RECT 429.415 -13.170 430.685 -12.940 ;
        RECT 431.125 -13.050 431.465 -11.250 ;
        RECT 432.530 -11.480 432.760 -10.880 ;
        RECT 431.760 -11.710 432.760 -11.480 ;
        RECT 431.760 -12.645 431.990 -11.710 ;
        RECT 432.990 -11.940 433.330 -11.120 ;
        RECT 433.725 -11.710 433.955 -10.880 ;
        RECT 434.550 -11.730 434.890 -11.120 ;
        RECT 435.650 -11.270 435.880 -10.880 ;
        RECT 435.650 -11.500 438.835 -11.270 ;
        RECT 438.605 -11.710 438.835 -11.500 ;
        RECT 432.440 -12.170 433.330 -11.940 ;
        RECT 434.210 -11.960 438.190 -11.730 ;
        RECT 429.415 -13.280 429.645 -13.170 ;
        RECT 428.460 -13.510 429.645 -13.280 ;
        RECT 430.455 -13.280 430.685 -13.170 ;
        RECT 432.440 -13.280 432.670 -12.170 ;
        RECT 434.210 -12.965 434.440 -11.960 ;
        RECT 439.185 -12.190 439.415 -10.910 ;
        RECT 446.150 -10.930 446.410 -10.770 ;
        RECT 440.250 -11.195 440.655 -10.965 ;
        RECT 434.725 -12.420 439.735 -12.190 ;
        RECT 434.725 -12.645 435.025 -12.420 ;
        RECT 433.800 -13.195 434.440 -12.965 ;
        RECT 435.885 -12.880 438.715 -12.650 ;
        RECT 439.505 -12.880 439.735 -12.420 ;
        RECT 435.885 -13.250 436.115 -12.880 ;
        RECT 438.485 -13.075 438.715 -12.880 ;
        RECT 439.965 -13.110 440.195 -12.030 ;
        RECT 440.425 -12.540 440.655 -11.195 ;
        RECT 442.110 -11.215 442.615 -10.985 ;
        RECT 440.960 -12.270 441.990 -11.890 ;
        RECT 442.385 -12.505 442.615 -11.215 ;
        RECT 444.405 -11.400 444.635 -10.930 ;
        RECT 440.425 -12.880 440.755 -12.540 ;
        RECT 440.985 -12.735 442.615 -12.505 ;
        RECT 440.985 -13.110 441.215 -12.735 ;
        RECT 430.455 -13.510 432.670 -13.280 ;
        RECT 439.965 -13.340 441.215 -13.110 ;
        RECT 442.265 -13.335 442.615 -12.735 ;
        RECT 442.845 -11.630 444.635 -11.400 ;
        RECT 442.845 -12.525 443.075 -11.630 ;
        RECT 443.310 -12.270 444.600 -11.890 ;
        RECT 442.845 -12.755 444.535 -12.525 ;
        RECT 444.305 -13.345 444.535 -12.755 ;
        RECT 446.140 -12.830 446.475 -10.930 ;
        RECT 447.365 -11.675 448.640 -11.445 ;
        RECT 447.365 -13.510 447.595 -11.675 ;
        RECT 448.885 -12.080 449.115 -10.650 ;
        RECT 447.850 -12.310 449.115 -12.080 ;
        RECT 449.605 -11.675 450.880 -11.445 ;
        RECT 449.605 -13.510 449.835 -11.675 ;
        RECT 451.125 -12.080 451.355 -10.650 ;
        RECT 450.090 -12.310 451.355 -12.080 ;
        RECT 454.085 -11.675 455.360 -11.445 ;
        RECT 454.085 -13.510 454.315 -11.675 ;
        RECT 455.605 -12.080 455.835 -10.650 ;
        RECT 454.570 -12.310 455.835 -12.080 ;
        RECT 456.325 -11.675 457.600 -11.445 ;
        RECT 456.325 -13.510 456.555 -11.675 ;
        RECT 457.845 -12.080 458.075 -10.650 ;
        RECT 456.810 -12.310 458.075 -12.080 ;
        RECT 458.565 -11.675 459.840 -11.445 ;
        RECT 458.565 -13.510 458.795 -11.675 ;
        RECT 460.085 -12.080 460.315 -10.650 ;
        RECT 459.050 -12.310 460.315 -12.080 ;
        RECT 297.285 -16.405 297.515 -14.570 ;
        RECT 297.770 -16.000 299.035 -15.770 ;
        RECT 297.285 -16.635 298.560 -16.405 ;
        RECT 298.805 -17.430 299.035 -16.000 ;
        RECT 299.925 -17.430 300.255 -14.570 ;
        RECT 301.765 -15.145 302.150 -14.570 ;
        RECT 301.765 -15.380 303.775 -15.145 ;
        RECT 300.485 -16.760 300.810 -15.760 ;
        RECT 301.765 -17.160 301.995 -15.380 ;
        RECT 302.225 -16.330 303.110 -15.770 ;
        RECT 303.490 -16.130 303.775 -15.380 ;
        RECT 302.225 -17.310 302.740 -16.330 ;
        RECT 304.005 -16.360 304.475 -14.580 ;
        RECT 303.850 -17.385 304.475 -16.360 ;
        RECT 305.585 -16.990 305.910 -15.010 ;
        RECT 306.140 -17.360 306.475 -14.590 ;
        RECT 308.380 -17.150 308.715 -15.250 ;
        RECT 309.605 -16.405 309.835 -14.570 ;
        RECT 310.090 -16.000 311.355 -15.770 ;
        RECT 309.605 -16.635 310.880 -16.405 ;
        RECT 311.125 -17.430 311.355 -16.000 ;
        RECT 311.845 -16.405 312.075 -14.570 ;
        RECT 312.330 -16.000 313.595 -15.770 ;
        RECT 311.845 -16.635 313.120 -16.405 ;
        RECT 313.365 -17.430 313.595 -16.000 ;
        RECT 316.885 -16.405 317.115 -14.570 ;
        RECT 317.370 -16.000 318.635 -15.770 ;
        RECT 316.885 -16.635 318.160 -16.405 ;
        RECT 318.405 -17.430 318.635 -16.000 ;
        RECT 319.125 -16.405 319.355 -14.570 ;
        RECT 321.470 -15.670 322.100 -14.615 ;
        RECT 319.610 -16.000 320.875 -15.770 ;
        RECT 319.125 -16.635 320.400 -16.405 ;
        RECT 320.645 -17.430 320.875 -16.000 ;
        RECT 321.470 -16.920 321.800 -15.670 ;
        RECT 323.460 -16.220 323.820 -14.615 ;
        RECT 324.060 -14.830 325.265 -14.600 ;
        RECT 322.065 -16.450 322.920 -16.320 ;
        RECT 324.060 -16.450 324.290 -14.830 ;
        RECT 322.065 -16.680 324.290 -16.450 ;
        RECT 321.470 -17.350 322.235 -16.920 ;
        RECT 323.895 -17.430 324.290 -16.680 ;
        RECT 324.520 -16.885 324.940 -15.080 ;
        RECT 328.645 -15.145 329.030 -14.570 ;
        RECT 326.860 -17.150 327.195 -15.250 ;
        RECT 328.645 -15.380 330.655 -15.145 ;
        RECT 326.870 -17.310 327.130 -17.150 ;
        RECT 328.645 -17.160 328.875 -15.380 ;
        RECT 329.105 -16.330 329.990 -15.770 ;
        RECT 330.370 -16.130 330.655 -15.380 ;
        RECT 329.105 -17.310 329.620 -16.330 ;
        RECT 330.885 -16.360 331.355 -14.580 ;
        RECT 332.105 -15.325 332.335 -14.735 ;
        RECT 332.105 -15.555 333.795 -15.325 ;
        RECT 331.910 -16.190 333.330 -15.810 ;
        RECT 330.730 -17.385 331.355 -16.360 ;
        RECT 333.565 -16.450 333.795 -15.555 ;
        RECT 332.005 -16.680 333.795 -16.450 ;
        RECT 334.025 -15.345 334.375 -14.745 ;
        RECT 335.425 -14.970 336.675 -14.740 ;
        RECT 343.970 -14.800 346.185 -14.570 ;
        RECT 335.425 -15.345 335.655 -14.970 ;
        RECT 334.025 -15.575 335.655 -15.345 ;
        RECT 335.885 -15.540 336.215 -15.200 ;
        RECT 332.005 -17.150 332.235 -16.680 ;
        RECT 334.025 -16.865 334.255 -15.575 ;
        RECT 334.650 -16.190 335.680 -15.810 ;
        RECT 334.025 -17.095 334.530 -16.865 ;
        RECT 335.985 -16.885 336.215 -15.540 ;
        RECT 336.445 -16.050 336.675 -14.970 ;
        RECT 337.925 -15.200 338.155 -15.005 ;
        RECT 340.525 -15.200 340.755 -14.830 ;
        RECT 336.905 -15.660 337.135 -15.200 ;
        RECT 337.925 -15.430 340.755 -15.200 ;
        RECT 342.200 -15.115 342.840 -14.885 ;
        RECT 341.615 -15.660 341.915 -15.435 ;
        RECT 336.905 -15.890 341.915 -15.660 ;
        RECT 335.985 -17.115 336.390 -16.885 ;
        RECT 337.225 -17.170 337.455 -15.890 ;
        RECT 342.200 -16.120 342.430 -15.115 ;
        RECT 343.970 -15.910 344.200 -14.800 ;
        RECT 345.955 -14.910 346.185 -14.800 ;
        RECT 346.995 -14.800 348.180 -14.570 ;
        RECT 346.995 -14.910 347.225 -14.800 ;
        RECT 338.450 -16.350 342.430 -16.120 ;
        RECT 343.310 -16.140 344.200 -15.910 ;
        RECT 337.805 -16.580 338.035 -16.370 ;
        RECT 337.805 -16.810 340.990 -16.580 ;
        RECT 340.760 -17.200 340.990 -16.810 ;
        RECT 341.750 -16.960 342.090 -16.350 ;
        RECT 342.685 -17.200 342.915 -16.370 ;
        RECT 343.310 -16.960 343.650 -16.140 ;
        RECT 344.650 -16.370 344.880 -15.435 ;
        RECT 343.880 -16.600 344.880 -16.370 ;
        RECT 343.880 -17.200 344.110 -16.600 ;
        RECT 345.175 -16.830 345.515 -15.030 ;
        RECT 345.955 -15.140 347.225 -14.910 ;
        RECT 347.490 -15.555 347.720 -15.030 ;
        RECT 345.755 -15.785 347.720 -15.555 ;
        RECT 344.710 -17.170 345.515 -16.830 ;
        RECT 346.420 -16.940 346.965 -16.130 ;
        RECT 347.490 -16.280 347.720 -15.785 ;
        RECT 347.950 -16.050 348.180 -14.800 ;
        RECT 347.490 -16.510 349.990 -16.280 ;
        RECT 346.420 -16.990 348.055 -16.940 ;
        RECT 340.760 -17.430 344.110 -17.200 ;
        RECT 346.410 -17.250 348.055 -16.990 ;
        RECT 348.410 -17.170 348.640 -16.510 ;
        RECT 346.420 -17.300 348.055 -17.250 ;
        RECT 350.235 -17.410 350.670 -14.580 ;
        RECT 351.045 -15.145 351.430 -14.570 ;
        RECT 351.045 -15.380 353.055 -15.145 ;
        RECT 351.045 -17.160 351.275 -15.380 ;
        RECT 351.505 -16.330 352.390 -15.770 ;
        RECT 352.770 -16.130 353.055 -15.380 ;
        RECT 351.505 -17.310 352.020 -16.330 ;
        RECT 353.285 -16.360 353.755 -14.580 ;
        RECT 353.130 -17.385 353.755 -16.360 ;
        RECT 356.085 -16.405 356.315 -14.570 ;
        RECT 358.775 -15.280 359.055 -14.580 ;
        RECT 359.910 -15.280 360.170 -15.250 ;
        RECT 358.775 -15.600 360.200 -15.280 ;
        RECT 356.570 -16.000 357.835 -15.770 ;
        RECT 356.085 -16.635 357.360 -16.405 ;
        RECT 357.605 -17.430 357.835 -16.000 ;
        RECT 358.585 -16.170 359.615 -15.830 ;
        RECT 359.310 -17.360 359.615 -16.170 ;
        RECT 359.845 -17.360 360.200 -15.600 ;
        RECT 360.430 -16.780 360.735 -14.640 ;
        RECT 362.715 -14.750 364.650 -14.590 ;
        RECT 362.650 -14.820 364.650 -14.750 ;
        RECT 362.650 -14.925 363.030 -14.820 ;
        RECT 362.145 -15.010 363.030 -14.925 ;
        RECT 362.145 -15.160 362.945 -15.010 ;
        RECT 362.145 -16.640 362.415 -15.160 ;
        RECT 363.260 -15.580 366.230 -15.260 ;
        RECT 363.260 -15.810 363.560 -15.580 ;
        RECT 362.650 -16.190 363.560 -15.810 ;
        RECT 363.820 -16.190 365.560 -15.810 ;
        RECT 365.980 -16.380 366.230 -15.580 ;
        RECT 367.285 -16.405 367.515 -14.570 ;
        RECT 367.770 -16.000 369.035 -15.770 ;
        RECT 367.285 -16.635 368.560 -16.405 ;
        RECT 362.145 -16.910 365.675 -16.640 ;
        RECT 363.205 -17.430 363.435 -16.910 ;
        RECT 365.445 -17.430 365.675 -16.910 ;
        RECT 368.805 -17.430 369.035 -16.000 ;
        RECT 370.545 -16.780 370.850 -14.640 ;
        RECT 372.225 -15.280 372.505 -14.580 ;
        RECT 371.080 -15.600 372.505 -15.280 ;
        RECT 371.080 -17.360 371.435 -15.600 ;
        RECT 371.665 -16.170 372.695 -15.830 ;
        RECT 371.665 -17.360 371.970 -16.170 ;
        RECT 373.445 -16.405 373.675 -14.570 ;
        RECT 375.790 -15.670 376.420 -14.615 ;
        RECT 373.930 -16.000 375.195 -15.770 ;
        RECT 373.445 -16.635 374.720 -16.405 ;
        RECT 374.965 -17.430 375.195 -16.000 ;
        RECT 375.790 -16.920 376.120 -15.670 ;
        RECT 377.780 -16.220 378.140 -14.615 ;
        RECT 378.380 -14.830 379.585 -14.600 ;
        RECT 376.385 -16.450 377.240 -16.320 ;
        RECT 378.380 -16.450 378.610 -14.830 ;
        RECT 376.385 -16.680 378.610 -16.450 ;
        RECT 375.790 -17.350 376.555 -16.920 ;
        RECT 378.215 -17.430 378.610 -16.680 ;
        RECT 378.840 -16.885 379.260 -15.080 ;
        RECT 380.165 -15.145 380.550 -14.570 ;
        RECT 380.165 -15.380 382.175 -15.145 ;
        RECT 380.165 -17.160 380.395 -15.380 ;
        RECT 380.625 -16.330 381.510 -15.770 ;
        RECT 381.890 -16.130 382.175 -15.380 ;
        RECT 380.625 -17.310 381.140 -16.330 ;
        RECT 382.405 -16.360 382.875 -14.580 ;
        RECT 382.250 -17.385 382.875 -16.360 ;
        RECT 383.525 -16.405 383.755 -14.570 ;
        RECT 384.010 -16.000 385.275 -15.770 ;
        RECT 383.525 -16.635 384.800 -16.405 ;
        RECT 385.045 -17.430 385.275 -16.000 ;
        RECT 385.765 -16.405 385.995 -14.570 ;
        RECT 390.845 -14.800 393.165 -14.570 ;
        RECT 390.845 -15.600 391.075 -14.800 ;
        RECT 391.305 -15.370 392.690 -15.030 ;
        RECT 386.250 -16.000 387.515 -15.770 ;
        RECT 385.765 -16.635 387.040 -16.405 ;
        RECT 387.285 -17.430 387.515 -16.000 ;
        RECT 389.570 -16.060 390.545 -15.810 ;
        RECT 390.845 -15.830 391.435 -15.600 ;
        RECT 389.570 -16.360 390.975 -16.060 ;
        RECT 390.640 -17.410 390.975 -16.360 ;
        RECT 391.205 -17.410 391.435 -15.830 ;
        RECT 391.760 -17.410 392.095 -15.640 ;
        RECT 392.325 -17.410 392.690 -15.370 ;
        RECT 392.935 -15.270 393.165 -14.800 ;
        RECT 392.935 -15.500 393.675 -15.270 ;
        RECT 396.725 -15.280 396.955 -14.570 ;
        RECT 398.865 -15.280 399.095 -14.570 ;
        RECT 401.385 -15.140 401.615 -14.570 ;
        RECT 426.770 -14.720 427.110 -14.635 ;
        RECT 412.310 -14.905 413.360 -14.720 ;
        RECT 414.200 -14.905 415.400 -14.720 ;
        RECT 416.240 -14.905 417.440 -14.720 ;
        RECT 418.280 -14.905 419.585 -14.720 ;
        RECT 412.310 -14.935 419.585 -14.905 ;
        RECT 420.420 -14.935 424.285 -14.720 ;
        RECT 425.120 -14.935 427.110 -14.720 ;
        RECT 392.920 -17.410 393.215 -15.730 ;
        RECT 393.445 -17.410 393.675 -15.500 ;
        RECT 396.280 -15.600 399.095 -15.280 ;
        RECT 399.695 -15.370 401.615 -15.140 ;
        RECT 403.010 -15.245 408.605 -15.010 ;
        RECT 412.310 -15.040 427.110 -14.935 ;
        RECT 412.310 -15.165 420.670 -15.040 ;
        RECT 424.035 -15.165 425.370 -15.040 ;
        RECT 396.280 -16.450 396.600 -15.600 ;
        RECT 399.695 -15.920 399.925 -15.370 ;
        RECT 396.935 -16.220 399.925 -15.920 ;
        RECT 400.540 -16.220 402.260 -15.840 ;
        RECT 396.280 -16.680 399.095 -16.450 ;
        RECT 396.625 -17.270 396.855 -16.680 ;
        RECT 398.865 -17.270 399.095 -16.680 ;
        RECT 399.695 -16.460 399.925 -16.220 ;
        RECT 399.695 -16.690 401.515 -16.460 ;
        RECT 401.285 -17.270 401.515 -16.690 ;
        RECT 403.010 -16.860 403.310 -15.245 ;
        RECT 404.145 -15.710 409.055 -15.475 ;
        RECT 404.145 -15.810 404.420 -15.710 ;
        RECT 403.660 -16.190 404.420 -15.810 ;
        RECT 408.570 -15.810 409.055 -15.710 ;
        RECT 404.650 -16.175 407.930 -15.940 ;
        RECT 408.570 -16.175 409.550 -15.810 ;
        RECT 412.920 -16.160 419.010 -15.840 ;
        RECT 404.830 -16.430 407.080 -16.405 ;
        RECT 404.650 -16.690 407.080 -16.430 ;
        RECT 404.830 -16.695 407.080 -16.690 ;
        RECT 407.410 -16.425 407.930 -16.175 ;
        RECT 419.240 -16.405 419.560 -15.535 ;
        RECT 407.410 -16.700 409.125 -16.425 ;
        RECT 412.000 -16.635 419.560 -16.405 ;
        RECT 414.680 -16.740 416.830 -16.635 ;
        RECT 419.800 -16.740 420.120 -15.165 ;
        RECT 420.880 -15.600 423.805 -15.280 ;
        RECT 426.770 -15.485 427.110 -15.040 ;
        RECT 420.880 -15.840 421.220 -15.600 ;
        RECT 423.555 -15.820 423.805 -15.600 ;
        RECT 420.350 -16.190 421.220 -15.840 ;
        RECT 421.450 -16.190 423.220 -15.840 ;
        RECT 423.555 -16.050 429.140 -15.820 ;
        RECT 422.970 -16.280 423.220 -16.190 ;
        RECT 422.970 -16.510 427.800 -16.280 ;
        RECT 430.005 -16.405 430.235 -14.570 ;
        RECT 430.490 -16.000 431.755 -15.770 ;
        RECT 430.005 -16.635 431.280 -16.405 ;
        RECT 403.010 -16.985 404.250 -16.860 ;
        RECT 403.010 -17.095 406.875 -16.985 ;
        RECT 411.560 -17.095 414.430 -16.865 ;
        RECT 403.920 -17.255 406.875 -17.095 ;
        RECT 414.200 -17.200 414.430 -17.095 ;
        RECT 417.210 -17.095 419.105 -16.865 ;
        RECT 419.800 -16.970 428.240 -16.740 ;
        RECT 417.210 -17.200 417.440 -17.095 ;
        RECT 414.200 -17.430 417.440 -17.200 ;
        RECT 418.875 -17.200 419.105 -17.095 ;
        RECT 418.875 -17.430 429.580 -17.200 ;
        RECT 431.525 -17.430 431.755 -16.000 ;
        RECT 434.485 -16.405 434.715 -14.570 ;
        RECT 434.970 -16.000 436.235 -15.770 ;
        RECT 434.485 -16.635 435.760 -16.405 ;
        RECT 436.005 -17.430 436.235 -16.000 ;
        RECT 436.725 -16.405 436.955 -14.570 ;
        RECT 437.210 -16.000 438.475 -15.770 ;
        RECT 436.725 -16.635 438.000 -16.405 ;
        RECT 438.245 -17.430 438.475 -16.000 ;
        RECT 438.965 -16.405 439.195 -14.570 ;
        RECT 439.450 -16.000 440.715 -15.770 ;
        RECT 438.965 -16.635 440.240 -16.405 ;
        RECT 440.485 -17.430 440.715 -16.000 ;
        RECT 441.205 -16.405 441.435 -14.570 ;
        RECT 441.690 -16.000 442.955 -15.770 ;
        RECT 441.205 -16.635 442.480 -16.405 ;
        RECT 442.725 -17.430 442.955 -16.000 ;
        RECT 443.445 -16.405 443.675 -14.570 ;
        RECT 447.825 -15.200 448.055 -14.580 ;
        RECT 450.065 -15.200 450.295 -14.580 ;
        RECT 447.825 -15.430 450.875 -15.200 ;
        RECT 443.930 -16.000 445.195 -15.770 ;
        RECT 443.445 -16.635 444.720 -16.405 ;
        RECT 444.965 -17.430 445.195 -16.000 ;
        RECT 447.210 -16.245 450.070 -15.810 ;
        RECT 450.540 -15.935 450.875 -15.430 ;
        RECT 450.540 -16.275 454.830 -15.935 ;
        RECT 456.900 -16.275 460.100 -15.930 ;
        RECT 450.540 -16.710 450.875 -16.275 ;
        RECT 447.925 -16.945 450.875 -16.710 ;
        RECT 447.925 -17.285 448.155 -16.945 ;
        RECT 450.165 -17.285 450.395 -16.945 ;
        RECT 298.625 -19.240 298.855 -18.760 ;
        RECT 297.710 -19.470 298.855 -19.240 ;
        RECT 297.710 -20.320 298.050 -19.470 ;
        RECT 300.440 -19.700 300.815 -18.510 ;
        RECT 312.200 -18.720 315.550 -18.490 ;
        RECT 298.310 -20.000 299.630 -19.700 ;
        RECT 297.710 -20.670 298.855 -20.320 ;
        RECT 298.625 -21.350 298.855 -20.670 ;
        RECT 299.305 -20.550 299.630 -20.000 ;
        RECT 299.870 -20.110 300.815 -19.700 ;
        RECT 301.045 -20.550 301.275 -18.765 ;
        RECT 303.445 -19.240 303.675 -18.770 ;
        RECT 305.465 -19.055 305.970 -18.825 ;
        RECT 307.425 -19.035 307.830 -18.805 ;
        RECT 303.445 -19.470 305.235 -19.240 ;
        RECT 303.480 -20.110 304.770 -19.730 ;
        RECT 305.005 -20.365 305.235 -19.470 ;
        RECT 299.305 -20.780 301.275 -20.550 ;
        RECT 301.045 -21.350 301.275 -20.780 ;
        RECT 303.545 -20.595 305.235 -20.365 ;
        RECT 305.465 -20.345 305.695 -19.055 ;
        RECT 306.090 -20.110 307.120 -19.730 ;
        RECT 305.465 -20.575 307.095 -20.345 ;
        RECT 307.425 -20.380 307.655 -19.035 ;
        RECT 303.545 -21.185 303.775 -20.595 ;
        RECT 305.465 -21.175 305.815 -20.575 ;
        RECT 306.865 -20.950 307.095 -20.575 ;
        RECT 307.325 -20.720 307.655 -20.380 ;
        RECT 307.885 -20.950 308.115 -19.870 ;
        RECT 308.665 -20.030 308.895 -18.750 ;
        RECT 312.200 -19.110 312.430 -18.720 ;
        RECT 309.245 -19.340 312.430 -19.110 ;
        RECT 309.245 -19.550 309.475 -19.340 ;
        RECT 313.190 -19.570 313.530 -18.960 ;
        RECT 314.125 -19.550 314.355 -18.720 ;
        RECT 309.890 -19.800 313.870 -19.570 ;
        RECT 308.345 -20.260 313.355 -20.030 ;
        RECT 308.345 -20.720 308.575 -20.260 ;
        RECT 313.055 -20.485 313.355 -20.260 ;
        RECT 309.365 -20.720 312.195 -20.490 ;
        RECT 309.365 -20.915 309.595 -20.720 ;
        RECT 306.865 -21.180 308.115 -20.950 ;
        RECT 311.965 -21.090 312.195 -20.720 ;
        RECT 313.640 -20.805 313.870 -19.800 ;
        RECT 314.750 -19.780 315.090 -18.960 ;
        RECT 315.320 -19.320 315.550 -18.720 ;
        RECT 316.150 -19.090 316.955 -18.750 ;
        RECT 315.320 -19.550 316.320 -19.320 ;
        RECT 314.750 -20.010 315.640 -19.780 ;
        RECT 313.640 -21.035 314.280 -20.805 ;
        RECT 315.410 -21.120 315.640 -20.010 ;
        RECT 316.090 -20.485 316.320 -19.550 ;
        RECT 316.615 -20.890 316.955 -19.090 ;
        RECT 317.860 -18.980 319.495 -18.620 ;
        RECT 317.860 -19.790 318.405 -18.980 ;
        RECT 319.850 -19.410 320.080 -18.750 ;
        RECT 318.930 -19.640 321.430 -19.410 ;
        RECT 318.930 -20.135 319.160 -19.640 ;
        RECT 317.195 -20.365 319.160 -20.135 ;
        RECT 317.395 -21.010 318.665 -20.780 ;
        RECT 318.930 -20.890 319.160 -20.365 ;
        RECT 317.395 -21.120 317.625 -21.010 ;
        RECT 315.410 -21.350 317.625 -21.120 ;
        RECT 318.435 -21.120 318.665 -21.010 ;
        RECT 319.390 -21.120 319.620 -19.870 ;
        RECT 318.435 -21.350 319.620 -21.120 ;
        RECT 321.675 -21.340 322.110 -18.510 ;
        RECT 323.480 -18.830 324.820 -18.510 ;
        RECT 322.900 -19.730 323.250 -19.120 ;
        RECT 322.355 -20.110 323.250 -19.730 ;
        RECT 322.430 -21.120 322.770 -20.455 ;
        RECT 323.480 -20.685 323.785 -18.830 ;
        RECT 324.580 -19.730 324.920 -19.120 ;
        RECT 325.715 -19.730 326.055 -19.120 ;
        RECT 324.015 -20.110 324.920 -19.730 ;
        RECT 325.150 -20.110 326.055 -19.730 ;
        RECT 324.470 -21.120 324.810 -20.455 ;
        RECT 327.980 -20.670 328.315 -18.770 ;
        RECT 329.205 -19.515 330.480 -19.285 ;
        RECT 322.430 -21.350 324.810 -21.120 ;
        RECT 329.205 -21.350 329.435 -19.515 ;
        RECT 330.725 -19.920 330.955 -18.490 ;
        RECT 329.690 -20.150 330.955 -19.920 ;
        RECT 331.445 -19.515 332.720 -19.285 ;
        RECT 331.445 -21.350 331.675 -19.515 ;
        RECT 332.965 -19.920 333.195 -18.490 ;
        RECT 331.930 -20.150 333.195 -19.920 ;
        RECT 336.485 -19.515 337.760 -19.285 ;
        RECT 336.485 -21.350 336.715 -19.515 ;
        RECT 338.005 -19.920 338.235 -18.490 ;
        RECT 336.970 -20.150 338.235 -19.920 ;
        RECT 338.725 -19.515 340.000 -19.285 ;
        RECT 338.725 -21.350 338.955 -19.515 ;
        RECT 340.245 -19.920 340.475 -18.490 ;
        RECT 339.210 -20.150 340.475 -19.920 ;
        RECT 340.965 -19.515 342.240 -19.285 ;
        RECT 340.965 -21.350 341.195 -19.515 ;
        RECT 342.485 -19.920 342.715 -18.490 ;
        RECT 341.450 -20.150 342.715 -19.920 ;
        RECT 343.205 -19.515 344.480 -19.285 ;
        RECT 343.205 -21.350 343.435 -19.515 ;
        RECT 344.725 -19.920 344.955 -18.490 ;
        RECT 343.690 -20.150 344.955 -19.920 ;
        RECT 345.445 -19.515 346.720 -19.285 ;
        RECT 345.445 -21.350 345.675 -19.515 ;
        RECT 346.965 -19.920 347.195 -18.490 ;
        RECT 345.930 -20.150 347.195 -19.920 ;
        RECT 347.685 -19.515 348.960 -19.285 ;
        RECT 347.685 -21.350 347.915 -19.515 ;
        RECT 349.205 -19.920 349.435 -18.490 ;
        RECT 348.170 -20.150 349.435 -19.920 ;
        RECT 349.925 -19.515 351.200 -19.285 ;
        RECT 349.925 -21.350 350.155 -19.515 ;
        RECT 351.445 -19.920 351.675 -18.490 ;
        RECT 350.410 -20.150 351.675 -19.920 ;
        RECT 352.165 -19.515 353.440 -19.285 ;
        RECT 352.165 -21.350 352.395 -19.515 ;
        RECT 353.685 -19.920 353.915 -18.490 ;
        RECT 352.650 -20.150 353.915 -19.920 ;
        RECT 354.405 -19.515 355.680 -19.285 ;
        RECT 354.405 -21.350 354.635 -19.515 ;
        RECT 355.925 -19.920 356.155 -18.490 ;
        RECT 354.890 -20.150 356.155 -19.920 ;
        RECT 356.645 -19.515 357.920 -19.285 ;
        RECT 356.645 -21.350 356.875 -19.515 ;
        RECT 358.165 -19.920 358.395 -18.490 ;
        RECT 357.130 -20.150 358.395 -19.920 ;
        RECT 358.885 -19.515 360.160 -19.285 ;
        RECT 358.885 -21.350 359.115 -19.515 ;
        RECT 360.405 -19.920 360.635 -18.490 ;
        RECT 359.370 -20.150 360.635 -19.920 ;
        RECT 361.125 -19.515 362.400 -19.285 ;
        RECT 361.125 -21.350 361.355 -19.515 ;
        RECT 362.645 -19.920 362.875 -18.490 ;
        RECT 366.330 -18.830 366.670 -18.520 ;
        RECT 368.570 -18.830 368.910 -18.520 ;
        RECT 366.330 -19.060 369.405 -18.830 ;
        RECT 369.175 -19.200 369.405 -19.060 ;
        RECT 370.405 -18.960 372.170 -18.640 ;
        RECT 370.405 -19.200 370.665 -18.960 ;
        RECT 369.175 -19.520 370.665 -19.200 ;
        RECT 371.010 -19.520 373.160 -19.200 ;
        RECT 361.610 -20.150 362.875 -19.920 ;
        RECT 365.295 -20.080 366.435 -19.760 ;
        RECT 366.925 -20.080 368.670 -19.760 ;
        RECT 365.890 -20.320 366.435 -20.080 ;
        RECT 369.100 -20.320 369.720 -19.760 ;
        RECT 365.365 -20.785 365.595 -20.460 ;
        RECT 365.890 -20.555 369.720 -20.320 ;
        RECT 368.655 -20.670 369.720 -20.555 ;
        RECT 369.960 -20.320 370.280 -19.520 ;
        RECT 370.550 -20.080 373.900 -19.760 ;
        RECT 369.960 -20.740 373.150 -20.320 ;
        RECT 365.365 -21.015 368.410 -20.785 ;
        RECT 365.365 -21.350 365.595 -21.015 ;
        RECT 368.180 -21.120 368.410 -21.015 ;
        RECT 373.845 -21.120 374.075 -20.460 ;
        RECT 368.180 -21.350 374.075 -21.120 ;
        RECT 376.085 -21.350 376.415 -18.490 ;
        RECT 376.645 -20.160 376.970 -19.160 ;
        RECT 377.925 -19.515 379.200 -19.285 ;
        RECT 377.925 -21.350 378.155 -19.515 ;
        RECT 379.445 -19.920 379.675 -18.490 ;
        RECT 383.750 -18.960 385.420 -18.640 ;
        RECT 382.220 -19.520 384.760 -19.200 ;
        RECT 385.060 -19.225 385.420 -18.960 ;
        RECT 385.060 -19.495 386.090 -19.225 ;
        RECT 378.410 -20.150 379.675 -19.920 ;
        RECT 382.220 -20.080 385.630 -19.760 ;
        RECT 385.860 -20.320 386.090 -19.495 ;
        RECT 382.820 -20.640 386.090 -20.320 ;
        RECT 386.885 -19.515 388.160 -19.285 ;
        RECT 382.820 -21.340 383.180 -20.640 ;
        RECT 384.905 -21.340 385.135 -20.640 ;
        RECT 386.885 -21.350 387.115 -19.515 ;
        RECT 388.405 -19.920 388.635 -18.490 ;
        RECT 390.645 -19.010 390.875 -18.490 ;
        RECT 392.885 -19.010 393.115 -18.490 ;
        RECT 396.380 -18.720 404.420 -18.490 ;
        RECT 396.380 -18.825 396.610 -18.720 ;
        RECT 387.370 -20.150 388.635 -19.920 ;
        RECT 389.585 -19.280 393.115 -19.010 ;
        RECT 394.660 -19.055 396.610 -18.825 ;
        RECT 396.840 -19.180 403.080 -18.950 ;
        RECT 389.585 -20.760 389.855 -19.280 ;
        RECT 390.090 -20.110 391.000 -19.730 ;
        RECT 391.260 -20.110 393.000 -19.730 ;
        RECT 390.700 -20.340 391.000 -20.110 ;
        RECT 393.420 -20.340 393.670 -19.540 ;
        RECT 394.630 -20.110 396.610 -19.730 ;
        RECT 390.700 -20.660 393.670 -20.340 ;
        RECT 396.840 -20.490 397.160 -19.180 ;
        RECT 403.450 -19.410 404.460 -19.170 ;
        RECT 401.225 -19.625 404.460 -19.410 ;
        RECT 399.900 -19.640 404.460 -19.625 ;
        RECT 397.450 -20.080 398.280 -19.730 ;
        RECT 390.710 -20.670 390.970 -20.660 ;
        RECT 395.845 -20.720 397.680 -20.490 ;
        RECT 389.585 -20.910 390.385 -20.760 ;
        RECT 395.845 -20.850 396.075 -20.720 ;
        RECT 389.585 -20.995 390.470 -20.910 ;
        RECT 390.090 -21.100 390.470 -20.995 ;
        RECT 390.090 -21.170 392.090 -21.100 ;
        RECT 390.155 -21.330 392.090 -21.170 ;
        RECT 395.750 -21.230 396.075 -20.850 ;
        RECT 395.845 -21.335 396.075 -21.230 ;
        RECT 397.450 -21.120 397.680 -20.720 ;
        RECT 397.950 -20.655 398.280 -20.080 ;
        RECT 398.510 -20.110 399.470 -19.730 ;
        RECT 399.900 -19.945 401.455 -19.640 ;
        RECT 398.940 -20.195 399.470 -20.110 ;
        RECT 402.150 -20.195 402.830 -19.870 ;
        RECT 398.940 -20.425 402.830 -20.195 ;
        RECT 401.735 -20.650 402.830 -20.425 ;
        RECT 397.950 -20.880 401.330 -20.655 ;
        RECT 403.490 -20.880 403.720 -19.870 ;
        RECT 404.100 -20.240 404.460 -19.640 ;
        RECT 405.365 -19.515 406.640 -19.285 ;
        RECT 397.950 -20.890 403.720 -20.880 ;
        RECT 397.450 -21.350 400.830 -21.120 ;
        RECT 401.080 -21.220 403.720 -20.890 ;
        RECT 405.365 -21.350 405.595 -19.515 ;
        RECT 406.885 -19.920 407.115 -18.490 ;
        RECT 410.350 -19.010 410.690 -18.655 ;
        RECT 412.590 -19.010 412.930 -18.655 ;
        RECT 410.350 -19.245 412.930 -19.010 ;
        RECT 416.910 -18.845 417.255 -18.490 ;
        RECT 418.610 -18.845 420.030 -18.490 ;
        RECT 420.850 -18.845 422.270 -18.490 ;
        RECT 423.630 -18.845 424.015 -18.490 ;
        RECT 416.910 -19.075 424.015 -18.845 ;
        RECT 405.850 -20.150 407.115 -19.920 ;
        RECT 409.530 -20.150 410.600 -19.720 ;
        RECT 410.260 -21.350 410.600 -20.150 ;
        RECT 410.830 -21.350 411.170 -19.535 ;
        RECT 411.950 -21.350 412.290 -19.535 ;
        RECT 412.530 -21.350 412.930 -19.245 ;
        RECT 419.265 -19.550 421.775 -19.320 ;
        RECT 417.530 -20.340 417.910 -19.690 ;
        RECT 419.265 -19.730 419.535 -19.550 ;
        RECT 418.510 -20.110 419.535 -19.730 ;
        RECT 421.450 -19.730 421.775 -19.550 ;
        RECT 422.580 -19.625 423.455 -19.350 ;
        RECT 419.770 -20.055 421.205 -19.785 ;
        RECT 421.450 -20.055 422.225 -19.730 ;
        RECT 422.580 -20.340 422.855 -19.625 ;
        RECT 423.740 -19.980 424.015 -19.075 ;
        RECT 417.530 -20.615 422.855 -20.340 ;
        RECT 423.105 -20.210 424.015 -19.980 ;
        RECT 423.105 -20.900 423.335 -20.210 ;
        RECT 425.420 -20.670 425.755 -18.770 ;
        RECT 426.645 -19.515 427.920 -19.285 ;
        RECT 420.320 -21.195 423.335 -20.900 ;
        RECT 426.645 -21.350 426.875 -19.515 ;
        RECT 428.165 -19.920 428.395 -18.490 ;
        RECT 427.130 -20.150 428.395 -19.920 ;
        RECT 430.565 -20.480 430.795 -18.525 ;
        RECT 431.025 -19.700 431.400 -18.995 ;
        RECT 432.660 -19.565 433.250 -18.525 ;
        RECT 442.680 -18.720 446.030 -18.490 ;
        RECT 433.925 -19.240 434.155 -18.770 ;
        RECT 435.945 -19.055 436.450 -18.825 ;
        RECT 437.905 -19.035 438.310 -18.805 ;
        RECT 433.925 -19.470 435.715 -19.240 ;
        RECT 431.025 -20.110 431.910 -19.700 ;
        RECT 432.250 -20.480 432.590 -19.840 ;
        RECT 430.565 -20.715 432.590 -20.480 ;
        RECT 430.565 -21.340 430.895 -20.715 ;
        RECT 432.885 -21.280 433.250 -19.565 ;
        RECT 433.830 -20.110 435.250 -19.730 ;
        RECT 435.485 -20.365 435.715 -19.470 ;
        RECT 434.025 -20.595 435.715 -20.365 ;
        RECT 435.945 -20.345 436.175 -19.055 ;
        RECT 436.570 -20.110 437.600 -19.730 ;
        RECT 435.945 -20.575 437.575 -20.345 ;
        RECT 437.905 -20.380 438.135 -19.035 ;
        RECT 434.025 -21.185 434.255 -20.595 ;
        RECT 435.945 -21.175 436.295 -20.575 ;
        RECT 437.345 -20.950 437.575 -20.575 ;
        RECT 437.805 -20.720 438.135 -20.380 ;
        RECT 438.365 -20.950 438.595 -19.870 ;
        RECT 439.145 -20.030 439.375 -18.750 ;
        RECT 442.680 -19.110 442.910 -18.720 ;
        RECT 439.725 -19.340 442.910 -19.110 ;
        RECT 439.725 -19.550 439.955 -19.340 ;
        RECT 443.670 -19.570 444.010 -18.960 ;
        RECT 444.605 -19.550 444.835 -18.720 ;
        RECT 440.370 -19.800 444.350 -19.570 ;
        RECT 438.825 -20.260 443.835 -20.030 ;
        RECT 438.825 -20.720 439.055 -20.260 ;
        RECT 443.535 -20.485 443.835 -20.260 ;
        RECT 439.845 -20.720 442.675 -20.490 ;
        RECT 439.845 -20.915 440.075 -20.720 ;
        RECT 437.345 -21.180 438.595 -20.950 ;
        RECT 442.445 -21.090 442.675 -20.720 ;
        RECT 444.120 -20.805 444.350 -19.800 ;
        RECT 445.230 -19.780 445.570 -18.960 ;
        RECT 445.800 -19.320 446.030 -18.720 ;
        RECT 446.630 -19.090 447.435 -18.750 ;
        RECT 445.800 -19.550 446.800 -19.320 ;
        RECT 445.230 -20.010 446.120 -19.780 ;
        RECT 444.120 -21.035 444.760 -20.805 ;
        RECT 445.890 -21.120 446.120 -20.010 ;
        RECT 446.570 -20.485 446.800 -19.550 ;
        RECT 447.095 -20.890 447.435 -19.090 ;
        RECT 448.340 -18.980 449.975 -18.620 ;
        RECT 448.340 -19.790 448.885 -18.980 ;
        RECT 450.330 -19.410 450.560 -18.750 ;
        RECT 449.410 -19.640 451.910 -19.410 ;
        RECT 449.410 -20.135 449.640 -19.640 ;
        RECT 447.675 -20.365 449.640 -20.135 ;
        RECT 447.875 -21.010 449.145 -20.780 ;
        RECT 449.410 -20.890 449.640 -20.365 ;
        RECT 447.875 -21.120 448.105 -21.010 ;
        RECT 445.890 -21.350 448.105 -21.120 ;
        RECT 448.915 -21.120 449.145 -21.010 ;
        RECT 449.870 -21.120 450.100 -19.870 ;
        RECT 448.915 -21.350 450.100 -21.120 ;
        RECT 452.155 -21.340 452.590 -18.510 ;
        RECT 454.805 -19.560 455.430 -18.535 ;
        RECT 454.805 -21.340 455.275 -19.560 ;
        RECT 456.540 -19.590 457.055 -18.610 ;
        RECT 455.505 -20.540 455.790 -19.790 ;
        RECT 456.170 -20.150 457.055 -19.590 ;
        RECT 457.285 -20.540 457.515 -18.760 ;
        RECT 455.505 -20.775 457.515 -20.540 ;
        RECT 457.130 -21.350 457.515 -20.775 ;
        RECT 458.190 -19.565 458.780 -18.525 ;
        RECT 458.190 -21.280 458.555 -19.565 ;
        RECT 460.040 -19.700 460.415 -18.995 ;
        RECT 458.850 -20.480 459.190 -19.840 ;
        RECT 459.530 -20.110 460.415 -19.700 ;
        RECT 460.645 -20.480 460.875 -18.525 ;
        RECT 458.850 -20.715 460.875 -20.480 ;
        RECT 460.545 -21.340 460.875 -20.715 ;
        RECT 170.750 -22.950 171.130 -22.350 ;
        RECT 172.990 -22.950 173.370 -22.350 ;
        RECT 175.230 -22.950 175.610 -22.350 ;
        RECT 177.470 -22.950 177.850 -22.350 ;
        RECT 180.830 -22.950 181.210 -22.350 ;
        RECT 183.070 -22.950 183.450 -22.350 ;
        RECT 185.310 -22.950 185.690 -22.350 ;
        RECT 187.550 -22.950 187.930 -22.350 ;
        RECT 170.750 -23.250 189.320 -22.950 ;
        RECT 298.905 -23.090 299.135 -22.420 ;
        RECT 301.145 -23.090 301.375 -22.420 ;
        RECT 303.385 -23.090 303.615 -22.420 ;
        RECT 305.525 -23.090 305.755 -22.420 ;
        RECT 307.865 -23.040 308.095 -22.420 ;
        RECT 310.105 -23.040 310.335 -22.420 ;
        RECT 171.870 -24.950 172.250 -24.350 ;
        RECT 176.350 -24.950 176.730 -24.350 ;
        RECT 181.950 -24.950 182.330 -24.350 ;
        RECT 186.430 -24.950 186.810 -24.350 ;
        RECT 166.590 -25.250 186.810 -24.950 ;
        RECT 166.590 -30.510 166.890 -25.250 ;
        RECT 174.110 -26.950 174.490 -26.350 ;
        RECT 184.190 -26.950 184.570 -26.350 ;
        RECT 173.390 -27.250 184.570 -26.950 ;
        RECT 173.390 -30.510 173.690 -27.250 ;
        RECT 178.355 -29.640 178.970 -28.740 ;
        RECT 179.710 -29.640 180.255 -28.740 ;
        RECT 166.590 -30.810 170.020 -30.510 ;
        RECT 166.590 -33.790 166.820 -30.810 ;
        RECT 168.190 -33.790 168.420 -30.810 ;
        RECT 169.790 -33.790 170.020 -30.810 ;
        RECT 173.390 -30.810 175.220 -30.510 ;
        RECT 173.390 -33.790 173.620 -30.810 ;
        RECT 174.990 -33.790 175.220 -30.810 ;
        RECT 178.355 -33.790 178.655 -29.640 ;
        RECT 179.955 -33.790 180.255 -29.640 ;
        RECT 189.020 -30.510 189.320 -23.250 ;
        RECT 298.870 -23.470 305.755 -23.090 ;
        RECT 307.285 -23.270 310.335 -23.040 ;
        RECT 298.060 -24.115 301.260 -23.770 ;
        RECT 301.960 -24.380 302.760 -23.470 ;
        RECT 307.285 -23.775 307.620 -23.270 ;
        RECT 303.330 -24.115 307.620 -23.775 ;
        RECT 308.090 -24.085 310.950 -23.650 ;
        RECT 298.805 -24.760 305.755 -24.380 ;
        RECT 298.805 -25.125 299.035 -24.760 ;
        RECT 301.045 -25.125 301.275 -24.760 ;
        RECT 303.285 -25.125 303.515 -24.760 ;
        RECT 305.495 -25.125 305.755 -24.760 ;
        RECT 307.285 -24.550 307.620 -24.115 ;
        RECT 312.005 -24.200 312.475 -22.420 ;
        RECT 314.330 -22.985 314.715 -22.410 ;
        RECT 312.705 -23.220 314.715 -22.985 ;
        RECT 312.705 -23.970 312.990 -23.220 ;
        RECT 313.370 -24.170 314.255 -23.610 ;
        RECT 307.285 -24.785 310.235 -24.550 ;
        RECT 307.765 -25.125 307.995 -24.785 ;
        RECT 310.005 -25.125 310.235 -24.785 ;
        RECT 312.005 -25.225 312.630 -24.200 ;
        RECT 313.740 -25.150 314.255 -24.170 ;
        RECT 314.485 -25.000 314.715 -23.220 ;
        RECT 316.885 -24.245 317.115 -22.410 ;
        RECT 319.575 -23.120 319.855 -22.420 ;
        RECT 319.575 -23.150 321.000 -23.120 ;
        RECT 319.530 -23.410 321.000 -23.150 ;
        RECT 319.575 -23.440 321.000 -23.410 ;
        RECT 317.370 -23.840 318.635 -23.610 ;
        RECT 316.885 -24.475 318.160 -24.245 ;
        RECT 318.405 -25.270 318.635 -23.840 ;
        RECT 319.385 -24.010 320.415 -23.670 ;
        RECT 320.110 -25.200 320.415 -24.010 ;
        RECT 320.645 -25.200 321.000 -23.440 ;
        RECT 321.230 -24.620 321.535 -22.480 ;
        RECT 322.485 -24.245 322.715 -22.410 ;
        RECT 322.970 -23.840 324.235 -23.610 ;
        RECT 322.485 -24.475 323.760 -24.245 ;
        RECT 324.005 -25.270 324.235 -23.840 ;
        RECT 324.725 -24.245 324.955 -22.410 ;
        RECT 325.210 -23.840 326.475 -23.610 ;
        RECT 324.725 -24.475 326.000 -24.245 ;
        RECT 326.245 -25.270 326.475 -23.840 ;
        RECT 326.965 -24.245 327.195 -22.410 ;
        RECT 327.450 -23.840 328.715 -23.610 ;
        RECT 326.965 -24.475 328.240 -24.245 ;
        RECT 328.485 -25.270 328.715 -23.840 ;
        RECT 329.205 -24.245 329.435 -22.410 ;
        RECT 329.690 -23.840 330.955 -23.610 ;
        RECT 329.205 -24.475 330.480 -24.245 ;
        RECT 330.725 -25.270 330.955 -23.840 ;
        RECT 331.445 -24.245 331.675 -22.410 ;
        RECT 331.930 -23.840 333.195 -23.610 ;
        RECT 331.445 -24.475 332.720 -24.245 ;
        RECT 332.965 -25.270 333.195 -23.840 ;
        RECT 333.685 -24.245 333.915 -22.410 ;
        RECT 334.170 -23.840 335.435 -23.610 ;
        RECT 333.685 -24.475 334.960 -24.245 ;
        RECT 335.205 -25.270 335.435 -23.840 ;
        RECT 335.925 -24.245 336.155 -22.410 ;
        RECT 336.410 -23.840 337.675 -23.610 ;
        RECT 335.925 -24.475 337.200 -24.245 ;
        RECT 337.445 -25.270 337.675 -23.840 ;
        RECT 338.165 -24.245 338.395 -22.410 ;
        RECT 338.650 -23.840 339.915 -23.610 ;
        RECT 338.165 -24.475 339.440 -24.245 ;
        RECT 339.685 -25.270 339.915 -23.840 ;
        RECT 340.405 -24.245 340.635 -22.410 ;
        RECT 340.890 -23.840 342.155 -23.610 ;
        RECT 340.405 -24.475 341.680 -24.245 ;
        RECT 341.925 -25.270 342.155 -23.840 ;
        RECT 343.365 -24.200 343.835 -22.420 ;
        RECT 345.690 -22.985 346.075 -22.410 ;
        RECT 344.065 -23.220 346.075 -22.985 ;
        RECT 344.065 -23.970 344.350 -23.220 ;
        RECT 344.730 -24.170 345.615 -23.610 ;
        RECT 343.365 -25.225 343.990 -24.200 ;
        RECT 345.100 -25.150 345.615 -24.170 ;
        RECT 345.845 -25.000 346.075 -23.220 ;
        RECT 346.565 -24.245 346.795 -22.410 ;
        RECT 347.050 -23.840 348.315 -23.610 ;
        RECT 346.565 -24.475 347.840 -24.245 ;
        RECT 348.085 -25.270 348.315 -23.840 ;
        RECT 348.805 -24.245 349.035 -22.410 ;
        RECT 349.290 -23.840 350.555 -23.610 ;
        RECT 348.805 -24.475 350.080 -24.245 ;
        RECT 350.325 -25.270 350.555 -23.840 ;
        RECT 351.500 -24.990 351.835 -23.090 ;
        RECT 353.185 -24.830 353.510 -22.850 ;
        RECT 353.740 -25.200 354.075 -22.430 ;
        RECT 356.545 -24.190 356.870 -22.480 ;
        RECT 357.160 -22.660 360.205 -22.430 ;
        RECT 357.160 -24.705 357.390 -22.660 ;
        RECT 357.640 -23.610 358.000 -22.955 ;
        RECT 358.280 -23.120 359.675 -22.890 ;
        RECT 357.640 -24.115 358.555 -23.610 ;
        RECT 356.085 -24.935 358.555 -24.705 ;
        RECT 356.085 -25.250 356.315 -24.935 ;
        RECT 358.325 -25.250 358.555 -24.935 ;
        RECT 358.785 -25.250 359.080 -23.580 ;
        RECT 359.320 -25.250 359.675 -23.120 ;
        RECT 359.975 -23.120 360.205 -22.660 ;
        RECT 359.975 -23.350 360.795 -23.120 ;
        RECT 359.905 -25.250 360.220 -23.580 ;
        RECT 360.565 -25.250 360.795 -23.350 ;
        RECT 362.740 -23.500 362.970 -22.420 ;
        RECT 365.100 -22.640 373.650 -22.410 ;
        RECT 373.310 -22.745 373.650 -22.640 ;
        RECT 383.765 -22.745 383.995 -22.420 ;
        RECT 373.310 -22.975 383.995 -22.745 ;
        RECT 361.560 -23.730 362.970 -23.500 ;
        RECT 365.220 -23.440 372.580 -23.120 ;
        RECT 373.310 -23.270 373.650 -22.975 ;
        RECT 374.580 -23.440 383.040 -23.205 ;
        RECT 383.765 -23.270 383.995 -22.975 ;
        RECT 385.805 -22.640 388.125 -22.410 ;
        RECT 361.560 -25.270 361.950 -23.730 ;
        RECT 362.185 -24.360 363.000 -23.980 ;
        RECT 362.635 -25.245 363.000 -24.360 ;
        RECT 363.240 -24.740 363.605 -23.610 ;
        RECT 365.220 -24.615 365.450 -23.440 ;
        RECT 374.580 -23.680 374.810 -23.440 ;
        RECT 365.680 -24.000 373.275 -23.680 ;
        RECT 373.790 -24.000 374.810 -23.680 ;
        RECT 377.770 -23.835 378.110 -23.440 ;
        RECT 379.445 -23.835 379.785 -23.440 ;
        RECT 380.320 -24.065 382.490 -23.670 ;
        RECT 382.810 -23.680 383.040 -23.440 ;
        RECT 385.805 -23.440 386.035 -22.640 ;
        RECT 386.265 -23.210 387.650 -22.870 ;
        RECT 382.810 -24.000 383.830 -23.680 ;
        RECT 384.530 -23.900 385.505 -23.650 ;
        RECT 385.805 -23.670 386.395 -23.440 ;
        RECT 365.950 -24.460 372.175 -24.230 ;
        RECT 375.080 -24.295 382.490 -24.065 ;
        RECT 384.530 -24.200 385.935 -23.900 ;
        RECT 365.950 -24.590 368.070 -24.460 ;
        RECT 365.220 -24.770 365.660 -24.615 ;
        RECT 372.745 -24.700 382.980 -24.525 ;
        RECT 368.720 -24.755 382.980 -24.700 ;
        RECT 365.220 -24.845 365.770 -24.770 ;
        RECT 365.430 -24.870 365.770 -24.845 ;
        RECT 368.720 -24.870 372.975 -24.755 ;
        RECT 365.430 -24.930 372.975 -24.870 ;
        RECT 365.430 -25.100 368.950 -24.930 ;
        RECT 365.510 -25.150 365.770 -25.100 ;
        RECT 367.140 -25.270 367.480 -25.100 ;
        RECT 371.220 -25.225 371.560 -24.930 ;
        RECT 374.600 -25.025 374.940 -24.755 ;
        RECT 377.280 -25.025 377.620 -24.755 ;
        RECT 379.960 -25.025 380.300 -24.755 ;
        RECT 382.640 -25.025 382.980 -24.755 ;
        RECT 385.600 -25.250 385.935 -24.200 ;
        RECT 386.165 -25.250 386.395 -23.670 ;
        RECT 386.720 -25.250 387.055 -23.480 ;
        RECT 387.285 -25.250 387.650 -23.210 ;
        RECT 387.895 -23.110 388.125 -22.640 ;
        RECT 387.895 -23.340 388.635 -23.110 ;
        RECT 387.880 -25.250 388.175 -23.570 ;
        RECT 388.405 -25.250 388.635 -23.340 ;
        RECT 390.645 -24.990 390.980 -23.090 ;
        RECT 392.380 -24.990 392.715 -23.090 ;
        RECT 395.285 -24.245 395.515 -22.410 ;
        RECT 395.770 -23.840 397.035 -23.610 ;
        RECT 395.285 -24.475 396.560 -24.245 ;
        RECT 392.390 -25.150 392.650 -24.990 ;
        RECT 396.805 -25.270 397.035 -23.840 ;
        RECT 397.525 -24.245 397.755 -22.410 ;
        RECT 399.865 -23.165 400.095 -22.575 ;
        RECT 399.865 -23.395 401.555 -23.165 ;
        RECT 398.010 -23.840 399.275 -23.610 ;
        RECT 397.525 -24.475 398.800 -24.245 ;
        RECT 399.045 -25.270 399.275 -23.840 ;
        RECT 399.670 -24.030 401.090 -23.650 ;
        RECT 401.325 -24.290 401.555 -23.395 ;
        RECT 399.765 -24.520 401.555 -24.290 ;
        RECT 401.785 -23.185 402.135 -22.585 ;
        RECT 403.185 -22.810 404.435 -22.580 ;
        RECT 411.730 -22.640 413.945 -22.410 ;
        RECT 403.185 -23.185 403.415 -22.810 ;
        RECT 401.785 -23.415 403.415 -23.185 ;
        RECT 403.645 -23.380 403.975 -23.040 ;
        RECT 399.765 -24.990 399.995 -24.520 ;
        RECT 401.785 -24.705 402.015 -23.415 ;
        RECT 402.410 -24.030 403.440 -23.650 ;
        RECT 401.785 -24.935 402.290 -24.705 ;
        RECT 403.745 -24.725 403.975 -23.380 ;
        RECT 404.205 -23.890 404.435 -22.810 ;
        RECT 405.685 -23.040 405.915 -22.845 ;
        RECT 408.285 -23.040 408.515 -22.670 ;
        RECT 404.665 -23.500 404.895 -23.040 ;
        RECT 405.685 -23.270 408.515 -23.040 ;
        RECT 409.960 -22.955 410.600 -22.725 ;
        RECT 409.375 -23.500 409.675 -23.275 ;
        RECT 404.665 -23.730 409.675 -23.500 ;
        RECT 403.745 -24.955 404.150 -24.725 ;
        RECT 404.985 -25.010 405.215 -23.730 ;
        RECT 409.960 -23.960 410.190 -22.955 ;
        RECT 411.730 -23.750 411.960 -22.640 ;
        RECT 413.715 -22.750 413.945 -22.640 ;
        RECT 414.755 -22.640 415.940 -22.410 ;
        RECT 414.755 -22.750 414.985 -22.640 ;
        RECT 406.210 -24.190 410.190 -23.960 ;
        RECT 411.070 -23.980 411.960 -23.750 ;
        RECT 405.565 -24.420 405.795 -24.210 ;
        RECT 405.565 -24.650 408.750 -24.420 ;
        RECT 408.520 -25.040 408.750 -24.650 ;
        RECT 409.510 -24.800 409.850 -24.190 ;
        RECT 410.445 -25.040 410.675 -24.210 ;
        RECT 411.070 -24.800 411.410 -23.980 ;
        RECT 412.410 -24.210 412.640 -23.275 ;
        RECT 411.640 -24.440 412.640 -24.210 ;
        RECT 411.640 -25.040 411.870 -24.440 ;
        RECT 412.935 -24.670 413.275 -22.870 ;
        RECT 413.715 -22.980 414.985 -22.750 ;
        RECT 415.250 -23.395 415.480 -22.870 ;
        RECT 413.515 -23.625 415.480 -23.395 ;
        RECT 412.470 -25.010 413.275 -24.670 ;
        RECT 414.180 -24.780 414.725 -23.970 ;
        RECT 415.250 -24.120 415.480 -23.625 ;
        RECT 415.710 -23.890 415.940 -22.640 ;
        RECT 415.250 -24.350 417.750 -24.120 ;
        RECT 408.520 -25.270 411.870 -25.040 ;
        RECT 414.180 -25.140 415.815 -24.780 ;
        RECT 416.170 -25.010 416.400 -24.350 ;
        RECT 417.995 -25.250 418.430 -22.420 ;
        RECT 418.750 -22.640 421.130 -22.410 ;
        RECT 418.750 -23.305 419.090 -22.640 ;
        RECT 418.675 -24.030 419.570 -23.650 ;
        RECT 419.220 -24.640 419.570 -24.030 ;
        RECT 419.800 -24.930 420.105 -23.075 ;
        RECT 420.790 -23.305 421.130 -22.640 ;
        RECT 420.335 -24.030 421.240 -23.650 ;
        RECT 421.470 -24.030 422.375 -23.650 ;
        RECT 420.900 -24.640 421.240 -24.030 ;
        RECT 422.035 -24.640 422.375 -24.030 ;
        RECT 420.390 -24.930 420.650 -24.770 ;
        RECT 419.800 -25.250 421.140 -24.930 ;
        RECT 424.300 -24.990 424.635 -23.090 ;
        RECT 425.525 -24.245 425.755 -22.410 ;
        RECT 426.010 -23.840 427.275 -23.610 ;
        RECT 425.525 -24.475 426.800 -24.245 ;
        RECT 427.045 -25.270 427.275 -23.840 ;
        RECT 427.765 -24.245 427.995 -22.410 ;
        RECT 428.250 -23.840 429.515 -23.610 ;
        RECT 427.765 -24.475 429.040 -24.245 ;
        RECT 429.285 -25.270 429.515 -23.840 ;
        RECT 430.005 -24.245 430.235 -22.410 ;
        RECT 430.490 -23.840 431.755 -23.610 ;
        RECT 430.005 -24.475 431.280 -24.245 ;
        RECT 431.525 -25.270 431.755 -23.840 ;
        RECT 435.490 -25.260 435.890 -22.420 ;
        RECT 436.185 -24.485 436.415 -24.020 ;
        RECT 437.120 -24.255 437.470 -22.515 ;
        RECT 437.700 -22.835 439.500 -22.605 ;
        RECT 437.700 -24.485 437.930 -22.835 ;
        RECT 441.905 -23.075 442.290 -22.410 ;
        RECT 438.560 -23.310 442.290 -23.075 ;
        RECT 438.560 -23.840 438.900 -23.310 ;
        RECT 439.150 -23.990 441.610 -23.605 ;
        RECT 439.150 -24.150 439.460 -23.990 ;
        RECT 436.185 -24.715 437.930 -24.485 ;
        RECT 438.160 -24.550 439.460 -24.150 ;
        RECT 439.815 -24.550 441.465 -24.220 ;
        RECT 437.700 -25.020 437.930 -24.715 ;
        RECT 437.700 -25.250 439.060 -25.020 ;
        RECT 441.950 -25.260 442.290 -23.310 ;
        RECT 443.630 -24.195 443.995 -22.480 ;
        RECT 445.985 -23.045 446.315 -22.420 ;
        RECT 444.290 -23.280 446.315 -23.045 ;
        RECT 447.825 -23.040 448.055 -22.420 ;
        RECT 450.065 -23.040 450.295 -22.420 ;
        RECT 447.825 -23.270 450.875 -23.040 ;
        RECT 444.290 -23.920 444.630 -23.280 ;
        RECT 444.970 -24.060 445.855 -23.650 ;
        RECT 443.630 -25.235 444.220 -24.195 ;
        RECT 445.480 -24.765 445.855 -24.060 ;
        RECT 446.085 -25.235 446.315 -23.280 ;
        RECT 447.210 -24.085 450.070 -23.650 ;
        RECT 450.540 -23.775 450.875 -23.270 ;
        RECT 452.405 -23.090 452.635 -22.420 ;
        RECT 454.545 -23.090 454.775 -22.420 ;
        RECT 456.785 -23.090 457.015 -22.420 ;
        RECT 459.025 -22.530 459.255 -22.420 ;
        RECT 459.025 -22.910 459.290 -22.530 ;
        RECT 459.025 -23.090 459.255 -22.910 ;
        RECT 452.405 -23.470 459.255 -23.090 ;
        RECT 450.540 -24.115 454.830 -23.775 ;
        RECT 450.540 -24.550 450.875 -24.115 ;
        RECT 455.400 -24.380 456.200 -23.470 ;
        RECT 456.900 -24.115 460.100 -23.770 ;
        RECT 447.925 -24.785 450.875 -24.550 ;
        RECT 452.405 -24.760 459.355 -24.380 ;
        RECT 447.925 -25.125 448.155 -24.785 ;
        RECT 450.165 -25.125 450.395 -24.785 ;
        RECT 452.405 -25.125 452.665 -24.760 ;
        RECT 454.645 -25.125 454.875 -24.760 ;
        RECT 456.885 -25.125 457.115 -24.760 ;
        RECT 459.125 -25.125 459.355 -24.760 ;
        RECT 307.160 -26.560 310.510 -26.330 ;
        RECT 298.405 -27.080 298.635 -26.610 ;
        RECT 300.425 -26.895 300.930 -26.665 ;
        RECT 302.385 -26.875 302.790 -26.645 ;
        RECT 298.405 -27.310 300.195 -27.080 ;
        RECT 298.440 -27.950 299.730 -27.570 ;
        RECT 299.965 -28.205 300.195 -27.310 ;
        RECT 298.505 -28.435 300.195 -28.205 ;
        RECT 300.425 -28.185 300.655 -26.895 ;
        RECT 301.050 -27.950 302.080 -27.570 ;
        RECT 300.425 -28.415 302.055 -28.185 ;
        RECT 302.385 -28.220 302.615 -26.875 ;
        RECT 298.505 -29.025 298.735 -28.435 ;
        RECT 300.425 -29.015 300.775 -28.415 ;
        RECT 301.825 -28.790 302.055 -28.415 ;
        RECT 302.285 -28.560 302.615 -28.220 ;
        RECT 302.845 -28.790 303.075 -27.710 ;
        RECT 303.625 -27.870 303.855 -26.590 ;
        RECT 307.160 -26.950 307.390 -26.560 ;
        RECT 304.205 -27.180 307.390 -26.950 ;
        RECT 304.205 -27.390 304.435 -27.180 ;
        RECT 308.150 -27.410 308.490 -26.800 ;
        RECT 309.085 -27.390 309.315 -26.560 ;
        RECT 304.850 -27.640 308.830 -27.410 ;
        RECT 303.305 -28.100 308.315 -27.870 ;
        RECT 303.305 -28.560 303.535 -28.100 ;
        RECT 308.015 -28.325 308.315 -28.100 ;
        RECT 304.325 -28.560 307.155 -28.330 ;
        RECT 304.325 -28.755 304.555 -28.560 ;
        RECT 301.825 -29.020 303.075 -28.790 ;
        RECT 306.925 -28.930 307.155 -28.560 ;
        RECT 308.600 -28.645 308.830 -27.640 ;
        RECT 309.710 -27.620 310.050 -26.800 ;
        RECT 310.280 -27.160 310.510 -26.560 ;
        RECT 311.110 -26.930 311.915 -26.590 ;
        RECT 310.280 -27.390 311.280 -27.160 ;
        RECT 309.710 -27.850 310.600 -27.620 ;
        RECT 308.600 -28.875 309.240 -28.645 ;
        RECT 310.370 -28.960 310.600 -27.850 ;
        RECT 311.050 -28.325 311.280 -27.390 ;
        RECT 311.575 -28.730 311.915 -26.930 ;
        RECT 312.820 -26.820 314.455 -26.460 ;
        RECT 312.820 -27.630 313.365 -26.820 ;
        RECT 314.810 -27.250 315.040 -26.590 ;
        RECT 313.890 -27.480 316.390 -27.250 ;
        RECT 313.890 -27.975 314.120 -27.480 ;
        RECT 312.155 -28.205 314.120 -27.975 ;
        RECT 312.355 -28.850 313.625 -28.620 ;
        RECT 313.890 -28.730 314.120 -28.205 ;
        RECT 312.355 -28.960 312.585 -28.850 ;
        RECT 310.370 -29.190 312.585 -28.960 ;
        RECT 313.395 -28.960 313.625 -28.850 ;
        RECT 314.350 -28.960 314.580 -27.710 ;
        RECT 313.395 -29.190 314.580 -28.960 ;
        RECT 316.635 -29.180 317.070 -26.350 ;
        RECT 319.100 -26.670 320.440 -26.350 ;
        RECT 319.590 -26.830 319.850 -26.670 ;
        RECT 317.865 -27.570 318.205 -26.960 ;
        RECT 319.000 -27.570 319.340 -26.960 ;
        RECT 317.865 -27.950 318.770 -27.570 ;
        RECT 319.000 -27.950 319.905 -27.570 ;
        RECT 319.110 -28.960 319.450 -28.295 ;
        RECT 320.135 -28.525 320.440 -26.670 ;
        RECT 322.030 -26.840 322.795 -26.410 ;
        RECT 320.670 -27.570 321.020 -26.960 ;
        RECT 320.670 -27.950 321.565 -27.570 ;
        RECT 322.030 -28.090 322.360 -26.840 ;
        RECT 324.455 -27.080 324.850 -26.330 ;
        RECT 322.625 -27.310 324.850 -27.080 ;
        RECT 322.625 -27.440 323.480 -27.310 ;
        RECT 321.150 -28.960 321.490 -28.295 ;
        RECT 319.110 -29.190 321.490 -28.960 ;
        RECT 322.030 -29.145 322.660 -28.090 ;
        RECT 324.020 -29.145 324.380 -27.540 ;
        RECT 324.620 -28.930 324.850 -27.310 ;
        RECT 325.080 -28.680 325.500 -26.875 ;
        RECT 326.405 -27.355 327.680 -27.125 ;
        RECT 324.620 -29.160 325.825 -28.930 ;
        RECT 326.405 -29.190 326.635 -27.355 ;
        RECT 327.925 -27.760 328.155 -26.330 ;
        RECT 326.890 -27.990 328.155 -27.760 ;
        RECT 328.645 -27.355 329.920 -27.125 ;
        RECT 328.645 -29.190 328.875 -27.355 ;
        RECT 330.165 -27.760 330.395 -26.330 ;
        RECT 329.130 -27.990 330.395 -27.760 ;
        RECT 330.885 -27.355 332.160 -27.125 ;
        RECT 330.885 -29.190 331.115 -27.355 ;
        RECT 332.405 -27.760 332.635 -26.330 ;
        RECT 331.370 -27.990 332.635 -27.760 ;
        RECT 333.125 -27.355 334.400 -27.125 ;
        RECT 333.125 -29.190 333.355 -27.355 ;
        RECT 334.645 -27.760 334.875 -26.330 ;
        RECT 333.610 -27.990 334.875 -27.760 ;
        RECT 336.485 -27.355 337.760 -27.125 ;
        RECT 336.485 -29.190 336.715 -27.355 ;
        RECT 338.005 -27.760 338.235 -26.330 ;
        RECT 336.970 -27.990 338.235 -27.760 ;
        RECT 338.725 -27.355 340.000 -27.125 ;
        RECT 338.725 -29.190 338.955 -27.355 ;
        RECT 340.245 -27.760 340.475 -26.330 ;
        RECT 339.210 -27.990 340.475 -27.760 ;
        RECT 340.965 -27.355 342.240 -27.125 ;
        RECT 340.965 -29.190 341.195 -27.355 ;
        RECT 342.485 -27.760 342.715 -26.330 ;
        RECT 341.450 -27.990 342.715 -27.760 ;
        RECT 343.205 -27.355 344.480 -27.125 ;
        RECT 343.205 -29.190 343.435 -27.355 ;
        RECT 344.725 -27.760 344.955 -26.330 ;
        RECT 343.690 -27.990 344.955 -27.760 ;
        RECT 345.445 -27.355 346.720 -27.125 ;
        RECT 345.445 -29.190 345.675 -27.355 ;
        RECT 346.965 -27.760 347.195 -26.330 ;
        RECT 345.930 -27.990 347.195 -27.760 ;
        RECT 349.265 -28.750 349.590 -26.770 ;
        RECT 349.820 -29.170 350.155 -26.400 ;
        RECT 351.605 -26.665 351.835 -26.350 ;
        RECT 353.845 -26.665 354.075 -26.350 ;
        RECT 351.605 -26.895 354.075 -26.665 ;
        RECT 352.065 -29.120 352.390 -27.410 ;
        RECT 352.680 -28.940 352.910 -26.895 ;
        RECT 353.160 -27.990 354.075 -27.485 ;
        RECT 353.160 -28.645 353.520 -27.990 ;
        RECT 354.305 -28.020 354.600 -26.350 ;
        RECT 354.840 -28.480 355.195 -26.350 ;
        RECT 355.425 -28.020 355.740 -26.350 ;
        RECT 356.085 -28.250 356.315 -26.350 ;
        RECT 353.800 -28.710 355.195 -28.480 ;
        RECT 355.495 -28.480 356.315 -28.250 ;
        RECT 357.205 -27.355 358.480 -27.125 ;
        RECT 355.495 -28.940 355.725 -28.480 ;
        RECT 352.680 -29.170 355.725 -28.940 ;
        RECT 357.205 -29.190 357.435 -27.355 ;
        RECT 358.725 -27.760 358.955 -26.330 ;
        RECT 357.690 -27.990 358.955 -27.760 ;
        RECT 359.445 -27.355 360.720 -27.125 ;
        RECT 359.445 -29.190 359.675 -27.355 ;
        RECT 360.965 -27.760 361.195 -26.330 ;
        RECT 359.930 -27.990 361.195 -27.760 ;
        RECT 361.685 -27.355 362.960 -27.125 ;
        RECT 361.685 -29.190 361.915 -27.355 ;
        RECT 363.205 -27.760 363.435 -26.330 ;
        RECT 362.170 -27.990 363.435 -27.760 ;
        RECT 364.645 -27.400 365.270 -26.375 ;
        RECT 364.645 -29.180 365.115 -27.400 ;
        RECT 366.380 -27.430 366.895 -26.450 ;
        RECT 365.345 -28.380 365.630 -27.630 ;
        RECT 366.010 -27.990 366.895 -27.430 ;
        RECT 367.125 -28.380 367.355 -26.600 ;
        RECT 365.345 -28.615 367.355 -28.380 ;
        RECT 366.970 -29.190 367.355 -28.615 ;
        RECT 367.845 -27.355 369.120 -27.125 ;
        RECT 367.845 -29.190 368.075 -27.355 ;
        RECT 369.365 -27.760 369.595 -26.330 ;
        RECT 368.330 -27.990 369.595 -27.760 ;
        RECT 370.085 -27.355 371.360 -27.125 ;
        RECT 370.085 -29.190 370.315 -27.355 ;
        RECT 371.605 -27.760 371.835 -26.330 ;
        RECT 370.570 -27.990 371.835 -27.760 ;
        RECT 372.325 -27.355 373.600 -27.125 ;
        RECT 372.325 -29.190 372.555 -27.355 ;
        RECT 373.845 -27.760 374.075 -26.330 ;
        RECT 372.810 -27.990 374.075 -27.760 ;
        RECT 375.845 -27.400 376.470 -26.375 ;
        RECT 375.845 -29.180 376.315 -27.400 ;
        RECT 377.580 -27.430 378.095 -26.450 ;
        RECT 376.545 -28.380 376.830 -27.630 ;
        RECT 377.210 -27.990 378.095 -27.430 ;
        RECT 378.325 -28.380 378.555 -26.600 ;
        RECT 376.545 -28.615 378.555 -28.380 ;
        RECT 378.170 -29.190 378.555 -28.615 ;
        RECT 379.045 -27.355 380.320 -27.125 ;
        RECT 379.045 -29.190 379.275 -27.355 ;
        RECT 380.565 -27.760 380.795 -26.330 ;
        RECT 379.530 -27.990 380.795 -27.760 ;
        RECT 381.285 -27.355 382.560 -27.125 ;
        RECT 381.285 -29.190 381.515 -27.355 ;
        RECT 382.805 -27.760 383.035 -26.330 ;
        RECT 384.865 -27.080 385.095 -26.600 ;
        RECT 381.770 -27.990 383.035 -27.760 ;
        RECT 383.950 -27.310 385.095 -27.080 ;
        RECT 383.950 -28.160 384.290 -27.310 ;
        RECT 386.680 -27.540 387.055 -26.350 ;
        RECT 384.550 -27.840 385.870 -27.540 ;
        RECT 383.950 -28.510 385.095 -28.160 ;
        RECT 384.865 -29.190 385.095 -28.510 ;
        RECT 385.545 -28.390 385.870 -27.840 ;
        RECT 386.110 -27.950 387.055 -27.540 ;
        RECT 387.285 -28.390 387.515 -26.605 ;
        RECT 385.545 -28.620 387.515 -28.390 ;
        RECT 387.285 -29.190 387.515 -28.620 ;
        RECT 388.005 -27.355 389.280 -27.125 ;
        RECT 388.005 -29.190 388.235 -27.355 ;
        RECT 389.525 -27.760 389.755 -26.330 ;
        RECT 388.490 -27.990 389.755 -27.760 ;
        RECT 390.245 -27.355 391.520 -27.125 ;
        RECT 390.245 -29.190 390.475 -27.355 ;
        RECT 391.765 -27.760 391.995 -26.330 ;
        RECT 390.730 -27.990 391.995 -27.760 ;
        RECT 392.485 -27.355 393.760 -27.125 ;
        RECT 392.485 -29.190 392.715 -27.355 ;
        RECT 394.005 -27.760 394.235 -26.330 ;
        RECT 392.970 -27.990 394.235 -27.760 ;
        RECT 395.115 -27.990 395.480 -26.860 ;
        RECT 395.720 -27.240 396.085 -26.355 ;
        RECT 395.720 -27.620 396.535 -27.240 ;
        RECT 396.770 -27.870 397.160 -26.330 ;
        RECT 395.750 -28.100 397.160 -27.870 ;
        RECT 397.525 -27.355 398.800 -27.125 ;
        RECT 395.750 -29.180 395.980 -28.100 ;
        RECT 397.525 -29.190 397.755 -27.355 ;
        RECT 399.045 -27.760 399.275 -26.330 ;
        RECT 401.320 -26.670 402.660 -26.350 ;
        RECT 400.740 -27.570 401.090 -26.960 ;
        RECT 398.010 -27.990 399.275 -27.760 ;
        RECT 400.195 -27.950 401.090 -27.570 ;
        RECT 400.270 -28.960 400.610 -28.295 ;
        RECT 401.320 -28.525 401.625 -26.670 ;
        RECT 401.910 -26.830 402.170 -26.670 ;
        RECT 402.420 -27.570 402.760 -26.960 ;
        RECT 403.555 -27.570 403.895 -26.960 ;
        RECT 401.855 -27.950 402.760 -27.570 ;
        RECT 402.990 -27.950 403.895 -27.570 ;
        RECT 402.310 -28.960 402.650 -28.295 ;
        RECT 400.270 -29.190 402.650 -28.960 ;
        RECT 405.205 -29.170 405.540 -26.400 ;
        RECT 405.770 -28.750 406.095 -26.770 ;
        RECT 407.045 -27.355 408.320 -27.125 ;
        RECT 407.045 -29.190 407.275 -27.355 ;
        RECT 408.565 -27.760 408.795 -26.330 ;
        RECT 407.530 -27.990 408.795 -27.760 ;
        RECT 409.285 -27.355 410.560 -27.125 ;
        RECT 409.285 -29.190 409.515 -27.355 ;
        RECT 410.805 -27.760 411.035 -26.330 ;
        RECT 409.770 -27.990 411.035 -27.760 ;
        RECT 411.525 -27.355 412.800 -27.125 ;
        RECT 411.525 -29.190 411.755 -27.355 ;
        RECT 413.045 -27.760 413.275 -26.330 ;
        RECT 412.010 -27.990 413.275 -27.760 ;
        RECT 414.885 -27.355 416.160 -27.125 ;
        RECT 414.885 -29.190 415.115 -27.355 ;
        RECT 416.405 -27.760 416.635 -26.330 ;
        RECT 418.150 -26.610 418.410 -26.450 ;
        RECT 415.370 -27.990 416.635 -27.760 ;
        RECT 418.085 -28.510 418.420 -26.610 ;
        RECT 419.820 -28.510 420.155 -26.610 ;
        RECT 422.020 -27.560 422.425 -26.855 ;
        RECT 421.480 -27.950 422.425 -27.560 ;
        RECT 423.140 -27.760 423.500 -26.350 ;
        RECT 424.260 -27.760 424.570 -26.350 ;
        RECT 424.800 -28.160 425.030 -26.455 ;
        RECT 422.760 -28.580 425.030 -28.160 ;
        RECT 422.760 -29.180 422.990 -28.580 ;
        RECT 424.740 -28.690 425.030 -28.580 ;
        RECT 425.525 -28.380 425.755 -26.600 ;
        RECT 425.985 -27.430 426.500 -26.450 ;
        RECT 427.610 -27.400 428.235 -26.375 ;
        RECT 425.985 -27.990 426.870 -27.430 ;
        RECT 427.250 -28.380 427.535 -27.630 ;
        RECT 425.525 -28.615 427.535 -28.380 ;
        RECT 424.740 -29.070 425.130 -28.690 ;
        RECT 424.740 -29.180 425.030 -29.070 ;
        RECT 425.525 -29.190 425.910 -28.615 ;
        RECT 427.765 -29.180 428.235 -27.400 ;
        RECT 430.565 -28.320 430.795 -26.365 ;
        RECT 431.025 -27.540 431.400 -26.835 ;
        RECT 432.660 -27.405 433.250 -26.365 ;
        RECT 433.925 -26.855 434.155 -26.605 ;
        RECT 433.925 -27.090 436.855 -26.855 ;
        RECT 431.025 -27.950 431.910 -27.540 ;
        RECT 432.250 -28.320 432.590 -27.680 ;
        RECT 430.565 -28.555 432.590 -28.320 ;
        RECT 430.565 -29.180 430.895 -28.555 ;
        RECT 432.885 -29.120 433.250 -27.405 ;
        RECT 434.340 -28.610 434.700 -27.340 ;
        RECT 434.945 -29.125 435.175 -27.090 ;
        RECT 435.460 -29.170 435.820 -27.340 ;
        RECT 436.625 -27.785 436.855 -27.090 ;
        RECT 437.130 -29.180 437.550 -26.355 ;
        RECT 439.525 -26.815 439.755 -26.475 ;
        RECT 441.765 -26.815 441.995 -26.475 ;
        RECT 439.525 -27.050 442.475 -26.815 ;
        RECT 442.140 -27.485 442.475 -27.050 ;
        RECT 438.810 -27.950 441.670 -27.515 ;
        RECT 442.140 -27.825 446.430 -27.485 ;
        RECT 442.140 -28.330 442.475 -27.825 ;
        RECT 448.500 -27.830 451.700 -27.485 ;
        RECT 439.425 -28.560 442.475 -28.330 ;
        RECT 456.885 -28.390 457.115 -26.605 ;
        RECT 457.345 -27.540 457.720 -26.350 ;
        RECT 459.305 -27.080 459.535 -26.600 ;
        RECT 459.305 -27.310 460.450 -27.080 ;
        RECT 457.345 -27.950 458.290 -27.540 ;
        RECT 458.530 -27.840 459.850 -27.540 ;
        RECT 458.530 -28.390 458.855 -27.840 ;
        RECT 460.110 -28.160 460.450 -27.310 ;
        RECT 439.425 -29.180 439.655 -28.560 ;
        RECT 441.665 -29.180 441.895 -28.560 ;
        RECT 456.885 -28.620 458.855 -28.390 ;
        RECT 459.305 -28.510 460.450 -28.160 ;
        RECT 456.885 -29.190 457.115 -28.620 ;
        RECT 459.305 -29.190 459.535 -28.510 ;
        RECT 184.290 -30.810 189.320 -30.510 ;
        RECT 184.290 -33.790 184.520 -30.810 ;
        RECT 185.890 -33.790 186.120 -30.810 ;
        RECT 187.490 -33.790 187.720 -30.810 ;
        RECT 189.090 -33.790 189.320 -30.810 ;
        RECT 298.905 -30.930 299.135 -30.260 ;
        RECT 301.145 -30.930 301.375 -30.260 ;
        RECT 303.385 -30.930 303.615 -30.260 ;
        RECT 305.525 -30.930 305.755 -30.260 ;
        RECT 307.865 -30.880 308.095 -30.260 ;
        RECT 310.105 -30.880 310.335 -30.260 ;
        RECT 313.370 -30.445 313.750 -30.430 ;
        RECT 313.370 -30.675 314.235 -30.445 ;
        RECT 313.370 -30.690 313.750 -30.675 ;
        RECT 298.905 -31.310 305.755 -30.930 ;
        RECT 307.285 -31.110 310.335 -30.880 ;
        RECT 298.060 -31.955 301.260 -31.610 ;
        RECT 301.960 -32.110 302.760 -31.310 ;
        RECT 307.285 -31.615 307.620 -31.110 ;
        RECT 303.330 -31.955 307.620 -31.615 ;
        RECT 308.090 -31.925 310.950 -31.490 ;
        RECT 301.610 -32.220 302.760 -32.110 ;
        RECT 298.805 -32.600 305.755 -32.220 ;
        RECT 298.805 -32.965 299.035 -32.600 ;
        RECT 301.045 -32.965 301.275 -32.600 ;
        RECT 303.285 -32.965 303.515 -32.600 ;
        RECT 305.495 -32.965 305.755 -32.600 ;
        RECT 307.285 -32.390 307.620 -31.955 ;
        RECT 307.285 -32.625 310.235 -32.390 ;
        RECT 307.765 -32.965 307.995 -32.625 ;
        RECT 310.005 -32.965 310.235 -32.625 ;
        RECT 312.860 -32.830 313.195 -30.930 ;
        RECT 314.005 -31.565 314.235 -30.675 ;
        RECT 317.335 -30.960 317.615 -30.260 ;
        RECT 317.335 -31.280 318.760 -30.960 ;
        RECT 315.050 -31.565 315.430 -31.550 ;
        RECT 314.005 -31.795 315.430 -31.565 ;
        RECT 315.050 -31.810 315.430 -31.795 ;
        RECT 317.145 -31.850 318.175 -31.510 ;
        RECT 317.870 -33.040 318.175 -31.850 ;
        RECT 318.405 -33.040 318.760 -31.280 ;
        RECT 318.990 -32.460 319.295 -30.320 ;
        RECT 320.695 -30.960 320.975 -30.260 ;
        RECT 320.695 -30.990 322.120 -30.960 ;
        RECT 320.650 -31.250 322.120 -30.990 ;
        RECT 320.695 -31.280 322.120 -31.250 ;
        RECT 320.505 -31.850 321.535 -31.510 ;
        RECT 321.230 -33.040 321.535 -31.850 ;
        RECT 321.765 -33.040 322.120 -31.280 ;
        RECT 322.350 -32.460 322.655 -30.320 ;
        RECT 323.605 -32.085 323.835 -30.250 ;
        RECT 324.090 -31.680 325.355 -31.450 ;
        RECT 323.605 -32.315 324.880 -32.085 ;
        RECT 325.125 -33.110 325.355 -31.680 ;
        RECT 325.845 -32.085 326.075 -30.250 ;
        RECT 328.185 -31.005 328.415 -30.415 ;
        RECT 328.185 -31.235 329.875 -31.005 ;
        RECT 326.330 -31.680 327.595 -31.450 ;
        RECT 325.845 -32.315 327.120 -32.085 ;
        RECT 327.365 -33.110 327.595 -31.680 ;
        RECT 327.990 -31.870 329.410 -31.490 ;
        RECT 329.645 -32.130 329.875 -31.235 ;
        RECT 328.085 -32.360 329.875 -32.130 ;
        RECT 330.105 -31.025 330.455 -30.425 ;
        RECT 331.505 -30.650 332.755 -30.420 ;
        RECT 340.050 -30.480 342.265 -30.250 ;
        RECT 331.505 -31.025 331.735 -30.650 ;
        RECT 330.105 -31.255 331.735 -31.025 ;
        RECT 331.965 -31.220 332.295 -30.880 ;
        RECT 328.085 -32.830 328.315 -32.360 ;
        RECT 330.105 -32.545 330.335 -31.255 ;
        RECT 330.730 -31.870 331.760 -31.490 ;
        RECT 330.105 -32.775 330.610 -32.545 ;
        RECT 332.065 -32.565 332.295 -31.220 ;
        RECT 332.525 -31.730 332.755 -30.650 ;
        RECT 334.005 -30.880 334.235 -30.685 ;
        RECT 336.605 -30.880 336.835 -30.510 ;
        RECT 332.985 -31.340 333.215 -30.880 ;
        RECT 334.005 -31.110 336.835 -30.880 ;
        RECT 338.280 -30.795 338.920 -30.565 ;
        RECT 337.695 -31.340 337.995 -31.115 ;
        RECT 332.985 -31.570 337.995 -31.340 ;
        RECT 332.065 -32.795 332.470 -32.565 ;
        RECT 333.305 -32.850 333.535 -31.570 ;
        RECT 338.280 -31.800 338.510 -30.795 ;
        RECT 340.050 -31.590 340.280 -30.480 ;
        RECT 342.035 -30.590 342.265 -30.480 ;
        RECT 343.075 -30.480 344.260 -30.250 ;
        RECT 343.075 -30.590 343.305 -30.480 ;
        RECT 334.530 -32.030 338.510 -31.800 ;
        RECT 339.390 -31.820 340.280 -31.590 ;
        RECT 333.885 -32.260 334.115 -32.050 ;
        RECT 333.885 -32.490 337.070 -32.260 ;
        RECT 336.840 -32.880 337.070 -32.490 ;
        RECT 337.830 -32.640 338.170 -32.030 ;
        RECT 338.765 -32.880 338.995 -32.050 ;
        RECT 339.390 -32.640 339.730 -31.820 ;
        RECT 340.730 -32.050 340.960 -31.115 ;
        RECT 339.960 -32.280 340.960 -32.050 ;
        RECT 339.960 -32.880 340.190 -32.280 ;
        RECT 341.255 -32.510 341.595 -30.710 ;
        RECT 342.035 -30.820 343.305 -30.590 ;
        RECT 343.570 -31.235 343.800 -30.710 ;
        RECT 341.835 -31.465 343.800 -31.235 ;
        RECT 340.790 -32.850 341.595 -32.510 ;
        RECT 342.500 -32.620 343.045 -31.810 ;
        RECT 343.570 -31.960 343.800 -31.465 ;
        RECT 344.030 -31.730 344.260 -30.480 ;
        RECT 343.570 -32.190 346.070 -31.960 ;
        RECT 342.500 -32.670 344.135 -32.620 ;
        RECT 336.840 -33.110 340.190 -32.880 ;
        RECT 342.490 -32.930 344.135 -32.670 ;
        RECT 344.490 -32.850 344.720 -32.190 ;
        RECT 342.500 -32.980 344.135 -32.930 ;
        RECT 346.315 -33.090 346.750 -30.260 ;
        RECT 347.125 -32.085 347.355 -30.250 ;
        RECT 347.610 -31.680 348.875 -31.450 ;
        RECT 347.125 -32.315 348.400 -32.085 ;
        RECT 348.645 -33.110 348.875 -31.680 ;
        RECT 349.365 -32.085 349.595 -30.250 ;
        RECT 349.850 -31.680 351.115 -31.450 ;
        RECT 349.365 -32.315 350.640 -32.085 ;
        RECT 350.885 -33.110 351.115 -31.680 ;
        RECT 351.605 -32.085 351.835 -30.250 ;
        RECT 352.090 -31.680 353.355 -31.450 ;
        RECT 351.605 -32.315 352.880 -32.085 ;
        RECT 353.125 -33.110 353.355 -31.680 ;
        RECT 356.085 -32.085 356.315 -30.250 ;
        RECT 356.570 -31.680 357.835 -31.450 ;
        RECT 356.085 -32.315 357.360 -32.085 ;
        RECT 357.605 -33.110 357.835 -31.680 ;
        RECT 358.325 -32.085 358.555 -30.250 ;
        RECT 358.810 -31.680 360.075 -31.450 ;
        RECT 358.325 -32.315 359.600 -32.085 ;
        RECT 359.845 -33.110 360.075 -31.680 ;
        RECT 360.565 -32.085 360.795 -30.250 ;
        RECT 361.050 -31.680 362.315 -31.450 ;
        RECT 360.565 -32.315 361.840 -32.085 ;
        RECT 362.085 -33.110 362.315 -31.680 ;
        RECT 362.805 -32.085 363.035 -30.250 ;
        RECT 363.290 -31.680 364.555 -31.450 ;
        RECT 362.805 -32.315 364.080 -32.085 ;
        RECT 364.325 -33.110 364.555 -31.680 ;
        RECT 365.045 -32.085 365.275 -30.250 ;
        RECT 365.530 -31.680 366.795 -31.450 ;
        RECT 365.045 -32.315 366.320 -32.085 ;
        RECT 366.565 -33.110 366.795 -31.680 ;
        RECT 369.410 -33.100 369.810 -30.260 ;
        RECT 370.105 -32.325 370.335 -31.860 ;
        RECT 371.040 -32.095 371.390 -30.355 ;
        RECT 371.620 -30.675 373.420 -30.445 ;
        RECT 371.620 -32.325 371.850 -30.675 ;
        RECT 375.825 -30.915 376.210 -30.250 ;
        RECT 372.480 -31.150 376.210 -30.915 ;
        RECT 372.480 -31.680 372.820 -31.150 ;
        RECT 373.070 -31.830 375.530 -31.445 ;
        RECT 373.070 -31.990 373.380 -31.830 ;
        RECT 370.105 -32.555 371.850 -32.325 ;
        RECT 372.080 -32.390 373.380 -31.990 ;
        RECT 373.735 -32.390 375.385 -32.060 ;
        RECT 371.620 -32.860 371.850 -32.555 ;
        RECT 371.620 -33.090 372.980 -32.860 ;
        RECT 375.870 -33.100 376.210 -31.150 ;
        RECT 376.805 -32.085 377.035 -30.250 ;
        RECT 377.290 -31.680 378.555 -31.450 ;
        RECT 376.805 -32.315 378.080 -32.085 ;
        RECT 378.325 -33.110 378.555 -31.680 ;
        RECT 379.045 -32.085 379.275 -30.250 ;
        RECT 379.530 -31.680 380.795 -31.450 ;
        RECT 379.045 -32.315 380.320 -32.085 ;
        RECT 380.565 -33.110 380.795 -31.680 ;
        RECT 381.285 -32.085 381.515 -30.250 ;
        RECT 381.770 -31.680 383.035 -31.450 ;
        RECT 381.285 -32.315 382.560 -32.085 ;
        RECT 382.805 -33.110 383.035 -31.680 ;
        RECT 385.090 -33.100 385.490 -30.260 ;
        RECT 385.785 -32.325 386.015 -31.860 ;
        RECT 386.720 -32.095 387.070 -30.355 ;
        RECT 387.300 -30.675 389.100 -30.445 ;
        RECT 387.300 -32.325 387.530 -30.675 ;
        RECT 391.505 -30.915 391.890 -30.250 ;
        RECT 388.160 -31.150 391.890 -30.915 ;
        RECT 388.160 -31.680 388.500 -31.150 ;
        RECT 388.750 -31.830 391.210 -31.445 ;
        RECT 388.750 -31.990 389.060 -31.830 ;
        RECT 385.785 -32.555 387.530 -32.325 ;
        RECT 387.760 -32.390 389.060 -31.990 ;
        RECT 389.415 -32.390 391.065 -32.060 ;
        RECT 387.300 -32.860 387.530 -32.555 ;
        RECT 387.300 -33.090 388.660 -32.860 ;
        RECT 391.550 -33.100 391.890 -31.150 ;
        RECT 395.285 -32.085 395.515 -30.250 ;
        RECT 395.770 -31.680 397.035 -31.450 ;
        RECT 395.285 -32.315 396.560 -32.085 ;
        RECT 396.805 -33.110 397.035 -31.680 ;
        RECT 397.525 -32.085 397.755 -30.250 ;
        RECT 398.010 -31.680 399.275 -31.450 ;
        RECT 397.525 -32.315 398.800 -32.085 ;
        RECT 399.045 -33.110 399.275 -31.680 ;
        RECT 399.765 -32.085 399.995 -30.250 ;
        RECT 401.950 -30.480 404.330 -30.250 ;
        RECT 401.950 -31.145 402.290 -30.480 ;
        RECT 400.250 -31.680 401.515 -31.450 ;
        RECT 399.765 -32.315 401.040 -32.085 ;
        RECT 401.285 -33.110 401.515 -31.680 ;
        RECT 401.875 -31.870 402.770 -31.490 ;
        RECT 402.420 -32.480 402.770 -31.870 ;
        RECT 403.000 -32.770 403.305 -30.915 ;
        RECT 403.990 -31.145 404.330 -30.480 ;
        RECT 403.535 -31.870 404.440 -31.490 ;
        RECT 404.670 -31.870 405.575 -31.490 ;
        RECT 404.100 -32.480 404.440 -31.870 ;
        RECT 405.235 -32.480 405.575 -31.870 ;
        RECT 406.485 -32.085 406.715 -30.250 ;
        RECT 406.970 -31.680 408.235 -31.450 ;
        RECT 406.485 -32.315 407.760 -32.085 ;
        RECT 403.000 -33.090 404.340 -32.770 ;
        RECT 408.005 -33.110 408.235 -31.680 ;
        RECT 408.725 -32.085 408.955 -30.250 ;
        RECT 409.210 -31.680 410.475 -31.450 ;
        RECT 408.725 -32.315 410.000 -32.085 ;
        RECT 410.245 -33.110 410.475 -31.680 ;
        RECT 410.965 -32.085 411.195 -30.250 ;
        RECT 411.450 -31.680 412.715 -31.450 ;
        RECT 410.965 -32.315 412.240 -32.085 ;
        RECT 412.485 -33.110 412.715 -31.680 ;
        RECT 413.205 -32.085 413.435 -30.250 ;
        RECT 413.690 -31.680 414.955 -31.450 ;
        RECT 413.205 -32.315 414.480 -32.085 ;
        RECT 414.725 -33.110 414.955 -31.680 ;
        RECT 415.445 -32.085 415.675 -30.250 ;
        RECT 415.930 -31.680 417.195 -31.450 ;
        RECT 415.445 -32.315 416.720 -32.085 ;
        RECT 416.965 -33.110 417.195 -31.680 ;
        RECT 417.685 -32.085 417.915 -30.250 ;
        RECT 420.990 -30.480 423.370 -30.250 ;
        RECT 420.990 -31.145 421.330 -30.480 ;
        RECT 418.170 -31.680 419.435 -31.450 ;
        RECT 417.685 -32.315 418.960 -32.085 ;
        RECT 419.205 -33.110 419.435 -31.680 ;
        RECT 420.915 -31.870 421.810 -31.490 ;
        RECT 421.460 -32.480 421.810 -31.870 ;
        RECT 422.040 -32.770 422.345 -30.915 ;
        RECT 423.030 -31.145 423.370 -30.480 ;
        RECT 426.685 -30.480 429.005 -30.250 ;
        RECT 426.685 -31.280 426.915 -30.480 ;
        RECT 427.145 -31.050 428.530 -30.710 ;
        RECT 422.575 -31.870 423.480 -31.490 ;
        RECT 423.710 -31.870 424.615 -31.490 ;
        RECT 423.140 -32.480 423.480 -31.870 ;
        RECT 424.275 -32.480 424.615 -31.870 ;
        RECT 425.410 -31.740 426.385 -31.490 ;
        RECT 426.685 -31.510 427.275 -31.280 ;
        RECT 425.410 -32.040 426.815 -31.740 ;
        RECT 422.040 -33.090 423.380 -32.770 ;
        RECT 426.480 -33.090 426.815 -32.040 ;
        RECT 427.045 -33.090 427.275 -31.510 ;
        RECT 427.600 -33.090 427.935 -31.320 ;
        RECT 428.165 -33.090 428.530 -31.050 ;
        RECT 428.775 -30.950 429.005 -30.480 ;
        RECT 428.775 -31.180 429.515 -30.950 ;
        RECT 430.455 -30.960 430.735 -30.260 ;
        RECT 430.455 -30.990 431.880 -30.960 ;
        RECT 428.760 -33.090 429.055 -31.410 ;
        RECT 429.285 -33.090 429.515 -31.180 ;
        RECT 430.410 -31.250 431.880 -30.990 ;
        RECT 430.455 -31.280 431.880 -31.250 ;
        RECT 430.265 -31.850 431.295 -31.510 ;
        RECT 430.990 -33.040 431.295 -31.850 ;
        RECT 431.525 -33.040 431.880 -31.280 ;
        RECT 432.110 -32.460 432.415 -30.320 ;
        RECT 436.065 -31.990 436.360 -30.330 ;
        RECT 437.160 -31.990 437.480 -30.330 ;
        RECT 437.810 -30.590 440.810 -30.360 ;
        RECT 437.810 -32.240 438.040 -30.590 ;
        RECT 440.580 -30.770 440.810 -30.590 ;
        RECT 438.280 -31.490 438.600 -30.890 ;
        RECT 438.830 -31.260 440.315 -30.940 ;
        RECT 440.580 -31.000 441.435 -30.770 ;
        RECT 438.280 -31.910 439.190 -31.490 ;
        RECT 436.725 -32.475 439.195 -32.240 ;
        RECT 436.725 -33.030 436.955 -32.475 ;
        RECT 438.965 -33.030 439.195 -32.475 ;
        RECT 439.425 -33.030 439.730 -31.490 ;
        RECT 439.960 -33.030 440.315 -31.260 ;
        RECT 440.545 -33.030 440.850 -31.450 ;
        RECT 441.205 -33.030 441.435 -31.000 ;
        RECT 442.425 -31.005 442.655 -30.415 ;
        RECT 442.425 -31.235 444.115 -31.005 ;
        RECT 442.230 -31.870 443.650 -31.490 ;
        RECT 443.885 -32.130 444.115 -31.235 ;
        RECT 442.325 -32.360 444.115 -32.130 ;
        RECT 444.345 -31.025 444.695 -30.425 ;
        RECT 445.745 -30.650 446.995 -30.420 ;
        RECT 454.290 -30.480 456.505 -30.250 ;
        RECT 445.745 -31.025 445.975 -30.650 ;
        RECT 444.345 -31.255 445.975 -31.025 ;
        RECT 446.205 -31.220 446.535 -30.880 ;
        RECT 442.325 -32.830 442.555 -32.360 ;
        RECT 444.345 -32.545 444.575 -31.255 ;
        RECT 444.970 -31.870 446.000 -31.490 ;
        RECT 444.345 -32.775 444.850 -32.545 ;
        RECT 446.305 -32.565 446.535 -31.220 ;
        RECT 446.765 -31.730 446.995 -30.650 ;
        RECT 448.245 -30.880 448.475 -30.685 ;
        RECT 450.845 -30.880 451.075 -30.510 ;
        RECT 447.225 -31.340 447.455 -30.880 ;
        RECT 448.245 -31.110 451.075 -30.880 ;
        RECT 452.520 -30.795 453.160 -30.565 ;
        RECT 451.935 -31.340 452.235 -31.115 ;
        RECT 447.225 -31.570 452.235 -31.340 ;
        RECT 446.305 -32.795 446.710 -32.565 ;
        RECT 447.545 -32.850 447.775 -31.570 ;
        RECT 452.520 -31.800 452.750 -30.795 ;
        RECT 454.290 -31.590 454.520 -30.480 ;
        RECT 456.275 -30.590 456.505 -30.480 ;
        RECT 457.315 -30.480 458.500 -30.250 ;
        RECT 457.315 -30.590 457.545 -30.480 ;
        RECT 448.770 -32.030 452.750 -31.800 ;
        RECT 453.630 -31.820 454.520 -31.590 ;
        RECT 448.125 -32.260 448.355 -32.050 ;
        RECT 448.125 -32.490 451.310 -32.260 ;
        RECT 451.080 -32.880 451.310 -32.490 ;
        RECT 452.070 -32.640 452.410 -32.030 ;
        RECT 453.005 -32.880 453.235 -32.050 ;
        RECT 453.630 -32.640 453.970 -31.820 ;
        RECT 454.970 -32.050 455.200 -31.115 ;
        RECT 454.200 -32.280 455.200 -32.050 ;
        RECT 454.200 -32.880 454.430 -32.280 ;
        RECT 455.495 -32.510 455.835 -30.710 ;
        RECT 456.275 -30.820 457.545 -30.590 ;
        RECT 457.810 -31.235 458.040 -30.710 ;
        RECT 456.075 -31.465 458.040 -31.235 ;
        RECT 455.030 -32.850 455.835 -32.510 ;
        RECT 456.740 -32.620 457.285 -31.810 ;
        RECT 457.810 -31.960 458.040 -31.465 ;
        RECT 458.270 -31.730 458.500 -30.480 ;
        RECT 457.810 -32.190 460.310 -31.960 ;
        RECT 451.080 -33.110 454.430 -32.880 ;
        RECT 456.740 -32.980 458.375 -32.620 ;
        RECT 458.730 -32.850 458.960 -32.190 ;
        RECT 460.555 -33.090 460.990 -30.260 ;
        RECT 166.935 -34.250 169.675 -34.020 ;
        RECT 173.735 -34.250 174.875 -34.020 ;
        RECT 168.115 -35.150 168.495 -34.250 ;
        RECT 174.115 -35.150 174.495 -34.250 ;
        RECT 178.045 -34.355 179.075 -34.020 ;
        RECT 179.535 -34.355 180.565 -34.020 ;
        RECT 183.835 -34.250 189.775 -34.020 ;
        RECT 178.045 -35.215 178.425 -34.355 ;
        RECT 180.185 -35.215 180.565 -34.355 ;
        RECT 186.615 -35.150 186.995 -34.250 ;
        RECT 297.285 -35.195 298.560 -34.965 ;
        RECT 297.285 -37.030 297.515 -35.195 ;
        RECT 298.805 -35.600 299.035 -34.170 ;
        RECT 309.400 -34.400 312.750 -34.170 ;
        RECT 315.060 -34.350 316.695 -34.300 ;
        RECT 300.645 -34.920 300.875 -34.450 ;
        RECT 302.665 -34.735 303.170 -34.505 ;
        RECT 304.625 -34.715 305.030 -34.485 ;
        RECT 300.645 -35.150 302.435 -34.920 ;
        RECT 297.770 -35.830 299.035 -35.600 ;
        RECT 300.550 -35.790 301.970 -35.410 ;
        RECT 302.205 -36.045 302.435 -35.150 ;
        RECT 300.745 -36.275 302.435 -36.045 ;
        RECT 302.665 -36.025 302.895 -34.735 ;
        RECT 303.290 -35.790 304.320 -35.410 ;
        RECT 302.665 -36.255 304.295 -36.025 ;
        RECT 304.625 -36.060 304.855 -34.715 ;
        RECT 300.745 -36.865 300.975 -36.275 ;
        RECT 302.665 -36.855 303.015 -36.255 ;
        RECT 304.065 -36.630 304.295 -36.255 ;
        RECT 304.525 -36.400 304.855 -36.060 ;
        RECT 305.085 -36.630 305.315 -35.550 ;
        RECT 305.865 -35.710 306.095 -34.430 ;
        RECT 309.400 -34.790 309.630 -34.400 ;
        RECT 306.445 -35.020 309.630 -34.790 ;
        RECT 306.445 -35.230 306.675 -35.020 ;
        RECT 310.390 -35.250 310.730 -34.640 ;
        RECT 311.325 -35.230 311.555 -34.400 ;
        RECT 307.090 -35.480 311.070 -35.250 ;
        RECT 305.545 -35.940 310.555 -35.710 ;
        RECT 305.545 -36.400 305.775 -35.940 ;
        RECT 310.255 -36.165 310.555 -35.940 ;
        RECT 306.565 -36.400 309.395 -36.170 ;
        RECT 306.565 -36.595 306.795 -36.400 ;
        RECT 304.065 -36.860 305.315 -36.630 ;
        RECT 309.165 -36.770 309.395 -36.400 ;
        RECT 310.840 -36.485 311.070 -35.480 ;
        RECT 311.950 -35.460 312.290 -34.640 ;
        RECT 312.520 -35.000 312.750 -34.400 ;
        RECT 313.350 -34.770 314.155 -34.430 ;
        RECT 315.050 -34.610 316.695 -34.350 ;
        RECT 312.520 -35.230 313.520 -35.000 ;
        RECT 311.950 -35.690 312.840 -35.460 ;
        RECT 310.840 -36.715 311.480 -36.485 ;
        RECT 312.610 -36.800 312.840 -35.690 ;
        RECT 313.290 -36.165 313.520 -35.230 ;
        RECT 313.815 -36.570 314.155 -34.770 ;
        RECT 315.060 -34.660 316.695 -34.610 ;
        RECT 315.060 -35.470 315.605 -34.660 ;
        RECT 317.050 -35.090 317.280 -34.430 ;
        RECT 316.130 -35.320 318.630 -35.090 ;
        RECT 316.130 -35.815 316.360 -35.320 ;
        RECT 314.395 -36.045 316.360 -35.815 ;
        RECT 314.595 -36.690 315.865 -36.460 ;
        RECT 316.130 -36.570 316.360 -36.045 ;
        RECT 314.595 -36.800 314.825 -36.690 ;
        RECT 312.610 -37.030 314.825 -36.800 ;
        RECT 315.635 -36.800 315.865 -36.690 ;
        RECT 316.590 -36.800 316.820 -35.550 ;
        RECT 315.635 -37.030 316.820 -36.800 ;
        RECT 318.875 -37.020 319.310 -34.190 ;
        RECT 321.340 -34.510 322.680 -34.190 ;
        RECT 320.105 -35.410 320.445 -34.800 ;
        RECT 321.240 -35.410 321.580 -34.800 ;
        RECT 320.105 -35.790 321.010 -35.410 ;
        RECT 321.240 -35.790 322.145 -35.410 ;
        RECT 321.350 -36.800 321.690 -36.135 ;
        RECT 322.375 -36.365 322.680 -34.510 ;
        RECT 322.910 -35.410 323.260 -34.800 ;
        RECT 322.910 -35.790 323.805 -35.410 ;
        RECT 323.390 -36.800 323.730 -36.135 ;
        RECT 325.180 -36.350 325.515 -34.450 ;
        RECT 326.405 -35.195 327.680 -34.965 ;
        RECT 321.350 -37.030 323.730 -36.800 ;
        RECT 326.405 -37.030 326.635 -35.195 ;
        RECT 327.925 -35.600 328.155 -34.170 ;
        RECT 326.890 -35.830 328.155 -35.600 ;
        RECT 330.510 -35.245 331.100 -34.205 ;
        RECT 330.510 -36.960 330.875 -35.245 ;
        RECT 332.360 -35.380 332.735 -34.675 ;
        RECT 331.170 -36.160 331.510 -35.520 ;
        RECT 331.850 -35.790 332.735 -35.380 ;
        RECT 332.965 -36.160 333.195 -34.205 ;
        RECT 337.470 -35.430 337.775 -34.240 ;
        RECT 336.745 -35.770 337.775 -35.430 ;
        RECT 338.005 -36.000 338.360 -34.240 ;
        RECT 331.170 -36.395 333.195 -36.160 ;
        RECT 332.865 -37.020 333.195 -36.395 ;
        RECT 336.935 -36.320 338.360 -36.000 ;
        RECT 336.935 -37.020 337.215 -36.320 ;
        RECT 338.590 -36.960 338.895 -34.820 ;
        RECT 339.845 -35.195 341.120 -34.965 ;
        RECT 339.845 -37.030 340.075 -35.195 ;
        RECT 341.365 -35.600 341.595 -34.170 ;
        RECT 340.330 -35.830 341.595 -35.600 ;
        RECT 342.085 -35.195 343.360 -34.965 ;
        RECT 342.085 -37.030 342.315 -35.195 ;
        RECT 343.605 -35.600 343.835 -34.170 ;
        RECT 345.665 -34.920 345.895 -34.440 ;
        RECT 342.570 -35.830 343.835 -35.600 ;
        RECT 344.750 -35.150 345.895 -34.920 ;
        RECT 344.750 -36.000 345.090 -35.150 ;
        RECT 347.480 -35.380 347.855 -34.190 ;
        RECT 345.350 -35.680 346.670 -35.380 ;
        RECT 344.750 -36.350 345.895 -36.000 ;
        RECT 345.665 -37.030 345.895 -36.350 ;
        RECT 346.345 -36.230 346.670 -35.680 ;
        RECT 346.910 -35.790 347.855 -35.380 ;
        RECT 348.085 -36.230 348.315 -34.445 ;
        RECT 346.345 -36.460 348.315 -36.230 ;
        RECT 348.085 -37.030 348.315 -36.460 ;
        RECT 349.265 -36.590 349.590 -34.610 ;
        RECT 349.820 -37.010 350.155 -34.240 ;
        RECT 351.445 -36.090 351.675 -34.190 ;
        RECT 352.020 -35.860 352.335 -34.190 ;
        RECT 351.445 -36.320 352.265 -36.090 ;
        RECT 352.035 -36.780 352.265 -36.320 ;
        RECT 352.565 -36.320 352.920 -34.190 ;
        RECT 353.160 -35.860 353.455 -34.190 ;
        RECT 353.685 -34.505 353.915 -34.190 ;
        RECT 355.925 -34.505 356.155 -34.190 ;
        RECT 353.685 -34.735 356.155 -34.505 ;
        RECT 353.685 -35.830 354.600 -35.325 ;
        RECT 352.565 -36.550 353.960 -36.320 ;
        RECT 354.240 -36.485 354.600 -35.830 ;
        RECT 354.850 -36.780 355.080 -34.735 ;
        RECT 352.035 -37.010 355.080 -36.780 ;
        RECT 355.370 -36.960 355.695 -35.250 ;
        RECT 357.045 -36.090 357.275 -34.190 ;
        RECT 357.620 -35.860 357.935 -34.190 ;
        RECT 357.045 -36.320 357.865 -36.090 ;
        RECT 357.635 -36.780 357.865 -36.320 ;
        RECT 358.165 -36.320 358.520 -34.190 ;
        RECT 358.760 -35.860 359.055 -34.190 ;
        RECT 359.285 -34.505 359.515 -34.190 ;
        RECT 361.525 -34.505 361.755 -34.190 ;
        RECT 359.285 -34.735 361.755 -34.505 ;
        RECT 359.285 -35.830 360.200 -35.325 ;
        RECT 358.165 -36.550 359.560 -36.320 ;
        RECT 359.840 -36.485 360.200 -35.830 ;
        RECT 360.450 -36.780 360.680 -34.735 ;
        RECT 357.635 -37.010 360.680 -36.780 ;
        RECT 360.970 -36.960 361.295 -35.250 ;
        RECT 362.645 -37.010 362.980 -34.240 ;
        RECT 363.210 -36.590 363.535 -34.610 ;
        RECT 364.670 -35.245 365.260 -34.205 ;
        RECT 364.670 -36.960 365.035 -35.245 ;
        RECT 366.520 -35.380 366.895 -34.675 ;
        RECT 365.330 -36.160 365.670 -35.520 ;
        RECT 366.010 -35.790 366.895 -35.380 ;
        RECT 367.125 -36.160 367.355 -34.205 ;
        RECT 365.330 -36.395 367.355 -36.160 ;
        RECT 367.025 -37.020 367.355 -36.395 ;
        RECT 367.845 -36.160 368.075 -34.205 ;
        RECT 368.305 -35.380 368.680 -34.675 ;
        RECT 369.940 -35.245 370.530 -34.205 ;
        RECT 368.305 -35.790 369.190 -35.380 ;
        RECT 369.530 -36.160 369.870 -35.520 ;
        RECT 367.845 -36.395 369.870 -36.160 ;
        RECT 367.845 -37.020 368.175 -36.395 ;
        RECT 370.165 -36.960 370.530 -35.245 ;
        RECT 371.390 -35.245 371.980 -34.205 ;
        RECT 371.390 -36.960 371.755 -35.245 ;
        RECT 373.240 -35.380 373.615 -34.675 ;
        RECT 372.050 -36.160 372.390 -35.520 ;
        RECT 372.730 -35.790 373.615 -35.380 ;
        RECT 373.845 -36.160 374.075 -34.205 ;
        RECT 372.050 -36.395 374.075 -36.160 ;
        RECT 373.745 -37.020 374.075 -36.395 ;
        RECT 375.685 -35.195 376.960 -34.965 ;
        RECT 375.685 -37.030 375.915 -35.195 ;
        RECT 377.205 -35.600 377.435 -34.170 ;
        RECT 377.830 -34.450 378.090 -34.290 ;
        RECT 376.170 -35.830 377.435 -35.600 ;
        RECT 377.820 -36.350 378.155 -34.450 ;
        RECT 380.060 -36.350 380.395 -34.450 ;
        RECT 381.285 -36.230 381.515 -34.445 ;
        RECT 381.745 -35.380 382.120 -34.190 ;
        RECT 383.705 -34.920 383.935 -34.440 ;
        RECT 383.705 -35.150 384.850 -34.920 ;
        RECT 381.745 -35.790 382.690 -35.380 ;
        RECT 382.930 -35.680 384.250 -35.380 ;
        RECT 382.930 -36.230 383.255 -35.680 ;
        RECT 384.510 -36.000 384.850 -35.150 ;
        RECT 386.750 -35.430 387.055 -34.240 ;
        RECT 386.025 -35.770 387.055 -35.430 ;
        RECT 387.285 -36.000 387.640 -34.240 ;
        RECT 381.285 -36.460 383.255 -36.230 ;
        RECT 383.705 -36.350 384.850 -36.000 ;
        RECT 386.215 -36.030 387.640 -36.000 ;
        RECT 386.170 -36.290 387.640 -36.030 ;
        RECT 386.215 -36.320 387.640 -36.290 ;
        RECT 381.285 -37.030 381.515 -36.460 ;
        RECT 383.705 -37.030 383.935 -36.350 ;
        RECT 386.215 -37.020 386.495 -36.320 ;
        RECT 387.870 -36.960 388.175 -34.820 ;
        RECT 389.310 -35.245 389.900 -34.205 ;
        RECT 389.310 -36.960 389.675 -35.245 ;
        RECT 391.160 -35.380 391.535 -34.675 ;
        RECT 389.970 -36.160 390.310 -35.520 ;
        RECT 390.650 -35.790 391.535 -35.380 ;
        RECT 391.765 -36.160 391.995 -34.205 ;
        RECT 389.970 -36.395 391.995 -36.160 ;
        RECT 391.665 -37.020 391.995 -36.395 ;
        RECT 392.485 -35.195 393.760 -34.965 ;
        RECT 392.485 -37.030 392.715 -35.195 ;
        RECT 394.005 -35.600 394.235 -34.170 ;
        RECT 392.970 -35.830 394.235 -35.600 ;
        RECT 394.725 -35.195 396.000 -34.965 ;
        RECT 394.725 -37.030 394.955 -35.195 ;
        RECT 396.245 -35.600 396.475 -34.170 ;
        RECT 395.210 -35.830 396.475 -35.600 ;
        RECT 396.965 -35.195 398.240 -34.965 ;
        RECT 396.965 -37.030 397.195 -35.195 ;
        RECT 398.485 -35.600 398.715 -34.170 ;
        RECT 397.450 -35.830 398.715 -35.600 ;
        RECT 399.205 -35.195 400.480 -34.965 ;
        RECT 399.205 -37.030 399.435 -35.195 ;
        RECT 400.725 -35.600 400.955 -34.170 ;
        RECT 399.690 -35.830 400.955 -35.600 ;
        RECT 401.445 -35.195 402.720 -34.965 ;
        RECT 401.445 -37.030 401.675 -35.195 ;
        RECT 402.965 -35.600 403.195 -34.170 ;
        RECT 401.930 -35.830 403.195 -35.600 ;
        RECT 403.685 -35.195 404.960 -34.965 ;
        RECT 403.685 -37.030 403.915 -35.195 ;
        RECT 405.205 -35.600 405.435 -34.170 ;
        RECT 404.170 -35.830 405.435 -35.600 ;
        RECT 405.925 -35.195 407.200 -34.965 ;
        RECT 405.925 -37.030 406.155 -35.195 ;
        RECT 407.445 -35.600 407.675 -34.170 ;
        RECT 406.410 -35.830 407.675 -35.600 ;
        RECT 408.165 -35.195 409.440 -34.965 ;
        RECT 408.165 -37.030 408.395 -35.195 ;
        RECT 409.685 -35.600 409.915 -34.170 ;
        RECT 408.650 -35.830 409.915 -35.600 ;
        RECT 410.405 -35.195 411.680 -34.965 ;
        RECT 410.405 -37.030 410.635 -35.195 ;
        RECT 411.925 -35.600 412.155 -34.170 ;
        RECT 410.890 -35.830 412.155 -35.600 ;
        RECT 414.885 -35.195 416.160 -34.965 ;
        RECT 414.885 -37.030 415.115 -35.195 ;
        RECT 416.405 -35.600 416.635 -34.170 ;
        RECT 418.710 -34.450 418.970 -34.290 ;
        RECT 415.370 -35.830 416.635 -35.600 ;
        RECT 418.700 -36.350 419.035 -34.450 ;
        RECT 419.925 -35.195 421.200 -34.965 ;
        RECT 419.925 -37.030 420.155 -35.195 ;
        RECT 421.445 -35.600 421.675 -34.170 ;
        RECT 420.410 -35.830 421.675 -35.600 ;
        RECT 422.165 -35.195 423.440 -34.965 ;
        RECT 422.165 -37.030 422.395 -35.195 ;
        RECT 423.685 -35.600 423.915 -34.170 ;
        RECT 422.650 -35.830 423.915 -35.600 ;
        RECT 424.405 -35.195 425.680 -34.965 ;
        RECT 424.405 -37.030 424.635 -35.195 ;
        RECT 425.925 -35.600 426.155 -34.170 ;
        RECT 424.890 -35.830 426.155 -35.600 ;
        RECT 426.645 -35.195 427.920 -34.965 ;
        RECT 426.645 -37.030 426.875 -35.195 ;
        RECT 428.165 -35.600 428.395 -34.170 ;
        RECT 432.145 -34.400 435.565 -34.170 ;
        RECT 432.145 -34.505 432.375 -34.400 ;
        RECT 429.380 -34.735 432.375 -34.505 ;
        RECT 435.335 -34.505 435.565 -34.400 ;
        RECT 436.950 -34.400 443.560 -34.170 ;
        RECT 436.950 -34.505 437.180 -34.400 ;
        RECT 435.335 -34.740 437.180 -34.505 ;
        RECT 432.650 -34.970 434.860 -34.850 ;
        RECT 438.880 -34.860 442.550 -34.630 ;
        RECT 430.910 -35.200 436.740 -34.970 ;
        RECT 427.130 -35.830 428.395 -35.600 ;
        RECT 429.850 -35.790 437.730 -35.430 ;
        RECT 438.250 -35.770 441.870 -35.430 ;
        RECT 442.170 -36.020 442.550 -34.860 ;
        RECT 430.410 -36.395 442.550 -36.020 ;
        RECT 430.410 -37.000 430.750 -36.395 ;
        RECT 432.550 -37.000 432.890 -36.395 ;
        RECT 434.690 -37.000 435.030 -36.395 ;
        RECT 436.830 -37.000 437.170 -36.395 ;
        RECT 439.190 -37.000 439.530 -36.395 ;
        RECT 441.860 -37.000 442.550 -36.395 ;
        RECT 444.405 -37.010 444.740 -34.240 ;
        RECT 444.970 -36.590 445.295 -34.610 ;
        RECT 446.245 -36.220 446.475 -34.440 ;
        RECT 446.705 -35.270 447.220 -34.290 ;
        RECT 448.330 -35.240 448.955 -34.215 ;
        RECT 446.705 -35.830 447.590 -35.270 ;
        RECT 447.970 -36.220 448.255 -35.470 ;
        RECT 446.245 -36.455 448.255 -36.220 ;
        RECT 446.245 -37.030 446.630 -36.455 ;
        RECT 448.485 -37.020 448.955 -35.240 ;
        RECT 449.765 -35.240 450.390 -34.215 ;
        RECT 449.765 -37.020 450.235 -35.240 ;
        RECT 451.500 -35.270 452.015 -34.290 ;
        RECT 450.465 -36.220 450.750 -35.470 ;
        RECT 451.130 -35.830 452.015 -35.270 ;
        RECT 452.245 -36.220 452.475 -34.440 ;
        RECT 455.110 -34.450 455.370 -34.290 ;
        RECT 450.465 -36.455 452.475 -36.220 ;
        RECT 455.100 -36.350 455.435 -34.450 ;
        RECT 458.225 -34.920 458.455 -34.440 ;
        RECT 457.310 -35.150 458.455 -34.920 ;
        RECT 457.310 -36.000 457.650 -35.150 ;
        RECT 460.040 -35.380 460.415 -34.190 ;
        RECT 457.910 -35.680 459.230 -35.380 ;
        RECT 457.310 -36.350 458.455 -36.000 ;
        RECT 452.090 -37.030 452.475 -36.455 ;
        RECT 458.225 -37.030 458.455 -36.350 ;
        RECT 458.905 -36.230 459.230 -35.680 ;
        RECT 459.470 -35.790 460.415 -35.380 ;
        RECT 460.645 -36.230 460.875 -34.445 ;
        RECT 458.905 -36.460 460.875 -36.230 ;
        RECT 460.645 -37.030 460.875 -36.460 ;
        RECT 298.905 -38.770 299.135 -38.100 ;
        RECT 301.145 -38.770 301.375 -38.100 ;
        RECT 303.385 -38.770 303.615 -38.100 ;
        RECT 305.525 -38.770 305.755 -38.100 ;
        RECT 307.865 -38.720 308.095 -38.100 ;
        RECT 310.105 -38.720 310.335 -38.100 ;
        RECT 298.905 -39.150 305.755 -38.770 ;
        RECT 307.285 -38.950 310.335 -38.720 ;
        RECT 298.060 -39.795 301.260 -39.450 ;
        RECT 301.960 -40.060 302.760 -39.150 ;
        RECT 307.285 -39.455 307.620 -38.950 ;
        RECT 303.330 -39.795 307.620 -39.455 ;
        RECT 308.090 -39.765 310.950 -39.330 ;
        RECT 298.805 -40.440 305.755 -40.060 ;
        RECT 298.805 -40.805 299.035 -40.440 ;
        RECT 301.045 -40.805 301.275 -40.440 ;
        RECT 303.285 -40.805 303.515 -40.440 ;
        RECT 305.495 -40.450 305.755 -40.440 ;
        RECT 307.285 -40.230 307.620 -39.795 ;
        RECT 305.495 -40.805 305.850 -40.450 ;
        RECT 307.285 -40.465 310.235 -40.230 ;
        RECT 307.765 -40.805 307.995 -40.465 ;
        RECT 310.005 -40.805 310.235 -40.465 ;
        RECT 305.590 -40.830 305.850 -40.805 ;
        RECT 312.245 -40.880 312.580 -38.110 ;
        RECT 312.810 -40.510 313.135 -38.530 ;
        RECT 317.550 -39.190 318.180 -38.135 ;
        RECT 317.550 -40.440 317.880 -39.190 ;
        RECT 319.540 -39.740 319.900 -38.135 ;
        RECT 320.140 -38.350 321.345 -38.120 ;
        RECT 318.145 -39.970 319.000 -39.840 ;
        RECT 320.140 -39.970 320.370 -38.350 ;
        RECT 318.145 -40.200 320.370 -39.970 ;
        RECT 317.550 -40.870 318.315 -40.440 ;
        RECT 319.975 -40.950 320.370 -40.200 ;
        RECT 320.600 -40.405 321.020 -38.600 ;
        RECT 322.940 -40.670 323.275 -38.770 ;
        RECT 326.030 -39.875 326.395 -38.160 ;
        RECT 328.385 -38.725 328.715 -38.100 ;
        RECT 326.690 -38.960 328.715 -38.725 ;
        RECT 326.690 -39.600 327.030 -38.960 ;
        RECT 327.370 -39.740 328.255 -39.330 ;
        RECT 326.030 -40.915 326.620 -39.875 ;
        RECT 327.880 -40.445 328.255 -39.740 ;
        RECT 328.485 -40.915 328.715 -38.960 ;
        RECT 329.305 -38.845 329.535 -38.255 ;
        RECT 329.305 -39.075 330.995 -38.845 ;
        RECT 329.240 -39.710 330.530 -39.330 ;
        RECT 330.765 -39.970 330.995 -39.075 ;
        RECT 329.205 -40.200 330.995 -39.970 ;
        RECT 331.225 -38.865 331.575 -38.265 ;
        RECT 332.625 -38.490 333.875 -38.260 ;
        RECT 341.170 -38.320 343.385 -38.090 ;
        RECT 332.625 -38.865 332.855 -38.490 ;
        RECT 331.225 -39.095 332.855 -38.865 ;
        RECT 333.085 -39.060 333.415 -38.720 ;
        RECT 329.205 -40.670 329.435 -40.200 ;
        RECT 331.225 -40.385 331.455 -39.095 ;
        RECT 331.850 -39.710 332.880 -39.330 ;
        RECT 331.225 -40.615 331.730 -40.385 ;
        RECT 333.185 -40.405 333.415 -39.060 ;
        RECT 333.645 -39.570 333.875 -38.490 ;
        RECT 335.125 -38.720 335.355 -38.525 ;
        RECT 337.725 -38.720 337.955 -38.350 ;
        RECT 334.105 -39.180 334.335 -38.720 ;
        RECT 335.125 -38.950 337.955 -38.720 ;
        RECT 339.400 -38.635 340.040 -38.405 ;
        RECT 338.815 -39.180 339.115 -38.955 ;
        RECT 334.105 -39.410 339.115 -39.180 ;
        RECT 333.185 -40.635 333.590 -40.405 ;
        RECT 334.425 -40.690 334.655 -39.410 ;
        RECT 339.400 -39.640 339.630 -38.635 ;
        RECT 341.170 -39.430 341.400 -38.320 ;
        RECT 343.155 -38.430 343.385 -38.320 ;
        RECT 344.195 -38.320 345.380 -38.090 ;
        RECT 344.195 -38.430 344.425 -38.320 ;
        RECT 335.650 -39.870 339.630 -39.640 ;
        RECT 340.510 -39.660 341.400 -39.430 ;
        RECT 335.005 -40.100 335.235 -39.890 ;
        RECT 335.005 -40.330 338.190 -40.100 ;
        RECT 337.960 -40.720 338.190 -40.330 ;
        RECT 338.950 -40.480 339.290 -39.870 ;
        RECT 339.885 -40.720 340.115 -39.890 ;
        RECT 340.510 -40.480 340.850 -39.660 ;
        RECT 341.850 -39.890 342.080 -38.955 ;
        RECT 341.080 -40.120 342.080 -39.890 ;
        RECT 341.080 -40.720 341.310 -40.120 ;
        RECT 342.375 -40.350 342.715 -38.550 ;
        RECT 343.155 -38.660 344.425 -38.430 ;
        RECT 344.690 -39.075 344.920 -38.550 ;
        RECT 342.955 -39.305 344.920 -39.075 ;
        RECT 341.910 -40.690 342.715 -40.350 ;
        RECT 343.620 -40.460 344.165 -39.650 ;
        RECT 344.690 -39.800 344.920 -39.305 ;
        RECT 345.150 -39.570 345.380 -38.320 ;
        RECT 344.690 -40.030 347.190 -39.800 ;
        RECT 337.960 -40.950 341.310 -40.720 ;
        RECT 343.620 -40.820 345.255 -40.460 ;
        RECT 345.610 -40.690 345.840 -40.030 ;
        RECT 347.435 -40.930 347.870 -38.100 ;
        RECT 348.245 -39.925 348.475 -38.090 ;
        RECT 348.730 -39.520 349.995 -39.290 ;
        RECT 348.245 -40.155 349.520 -39.925 ;
        RECT 349.765 -40.950 349.995 -39.520 ;
        RECT 350.485 -39.925 350.715 -38.090 ;
        RECT 350.970 -39.520 352.235 -39.290 ;
        RECT 350.485 -40.155 351.760 -39.925 ;
        RECT 352.005 -40.950 352.235 -39.520 ;
        RECT 352.725 -39.925 352.955 -38.090 ;
        RECT 353.210 -39.520 354.475 -39.290 ;
        RECT 352.725 -40.155 354.000 -39.925 ;
        RECT 354.245 -40.950 354.475 -39.520 ;
        RECT 356.545 -40.510 356.870 -38.530 ;
        RECT 357.100 -40.880 357.435 -38.110 ;
        RECT 358.325 -39.925 358.555 -38.090 ;
        RECT 358.810 -39.520 360.075 -39.290 ;
        RECT 358.325 -40.155 359.600 -39.925 ;
        RECT 359.845 -40.950 360.075 -39.520 ;
        RECT 360.565 -39.925 360.795 -38.090 ;
        RECT 361.050 -39.520 362.315 -39.290 ;
        RECT 360.565 -40.155 361.840 -39.925 ;
        RECT 362.085 -40.950 362.315 -39.520 ;
        RECT 362.805 -39.925 363.035 -38.090 ;
        RECT 363.290 -39.520 364.555 -39.290 ;
        RECT 362.805 -40.155 364.080 -39.925 ;
        RECT 364.325 -40.950 364.555 -39.520 ;
        RECT 365.045 -39.925 365.275 -38.090 ;
        RECT 365.530 -39.520 366.795 -39.290 ;
        RECT 365.045 -40.155 366.320 -39.925 ;
        RECT 366.565 -40.950 366.795 -39.520 ;
        RECT 367.285 -39.925 367.515 -38.090 ;
        RECT 369.625 -38.845 369.855 -38.255 ;
        RECT 369.625 -39.075 371.315 -38.845 ;
        RECT 367.770 -39.520 369.035 -39.290 ;
        RECT 367.285 -40.155 368.560 -39.925 ;
        RECT 368.805 -40.950 369.035 -39.520 ;
        RECT 369.430 -39.710 370.850 -39.330 ;
        RECT 371.085 -39.970 371.315 -39.075 ;
        RECT 369.525 -40.200 371.315 -39.970 ;
        RECT 371.545 -38.865 371.895 -38.265 ;
        RECT 372.945 -38.490 374.195 -38.260 ;
        RECT 381.490 -38.320 383.705 -38.090 ;
        RECT 372.945 -38.865 373.175 -38.490 ;
        RECT 371.545 -39.095 373.175 -38.865 ;
        RECT 373.405 -39.060 373.735 -38.720 ;
        RECT 369.525 -40.670 369.755 -40.200 ;
        RECT 371.545 -40.385 371.775 -39.095 ;
        RECT 372.170 -39.710 373.200 -39.330 ;
        RECT 371.545 -40.615 372.050 -40.385 ;
        RECT 373.505 -40.405 373.735 -39.060 ;
        RECT 373.965 -39.570 374.195 -38.490 ;
        RECT 375.445 -38.720 375.675 -38.525 ;
        RECT 378.045 -38.720 378.275 -38.350 ;
        RECT 374.425 -39.180 374.655 -38.720 ;
        RECT 375.445 -38.950 378.275 -38.720 ;
        RECT 379.720 -38.635 380.360 -38.405 ;
        RECT 379.135 -39.180 379.435 -38.955 ;
        RECT 374.425 -39.410 379.435 -39.180 ;
        RECT 373.505 -40.635 373.910 -40.405 ;
        RECT 374.745 -40.690 374.975 -39.410 ;
        RECT 379.720 -39.640 379.950 -38.635 ;
        RECT 381.490 -39.430 381.720 -38.320 ;
        RECT 383.475 -38.430 383.705 -38.320 ;
        RECT 384.515 -38.320 385.700 -38.090 ;
        RECT 384.515 -38.430 384.745 -38.320 ;
        RECT 375.970 -39.870 379.950 -39.640 ;
        RECT 380.830 -39.660 381.720 -39.430 ;
        RECT 375.325 -40.100 375.555 -39.890 ;
        RECT 375.325 -40.330 378.510 -40.100 ;
        RECT 378.280 -40.720 378.510 -40.330 ;
        RECT 379.270 -40.480 379.610 -39.870 ;
        RECT 380.205 -40.720 380.435 -39.890 ;
        RECT 380.830 -40.480 381.170 -39.660 ;
        RECT 382.170 -39.890 382.400 -38.955 ;
        RECT 381.400 -40.120 382.400 -39.890 ;
        RECT 381.400 -40.720 381.630 -40.120 ;
        RECT 382.695 -40.350 383.035 -38.550 ;
        RECT 383.475 -38.660 384.745 -38.430 ;
        RECT 385.010 -39.075 385.240 -38.550 ;
        RECT 383.275 -39.305 385.240 -39.075 ;
        RECT 382.230 -40.690 383.035 -40.350 ;
        RECT 383.940 -40.460 384.485 -39.650 ;
        RECT 385.010 -39.800 385.240 -39.305 ;
        RECT 385.470 -39.570 385.700 -38.320 ;
        RECT 385.010 -40.030 387.510 -39.800 ;
        RECT 383.940 -40.510 385.575 -40.460 ;
        RECT 378.280 -40.950 381.630 -40.720 ;
        RECT 383.930 -40.770 385.575 -40.510 ;
        RECT 385.930 -40.690 386.160 -40.030 ;
        RECT 383.940 -40.820 385.575 -40.770 ;
        RECT 387.755 -40.930 388.190 -38.100 ;
        RECT 388.565 -39.925 388.795 -38.090 ;
        RECT 389.050 -39.520 390.315 -39.290 ;
        RECT 388.565 -40.155 389.840 -39.925 ;
        RECT 390.085 -40.950 390.315 -39.520 ;
        RECT 390.700 -40.670 391.035 -38.770 ;
        RECT 391.925 -39.925 392.155 -38.090 ;
        RECT 392.410 -39.520 393.675 -39.290 ;
        RECT 391.925 -40.155 393.200 -39.925 ;
        RECT 393.445 -40.950 393.675 -39.520 ;
        RECT 395.285 -39.925 395.515 -38.090 ;
        RECT 395.770 -39.520 397.035 -39.290 ;
        RECT 395.285 -40.155 396.560 -39.925 ;
        RECT 396.805 -40.950 397.035 -39.520 ;
        RECT 397.525 -39.925 397.755 -38.090 ;
        RECT 399.865 -38.845 400.095 -38.255 ;
        RECT 399.865 -39.075 401.555 -38.845 ;
        RECT 398.010 -39.520 399.275 -39.290 ;
        RECT 397.525 -40.155 398.800 -39.925 ;
        RECT 399.045 -40.950 399.275 -39.520 ;
        RECT 399.800 -39.710 401.090 -39.330 ;
        RECT 401.325 -39.970 401.555 -39.075 ;
        RECT 399.765 -40.200 401.555 -39.970 ;
        RECT 401.785 -38.865 402.135 -38.265 ;
        RECT 403.185 -38.490 404.435 -38.260 ;
        RECT 411.730 -38.320 413.945 -38.090 ;
        RECT 403.185 -38.865 403.415 -38.490 ;
        RECT 401.785 -39.095 403.415 -38.865 ;
        RECT 403.645 -39.060 403.975 -38.720 ;
        RECT 399.765 -40.670 399.995 -40.200 ;
        RECT 401.785 -40.385 402.015 -39.095 ;
        RECT 402.410 -39.710 403.440 -39.330 ;
        RECT 401.785 -40.615 402.290 -40.385 ;
        RECT 403.745 -40.405 403.975 -39.060 ;
        RECT 404.205 -39.570 404.435 -38.490 ;
        RECT 405.685 -38.720 405.915 -38.525 ;
        RECT 408.285 -38.720 408.515 -38.350 ;
        RECT 404.665 -39.180 404.895 -38.720 ;
        RECT 405.685 -38.950 408.515 -38.720 ;
        RECT 409.960 -38.635 410.600 -38.405 ;
        RECT 409.375 -39.180 409.675 -38.955 ;
        RECT 404.665 -39.410 409.675 -39.180 ;
        RECT 403.745 -40.635 404.150 -40.405 ;
        RECT 404.985 -40.690 405.215 -39.410 ;
        RECT 409.960 -39.640 410.190 -38.635 ;
        RECT 411.730 -39.430 411.960 -38.320 ;
        RECT 413.715 -38.430 413.945 -38.320 ;
        RECT 414.755 -38.320 415.940 -38.090 ;
        RECT 414.755 -38.430 414.985 -38.320 ;
        RECT 406.210 -39.870 410.190 -39.640 ;
        RECT 411.070 -39.660 411.960 -39.430 ;
        RECT 405.565 -40.100 405.795 -39.890 ;
        RECT 405.565 -40.330 408.750 -40.100 ;
        RECT 408.520 -40.720 408.750 -40.330 ;
        RECT 409.510 -40.480 409.850 -39.870 ;
        RECT 410.445 -40.720 410.675 -39.890 ;
        RECT 411.070 -40.480 411.410 -39.660 ;
        RECT 412.410 -39.890 412.640 -38.955 ;
        RECT 411.640 -40.120 412.640 -39.890 ;
        RECT 411.640 -40.720 411.870 -40.120 ;
        RECT 412.935 -40.350 413.275 -38.550 ;
        RECT 413.715 -38.660 414.985 -38.430 ;
        RECT 415.250 -39.075 415.480 -38.550 ;
        RECT 413.515 -39.305 415.480 -39.075 ;
        RECT 412.470 -40.690 413.275 -40.350 ;
        RECT 414.180 -40.460 414.725 -39.650 ;
        RECT 415.250 -39.800 415.480 -39.305 ;
        RECT 415.710 -39.570 415.940 -38.320 ;
        RECT 415.250 -40.030 417.750 -39.800 ;
        RECT 408.520 -40.950 411.870 -40.720 ;
        RECT 414.180 -40.820 415.815 -40.460 ;
        RECT 416.170 -40.690 416.400 -40.030 ;
        RECT 417.995 -40.930 418.430 -38.100 ;
        RECT 420.425 -38.770 420.655 -38.100 ;
        RECT 422.665 -38.770 422.895 -38.100 ;
        RECT 424.905 -38.770 425.135 -38.100 ;
        RECT 427.045 -38.770 427.275 -38.100 ;
        RECT 429.385 -38.720 429.615 -38.100 ;
        RECT 431.625 -38.720 431.855 -38.100 ;
        RECT 420.425 -39.150 427.275 -38.770 ;
        RECT 428.805 -38.950 431.855 -38.720 ;
        RECT 419.580 -39.795 422.780 -39.450 ;
        RECT 423.480 -40.060 424.280 -39.150 ;
        RECT 428.805 -39.455 429.140 -38.950 ;
        RECT 424.850 -39.795 429.140 -39.455 ;
        RECT 429.610 -39.765 432.470 -39.330 ;
        RECT 420.325 -40.440 427.275 -40.060 ;
        RECT 420.325 -40.805 420.555 -40.440 ;
        RECT 422.565 -40.805 422.795 -40.440 ;
        RECT 424.805 -40.805 425.035 -40.440 ;
        RECT 427.015 -40.450 427.275 -40.440 ;
        RECT 428.805 -40.230 429.140 -39.795 ;
        RECT 427.015 -40.805 427.370 -40.450 ;
        RECT 428.805 -40.465 431.755 -40.230 ;
        RECT 435.505 -40.300 435.810 -38.160 ;
        RECT 436.070 -38.800 436.330 -38.770 ;
        RECT 437.185 -38.800 437.465 -38.100 ;
        RECT 436.040 -39.120 437.465 -38.800 ;
        RECT 429.285 -40.805 429.515 -40.465 ;
        RECT 431.525 -40.805 431.755 -40.465 ;
        RECT 427.110 -40.830 427.370 -40.805 ;
        RECT 436.040 -40.880 436.395 -39.120 ;
        RECT 436.625 -39.690 437.655 -39.350 ;
        RECT 436.625 -40.880 436.930 -39.690 ;
        RECT 438.805 -40.880 439.140 -38.110 ;
        RECT 439.370 -40.510 439.695 -38.530 ;
        RECT 443.345 -38.720 443.575 -38.100 ;
        RECT 445.585 -38.720 445.815 -38.100 ;
        RECT 443.345 -38.950 446.395 -38.720 ;
        RECT 442.730 -39.765 445.590 -39.330 ;
        RECT 446.060 -39.455 446.395 -38.950 ;
        RECT 447.925 -38.770 448.155 -38.100 ;
        RECT 450.065 -38.770 450.295 -38.100 ;
        RECT 452.305 -38.770 452.535 -38.100 ;
        RECT 454.545 -38.770 454.775 -38.100 ;
        RECT 447.925 -39.150 454.775 -38.770 ;
        RECT 457.350 -38.780 457.610 -38.770 ;
        RECT 458.215 -38.780 458.445 -38.090 ;
        RECT 446.060 -39.795 450.350 -39.455 ;
        RECT 446.060 -40.230 446.395 -39.795 ;
        RECT 450.920 -40.060 451.720 -39.150 ;
        RECT 457.320 -39.270 458.445 -38.780 ;
        RECT 460.645 -38.855 460.875 -38.090 ;
        RECT 458.990 -39.090 460.875 -38.855 ;
        RECT 452.420 -39.795 455.620 -39.450 ;
        RECT 443.445 -40.465 446.395 -40.230 ;
        RECT 447.925 -40.440 454.875 -40.060 ;
        RECT 457.320 -40.180 457.640 -39.270 ;
        RECT 458.990 -39.590 459.220 -39.090 ;
        RECT 457.880 -39.930 459.220 -39.590 ;
        RECT 457.320 -40.415 458.445 -40.180 ;
        RECT 447.925 -40.450 448.185 -40.440 ;
        RECT 443.445 -40.805 443.675 -40.465 ;
        RECT 445.685 -40.805 445.915 -40.465 ;
        RECT 447.830 -40.805 448.185 -40.450 ;
        RECT 450.165 -40.805 450.395 -40.440 ;
        RECT 452.405 -40.805 452.635 -40.440 ;
        RECT 454.645 -40.805 454.875 -40.440 ;
        RECT 447.830 -40.830 448.090 -40.805 ;
        RECT 458.215 -40.910 458.445 -40.415 ;
        RECT 460.645 -40.910 460.875 -39.090 ;
        RECT 298.805 -42.520 299.035 -42.155 ;
        RECT 301.045 -42.520 301.275 -42.155 ;
        RECT 303.285 -42.520 303.515 -42.155 ;
        RECT 305.495 -42.520 305.755 -42.155 ;
        RECT 307.765 -42.495 307.995 -42.155 ;
        RECT 310.005 -42.495 310.235 -42.155 ;
        RECT 298.805 -42.900 305.755 -42.520 ;
        RECT 307.285 -42.730 310.235 -42.495 ;
        RECT 298.060 -43.510 301.260 -43.165 ;
        RECT 301.960 -43.810 302.760 -42.900 ;
        RECT 307.285 -43.165 307.620 -42.730 ;
        RECT 313.185 -42.760 313.415 -42.280 ;
        RECT 303.330 -43.505 307.620 -43.165 ;
        RECT 312.270 -42.990 313.415 -42.760 ;
        RECT 298.905 -44.190 305.755 -43.810 ;
        RECT 298.905 -44.370 299.135 -44.190 ;
        RECT 298.870 -44.750 299.135 -44.370 ;
        RECT 298.905 -44.860 299.135 -44.750 ;
        RECT 301.145 -44.860 301.375 -44.190 ;
        RECT 303.385 -44.860 303.615 -44.190 ;
        RECT 305.525 -44.860 305.755 -44.190 ;
        RECT 307.285 -44.010 307.620 -43.505 ;
        RECT 308.090 -43.630 310.950 -43.195 ;
        RECT 312.270 -43.840 312.610 -42.990 ;
        RECT 315.000 -43.220 315.375 -42.030 ;
        RECT 325.080 -42.240 328.430 -42.010 ;
        RECT 312.870 -43.520 314.190 -43.220 ;
        RECT 307.285 -44.240 310.335 -44.010 ;
        RECT 312.270 -44.190 313.415 -43.840 ;
        RECT 307.865 -44.860 308.095 -44.240 ;
        RECT 310.105 -44.860 310.335 -44.240 ;
        RECT 313.185 -44.870 313.415 -44.190 ;
        RECT 313.865 -44.070 314.190 -43.520 ;
        RECT 314.430 -43.630 315.375 -43.220 ;
        RECT 315.605 -44.070 315.835 -42.285 ;
        RECT 316.325 -42.760 316.555 -42.290 ;
        RECT 318.345 -42.575 318.850 -42.345 ;
        RECT 320.305 -42.555 320.710 -42.325 ;
        RECT 316.325 -42.990 318.115 -42.760 ;
        RECT 316.360 -43.630 317.650 -43.250 ;
        RECT 317.885 -43.885 318.115 -42.990 ;
        RECT 313.865 -44.300 315.835 -44.070 ;
        RECT 315.605 -44.870 315.835 -44.300 ;
        RECT 316.425 -44.115 318.115 -43.885 ;
        RECT 318.345 -43.865 318.575 -42.575 ;
        RECT 318.970 -43.630 320.000 -43.250 ;
        RECT 318.345 -44.095 319.975 -43.865 ;
        RECT 320.305 -43.900 320.535 -42.555 ;
        RECT 316.425 -44.705 316.655 -44.115 ;
        RECT 318.345 -44.695 318.695 -44.095 ;
        RECT 319.745 -44.470 319.975 -44.095 ;
        RECT 320.205 -44.240 320.535 -43.900 ;
        RECT 320.765 -44.470 320.995 -43.390 ;
        RECT 321.545 -43.550 321.775 -42.270 ;
        RECT 325.080 -42.630 325.310 -42.240 ;
        RECT 322.125 -42.860 325.310 -42.630 ;
        RECT 322.125 -43.070 322.355 -42.860 ;
        RECT 326.070 -43.090 326.410 -42.480 ;
        RECT 327.005 -43.070 327.235 -42.240 ;
        RECT 322.770 -43.320 326.750 -43.090 ;
        RECT 321.225 -43.780 326.235 -43.550 ;
        RECT 321.225 -44.240 321.455 -43.780 ;
        RECT 325.935 -44.005 326.235 -43.780 ;
        RECT 322.245 -44.240 325.075 -44.010 ;
        RECT 322.245 -44.435 322.475 -44.240 ;
        RECT 319.745 -44.700 320.995 -44.470 ;
        RECT 324.845 -44.610 325.075 -44.240 ;
        RECT 326.520 -44.325 326.750 -43.320 ;
        RECT 327.630 -43.300 327.970 -42.480 ;
        RECT 328.200 -42.840 328.430 -42.240 ;
        RECT 329.030 -42.610 329.835 -42.270 ;
        RECT 328.200 -43.070 329.200 -42.840 ;
        RECT 327.630 -43.530 328.520 -43.300 ;
        RECT 326.520 -44.555 327.160 -44.325 ;
        RECT 328.290 -44.640 328.520 -43.530 ;
        RECT 328.970 -44.005 329.200 -43.070 ;
        RECT 329.495 -44.410 329.835 -42.610 ;
        RECT 330.740 -42.500 332.375 -42.140 ;
        RECT 330.740 -43.310 331.285 -42.500 ;
        RECT 332.730 -42.930 332.960 -42.270 ;
        RECT 331.810 -43.160 334.310 -42.930 ;
        RECT 331.810 -43.655 332.040 -43.160 ;
        RECT 330.075 -43.885 332.040 -43.655 ;
        RECT 330.275 -44.530 331.545 -44.300 ;
        RECT 331.810 -44.410 332.040 -43.885 ;
        RECT 330.275 -44.640 330.505 -44.530 ;
        RECT 328.290 -44.870 330.505 -44.640 ;
        RECT 331.315 -44.640 331.545 -44.530 ;
        RECT 332.270 -44.640 332.500 -43.390 ;
        RECT 331.315 -44.870 332.500 -44.640 ;
        RECT 334.555 -44.860 334.990 -42.030 ;
        RECT 338.945 -42.760 339.175 -42.280 ;
        RECT 338.030 -42.990 339.175 -42.760 ;
        RECT 338.030 -43.840 338.370 -42.990 ;
        RECT 340.760 -43.220 341.135 -42.030 ;
        RECT 338.630 -43.520 339.950 -43.220 ;
        RECT 338.030 -44.190 339.175 -43.840 ;
        RECT 338.945 -44.870 339.175 -44.190 ;
        RECT 339.625 -44.070 339.950 -43.520 ;
        RECT 340.190 -43.630 341.135 -43.220 ;
        RECT 341.365 -44.070 341.595 -42.285 ;
        RECT 343.080 -42.350 344.420 -42.030 ;
        RECT 342.500 -43.250 342.850 -42.640 ;
        RECT 341.955 -43.630 342.850 -43.250 ;
        RECT 339.625 -44.300 341.595 -44.070 ;
        RECT 341.365 -44.870 341.595 -44.300 ;
        RECT 342.030 -44.640 342.370 -43.975 ;
        RECT 343.080 -44.205 343.385 -42.350 ;
        RECT 346.670 -42.520 347.435 -42.090 ;
        RECT 344.180 -43.250 344.520 -42.640 ;
        RECT 345.315 -43.250 345.655 -42.640 ;
        RECT 343.615 -43.630 344.520 -43.250 ;
        RECT 344.750 -43.630 345.655 -43.250 ;
        RECT 346.670 -43.770 347.000 -42.520 ;
        RECT 349.095 -42.760 349.490 -42.010 ;
        RECT 347.265 -42.990 349.490 -42.760 ;
        RECT 347.265 -43.120 348.120 -42.990 ;
        RECT 344.070 -44.640 344.410 -43.975 ;
        RECT 342.030 -44.870 344.410 -44.640 ;
        RECT 346.670 -44.825 347.300 -43.770 ;
        RECT 348.660 -44.825 349.020 -43.220 ;
        RECT 349.260 -44.610 349.490 -42.990 ;
        RECT 349.720 -44.360 350.140 -42.555 ;
        RECT 351.045 -43.035 352.320 -42.805 ;
        RECT 349.260 -44.840 350.465 -44.610 ;
        RECT 351.045 -44.870 351.275 -43.035 ;
        RECT 352.565 -43.440 352.795 -42.010 ;
        RECT 351.530 -43.670 352.795 -43.440 ;
        RECT 354.850 -44.860 355.285 -42.030 ;
        RECT 356.880 -42.930 357.110 -42.270 ;
        RECT 357.465 -42.500 359.100 -42.140 ;
        RECT 361.410 -42.240 364.760 -42.010 ;
        RECT 355.530 -43.160 358.030 -42.930 ;
        RECT 357.340 -44.640 357.570 -43.390 ;
        RECT 357.800 -43.655 358.030 -43.160 ;
        RECT 358.555 -43.310 359.100 -42.500 ;
        RECT 360.005 -42.610 360.810 -42.270 ;
        RECT 357.800 -43.885 359.765 -43.655 ;
        RECT 357.800 -44.410 358.030 -43.885 ;
        RECT 358.295 -44.530 359.565 -44.300 ;
        RECT 360.005 -44.410 360.345 -42.610 ;
        RECT 361.410 -42.840 361.640 -42.240 ;
        RECT 360.640 -43.070 361.640 -42.840 ;
        RECT 360.640 -44.005 360.870 -43.070 ;
        RECT 361.870 -43.300 362.210 -42.480 ;
        RECT 362.605 -43.070 362.835 -42.240 ;
        RECT 363.430 -43.090 363.770 -42.480 ;
        RECT 364.530 -42.630 364.760 -42.240 ;
        RECT 364.530 -42.860 367.715 -42.630 ;
        RECT 367.485 -43.070 367.715 -42.860 ;
        RECT 361.320 -43.530 362.210 -43.300 ;
        RECT 363.090 -43.320 367.070 -43.090 ;
        RECT 358.295 -44.640 358.525 -44.530 ;
        RECT 357.340 -44.870 358.525 -44.640 ;
        RECT 359.335 -44.640 359.565 -44.530 ;
        RECT 361.320 -44.640 361.550 -43.530 ;
        RECT 363.090 -44.325 363.320 -43.320 ;
        RECT 368.065 -43.550 368.295 -42.270 ;
        RECT 369.130 -42.555 369.535 -42.325 ;
        RECT 363.605 -43.780 368.615 -43.550 ;
        RECT 363.605 -44.005 363.905 -43.780 ;
        RECT 362.680 -44.555 363.320 -44.325 ;
        RECT 364.765 -44.240 367.595 -44.010 ;
        RECT 368.385 -44.240 368.615 -43.780 ;
        RECT 364.765 -44.610 364.995 -44.240 ;
        RECT 367.365 -44.435 367.595 -44.240 ;
        RECT 368.845 -44.470 369.075 -43.390 ;
        RECT 369.305 -43.900 369.535 -42.555 ;
        RECT 370.990 -42.575 371.495 -42.345 ;
        RECT 369.840 -43.630 370.870 -43.250 ;
        RECT 371.265 -43.865 371.495 -42.575 ;
        RECT 373.285 -42.760 373.515 -42.290 ;
        RECT 369.305 -44.240 369.635 -43.900 ;
        RECT 369.865 -44.095 371.495 -43.865 ;
        RECT 369.865 -44.470 370.095 -44.095 ;
        RECT 359.335 -44.870 361.550 -44.640 ;
        RECT 368.845 -44.700 370.095 -44.470 ;
        RECT 371.145 -44.695 371.495 -44.095 ;
        RECT 371.725 -42.990 373.515 -42.760 ;
        RECT 371.725 -43.885 371.955 -42.990 ;
        RECT 372.190 -43.630 373.480 -43.250 ;
        RECT 371.725 -44.115 373.415 -43.885 ;
        RECT 373.185 -44.705 373.415 -44.115 ;
        RECT 376.085 -44.850 376.420 -42.080 ;
        RECT 376.650 -44.430 376.975 -42.450 ;
        RECT 379.045 -44.000 379.275 -42.045 ;
        RECT 379.505 -43.220 379.880 -42.515 ;
        RECT 381.140 -43.085 381.730 -42.045 ;
        RECT 379.505 -43.630 380.390 -43.220 ;
        RECT 380.730 -44.000 381.070 -43.360 ;
        RECT 379.045 -44.235 381.070 -44.000 ;
        RECT 379.045 -44.860 379.375 -44.235 ;
        RECT 381.365 -44.800 381.730 -43.085 ;
        RECT 382.290 -44.860 382.725 -42.030 ;
        RECT 384.905 -42.190 386.540 -42.140 ;
        RECT 384.320 -42.930 384.550 -42.270 ;
        RECT 384.905 -42.450 386.550 -42.190 ;
        RECT 388.850 -42.240 392.200 -42.010 ;
        RECT 384.905 -42.500 386.540 -42.450 ;
        RECT 382.970 -43.160 385.470 -42.930 ;
        RECT 384.780 -44.640 385.010 -43.390 ;
        RECT 385.240 -43.655 385.470 -43.160 ;
        RECT 385.995 -43.310 386.540 -42.500 ;
        RECT 387.445 -42.610 388.250 -42.270 ;
        RECT 385.240 -43.885 387.205 -43.655 ;
        RECT 385.240 -44.410 385.470 -43.885 ;
        RECT 385.735 -44.530 387.005 -44.300 ;
        RECT 387.445 -44.410 387.785 -42.610 ;
        RECT 388.850 -42.840 389.080 -42.240 ;
        RECT 388.080 -43.070 389.080 -42.840 ;
        RECT 388.080 -44.005 388.310 -43.070 ;
        RECT 389.310 -43.300 389.650 -42.480 ;
        RECT 390.045 -43.070 390.275 -42.240 ;
        RECT 390.870 -43.090 391.210 -42.480 ;
        RECT 391.970 -42.630 392.200 -42.240 ;
        RECT 391.970 -42.860 395.155 -42.630 ;
        RECT 394.925 -43.070 395.155 -42.860 ;
        RECT 388.760 -43.530 389.650 -43.300 ;
        RECT 390.530 -43.320 394.510 -43.090 ;
        RECT 385.735 -44.640 385.965 -44.530 ;
        RECT 384.780 -44.870 385.965 -44.640 ;
        RECT 386.775 -44.640 387.005 -44.530 ;
        RECT 388.760 -44.640 388.990 -43.530 ;
        RECT 390.530 -44.325 390.760 -43.320 ;
        RECT 395.505 -43.550 395.735 -42.270 ;
        RECT 402.470 -42.290 402.730 -42.130 ;
        RECT 396.570 -42.555 396.975 -42.325 ;
        RECT 391.045 -43.780 396.055 -43.550 ;
        RECT 391.045 -44.005 391.345 -43.780 ;
        RECT 390.120 -44.555 390.760 -44.325 ;
        RECT 392.205 -44.240 395.035 -44.010 ;
        RECT 395.825 -44.240 396.055 -43.780 ;
        RECT 392.205 -44.610 392.435 -44.240 ;
        RECT 394.805 -44.435 395.035 -44.240 ;
        RECT 396.285 -44.470 396.515 -43.390 ;
        RECT 396.745 -43.900 396.975 -42.555 ;
        RECT 398.430 -42.575 398.935 -42.345 ;
        RECT 397.280 -43.630 398.310 -43.250 ;
        RECT 398.705 -43.865 398.935 -42.575 ;
        RECT 400.725 -42.760 400.955 -42.290 ;
        RECT 396.745 -44.240 397.075 -43.900 ;
        RECT 397.305 -44.095 398.935 -43.865 ;
        RECT 397.305 -44.470 397.535 -44.095 ;
        RECT 386.775 -44.870 388.990 -44.640 ;
        RECT 396.285 -44.700 397.535 -44.470 ;
        RECT 398.585 -44.695 398.935 -44.095 ;
        RECT 399.165 -42.990 400.955 -42.760 ;
        RECT 399.165 -43.885 399.395 -42.990 ;
        RECT 399.630 -43.630 401.050 -43.250 ;
        RECT 399.165 -44.115 400.855 -43.885 ;
        RECT 400.625 -44.705 400.855 -44.115 ;
        RECT 402.460 -44.190 402.795 -42.290 ;
        RECT 403.685 -43.035 404.960 -42.805 ;
        RECT 403.685 -44.870 403.915 -43.035 ;
        RECT 405.205 -43.440 405.435 -42.010 ;
        RECT 404.170 -43.670 405.435 -43.440 ;
        RECT 406.385 -44.430 406.710 -42.450 ;
        RECT 406.940 -44.850 407.275 -42.080 ;
        RECT 409.190 -42.290 409.450 -42.130 ;
        RECT 409.180 -44.190 409.515 -42.290 ;
        RECT 410.405 -43.035 411.680 -42.805 ;
        RECT 410.405 -44.870 410.635 -43.035 ;
        RECT 411.925 -43.440 412.155 -42.010 ;
        RECT 410.890 -43.670 412.155 -43.440 ;
        RECT 414.885 -43.035 416.160 -42.805 ;
        RECT 414.885 -44.870 415.115 -43.035 ;
        RECT 416.405 -43.440 416.635 -42.010 ;
        RECT 417.590 -42.290 417.850 -42.130 ;
        RECT 415.370 -43.670 416.635 -43.440 ;
        RECT 417.525 -44.190 417.860 -42.290 ;
        RECT 418.705 -44.430 419.030 -42.450 ;
        RECT 419.260 -44.850 419.595 -42.080 ;
        RECT 429.240 -42.240 432.590 -42.010 ;
        RECT 420.485 -42.760 420.715 -42.290 ;
        RECT 422.505 -42.575 423.010 -42.345 ;
        RECT 424.465 -42.555 424.870 -42.325 ;
        RECT 420.485 -42.990 422.275 -42.760 ;
        RECT 420.520 -43.630 421.810 -43.250 ;
        RECT 422.045 -43.885 422.275 -42.990 ;
        RECT 420.585 -44.115 422.275 -43.885 ;
        RECT 422.505 -43.865 422.735 -42.575 ;
        RECT 423.130 -43.630 424.160 -43.250 ;
        RECT 422.505 -44.095 424.135 -43.865 ;
        RECT 424.465 -43.900 424.695 -42.555 ;
        RECT 420.585 -44.705 420.815 -44.115 ;
        RECT 422.505 -44.695 422.855 -44.095 ;
        RECT 423.905 -44.470 424.135 -44.095 ;
        RECT 424.365 -44.240 424.695 -43.900 ;
        RECT 424.925 -44.470 425.155 -43.390 ;
        RECT 425.705 -43.550 425.935 -42.270 ;
        RECT 429.240 -42.630 429.470 -42.240 ;
        RECT 426.285 -42.860 429.470 -42.630 ;
        RECT 426.285 -43.070 426.515 -42.860 ;
        RECT 430.230 -43.090 430.570 -42.480 ;
        RECT 431.165 -43.070 431.395 -42.240 ;
        RECT 426.930 -43.320 430.910 -43.090 ;
        RECT 425.385 -43.780 430.395 -43.550 ;
        RECT 425.385 -44.240 425.615 -43.780 ;
        RECT 430.095 -44.005 430.395 -43.780 ;
        RECT 426.405 -44.240 429.235 -44.010 ;
        RECT 426.405 -44.435 426.635 -44.240 ;
        RECT 423.905 -44.700 425.155 -44.470 ;
        RECT 429.005 -44.610 429.235 -44.240 ;
        RECT 430.680 -44.325 430.910 -43.320 ;
        RECT 431.790 -43.300 432.130 -42.480 ;
        RECT 432.360 -42.840 432.590 -42.240 ;
        RECT 433.190 -42.610 433.995 -42.270 ;
        RECT 432.360 -43.070 433.360 -42.840 ;
        RECT 431.790 -43.530 432.680 -43.300 ;
        RECT 430.680 -44.555 431.320 -44.325 ;
        RECT 432.450 -44.640 432.680 -43.530 ;
        RECT 433.130 -44.005 433.360 -43.070 ;
        RECT 433.655 -44.410 433.995 -42.610 ;
        RECT 434.900 -42.500 436.535 -42.140 ;
        RECT 434.900 -43.310 435.445 -42.500 ;
        RECT 436.890 -42.930 437.120 -42.270 ;
        RECT 435.970 -43.160 438.470 -42.930 ;
        RECT 435.970 -43.655 436.200 -43.160 ;
        RECT 434.235 -43.885 436.200 -43.655 ;
        RECT 434.435 -44.530 435.705 -44.300 ;
        RECT 435.970 -44.410 436.200 -43.885 ;
        RECT 434.435 -44.640 434.665 -44.530 ;
        RECT 432.450 -44.870 434.665 -44.640 ;
        RECT 435.475 -44.640 435.705 -44.530 ;
        RECT 436.430 -44.640 436.660 -43.390 ;
        RECT 435.475 -44.870 436.660 -44.640 ;
        RECT 438.715 -44.860 439.150 -42.030 ;
        RECT 441.105 -44.430 441.430 -42.450 ;
        RECT 441.660 -44.850 441.995 -42.080 ;
        RECT 443.910 -42.290 444.170 -42.130 ;
        RECT 443.900 -44.190 444.235 -42.290 ;
        RECT 445.125 -43.035 446.400 -42.805 ;
        RECT 445.125 -44.870 445.355 -43.035 ;
        RECT 446.645 -43.440 446.875 -42.010 ;
        RECT 445.610 -43.670 446.875 -43.440 ;
        RECT 447.365 -43.035 448.640 -42.805 ;
        RECT 447.365 -44.870 447.595 -43.035 ;
        RECT 448.885 -43.440 449.115 -42.010 ;
        RECT 450.070 -42.290 450.330 -42.130 ;
        RECT 447.850 -43.670 449.115 -43.440 ;
        RECT 450.005 -44.190 450.340 -42.290 ;
        RECT 454.485 -44.870 454.815 -42.010 ;
        RECT 455.045 -43.680 455.370 -42.680 ;
        RECT 458.190 -43.085 458.780 -42.045 ;
        RECT 458.190 -44.800 458.555 -43.085 ;
        RECT 458.850 -44.000 459.190 -43.360 ;
        RECT 460.645 -44.000 460.875 -42.045 ;
        RECT 458.850 -44.235 460.875 -44.000 ;
        RECT 460.545 -44.860 460.875 -44.235 ;
        RECT 300.585 -46.610 300.815 -45.940 ;
        RECT 302.825 -46.610 303.055 -45.940 ;
        RECT 305.065 -46.610 305.295 -45.940 ;
        RECT 307.205 -46.610 307.435 -45.940 ;
        RECT 309.545 -46.560 309.775 -45.940 ;
        RECT 311.785 -46.560 312.015 -45.940 ;
        RECT 300.550 -46.990 307.435 -46.610 ;
        RECT 308.965 -46.790 312.015 -46.560 ;
        RECT 317.905 -46.560 318.135 -45.940 ;
        RECT 320.145 -46.560 320.375 -45.940 ;
        RECT 317.905 -46.790 320.955 -46.560 ;
        RECT 299.740 -47.635 302.940 -47.290 ;
        RECT 303.640 -47.900 304.440 -46.990 ;
        RECT 308.965 -47.295 309.300 -46.790 ;
        RECT 305.010 -47.635 309.300 -47.295 ;
        RECT 309.770 -47.605 312.630 -47.170 ;
        RECT 317.290 -47.605 320.150 -47.170 ;
        RECT 320.620 -47.295 320.955 -46.790 ;
        RECT 322.485 -46.610 322.715 -45.940 ;
        RECT 324.625 -46.610 324.855 -45.940 ;
        RECT 326.865 -46.610 327.095 -45.940 ;
        RECT 329.105 -46.610 329.335 -45.940 ;
        RECT 336.385 -46.560 336.615 -45.940 ;
        RECT 338.625 -46.560 338.855 -45.940 ;
        RECT 322.485 -46.990 329.335 -46.610 ;
        RECT 300.485 -48.280 307.435 -47.900 ;
        RECT 300.485 -48.645 300.715 -48.280 ;
        RECT 302.725 -48.645 302.955 -48.280 ;
        RECT 304.965 -48.645 305.195 -48.280 ;
        RECT 307.175 -48.645 307.435 -48.280 ;
        RECT 308.965 -48.070 309.300 -47.635 ;
        RECT 320.620 -47.635 324.910 -47.295 ;
        RECT 320.620 -48.070 320.955 -47.635 ;
        RECT 325.480 -47.900 326.280 -46.990 ;
        RECT 326.980 -47.635 330.180 -47.290 ;
        RECT 308.965 -48.305 311.915 -48.070 ;
        RECT 309.445 -48.645 309.675 -48.305 ;
        RECT 311.685 -48.645 311.915 -48.305 ;
        RECT 318.005 -48.305 320.955 -48.070 ;
        RECT 322.485 -48.280 329.435 -47.900 ;
        RECT 322.485 -48.290 322.745 -48.280 ;
        RECT 318.005 -48.645 318.235 -48.305 ;
        RECT 320.245 -48.645 320.475 -48.305 ;
        RECT 322.390 -48.645 322.745 -48.290 ;
        RECT 324.725 -48.645 324.955 -48.280 ;
        RECT 326.965 -48.645 327.195 -48.280 ;
        RECT 329.205 -48.645 329.435 -48.280 ;
        RECT 333.525 -48.510 333.860 -46.610 ;
        RECT 336.385 -46.790 339.435 -46.560 ;
        RECT 340.965 -46.610 341.195 -45.940 ;
        RECT 343.105 -46.610 343.335 -45.940 ;
        RECT 345.345 -46.610 345.575 -45.940 ;
        RECT 347.585 -46.610 347.815 -45.940 ;
        RECT 335.770 -47.605 338.630 -47.170 ;
        RECT 339.100 -47.295 339.435 -46.790 ;
        RECT 340.870 -46.990 347.815 -46.610 ;
        RECT 339.100 -47.635 343.390 -47.295 ;
        RECT 339.100 -48.070 339.435 -47.635 ;
        RECT 343.960 -47.900 344.760 -46.990 ;
        RECT 345.460 -47.635 348.660 -47.290 ;
        RECT 349.925 -47.765 350.155 -45.930 ;
        RECT 355.425 -46.560 355.655 -45.940 ;
        RECT 357.665 -46.560 357.895 -45.940 ;
        RECT 350.410 -47.360 351.675 -47.130 ;
        RECT 336.485 -48.305 339.435 -48.070 ;
        RECT 340.965 -48.280 347.915 -47.900 ;
        RECT 349.925 -47.995 351.200 -47.765 ;
        RECT 336.485 -48.645 336.715 -48.305 ;
        RECT 338.725 -48.645 338.955 -48.305 ;
        RECT 340.965 -48.645 341.225 -48.280 ;
        RECT 343.205 -48.645 343.435 -48.280 ;
        RECT 345.445 -48.645 345.675 -48.280 ;
        RECT 347.685 -48.645 347.915 -48.280 ;
        RECT 322.390 -48.670 322.650 -48.645 ;
        RECT 351.445 -48.790 351.675 -47.360 ;
        RECT 352.565 -48.510 352.900 -46.610 ;
        RECT 355.425 -46.790 358.475 -46.560 ;
        RECT 360.005 -46.610 360.235 -45.940 ;
        RECT 362.145 -46.610 362.375 -45.940 ;
        RECT 364.385 -46.610 364.615 -45.940 ;
        RECT 366.625 -46.610 366.855 -45.940 ;
        RECT 354.810 -47.605 357.670 -47.170 ;
        RECT 358.140 -47.295 358.475 -46.790 ;
        RECT 359.910 -46.990 366.855 -46.610 ;
        RECT 358.140 -47.635 362.430 -47.295 ;
        RECT 358.140 -48.070 358.475 -47.635 ;
        RECT 363.000 -47.900 363.800 -46.990 ;
        RECT 364.500 -47.635 367.700 -47.290 ;
        RECT 368.965 -47.765 369.195 -45.930 ;
        RECT 374.465 -46.560 374.695 -45.940 ;
        RECT 376.705 -46.560 376.935 -45.940 ;
        RECT 374.465 -46.790 377.515 -46.560 ;
        RECT 369.450 -47.360 370.715 -47.130 ;
        RECT 355.525 -48.305 358.475 -48.070 ;
        RECT 360.005 -48.280 366.955 -47.900 ;
        RECT 368.965 -47.995 370.240 -47.765 ;
        RECT 355.525 -48.645 355.755 -48.305 ;
        RECT 357.765 -48.645 357.995 -48.305 ;
        RECT 360.005 -48.645 360.265 -48.280 ;
        RECT 362.245 -48.645 362.475 -48.280 ;
        RECT 364.485 -48.645 364.715 -48.280 ;
        RECT 366.725 -48.645 366.955 -48.280 ;
        RECT 370.485 -48.790 370.715 -47.360 ;
        RECT 373.850 -47.605 376.710 -47.170 ;
        RECT 377.180 -47.295 377.515 -46.790 ;
        RECT 379.045 -46.610 379.275 -45.940 ;
        RECT 381.185 -46.610 381.415 -45.940 ;
        RECT 383.425 -46.610 383.655 -45.940 ;
        RECT 385.665 -46.610 385.895 -45.940 ;
        RECT 379.045 -46.990 385.895 -46.610 ;
        RECT 377.180 -47.635 381.470 -47.295 ;
        RECT 377.180 -48.070 377.515 -47.635 ;
        RECT 382.040 -47.790 382.840 -46.990 ;
        RECT 383.540 -47.635 386.740 -47.290 ;
        RECT 381.690 -47.900 382.840 -47.790 ;
        RECT 374.565 -48.305 377.515 -48.070 ;
        RECT 379.045 -48.280 385.995 -47.900 ;
        RECT 374.565 -48.645 374.795 -48.305 ;
        RECT 376.805 -48.645 377.035 -48.305 ;
        RECT 379.045 -48.645 379.305 -48.280 ;
        RECT 381.285 -48.645 381.515 -48.280 ;
        RECT 383.525 -48.645 383.755 -48.280 ;
        RECT 385.765 -48.645 385.995 -48.280 ;
        RECT 389.025 -48.350 389.350 -46.370 ;
        RECT 389.580 -48.720 389.915 -45.950 ;
        RECT 393.505 -46.560 393.735 -45.940 ;
        RECT 395.745 -46.560 395.975 -45.940 ;
        RECT 393.505 -46.790 396.555 -46.560 ;
        RECT 392.890 -47.605 395.750 -47.170 ;
        RECT 396.220 -47.295 396.555 -46.790 ;
        RECT 398.085 -46.610 398.315 -45.940 ;
        RECT 400.225 -46.610 400.455 -45.940 ;
        RECT 402.465 -46.610 402.695 -45.940 ;
        RECT 404.705 -46.610 404.935 -45.940 ;
        RECT 398.085 -46.990 404.935 -46.610 ;
        RECT 396.220 -47.635 400.510 -47.295 ;
        RECT 396.220 -48.070 396.555 -47.635 ;
        RECT 401.080 -47.900 401.880 -46.990 ;
        RECT 402.580 -47.635 405.780 -47.290 ;
        RECT 407.045 -47.765 407.275 -45.930 ;
        RECT 412.545 -46.560 412.775 -45.940 ;
        RECT 414.785 -46.560 415.015 -45.940 ;
        RECT 412.545 -46.790 415.595 -46.560 ;
        RECT 417.125 -46.610 417.355 -45.940 ;
        RECT 419.265 -46.610 419.495 -45.940 ;
        RECT 421.505 -46.610 421.735 -45.940 ;
        RECT 423.745 -46.610 423.975 -45.940 ;
        RECT 407.530 -47.360 408.795 -47.130 ;
        RECT 393.605 -48.305 396.555 -48.070 ;
        RECT 398.085 -48.280 405.035 -47.900 ;
        RECT 407.045 -47.995 408.320 -47.765 ;
        RECT 393.605 -48.645 393.835 -48.305 ;
        RECT 395.845 -48.645 396.075 -48.305 ;
        RECT 398.085 -48.645 398.345 -48.280 ;
        RECT 400.325 -48.645 400.555 -48.280 ;
        RECT 402.565 -48.645 402.795 -48.280 ;
        RECT 404.805 -48.645 405.035 -48.280 ;
        RECT 408.565 -48.790 408.795 -47.360 ;
        RECT 411.930 -47.605 414.790 -47.170 ;
        RECT 415.260 -47.295 415.595 -46.790 ;
        RECT 417.030 -46.990 423.975 -46.610 ;
        RECT 415.260 -47.635 419.550 -47.295 ;
        RECT 415.260 -48.070 415.595 -47.635 ;
        RECT 420.120 -47.900 420.920 -46.990 ;
        RECT 421.620 -47.635 424.820 -47.290 ;
        RECT 426.085 -47.765 426.315 -45.930 ;
        RECT 431.585 -46.560 431.815 -45.940 ;
        RECT 433.825 -46.560 434.055 -45.940 ;
        RECT 431.585 -46.790 434.635 -46.560 ;
        RECT 436.165 -46.610 436.395 -45.940 ;
        RECT 438.305 -46.610 438.535 -45.940 ;
        RECT 440.545 -46.610 440.775 -45.940 ;
        RECT 442.785 -46.610 443.015 -45.940 ;
        RECT 426.570 -47.360 427.835 -47.130 ;
        RECT 412.645 -48.305 415.595 -48.070 ;
        RECT 417.125 -48.280 424.075 -47.900 ;
        RECT 426.085 -47.995 427.360 -47.765 ;
        RECT 412.645 -48.645 412.875 -48.305 ;
        RECT 414.885 -48.645 415.115 -48.305 ;
        RECT 417.125 -48.645 417.385 -48.280 ;
        RECT 419.365 -48.645 419.595 -48.280 ;
        RECT 421.605 -48.645 421.835 -48.280 ;
        RECT 423.845 -48.645 424.075 -48.280 ;
        RECT 427.605 -48.790 427.835 -47.360 ;
        RECT 430.970 -47.605 433.830 -47.170 ;
        RECT 434.300 -47.295 434.635 -46.790 ;
        RECT 436.070 -46.990 443.015 -46.610 ;
        RECT 434.300 -47.635 438.590 -47.295 ;
        RECT 434.300 -48.070 434.635 -47.635 ;
        RECT 439.160 -47.900 439.960 -46.990 ;
        RECT 440.660 -47.635 443.860 -47.290 ;
        RECT 445.125 -47.765 445.355 -45.930 ;
        RECT 454.645 -46.565 454.975 -45.940 ;
        RECT 445.610 -47.360 446.875 -47.130 ;
        RECT 431.685 -48.305 434.635 -48.070 ;
        RECT 436.165 -48.280 443.115 -47.900 ;
        RECT 445.125 -47.995 446.400 -47.765 ;
        RECT 431.685 -48.645 431.915 -48.305 ;
        RECT 433.925 -48.645 434.155 -48.305 ;
        RECT 436.165 -48.645 436.425 -48.280 ;
        RECT 438.405 -48.645 438.635 -48.280 ;
        RECT 440.645 -48.645 440.875 -48.280 ;
        RECT 442.885 -48.645 443.115 -48.280 ;
        RECT 446.645 -48.790 446.875 -47.360 ;
        RECT 453.925 -48.510 454.260 -46.610 ;
        RECT 454.645 -46.800 456.670 -46.565 ;
        RECT 454.645 -48.755 454.875 -46.800 ;
        RECT 456.330 -47.440 456.670 -46.800 ;
        RECT 456.965 -47.715 457.330 -46.000 ;
        RECT 456.740 -48.755 457.330 -47.715 ;
        RECT 458.190 -47.715 458.555 -46.000 ;
        RECT 460.545 -46.565 460.875 -45.940 ;
        RECT 458.850 -46.800 460.875 -46.565 ;
        RECT 458.850 -47.440 459.190 -46.800 ;
        RECT 458.190 -48.755 458.780 -47.715 ;
        RECT 460.645 -48.755 460.875 -46.800 ;
        RECT 143.575 -64.140 144.605 -63.690 ;
        RECT 144.285 -64.850 144.605 -64.140 ;
        RECT 144.845 -64.620 145.260 -63.100 ;
        RECT 145.490 -64.095 146.435 -63.865 ;
        RECT 145.490 -64.850 145.745 -64.095 ;
        RECT 144.285 -65.150 145.745 -64.850 ;
        RECT 143.575 -67.500 144.605 -67.050 ;
        RECT 144.285 -68.210 144.605 -67.500 ;
        RECT 144.845 -67.980 145.260 -66.460 ;
        RECT 145.490 -67.455 146.435 -67.225 ;
        RECT 145.490 -68.210 145.745 -67.455 ;
        RECT 144.285 -68.510 145.745 -68.210 ;
        RECT 143.575 -70.860 144.605 -70.410 ;
        RECT 144.285 -71.570 144.605 -70.860 ;
        RECT 144.845 -71.340 145.260 -69.820 ;
        RECT 145.490 -70.815 146.435 -70.585 ;
        RECT 145.490 -71.570 145.745 -70.815 ;
        RECT 144.285 -71.870 145.745 -71.570 ;
        RECT 143.575 -74.220 144.605 -73.770 ;
        RECT 144.285 -74.930 144.605 -74.220 ;
        RECT 144.845 -74.700 145.260 -73.180 ;
        RECT 145.490 -74.175 146.435 -73.945 ;
        RECT 145.490 -74.930 145.745 -74.175 ;
        RECT 144.285 -75.230 145.745 -74.930 ;
        RECT 143.575 -77.580 144.605 -77.130 ;
        RECT 144.285 -78.290 144.605 -77.580 ;
        RECT 144.845 -78.060 145.260 -76.540 ;
        RECT 145.490 -77.535 146.435 -77.305 ;
        RECT 145.490 -78.290 145.745 -77.535 ;
        RECT 144.285 -78.590 145.745 -78.290 ;
        RECT -484.745 -79.315 -483.845 -79.275 ;
        RECT -494.430 -79.615 -483.845 -79.315 ;
        RECT -494.430 -81.640 -492.560 -79.615 ;
        RECT -484.745 -79.655 -483.845 -79.615 ;
        RECT 143.575 -80.940 144.605 -80.490 ;
        RECT -492.330 -82.430 -492.100 -81.795 ;
        RECT -492.330 -82.660 -489.660 -82.430 ;
        RECT -492.330 -83.295 -492.100 -82.660 ;
        RECT -497.595 -83.450 -495.515 -83.365 ;
        RECT -497.595 -83.680 -492.560 -83.450 ;
        RECT -497.595 -83.765 -495.515 -83.680 ;
        RECT -492.330 -84.395 -492.100 -83.835 ;
        RECT -492.330 -84.775 -491.430 -84.395 ;
        RECT -492.330 -85.335 -492.100 -84.775 ;
        RECT -494.430 -85.720 -492.560 -85.490 ;
        RECT -494.430 -86.965 -492.560 -86.510 ;
        RECT -491.110 -86.965 -490.880 -82.660 ;
        RECT -489.890 -85.335 -489.660 -82.660 ;
        RECT -486.955 -83.235 -486.555 -81.155 ;
        RECT 144.285 -81.650 144.605 -80.940 ;
        RECT 144.845 -81.420 145.260 -79.900 ;
        RECT 145.490 -80.895 146.435 -80.665 ;
        RECT 145.490 -81.650 145.745 -80.895 ;
        RECT 144.285 -81.950 145.745 -81.650 ;
        RECT -486.870 -85.490 -486.640 -83.235 ;
        RECT 143.575 -84.300 144.605 -83.850 ;
        RECT 144.285 -85.010 144.605 -84.300 ;
        RECT 144.845 -84.780 145.260 -83.260 ;
        RECT 145.490 -84.255 146.435 -84.025 ;
        RECT 145.490 -85.010 145.745 -84.255 ;
        RECT 144.285 -85.310 145.745 -85.010 ;
        RECT -490.615 -85.875 -490.235 -85.665 ;
        RECT -489.430 -85.720 -486.640 -85.490 ;
        RECT -490.615 -86.355 -489.660 -85.875 ;
        RECT -490.615 -86.565 -490.235 -86.355 ;
        RECT -489.430 -86.965 -487.560 -86.510 ;
        RECT -494.430 -87.265 -487.560 -86.965 ;
        RECT -486.870 -87.105 -486.640 -85.720 ;
        RECT 143.575 -87.660 144.605 -87.210 ;
        RECT 144.285 -88.370 144.605 -87.660 ;
        RECT 144.845 -88.140 145.260 -86.620 ;
        RECT 145.490 -87.615 146.435 -87.385 ;
        RECT 145.490 -88.370 145.745 -87.615 ;
        RECT 144.285 -88.670 145.745 -88.370 ;
        RECT 143.575 -91.020 144.605 -90.570 ;
        RECT 144.285 -91.730 144.605 -91.020 ;
        RECT 144.845 -91.500 145.260 -89.980 ;
        RECT 145.490 -90.975 146.435 -90.745 ;
        RECT 145.490 -91.730 145.745 -90.975 ;
        RECT 144.285 -92.030 145.745 -91.730 ;
        RECT 143.575 -94.380 144.605 -93.930 ;
        RECT 144.285 -95.090 144.605 -94.380 ;
        RECT 144.845 -94.860 145.260 -93.340 ;
        RECT 145.490 -94.335 146.435 -94.105 ;
        RECT 145.490 -95.090 145.745 -94.335 ;
        RECT 144.285 -95.390 145.745 -95.090 ;
        RECT -493.475 -95.830 -492.575 -95.450 ;
        RECT -489.445 -95.830 -488.545 -95.450 ;
        RECT -491.830 -95.945 -491.430 -95.830 ;
        RECT -492.345 -96.285 -489.675 -95.945 ;
        RECT -491.830 -98.115 -491.430 -96.285 ;
        RECT 143.575 -97.740 144.605 -97.290 ;
        RECT 144.285 -98.450 144.605 -97.740 ;
        RECT 145.490 -97.695 146.435 -97.465 ;
        RECT 145.490 -98.450 145.745 -97.695 ;
        RECT 144.285 -98.750 145.745 -98.450 ;
      LAYER Via1 ;
        RECT -491.760 97.205 -491.500 97.985 ;
        RECT 143.665 97.385 143.925 97.645 ;
        RECT -493.415 95.510 -492.635 95.770 ;
        RECT -489.385 95.510 -488.605 95.770 ;
        RECT 143.665 94.025 143.925 94.285 ;
        RECT 144.920 93.500 145.180 93.760 ;
        RECT 143.665 90.665 143.925 90.925 ;
        RECT 144.920 90.140 145.180 90.400 ;
        RECT 143.665 87.305 143.925 87.565 ;
        RECT -492.270 84.455 -491.490 84.715 ;
        RECT -497.465 83.435 -495.645 83.695 ;
        RECT -490.555 85.725 -490.295 86.505 ;
        RECT 144.920 86.780 145.180 87.040 ;
        RECT 143.665 83.945 143.925 84.205 ;
        RECT 144.920 83.420 145.180 83.680 ;
        RECT -486.885 81.285 -486.625 83.105 ;
        RECT 143.665 80.585 143.925 80.845 ;
        RECT 144.920 80.060 145.180 80.320 ;
        RECT -484.685 79.335 -483.905 79.595 ;
        RECT 143.665 77.225 143.925 77.485 ;
        RECT 144.920 76.700 145.180 76.960 ;
        RECT 143.665 73.865 143.925 74.125 ;
        RECT 144.920 73.340 145.180 73.600 ;
        RECT 143.665 70.505 143.925 70.765 ;
        RECT 144.920 69.980 145.180 70.240 ;
        RECT 143.665 67.145 143.925 67.405 ;
        RECT 144.920 66.620 145.180 66.880 ;
        RECT 143.665 63.785 143.925 64.045 ;
        RECT 144.920 63.260 145.180 63.520 ;
        RECT 300.550 47.710 300.810 47.970 ;
        RECT 322.390 47.710 322.650 47.970 ;
        RECT 310.070 46.590 310.330 46.850 ;
        RECT 319.030 46.590 319.290 46.850 ;
        RECT 336.950 47.710 337.210 47.970 ;
        RECT 346.470 46.590 346.730 46.850 ;
        RECT 359.910 47.710 360.170 47.970 ;
        RECT 354.870 46.590 355.130 46.850 ;
        RECT 375.030 47.710 375.290 47.970 ;
        RECT 394.070 47.710 394.330 47.970 ;
        RECT 384.550 46.590 384.810 46.850 ;
        RECT 417.030 47.710 417.290 47.970 ;
        RECT 405.830 46.590 406.090 46.850 ;
        RECT 389.030 45.470 389.290 45.730 ;
        RECT 411.990 46.590 412.250 46.850 ;
        RECT 432.150 47.710 432.410 47.970 ;
        RECT 408.070 45.470 408.330 45.730 ;
        RECT 426.550 46.030 426.810 46.290 ;
        RECT 427.110 45.470 427.370 45.730 ;
        RECT 428.230 46.590 428.490 46.850 ;
        RECT 443.910 46.590 444.170 46.850 ;
        RECT 446.150 45.470 446.410 45.730 ;
        RECT 298.870 42.110 299.130 42.370 ;
        RECT 310.630 42.670 310.890 42.930 ;
        RECT 312.310 42.670 312.570 42.930 ;
        RECT 312.870 42.110 313.130 42.370 ;
        RECT 315.110 42.110 315.370 42.370 ;
        RECT 317.350 42.110 317.610 42.370 ;
        RECT 319.590 42.110 319.850 42.370 ;
        RECT 314.550 41.550 314.810 41.810 ;
        RECT 334.150 43.230 334.410 43.490 ;
        RECT 338.070 42.110 338.330 42.370 ;
        RECT 340.870 43.790 341.130 44.050 ;
        RECT 333.590 41.550 333.850 41.810 ;
        RECT 339.190 41.550 339.450 41.810 ;
        RECT 342.550 43.790 342.810 44.050 ;
        RECT 344.230 43.790 344.490 44.050 ;
        RECT 349.830 43.230 350.090 43.490 ;
        RECT 350.390 41.550 350.650 41.810 ;
        RECT 352.070 43.790 352.330 44.050 ;
        RECT 353.750 43.790 354.010 44.050 ;
        RECT 355.430 42.670 355.690 42.930 ;
        RECT 358.790 42.670 359.050 42.930 ;
        RECT 369.990 43.230 370.250 43.490 ;
        RECT 373.910 41.550 374.170 41.810 ;
        RECT 376.150 43.790 376.410 44.050 ;
        RECT 377.830 41.550 378.090 41.810 ;
        RECT 378.950 42.110 379.210 42.370 ;
        RECT 381.750 42.110 382.010 42.370 ;
        RECT 383.990 42.670 384.250 42.930 ;
        RECT 385.670 42.670 385.930 42.930 ;
        RECT 386.790 42.670 387.050 42.930 ;
        RECT 387.910 42.670 388.170 42.930 ;
        RECT 392.390 43.790 392.650 44.050 ;
        RECT 389.030 42.670 389.290 42.930 ;
        RECT 387.350 42.110 387.610 42.370 ;
        RECT 391.830 42.110 392.090 42.370 ;
        RECT 394.070 42.670 394.330 42.930 ;
        RECT 396.870 42.670 397.130 42.930 ;
        RECT 408.630 43.230 408.890 43.490 ;
        RECT 415.350 42.670 415.610 42.930 ;
        RECT 416.470 42.670 416.730 42.930 ;
        RECT 422.070 43.790 422.330 44.050 ;
        RECT 418.710 42.670 418.970 42.930 ;
        RECT 419.830 42.670 420.090 42.930 ;
        RECT 420.950 42.670 421.210 42.930 ;
        RECT 412.550 41.550 412.810 41.810 ;
        RECT 417.590 42.110 417.850 42.370 ;
        RECT 423.190 42.670 423.450 42.930 ;
        RECT 424.870 41.550 425.130 41.810 ;
        RECT 428.790 43.230 429.050 43.490 ;
        RECT 439.990 42.670 440.250 42.930 ;
        RECT 443.350 42.670 443.610 42.930 ;
        RECT 444.470 42.110 444.730 42.370 ;
        RECT 445.590 43.230 445.850 43.490 ;
        RECT 448.390 42.110 448.650 42.370 ;
        RECT 446.150 41.550 446.410 41.810 ;
        RECT 298.870 39.310 299.130 39.570 ;
        RECT 312.870 39.310 313.130 39.570 ;
        RECT 308.390 38.750 308.650 39.010 ;
        RECT 318.470 38.750 318.730 39.010 ;
        RECT 321.830 38.750 322.090 39.010 ;
        RECT 336.950 39.310 337.210 39.570 ;
        RECT 333.030 37.630 333.290 37.890 ;
        RECT 338.070 38.750 338.330 39.010 ;
        RECT 339.190 38.750 339.450 39.010 ;
        RECT 339.750 37.630 340.010 37.890 ;
        RECT 341.430 38.750 341.690 39.010 ;
        RECT 343.670 37.630 343.930 37.890 ;
        RECT 361.030 39.870 361.290 40.130 ;
        RECT 361.590 38.190 361.850 38.450 ;
        RECT 363.270 38.750 363.530 39.010 ;
        RECT 364.390 37.630 364.650 37.890 ;
        RECT 364.950 38.190 365.210 38.450 ;
        RECT 365.510 38.750 365.770 39.010 ;
        RECT 366.070 37.630 366.330 37.890 ;
        RECT 386.230 39.870 386.490 40.130 ;
        RECT 387.910 38.750 388.170 39.010 ;
        RECT 389.030 39.310 389.290 39.570 ;
        RECT 390.710 38.190 390.970 38.450 ;
        RECT 391.270 37.630 391.530 37.890 ;
        RECT 404.710 38.750 404.970 39.010 ;
        RECT 427.110 39.310 427.370 39.570 ;
        RECT 437.190 39.310 437.450 39.570 ;
        RECT 431.590 38.750 431.850 39.010 ;
        RECT 434.950 38.750 435.210 39.010 ;
        RECT 436.070 38.750 436.330 39.010 ;
        RECT 439.430 39.310 439.690 39.570 ;
        RECT 437.750 38.190 438.010 38.450 ;
        RECT 439.990 39.310 440.250 39.570 ;
        RECT 441.110 38.750 441.370 39.010 ;
        RECT 442.230 37.630 442.490 37.890 ;
        RECT 446.150 37.630 446.410 37.890 ;
        RECT 457.350 38.750 457.610 39.010 ;
        RECT 459.590 38.750 459.850 39.010 ;
        RECT 168.175 34.310 168.435 35.090 ;
        RECT 174.175 34.310 174.435 35.090 ;
        RECT 178.105 34.375 178.365 35.155 ;
        RECT 180.245 34.375 180.505 35.155 ;
        RECT 186.675 34.310 186.935 35.090 ;
        RECT 299.430 34.270 299.690 34.530 ;
        RECT 310.630 34.830 310.890 35.090 ;
        RECT 337.510 35.390 337.770 35.650 ;
        RECT 338.070 35.390 338.330 35.650 ;
        RECT 338.630 35.390 338.890 35.650 ;
        RECT 341.990 34.830 342.250 35.090 ;
        RECT 340.870 34.270 341.130 34.530 ;
        RECT 345.350 34.830 345.610 35.090 ;
        RECT 356.550 35.390 356.810 35.650 ;
        RECT 360.470 35.950 360.730 36.210 ;
        RECT 361.590 34.830 361.850 35.090 ;
        RECT 362.710 34.830 362.970 35.090 ;
        RECT 363.830 35.950 364.090 36.210 ;
        RECT 364.390 34.830 364.650 35.090 ;
        RECT 363.270 34.270 363.530 34.530 ;
        RECT 384.550 34.830 384.810 35.090 ;
        RECT 385.670 34.830 385.930 35.090 ;
        RECT 386.230 35.390 386.490 35.650 ;
        RECT 387.910 35.390 388.170 35.650 ;
        RECT 386.790 34.830 387.050 35.090 ;
        RECT 391.270 34.830 391.530 35.090 ;
        RECT 392.950 34.830 393.210 35.090 ;
        RECT 404.710 35.950 404.970 36.210 ;
        RECT 410.310 34.270 410.570 34.530 ;
        RECT 408.630 33.710 408.890 33.970 ;
        RECT 417.030 34.830 417.290 35.090 ;
        RECT 415.350 33.710 415.610 33.970 ;
        RECT 433.830 35.390 434.090 35.650 ;
        RECT 422.070 34.830 422.330 35.090 ;
        RECT 418.150 34.270 418.410 34.530 ;
        RECT 437.750 35.390 438.010 35.650 ;
        RECT 448.950 34.830 449.210 35.090 ;
        RECT 452.310 34.830 452.570 35.090 ;
        RECT 455.670 34.270 455.930 34.530 ;
        RECT 178.650 28.800 178.910 29.580 ;
        RECT 179.770 28.800 180.030 29.580 ;
        RECT 174.170 26.410 174.430 27.190 ;
        RECT 184.250 26.410 184.510 27.190 ;
        RECT 171.930 24.410 172.190 25.190 ;
        RECT 176.410 24.410 176.670 25.190 ;
        RECT 182.010 24.410 182.270 25.190 ;
        RECT 186.490 24.410 186.750 25.190 ;
        RECT 302.790 32.030 303.050 32.290 ;
        RECT 303.350 30.350 303.610 30.610 ;
        RECT 317.350 30.910 317.610 31.170 ;
        RECT 320.150 30.910 320.410 31.170 ;
        RECT 332.470 29.790 332.730 30.050 ;
        RECT 335.270 30.350 335.530 30.610 ;
        RECT 337.510 30.910 337.770 31.170 ;
        RECT 336.390 30.350 336.650 30.610 ;
        RECT 341.430 31.470 341.690 31.730 ;
        RECT 339.750 30.910 340.010 31.170 ;
        RECT 338.630 29.790 338.890 30.050 ;
        RECT 349.270 32.030 349.530 32.290 ;
        RECT 343.670 29.790 343.930 30.050 ;
        RECT 349.830 31.470 350.090 31.730 ;
        RECT 360.470 30.350 360.730 30.610 ;
        RECT 362.150 30.350 362.410 30.610 ;
        RECT 363.270 30.910 363.530 31.170 ;
        RECT 366.630 30.910 366.890 31.170 ;
        RECT 377.830 30.350 378.090 30.610 ;
        RECT 381.750 30.350 382.010 30.610 ;
        RECT 383.430 29.790 383.690 30.050 ;
        RECT 383.990 29.790 384.250 30.050 ;
        RECT 384.550 29.790 384.810 30.050 ;
        RECT 385.110 30.910 385.370 31.170 ;
        RECT 386.230 30.350 386.490 30.610 ;
        RECT 389.590 30.910 389.850 31.170 ;
        RECT 387.910 29.790 388.170 30.050 ;
        RECT 409.190 31.470 409.450 31.730 ;
        RECT 411.430 31.470 411.690 31.730 ;
        RECT 413.670 30.910 413.930 31.170 ;
        RECT 415.910 30.910 416.170 31.170 ;
        RECT 427.110 32.030 427.370 32.290 ;
        RECT 417.590 30.350 417.850 30.610 ;
        RECT 431.590 30.910 431.850 31.170 ;
        RECT 434.390 29.790 434.650 30.050 ;
        RECT 438.310 29.790 438.570 30.050 ;
        RECT 449.510 30.910 449.770 31.170 ;
        RECT 452.870 30.910 453.130 31.170 ;
        RECT 455.110 30.910 455.370 31.170 ;
        RECT 453.990 29.790 454.250 30.050 ;
        RECT 458.470 30.350 458.730 30.610 ;
        RECT 460.150 30.350 460.410 30.610 ;
        RECT 299.990 26.990 300.250 27.250 ;
        RECT 302.790 25.870 303.050 26.130 ;
        RECT 319.030 28.110 319.290 28.370 ;
        RECT 317.910 26.990 318.170 27.250 ;
        RECT 321.270 26.990 321.530 27.250 ;
        RECT 320.710 25.870 320.970 26.130 ;
        RECT 337.510 28.110 337.770 28.370 ;
        RECT 333.030 26.990 333.290 27.250 ;
        RECT 331.350 26.430 331.610 26.690 ;
        RECT 334.150 27.550 334.410 27.810 ;
        RECT 340.310 26.990 340.570 27.250 ;
        RECT 342.550 26.990 342.810 27.250 ;
        RECT 354.870 28.110 355.130 28.370 ;
        RECT 357.670 26.990 357.930 27.250 ;
        RECT 363.270 28.110 363.530 28.370 ;
        RECT 364.950 28.110 365.210 28.370 ;
        RECT 369.430 28.110 369.690 28.370 ;
        RECT 369.990 26.990 370.250 27.250 ;
        RECT 378.950 26.990 379.210 27.250 ;
        RECT 381.190 26.990 381.450 27.250 ;
        RECT 389.030 28.110 389.290 28.370 ;
        RECT 390.710 26.990 390.970 27.250 ;
        RECT 409.190 26.430 409.450 26.690 ;
        RECT 411.430 26.990 411.690 27.250 ;
        RECT 417.030 26.990 417.290 27.250 ;
        RECT 415.350 26.430 415.610 26.690 ;
        RECT 420.390 26.990 420.650 27.250 ;
        RECT 421.510 26.990 421.770 27.250 ;
        RECT 418.150 26.430 418.410 26.690 ;
        RECT 423.190 26.990 423.450 27.250 ;
        RECT 424.870 26.990 425.130 27.250 ;
        RECT 422.070 26.430 422.330 26.690 ;
        RECT 438.870 26.990 439.130 27.250 ;
        RECT 457.910 28.110 458.170 28.370 ;
        RECT 456.230 26.990 456.490 27.250 ;
        RECT 454.550 25.870 454.810 26.130 ;
        RECT 456.230 25.870 456.490 26.130 ;
        RECT 459.030 26.990 459.290 27.250 ;
        RECT 170.810 22.410 171.070 23.190 ;
        RECT 173.050 22.410 173.310 23.190 ;
        RECT 175.290 22.410 175.550 23.190 ;
        RECT 177.530 22.410 177.790 23.190 ;
        RECT 180.890 22.410 181.150 23.190 ;
        RECT 183.130 22.410 183.390 23.190 ;
        RECT 185.370 22.410 185.630 23.190 ;
        RECT 187.610 22.410 187.870 23.190 ;
        RECT 335.270 24.190 335.530 24.450 ;
        RECT 334.150 23.630 334.410 23.890 ;
        RECT 334.150 22.510 334.410 22.770 ;
        RECT 337.510 22.510 337.770 22.770 ;
        RECT 343.670 24.190 343.930 24.450 ;
        RECT 344.230 23.070 344.490 23.330 ;
        RECT 346.470 23.070 346.730 23.330 ;
        RECT 347.590 23.070 347.850 23.330 ;
        RECT 348.150 23.070 348.410 23.330 ;
        RECT 349.270 23.070 349.530 23.330 ;
        RECT 350.950 21.950 351.210 22.210 ;
        RECT 385.670 23.070 385.930 23.330 ;
        RECT 386.230 21.950 386.490 22.210 ;
        RECT 386.790 23.070 387.050 23.330 ;
        RECT 387.350 21.950 387.610 22.210 ;
        RECT 390.150 23.070 390.410 23.330 ;
        RECT 387.910 21.950 388.170 22.210 ;
        RECT 390.710 21.950 390.970 22.210 ;
        RECT 419.830 23.070 420.090 23.330 ;
        RECT 418.710 21.950 418.970 22.210 ;
        RECT 422.070 23.070 422.330 23.330 ;
        RECT 427.110 23.630 427.370 23.890 ;
        RECT 423.750 21.950 424.010 22.210 ;
        RECT 429.350 21.950 429.610 22.210 ;
        RECT 432.150 21.950 432.410 22.210 ;
        RECT 434.950 21.950 435.210 22.210 ;
        RECT 436.630 22.510 436.890 22.770 ;
        RECT 438.870 24.190 439.130 24.450 ;
        RECT 439.430 21.950 439.690 22.210 ;
        RECT 440.550 23.070 440.810 23.330 ;
        RECT 442.230 21.950 442.490 22.210 ;
        RECT 446.150 21.950 446.410 22.210 ;
        RECT 457.350 23.070 457.610 23.330 ;
        RECT 459.590 23.070 459.850 23.330 ;
        RECT 302.790 19.150 303.050 19.410 ;
        RECT 297.750 18.030 298.010 18.290 ;
        RECT 313.990 19.150 314.250 19.410 ;
        RECT 316.790 19.150 317.050 19.410 ;
        RECT 323.510 19.150 323.770 19.410 ;
        RECT 324.070 19.150 324.330 19.410 ;
        RECT 325.190 19.150 325.450 19.410 ;
        RECT 326.310 19.150 326.570 19.410 ;
        RECT 365.510 20.270 365.770 20.530 ;
        RECT 367.190 19.710 367.450 19.970 ;
        RECT 369.430 19.150 369.690 19.410 ;
        RECT 368.870 18.030 369.130 18.290 ;
        RECT 382.310 19.150 382.570 19.410 ;
        RECT 382.870 19.150 383.130 19.410 ;
        RECT 385.110 19.710 385.370 19.970 ;
        RECT 383.990 19.150 384.250 19.410 ;
        RECT 383.430 18.590 383.690 18.850 ;
        RECT 389.590 19.150 389.850 19.410 ;
        RECT 391.830 19.150 392.090 19.410 ;
        RECT 404.710 20.270 404.970 20.530 ;
        RECT 407.510 20.270 407.770 20.530 ;
        RECT 415.350 19.150 415.610 19.410 ;
        RECT 416.470 20.270 416.730 20.530 ;
        RECT 417.030 18.030 417.290 18.290 ;
        RECT 425.990 18.590 426.250 18.850 ;
        RECT 427.110 20.270 427.370 20.530 ;
        RECT 429.910 20.270 430.170 20.530 ;
        RECT 434.950 20.270 435.210 20.530 ;
        RECT 427.670 18.590 427.930 18.850 ;
        RECT 431.590 18.590 431.850 18.850 ;
        RECT 432.710 19.710 432.970 19.970 ;
        RECT 434.390 19.150 434.650 19.410 ;
        RECT 437.190 19.710 437.450 19.970 ;
        RECT 435.510 19.150 435.770 19.410 ;
        RECT 438.870 19.150 439.130 19.410 ;
        RECT 460.150 20.270 460.410 20.530 ;
        RECT 457.350 19.150 457.610 19.410 ;
        RECT 298.870 15.790 299.130 16.050 ;
        RECT 310.630 15.230 310.890 15.490 ;
        RECT 312.870 15.230 313.130 15.490 ;
        RECT 320.150 14.670 320.410 14.930 ;
        RECT 326.310 15.790 326.570 16.050 ;
        RECT 320.710 14.110 320.970 14.370 ;
        RECT 321.270 14.110 321.530 14.370 ;
        RECT 325.750 14.110 326.010 14.370 ;
        RECT 326.870 14.670 327.130 14.930 ;
        RECT 341.430 15.230 341.690 15.490 ;
        RECT 343.110 15.230 343.370 15.490 ;
        RECT 344.230 15.230 344.490 15.490 ;
        RECT 343.110 14.110 343.370 14.370 ;
        RECT 363.270 15.230 363.530 15.490 ;
        RECT 366.630 15.230 366.890 15.490 ;
        RECT 377.830 14.110 378.090 14.370 ;
        RECT 381.750 14.110 382.010 14.370 ;
        RECT 391.270 14.110 391.530 14.370 ;
        RECT 396.310 15.230 396.570 15.490 ;
        RECT 401.910 15.790 402.170 16.050 ;
        RECT 400.230 15.230 400.490 15.490 ;
        RECT 399.110 14.670 399.370 14.930 ;
        RECT 397.430 14.110 397.690 14.370 ;
        RECT 401.350 14.110 401.610 14.370 ;
        RECT 404.150 15.230 404.410 15.490 ;
        RECT 401.910 14.110 402.170 14.370 ;
        RECT 406.950 15.230 407.210 15.490 ;
        RECT 419.830 14.110 420.090 14.370 ;
        RECT 423.750 15.230 424.010 15.490 ;
        RECT 422.630 14.110 422.890 14.370 ;
        RECT 426.550 14.110 426.810 14.370 ;
        RECT 428.230 14.110 428.490 14.370 ;
        RECT 435.510 15.790 435.770 16.050 ;
        RECT 429.910 14.110 430.170 14.370 ;
        RECT 434.950 14.670 435.210 14.930 ;
        RECT 436.070 15.230 436.330 15.490 ;
        RECT 437.750 14.670 438.010 14.930 ;
        RECT 442.230 14.670 442.490 14.930 ;
        RECT 446.150 14.110 446.410 14.370 ;
        RECT 457.350 15.230 457.610 15.490 ;
        RECT 459.590 15.230 459.850 15.490 ;
        RECT 183.965 10.365 184.745 10.625 ;
        RECT 181.465 5.970 182.245 6.230 ;
        RECT 179.725 4.110 179.985 4.890 ;
        RECT 171.465 2.870 172.245 3.130 ;
        RECT 175.965 2.870 176.745 3.130 ;
        RECT 173.260 1.070 174.040 1.330 ;
        RECT 175.965 1.070 176.745 1.330 ;
        RECT 173.260 -1.330 174.040 -1.070 ;
        RECT 181.965 2.870 182.745 3.130 ;
        RECT 180.685 1.070 181.465 1.330 ;
        RECT 185.465 5.975 186.245 6.235 ;
        RECT 230.320 9.565 231.100 9.825 ;
        RECT 234.350 9.565 235.130 9.825 ;
        RECT 235.920 9.780 236.180 10.560 ;
        RECT 306.150 11.870 306.410 12.130 ;
        RECT 307.270 10.750 307.530 11.010 ;
        RECT 308.390 11.310 308.650 11.570 ;
        RECT 310.070 10.190 310.330 10.450 ;
        RECT 313.990 11.310 314.250 11.570 ;
        RECT 312.310 10.750 312.570 11.010 ;
        RECT 323.510 11.870 323.770 12.130 ;
        RECT 321.270 11.310 321.530 11.570 ;
        RECT 325.190 12.430 325.450 12.690 ;
        RECT 325.750 11.310 326.010 11.570 ;
        RECT 326.310 11.310 326.570 11.570 ;
        RECT 327.430 11.870 327.690 12.130 ;
        RECT 346.470 11.310 346.730 11.570 ;
        RECT 341.430 10.190 341.690 10.450 ;
        RECT 357.110 11.310 357.370 11.570 ;
        RECT 359.350 11.310 359.610 11.570 ;
        RECT 367.190 11.870 367.450 12.130 ;
        RECT 368.870 11.870 369.130 12.130 ;
        RECT 370.550 11.870 370.810 12.130 ;
        RECT 371.670 11.310 371.930 11.570 ;
        RECT 383.990 10.750 384.250 11.010 ;
        RECT 386.230 11.310 386.490 11.570 ;
        RECT 388.470 12.430 388.730 12.690 ;
        RECT 389.590 11.310 389.850 11.570 ;
        RECT 392.390 12.430 392.650 12.690 ;
        RECT 391.830 11.310 392.090 11.570 ;
        RECT 393.510 11.310 393.770 11.570 ;
        RECT 404.150 12.430 404.410 12.690 ;
        RECT 403.590 11.870 403.850 12.130 ;
        RECT 405.830 12.430 406.090 12.690 ;
        RECT 407.510 11.310 407.770 11.570 ;
        RECT 409.750 10.750 410.010 11.010 ;
        RECT 426.550 12.430 426.810 12.690 ;
        RECT 432.710 12.430 432.970 12.690 ;
        RECT 434.390 11.870 434.650 12.130 ;
        RECT 435.510 11.310 435.770 11.570 ;
        RECT 438.870 11.310 439.130 11.570 ;
        RECT 437.190 10.190 437.450 10.450 ;
        RECT 232.355 9.175 233.135 9.435 ;
        RECT 230.320 5.205 231.100 5.465 ;
        RECT 232.315 5.010 233.095 5.270 ;
        RECT 234.350 5.205 235.130 5.465 ;
        RECT 235.920 5.420 236.180 6.200 ;
        RECT 298.310 7.390 298.570 7.650 ;
        RECT 299.430 6.830 299.690 7.090 ;
        RECT 302.230 7.390 302.490 7.650 ;
        RECT 303.910 6.830 304.170 7.090 ;
        RECT 305.590 7.390 305.850 7.650 ;
        RECT 308.390 7.390 308.650 7.650 ;
        RECT 310.070 6.830 310.330 7.090 ;
        RECT 311.190 8.510 311.450 8.770 ;
        RECT 316.790 7.390 317.050 7.650 ;
        RECT 312.870 6.270 313.130 6.530 ;
        RECT 318.470 7.390 318.730 7.650 ;
        RECT 319.590 7.390 319.850 7.650 ;
        RECT 321.830 7.390 322.090 7.650 ;
        RECT 323.510 7.390 323.770 7.650 ;
        RECT 322.390 6.830 322.650 7.090 ;
        RECT 317.910 6.270 318.170 6.530 ;
        RECT 329.670 7.950 329.930 8.210 ;
        RECT 331.910 6.830 332.170 7.090 ;
        RECT 327.430 6.270 327.690 6.530 ;
        RECT 340.310 7.950 340.570 8.210 ;
        RECT 339.190 6.830 339.450 7.090 ;
        RECT 344.230 8.510 344.490 8.770 ;
        RECT 344.790 6.830 345.050 7.090 ;
        RECT 345.910 6.830 346.170 7.090 ;
        RECT 368.310 7.390 368.570 7.650 ;
        RECT 371.110 7.390 371.370 7.650 ;
        RECT 382.870 6.830 383.130 7.090 ;
        RECT 391.830 7.950 392.090 8.210 ;
        RECT 386.790 6.270 387.050 6.530 ;
        RECT 391.270 6.270 391.530 6.530 ;
        RECT 392.390 6.830 392.650 7.090 ;
        RECT 403.590 7.950 403.850 8.210 ;
        RECT 396.310 6.270 396.570 6.530 ;
        RECT 401.350 7.390 401.610 7.650 ;
        RECT 401.910 7.390 402.170 7.650 ;
        RECT 403.030 6.270 403.290 6.530 ;
        RECT 404.150 7.390 404.410 7.650 ;
        RECT 406.950 7.390 407.210 7.650 ;
        RECT 409.190 7.390 409.450 7.650 ;
        RECT 407.510 6.830 407.770 7.090 ;
        RECT 411.430 7.390 411.690 7.650 ;
        RECT 423.190 6.830 423.450 7.090 ;
        RECT 427.110 6.270 427.370 6.530 ;
        RECT 434.390 7.390 434.650 7.650 ;
        RECT 436.630 6.830 436.890 7.090 ;
        RECT 437.750 6.830 438.010 7.090 ;
        RECT 435.510 6.270 435.770 6.530 ;
        RECT 439.430 7.390 439.690 7.650 ;
        RECT 442.230 7.390 442.490 7.650 ;
        RECT 447.830 7.390 448.090 7.650 ;
        RECT 287.260 4.870 287.520 5.130 ;
        RECT 287.820 4.870 288.080 5.130 ;
        RECT 288.380 4.870 288.640 5.130 ;
        RECT 230.320 3.975 231.100 4.235 ;
        RECT 232.355 4.170 233.135 4.430 ;
        RECT 234.350 3.975 235.130 4.235 ;
        RECT 287.260 4.310 287.520 4.570 ;
        RECT 287.820 4.310 288.080 4.570 ;
        RECT 288.380 4.310 288.640 4.570 ;
        RECT 298.310 4.590 298.570 4.850 ;
        RECT 223.390 2.870 223.650 3.130 ;
        RECT 223.950 2.870 224.210 3.130 ;
        RECT 235.920 3.240 236.180 4.020 ;
        RECT 303.910 4.590 304.170 4.850 ;
        RECT 301.670 2.910 301.930 3.170 ;
        RECT 306.150 4.030 306.410 4.290 ;
        RECT 311.190 4.030 311.450 4.290 ;
        RECT 321.830 4.590 322.090 4.850 ;
        RECT 312.310 3.470 312.570 3.730 ;
        RECT 317.910 4.030 318.170 4.290 ;
        RECT 319.030 2.910 319.290 3.170 ;
        RECT 321.270 2.910 321.530 3.170 ;
        RECT 324.630 2.910 324.890 3.170 ;
        RECT 326.870 4.590 327.130 4.850 ;
        RECT 329.670 4.590 329.930 4.850 ;
        RECT 330.790 3.470 331.050 3.730 ;
        RECT 343.670 3.470 343.930 3.730 ;
        RECT 346.470 3.470 346.730 3.730 ;
        RECT 348.710 3.470 348.970 3.730 ;
        RECT 350.950 2.910 351.210 3.170 ;
        RECT 348.150 2.350 348.410 2.610 ;
        RECT 355.990 3.470 356.250 3.730 ;
        RECT 358.790 3.470 359.050 3.730 ;
        RECT 369.990 4.590 370.250 4.850 ;
        RECT 373.910 2.350 374.170 2.610 ;
        RECT 388.470 4.030 388.730 4.290 ;
        RECT 386.790 3.470 387.050 3.730 ;
        RECT 397.990 4.590 398.250 4.850 ;
        RECT 400.230 4.030 400.490 4.290 ;
        RECT 392.390 3.470 392.650 3.730 ;
        RECT 394.630 3.470 394.890 3.730 ;
        RECT 391.830 2.910 392.090 3.170 ;
        RECT 397.990 3.470 398.250 3.730 ;
        RECT 406.390 3.470 406.650 3.730 ;
        RECT 426.550 4.590 426.810 4.850 ;
        RECT 428.230 3.470 428.490 3.730 ;
        RECT 432.150 4.030 432.410 4.290 ;
        RECT 431.590 3.470 431.850 3.730 ;
        RECT 429.350 2.910 429.610 3.170 ;
        RECT 435.510 4.030 435.770 4.290 ;
        RECT 434.390 3.470 434.650 3.730 ;
        RECT 433.270 2.910 433.530 3.170 ;
        RECT 436.630 4.590 436.890 4.850 ;
        RECT 439.990 3.470 440.250 3.730 ;
        RECT 437.190 2.350 437.450 2.610 ;
        RECT 454.550 3.470 454.810 3.730 ;
        RECT 456.790 2.910 457.050 3.170 ;
        RECT 175.965 -1.330 176.745 -1.070 ;
        RECT 171.465 -3.130 172.245 -2.870 ;
        RECT 175.965 -3.130 176.745 -2.870 ;
        RECT 232.355 0.005 233.135 0.265 ;
        RECT 180.685 -1.330 181.465 -1.070 ;
        RECT 181.965 -3.130 182.745 -2.870 ;
        RECT 179.725 -4.890 179.985 -4.110 ;
        RECT 181.465 -6.230 182.245 -5.970 ;
        RECT 185.465 -6.230 186.245 -5.970 ;
        RECT 230.320 -0.385 231.100 -0.125 ;
        RECT 234.350 -0.385 235.130 -0.125 ;
        RECT 235.920 -1.120 236.180 -0.340 ;
        RECT 304.470 0.110 304.730 0.370 ;
        RECT 305.030 -0.450 305.290 -0.190 ;
        RECT 305.590 -1.570 305.850 -1.310 ;
        RECT 317.350 -0.450 317.610 -0.190 ;
        RECT 319.590 -0.450 319.850 -0.190 ;
        RECT 320.150 -1.570 320.410 -1.310 ;
        RECT 320.710 -1.570 320.970 -1.310 ;
        RECT 323.510 -1.570 323.770 -1.310 ;
        RECT 329.110 -0.450 329.370 -0.190 ;
        RECT 331.350 -0.450 331.610 -0.190 ;
        RECT 346.470 0.670 346.730 0.930 ;
        RECT 343.670 -1.570 343.930 -1.310 ;
        RECT 347.590 0.670 347.850 0.930 ;
        RECT 349.270 -0.450 349.530 -0.190 ;
        RECT 349.830 -1.570 350.090 -1.310 ;
        RECT 350.390 -1.570 350.650 -1.310 ;
        RECT 350.950 -0.450 351.210 -0.190 ;
        RECT 353.750 -1.570 354.010 -1.310 ;
        RECT 362.150 0.110 362.410 0.370 ;
        RECT 356.550 -1.010 356.810 -0.750 ;
        RECT 358.230 -1.010 358.490 -0.750 ;
        RECT 361.590 -1.010 361.850 -0.750 ;
        RECT 363.830 -0.450 364.090 -0.190 ;
        RECT 363.270 -1.010 363.530 -0.750 ;
        RECT 370.550 0.110 370.810 0.370 ;
        RECT 368.310 -0.450 368.570 -0.190 ;
        RECT 369.430 -1.010 369.690 -0.750 ;
        RECT 371.110 -1.010 371.370 -0.750 ;
        RECT 382.310 -0.450 382.570 -0.190 ;
        RECT 382.870 -1.570 383.130 -1.310 ;
        RECT 384.550 -1.570 384.810 -1.310 ;
        RECT 387.350 -1.010 387.610 -0.750 ;
        RECT 392.950 0.110 393.210 0.370 ;
        RECT 390.150 -1.570 390.410 -1.310 ;
        RECT 396.870 -0.450 397.130 -0.190 ;
        RECT 395.750 -1.010 396.010 -0.750 ;
        RECT 401.350 0.110 401.610 0.370 ;
        RECT 399.670 -0.450 399.930 -0.190 ;
        RECT 402.470 -1.010 402.730 -0.750 ;
        RECT 404.710 -1.570 404.970 -1.310 ;
        RECT 408.630 -0.450 408.890 -0.190 ;
        RECT 409.190 -1.570 409.450 -1.310 ;
        RECT 412.550 -1.010 412.810 -0.750 ;
        RECT 411.990 -1.570 412.250 -1.310 ;
        RECT 415.350 -1.570 415.610 -1.310 ;
        RECT 418.150 -1.010 418.410 -0.750 ;
        RECT 434.950 0.670 435.210 0.930 ;
        RECT 436.630 0.110 436.890 0.370 ;
        RECT 438.310 0.110 438.570 0.370 ;
        RECT 436.070 -1.010 436.330 -0.750 ;
        RECT 439.430 0.670 439.690 0.930 ;
        RECT 441.110 0.670 441.370 0.930 ;
        RECT 442.230 -0.450 442.490 -0.190 ;
        RECT 446.150 -1.010 446.410 -0.750 ;
        RECT 457.350 -0.450 457.610 -0.190 ;
        RECT 459.590 -0.450 459.850 -0.190 ;
        RECT 223.510 -3.130 223.770 -2.870 ;
        RECT 224.070 -3.130 224.330 -2.870 ;
        RECT 298.310 -4.370 298.570 -4.110 ;
        RECT 287.260 -5.210 287.520 -4.950 ;
        RECT 287.820 -5.210 288.080 -4.950 ;
        RECT 288.380 -5.210 288.640 -4.950 ;
        RECT 230.550 -5.805 231.330 -5.545 ;
        RECT 234.065 -5.805 234.845 -5.545 ;
        RECT 300.550 -4.370 300.810 -4.110 ;
        RECT 230.335 -7.375 230.595 -6.595 ;
        RECT 233.850 -7.375 234.110 -6.595 ;
        RECT 229.955 -9.390 230.215 -8.610 ;
        RECT 233.470 -9.390 233.730 -8.610 ;
        RECT 287.260 -5.770 287.520 -5.510 ;
        RECT 287.820 -5.770 288.080 -5.510 ;
        RECT 288.380 -5.770 288.640 -5.510 ;
        RECT 316.230 -3.250 316.490 -2.990 ;
        RECT 311.750 -4.370 312.010 -4.110 ;
        RECT 317.350 -3.250 317.610 -2.990 ;
        RECT 318.470 -3.250 318.730 -2.990 ;
        RECT 319.030 -3.810 319.290 -3.550 ;
        RECT 320.710 -4.370 320.970 -4.110 ;
        RECT 321.830 -3.810 322.090 -3.550 ;
        RECT 324.630 -3.810 324.890 -3.550 ;
        RECT 325.750 -3.250 326.010 -2.990 ;
        RECT 328.550 -3.250 328.810 -2.990 ;
        RECT 324.070 -4.370 324.330 -4.110 ;
        RECT 326.310 -4.370 326.570 -4.110 ;
        RECT 321.270 -4.930 321.530 -4.670 ;
        RECT 330.790 -4.930 331.050 -4.670 ;
        RECT 336.950 -3.810 337.210 -3.550 ;
        RECT 338.630 -4.370 338.890 -4.110 ;
        RECT 345.910 -4.370 346.170 -4.110 ;
        RECT 346.470 -3.810 346.730 -3.550 ;
        RECT 347.030 -4.370 347.290 -4.110 ;
        RECT 349.270 -3.250 349.530 -2.990 ;
        RECT 350.950 -4.370 351.210 -4.110 ;
        RECT 351.510 -3.810 351.770 -3.550 ;
        RECT 362.150 -3.250 362.410 -2.990 ;
        RECT 361.590 -4.370 361.850 -4.110 ;
        RECT 362.710 -4.370 362.970 -4.110 ;
        RECT 363.830 -5.490 364.090 -5.230 ;
        RECT 369.430 -3.810 369.690 -3.550 ;
        RECT 369.990 -3.250 370.250 -2.990 ;
        RECT 370.550 -5.490 370.810 -5.230 ;
        RECT 388.470 -3.810 388.730 -3.550 ;
        RECT 383.990 -4.370 384.250 -4.110 ;
        RECT 386.230 -4.370 386.490 -4.110 ;
        RECT 394.630 -4.370 394.890 -4.110 ;
        RECT 382.310 -5.490 382.570 -5.230 ;
        RECT 383.990 -5.490 384.250 -5.230 ;
        RECT 397.430 -4.930 397.690 -4.670 ;
        RECT 407.510 -3.810 407.770 -3.550 ;
        RECT 400.790 -4.370 401.050 -4.110 ;
        RECT 403.590 -4.370 403.850 -4.110 ;
        RECT 406.390 -4.370 406.650 -4.110 ;
        RECT 409.190 -3.250 409.450 -2.990 ;
        RECT 435.510 -3.250 435.770 -2.990 ;
        RECT 418.150 -3.810 418.410 -3.550 ;
        RECT 411.990 -4.370 412.250 -4.110 ;
        RECT 419.830 -4.370 420.090 -4.110 ;
        RECT 401.910 -5.490 402.170 -5.230 ;
        RECT 423.750 -4.370 424.010 -4.110 ;
        RECT 424.870 -4.370 425.130 -4.110 ;
        RECT 417.590 -5.490 417.850 -5.230 ;
        RECT 437.190 -4.370 437.450 -4.110 ;
        RECT 440.550 -4.370 440.810 -4.110 ;
        RECT 457.350 -4.370 457.610 -4.110 ;
        RECT 460.150 -4.370 460.410 -4.110 ;
        RECT 298.870 -7.170 299.130 -6.910 ;
        RECT 308.390 -8.290 308.650 -8.030 ;
        RECT 321.830 -8.290 322.090 -8.030 ;
        RECT 323.510 -8.290 323.770 -8.030 ;
        RECT 335.270 -8.850 335.530 -8.590 ;
        RECT 339.190 -7.170 339.450 -6.910 ;
        RECT 362.150 -8.850 362.410 -8.590 ;
        RECT 364.950 -8.290 365.210 -8.030 ;
        RECT 367.750 -8.290 368.010 -8.030 ;
        RECT 363.270 -8.850 363.530 -8.590 ;
        RECT 375.590 -8.290 375.850 -8.030 ;
        RECT 362.710 -9.410 362.970 -9.150 ;
        RECT 382.310 -8.850 382.570 -8.590 ;
        RECT 385.110 -8.290 385.370 -8.030 ;
        RECT 387.910 -8.290 388.170 -8.030 ;
        RECT 389.590 -7.730 389.850 -7.470 ;
        RECT 391.830 -8.290 392.090 -8.030 ;
        RECT 377.270 -9.410 377.530 -9.150 ;
        RECT 391.270 -8.850 391.530 -8.590 ;
        RECT 403.590 -7.730 403.850 -7.470 ;
        RECT 399.670 -8.290 399.930 -8.030 ;
        RECT 401.350 -8.290 401.610 -8.030 ;
        RECT 404.150 -8.850 404.410 -8.590 ;
        RECT 406.950 -8.290 407.210 -8.030 ;
        RECT 396.310 -9.410 396.570 -9.150 ;
        RECT 408.630 -8.850 408.890 -8.590 ;
        RECT 406.390 -9.410 406.650 -9.150 ;
        RECT 411.990 -8.290 412.250 -8.030 ;
        RECT 414.230 -7.730 414.490 -7.470 ;
        RECT 419.830 -7.730 420.090 -7.470 ;
        RECT 422.630 -8.290 422.890 -8.030 ;
        RECT 424.310 -8.290 424.570 -8.030 ;
        RECT 427.110 -8.290 427.370 -8.030 ;
        RECT 428.790 -8.850 429.050 -8.590 ;
        RECT 438.310 -7.730 438.570 -7.470 ;
        RECT 430.470 -9.410 430.730 -9.150 ;
        RECT 442.790 -8.290 443.050 -8.030 ;
        RECT 445.030 -8.290 445.290 -8.030 ;
        RECT 456.790 -9.410 457.050 -9.150 ;
        RECT 460.710 -9.410 460.970 -9.150 ;
        RECT 183.965 -10.625 184.745 -10.365 ;
        RECT 230.335 -11.405 230.595 -10.625 ;
        RECT 233.850 -11.405 234.110 -10.625 ;
        RECT 298.870 -13.330 299.130 -13.070 ;
        RECT 308.390 -12.210 308.650 -11.950 ;
        RECT 347.590 -11.090 347.850 -10.830 ;
        RECT 349.270 -12.210 349.530 -11.950 ;
        RECT 352.070 -11.650 352.330 -11.390 ;
        RECT 353.190 -12.210 353.450 -11.950 ;
        RECT 363.270 -11.090 363.530 -10.830 ;
        RECT 360.470 -12.770 360.730 -12.510 ;
        RECT 366.630 -11.090 366.890 -10.830 ;
        RECT 368.310 -12.210 368.570 -11.950 ;
        RECT 371.110 -11.650 371.370 -11.390 ;
        RECT 372.230 -12.210 372.490 -11.950 ;
        RECT 379.510 -12.210 379.770 -11.950 ;
        RECT 396.310 -11.650 396.570 -11.390 ;
        RECT 383.430 -12.210 383.690 -11.950 ;
        RECT 384.550 -12.210 384.810 -11.950 ;
        RECT 398.550 -12.210 398.810 -11.950 ;
        RECT 381.190 -12.770 381.450 -12.510 ;
        RECT 403.590 -11.650 403.850 -11.390 ;
        RECT 400.790 -12.210 401.050 -11.950 ;
        RECT 383.990 -13.330 384.250 -13.070 ;
        RECT 392.390 -12.770 392.650 -12.510 ;
        RECT 411.990 -11.650 412.250 -11.390 ;
        RECT 417.030 -11.650 417.290 -11.390 ;
        RECT 412.550 -12.770 412.810 -12.510 ;
        RECT 410.870 -13.330 411.130 -13.070 ;
        RECT 419.270 -12.770 419.530 -12.510 ;
        RECT 425.990 -11.090 426.250 -10.830 ;
        RECT 429.350 -11.090 429.610 -10.830 ;
        RECT 441.110 -12.210 441.370 -11.950 ;
        RECT 446.150 -11.090 446.410 -10.830 ;
        RECT 443.350 -12.210 443.610 -11.950 ;
        RECT 299.990 -15.010 300.250 -14.750 ;
        RECT 300.550 -16.690 300.810 -16.430 ;
        RECT 302.790 -16.130 303.050 -15.870 ;
        RECT 306.150 -15.010 306.410 -14.750 ;
        RECT 303.910 -16.690 304.170 -16.430 ;
        RECT 305.590 -15.570 305.850 -15.310 ;
        RECT 308.390 -15.570 308.650 -15.310 ;
        RECT 323.510 -16.130 323.770 -15.870 ;
        RECT 321.830 -17.250 322.090 -16.990 ;
        RECT 324.630 -16.690 324.890 -16.430 ;
        RECT 326.870 -17.250 327.130 -16.990 ;
        RECT 329.110 -16.130 329.370 -15.870 ;
        RECT 331.910 -16.130 332.170 -15.870 ;
        RECT 330.790 -17.250 331.050 -16.990 ;
        RECT 335.270 -16.130 335.530 -15.870 ;
        RECT 350.390 -15.570 350.650 -15.310 ;
        RECT 346.470 -17.250 346.730 -16.990 ;
        RECT 352.070 -16.130 352.330 -15.870 ;
        RECT 359.910 -15.570 360.170 -15.310 ;
        RECT 353.190 -17.250 353.450 -16.990 ;
        RECT 359.350 -17.250 359.610 -16.990 ;
        RECT 360.470 -16.690 360.730 -16.430 ;
        RECT 362.710 -15.010 362.970 -14.750 ;
        RECT 363.270 -16.130 363.530 -15.870 ;
        RECT 363.830 -16.130 364.090 -15.870 ;
        RECT 370.550 -16.690 370.810 -16.430 ;
        RECT 371.670 -15.570 371.930 -15.310 ;
        RECT 372.230 -16.130 372.490 -15.870 ;
        RECT 376.150 -15.010 376.410 -14.750 ;
        RECT 377.830 -15.010 378.090 -14.750 ;
        RECT 378.950 -16.690 379.210 -16.430 ;
        RECT 380.630 -16.130 380.890 -15.870 ;
        RECT 382.310 -16.690 382.570 -16.430 ;
        RECT 390.710 -16.690 390.970 -16.430 ;
        RECT 391.830 -17.250 392.090 -16.990 ;
        RECT 417.030 -15.010 417.290 -14.750 ;
        RECT 392.390 -17.250 392.650 -16.990 ;
        RECT 392.950 -16.130 393.210 -15.870 ;
        RECT 397.990 -15.570 398.250 -15.310 ;
        RECT 401.910 -16.130 402.170 -15.870 ;
        RECT 404.150 -16.130 404.410 -15.870 ;
        RECT 415.350 -16.130 415.610 -15.870 ;
        RECT 403.030 -16.690 403.290 -16.430 ;
        RECT 404.710 -16.690 404.970 -16.430 ;
        RECT 408.630 -16.690 408.890 -16.430 ;
        RECT 414.790 -16.690 415.050 -16.430 ;
        RECT 420.950 -16.130 421.210 -15.870 ;
        RECT 422.630 -16.130 422.890 -15.870 ;
        RECT 448.390 -16.130 448.650 -15.870 ;
        RECT 298.310 -20.610 298.570 -20.350 ;
        RECT 300.550 -20.050 300.810 -19.790 ;
        RECT 304.470 -20.050 304.730 -19.790 ;
        RECT 306.710 -20.050 306.970 -19.790 ;
        RECT 319.030 -18.930 319.290 -18.670 ;
        RECT 323.510 -18.930 323.770 -18.670 ;
        RECT 321.830 -19.490 322.090 -19.230 ;
        RECT 322.950 -20.050 323.210 -19.790 ;
        RECT 324.630 -20.050 324.890 -19.790 ;
        RECT 325.190 -20.050 325.450 -19.790 ;
        RECT 327.990 -20.610 328.250 -20.350 ;
        RECT 372.790 -19.490 373.050 -19.230 ;
        RECT 365.510 -20.050 365.770 -19.790 ;
        RECT 368.310 -20.050 368.570 -19.790 ;
        RECT 371.670 -20.050 371.930 -19.790 ;
        RECT 372.230 -20.610 372.490 -20.350 ;
        RECT 376.710 -19.490 376.970 -19.230 ;
        RECT 376.150 -20.610 376.410 -20.350 ;
        RECT 382.870 -19.490 383.130 -19.230 ;
        RECT 385.110 -20.050 385.370 -19.790 ;
        RECT 385.670 -20.610 385.930 -20.350 ;
        RECT 391.830 -20.050 392.090 -19.790 ;
        RECT 394.630 -20.050 394.890 -19.790 ;
        RECT 390.710 -20.610 390.970 -20.350 ;
        RECT 403.590 -19.490 403.850 -19.230 ;
        RECT 390.150 -21.170 390.410 -20.910 ;
        RECT 395.750 -21.170 396.010 -20.910 ;
        RECT 401.910 -20.610 402.170 -20.350 ;
        RECT 402.470 -21.170 402.730 -20.910 ;
        RECT 410.310 -21.170 410.570 -20.910 ;
        RECT 410.870 -20.610 411.130 -20.350 ;
        RECT 411.990 -20.050 412.250 -19.790 ;
        RECT 418.710 -20.050 418.970 -19.790 ;
        RECT 419.830 -20.050 420.090 -19.790 ;
        RECT 418.150 -20.610 418.410 -20.350 ;
        RECT 425.430 -19.490 425.690 -19.230 ;
        RECT 412.550 -21.170 412.810 -20.910 ;
        RECT 421.510 -21.170 421.770 -20.910 ;
        RECT 432.710 -18.930 432.970 -18.670 ;
        RECT 431.590 -20.050 431.850 -19.790 ;
        RECT 433.830 -20.050 434.090 -19.790 ;
        RECT 436.630 -20.050 436.890 -19.790 ;
        RECT 449.510 -18.930 449.770 -18.670 ;
        RECT 452.310 -18.930 452.570 -18.670 ;
        RECT 455.110 -18.930 455.370 -18.670 ;
        RECT 456.230 -20.050 456.490 -19.790 ;
        RECT 458.470 -19.490 458.730 -19.230 ;
        RECT 459.590 -20.050 459.850 -19.790 ;
        RECT 170.810 -23.190 171.070 -22.410 ;
        RECT 173.050 -23.190 173.310 -22.410 ;
        RECT 175.290 -23.190 175.550 -22.410 ;
        RECT 177.530 -23.190 177.790 -22.410 ;
        RECT 180.890 -23.190 181.150 -22.410 ;
        RECT 183.130 -23.190 183.390 -22.410 ;
        RECT 185.370 -23.190 185.630 -22.410 ;
        RECT 187.610 -23.190 187.870 -22.410 ;
        RECT 171.930 -25.190 172.190 -24.410 ;
        RECT 176.410 -25.190 176.670 -24.410 ;
        RECT 182.010 -25.190 182.270 -24.410 ;
        RECT 186.490 -25.190 186.750 -24.410 ;
        RECT 174.170 -27.190 174.430 -26.410 ;
        RECT 184.250 -27.190 184.510 -26.410 ;
        RECT 178.650 -29.580 178.910 -28.800 ;
        RECT 179.770 -29.580 180.030 -28.800 ;
        RECT 298.870 -23.410 299.130 -23.150 ;
        RECT 308.390 -23.970 308.650 -23.710 ;
        RECT 312.310 -24.530 312.570 -24.270 ;
        RECT 313.990 -25.090 314.250 -24.830 ;
        RECT 319.590 -23.410 319.850 -23.150 ;
        RECT 320.150 -25.090 320.410 -24.830 ;
        RECT 321.270 -23.410 321.530 -23.150 ;
        RECT 343.670 -25.090 343.930 -24.830 ;
        RECT 345.350 -25.090 345.610 -24.830 ;
        RECT 351.510 -24.530 351.770 -24.270 ;
        RECT 353.190 -24.530 353.450 -24.270 ;
        RECT 356.550 -23.970 356.810 -23.710 ;
        RECT 359.350 -23.410 359.610 -23.150 ;
        RECT 358.230 -23.970 358.490 -23.710 ;
        RECT 353.750 -25.090 354.010 -24.830 ;
        RECT 358.790 -25.090 359.050 -24.830 ;
        RECT 359.910 -25.090 360.170 -24.830 ;
        RECT 361.590 -23.970 361.850 -23.710 ;
        RECT 363.270 -23.970 363.530 -23.710 ;
        RECT 362.710 -24.530 362.970 -24.270 ;
        RECT 372.790 -23.970 373.050 -23.710 ;
        RECT 374.470 -23.970 374.730 -23.710 ;
        RECT 380.630 -23.970 380.890 -23.710 ;
        RECT 367.190 -24.530 367.450 -24.270 ;
        RECT 365.510 -25.090 365.770 -24.830 ;
        RECT 385.670 -25.090 385.930 -24.830 ;
        RECT 386.790 -25.090 387.050 -24.830 ;
        RECT 387.350 -25.090 387.610 -24.830 ;
        RECT 387.910 -25.090 388.170 -24.830 ;
        RECT 390.710 -23.970 390.970 -23.710 ;
        RECT 392.390 -25.090 392.650 -24.830 ;
        RECT 399.670 -23.970 399.930 -23.710 ;
        RECT 402.470 -23.970 402.730 -23.710 ;
        RECT 418.150 -23.410 418.410 -23.150 ;
        RECT 415.350 -25.090 415.610 -24.830 ;
        RECT 418.710 -23.970 418.970 -23.710 ;
        RECT 424.310 -23.410 424.570 -23.150 ;
        RECT 420.390 -23.970 420.650 -23.710 ;
        RECT 421.510 -23.970 421.770 -23.710 ;
        RECT 420.390 -25.090 420.650 -24.830 ;
        RECT 435.510 -23.410 435.770 -23.150 ;
        RECT 437.190 -23.410 437.450 -23.150 ;
        RECT 438.310 -24.530 438.570 -24.270 ;
        RECT 439.990 -24.530 440.250 -24.270 ;
        RECT 445.590 -24.530 445.850 -24.270 ;
        RECT 443.910 -25.090 444.170 -24.830 ;
        RECT 447.270 -23.970 447.530 -23.710 ;
        RECT 459.030 -22.850 459.290 -22.590 ;
        RECT 299.430 -27.890 299.690 -27.630 ;
        RECT 301.670 -27.890 301.930 -27.630 ;
        RECT 313.430 -26.770 313.690 -26.510 ;
        RECT 319.590 -26.770 319.850 -26.510 ;
        RECT 316.790 -27.890 317.050 -27.630 ;
        RECT 319.030 -27.330 319.290 -27.070 ;
        RECT 318.470 -27.890 318.730 -27.630 ;
        RECT 322.390 -26.770 322.650 -26.510 ;
        RECT 321.270 -27.890 321.530 -27.630 ;
        RECT 324.070 -27.890 324.330 -27.630 ;
        RECT 325.190 -27.330 325.450 -27.070 ;
        RECT 349.830 -26.770 350.090 -26.510 ;
        RECT 349.270 -27.330 349.530 -27.070 ;
        RECT 354.310 -26.770 354.570 -26.510 ;
        RECT 352.070 -29.010 352.330 -28.750 ;
        RECT 353.750 -27.890 354.010 -27.630 ;
        RECT 355.430 -27.890 355.690 -27.630 ;
        RECT 354.870 -28.450 355.130 -28.190 ;
        RECT 364.950 -27.330 365.210 -27.070 ;
        RECT 366.630 -27.890 366.890 -27.630 ;
        RECT 376.150 -27.330 376.410 -27.070 ;
        RECT 377.830 -26.770 378.090 -26.510 ;
        RECT 383.990 -28.450 384.250 -28.190 ;
        RECT 386.230 -27.890 386.490 -27.630 ;
        RECT 395.750 -26.770 396.010 -26.510 ;
        RECT 395.190 -27.330 395.450 -27.070 ;
        RECT 396.870 -27.890 397.130 -27.630 ;
        RECT 400.230 -27.890 400.490 -27.630 ;
        RECT 401.910 -26.770 402.170 -26.510 ;
        RECT 402.470 -27.890 402.730 -27.630 ;
        RECT 403.590 -27.890 403.850 -27.630 ;
        RECT 405.270 -27.890 405.530 -27.630 ;
        RECT 405.830 -27.330 406.090 -27.070 ;
        RECT 418.150 -26.770 418.410 -26.510 ;
        RECT 423.190 -26.770 423.450 -26.510 ;
        RECT 422.070 -27.330 422.330 -27.070 ;
        RECT 424.310 -27.330 424.570 -27.070 ;
        RECT 419.830 -28.450 420.090 -28.190 ;
        RECT 425.990 -27.330 426.250 -27.070 ;
        RECT 427.670 -27.330 427.930 -27.070 ;
        RECT 424.870 -29.010 425.130 -28.750 ;
        RECT 432.710 -27.330 432.970 -27.070 ;
        RECT 437.190 -26.770 437.450 -26.510 ;
        RECT 431.590 -27.890 431.850 -27.630 ;
        RECT 434.390 -28.450 434.650 -28.190 ;
        RECT 435.510 -27.890 435.770 -27.630 ;
        RECT 438.870 -27.890 439.130 -27.630 ;
        RECT 457.350 -26.770 457.610 -26.510 ;
        RECT 460.150 -28.450 460.410 -28.190 ;
        RECT 313.430 -30.690 313.690 -30.430 ;
        RECT 309.510 -31.810 309.770 -31.550 ;
        RECT 312.870 -31.810 313.130 -31.550 ;
        RECT 317.350 -30.690 317.610 -30.430 ;
        RECT 319.030 -30.690 319.290 -30.430 ;
        RECT 315.110 -31.810 315.370 -31.550 ;
        RECT 301.670 -32.370 301.930 -32.110 ;
        RECT 317.910 -32.930 318.170 -32.670 ;
        RECT 320.710 -31.250 320.970 -30.990 ;
        RECT 321.270 -32.930 321.530 -32.670 ;
        RECT 322.390 -32.370 322.650 -32.110 ;
        RECT 327.990 -31.810 328.250 -31.550 ;
        RECT 331.350 -31.810 331.610 -31.550 ;
        RECT 346.470 -31.810 346.730 -31.550 ;
        RECT 342.550 -32.930 342.810 -32.670 ;
        RECT 371.110 -30.690 371.370 -30.430 ;
        RECT 372.230 -32.370 372.490 -32.110 ;
        RECT 373.910 -32.370 374.170 -32.110 ;
        RECT 369.430 -32.930 369.690 -32.670 ;
        RECT 386.790 -30.690 387.050 -30.430 ;
        RECT 389.590 -31.810 389.850 -31.550 ;
        RECT 390.150 -32.370 390.410 -32.110 ;
        RECT 385.110 -32.930 385.370 -32.670 ;
        RECT 401.910 -31.810 402.170 -31.550 ;
        RECT 403.590 -31.810 403.850 -31.550 ;
        RECT 405.270 -32.370 405.530 -32.110 ;
        RECT 403.030 -32.930 403.290 -32.670 ;
        RECT 421.510 -31.810 421.770 -31.550 ;
        RECT 423.190 -31.810 423.450 -31.550 ;
        RECT 423.750 -31.810 424.010 -31.550 ;
        RECT 422.070 -32.370 422.330 -32.110 ;
        RECT 425.430 -31.810 425.690 -31.550 ;
        RECT 427.670 -32.930 427.930 -32.670 ;
        RECT 428.230 -32.930 428.490 -32.670 ;
        RECT 428.790 -31.810 429.050 -31.550 ;
        RECT 430.470 -31.250 430.730 -30.990 ;
        RECT 431.030 -32.930 431.290 -32.670 ;
        RECT 436.070 -31.810 436.330 -31.550 ;
        RECT 437.190 -31.250 437.450 -30.990 ;
        RECT 432.150 -32.370 432.410 -32.110 ;
        RECT 438.310 -31.250 438.570 -30.990 ;
        RECT 439.430 -32.370 439.690 -32.110 ;
        RECT 439.990 -31.810 440.250 -31.550 ;
        RECT 440.550 -32.370 440.810 -32.110 ;
        RECT 442.230 -31.810 442.490 -31.550 ;
        RECT 445.030 -31.810 445.290 -31.550 ;
        RECT 456.790 -32.370 457.050 -32.110 ;
        RECT 460.710 -32.930 460.970 -32.670 ;
        RECT 168.175 -35.090 168.435 -34.310 ;
        RECT 174.175 -35.090 174.435 -34.310 ;
        RECT 178.105 -35.155 178.365 -34.375 ;
        RECT 180.245 -35.155 180.505 -34.375 ;
        RECT 186.675 -35.090 186.935 -34.310 ;
        RECT 300.550 -35.730 300.810 -35.470 ;
        RECT 303.910 -35.730 304.170 -35.470 ;
        RECT 315.110 -34.610 315.370 -34.350 ;
        RECT 322.390 -34.610 322.650 -34.350 ;
        RECT 319.030 -35.730 319.290 -35.470 ;
        RECT 320.150 -35.730 320.410 -35.470 ;
        RECT 321.830 -35.730 322.090 -35.470 ;
        RECT 323.510 -35.730 323.770 -35.470 ;
        RECT 325.190 -36.290 325.450 -36.030 ;
        RECT 330.790 -34.610 331.050 -34.350 ;
        RECT 331.910 -35.730 332.170 -35.470 ;
        RECT 337.510 -34.610 337.770 -34.350 ;
        RECT 336.950 -36.850 337.210 -36.590 ;
        RECT 338.630 -36.850 338.890 -36.590 ;
        RECT 344.790 -35.730 345.050 -35.470 ;
        RECT 347.030 -35.730 347.290 -35.470 ;
        RECT 349.270 -36.290 349.530 -36.030 ;
        RECT 349.830 -35.170 350.090 -34.910 ;
        RECT 352.070 -35.730 352.330 -35.470 ;
        RECT 353.190 -34.610 353.450 -34.350 ;
        RECT 354.310 -35.730 354.570 -35.470 ;
        RECT 352.630 -36.290 352.890 -36.030 ;
        RECT 355.430 -35.730 355.690 -35.470 ;
        RECT 357.670 -34.610 357.930 -34.350 ;
        RECT 358.790 -35.730 359.050 -35.470 ;
        RECT 359.350 -35.730 359.610 -35.470 ;
        RECT 358.230 -36.290 358.490 -36.030 ;
        RECT 361.030 -36.850 361.290 -36.590 ;
        RECT 363.270 -35.170 363.530 -34.910 ;
        RECT 364.950 -35.170 365.210 -34.910 ;
        RECT 362.710 -36.850 362.970 -36.590 ;
        RECT 366.630 -35.730 366.890 -35.470 ;
        RECT 369.990 -35.170 370.250 -34.910 ;
        RECT 368.870 -35.730 369.130 -35.470 ;
        RECT 371.670 -34.610 371.930 -34.350 ;
        RECT 372.790 -35.730 373.050 -35.470 ;
        RECT 377.830 -34.610 378.090 -34.350 ;
        RECT 380.070 -35.170 380.330 -34.910 ;
        RECT 386.790 -34.610 387.050 -34.350 ;
        RECT 382.310 -35.730 382.570 -35.470 ;
        RECT 389.590 -34.610 389.850 -34.350 ;
        RECT 383.990 -36.290 384.250 -36.030 ;
        RECT 386.230 -36.290 386.490 -36.030 ;
        RECT 387.910 -36.850 388.170 -36.590 ;
        RECT 391.270 -35.730 391.530 -35.470 ;
        RECT 418.710 -34.610 418.970 -34.350 ;
        RECT 444.470 -34.610 444.730 -34.350 ;
        RECT 432.710 -35.170 432.970 -34.910 ;
        RECT 437.190 -35.730 437.450 -35.470 ;
        RECT 439.430 -35.730 439.690 -35.470 ;
        RECT 433.270 -36.290 433.530 -36.030 ;
        RECT 445.030 -35.170 445.290 -34.910 ;
        RECT 448.390 -34.610 448.650 -34.350 ;
        RECT 446.710 -35.730 446.970 -35.470 ;
        RECT 450.070 -34.610 450.330 -34.350 ;
        RECT 451.190 -35.730 451.450 -35.470 ;
        RECT 455.110 -34.610 455.370 -34.350 ;
        RECT 460.150 -34.610 460.410 -34.350 ;
        RECT 457.350 -35.730 457.610 -35.470 ;
        RECT 310.630 -39.650 310.890 -39.390 ;
        RECT 305.590 -40.770 305.850 -40.510 ;
        RECT 317.910 -38.530 318.170 -38.270 ;
        RECT 312.870 -39.090 313.130 -38.830 ;
        RECT 319.590 -38.530 319.850 -38.270 ;
        RECT 312.310 -40.770 312.570 -40.510 ;
        RECT 320.710 -39.090 320.970 -38.830 ;
        RECT 322.950 -39.090 323.210 -38.830 ;
        RECT 327.990 -39.650 328.250 -39.390 ;
        RECT 326.310 -40.210 326.570 -39.950 ;
        RECT 330.230 -39.650 330.490 -39.390 ;
        RECT 332.470 -39.650 332.730 -39.390 ;
        RECT 347.590 -38.530 347.850 -38.270 ;
        RECT 344.790 -40.770 345.050 -40.510 ;
        RECT 357.110 -38.530 357.370 -38.270 ;
        RECT 356.550 -40.210 356.810 -39.950 ;
        RECT 369.430 -39.650 369.690 -39.390 ;
        RECT 372.230 -39.650 372.490 -39.390 ;
        RECT 387.910 -38.530 388.170 -38.270 ;
        RECT 383.990 -40.770 384.250 -40.510 ;
        RECT 390.710 -39.090 390.970 -38.830 ;
        RECT 400.790 -39.650 401.050 -39.390 ;
        RECT 403.030 -39.650 403.290 -39.390 ;
        RECT 418.150 -38.530 418.410 -38.270 ;
        RECT 414.790 -40.770 415.050 -40.510 ;
        RECT 435.510 -38.530 435.770 -38.270 ;
        RECT 431.590 -39.650 431.850 -39.390 ;
        RECT 436.070 -39.090 436.330 -38.830 ;
        RECT 427.110 -40.770 427.370 -40.510 ;
        RECT 437.190 -39.650 437.450 -39.390 ;
        RECT 438.870 -40.210 439.130 -39.950 ;
        RECT 439.430 -39.090 439.690 -38.830 ;
        RECT 442.790 -39.650 443.050 -39.390 ;
        RECT 457.350 -39.090 457.610 -38.830 ;
        RECT 447.830 -40.770 448.090 -40.510 ;
        RECT 298.870 -44.690 299.130 -44.430 ;
        RECT 308.950 -43.570 309.210 -43.310 ;
        RECT 312.310 -43.570 312.570 -43.310 ;
        RECT 315.110 -43.570 315.370 -43.310 ;
        RECT 317.350 -43.570 317.610 -43.310 ;
        RECT 319.030 -43.570 319.290 -43.310 ;
        RECT 331.910 -42.450 332.170 -42.190 ;
        RECT 334.710 -43.570 334.970 -43.310 ;
        RECT 338.630 -44.130 338.890 -43.870 ;
        RECT 340.310 -43.570 340.570 -43.310 ;
        RECT 343.110 -42.450 343.370 -42.190 ;
        RECT 342.550 -43.010 342.810 -42.750 ;
        RECT 344.230 -43.010 344.490 -42.750 ;
        RECT 344.790 -43.570 345.050 -43.310 ;
        RECT 348.710 -43.570 348.970 -43.310 ;
        RECT 347.030 -44.130 347.290 -43.870 ;
        RECT 349.830 -43.010 350.090 -42.750 ;
        RECT 354.870 -42.450 355.130 -42.190 ;
        RECT 357.670 -42.450 357.930 -42.190 ;
        RECT 369.990 -43.570 370.250 -43.310 ;
        RECT 372.790 -43.570 373.050 -43.310 ;
        RECT 376.710 -43.010 376.970 -42.750 ;
        RECT 381.190 -43.010 381.450 -42.750 ;
        RECT 380.070 -43.570 380.330 -43.310 ;
        RECT 376.150 -44.690 376.410 -44.430 ;
        RECT 382.310 -42.450 382.570 -42.190 ;
        RECT 386.230 -42.450 386.490 -42.190 ;
        RECT 397.430 -43.570 397.690 -43.310 ;
        RECT 402.470 -42.450 402.730 -42.190 ;
        RECT 400.790 -43.570 401.050 -43.310 ;
        RECT 406.390 -43.010 406.650 -42.750 ;
        RECT 409.190 -42.450 409.450 -42.190 ;
        RECT 406.950 -44.690 407.210 -44.430 ;
        RECT 417.590 -42.450 417.850 -42.190 ;
        RECT 418.710 -43.010 418.970 -42.750 ;
        RECT 421.510 -43.570 421.770 -43.310 ;
        RECT 419.270 -44.690 419.530 -44.430 ;
        RECT 423.750 -43.570 424.010 -43.310 ;
        RECT 436.070 -42.450 436.330 -42.190 ;
        RECT 438.870 -42.450 439.130 -42.190 ;
        RECT 441.670 -42.450 441.930 -42.190 ;
        RECT 441.110 -43.570 441.370 -43.310 ;
        RECT 443.910 -42.450 444.170 -42.190 ;
        RECT 450.070 -42.450 450.330 -42.190 ;
        RECT 458.470 -42.450 458.730 -42.190 ;
        RECT 455.110 -43.010 455.370 -42.750 ;
        RECT 454.550 -44.130 454.810 -43.870 ;
        RECT 300.550 -46.930 300.810 -46.670 ;
        RECT 312.310 -47.490 312.570 -47.230 ;
        RECT 319.030 -47.490 319.290 -47.230 ;
        RECT 333.590 -46.930 333.850 -46.670 ;
        RECT 322.390 -48.610 322.650 -48.350 ;
        RECT 335.830 -47.490 336.090 -47.230 ;
        RECT 340.870 -46.930 341.130 -46.670 ;
        RECT 352.630 -46.930 352.890 -46.670 ;
        RECT 354.870 -47.490 355.130 -47.230 ;
        RECT 359.910 -46.930 360.170 -46.670 ;
        RECT 376.150 -47.490 376.410 -47.230 ;
        RECT 389.030 -46.930 389.290 -46.670 ;
        RECT 381.750 -48.050 382.010 -47.790 ;
        RECT 389.590 -47.490 389.850 -47.230 ;
        RECT 392.950 -47.490 393.210 -47.230 ;
        RECT 398.550 -46.930 398.810 -46.670 ;
        RECT 411.990 -47.490 412.250 -47.230 ;
        RECT 417.030 -46.930 417.290 -46.670 ;
        RECT 432.150 -47.490 432.410 -47.230 ;
        RECT 436.070 -46.930 436.330 -46.670 ;
        RECT 453.990 -46.930 454.250 -46.670 ;
        RECT 456.790 -48.050 457.050 -47.790 ;
        RECT 458.470 -48.050 458.730 -47.790 ;
        RECT 144.920 -63.520 145.180 -63.260 ;
        RECT 143.665 -64.045 143.925 -63.785 ;
        RECT 144.920 -66.880 145.180 -66.620 ;
        RECT 143.665 -67.405 143.925 -67.145 ;
        RECT 144.920 -70.240 145.180 -69.980 ;
        RECT 143.665 -70.765 143.925 -70.505 ;
        RECT 144.920 -73.600 145.180 -73.340 ;
        RECT 143.665 -74.125 143.925 -73.865 ;
        RECT 144.920 -76.960 145.180 -76.700 ;
        RECT 143.665 -77.485 143.925 -77.225 ;
        RECT -484.685 -79.595 -483.905 -79.335 ;
        RECT 144.920 -80.320 145.180 -80.060 ;
        RECT 143.665 -80.845 143.925 -80.585 ;
        RECT -497.465 -83.695 -495.645 -83.435 ;
        RECT -492.270 -84.715 -491.490 -84.455 ;
        RECT -486.885 -83.105 -486.625 -81.285 ;
        RECT 144.920 -83.680 145.180 -83.420 ;
        RECT 143.665 -84.205 143.925 -83.945 ;
        RECT -490.555 -86.505 -490.295 -85.725 ;
        RECT 144.920 -87.040 145.180 -86.780 ;
        RECT 143.665 -87.565 143.925 -87.305 ;
        RECT 144.920 -90.400 145.180 -90.140 ;
        RECT 143.665 -90.925 143.925 -90.665 ;
        RECT 144.920 -93.760 145.180 -93.500 ;
        RECT 143.665 -94.285 143.925 -94.025 ;
        RECT -493.415 -95.770 -492.635 -95.510 ;
        RECT -489.385 -95.770 -488.605 -95.510 ;
        RECT -491.760 -97.985 -491.500 -97.205 ;
        RECT 143.665 -97.645 143.925 -97.385 ;
      LAYER Metal2 ;
        RECT -492.150 105.625 -491.110 106.425 ;
        RECT -491.830 97.075 -491.430 105.625 ;
        RECT 466.700 105.525 469.200 106.525 ;
        RECT -189.405 96.915 -189.005 98.115 ;
        RECT 120.925 97.715 121.925 97.765 ;
        RECT 120.925 97.315 143.995 97.715 ;
        RECT 120.925 97.265 121.925 97.315 ;
        RECT -493.475 95.450 -488.545 95.830 ;
        RECT -490.615 90.515 -490.235 95.450 ;
        RECT -490.615 90.135 -490.225 90.515 ;
        RECT -332.765 90.195 -332.365 91.395 ;
        RECT -490.615 84.775 -490.235 90.135 ;
        RECT -404.445 86.835 -404.045 88.035 ;
        RECT -492.330 84.395 -490.235 84.775 ;
        RECT -497.595 83.365 -495.515 83.765 ;
        RECT -440.285 83.475 -439.885 84.675 ;
        RECT -486.955 81.155 -486.555 83.235 ;
        RECT -458.205 80.115 -457.805 81.315 ;
        RECT -484.745 79.275 -482.495 79.655 ;
        RECT -483.245 56.095 -482.495 79.275 ;
        RECT -467.165 76.755 -466.765 77.955 ;
        RECT -471.645 73.395 -471.245 74.595 ;
        RECT -473.885 70.035 -473.485 71.235 ;
        RECT -477.745 66.285 -475.785 66.685 ;
        RECT -475.005 66.675 -474.605 67.875 ;
        RECT -477.745 56.255 -477.465 66.285 ;
        RECT -477.185 56.695 -476.905 66.285 ;
        RECT -476.625 56.255 -476.345 65.695 ;
        RECT -476.065 56.695 -475.785 66.285 ;
        RECT -475.505 56.255 -475.225 65.695 ;
        RECT -474.945 56.535 -474.665 66.675 ;
        RECT -474.385 56.255 -474.105 65.695 ;
        RECT -473.825 56.535 -473.545 70.035 ;
        RECT -472.765 66.675 -472.365 67.875 ;
        RECT -473.265 56.255 -472.985 65.695 ;
        RECT -472.705 56.535 -472.425 66.675 ;
        RECT -472.145 56.255 -471.865 65.695 ;
        RECT -471.585 56.535 -471.305 73.395 ;
        RECT -469.405 70.035 -469.005 71.235 ;
        RECT -470.525 66.675 -470.125 67.875 ;
        RECT -471.025 56.255 -470.745 65.695 ;
        RECT -470.465 56.535 -470.185 66.675 ;
        RECT -469.905 56.255 -469.625 65.695 ;
        RECT -469.345 56.535 -469.065 70.035 ;
        RECT -468.285 66.675 -467.885 67.875 ;
        RECT -468.785 56.255 -468.505 65.695 ;
        RECT -468.225 56.535 -467.945 66.675 ;
        RECT -467.665 56.255 -467.385 65.695 ;
        RECT -467.105 56.535 -466.825 76.755 ;
        RECT -462.685 73.395 -462.285 74.595 ;
        RECT -464.925 70.035 -464.525 71.235 ;
        RECT -466.045 66.675 -465.645 67.875 ;
        RECT -466.545 56.255 -466.265 65.695 ;
        RECT -465.985 56.535 -465.705 66.675 ;
        RECT -465.425 56.255 -465.145 65.695 ;
        RECT -464.865 56.535 -464.585 70.035 ;
        RECT -463.805 66.675 -463.405 67.875 ;
        RECT -464.305 56.255 -464.025 65.695 ;
        RECT -463.745 56.535 -463.465 66.675 ;
        RECT -463.185 56.255 -462.905 65.695 ;
        RECT -462.625 56.535 -462.345 73.395 ;
        RECT -460.445 70.035 -460.045 71.235 ;
        RECT -461.565 66.675 -461.165 67.875 ;
        RECT -462.065 56.255 -461.785 65.695 ;
        RECT -461.505 56.535 -461.225 66.675 ;
        RECT -460.945 56.255 -460.665 65.695 ;
        RECT -460.385 56.535 -460.105 70.035 ;
        RECT -459.325 66.675 -458.925 67.875 ;
        RECT -459.825 56.255 -459.545 65.695 ;
        RECT -459.265 56.535 -458.985 66.675 ;
        RECT -458.705 56.255 -458.425 65.695 ;
        RECT -458.145 56.535 -457.865 80.115 ;
        RECT -449.245 76.755 -448.845 77.955 ;
        RECT -453.725 73.395 -453.325 74.595 ;
        RECT -455.965 70.035 -455.565 71.235 ;
        RECT -457.085 66.675 -456.685 67.875 ;
        RECT -457.585 56.255 -457.305 65.695 ;
        RECT -457.025 56.535 -456.745 66.675 ;
        RECT -456.465 56.255 -456.185 65.695 ;
        RECT -455.905 56.535 -455.625 70.035 ;
        RECT -454.845 66.675 -454.445 67.875 ;
        RECT -455.345 56.255 -455.065 65.695 ;
        RECT -454.785 56.535 -454.505 66.675 ;
        RECT -454.225 56.255 -453.945 65.695 ;
        RECT -453.665 56.535 -453.385 73.395 ;
        RECT -451.485 70.035 -451.085 71.235 ;
        RECT -452.605 66.675 -452.205 67.875 ;
        RECT -453.105 56.255 -452.825 65.695 ;
        RECT -452.545 56.535 -452.265 66.675 ;
        RECT -451.985 56.255 -451.705 65.695 ;
        RECT -451.425 56.535 -451.145 70.035 ;
        RECT -450.365 66.675 -449.965 67.875 ;
        RECT -450.865 56.255 -450.585 65.695 ;
        RECT -450.305 56.535 -450.025 66.675 ;
        RECT -449.745 56.255 -449.465 65.695 ;
        RECT -449.185 56.535 -448.905 76.755 ;
        RECT -444.765 73.395 -444.365 74.595 ;
        RECT -447.005 70.035 -446.605 71.235 ;
        RECT -448.125 66.675 -447.725 67.875 ;
        RECT -448.625 56.255 -448.345 65.695 ;
        RECT -448.065 56.535 -447.785 66.675 ;
        RECT -447.505 56.255 -447.225 65.695 ;
        RECT -446.945 56.535 -446.665 70.035 ;
        RECT -445.885 66.675 -445.485 67.875 ;
        RECT -446.385 56.255 -446.105 65.695 ;
        RECT -445.825 56.535 -445.545 66.675 ;
        RECT -445.265 56.255 -444.985 65.695 ;
        RECT -444.705 56.535 -444.425 73.395 ;
        RECT -442.525 70.035 -442.125 71.235 ;
        RECT -443.645 66.675 -443.245 67.875 ;
        RECT -444.145 56.255 -443.865 65.695 ;
        RECT -443.585 56.535 -443.305 66.675 ;
        RECT -443.025 56.255 -442.745 65.695 ;
        RECT -442.465 56.535 -442.185 70.035 ;
        RECT -441.405 66.675 -441.005 67.875 ;
        RECT -441.905 56.255 -441.625 65.695 ;
        RECT -441.345 56.535 -441.065 66.675 ;
        RECT -440.785 56.255 -440.505 65.695 ;
        RECT -440.225 56.535 -439.945 83.475 ;
        RECT -422.365 80.115 -421.965 81.315 ;
        RECT -431.325 76.755 -430.925 77.955 ;
        RECT -435.805 73.395 -435.405 74.595 ;
        RECT -438.045 70.035 -437.645 71.235 ;
        RECT -439.165 66.675 -438.765 67.875 ;
        RECT -439.665 56.255 -439.385 65.695 ;
        RECT -439.105 56.535 -438.825 66.675 ;
        RECT -438.545 56.255 -438.265 65.695 ;
        RECT -437.985 56.535 -437.705 70.035 ;
        RECT -436.925 66.675 -436.525 67.875 ;
        RECT -437.425 56.255 -437.145 65.695 ;
        RECT -436.865 56.535 -436.585 66.675 ;
        RECT -436.305 56.255 -436.025 65.695 ;
        RECT -435.745 56.535 -435.465 73.395 ;
        RECT -433.565 70.035 -433.165 71.235 ;
        RECT -434.685 66.675 -434.285 67.875 ;
        RECT -435.185 56.255 -434.905 65.695 ;
        RECT -434.625 56.535 -434.345 66.675 ;
        RECT -434.065 56.255 -433.785 65.695 ;
        RECT -433.505 56.535 -433.225 70.035 ;
        RECT -432.445 66.675 -432.045 67.875 ;
        RECT -432.945 56.255 -432.665 65.695 ;
        RECT -432.385 56.535 -432.105 66.675 ;
        RECT -431.825 56.255 -431.545 65.695 ;
        RECT -431.265 56.535 -430.985 76.755 ;
        RECT -426.845 73.395 -426.445 74.595 ;
        RECT -429.085 70.035 -428.685 71.235 ;
        RECT -430.205 66.675 -429.805 67.875 ;
        RECT -430.705 56.255 -430.425 65.695 ;
        RECT -430.145 56.535 -429.865 66.675 ;
        RECT -429.585 56.255 -429.305 65.695 ;
        RECT -429.025 56.535 -428.745 70.035 ;
        RECT -427.965 66.675 -427.565 67.875 ;
        RECT -428.465 56.255 -428.185 65.695 ;
        RECT -427.905 56.535 -427.625 66.675 ;
        RECT -427.345 56.255 -427.065 65.695 ;
        RECT -426.785 56.535 -426.505 73.395 ;
        RECT -424.605 70.035 -424.205 71.235 ;
        RECT -425.725 66.675 -425.325 67.875 ;
        RECT -426.225 56.255 -425.945 65.695 ;
        RECT -425.665 56.535 -425.385 66.675 ;
        RECT -425.105 56.255 -424.825 65.695 ;
        RECT -424.545 56.535 -424.265 70.035 ;
        RECT -423.485 66.675 -423.085 67.875 ;
        RECT -423.985 56.255 -423.705 65.695 ;
        RECT -423.425 56.535 -423.145 66.675 ;
        RECT -422.865 56.255 -422.585 65.695 ;
        RECT -422.305 56.535 -422.025 80.115 ;
        RECT -413.405 76.755 -413.005 77.955 ;
        RECT -417.885 73.395 -417.485 74.595 ;
        RECT -420.125 70.035 -419.725 71.235 ;
        RECT -421.245 66.675 -420.845 67.875 ;
        RECT -421.745 56.255 -421.465 65.695 ;
        RECT -421.185 56.535 -420.905 66.675 ;
        RECT -420.625 56.255 -420.345 65.695 ;
        RECT -420.065 56.535 -419.785 70.035 ;
        RECT -419.005 66.675 -418.605 67.875 ;
        RECT -419.505 56.255 -419.225 65.695 ;
        RECT -418.945 56.535 -418.665 66.675 ;
        RECT -418.385 56.255 -418.105 65.695 ;
        RECT -417.825 56.535 -417.545 73.395 ;
        RECT -415.645 70.035 -415.245 71.235 ;
        RECT -416.765 66.675 -416.365 67.875 ;
        RECT -417.265 56.255 -416.985 65.695 ;
        RECT -416.705 56.535 -416.425 66.675 ;
        RECT -416.145 56.255 -415.865 65.695 ;
        RECT -415.585 56.535 -415.305 70.035 ;
        RECT -414.525 66.675 -414.125 67.875 ;
        RECT -415.025 56.255 -414.745 65.695 ;
        RECT -414.465 56.535 -414.185 66.675 ;
        RECT -413.905 56.255 -413.625 65.695 ;
        RECT -413.345 56.535 -413.065 76.755 ;
        RECT -408.925 73.395 -408.525 74.595 ;
        RECT -411.165 70.035 -410.765 71.235 ;
        RECT -412.285 66.675 -411.885 67.875 ;
        RECT -412.785 56.255 -412.505 65.695 ;
        RECT -412.225 56.535 -411.945 66.675 ;
        RECT -411.665 56.255 -411.385 65.695 ;
        RECT -411.105 56.535 -410.825 70.035 ;
        RECT -410.045 66.675 -409.645 67.875 ;
        RECT -410.545 56.255 -410.265 65.695 ;
        RECT -409.985 56.535 -409.705 66.675 ;
        RECT -409.425 56.255 -409.145 65.695 ;
        RECT -408.865 56.535 -408.585 73.395 ;
        RECT -406.685 70.035 -406.285 71.235 ;
        RECT -407.805 66.675 -407.405 67.875 ;
        RECT -408.305 56.255 -408.025 65.695 ;
        RECT -407.745 56.535 -407.465 66.675 ;
        RECT -407.185 56.255 -406.905 65.695 ;
        RECT -406.625 56.535 -406.345 70.035 ;
        RECT -405.565 66.675 -405.165 67.875 ;
        RECT -406.065 56.255 -405.785 65.695 ;
        RECT -405.505 56.535 -405.225 66.675 ;
        RECT -404.945 56.255 -404.665 65.695 ;
        RECT -404.385 56.535 -404.105 86.835 ;
        RECT -368.605 83.475 -368.205 84.675 ;
        RECT -386.525 80.115 -386.125 81.315 ;
        RECT -395.485 76.755 -395.085 77.955 ;
        RECT -399.965 73.395 -399.565 74.595 ;
        RECT -402.205 70.035 -401.805 71.235 ;
        RECT -403.325 66.675 -402.925 67.875 ;
        RECT -403.825 56.255 -403.545 65.695 ;
        RECT -403.265 56.535 -402.985 66.675 ;
        RECT -402.705 56.255 -402.425 65.695 ;
        RECT -402.145 56.535 -401.865 70.035 ;
        RECT -401.085 66.675 -400.685 67.875 ;
        RECT -401.585 56.255 -401.305 65.695 ;
        RECT -401.025 56.535 -400.745 66.675 ;
        RECT -400.465 56.255 -400.185 65.695 ;
        RECT -399.905 56.535 -399.625 73.395 ;
        RECT -397.725 70.035 -397.325 71.235 ;
        RECT -398.845 66.675 -398.445 67.875 ;
        RECT -399.345 56.255 -399.065 65.695 ;
        RECT -398.785 56.535 -398.505 66.675 ;
        RECT -398.225 56.255 -397.945 65.695 ;
        RECT -397.665 56.535 -397.385 70.035 ;
        RECT -396.605 66.675 -396.205 67.875 ;
        RECT -397.105 56.255 -396.825 65.695 ;
        RECT -396.545 56.535 -396.265 66.675 ;
        RECT -395.985 56.255 -395.705 65.695 ;
        RECT -395.425 56.535 -395.145 76.755 ;
        RECT -391.005 73.395 -390.605 74.595 ;
        RECT -393.245 70.035 -392.845 71.235 ;
        RECT -394.365 66.675 -393.965 67.875 ;
        RECT -394.865 56.255 -394.585 65.695 ;
        RECT -394.305 56.535 -394.025 66.675 ;
        RECT -393.745 56.255 -393.465 65.695 ;
        RECT -393.185 56.535 -392.905 70.035 ;
        RECT -392.125 66.675 -391.725 67.875 ;
        RECT -392.625 56.255 -392.345 65.695 ;
        RECT -392.065 56.535 -391.785 66.675 ;
        RECT -391.505 56.255 -391.225 65.695 ;
        RECT -390.945 56.535 -390.665 73.395 ;
        RECT -388.765 70.035 -388.365 71.235 ;
        RECT -389.885 66.675 -389.485 67.875 ;
        RECT -390.385 56.255 -390.105 65.695 ;
        RECT -389.825 56.535 -389.545 66.675 ;
        RECT -389.265 56.255 -388.985 65.695 ;
        RECT -388.705 56.535 -388.425 70.035 ;
        RECT -387.645 66.675 -387.245 67.875 ;
        RECT -388.145 56.255 -387.865 65.695 ;
        RECT -387.585 56.535 -387.305 66.675 ;
        RECT -387.025 56.255 -386.745 65.695 ;
        RECT -386.465 56.535 -386.185 80.115 ;
        RECT -377.565 76.755 -377.165 77.955 ;
        RECT -382.045 73.395 -381.645 74.595 ;
        RECT -384.285 70.035 -383.885 71.235 ;
        RECT -385.405 66.675 -385.005 67.875 ;
        RECT -385.905 56.255 -385.625 65.695 ;
        RECT -385.345 56.535 -385.065 66.675 ;
        RECT -384.785 56.255 -384.505 65.695 ;
        RECT -384.225 56.535 -383.945 70.035 ;
        RECT -383.165 66.675 -382.765 67.875 ;
        RECT -383.665 56.255 -383.385 65.695 ;
        RECT -383.105 56.535 -382.825 66.675 ;
        RECT -382.545 56.255 -382.265 65.695 ;
        RECT -381.985 56.535 -381.705 73.395 ;
        RECT -379.805 70.035 -379.405 71.235 ;
        RECT -380.925 66.675 -380.525 67.875 ;
        RECT -381.425 56.255 -381.145 65.695 ;
        RECT -380.865 56.535 -380.585 66.675 ;
        RECT -380.305 56.255 -380.025 65.695 ;
        RECT -379.745 56.535 -379.465 70.035 ;
        RECT -378.685 66.675 -378.285 67.875 ;
        RECT -379.185 56.255 -378.905 65.695 ;
        RECT -378.625 56.535 -378.345 66.675 ;
        RECT -378.065 56.255 -377.785 65.695 ;
        RECT -377.505 56.535 -377.225 76.755 ;
        RECT -373.085 73.395 -372.685 74.595 ;
        RECT -375.325 70.035 -374.925 71.235 ;
        RECT -376.445 66.675 -376.045 67.875 ;
        RECT -376.945 56.255 -376.665 65.695 ;
        RECT -376.385 56.535 -376.105 66.675 ;
        RECT -375.825 56.255 -375.545 65.695 ;
        RECT -375.265 56.535 -374.985 70.035 ;
        RECT -374.205 66.675 -373.805 67.875 ;
        RECT -374.705 56.255 -374.425 65.695 ;
        RECT -374.145 56.535 -373.865 66.675 ;
        RECT -373.585 56.255 -373.305 65.695 ;
        RECT -373.025 56.535 -372.745 73.395 ;
        RECT -370.845 70.035 -370.445 71.235 ;
        RECT -371.965 66.675 -371.565 67.875 ;
        RECT -372.465 56.255 -372.185 65.695 ;
        RECT -371.905 56.535 -371.625 66.675 ;
        RECT -371.345 56.255 -371.065 65.695 ;
        RECT -370.785 56.535 -370.505 70.035 ;
        RECT -369.725 66.675 -369.325 67.875 ;
        RECT -370.225 56.255 -369.945 65.695 ;
        RECT -369.665 56.535 -369.385 66.675 ;
        RECT -369.105 56.255 -368.825 65.695 ;
        RECT -368.545 56.535 -368.265 83.475 ;
        RECT -350.685 80.115 -350.285 81.315 ;
        RECT -359.645 76.755 -359.245 77.955 ;
        RECT -364.125 73.395 -363.725 74.595 ;
        RECT -366.365 70.035 -365.965 71.235 ;
        RECT -367.485 66.675 -367.085 67.875 ;
        RECT -367.985 56.255 -367.705 65.695 ;
        RECT -367.425 56.535 -367.145 66.675 ;
        RECT -366.865 56.255 -366.585 65.695 ;
        RECT -366.305 56.535 -366.025 70.035 ;
        RECT -365.245 66.675 -364.845 67.875 ;
        RECT -365.745 56.255 -365.465 65.695 ;
        RECT -365.185 56.535 -364.905 66.675 ;
        RECT -364.625 56.255 -364.345 65.695 ;
        RECT -364.065 56.535 -363.785 73.395 ;
        RECT -361.885 70.035 -361.485 71.235 ;
        RECT -363.005 66.675 -362.605 67.875 ;
        RECT -363.505 56.255 -363.225 65.695 ;
        RECT -362.945 56.535 -362.665 66.675 ;
        RECT -362.385 56.255 -362.105 65.695 ;
        RECT -361.825 56.535 -361.545 70.035 ;
        RECT -360.765 66.675 -360.365 67.875 ;
        RECT -361.265 56.255 -360.985 65.695 ;
        RECT -360.705 56.535 -360.425 66.675 ;
        RECT -360.145 56.255 -359.865 65.695 ;
        RECT -359.585 56.535 -359.305 76.755 ;
        RECT -355.165 73.395 -354.765 74.595 ;
        RECT -357.405 70.035 -357.005 71.235 ;
        RECT -358.525 66.675 -358.125 67.875 ;
        RECT -359.025 56.255 -358.745 65.695 ;
        RECT -358.465 56.535 -358.185 66.675 ;
        RECT -357.905 56.255 -357.625 65.695 ;
        RECT -357.345 56.535 -357.065 70.035 ;
        RECT -356.285 66.675 -355.885 67.875 ;
        RECT -356.785 56.255 -356.505 65.695 ;
        RECT -356.225 56.535 -355.945 66.675 ;
        RECT -355.665 56.255 -355.385 65.695 ;
        RECT -355.105 56.535 -354.825 73.395 ;
        RECT -352.925 70.035 -352.525 71.235 ;
        RECT -354.045 66.675 -353.645 67.875 ;
        RECT -354.545 56.255 -354.265 65.695 ;
        RECT -353.985 56.535 -353.705 66.675 ;
        RECT -353.425 56.255 -353.145 65.695 ;
        RECT -352.865 56.535 -352.585 70.035 ;
        RECT -351.805 66.675 -351.405 67.875 ;
        RECT -352.305 56.255 -352.025 65.695 ;
        RECT -351.745 56.535 -351.465 66.675 ;
        RECT -351.185 56.255 -350.905 65.695 ;
        RECT -350.625 56.535 -350.345 80.115 ;
        RECT -341.725 76.755 -341.325 77.955 ;
        RECT -346.205 73.395 -345.805 74.595 ;
        RECT -348.445 70.035 -348.045 71.235 ;
        RECT -349.565 66.675 -349.165 67.875 ;
        RECT -350.065 56.255 -349.785 65.695 ;
        RECT -349.505 56.535 -349.225 66.675 ;
        RECT -348.945 56.255 -348.665 65.695 ;
        RECT -348.385 56.535 -348.105 70.035 ;
        RECT -347.325 66.675 -346.925 67.875 ;
        RECT -347.825 56.255 -347.545 65.695 ;
        RECT -347.265 56.535 -346.985 66.675 ;
        RECT -346.705 56.255 -346.425 65.695 ;
        RECT -346.145 56.535 -345.865 73.395 ;
        RECT -343.965 70.035 -343.565 71.235 ;
        RECT -345.085 66.675 -344.685 67.875 ;
        RECT -345.585 56.255 -345.305 65.695 ;
        RECT -345.025 56.535 -344.745 66.675 ;
        RECT -344.465 56.255 -344.185 65.695 ;
        RECT -343.905 56.535 -343.625 70.035 ;
        RECT -342.845 66.675 -342.445 67.875 ;
        RECT -343.345 56.255 -343.065 65.695 ;
        RECT -342.785 56.535 -342.505 66.675 ;
        RECT -342.225 56.255 -341.945 65.695 ;
        RECT -341.665 56.535 -341.385 76.755 ;
        RECT -337.245 73.395 -336.845 74.595 ;
        RECT -339.485 70.035 -339.085 71.235 ;
        RECT -340.605 66.675 -340.205 67.875 ;
        RECT -341.105 56.255 -340.825 65.695 ;
        RECT -340.545 56.535 -340.265 66.675 ;
        RECT -339.985 56.255 -339.705 65.695 ;
        RECT -339.425 56.535 -339.145 70.035 ;
        RECT -338.365 66.675 -337.965 67.875 ;
        RECT -338.865 56.255 -338.585 65.695 ;
        RECT -338.305 56.535 -338.025 66.675 ;
        RECT -337.745 56.255 -337.465 65.695 ;
        RECT -337.185 56.535 -336.905 73.395 ;
        RECT -335.005 70.035 -334.605 71.235 ;
        RECT -336.125 66.675 -335.725 67.875 ;
        RECT -336.625 56.255 -336.345 65.695 ;
        RECT -336.065 56.535 -335.785 66.675 ;
        RECT -335.505 56.255 -335.225 65.695 ;
        RECT -334.945 56.535 -334.665 70.035 ;
        RECT -333.885 66.675 -333.485 67.875 ;
        RECT -334.385 56.255 -334.105 65.695 ;
        RECT -333.825 56.535 -333.545 66.675 ;
        RECT -333.265 56.255 -332.985 65.695 ;
        RECT -332.705 56.535 -332.425 90.195 ;
        RECT -261.085 86.835 -260.685 88.035 ;
        RECT -296.925 83.475 -296.525 84.675 ;
        RECT -314.845 80.115 -314.445 81.315 ;
        RECT -323.805 76.755 -323.405 77.955 ;
        RECT -328.285 73.395 -327.885 74.595 ;
        RECT -330.525 70.035 -330.125 71.235 ;
        RECT -331.645 66.675 -331.245 67.875 ;
        RECT -332.145 56.255 -331.865 65.695 ;
        RECT -331.585 56.535 -331.305 66.675 ;
        RECT -331.025 56.255 -330.745 65.695 ;
        RECT -330.465 56.535 -330.185 70.035 ;
        RECT -329.405 66.675 -329.005 67.875 ;
        RECT -329.905 56.255 -329.625 65.695 ;
        RECT -329.345 56.535 -329.065 66.675 ;
        RECT -328.785 56.255 -328.505 65.695 ;
        RECT -328.225 56.535 -327.945 73.395 ;
        RECT -326.045 70.035 -325.645 71.235 ;
        RECT -327.165 66.675 -326.765 67.875 ;
        RECT -327.665 56.255 -327.385 65.695 ;
        RECT -327.105 56.535 -326.825 66.675 ;
        RECT -326.545 56.255 -326.265 65.695 ;
        RECT -325.985 56.535 -325.705 70.035 ;
        RECT -324.925 66.675 -324.525 67.875 ;
        RECT -325.425 56.255 -325.145 65.695 ;
        RECT -324.865 56.535 -324.585 66.675 ;
        RECT -324.305 56.255 -324.025 65.695 ;
        RECT -323.745 56.535 -323.465 76.755 ;
        RECT -319.325 73.395 -318.925 74.595 ;
        RECT -321.565 70.035 -321.165 71.235 ;
        RECT -322.685 66.675 -322.285 67.875 ;
        RECT -323.185 56.255 -322.905 65.695 ;
        RECT -322.625 56.535 -322.345 66.675 ;
        RECT -322.065 56.255 -321.785 65.695 ;
        RECT -321.505 56.535 -321.225 70.035 ;
        RECT -320.445 66.675 -320.045 67.875 ;
        RECT -320.945 56.255 -320.665 65.695 ;
        RECT -320.385 56.535 -320.105 66.675 ;
        RECT -319.825 56.255 -319.545 65.695 ;
        RECT -319.265 56.535 -318.985 73.395 ;
        RECT -317.085 70.035 -316.685 71.235 ;
        RECT -318.205 66.675 -317.805 67.875 ;
        RECT -318.705 56.255 -318.425 65.695 ;
        RECT -318.145 56.535 -317.865 66.675 ;
        RECT -317.585 56.255 -317.305 65.695 ;
        RECT -317.025 56.535 -316.745 70.035 ;
        RECT -315.965 66.675 -315.565 67.875 ;
        RECT -316.465 56.255 -316.185 65.695 ;
        RECT -315.905 56.535 -315.625 66.675 ;
        RECT -315.345 56.255 -315.065 65.695 ;
        RECT -314.785 56.535 -314.505 80.115 ;
        RECT -305.885 76.755 -305.485 77.955 ;
        RECT -310.365 73.395 -309.965 74.595 ;
        RECT -312.605 70.035 -312.205 71.235 ;
        RECT -313.725 66.675 -313.325 67.875 ;
        RECT -314.225 56.255 -313.945 65.695 ;
        RECT -313.665 56.535 -313.385 66.675 ;
        RECT -313.105 56.255 -312.825 65.695 ;
        RECT -312.545 56.535 -312.265 70.035 ;
        RECT -311.485 66.675 -311.085 67.875 ;
        RECT -311.985 56.255 -311.705 65.695 ;
        RECT -311.425 56.535 -311.145 66.675 ;
        RECT -310.865 56.255 -310.585 65.695 ;
        RECT -310.305 56.535 -310.025 73.395 ;
        RECT -308.125 70.035 -307.725 71.235 ;
        RECT -309.245 66.675 -308.845 67.875 ;
        RECT -309.745 56.255 -309.465 65.695 ;
        RECT -309.185 56.535 -308.905 66.675 ;
        RECT -308.625 56.255 -308.345 65.695 ;
        RECT -308.065 56.535 -307.785 70.035 ;
        RECT -307.005 66.675 -306.605 67.875 ;
        RECT -307.505 56.255 -307.225 65.695 ;
        RECT -306.945 56.535 -306.665 66.675 ;
        RECT -306.385 56.255 -306.105 65.695 ;
        RECT -305.825 56.535 -305.545 76.755 ;
        RECT -301.405 73.395 -301.005 74.595 ;
        RECT -303.645 70.035 -303.245 71.235 ;
        RECT -304.765 66.675 -304.365 67.875 ;
        RECT -305.265 56.255 -304.985 65.695 ;
        RECT -304.705 56.535 -304.425 66.675 ;
        RECT -304.145 56.255 -303.865 65.695 ;
        RECT -303.585 56.535 -303.305 70.035 ;
        RECT -302.525 66.675 -302.125 67.875 ;
        RECT -303.025 56.255 -302.745 65.695 ;
        RECT -302.465 56.535 -302.185 66.675 ;
        RECT -301.905 56.255 -301.625 65.695 ;
        RECT -301.345 56.535 -301.065 73.395 ;
        RECT -299.165 70.035 -298.765 71.235 ;
        RECT -300.285 66.675 -299.885 67.875 ;
        RECT -300.785 56.255 -300.505 65.695 ;
        RECT -300.225 56.535 -299.945 66.675 ;
        RECT -299.665 56.255 -299.385 65.695 ;
        RECT -299.105 56.535 -298.825 70.035 ;
        RECT -298.045 66.675 -297.645 67.875 ;
        RECT -298.545 56.255 -298.265 65.695 ;
        RECT -297.985 56.535 -297.705 66.675 ;
        RECT -297.425 56.255 -297.145 65.695 ;
        RECT -296.865 56.535 -296.585 83.475 ;
        RECT -279.005 80.115 -278.605 81.315 ;
        RECT -287.965 76.755 -287.565 77.955 ;
        RECT -292.445 73.395 -292.045 74.595 ;
        RECT -294.685 70.035 -294.285 71.235 ;
        RECT -295.805 66.675 -295.405 67.875 ;
        RECT -296.305 56.255 -296.025 65.695 ;
        RECT -295.745 56.535 -295.465 66.675 ;
        RECT -295.185 56.255 -294.905 65.695 ;
        RECT -294.625 56.535 -294.345 70.035 ;
        RECT -293.565 66.675 -293.165 67.875 ;
        RECT -294.065 56.255 -293.785 65.695 ;
        RECT -293.505 56.535 -293.225 66.675 ;
        RECT -292.945 56.255 -292.665 65.695 ;
        RECT -292.385 56.535 -292.105 73.395 ;
        RECT -290.205 70.035 -289.805 71.235 ;
        RECT -291.325 66.675 -290.925 67.875 ;
        RECT -291.825 56.255 -291.545 65.695 ;
        RECT -291.265 56.535 -290.985 66.675 ;
        RECT -290.705 56.255 -290.425 65.695 ;
        RECT -290.145 56.535 -289.865 70.035 ;
        RECT -289.085 66.675 -288.685 67.875 ;
        RECT -289.585 56.255 -289.305 65.695 ;
        RECT -289.025 56.535 -288.745 66.675 ;
        RECT -288.465 56.255 -288.185 65.695 ;
        RECT -287.905 56.535 -287.625 76.755 ;
        RECT -283.485 73.395 -283.085 74.595 ;
        RECT -285.725 70.035 -285.325 71.235 ;
        RECT -286.845 66.675 -286.445 67.875 ;
        RECT -287.345 56.255 -287.065 65.695 ;
        RECT -286.785 56.535 -286.505 66.675 ;
        RECT -286.225 56.255 -285.945 65.695 ;
        RECT -285.665 56.535 -285.385 70.035 ;
        RECT -284.605 66.675 -284.205 67.875 ;
        RECT -285.105 56.255 -284.825 65.695 ;
        RECT -284.545 56.535 -284.265 66.675 ;
        RECT -283.985 56.255 -283.705 65.695 ;
        RECT -283.425 56.535 -283.145 73.395 ;
        RECT -281.245 70.035 -280.845 71.235 ;
        RECT -282.365 66.675 -281.965 67.875 ;
        RECT -282.865 56.255 -282.585 65.695 ;
        RECT -282.305 56.535 -282.025 66.675 ;
        RECT -281.745 56.255 -281.465 65.695 ;
        RECT -281.185 56.535 -280.905 70.035 ;
        RECT -280.125 66.675 -279.725 67.875 ;
        RECT -280.625 56.255 -280.345 65.695 ;
        RECT -280.065 56.535 -279.785 66.675 ;
        RECT -279.505 56.255 -279.225 65.695 ;
        RECT -278.945 56.535 -278.665 80.115 ;
        RECT -270.045 76.755 -269.645 77.955 ;
        RECT -274.525 73.395 -274.125 74.595 ;
        RECT -276.765 70.035 -276.365 71.235 ;
        RECT -277.885 66.675 -277.485 67.875 ;
        RECT -278.385 56.255 -278.105 65.695 ;
        RECT -277.825 56.535 -277.545 66.675 ;
        RECT -277.265 56.255 -276.985 65.695 ;
        RECT -276.705 56.535 -276.425 70.035 ;
        RECT -275.645 66.675 -275.245 67.875 ;
        RECT -276.145 56.255 -275.865 65.695 ;
        RECT -275.585 56.535 -275.305 66.675 ;
        RECT -275.025 56.255 -274.745 65.695 ;
        RECT -274.465 56.535 -274.185 73.395 ;
        RECT -272.285 70.035 -271.885 71.235 ;
        RECT -273.405 66.675 -273.005 67.875 ;
        RECT -273.905 56.255 -273.625 65.695 ;
        RECT -273.345 56.535 -273.065 66.675 ;
        RECT -272.785 56.255 -272.505 65.695 ;
        RECT -272.225 56.535 -271.945 70.035 ;
        RECT -271.165 66.675 -270.765 67.875 ;
        RECT -271.665 56.255 -271.385 65.695 ;
        RECT -271.105 56.535 -270.825 66.675 ;
        RECT -270.545 56.255 -270.265 65.695 ;
        RECT -269.985 56.535 -269.705 76.755 ;
        RECT -265.565 73.395 -265.165 74.595 ;
        RECT -267.805 70.035 -267.405 71.235 ;
        RECT -268.925 66.675 -268.525 67.875 ;
        RECT -269.425 56.255 -269.145 65.695 ;
        RECT -268.865 56.535 -268.585 66.675 ;
        RECT -268.305 56.255 -268.025 65.695 ;
        RECT -267.745 56.535 -267.465 70.035 ;
        RECT -266.685 66.675 -266.285 67.875 ;
        RECT -267.185 56.255 -266.905 65.695 ;
        RECT -266.625 56.535 -266.345 66.675 ;
        RECT -266.065 56.255 -265.785 65.695 ;
        RECT -265.505 56.535 -265.225 73.395 ;
        RECT -263.325 70.035 -262.925 71.235 ;
        RECT -264.445 66.675 -264.045 67.875 ;
        RECT -264.945 56.255 -264.665 65.695 ;
        RECT -264.385 56.535 -264.105 66.675 ;
        RECT -263.825 56.255 -263.545 65.695 ;
        RECT -263.265 56.535 -262.985 70.035 ;
        RECT -262.205 66.675 -261.805 67.875 ;
        RECT -262.705 56.255 -262.425 65.695 ;
        RECT -262.145 56.535 -261.865 66.675 ;
        RECT -261.585 56.255 -261.305 65.695 ;
        RECT -261.025 56.535 -260.745 86.835 ;
        RECT -225.245 83.475 -224.845 84.675 ;
        RECT -243.165 80.115 -242.765 81.315 ;
        RECT -252.125 76.755 -251.725 77.955 ;
        RECT -256.605 73.395 -256.205 74.595 ;
        RECT -258.845 70.035 -258.445 71.235 ;
        RECT -259.965 66.675 -259.565 67.875 ;
        RECT -260.465 56.255 -260.185 65.695 ;
        RECT -259.905 56.535 -259.625 66.675 ;
        RECT -259.345 56.255 -259.065 65.695 ;
        RECT -258.785 56.535 -258.505 70.035 ;
        RECT -257.725 66.675 -257.325 67.875 ;
        RECT -258.225 56.255 -257.945 65.695 ;
        RECT -257.665 56.535 -257.385 66.675 ;
        RECT -257.105 56.255 -256.825 65.695 ;
        RECT -256.545 56.535 -256.265 73.395 ;
        RECT -254.365 70.035 -253.965 71.235 ;
        RECT -255.485 66.675 -255.085 67.875 ;
        RECT -255.985 56.255 -255.705 65.695 ;
        RECT -255.425 56.535 -255.145 66.675 ;
        RECT -254.865 56.255 -254.585 65.695 ;
        RECT -254.305 56.535 -254.025 70.035 ;
        RECT -253.245 66.675 -252.845 67.875 ;
        RECT -253.745 56.255 -253.465 65.695 ;
        RECT -253.185 56.535 -252.905 66.675 ;
        RECT -252.625 56.255 -252.345 65.695 ;
        RECT -252.065 56.535 -251.785 76.755 ;
        RECT -247.645 73.395 -247.245 74.595 ;
        RECT -249.885 70.035 -249.485 71.235 ;
        RECT -251.005 66.675 -250.605 67.875 ;
        RECT -251.505 56.255 -251.225 65.695 ;
        RECT -250.945 56.535 -250.665 66.675 ;
        RECT -250.385 56.255 -250.105 65.695 ;
        RECT -249.825 56.535 -249.545 70.035 ;
        RECT -248.765 66.675 -248.365 67.875 ;
        RECT -249.265 56.255 -248.985 65.695 ;
        RECT -248.705 56.535 -248.425 66.675 ;
        RECT -248.145 56.255 -247.865 65.695 ;
        RECT -247.585 56.535 -247.305 73.395 ;
        RECT -245.405 70.035 -245.005 71.235 ;
        RECT -246.525 66.675 -246.125 67.875 ;
        RECT -247.025 56.255 -246.745 65.695 ;
        RECT -246.465 56.535 -246.185 66.675 ;
        RECT -245.905 56.255 -245.625 65.695 ;
        RECT -245.345 56.535 -245.065 70.035 ;
        RECT -244.285 66.675 -243.885 67.875 ;
        RECT -244.785 56.255 -244.505 65.695 ;
        RECT -244.225 56.535 -243.945 66.675 ;
        RECT -243.665 56.255 -243.385 65.695 ;
        RECT -243.105 56.535 -242.825 80.115 ;
        RECT -234.205 76.755 -233.805 77.955 ;
        RECT -238.685 73.395 -238.285 74.595 ;
        RECT -240.925 70.035 -240.525 71.235 ;
        RECT -242.045 66.675 -241.645 67.875 ;
        RECT -242.545 56.255 -242.265 65.695 ;
        RECT -241.985 56.535 -241.705 66.675 ;
        RECT -241.425 56.255 -241.145 65.695 ;
        RECT -240.865 56.535 -240.585 70.035 ;
        RECT -239.805 66.675 -239.405 67.875 ;
        RECT -240.305 56.255 -240.025 65.695 ;
        RECT -239.745 56.535 -239.465 66.675 ;
        RECT -239.185 56.255 -238.905 65.695 ;
        RECT -238.625 56.535 -238.345 73.395 ;
        RECT -236.445 70.035 -236.045 71.235 ;
        RECT -237.565 66.675 -237.165 67.875 ;
        RECT -238.065 56.255 -237.785 65.695 ;
        RECT -237.505 56.535 -237.225 66.675 ;
        RECT -236.945 56.255 -236.665 65.695 ;
        RECT -236.385 56.535 -236.105 70.035 ;
        RECT -235.325 66.675 -234.925 67.875 ;
        RECT -235.825 56.255 -235.545 65.695 ;
        RECT -235.265 56.535 -234.985 66.675 ;
        RECT -234.705 56.255 -234.425 65.695 ;
        RECT -234.145 56.535 -233.865 76.755 ;
        RECT -229.725 73.395 -229.325 74.595 ;
        RECT -231.965 70.035 -231.565 71.235 ;
        RECT -233.085 66.675 -232.685 67.875 ;
        RECT -233.585 56.255 -233.305 65.695 ;
        RECT -233.025 56.535 -232.745 66.675 ;
        RECT -232.465 56.255 -232.185 65.695 ;
        RECT -231.905 56.535 -231.625 70.035 ;
        RECT -230.845 66.675 -230.445 67.875 ;
        RECT -231.345 56.255 -231.065 65.695 ;
        RECT -230.785 56.535 -230.505 66.675 ;
        RECT -230.225 56.255 -229.945 65.695 ;
        RECT -229.665 56.535 -229.385 73.395 ;
        RECT -227.485 70.035 -227.085 71.235 ;
        RECT -228.605 66.675 -228.205 67.875 ;
        RECT -229.105 56.255 -228.825 65.695 ;
        RECT -228.545 56.535 -228.265 66.675 ;
        RECT -227.985 56.255 -227.705 65.695 ;
        RECT -227.425 56.535 -227.145 70.035 ;
        RECT -226.365 66.675 -225.965 67.875 ;
        RECT -226.865 56.255 -226.585 65.695 ;
        RECT -226.305 56.535 -226.025 66.675 ;
        RECT -225.745 56.255 -225.465 65.695 ;
        RECT -225.185 56.535 -224.905 83.475 ;
        RECT -207.325 80.115 -206.925 81.315 ;
        RECT -216.285 76.755 -215.885 77.955 ;
        RECT -220.765 73.395 -220.365 74.595 ;
        RECT -223.005 70.035 -222.605 71.235 ;
        RECT -224.125 66.675 -223.725 67.875 ;
        RECT -224.625 56.255 -224.345 65.695 ;
        RECT -224.065 56.535 -223.785 66.675 ;
        RECT -223.505 56.255 -223.225 65.695 ;
        RECT -222.945 56.535 -222.665 70.035 ;
        RECT -221.885 66.675 -221.485 67.875 ;
        RECT -222.385 56.255 -222.105 65.695 ;
        RECT -221.825 56.535 -221.545 66.675 ;
        RECT -221.265 56.255 -220.985 65.695 ;
        RECT -220.705 56.535 -220.425 73.395 ;
        RECT -218.525 70.035 -218.125 71.235 ;
        RECT -219.645 66.675 -219.245 67.875 ;
        RECT -220.145 56.255 -219.865 65.695 ;
        RECT -219.585 56.535 -219.305 66.675 ;
        RECT -219.025 56.255 -218.745 65.695 ;
        RECT -218.465 56.535 -218.185 70.035 ;
        RECT -217.405 66.675 -217.005 67.875 ;
        RECT -217.905 56.255 -217.625 65.695 ;
        RECT -217.345 56.535 -217.065 66.675 ;
        RECT -216.785 56.255 -216.505 65.695 ;
        RECT -216.225 56.535 -215.945 76.755 ;
        RECT -211.805 73.395 -211.405 74.595 ;
        RECT -214.045 70.035 -213.645 71.235 ;
        RECT -215.165 66.675 -214.765 67.875 ;
        RECT -215.665 56.255 -215.385 65.695 ;
        RECT -215.105 56.535 -214.825 66.675 ;
        RECT -214.545 56.255 -214.265 65.695 ;
        RECT -213.985 56.535 -213.705 70.035 ;
        RECT -212.925 66.675 -212.525 67.875 ;
        RECT -213.425 56.255 -213.145 65.695 ;
        RECT -212.865 56.535 -212.585 66.675 ;
        RECT -212.305 56.255 -212.025 65.695 ;
        RECT -211.745 56.535 -211.465 73.395 ;
        RECT -209.565 70.035 -209.165 71.235 ;
        RECT -210.685 66.675 -210.285 67.875 ;
        RECT -211.185 56.255 -210.905 65.695 ;
        RECT -210.625 56.535 -210.345 66.675 ;
        RECT -210.065 56.255 -209.785 65.695 ;
        RECT -209.505 56.535 -209.225 70.035 ;
        RECT -208.445 66.675 -208.045 67.875 ;
        RECT -208.945 56.255 -208.665 65.695 ;
        RECT -208.385 56.535 -208.105 66.675 ;
        RECT -207.825 56.255 -207.545 65.695 ;
        RECT -207.265 56.535 -206.985 80.115 ;
        RECT -198.365 76.755 -197.965 77.955 ;
        RECT -202.845 73.395 -202.445 74.595 ;
        RECT -205.085 70.035 -204.685 71.235 ;
        RECT -206.205 66.675 -205.805 67.875 ;
        RECT -206.705 56.255 -206.425 65.695 ;
        RECT -206.145 56.535 -205.865 66.675 ;
        RECT -205.585 56.255 -205.305 65.695 ;
        RECT -205.025 56.535 -204.745 70.035 ;
        RECT -203.965 66.675 -203.565 67.875 ;
        RECT -204.465 56.255 -204.185 65.695 ;
        RECT -203.905 56.535 -203.625 66.675 ;
        RECT -203.345 56.255 -203.065 65.695 ;
        RECT -202.785 56.535 -202.505 73.395 ;
        RECT -200.605 70.035 -200.205 71.235 ;
        RECT -201.725 66.675 -201.325 67.875 ;
        RECT -202.225 56.255 -201.945 65.695 ;
        RECT -201.665 56.535 -201.385 66.675 ;
        RECT -201.105 56.255 -200.825 65.695 ;
        RECT -200.545 56.535 -200.265 70.035 ;
        RECT -199.485 66.675 -199.085 67.875 ;
        RECT -199.985 56.255 -199.705 65.695 ;
        RECT -199.425 56.535 -199.145 66.675 ;
        RECT -198.865 56.255 -198.585 65.695 ;
        RECT -198.305 56.535 -198.025 76.755 ;
        RECT -193.885 73.395 -193.485 74.595 ;
        RECT -196.125 70.035 -195.725 71.235 ;
        RECT -197.245 66.675 -196.845 67.875 ;
        RECT -197.745 56.255 -197.465 65.695 ;
        RECT -197.185 56.535 -196.905 66.675 ;
        RECT -196.625 56.255 -196.345 65.695 ;
        RECT -196.065 56.535 -195.785 70.035 ;
        RECT -195.005 66.675 -194.605 67.875 ;
        RECT -195.505 56.255 -195.225 65.695 ;
        RECT -194.945 56.535 -194.665 66.675 ;
        RECT -194.385 56.255 -194.105 65.695 ;
        RECT -193.825 56.535 -193.545 73.395 ;
        RECT -191.645 70.035 -191.245 71.235 ;
        RECT -192.765 66.675 -192.365 67.875 ;
        RECT -193.265 56.255 -192.985 65.695 ;
        RECT -192.705 56.535 -192.425 66.675 ;
        RECT -192.145 56.255 -191.865 65.695 ;
        RECT -191.585 56.535 -191.305 70.035 ;
        RECT -190.525 66.675 -190.125 67.875 ;
        RECT -191.025 56.255 -190.745 65.695 ;
        RECT -190.465 56.535 -190.185 66.675 ;
        RECT -189.905 56.255 -189.625 65.695 ;
        RECT -189.345 56.535 -189.065 96.915 ;
        RECT -188.285 93.555 -187.885 94.755 ;
        RECT 120.925 94.355 121.925 94.405 ;
        RECT 120.925 93.955 143.995 94.355 ;
        RECT 120.925 93.905 121.925 93.955 ;
        RECT -188.785 56.255 -188.505 65.695 ;
        RECT -188.225 56.535 -187.945 93.555 ;
        RECT 144.850 93.430 460.000 93.830 ;
        RECT -44.925 90.195 -44.525 91.395 ;
        RECT 120.925 90.995 121.925 91.045 ;
        RECT 120.925 90.595 143.995 90.995 ;
        RECT 120.925 90.545 121.925 90.595 ;
        RECT -116.605 86.835 -116.205 88.035 ;
        RECT -152.445 83.475 -152.045 84.675 ;
        RECT -170.365 80.115 -169.965 81.315 ;
        RECT -179.325 76.755 -178.925 77.955 ;
        RECT -183.805 73.395 -183.405 74.595 ;
        RECT -186.045 70.035 -185.645 71.235 ;
        RECT -187.165 66.675 -186.765 67.875 ;
        RECT -187.665 56.255 -187.385 65.695 ;
        RECT -187.105 56.535 -186.825 66.675 ;
        RECT -186.545 56.255 -186.265 65.695 ;
        RECT -185.985 56.535 -185.705 70.035 ;
        RECT -184.925 66.675 -184.525 67.875 ;
        RECT -185.425 56.255 -185.145 65.695 ;
        RECT -184.865 56.535 -184.585 66.675 ;
        RECT -184.305 56.255 -184.025 65.695 ;
        RECT -183.745 56.535 -183.465 73.395 ;
        RECT -181.565 70.035 -181.165 71.235 ;
        RECT -182.685 66.675 -182.285 67.875 ;
        RECT -183.185 56.255 -182.905 65.695 ;
        RECT -182.625 56.535 -182.345 66.675 ;
        RECT -182.065 56.255 -181.785 65.695 ;
        RECT -181.505 56.535 -181.225 70.035 ;
        RECT -180.445 66.675 -180.045 67.875 ;
        RECT -180.945 56.255 -180.665 65.695 ;
        RECT -180.385 56.535 -180.105 66.675 ;
        RECT -179.825 56.255 -179.545 65.695 ;
        RECT -179.265 56.535 -178.985 76.755 ;
        RECT -174.845 73.395 -174.445 74.595 ;
        RECT -177.085 70.035 -176.685 71.235 ;
        RECT -178.205 66.675 -177.805 67.875 ;
        RECT -178.705 56.255 -178.425 65.695 ;
        RECT -178.145 56.535 -177.865 66.675 ;
        RECT -177.585 56.255 -177.305 65.695 ;
        RECT -177.025 56.535 -176.745 70.035 ;
        RECT -175.965 66.675 -175.565 67.875 ;
        RECT -176.465 56.255 -176.185 65.695 ;
        RECT -175.905 56.535 -175.625 66.675 ;
        RECT -175.345 56.255 -175.065 65.695 ;
        RECT -174.785 56.535 -174.505 73.395 ;
        RECT -172.605 70.035 -172.205 71.235 ;
        RECT -173.725 66.675 -173.325 67.875 ;
        RECT -174.225 56.255 -173.945 65.695 ;
        RECT -173.665 56.535 -173.385 66.675 ;
        RECT -173.105 56.255 -172.825 65.695 ;
        RECT -172.545 56.535 -172.265 70.035 ;
        RECT -171.485 66.675 -171.085 67.875 ;
        RECT -171.985 56.255 -171.705 65.695 ;
        RECT -171.425 56.535 -171.145 66.675 ;
        RECT -170.865 56.255 -170.585 65.695 ;
        RECT -170.305 56.535 -170.025 80.115 ;
        RECT -161.405 76.755 -161.005 77.955 ;
        RECT -165.885 73.395 -165.485 74.595 ;
        RECT -168.125 70.035 -167.725 71.235 ;
        RECT -169.245 66.675 -168.845 67.875 ;
        RECT -169.745 56.255 -169.465 65.695 ;
        RECT -169.185 56.535 -168.905 66.675 ;
        RECT -168.625 56.255 -168.345 65.695 ;
        RECT -168.065 56.535 -167.785 70.035 ;
        RECT -167.005 66.675 -166.605 67.875 ;
        RECT -167.505 56.255 -167.225 65.695 ;
        RECT -166.945 56.535 -166.665 66.675 ;
        RECT -166.385 56.255 -166.105 65.695 ;
        RECT -165.825 56.535 -165.545 73.395 ;
        RECT -163.645 70.035 -163.245 71.235 ;
        RECT -164.765 66.675 -164.365 67.875 ;
        RECT -165.265 56.255 -164.985 65.695 ;
        RECT -164.705 56.535 -164.425 66.675 ;
        RECT -164.145 56.255 -163.865 65.695 ;
        RECT -163.585 56.535 -163.305 70.035 ;
        RECT -162.525 66.675 -162.125 67.875 ;
        RECT -163.025 56.255 -162.745 65.695 ;
        RECT -162.465 56.535 -162.185 66.675 ;
        RECT -161.905 56.255 -161.625 65.695 ;
        RECT -161.345 56.535 -161.065 76.755 ;
        RECT -156.925 73.395 -156.525 74.595 ;
        RECT -159.165 70.035 -158.765 71.235 ;
        RECT -160.285 66.675 -159.885 67.875 ;
        RECT -160.785 56.255 -160.505 65.695 ;
        RECT -160.225 56.535 -159.945 66.675 ;
        RECT -159.665 56.255 -159.385 65.695 ;
        RECT -159.105 56.535 -158.825 70.035 ;
        RECT -158.045 66.675 -157.645 67.875 ;
        RECT -158.545 56.255 -158.265 65.695 ;
        RECT -157.985 56.535 -157.705 66.675 ;
        RECT -157.425 56.255 -157.145 65.695 ;
        RECT -156.865 56.535 -156.585 73.395 ;
        RECT -154.685 70.035 -154.285 71.235 ;
        RECT -155.805 66.675 -155.405 67.875 ;
        RECT -156.305 56.255 -156.025 65.695 ;
        RECT -155.745 56.535 -155.465 66.675 ;
        RECT -155.185 56.255 -154.905 65.695 ;
        RECT -154.625 56.535 -154.345 70.035 ;
        RECT -153.565 66.675 -153.165 67.875 ;
        RECT -154.065 56.255 -153.785 65.695 ;
        RECT -153.505 56.535 -153.225 66.675 ;
        RECT -152.945 56.255 -152.665 65.695 ;
        RECT -152.385 56.535 -152.105 83.475 ;
        RECT -134.525 80.115 -134.125 81.315 ;
        RECT -143.485 76.755 -143.085 77.955 ;
        RECT -147.965 73.395 -147.565 74.595 ;
        RECT -150.205 70.035 -149.805 71.235 ;
        RECT -151.325 66.675 -150.925 67.875 ;
        RECT -151.825 56.255 -151.545 65.695 ;
        RECT -151.265 56.535 -150.985 66.675 ;
        RECT -150.705 56.255 -150.425 65.695 ;
        RECT -150.145 56.535 -149.865 70.035 ;
        RECT -149.085 66.675 -148.685 67.875 ;
        RECT -149.585 56.255 -149.305 65.695 ;
        RECT -149.025 56.535 -148.745 66.675 ;
        RECT -148.465 56.255 -148.185 65.695 ;
        RECT -147.905 56.535 -147.625 73.395 ;
        RECT -145.725 70.035 -145.325 71.235 ;
        RECT -146.845 66.675 -146.445 67.875 ;
        RECT -147.345 56.255 -147.065 65.695 ;
        RECT -146.785 56.535 -146.505 66.675 ;
        RECT -146.225 56.255 -145.945 65.695 ;
        RECT -145.665 56.535 -145.385 70.035 ;
        RECT -144.605 66.675 -144.205 67.875 ;
        RECT -145.105 56.255 -144.825 65.695 ;
        RECT -144.545 56.535 -144.265 66.675 ;
        RECT -143.985 56.255 -143.705 65.695 ;
        RECT -143.425 56.535 -143.145 76.755 ;
        RECT -139.005 73.395 -138.605 74.595 ;
        RECT -141.245 70.035 -140.845 71.235 ;
        RECT -142.365 66.675 -141.965 67.875 ;
        RECT -142.865 56.255 -142.585 65.695 ;
        RECT -142.305 56.535 -142.025 66.675 ;
        RECT -141.745 56.255 -141.465 65.695 ;
        RECT -141.185 56.535 -140.905 70.035 ;
        RECT -140.125 66.675 -139.725 67.875 ;
        RECT -140.625 56.255 -140.345 65.695 ;
        RECT -140.065 56.535 -139.785 66.675 ;
        RECT -139.505 56.255 -139.225 65.695 ;
        RECT -138.945 56.535 -138.665 73.395 ;
        RECT -136.765 70.035 -136.365 71.235 ;
        RECT -137.885 66.675 -137.485 67.875 ;
        RECT -138.385 56.255 -138.105 65.695 ;
        RECT -137.825 56.535 -137.545 66.675 ;
        RECT -137.265 56.255 -136.985 65.695 ;
        RECT -136.705 56.535 -136.425 70.035 ;
        RECT -135.645 66.675 -135.245 67.875 ;
        RECT -136.145 56.255 -135.865 65.695 ;
        RECT -135.585 56.535 -135.305 66.675 ;
        RECT -135.025 56.255 -134.745 65.695 ;
        RECT -134.465 56.535 -134.185 80.115 ;
        RECT -125.565 76.755 -125.165 77.955 ;
        RECT -130.045 73.395 -129.645 74.595 ;
        RECT -132.285 70.035 -131.885 71.235 ;
        RECT -133.405 66.675 -133.005 67.875 ;
        RECT -133.905 56.255 -133.625 65.695 ;
        RECT -133.345 56.535 -133.065 66.675 ;
        RECT -132.785 56.255 -132.505 65.695 ;
        RECT -132.225 56.535 -131.945 70.035 ;
        RECT -131.165 66.675 -130.765 67.875 ;
        RECT -131.665 56.255 -131.385 65.695 ;
        RECT -131.105 56.535 -130.825 66.675 ;
        RECT -130.545 56.255 -130.265 65.695 ;
        RECT -129.985 56.535 -129.705 73.395 ;
        RECT -127.805 70.035 -127.405 71.235 ;
        RECT -128.925 66.675 -128.525 67.875 ;
        RECT -129.425 56.255 -129.145 65.695 ;
        RECT -128.865 56.535 -128.585 66.675 ;
        RECT -128.305 56.255 -128.025 65.695 ;
        RECT -127.745 56.535 -127.465 70.035 ;
        RECT -126.685 66.675 -126.285 67.875 ;
        RECT -127.185 56.255 -126.905 65.695 ;
        RECT -126.625 56.535 -126.345 66.675 ;
        RECT -126.065 56.255 -125.785 65.695 ;
        RECT -125.505 56.535 -125.225 76.755 ;
        RECT -121.085 73.395 -120.685 74.595 ;
        RECT -123.325 70.035 -122.925 71.235 ;
        RECT -124.445 66.675 -124.045 67.875 ;
        RECT -124.945 56.255 -124.665 65.695 ;
        RECT -124.385 56.535 -124.105 66.675 ;
        RECT -123.825 56.255 -123.545 65.695 ;
        RECT -123.265 56.535 -122.985 70.035 ;
        RECT -122.205 66.675 -121.805 67.875 ;
        RECT -122.705 56.255 -122.425 65.695 ;
        RECT -122.145 56.535 -121.865 66.675 ;
        RECT -121.585 56.255 -121.305 65.695 ;
        RECT -121.025 56.535 -120.745 73.395 ;
        RECT -118.845 70.035 -118.445 71.235 ;
        RECT -119.965 66.675 -119.565 67.875 ;
        RECT -120.465 56.255 -120.185 65.695 ;
        RECT -119.905 56.535 -119.625 66.675 ;
        RECT -119.345 56.255 -119.065 65.695 ;
        RECT -118.785 56.535 -118.505 70.035 ;
        RECT -117.725 66.675 -117.325 67.875 ;
        RECT -118.225 56.255 -117.945 65.695 ;
        RECT -117.665 56.535 -117.385 66.675 ;
        RECT -117.105 56.255 -116.825 65.695 ;
        RECT -116.545 56.535 -116.265 86.835 ;
        RECT -80.765 83.475 -80.365 84.675 ;
        RECT -98.685 80.115 -98.285 81.315 ;
        RECT -107.645 76.755 -107.245 77.955 ;
        RECT -112.125 73.395 -111.725 74.595 ;
        RECT -114.365 70.035 -113.965 71.235 ;
        RECT -115.485 66.675 -115.085 67.875 ;
        RECT -115.985 56.255 -115.705 65.695 ;
        RECT -115.425 56.535 -115.145 66.675 ;
        RECT -114.865 56.255 -114.585 65.695 ;
        RECT -114.305 56.535 -114.025 70.035 ;
        RECT -113.245 66.675 -112.845 67.875 ;
        RECT -113.745 56.255 -113.465 65.695 ;
        RECT -113.185 56.535 -112.905 66.675 ;
        RECT -112.625 56.255 -112.345 65.695 ;
        RECT -112.065 56.535 -111.785 73.395 ;
        RECT -109.885 70.035 -109.485 71.235 ;
        RECT -111.005 66.675 -110.605 67.875 ;
        RECT -111.505 56.255 -111.225 65.695 ;
        RECT -110.945 56.535 -110.665 66.675 ;
        RECT -110.385 56.255 -110.105 65.695 ;
        RECT -109.825 56.535 -109.545 70.035 ;
        RECT -108.765 66.675 -108.365 67.875 ;
        RECT -109.265 56.255 -108.985 65.695 ;
        RECT -108.705 56.535 -108.425 66.675 ;
        RECT -108.145 56.255 -107.865 65.695 ;
        RECT -107.585 56.535 -107.305 76.755 ;
        RECT -103.165 73.395 -102.765 74.595 ;
        RECT -105.405 70.035 -105.005 71.235 ;
        RECT -106.525 66.675 -106.125 67.875 ;
        RECT -107.025 56.255 -106.745 65.695 ;
        RECT -106.465 56.535 -106.185 66.675 ;
        RECT -105.905 56.255 -105.625 65.695 ;
        RECT -105.345 56.535 -105.065 70.035 ;
        RECT -104.285 66.675 -103.885 67.875 ;
        RECT -104.785 56.255 -104.505 65.695 ;
        RECT -104.225 56.535 -103.945 66.675 ;
        RECT -103.665 56.255 -103.385 65.695 ;
        RECT -103.105 56.535 -102.825 73.395 ;
        RECT -100.925 70.035 -100.525 71.235 ;
        RECT -102.045 66.675 -101.645 67.875 ;
        RECT -102.545 56.255 -102.265 65.695 ;
        RECT -101.985 56.535 -101.705 66.675 ;
        RECT -101.425 56.255 -101.145 65.695 ;
        RECT -100.865 56.535 -100.585 70.035 ;
        RECT -99.805 66.675 -99.405 67.875 ;
        RECT -100.305 56.255 -100.025 65.695 ;
        RECT -99.745 56.535 -99.465 66.675 ;
        RECT -99.185 56.255 -98.905 65.695 ;
        RECT -98.625 56.535 -98.345 80.115 ;
        RECT -89.725 76.755 -89.325 77.955 ;
        RECT -94.205 73.395 -93.805 74.595 ;
        RECT -96.445 70.035 -96.045 71.235 ;
        RECT -97.565 66.675 -97.165 67.875 ;
        RECT -98.065 56.255 -97.785 65.695 ;
        RECT -97.505 56.535 -97.225 66.675 ;
        RECT -96.945 56.255 -96.665 65.695 ;
        RECT -96.385 56.535 -96.105 70.035 ;
        RECT -95.325 66.675 -94.925 67.875 ;
        RECT -95.825 56.255 -95.545 65.695 ;
        RECT -95.265 56.535 -94.985 66.675 ;
        RECT -94.705 56.255 -94.425 65.695 ;
        RECT -94.145 56.535 -93.865 73.395 ;
        RECT -91.965 70.035 -91.565 71.235 ;
        RECT -93.085 66.675 -92.685 67.875 ;
        RECT -93.585 56.255 -93.305 65.695 ;
        RECT -93.025 56.535 -92.745 66.675 ;
        RECT -92.465 56.255 -92.185 65.695 ;
        RECT -91.905 56.535 -91.625 70.035 ;
        RECT -90.845 66.675 -90.445 67.875 ;
        RECT -91.345 56.255 -91.065 65.695 ;
        RECT -90.785 56.535 -90.505 66.675 ;
        RECT -90.225 56.255 -89.945 65.695 ;
        RECT -89.665 56.535 -89.385 76.755 ;
        RECT -85.245 73.395 -84.845 74.595 ;
        RECT -87.485 70.035 -87.085 71.235 ;
        RECT -88.605 66.675 -88.205 67.875 ;
        RECT -89.105 56.255 -88.825 65.695 ;
        RECT -88.545 56.535 -88.265 66.675 ;
        RECT -87.985 56.255 -87.705 65.695 ;
        RECT -87.425 56.535 -87.145 70.035 ;
        RECT -86.365 66.675 -85.965 67.875 ;
        RECT -86.865 56.255 -86.585 65.695 ;
        RECT -86.305 56.535 -86.025 66.675 ;
        RECT -85.745 56.255 -85.465 65.695 ;
        RECT -85.185 56.535 -84.905 73.395 ;
        RECT -83.005 70.035 -82.605 71.235 ;
        RECT -84.125 66.675 -83.725 67.875 ;
        RECT -84.625 56.255 -84.345 65.695 ;
        RECT -84.065 56.535 -83.785 66.675 ;
        RECT -83.505 56.255 -83.225 65.695 ;
        RECT -82.945 56.535 -82.665 70.035 ;
        RECT -81.885 66.675 -81.485 67.875 ;
        RECT -82.385 56.255 -82.105 65.695 ;
        RECT -81.825 56.535 -81.545 66.675 ;
        RECT -81.265 56.255 -80.985 65.695 ;
        RECT -80.705 56.535 -80.425 83.475 ;
        RECT -62.845 80.115 -62.445 81.315 ;
        RECT -71.805 76.755 -71.405 77.955 ;
        RECT -76.285 73.395 -75.885 74.595 ;
        RECT -78.525 70.035 -78.125 71.235 ;
        RECT -79.645 66.675 -79.245 67.875 ;
        RECT -80.145 56.255 -79.865 65.695 ;
        RECT -79.585 56.535 -79.305 66.675 ;
        RECT -79.025 56.255 -78.745 65.695 ;
        RECT -78.465 56.535 -78.185 70.035 ;
        RECT -77.405 66.675 -77.005 67.875 ;
        RECT -77.905 56.255 -77.625 65.695 ;
        RECT -77.345 56.535 -77.065 66.675 ;
        RECT -76.785 56.255 -76.505 65.695 ;
        RECT -76.225 56.535 -75.945 73.395 ;
        RECT -74.045 70.035 -73.645 71.235 ;
        RECT -75.165 66.675 -74.765 67.875 ;
        RECT -75.665 56.255 -75.385 65.695 ;
        RECT -75.105 56.535 -74.825 66.675 ;
        RECT -74.545 56.255 -74.265 65.695 ;
        RECT -73.985 56.535 -73.705 70.035 ;
        RECT -72.925 66.675 -72.525 67.875 ;
        RECT -73.425 56.255 -73.145 65.695 ;
        RECT -72.865 56.535 -72.585 66.675 ;
        RECT -72.305 56.255 -72.025 65.695 ;
        RECT -71.745 56.535 -71.465 76.755 ;
        RECT -67.325 73.395 -66.925 74.595 ;
        RECT -69.565 70.035 -69.165 71.235 ;
        RECT -70.685 66.675 -70.285 67.875 ;
        RECT -71.185 56.255 -70.905 65.695 ;
        RECT -70.625 56.535 -70.345 66.675 ;
        RECT -70.065 56.255 -69.785 65.695 ;
        RECT -69.505 56.535 -69.225 70.035 ;
        RECT -68.445 66.675 -68.045 67.875 ;
        RECT -68.945 56.255 -68.665 65.695 ;
        RECT -68.385 56.535 -68.105 66.675 ;
        RECT -67.825 56.255 -67.545 65.695 ;
        RECT -67.265 56.535 -66.985 73.395 ;
        RECT -65.085 70.035 -64.685 71.235 ;
        RECT -66.205 66.675 -65.805 67.875 ;
        RECT -66.705 56.255 -66.425 65.695 ;
        RECT -66.145 56.535 -65.865 66.675 ;
        RECT -65.585 56.255 -65.305 65.695 ;
        RECT -65.025 56.535 -64.745 70.035 ;
        RECT -63.965 66.675 -63.565 67.875 ;
        RECT -64.465 56.255 -64.185 65.695 ;
        RECT -63.905 56.535 -63.625 66.675 ;
        RECT -63.345 56.255 -63.065 65.695 ;
        RECT -62.785 56.535 -62.505 80.115 ;
        RECT -53.885 76.755 -53.485 77.955 ;
        RECT -58.365 73.395 -57.965 74.595 ;
        RECT -60.605 70.035 -60.205 71.235 ;
        RECT -61.725 66.675 -61.325 67.875 ;
        RECT -62.225 56.255 -61.945 65.695 ;
        RECT -61.665 56.535 -61.385 66.675 ;
        RECT -61.105 56.255 -60.825 65.695 ;
        RECT -60.545 56.535 -60.265 70.035 ;
        RECT -59.485 66.675 -59.085 67.875 ;
        RECT -59.985 56.255 -59.705 65.695 ;
        RECT -59.425 56.535 -59.145 66.675 ;
        RECT -58.865 56.255 -58.585 65.695 ;
        RECT -58.305 56.535 -58.025 73.395 ;
        RECT -56.125 70.035 -55.725 71.235 ;
        RECT -57.245 66.675 -56.845 67.875 ;
        RECT -57.745 56.255 -57.465 65.695 ;
        RECT -57.185 56.535 -56.905 66.675 ;
        RECT -56.625 56.255 -56.345 65.695 ;
        RECT -56.065 56.535 -55.785 70.035 ;
        RECT -55.005 66.675 -54.605 67.875 ;
        RECT -55.505 56.255 -55.225 65.695 ;
        RECT -54.945 56.535 -54.665 66.675 ;
        RECT -54.385 56.255 -54.105 65.695 ;
        RECT -53.825 56.535 -53.545 76.755 ;
        RECT -49.405 73.395 -49.005 74.595 ;
        RECT -51.645 70.035 -51.245 71.235 ;
        RECT -52.765 66.675 -52.365 67.875 ;
        RECT -53.265 56.255 -52.985 65.695 ;
        RECT -52.705 56.535 -52.425 66.675 ;
        RECT -52.145 56.255 -51.865 65.695 ;
        RECT -51.585 56.535 -51.305 70.035 ;
        RECT -50.525 66.675 -50.125 67.875 ;
        RECT -51.025 56.255 -50.745 65.695 ;
        RECT -50.465 56.535 -50.185 66.675 ;
        RECT -49.905 56.255 -49.625 65.695 ;
        RECT -49.345 56.535 -49.065 73.395 ;
        RECT -47.165 70.035 -46.765 71.235 ;
        RECT -48.285 66.675 -47.885 67.875 ;
        RECT -48.785 56.255 -48.505 65.695 ;
        RECT -48.225 56.535 -47.945 66.675 ;
        RECT -47.665 56.255 -47.385 65.695 ;
        RECT -47.105 56.535 -46.825 70.035 ;
        RECT -46.045 66.675 -45.645 67.875 ;
        RECT -46.545 56.255 -46.265 65.695 ;
        RECT -45.985 56.535 -45.705 66.675 ;
        RECT -45.425 56.255 -45.145 65.695 ;
        RECT -44.865 56.535 -44.585 90.195 ;
        RECT 144.850 90.070 442.080 90.470 ;
        RECT 26.755 86.835 27.155 88.035 ;
        RECT 120.925 87.635 121.925 87.685 ;
        RECT 120.925 87.235 143.995 87.635 ;
        RECT 120.925 87.185 121.925 87.235 ;
        RECT -9.085 83.475 -8.685 84.675 ;
        RECT -27.005 80.115 -26.605 81.315 ;
        RECT -35.965 76.755 -35.565 77.955 ;
        RECT -40.445 73.395 -40.045 74.595 ;
        RECT -42.685 70.035 -42.285 71.235 ;
        RECT -43.805 66.675 -43.405 67.875 ;
        RECT -44.305 56.255 -44.025 65.695 ;
        RECT -43.745 56.535 -43.465 66.675 ;
        RECT -43.185 56.255 -42.905 65.695 ;
        RECT -42.625 56.535 -42.345 70.035 ;
        RECT -41.565 66.675 -41.165 67.875 ;
        RECT -42.065 56.255 -41.785 65.695 ;
        RECT -41.505 56.535 -41.225 66.675 ;
        RECT -40.945 56.255 -40.665 65.695 ;
        RECT -40.385 56.535 -40.105 73.395 ;
        RECT -38.205 70.035 -37.805 71.235 ;
        RECT -39.325 66.675 -38.925 67.875 ;
        RECT -39.825 56.255 -39.545 65.695 ;
        RECT -39.265 56.535 -38.985 66.675 ;
        RECT -38.705 56.255 -38.425 65.695 ;
        RECT -38.145 56.535 -37.865 70.035 ;
        RECT -37.085 66.675 -36.685 67.875 ;
        RECT -37.585 56.255 -37.305 65.695 ;
        RECT -37.025 56.535 -36.745 66.675 ;
        RECT -36.465 56.255 -36.185 65.695 ;
        RECT -35.905 56.535 -35.625 76.755 ;
        RECT -31.485 73.395 -31.085 74.595 ;
        RECT -33.725 70.035 -33.325 71.235 ;
        RECT -34.845 66.675 -34.445 67.875 ;
        RECT -35.345 56.255 -35.065 65.695 ;
        RECT -34.785 56.535 -34.505 66.675 ;
        RECT -34.225 56.255 -33.945 65.695 ;
        RECT -33.665 56.535 -33.385 70.035 ;
        RECT -32.605 66.675 -32.205 67.875 ;
        RECT -33.105 56.255 -32.825 65.695 ;
        RECT -32.545 56.535 -32.265 66.675 ;
        RECT -31.985 56.255 -31.705 65.695 ;
        RECT -31.425 56.535 -31.145 73.395 ;
        RECT -29.245 70.035 -28.845 71.235 ;
        RECT -30.365 66.675 -29.965 67.875 ;
        RECT -30.865 56.255 -30.585 65.695 ;
        RECT -30.305 56.535 -30.025 66.675 ;
        RECT -29.745 56.255 -29.465 65.695 ;
        RECT -29.185 56.535 -28.905 70.035 ;
        RECT -28.125 66.675 -27.725 67.875 ;
        RECT -28.625 56.255 -28.345 65.695 ;
        RECT -28.065 56.535 -27.785 66.675 ;
        RECT -27.505 56.255 -27.225 65.695 ;
        RECT -26.945 56.535 -26.665 80.115 ;
        RECT -18.045 76.755 -17.645 77.955 ;
        RECT -22.525 73.395 -22.125 74.595 ;
        RECT -24.765 70.035 -24.365 71.235 ;
        RECT -25.885 66.675 -25.485 67.875 ;
        RECT -26.385 56.255 -26.105 65.695 ;
        RECT -25.825 56.535 -25.545 66.675 ;
        RECT -25.265 56.255 -24.985 65.695 ;
        RECT -24.705 56.535 -24.425 70.035 ;
        RECT -23.645 66.675 -23.245 67.875 ;
        RECT -24.145 56.255 -23.865 65.695 ;
        RECT -23.585 56.535 -23.305 66.675 ;
        RECT -23.025 56.255 -22.745 65.695 ;
        RECT -22.465 56.535 -22.185 73.395 ;
        RECT -20.285 70.035 -19.885 71.235 ;
        RECT -21.405 66.675 -21.005 67.875 ;
        RECT -21.905 56.255 -21.625 65.695 ;
        RECT -21.345 56.535 -21.065 66.675 ;
        RECT -20.785 56.255 -20.505 65.695 ;
        RECT -20.225 56.535 -19.945 70.035 ;
        RECT -19.165 66.675 -18.765 67.875 ;
        RECT -19.665 56.255 -19.385 65.695 ;
        RECT -19.105 56.535 -18.825 66.675 ;
        RECT -18.545 56.255 -18.265 65.695 ;
        RECT -17.985 56.535 -17.705 76.755 ;
        RECT -13.565 73.395 -13.165 74.595 ;
        RECT -15.805 70.035 -15.405 71.235 ;
        RECT -16.925 66.675 -16.525 67.875 ;
        RECT -17.425 56.255 -17.145 65.695 ;
        RECT -16.865 56.535 -16.585 66.675 ;
        RECT -16.305 56.255 -16.025 65.695 ;
        RECT -15.745 56.535 -15.465 70.035 ;
        RECT -14.685 66.675 -14.285 67.875 ;
        RECT -15.185 56.255 -14.905 65.695 ;
        RECT -14.625 56.535 -14.345 66.675 ;
        RECT -14.065 56.255 -13.785 65.695 ;
        RECT -13.505 56.535 -13.225 73.395 ;
        RECT -11.325 70.035 -10.925 71.235 ;
        RECT -12.445 66.675 -12.045 67.875 ;
        RECT -12.945 56.255 -12.665 65.695 ;
        RECT -12.385 56.535 -12.105 66.675 ;
        RECT -11.825 56.255 -11.545 65.695 ;
        RECT -11.265 56.535 -10.985 70.035 ;
        RECT -10.205 66.675 -9.805 67.875 ;
        RECT -10.705 56.255 -10.425 65.695 ;
        RECT -10.145 56.535 -9.865 66.675 ;
        RECT -9.585 56.255 -9.305 65.695 ;
        RECT -9.025 56.535 -8.745 83.475 ;
        RECT 8.835 80.115 9.235 81.315 ;
        RECT -0.125 76.755 0.275 77.955 ;
        RECT -4.605 73.395 -4.205 74.595 ;
        RECT -6.845 70.035 -6.445 71.235 ;
        RECT -7.965 66.675 -7.565 67.875 ;
        RECT -8.465 56.255 -8.185 65.695 ;
        RECT -7.905 56.535 -7.625 66.675 ;
        RECT -7.345 56.255 -7.065 65.695 ;
        RECT -6.785 56.535 -6.505 70.035 ;
        RECT -5.725 66.675 -5.325 67.875 ;
        RECT -6.225 56.255 -5.945 65.695 ;
        RECT -5.665 56.535 -5.385 66.675 ;
        RECT -5.105 56.255 -4.825 65.695 ;
        RECT -4.545 56.535 -4.265 73.395 ;
        RECT -2.365 70.035 -1.965 71.235 ;
        RECT -3.485 66.675 -3.085 67.875 ;
        RECT -3.985 56.255 -3.705 65.695 ;
        RECT -3.425 56.535 -3.145 66.675 ;
        RECT -2.865 56.255 -2.585 65.695 ;
        RECT -2.305 56.535 -2.025 70.035 ;
        RECT -1.245 66.675 -0.845 67.875 ;
        RECT -1.745 56.255 -1.465 65.695 ;
        RECT -1.185 56.535 -0.905 66.675 ;
        RECT -0.625 56.255 -0.345 65.695 ;
        RECT -0.065 56.535 0.215 76.755 ;
        RECT 4.355 73.395 4.755 74.595 ;
        RECT 2.115 70.035 2.515 71.235 ;
        RECT 0.995 66.675 1.395 67.875 ;
        RECT 0.495 56.255 0.775 65.695 ;
        RECT 1.055 56.535 1.335 66.675 ;
        RECT 1.615 56.255 1.895 65.695 ;
        RECT 2.175 56.535 2.455 70.035 ;
        RECT 3.235 66.675 3.635 67.875 ;
        RECT 2.735 56.255 3.015 65.695 ;
        RECT 3.295 56.535 3.575 66.675 ;
        RECT 3.855 56.255 4.135 65.695 ;
        RECT 4.415 56.535 4.695 73.395 ;
        RECT 6.595 70.035 6.995 71.235 ;
        RECT 5.475 66.675 5.875 67.875 ;
        RECT 4.975 56.255 5.255 65.695 ;
        RECT 5.535 56.535 5.815 66.675 ;
        RECT 6.095 56.255 6.375 65.695 ;
        RECT 6.655 56.535 6.935 70.035 ;
        RECT 7.715 66.675 8.115 67.875 ;
        RECT 7.215 56.255 7.495 65.695 ;
        RECT 7.775 56.535 8.055 66.675 ;
        RECT 8.335 56.255 8.615 65.695 ;
        RECT 8.895 56.535 9.175 80.115 ;
        RECT 17.795 76.755 18.195 77.955 ;
        RECT 13.315 73.395 13.715 74.595 ;
        RECT 11.075 70.035 11.475 71.235 ;
        RECT 9.955 66.675 10.355 67.875 ;
        RECT 9.455 56.255 9.735 65.695 ;
        RECT 10.015 56.535 10.295 66.675 ;
        RECT 10.575 56.255 10.855 65.695 ;
        RECT 11.135 56.535 11.415 70.035 ;
        RECT 12.195 66.675 12.595 67.875 ;
        RECT 11.695 56.255 11.975 65.695 ;
        RECT 12.255 56.535 12.535 66.675 ;
        RECT 12.815 56.255 13.095 65.695 ;
        RECT 13.375 56.535 13.655 73.395 ;
        RECT 15.555 70.035 15.955 71.235 ;
        RECT 14.435 66.675 14.835 67.875 ;
        RECT 13.935 56.255 14.215 65.695 ;
        RECT 14.495 56.535 14.775 66.675 ;
        RECT 15.055 56.255 15.335 65.695 ;
        RECT 15.615 56.535 15.895 70.035 ;
        RECT 16.675 66.675 17.075 67.875 ;
        RECT 16.175 56.255 16.455 65.695 ;
        RECT 16.735 56.535 17.015 66.675 ;
        RECT 17.295 56.255 17.575 65.695 ;
        RECT 17.855 56.535 18.135 76.755 ;
        RECT 22.275 73.395 22.675 74.595 ;
        RECT 20.035 70.035 20.435 71.235 ;
        RECT 18.915 66.675 19.315 67.875 ;
        RECT 18.415 56.255 18.695 65.695 ;
        RECT 18.975 56.535 19.255 66.675 ;
        RECT 19.535 56.255 19.815 65.695 ;
        RECT 20.095 56.535 20.375 70.035 ;
        RECT 21.155 66.675 21.555 67.875 ;
        RECT 20.655 56.255 20.935 65.695 ;
        RECT 21.215 56.535 21.495 66.675 ;
        RECT 21.775 56.255 22.055 65.695 ;
        RECT 22.335 56.535 22.615 73.395 ;
        RECT 24.515 70.035 24.915 71.235 ;
        RECT 23.395 66.675 23.795 67.875 ;
        RECT 22.895 56.255 23.175 65.695 ;
        RECT 23.455 56.535 23.735 66.675 ;
        RECT 24.015 56.255 24.295 65.695 ;
        RECT 24.575 56.535 24.855 70.035 ;
        RECT 25.635 66.675 26.035 67.875 ;
        RECT 25.135 56.255 25.415 65.695 ;
        RECT 25.695 56.535 25.975 66.675 ;
        RECT 26.255 56.255 26.535 65.695 ;
        RECT 26.815 56.535 27.095 86.835 ;
        RECT 144.850 86.710 424.160 87.110 ;
        RECT 62.595 83.475 62.995 84.675 ;
        RECT 120.925 84.275 121.925 84.325 ;
        RECT 120.925 83.875 143.995 84.275 ;
        RECT 120.925 83.825 121.925 83.875 ;
        RECT 44.675 80.115 45.075 81.315 ;
        RECT 35.715 76.755 36.115 77.955 ;
        RECT 31.235 73.395 31.635 74.595 ;
        RECT 28.995 70.035 29.395 71.235 ;
        RECT 27.875 66.675 28.275 67.875 ;
        RECT 27.375 56.255 27.655 65.695 ;
        RECT 27.935 56.535 28.215 66.675 ;
        RECT 28.495 56.255 28.775 65.695 ;
        RECT 29.055 56.535 29.335 70.035 ;
        RECT 30.115 66.675 30.515 67.875 ;
        RECT 29.615 56.255 29.895 65.695 ;
        RECT 30.175 56.535 30.455 66.675 ;
        RECT 30.735 56.255 31.015 65.695 ;
        RECT 31.295 56.535 31.575 73.395 ;
        RECT 33.475 70.035 33.875 71.235 ;
        RECT 32.355 66.675 32.755 67.875 ;
        RECT 31.855 56.255 32.135 65.695 ;
        RECT 32.415 56.535 32.695 66.675 ;
        RECT 32.975 56.255 33.255 65.695 ;
        RECT 33.535 56.535 33.815 70.035 ;
        RECT 34.595 66.675 34.995 67.875 ;
        RECT 34.095 56.255 34.375 65.695 ;
        RECT 34.655 56.535 34.935 66.675 ;
        RECT 35.215 56.255 35.495 65.695 ;
        RECT 35.775 56.535 36.055 76.755 ;
        RECT 40.195 73.395 40.595 74.595 ;
        RECT 37.955 70.035 38.355 71.235 ;
        RECT 36.835 66.675 37.235 67.875 ;
        RECT 36.335 56.255 36.615 65.695 ;
        RECT 36.895 56.535 37.175 66.675 ;
        RECT 37.455 56.255 37.735 65.695 ;
        RECT 38.015 56.535 38.295 70.035 ;
        RECT 39.075 66.675 39.475 67.875 ;
        RECT 38.575 56.255 38.855 65.695 ;
        RECT 39.135 56.535 39.415 66.675 ;
        RECT 39.695 56.255 39.975 65.695 ;
        RECT 40.255 56.535 40.535 73.395 ;
        RECT 42.435 70.035 42.835 71.235 ;
        RECT 41.315 66.675 41.715 67.875 ;
        RECT 40.815 56.255 41.095 65.695 ;
        RECT 41.375 56.535 41.655 66.675 ;
        RECT 41.935 56.255 42.215 65.695 ;
        RECT 42.495 56.535 42.775 70.035 ;
        RECT 43.555 66.675 43.955 67.875 ;
        RECT 43.055 56.255 43.335 65.695 ;
        RECT 43.615 56.535 43.895 66.675 ;
        RECT 44.175 56.255 44.455 65.695 ;
        RECT 44.735 56.535 45.015 80.115 ;
        RECT 53.635 76.755 54.035 77.955 ;
        RECT 49.155 73.395 49.555 74.595 ;
        RECT 46.915 70.035 47.315 71.235 ;
        RECT 45.795 66.675 46.195 67.875 ;
        RECT 45.295 56.255 45.575 65.695 ;
        RECT 45.855 56.535 46.135 66.675 ;
        RECT 46.415 56.255 46.695 65.695 ;
        RECT 46.975 56.535 47.255 70.035 ;
        RECT 48.035 66.675 48.435 67.875 ;
        RECT 47.535 56.255 47.815 65.695 ;
        RECT 48.095 56.535 48.375 66.675 ;
        RECT 48.655 56.255 48.935 65.695 ;
        RECT 49.215 56.535 49.495 73.395 ;
        RECT 51.395 70.035 51.795 71.235 ;
        RECT 50.275 66.675 50.675 67.875 ;
        RECT 49.775 56.255 50.055 65.695 ;
        RECT 50.335 56.535 50.615 66.675 ;
        RECT 50.895 56.255 51.175 65.695 ;
        RECT 51.455 56.535 51.735 70.035 ;
        RECT 52.515 66.675 52.915 67.875 ;
        RECT 52.015 56.255 52.295 65.695 ;
        RECT 52.575 56.535 52.855 66.675 ;
        RECT 53.135 56.255 53.415 65.695 ;
        RECT 53.695 56.535 53.975 76.755 ;
        RECT 58.115 73.395 58.515 74.595 ;
        RECT 55.875 70.035 56.275 71.235 ;
        RECT 54.755 66.675 55.155 67.875 ;
        RECT 54.255 56.255 54.535 65.695 ;
        RECT 54.815 56.535 55.095 66.675 ;
        RECT 55.375 56.255 55.655 65.695 ;
        RECT 55.935 56.535 56.215 70.035 ;
        RECT 56.995 66.675 57.395 67.875 ;
        RECT 56.495 56.255 56.775 65.695 ;
        RECT 57.055 56.535 57.335 66.675 ;
        RECT 57.615 56.255 57.895 65.695 ;
        RECT 58.175 56.535 58.455 73.395 ;
        RECT 60.355 70.035 60.755 71.235 ;
        RECT 59.235 66.675 59.635 67.875 ;
        RECT 58.735 56.255 59.015 65.695 ;
        RECT 59.295 56.535 59.575 66.675 ;
        RECT 59.855 56.255 60.135 65.695 ;
        RECT 60.415 56.535 60.695 70.035 ;
        RECT 61.475 66.675 61.875 67.875 ;
        RECT 60.975 56.255 61.255 65.695 ;
        RECT 61.535 56.535 61.815 66.675 ;
        RECT 62.095 56.255 62.375 65.695 ;
        RECT 62.655 56.535 62.935 83.475 ;
        RECT 144.850 83.350 406.240 83.750 ;
        RECT 80.515 80.115 80.915 81.315 ;
        RECT 120.925 80.915 121.925 80.965 ;
        RECT 120.925 80.515 143.995 80.915 ;
        RECT 120.925 80.465 121.925 80.515 ;
        RECT 71.555 76.755 71.955 77.955 ;
        RECT 67.075 73.395 67.475 74.595 ;
        RECT 64.835 70.035 65.235 71.235 ;
        RECT 63.715 66.675 64.115 67.875 ;
        RECT 63.215 56.255 63.495 65.695 ;
        RECT 63.775 56.535 64.055 66.675 ;
        RECT 64.335 56.255 64.615 65.695 ;
        RECT 64.895 56.535 65.175 70.035 ;
        RECT 65.955 66.675 66.355 67.875 ;
        RECT 65.455 56.255 65.735 65.695 ;
        RECT 66.015 56.535 66.295 66.675 ;
        RECT 66.575 56.255 66.855 65.695 ;
        RECT 67.135 56.535 67.415 73.395 ;
        RECT 69.315 70.035 69.715 71.235 ;
        RECT 68.195 66.675 68.595 67.875 ;
        RECT 67.695 56.255 67.975 65.695 ;
        RECT 68.255 56.535 68.535 66.675 ;
        RECT 68.815 56.255 69.095 65.695 ;
        RECT 69.375 56.535 69.655 70.035 ;
        RECT 70.435 66.675 70.835 67.875 ;
        RECT 69.935 56.255 70.215 65.695 ;
        RECT 70.495 56.535 70.775 66.675 ;
        RECT 71.055 56.255 71.335 65.695 ;
        RECT 71.615 56.535 71.895 76.755 ;
        RECT 76.035 73.395 76.435 74.595 ;
        RECT 73.795 70.035 74.195 71.235 ;
        RECT 72.675 66.675 73.075 67.875 ;
        RECT 72.175 56.255 72.455 65.695 ;
        RECT 72.735 56.535 73.015 66.675 ;
        RECT 73.295 56.255 73.575 65.695 ;
        RECT 73.855 56.535 74.135 70.035 ;
        RECT 74.915 66.675 75.315 67.875 ;
        RECT 74.415 56.255 74.695 65.695 ;
        RECT 74.975 56.535 75.255 66.675 ;
        RECT 75.535 56.255 75.815 65.695 ;
        RECT 76.095 56.535 76.375 73.395 ;
        RECT 78.275 70.035 78.675 71.235 ;
        RECT 77.155 66.675 77.555 67.875 ;
        RECT 76.655 56.255 76.935 65.695 ;
        RECT 77.215 56.535 77.495 66.675 ;
        RECT 77.775 56.255 78.055 65.695 ;
        RECT 78.335 56.535 78.615 70.035 ;
        RECT 79.395 66.675 79.795 67.875 ;
        RECT 78.895 56.255 79.175 65.695 ;
        RECT 79.455 56.535 79.735 66.675 ;
        RECT 80.015 56.255 80.295 65.695 ;
        RECT 80.575 56.535 80.855 80.115 ;
        RECT 144.850 79.990 388.320 80.390 ;
        RECT 89.475 76.755 89.875 77.955 ;
        RECT 120.925 77.555 121.925 77.605 ;
        RECT 120.925 77.155 143.995 77.555 ;
        RECT 120.925 77.105 121.925 77.155 ;
        RECT 84.995 73.395 85.395 74.595 ;
        RECT 82.755 70.035 83.155 71.235 ;
        RECT 81.635 66.675 82.035 67.875 ;
        RECT 81.135 56.255 81.415 65.695 ;
        RECT 81.695 56.535 81.975 66.675 ;
        RECT 82.255 56.255 82.535 65.695 ;
        RECT 82.815 56.535 83.095 70.035 ;
        RECT 83.875 66.675 84.275 67.875 ;
        RECT 83.375 56.255 83.655 65.695 ;
        RECT 83.935 56.535 84.215 66.675 ;
        RECT 84.495 56.255 84.775 65.695 ;
        RECT 85.055 56.535 85.335 73.395 ;
        RECT 87.235 70.035 87.635 71.235 ;
        RECT 86.115 66.675 86.515 67.875 ;
        RECT 85.615 56.255 85.895 65.695 ;
        RECT 86.175 56.535 86.455 66.675 ;
        RECT 86.735 56.255 87.015 65.695 ;
        RECT 87.295 56.535 87.575 70.035 ;
        RECT 88.355 66.675 88.755 67.875 ;
        RECT 87.855 56.255 88.135 65.695 ;
        RECT 88.415 56.535 88.695 66.675 ;
        RECT 88.975 56.255 89.255 65.695 ;
        RECT 89.535 56.535 89.815 76.755 ;
        RECT 144.850 76.630 370.400 77.030 ;
        RECT 93.955 73.395 94.355 74.595 ;
        RECT 120.925 74.195 121.925 74.245 ;
        RECT 120.925 73.795 143.995 74.195 ;
        RECT 120.925 73.745 121.925 73.795 ;
        RECT 91.715 70.035 92.115 71.235 ;
        RECT 90.595 66.675 90.995 67.875 ;
        RECT 90.095 56.255 90.375 65.695 ;
        RECT 90.655 56.535 90.935 66.675 ;
        RECT 91.215 56.255 91.495 65.695 ;
        RECT 91.775 56.535 92.055 70.035 ;
        RECT 92.835 66.675 93.235 67.875 ;
        RECT 92.335 56.255 92.615 65.695 ;
        RECT 92.895 56.535 93.175 66.675 ;
        RECT 93.455 56.255 93.735 65.695 ;
        RECT 94.015 56.535 94.295 73.395 ;
        RECT 144.850 73.270 352.480 73.670 ;
        RECT 96.195 70.035 96.595 71.235 ;
        RECT 120.925 70.835 121.925 70.885 ;
        RECT 120.925 70.435 143.995 70.835 ;
        RECT 120.925 70.385 121.925 70.435 ;
        RECT 95.075 66.675 95.475 67.875 ;
        RECT 94.575 56.255 94.855 65.695 ;
        RECT 95.135 56.535 95.415 66.675 ;
        RECT 95.695 56.255 95.975 65.695 ;
        RECT 96.255 56.535 96.535 70.035 ;
        RECT 144.850 69.910 334.560 70.310 ;
        RECT 97.315 66.675 97.715 67.875 ;
        RECT 120.925 67.475 121.925 67.525 ;
        RECT 120.925 67.075 143.995 67.475 ;
        RECT 120.925 67.025 121.925 67.075 ;
        RECT 96.815 56.255 97.095 65.695 ;
        RECT 97.375 56.535 97.655 66.675 ;
        RECT 98.495 66.285 100.455 66.685 ;
        RECT 144.850 66.550 316.640 66.950 ;
        RECT 97.935 56.255 98.215 65.695 ;
        RECT 98.495 56.695 98.775 66.285 ;
        RECT 99.055 56.255 99.335 65.695 ;
        RECT 99.615 56.695 99.895 66.285 ;
        RECT 100.175 56.255 100.455 66.285 ;
        RECT 120.925 64.115 121.925 64.165 ;
        RECT 120.925 63.715 143.995 64.115 ;
        RECT 120.925 63.665 121.925 63.715 ;
        RECT 298.160 63.590 298.720 65.000 ;
        RECT 144.850 63.190 298.720 63.590 ;
        RECT 298.160 61.000 298.720 63.190 ;
        RECT 316.080 61.000 316.640 66.550 ;
        RECT 334.000 61.000 334.560 69.910 ;
        RECT 335.260 61.140 337.220 61.420 ;
        RECT -477.745 56.095 100.455 56.255 ;
        RECT 298.300 56.380 298.580 61.000 ;
        RECT 298.300 56.100 300.820 56.380 ;
        RECT -483.245 55.595 125.505 56.095 ;
        RECT -477.745 55.435 100.455 55.595 ;
        RECT -477.745 45.405 -477.465 55.435 ;
        RECT -477.185 45.405 -476.905 54.995 ;
        RECT -476.625 45.995 -476.345 55.435 ;
        RECT -476.065 45.405 -475.785 54.995 ;
        RECT -475.505 45.995 -475.225 55.435 ;
        RECT -477.745 45.005 -475.785 45.405 ;
        RECT -474.945 45.015 -474.665 55.155 ;
        RECT -474.385 45.995 -474.105 55.435 ;
        RECT -475.005 43.815 -474.605 45.015 ;
        RECT -473.825 41.655 -473.545 55.155 ;
        RECT -473.265 45.995 -472.985 55.435 ;
        RECT -472.705 45.015 -472.425 55.155 ;
        RECT -472.145 45.995 -471.865 55.435 ;
        RECT -472.765 43.815 -472.365 45.015 ;
        RECT -473.885 40.455 -473.485 41.655 ;
        RECT -471.585 38.295 -471.305 55.155 ;
        RECT -471.025 45.995 -470.745 55.435 ;
        RECT -470.465 45.015 -470.185 55.155 ;
        RECT -469.905 45.995 -469.625 55.435 ;
        RECT -470.525 43.815 -470.125 45.015 ;
        RECT -469.345 41.655 -469.065 55.155 ;
        RECT -468.785 45.995 -468.505 55.435 ;
        RECT -468.225 45.015 -467.945 55.155 ;
        RECT -467.665 45.995 -467.385 55.435 ;
        RECT -468.285 43.815 -467.885 45.015 ;
        RECT -469.405 40.455 -469.005 41.655 ;
        RECT -471.645 37.095 -471.245 38.295 ;
        RECT -467.105 34.935 -466.825 55.155 ;
        RECT -466.545 45.995 -466.265 55.435 ;
        RECT -465.985 45.015 -465.705 55.155 ;
        RECT -465.425 45.995 -465.145 55.435 ;
        RECT -466.045 43.815 -465.645 45.015 ;
        RECT -464.865 41.655 -464.585 55.155 ;
        RECT -464.305 45.995 -464.025 55.435 ;
        RECT -463.745 45.015 -463.465 55.155 ;
        RECT -463.185 45.995 -462.905 55.435 ;
        RECT -463.805 43.815 -463.405 45.015 ;
        RECT -464.925 40.455 -464.525 41.655 ;
        RECT -462.625 38.295 -462.345 55.155 ;
        RECT -462.065 45.995 -461.785 55.435 ;
        RECT -461.505 45.015 -461.225 55.155 ;
        RECT -460.945 45.995 -460.665 55.435 ;
        RECT -461.565 43.815 -461.165 45.015 ;
        RECT -460.385 41.655 -460.105 55.155 ;
        RECT -459.825 45.995 -459.545 55.435 ;
        RECT -459.265 45.015 -458.985 55.155 ;
        RECT -458.705 45.995 -458.425 55.435 ;
        RECT -459.325 43.815 -458.925 45.015 ;
        RECT -460.445 40.455 -460.045 41.655 ;
        RECT -462.685 37.095 -462.285 38.295 ;
        RECT -467.165 33.735 -466.765 34.935 ;
        RECT -458.145 31.575 -457.865 55.155 ;
        RECT -457.585 45.995 -457.305 55.435 ;
        RECT -457.025 45.015 -456.745 55.155 ;
        RECT -456.465 45.995 -456.185 55.435 ;
        RECT -457.085 43.815 -456.685 45.015 ;
        RECT -455.905 41.655 -455.625 55.155 ;
        RECT -455.345 45.995 -455.065 55.435 ;
        RECT -454.785 45.015 -454.505 55.155 ;
        RECT -454.225 45.995 -453.945 55.435 ;
        RECT -454.845 43.815 -454.445 45.015 ;
        RECT -455.965 40.455 -455.565 41.655 ;
        RECT -453.665 38.295 -453.385 55.155 ;
        RECT -453.105 45.995 -452.825 55.435 ;
        RECT -452.545 45.015 -452.265 55.155 ;
        RECT -451.985 45.995 -451.705 55.435 ;
        RECT -452.605 43.815 -452.205 45.015 ;
        RECT -451.425 41.655 -451.145 55.155 ;
        RECT -450.865 45.995 -450.585 55.435 ;
        RECT -450.305 45.015 -450.025 55.155 ;
        RECT -449.745 45.995 -449.465 55.435 ;
        RECT -450.365 43.815 -449.965 45.015 ;
        RECT -451.485 40.455 -451.085 41.655 ;
        RECT -453.725 37.095 -453.325 38.295 ;
        RECT -449.185 34.935 -448.905 55.155 ;
        RECT -448.625 45.995 -448.345 55.435 ;
        RECT -448.065 45.015 -447.785 55.155 ;
        RECT -447.505 45.995 -447.225 55.435 ;
        RECT -448.125 43.815 -447.725 45.015 ;
        RECT -446.945 41.655 -446.665 55.155 ;
        RECT -446.385 45.995 -446.105 55.435 ;
        RECT -445.825 45.015 -445.545 55.155 ;
        RECT -445.265 45.995 -444.985 55.435 ;
        RECT -445.885 43.815 -445.485 45.015 ;
        RECT -447.005 40.455 -446.605 41.655 ;
        RECT -444.705 38.295 -444.425 55.155 ;
        RECT -444.145 45.995 -443.865 55.435 ;
        RECT -443.585 45.015 -443.305 55.155 ;
        RECT -443.025 45.995 -442.745 55.435 ;
        RECT -443.645 43.815 -443.245 45.015 ;
        RECT -442.465 41.655 -442.185 55.155 ;
        RECT -441.905 45.995 -441.625 55.435 ;
        RECT -441.345 45.015 -441.065 55.155 ;
        RECT -440.785 45.995 -440.505 55.435 ;
        RECT -441.405 43.815 -441.005 45.015 ;
        RECT -442.525 40.455 -442.125 41.655 ;
        RECT -444.765 37.095 -444.365 38.295 ;
        RECT -449.245 33.735 -448.845 34.935 ;
        RECT -458.205 30.375 -457.805 31.575 ;
        RECT -440.225 28.215 -439.945 55.155 ;
        RECT -439.665 45.995 -439.385 55.435 ;
        RECT -439.105 45.015 -438.825 55.155 ;
        RECT -438.545 45.995 -438.265 55.435 ;
        RECT -439.165 43.815 -438.765 45.015 ;
        RECT -437.985 41.655 -437.705 55.155 ;
        RECT -437.425 45.995 -437.145 55.435 ;
        RECT -436.865 45.015 -436.585 55.155 ;
        RECT -436.305 45.995 -436.025 55.435 ;
        RECT -436.925 43.815 -436.525 45.015 ;
        RECT -438.045 40.455 -437.645 41.655 ;
        RECT -435.745 38.295 -435.465 55.155 ;
        RECT -435.185 45.995 -434.905 55.435 ;
        RECT -434.625 45.015 -434.345 55.155 ;
        RECT -434.065 45.995 -433.785 55.435 ;
        RECT -434.685 43.815 -434.285 45.015 ;
        RECT -433.505 41.655 -433.225 55.155 ;
        RECT -432.945 45.995 -432.665 55.435 ;
        RECT -432.385 45.015 -432.105 55.155 ;
        RECT -431.825 45.995 -431.545 55.435 ;
        RECT -432.445 43.815 -432.045 45.015 ;
        RECT -433.565 40.455 -433.165 41.655 ;
        RECT -435.805 37.095 -435.405 38.295 ;
        RECT -431.265 34.935 -430.985 55.155 ;
        RECT -430.705 45.995 -430.425 55.435 ;
        RECT -430.145 45.015 -429.865 55.155 ;
        RECT -429.585 45.995 -429.305 55.435 ;
        RECT -430.205 43.815 -429.805 45.015 ;
        RECT -429.025 41.655 -428.745 55.155 ;
        RECT -428.465 45.995 -428.185 55.435 ;
        RECT -427.905 45.015 -427.625 55.155 ;
        RECT -427.345 45.995 -427.065 55.435 ;
        RECT -427.965 43.815 -427.565 45.015 ;
        RECT -429.085 40.455 -428.685 41.655 ;
        RECT -426.785 38.295 -426.505 55.155 ;
        RECT -426.225 45.995 -425.945 55.435 ;
        RECT -425.665 45.015 -425.385 55.155 ;
        RECT -425.105 45.995 -424.825 55.435 ;
        RECT -425.725 43.815 -425.325 45.015 ;
        RECT -424.545 41.655 -424.265 55.155 ;
        RECT -423.985 45.995 -423.705 55.435 ;
        RECT -423.425 45.015 -423.145 55.155 ;
        RECT -422.865 45.995 -422.585 55.435 ;
        RECT -423.485 43.815 -423.085 45.015 ;
        RECT -424.605 40.455 -424.205 41.655 ;
        RECT -426.845 37.095 -426.445 38.295 ;
        RECT -431.325 33.735 -430.925 34.935 ;
        RECT -422.305 31.575 -422.025 55.155 ;
        RECT -421.745 45.995 -421.465 55.435 ;
        RECT -421.185 45.015 -420.905 55.155 ;
        RECT -420.625 45.995 -420.345 55.435 ;
        RECT -421.245 43.815 -420.845 45.015 ;
        RECT -420.065 41.655 -419.785 55.155 ;
        RECT -419.505 45.995 -419.225 55.435 ;
        RECT -418.945 45.015 -418.665 55.155 ;
        RECT -418.385 45.995 -418.105 55.435 ;
        RECT -419.005 43.815 -418.605 45.015 ;
        RECT -420.125 40.455 -419.725 41.655 ;
        RECT -417.825 38.295 -417.545 55.155 ;
        RECT -417.265 45.995 -416.985 55.435 ;
        RECT -416.705 45.015 -416.425 55.155 ;
        RECT -416.145 45.995 -415.865 55.435 ;
        RECT -416.765 43.815 -416.365 45.015 ;
        RECT -415.585 41.655 -415.305 55.155 ;
        RECT -415.025 45.995 -414.745 55.435 ;
        RECT -414.465 45.015 -414.185 55.155 ;
        RECT -413.905 45.995 -413.625 55.435 ;
        RECT -414.525 43.815 -414.125 45.015 ;
        RECT -415.645 40.455 -415.245 41.655 ;
        RECT -417.885 37.095 -417.485 38.295 ;
        RECT -413.345 34.935 -413.065 55.155 ;
        RECT -412.785 45.995 -412.505 55.435 ;
        RECT -412.225 45.015 -411.945 55.155 ;
        RECT -411.665 45.995 -411.385 55.435 ;
        RECT -412.285 43.815 -411.885 45.015 ;
        RECT -411.105 41.655 -410.825 55.155 ;
        RECT -410.545 45.995 -410.265 55.435 ;
        RECT -409.985 45.015 -409.705 55.155 ;
        RECT -409.425 45.995 -409.145 55.435 ;
        RECT -410.045 43.815 -409.645 45.015 ;
        RECT -411.165 40.455 -410.765 41.655 ;
        RECT -408.865 38.295 -408.585 55.155 ;
        RECT -408.305 45.995 -408.025 55.435 ;
        RECT -407.745 45.015 -407.465 55.155 ;
        RECT -407.185 45.995 -406.905 55.435 ;
        RECT -407.805 43.815 -407.405 45.015 ;
        RECT -406.625 41.655 -406.345 55.155 ;
        RECT -406.065 45.995 -405.785 55.435 ;
        RECT -405.505 45.015 -405.225 55.155 ;
        RECT -404.945 45.995 -404.665 55.435 ;
        RECT -405.565 43.815 -405.165 45.015 ;
        RECT -406.685 40.455 -406.285 41.655 ;
        RECT -408.925 37.095 -408.525 38.295 ;
        RECT -413.405 33.735 -413.005 34.935 ;
        RECT -422.365 30.375 -421.965 31.575 ;
        RECT -440.285 27.015 -439.885 28.215 ;
        RECT -404.385 24.855 -404.105 55.155 ;
        RECT -403.825 45.995 -403.545 55.435 ;
        RECT -403.265 45.015 -402.985 55.155 ;
        RECT -402.705 45.995 -402.425 55.435 ;
        RECT -403.325 43.815 -402.925 45.015 ;
        RECT -402.145 41.655 -401.865 55.155 ;
        RECT -401.585 45.995 -401.305 55.435 ;
        RECT -401.025 45.015 -400.745 55.155 ;
        RECT -400.465 45.995 -400.185 55.435 ;
        RECT -401.085 43.815 -400.685 45.015 ;
        RECT -402.205 40.455 -401.805 41.655 ;
        RECT -399.905 38.295 -399.625 55.155 ;
        RECT -399.345 45.995 -399.065 55.435 ;
        RECT -398.785 45.015 -398.505 55.155 ;
        RECT -398.225 45.995 -397.945 55.435 ;
        RECT -398.845 43.815 -398.445 45.015 ;
        RECT -397.665 41.655 -397.385 55.155 ;
        RECT -397.105 45.995 -396.825 55.435 ;
        RECT -396.545 45.015 -396.265 55.155 ;
        RECT -395.985 45.995 -395.705 55.435 ;
        RECT -396.605 43.815 -396.205 45.015 ;
        RECT -397.725 40.455 -397.325 41.655 ;
        RECT -399.965 37.095 -399.565 38.295 ;
        RECT -395.425 34.935 -395.145 55.155 ;
        RECT -394.865 45.995 -394.585 55.435 ;
        RECT -394.305 45.015 -394.025 55.155 ;
        RECT -393.745 45.995 -393.465 55.435 ;
        RECT -394.365 43.815 -393.965 45.015 ;
        RECT -393.185 41.655 -392.905 55.155 ;
        RECT -392.625 45.995 -392.345 55.435 ;
        RECT -392.065 45.015 -391.785 55.155 ;
        RECT -391.505 45.995 -391.225 55.435 ;
        RECT -392.125 43.815 -391.725 45.015 ;
        RECT -393.245 40.455 -392.845 41.655 ;
        RECT -390.945 38.295 -390.665 55.155 ;
        RECT -390.385 45.995 -390.105 55.435 ;
        RECT -389.825 45.015 -389.545 55.155 ;
        RECT -389.265 45.995 -388.985 55.435 ;
        RECT -389.885 43.815 -389.485 45.015 ;
        RECT -388.705 41.655 -388.425 55.155 ;
        RECT -388.145 45.995 -387.865 55.435 ;
        RECT -387.585 45.015 -387.305 55.155 ;
        RECT -387.025 45.995 -386.745 55.435 ;
        RECT -387.645 43.815 -387.245 45.015 ;
        RECT -388.765 40.455 -388.365 41.655 ;
        RECT -391.005 37.095 -390.605 38.295 ;
        RECT -395.485 33.735 -395.085 34.935 ;
        RECT -386.465 31.575 -386.185 55.155 ;
        RECT -385.905 45.995 -385.625 55.435 ;
        RECT -385.345 45.015 -385.065 55.155 ;
        RECT -384.785 45.995 -384.505 55.435 ;
        RECT -385.405 43.815 -385.005 45.015 ;
        RECT -384.225 41.655 -383.945 55.155 ;
        RECT -383.665 45.995 -383.385 55.435 ;
        RECT -383.105 45.015 -382.825 55.155 ;
        RECT -382.545 45.995 -382.265 55.435 ;
        RECT -383.165 43.815 -382.765 45.015 ;
        RECT -384.285 40.455 -383.885 41.655 ;
        RECT -381.985 38.295 -381.705 55.155 ;
        RECT -381.425 45.995 -381.145 55.435 ;
        RECT -380.865 45.015 -380.585 55.155 ;
        RECT -380.305 45.995 -380.025 55.435 ;
        RECT -380.925 43.815 -380.525 45.015 ;
        RECT -379.745 41.655 -379.465 55.155 ;
        RECT -379.185 45.995 -378.905 55.435 ;
        RECT -378.625 45.015 -378.345 55.155 ;
        RECT -378.065 45.995 -377.785 55.435 ;
        RECT -378.685 43.815 -378.285 45.015 ;
        RECT -379.805 40.455 -379.405 41.655 ;
        RECT -382.045 37.095 -381.645 38.295 ;
        RECT -377.505 34.935 -377.225 55.155 ;
        RECT -376.945 45.995 -376.665 55.435 ;
        RECT -376.385 45.015 -376.105 55.155 ;
        RECT -375.825 45.995 -375.545 55.435 ;
        RECT -376.445 43.815 -376.045 45.015 ;
        RECT -375.265 41.655 -374.985 55.155 ;
        RECT -374.705 45.995 -374.425 55.435 ;
        RECT -374.145 45.015 -373.865 55.155 ;
        RECT -373.585 45.995 -373.305 55.435 ;
        RECT -374.205 43.815 -373.805 45.015 ;
        RECT -375.325 40.455 -374.925 41.655 ;
        RECT -373.025 38.295 -372.745 55.155 ;
        RECT -372.465 45.995 -372.185 55.435 ;
        RECT -371.905 45.015 -371.625 55.155 ;
        RECT -371.345 45.995 -371.065 55.435 ;
        RECT -371.965 43.815 -371.565 45.015 ;
        RECT -370.785 41.655 -370.505 55.155 ;
        RECT -370.225 45.995 -369.945 55.435 ;
        RECT -369.665 45.015 -369.385 55.155 ;
        RECT -369.105 45.995 -368.825 55.435 ;
        RECT -369.725 43.815 -369.325 45.015 ;
        RECT -370.845 40.455 -370.445 41.655 ;
        RECT -373.085 37.095 -372.685 38.295 ;
        RECT -377.565 33.735 -377.165 34.935 ;
        RECT -386.525 30.375 -386.125 31.575 ;
        RECT -368.545 28.215 -368.265 55.155 ;
        RECT -367.985 45.995 -367.705 55.435 ;
        RECT -367.425 45.015 -367.145 55.155 ;
        RECT -366.865 45.995 -366.585 55.435 ;
        RECT -367.485 43.815 -367.085 45.015 ;
        RECT -366.305 41.655 -366.025 55.155 ;
        RECT -365.745 45.995 -365.465 55.435 ;
        RECT -365.185 45.015 -364.905 55.155 ;
        RECT -364.625 45.995 -364.345 55.435 ;
        RECT -365.245 43.815 -364.845 45.015 ;
        RECT -366.365 40.455 -365.965 41.655 ;
        RECT -364.065 38.295 -363.785 55.155 ;
        RECT -363.505 45.995 -363.225 55.435 ;
        RECT -362.945 45.015 -362.665 55.155 ;
        RECT -362.385 45.995 -362.105 55.435 ;
        RECT -363.005 43.815 -362.605 45.015 ;
        RECT -361.825 41.655 -361.545 55.155 ;
        RECT -361.265 45.995 -360.985 55.435 ;
        RECT -360.705 45.015 -360.425 55.155 ;
        RECT -360.145 45.995 -359.865 55.435 ;
        RECT -360.765 43.815 -360.365 45.015 ;
        RECT -361.885 40.455 -361.485 41.655 ;
        RECT -364.125 37.095 -363.725 38.295 ;
        RECT -359.585 34.935 -359.305 55.155 ;
        RECT -359.025 45.995 -358.745 55.435 ;
        RECT -358.465 45.015 -358.185 55.155 ;
        RECT -357.905 45.995 -357.625 55.435 ;
        RECT -358.525 43.815 -358.125 45.015 ;
        RECT -357.345 41.655 -357.065 55.155 ;
        RECT -356.785 45.995 -356.505 55.435 ;
        RECT -356.225 45.015 -355.945 55.155 ;
        RECT -355.665 45.995 -355.385 55.435 ;
        RECT -356.285 43.815 -355.885 45.015 ;
        RECT -357.405 40.455 -357.005 41.655 ;
        RECT -355.105 38.295 -354.825 55.155 ;
        RECT -354.545 45.995 -354.265 55.435 ;
        RECT -353.985 45.015 -353.705 55.155 ;
        RECT -353.425 45.995 -353.145 55.435 ;
        RECT -354.045 43.815 -353.645 45.015 ;
        RECT -352.865 41.655 -352.585 55.155 ;
        RECT -352.305 45.995 -352.025 55.435 ;
        RECT -351.745 45.015 -351.465 55.155 ;
        RECT -351.185 45.995 -350.905 55.435 ;
        RECT -351.805 43.815 -351.405 45.015 ;
        RECT -352.925 40.455 -352.525 41.655 ;
        RECT -355.165 37.095 -354.765 38.295 ;
        RECT -359.645 33.735 -359.245 34.935 ;
        RECT -350.625 31.575 -350.345 55.155 ;
        RECT -350.065 45.995 -349.785 55.435 ;
        RECT -349.505 45.015 -349.225 55.155 ;
        RECT -348.945 45.995 -348.665 55.435 ;
        RECT -349.565 43.815 -349.165 45.015 ;
        RECT -348.385 41.655 -348.105 55.155 ;
        RECT -347.825 45.995 -347.545 55.435 ;
        RECT -347.265 45.015 -346.985 55.155 ;
        RECT -346.705 45.995 -346.425 55.435 ;
        RECT -347.325 43.815 -346.925 45.015 ;
        RECT -348.445 40.455 -348.045 41.655 ;
        RECT -346.145 38.295 -345.865 55.155 ;
        RECT -345.585 45.995 -345.305 55.435 ;
        RECT -345.025 45.015 -344.745 55.155 ;
        RECT -344.465 45.995 -344.185 55.435 ;
        RECT -345.085 43.815 -344.685 45.015 ;
        RECT -343.905 41.655 -343.625 55.155 ;
        RECT -343.345 45.995 -343.065 55.435 ;
        RECT -342.785 45.015 -342.505 55.155 ;
        RECT -342.225 45.995 -341.945 55.435 ;
        RECT -342.845 43.815 -342.445 45.015 ;
        RECT -343.965 40.455 -343.565 41.655 ;
        RECT -346.205 37.095 -345.805 38.295 ;
        RECT -341.665 34.935 -341.385 55.155 ;
        RECT -341.105 45.995 -340.825 55.435 ;
        RECT -340.545 45.015 -340.265 55.155 ;
        RECT -339.985 45.995 -339.705 55.435 ;
        RECT -340.605 43.815 -340.205 45.015 ;
        RECT -339.425 41.655 -339.145 55.155 ;
        RECT -338.865 45.995 -338.585 55.435 ;
        RECT -338.305 45.015 -338.025 55.155 ;
        RECT -337.745 45.995 -337.465 55.435 ;
        RECT -338.365 43.815 -337.965 45.015 ;
        RECT -339.485 40.455 -339.085 41.655 ;
        RECT -337.185 38.295 -336.905 55.155 ;
        RECT -336.625 45.995 -336.345 55.435 ;
        RECT -336.065 45.015 -335.785 55.155 ;
        RECT -335.505 45.995 -335.225 55.435 ;
        RECT -336.125 43.815 -335.725 45.015 ;
        RECT -334.945 41.655 -334.665 55.155 ;
        RECT -334.385 45.995 -334.105 55.435 ;
        RECT -333.825 45.015 -333.545 55.155 ;
        RECT -333.265 45.995 -332.985 55.435 ;
        RECT -333.885 43.815 -333.485 45.015 ;
        RECT -335.005 40.455 -334.605 41.655 ;
        RECT -337.245 37.095 -336.845 38.295 ;
        RECT -341.725 33.735 -341.325 34.935 ;
        RECT -350.685 30.375 -350.285 31.575 ;
        RECT -368.605 27.015 -368.205 28.215 ;
        RECT -404.445 23.655 -404.045 24.855 ;
        RECT -332.705 21.495 -332.425 55.155 ;
        RECT -332.145 45.995 -331.865 55.435 ;
        RECT -331.585 45.015 -331.305 55.155 ;
        RECT -331.025 45.995 -330.745 55.435 ;
        RECT -331.645 43.815 -331.245 45.015 ;
        RECT -330.465 41.655 -330.185 55.155 ;
        RECT -329.905 45.995 -329.625 55.435 ;
        RECT -329.345 45.015 -329.065 55.155 ;
        RECT -328.785 45.995 -328.505 55.435 ;
        RECT -329.405 43.815 -329.005 45.015 ;
        RECT -330.525 40.455 -330.125 41.655 ;
        RECT -328.225 38.295 -327.945 55.155 ;
        RECT -327.665 45.995 -327.385 55.435 ;
        RECT -327.105 45.015 -326.825 55.155 ;
        RECT -326.545 45.995 -326.265 55.435 ;
        RECT -327.165 43.815 -326.765 45.015 ;
        RECT -325.985 41.655 -325.705 55.155 ;
        RECT -325.425 45.995 -325.145 55.435 ;
        RECT -324.865 45.015 -324.585 55.155 ;
        RECT -324.305 45.995 -324.025 55.435 ;
        RECT -324.925 43.815 -324.525 45.015 ;
        RECT -326.045 40.455 -325.645 41.655 ;
        RECT -328.285 37.095 -327.885 38.295 ;
        RECT -323.745 34.935 -323.465 55.155 ;
        RECT -323.185 45.995 -322.905 55.435 ;
        RECT -322.625 45.015 -322.345 55.155 ;
        RECT -322.065 45.995 -321.785 55.435 ;
        RECT -322.685 43.815 -322.285 45.015 ;
        RECT -321.505 41.655 -321.225 55.155 ;
        RECT -320.945 45.995 -320.665 55.435 ;
        RECT -320.385 45.015 -320.105 55.155 ;
        RECT -319.825 45.995 -319.545 55.435 ;
        RECT -320.445 43.815 -320.045 45.015 ;
        RECT -321.565 40.455 -321.165 41.655 ;
        RECT -319.265 38.295 -318.985 55.155 ;
        RECT -318.705 45.995 -318.425 55.435 ;
        RECT -318.145 45.015 -317.865 55.155 ;
        RECT -317.585 45.995 -317.305 55.435 ;
        RECT -318.205 43.815 -317.805 45.015 ;
        RECT -317.025 41.655 -316.745 55.155 ;
        RECT -316.465 45.995 -316.185 55.435 ;
        RECT -315.905 45.015 -315.625 55.155 ;
        RECT -315.345 45.995 -315.065 55.435 ;
        RECT -315.965 43.815 -315.565 45.015 ;
        RECT -317.085 40.455 -316.685 41.655 ;
        RECT -319.325 37.095 -318.925 38.295 ;
        RECT -323.805 33.735 -323.405 34.935 ;
        RECT -314.785 31.575 -314.505 55.155 ;
        RECT -314.225 45.995 -313.945 55.435 ;
        RECT -313.665 45.015 -313.385 55.155 ;
        RECT -313.105 45.995 -312.825 55.435 ;
        RECT -313.725 43.815 -313.325 45.015 ;
        RECT -312.545 41.655 -312.265 55.155 ;
        RECT -311.985 45.995 -311.705 55.435 ;
        RECT -311.425 45.015 -311.145 55.155 ;
        RECT -310.865 45.995 -310.585 55.435 ;
        RECT -311.485 43.815 -311.085 45.015 ;
        RECT -312.605 40.455 -312.205 41.655 ;
        RECT -310.305 38.295 -310.025 55.155 ;
        RECT -309.745 45.995 -309.465 55.435 ;
        RECT -309.185 45.015 -308.905 55.155 ;
        RECT -308.625 45.995 -308.345 55.435 ;
        RECT -309.245 43.815 -308.845 45.015 ;
        RECT -308.065 41.655 -307.785 55.155 ;
        RECT -307.505 45.995 -307.225 55.435 ;
        RECT -306.945 45.015 -306.665 55.155 ;
        RECT -306.385 45.995 -306.105 55.435 ;
        RECT -307.005 43.815 -306.605 45.015 ;
        RECT -308.125 40.455 -307.725 41.655 ;
        RECT -310.365 37.095 -309.965 38.295 ;
        RECT -305.825 34.935 -305.545 55.155 ;
        RECT -305.265 45.995 -304.985 55.435 ;
        RECT -304.705 45.015 -304.425 55.155 ;
        RECT -304.145 45.995 -303.865 55.435 ;
        RECT -304.765 43.815 -304.365 45.015 ;
        RECT -303.585 41.655 -303.305 55.155 ;
        RECT -303.025 45.995 -302.745 55.435 ;
        RECT -302.465 45.015 -302.185 55.155 ;
        RECT -301.905 45.995 -301.625 55.435 ;
        RECT -302.525 43.815 -302.125 45.015 ;
        RECT -303.645 40.455 -303.245 41.655 ;
        RECT -301.345 38.295 -301.065 55.155 ;
        RECT -300.785 45.995 -300.505 55.435 ;
        RECT -300.225 45.015 -299.945 55.155 ;
        RECT -299.665 45.995 -299.385 55.435 ;
        RECT -300.285 43.815 -299.885 45.015 ;
        RECT -299.105 41.655 -298.825 55.155 ;
        RECT -298.545 45.995 -298.265 55.435 ;
        RECT -297.985 45.015 -297.705 55.155 ;
        RECT -297.425 45.995 -297.145 55.435 ;
        RECT -298.045 43.815 -297.645 45.015 ;
        RECT -299.165 40.455 -298.765 41.655 ;
        RECT -301.405 37.095 -301.005 38.295 ;
        RECT -305.885 33.735 -305.485 34.935 ;
        RECT -314.845 30.375 -314.445 31.575 ;
        RECT -296.865 28.215 -296.585 55.155 ;
        RECT -296.305 45.995 -296.025 55.435 ;
        RECT -295.745 45.015 -295.465 55.155 ;
        RECT -295.185 45.995 -294.905 55.435 ;
        RECT -295.805 43.815 -295.405 45.015 ;
        RECT -294.625 41.655 -294.345 55.155 ;
        RECT -294.065 45.995 -293.785 55.435 ;
        RECT -293.505 45.015 -293.225 55.155 ;
        RECT -292.945 45.995 -292.665 55.435 ;
        RECT -293.565 43.815 -293.165 45.015 ;
        RECT -294.685 40.455 -294.285 41.655 ;
        RECT -292.385 38.295 -292.105 55.155 ;
        RECT -291.825 45.995 -291.545 55.435 ;
        RECT -291.265 45.015 -290.985 55.155 ;
        RECT -290.705 45.995 -290.425 55.435 ;
        RECT -291.325 43.815 -290.925 45.015 ;
        RECT -290.145 41.655 -289.865 55.155 ;
        RECT -289.585 45.995 -289.305 55.435 ;
        RECT -289.025 45.015 -288.745 55.155 ;
        RECT -288.465 45.995 -288.185 55.435 ;
        RECT -289.085 43.815 -288.685 45.015 ;
        RECT -290.205 40.455 -289.805 41.655 ;
        RECT -292.445 37.095 -292.045 38.295 ;
        RECT -287.905 34.935 -287.625 55.155 ;
        RECT -287.345 45.995 -287.065 55.435 ;
        RECT -286.785 45.015 -286.505 55.155 ;
        RECT -286.225 45.995 -285.945 55.435 ;
        RECT -286.845 43.815 -286.445 45.015 ;
        RECT -285.665 41.655 -285.385 55.155 ;
        RECT -285.105 45.995 -284.825 55.435 ;
        RECT -284.545 45.015 -284.265 55.155 ;
        RECT -283.985 45.995 -283.705 55.435 ;
        RECT -284.605 43.815 -284.205 45.015 ;
        RECT -285.725 40.455 -285.325 41.655 ;
        RECT -283.425 38.295 -283.145 55.155 ;
        RECT -282.865 45.995 -282.585 55.435 ;
        RECT -282.305 45.015 -282.025 55.155 ;
        RECT -281.745 45.995 -281.465 55.435 ;
        RECT -282.365 43.815 -281.965 45.015 ;
        RECT -281.185 41.655 -280.905 55.155 ;
        RECT -280.625 45.995 -280.345 55.435 ;
        RECT -280.065 45.015 -279.785 55.155 ;
        RECT -279.505 45.995 -279.225 55.435 ;
        RECT -280.125 43.815 -279.725 45.015 ;
        RECT -281.245 40.455 -280.845 41.655 ;
        RECT -283.485 37.095 -283.085 38.295 ;
        RECT -287.965 33.735 -287.565 34.935 ;
        RECT -278.945 31.575 -278.665 55.155 ;
        RECT -278.385 45.995 -278.105 55.435 ;
        RECT -277.825 45.015 -277.545 55.155 ;
        RECT -277.265 45.995 -276.985 55.435 ;
        RECT -277.885 43.815 -277.485 45.015 ;
        RECT -276.705 41.655 -276.425 55.155 ;
        RECT -276.145 45.995 -275.865 55.435 ;
        RECT -275.585 45.015 -275.305 55.155 ;
        RECT -275.025 45.995 -274.745 55.435 ;
        RECT -275.645 43.815 -275.245 45.015 ;
        RECT -276.765 40.455 -276.365 41.655 ;
        RECT -274.465 38.295 -274.185 55.155 ;
        RECT -273.905 45.995 -273.625 55.435 ;
        RECT -273.345 45.015 -273.065 55.155 ;
        RECT -272.785 45.995 -272.505 55.435 ;
        RECT -273.405 43.815 -273.005 45.015 ;
        RECT -272.225 41.655 -271.945 55.155 ;
        RECT -271.665 45.995 -271.385 55.435 ;
        RECT -271.105 45.015 -270.825 55.155 ;
        RECT -270.545 45.995 -270.265 55.435 ;
        RECT -271.165 43.815 -270.765 45.015 ;
        RECT -272.285 40.455 -271.885 41.655 ;
        RECT -274.525 37.095 -274.125 38.295 ;
        RECT -269.985 34.935 -269.705 55.155 ;
        RECT -269.425 45.995 -269.145 55.435 ;
        RECT -268.865 45.015 -268.585 55.155 ;
        RECT -268.305 45.995 -268.025 55.435 ;
        RECT -268.925 43.815 -268.525 45.015 ;
        RECT -267.745 41.655 -267.465 55.155 ;
        RECT -267.185 45.995 -266.905 55.435 ;
        RECT -266.625 45.015 -266.345 55.155 ;
        RECT -266.065 45.995 -265.785 55.435 ;
        RECT -266.685 43.815 -266.285 45.015 ;
        RECT -267.805 40.455 -267.405 41.655 ;
        RECT -265.505 38.295 -265.225 55.155 ;
        RECT -264.945 45.995 -264.665 55.435 ;
        RECT -264.385 45.015 -264.105 55.155 ;
        RECT -263.825 45.995 -263.545 55.435 ;
        RECT -264.445 43.815 -264.045 45.015 ;
        RECT -263.265 41.655 -262.985 55.155 ;
        RECT -262.705 45.995 -262.425 55.435 ;
        RECT -262.145 45.015 -261.865 55.155 ;
        RECT -261.585 45.995 -261.305 55.435 ;
        RECT -262.205 43.815 -261.805 45.015 ;
        RECT -263.325 40.455 -262.925 41.655 ;
        RECT -265.565 37.095 -265.165 38.295 ;
        RECT -270.045 33.735 -269.645 34.935 ;
        RECT -279.005 30.375 -278.605 31.575 ;
        RECT -296.925 27.015 -296.525 28.215 ;
        RECT -261.025 24.855 -260.745 55.155 ;
        RECT -260.465 45.995 -260.185 55.435 ;
        RECT -259.905 45.015 -259.625 55.155 ;
        RECT -259.345 45.995 -259.065 55.435 ;
        RECT -259.965 43.815 -259.565 45.015 ;
        RECT -258.785 41.655 -258.505 55.155 ;
        RECT -258.225 45.995 -257.945 55.435 ;
        RECT -257.665 45.015 -257.385 55.155 ;
        RECT -257.105 45.995 -256.825 55.435 ;
        RECT -257.725 43.815 -257.325 45.015 ;
        RECT -258.845 40.455 -258.445 41.655 ;
        RECT -256.545 38.295 -256.265 55.155 ;
        RECT -255.985 45.995 -255.705 55.435 ;
        RECT -255.425 45.015 -255.145 55.155 ;
        RECT -254.865 45.995 -254.585 55.435 ;
        RECT -255.485 43.815 -255.085 45.015 ;
        RECT -254.305 41.655 -254.025 55.155 ;
        RECT -253.745 45.995 -253.465 55.435 ;
        RECT -253.185 45.015 -252.905 55.155 ;
        RECT -252.625 45.995 -252.345 55.435 ;
        RECT -253.245 43.815 -252.845 45.015 ;
        RECT -254.365 40.455 -253.965 41.655 ;
        RECT -256.605 37.095 -256.205 38.295 ;
        RECT -252.065 34.935 -251.785 55.155 ;
        RECT -251.505 45.995 -251.225 55.435 ;
        RECT -250.945 45.015 -250.665 55.155 ;
        RECT -250.385 45.995 -250.105 55.435 ;
        RECT -251.005 43.815 -250.605 45.015 ;
        RECT -249.825 41.655 -249.545 55.155 ;
        RECT -249.265 45.995 -248.985 55.435 ;
        RECT -248.705 45.015 -248.425 55.155 ;
        RECT -248.145 45.995 -247.865 55.435 ;
        RECT -248.765 43.815 -248.365 45.015 ;
        RECT -249.885 40.455 -249.485 41.655 ;
        RECT -247.585 38.295 -247.305 55.155 ;
        RECT -247.025 45.995 -246.745 55.435 ;
        RECT -246.465 45.015 -246.185 55.155 ;
        RECT -245.905 45.995 -245.625 55.435 ;
        RECT -246.525 43.815 -246.125 45.015 ;
        RECT -245.345 41.655 -245.065 55.155 ;
        RECT -244.785 45.995 -244.505 55.435 ;
        RECT -244.225 45.015 -243.945 55.155 ;
        RECT -243.665 45.995 -243.385 55.435 ;
        RECT -244.285 43.815 -243.885 45.015 ;
        RECT -245.405 40.455 -245.005 41.655 ;
        RECT -247.645 37.095 -247.245 38.295 ;
        RECT -252.125 33.735 -251.725 34.935 ;
        RECT -243.105 31.575 -242.825 55.155 ;
        RECT -242.545 45.995 -242.265 55.435 ;
        RECT -241.985 45.015 -241.705 55.155 ;
        RECT -241.425 45.995 -241.145 55.435 ;
        RECT -242.045 43.815 -241.645 45.015 ;
        RECT -240.865 41.655 -240.585 55.155 ;
        RECT -240.305 45.995 -240.025 55.435 ;
        RECT -239.745 45.015 -239.465 55.155 ;
        RECT -239.185 45.995 -238.905 55.435 ;
        RECT -239.805 43.815 -239.405 45.015 ;
        RECT -240.925 40.455 -240.525 41.655 ;
        RECT -238.625 38.295 -238.345 55.155 ;
        RECT -238.065 45.995 -237.785 55.435 ;
        RECT -237.505 45.015 -237.225 55.155 ;
        RECT -236.945 45.995 -236.665 55.435 ;
        RECT -237.565 43.815 -237.165 45.015 ;
        RECT -236.385 41.655 -236.105 55.155 ;
        RECT -235.825 45.995 -235.545 55.435 ;
        RECT -235.265 45.015 -234.985 55.155 ;
        RECT -234.705 45.995 -234.425 55.435 ;
        RECT -235.325 43.815 -234.925 45.015 ;
        RECT -236.445 40.455 -236.045 41.655 ;
        RECT -238.685 37.095 -238.285 38.295 ;
        RECT -234.145 34.935 -233.865 55.155 ;
        RECT -233.585 45.995 -233.305 55.435 ;
        RECT -233.025 45.015 -232.745 55.155 ;
        RECT -232.465 45.995 -232.185 55.435 ;
        RECT -233.085 43.815 -232.685 45.015 ;
        RECT -231.905 41.655 -231.625 55.155 ;
        RECT -231.345 45.995 -231.065 55.435 ;
        RECT -230.785 45.015 -230.505 55.155 ;
        RECT -230.225 45.995 -229.945 55.435 ;
        RECT -230.845 43.815 -230.445 45.015 ;
        RECT -231.965 40.455 -231.565 41.655 ;
        RECT -229.665 38.295 -229.385 55.155 ;
        RECT -229.105 45.995 -228.825 55.435 ;
        RECT -228.545 45.015 -228.265 55.155 ;
        RECT -227.985 45.995 -227.705 55.435 ;
        RECT -228.605 43.815 -228.205 45.015 ;
        RECT -227.425 41.655 -227.145 55.155 ;
        RECT -226.865 45.995 -226.585 55.435 ;
        RECT -226.305 45.015 -226.025 55.155 ;
        RECT -225.745 45.995 -225.465 55.435 ;
        RECT -226.365 43.815 -225.965 45.015 ;
        RECT -227.485 40.455 -227.085 41.655 ;
        RECT -229.725 37.095 -229.325 38.295 ;
        RECT -234.205 33.735 -233.805 34.935 ;
        RECT -243.165 30.375 -242.765 31.575 ;
        RECT -225.185 28.215 -224.905 55.155 ;
        RECT -224.625 45.995 -224.345 55.435 ;
        RECT -224.065 45.015 -223.785 55.155 ;
        RECT -223.505 45.995 -223.225 55.435 ;
        RECT -224.125 43.815 -223.725 45.015 ;
        RECT -222.945 41.655 -222.665 55.155 ;
        RECT -222.385 45.995 -222.105 55.435 ;
        RECT -221.825 45.015 -221.545 55.155 ;
        RECT -221.265 45.995 -220.985 55.435 ;
        RECT -221.885 43.815 -221.485 45.015 ;
        RECT -223.005 40.455 -222.605 41.655 ;
        RECT -220.705 38.295 -220.425 55.155 ;
        RECT -220.145 45.995 -219.865 55.435 ;
        RECT -219.585 45.015 -219.305 55.155 ;
        RECT -219.025 45.995 -218.745 55.435 ;
        RECT -219.645 43.815 -219.245 45.015 ;
        RECT -218.465 41.655 -218.185 55.155 ;
        RECT -217.905 45.995 -217.625 55.435 ;
        RECT -217.345 45.015 -217.065 55.155 ;
        RECT -216.785 45.995 -216.505 55.435 ;
        RECT -217.405 43.815 -217.005 45.015 ;
        RECT -218.525 40.455 -218.125 41.655 ;
        RECT -220.765 37.095 -220.365 38.295 ;
        RECT -216.225 34.935 -215.945 55.155 ;
        RECT -215.665 45.995 -215.385 55.435 ;
        RECT -215.105 45.015 -214.825 55.155 ;
        RECT -214.545 45.995 -214.265 55.435 ;
        RECT -215.165 43.815 -214.765 45.015 ;
        RECT -213.985 41.655 -213.705 55.155 ;
        RECT -213.425 45.995 -213.145 55.435 ;
        RECT -212.865 45.015 -212.585 55.155 ;
        RECT -212.305 45.995 -212.025 55.435 ;
        RECT -212.925 43.815 -212.525 45.015 ;
        RECT -214.045 40.455 -213.645 41.655 ;
        RECT -211.745 38.295 -211.465 55.155 ;
        RECT -211.185 45.995 -210.905 55.435 ;
        RECT -210.625 45.015 -210.345 55.155 ;
        RECT -210.065 45.995 -209.785 55.435 ;
        RECT -210.685 43.815 -210.285 45.015 ;
        RECT -209.505 41.655 -209.225 55.155 ;
        RECT -208.945 45.995 -208.665 55.435 ;
        RECT -208.385 45.015 -208.105 55.155 ;
        RECT -207.825 45.995 -207.545 55.435 ;
        RECT -208.445 43.815 -208.045 45.015 ;
        RECT -209.565 40.455 -209.165 41.655 ;
        RECT -211.805 37.095 -211.405 38.295 ;
        RECT -216.285 33.735 -215.885 34.935 ;
        RECT -207.265 31.575 -206.985 55.155 ;
        RECT -206.705 45.995 -206.425 55.435 ;
        RECT -206.145 45.015 -205.865 55.155 ;
        RECT -205.585 45.995 -205.305 55.435 ;
        RECT -206.205 43.815 -205.805 45.015 ;
        RECT -205.025 41.655 -204.745 55.155 ;
        RECT -204.465 45.995 -204.185 55.435 ;
        RECT -203.905 45.015 -203.625 55.155 ;
        RECT -203.345 45.995 -203.065 55.435 ;
        RECT -203.965 43.815 -203.565 45.015 ;
        RECT -205.085 40.455 -204.685 41.655 ;
        RECT -202.785 38.295 -202.505 55.155 ;
        RECT -202.225 45.995 -201.945 55.435 ;
        RECT -201.665 45.015 -201.385 55.155 ;
        RECT -201.105 45.995 -200.825 55.435 ;
        RECT -201.725 43.815 -201.325 45.015 ;
        RECT -200.545 41.655 -200.265 55.155 ;
        RECT -199.985 45.995 -199.705 55.435 ;
        RECT -199.425 45.015 -199.145 55.155 ;
        RECT -198.865 45.995 -198.585 55.435 ;
        RECT -199.485 43.815 -199.085 45.015 ;
        RECT -200.605 40.455 -200.205 41.655 ;
        RECT -202.845 37.095 -202.445 38.295 ;
        RECT -198.305 34.935 -198.025 55.155 ;
        RECT -197.745 45.995 -197.465 55.435 ;
        RECT -197.185 45.015 -196.905 55.155 ;
        RECT -196.625 45.995 -196.345 55.435 ;
        RECT -197.245 43.815 -196.845 45.015 ;
        RECT -196.065 41.655 -195.785 55.155 ;
        RECT -195.505 45.995 -195.225 55.435 ;
        RECT -194.945 45.015 -194.665 55.155 ;
        RECT -194.385 45.995 -194.105 55.435 ;
        RECT -195.005 43.815 -194.605 45.015 ;
        RECT -196.125 40.455 -195.725 41.655 ;
        RECT -193.825 38.295 -193.545 55.155 ;
        RECT -193.265 45.995 -192.985 55.435 ;
        RECT -192.705 45.015 -192.425 55.155 ;
        RECT -192.145 45.995 -191.865 55.435 ;
        RECT -192.765 43.815 -192.365 45.015 ;
        RECT -191.585 41.655 -191.305 55.155 ;
        RECT -191.025 45.995 -190.745 55.435 ;
        RECT -190.465 45.015 -190.185 55.155 ;
        RECT -189.905 45.995 -189.625 55.435 ;
        RECT -190.525 43.815 -190.125 45.015 ;
        RECT -191.645 40.455 -191.245 41.655 ;
        RECT -193.885 37.095 -193.485 38.295 ;
        RECT -198.365 33.735 -197.965 34.935 ;
        RECT -207.325 30.375 -206.925 31.575 ;
        RECT -225.245 27.015 -224.845 28.215 ;
        RECT -261.085 23.655 -260.685 24.855 ;
        RECT -332.765 20.295 -332.365 21.495 ;
        RECT -189.345 14.775 -189.065 55.155 ;
        RECT -188.785 45.995 -188.505 55.435 ;
        RECT -188.225 18.135 -187.945 55.155 ;
        RECT -187.665 45.995 -187.385 55.435 ;
        RECT -187.105 45.015 -186.825 55.155 ;
        RECT -186.545 45.995 -186.265 55.435 ;
        RECT -187.165 43.815 -186.765 45.015 ;
        RECT -185.985 41.655 -185.705 55.155 ;
        RECT -185.425 45.995 -185.145 55.435 ;
        RECT -184.865 45.015 -184.585 55.155 ;
        RECT -184.305 45.995 -184.025 55.435 ;
        RECT -184.925 43.815 -184.525 45.015 ;
        RECT -186.045 40.455 -185.645 41.655 ;
        RECT -183.745 38.295 -183.465 55.155 ;
        RECT -183.185 45.995 -182.905 55.435 ;
        RECT -182.625 45.015 -182.345 55.155 ;
        RECT -182.065 45.995 -181.785 55.435 ;
        RECT -182.685 43.815 -182.285 45.015 ;
        RECT -181.505 41.655 -181.225 55.155 ;
        RECT -180.945 45.995 -180.665 55.435 ;
        RECT -180.385 45.015 -180.105 55.155 ;
        RECT -179.825 45.995 -179.545 55.435 ;
        RECT -180.445 43.815 -180.045 45.015 ;
        RECT -181.565 40.455 -181.165 41.655 ;
        RECT -183.805 37.095 -183.405 38.295 ;
        RECT -179.265 34.935 -178.985 55.155 ;
        RECT -178.705 45.995 -178.425 55.435 ;
        RECT -178.145 45.015 -177.865 55.155 ;
        RECT -177.585 45.995 -177.305 55.435 ;
        RECT -178.205 43.815 -177.805 45.015 ;
        RECT -177.025 41.655 -176.745 55.155 ;
        RECT -176.465 45.995 -176.185 55.435 ;
        RECT -175.905 45.015 -175.625 55.155 ;
        RECT -175.345 45.995 -175.065 55.435 ;
        RECT -175.965 43.815 -175.565 45.015 ;
        RECT -177.085 40.455 -176.685 41.655 ;
        RECT -174.785 38.295 -174.505 55.155 ;
        RECT -174.225 45.995 -173.945 55.435 ;
        RECT -173.665 45.015 -173.385 55.155 ;
        RECT -173.105 45.995 -172.825 55.435 ;
        RECT -173.725 43.815 -173.325 45.015 ;
        RECT -172.545 41.655 -172.265 55.155 ;
        RECT -171.985 45.995 -171.705 55.435 ;
        RECT -171.425 45.015 -171.145 55.155 ;
        RECT -170.865 45.995 -170.585 55.435 ;
        RECT -171.485 43.815 -171.085 45.015 ;
        RECT -172.605 40.455 -172.205 41.655 ;
        RECT -174.845 37.095 -174.445 38.295 ;
        RECT -179.325 33.735 -178.925 34.935 ;
        RECT -170.305 31.575 -170.025 55.155 ;
        RECT -169.745 45.995 -169.465 55.435 ;
        RECT -169.185 45.015 -168.905 55.155 ;
        RECT -168.625 45.995 -168.345 55.435 ;
        RECT -169.245 43.815 -168.845 45.015 ;
        RECT -168.065 41.655 -167.785 55.155 ;
        RECT -167.505 45.995 -167.225 55.435 ;
        RECT -166.945 45.015 -166.665 55.155 ;
        RECT -166.385 45.995 -166.105 55.435 ;
        RECT -167.005 43.815 -166.605 45.015 ;
        RECT -168.125 40.455 -167.725 41.655 ;
        RECT -165.825 38.295 -165.545 55.155 ;
        RECT -165.265 45.995 -164.985 55.435 ;
        RECT -164.705 45.015 -164.425 55.155 ;
        RECT -164.145 45.995 -163.865 55.435 ;
        RECT -164.765 43.815 -164.365 45.015 ;
        RECT -163.585 41.655 -163.305 55.155 ;
        RECT -163.025 45.995 -162.745 55.435 ;
        RECT -162.465 45.015 -162.185 55.155 ;
        RECT -161.905 45.995 -161.625 55.435 ;
        RECT -162.525 43.815 -162.125 45.015 ;
        RECT -163.645 40.455 -163.245 41.655 ;
        RECT -165.885 37.095 -165.485 38.295 ;
        RECT -161.345 34.935 -161.065 55.155 ;
        RECT -160.785 45.995 -160.505 55.435 ;
        RECT -160.225 45.015 -159.945 55.155 ;
        RECT -159.665 45.995 -159.385 55.435 ;
        RECT -160.285 43.815 -159.885 45.015 ;
        RECT -159.105 41.655 -158.825 55.155 ;
        RECT -158.545 45.995 -158.265 55.435 ;
        RECT -157.985 45.015 -157.705 55.155 ;
        RECT -157.425 45.995 -157.145 55.435 ;
        RECT -158.045 43.815 -157.645 45.015 ;
        RECT -159.165 40.455 -158.765 41.655 ;
        RECT -156.865 38.295 -156.585 55.155 ;
        RECT -156.305 45.995 -156.025 55.435 ;
        RECT -155.745 45.015 -155.465 55.155 ;
        RECT -155.185 45.995 -154.905 55.435 ;
        RECT -155.805 43.815 -155.405 45.015 ;
        RECT -154.625 41.655 -154.345 55.155 ;
        RECT -154.065 45.995 -153.785 55.435 ;
        RECT -153.505 45.015 -153.225 55.155 ;
        RECT -152.945 45.995 -152.665 55.435 ;
        RECT -153.565 43.815 -153.165 45.015 ;
        RECT -154.685 40.455 -154.285 41.655 ;
        RECT -156.925 37.095 -156.525 38.295 ;
        RECT -161.405 33.735 -161.005 34.935 ;
        RECT -170.365 30.375 -169.965 31.575 ;
        RECT -152.385 28.215 -152.105 55.155 ;
        RECT -151.825 45.995 -151.545 55.435 ;
        RECT -151.265 45.015 -150.985 55.155 ;
        RECT -150.705 45.995 -150.425 55.435 ;
        RECT -151.325 43.815 -150.925 45.015 ;
        RECT -150.145 41.655 -149.865 55.155 ;
        RECT -149.585 45.995 -149.305 55.435 ;
        RECT -149.025 45.015 -148.745 55.155 ;
        RECT -148.465 45.995 -148.185 55.435 ;
        RECT -149.085 43.815 -148.685 45.015 ;
        RECT -150.205 40.455 -149.805 41.655 ;
        RECT -147.905 38.295 -147.625 55.155 ;
        RECT -147.345 45.995 -147.065 55.435 ;
        RECT -146.785 45.015 -146.505 55.155 ;
        RECT -146.225 45.995 -145.945 55.435 ;
        RECT -146.845 43.815 -146.445 45.015 ;
        RECT -145.665 41.655 -145.385 55.155 ;
        RECT -145.105 45.995 -144.825 55.435 ;
        RECT -144.545 45.015 -144.265 55.155 ;
        RECT -143.985 45.995 -143.705 55.435 ;
        RECT -144.605 43.815 -144.205 45.015 ;
        RECT -145.725 40.455 -145.325 41.655 ;
        RECT -147.965 37.095 -147.565 38.295 ;
        RECT -143.425 34.935 -143.145 55.155 ;
        RECT -142.865 45.995 -142.585 55.435 ;
        RECT -142.305 45.015 -142.025 55.155 ;
        RECT -141.745 45.995 -141.465 55.435 ;
        RECT -142.365 43.815 -141.965 45.015 ;
        RECT -141.185 41.655 -140.905 55.155 ;
        RECT -140.625 45.995 -140.345 55.435 ;
        RECT -140.065 45.015 -139.785 55.155 ;
        RECT -139.505 45.995 -139.225 55.435 ;
        RECT -140.125 43.815 -139.725 45.015 ;
        RECT -141.245 40.455 -140.845 41.655 ;
        RECT -138.945 38.295 -138.665 55.155 ;
        RECT -138.385 45.995 -138.105 55.435 ;
        RECT -137.825 45.015 -137.545 55.155 ;
        RECT -137.265 45.995 -136.985 55.435 ;
        RECT -137.885 43.815 -137.485 45.015 ;
        RECT -136.705 41.655 -136.425 55.155 ;
        RECT -136.145 45.995 -135.865 55.435 ;
        RECT -135.585 45.015 -135.305 55.155 ;
        RECT -135.025 45.995 -134.745 55.435 ;
        RECT -135.645 43.815 -135.245 45.015 ;
        RECT -136.765 40.455 -136.365 41.655 ;
        RECT -139.005 37.095 -138.605 38.295 ;
        RECT -143.485 33.735 -143.085 34.935 ;
        RECT -134.465 31.575 -134.185 55.155 ;
        RECT -133.905 45.995 -133.625 55.435 ;
        RECT -133.345 45.015 -133.065 55.155 ;
        RECT -132.785 45.995 -132.505 55.435 ;
        RECT -133.405 43.815 -133.005 45.015 ;
        RECT -132.225 41.655 -131.945 55.155 ;
        RECT -131.665 45.995 -131.385 55.435 ;
        RECT -131.105 45.015 -130.825 55.155 ;
        RECT -130.545 45.995 -130.265 55.435 ;
        RECT -131.165 43.815 -130.765 45.015 ;
        RECT -132.285 40.455 -131.885 41.655 ;
        RECT -129.985 38.295 -129.705 55.155 ;
        RECT -129.425 45.995 -129.145 55.435 ;
        RECT -128.865 45.015 -128.585 55.155 ;
        RECT -128.305 45.995 -128.025 55.435 ;
        RECT -128.925 43.815 -128.525 45.015 ;
        RECT -127.745 41.655 -127.465 55.155 ;
        RECT -127.185 45.995 -126.905 55.435 ;
        RECT -126.625 45.015 -126.345 55.155 ;
        RECT -126.065 45.995 -125.785 55.435 ;
        RECT -126.685 43.815 -126.285 45.015 ;
        RECT -127.805 40.455 -127.405 41.655 ;
        RECT -130.045 37.095 -129.645 38.295 ;
        RECT -125.505 34.935 -125.225 55.155 ;
        RECT -124.945 45.995 -124.665 55.435 ;
        RECT -124.385 45.015 -124.105 55.155 ;
        RECT -123.825 45.995 -123.545 55.435 ;
        RECT -124.445 43.815 -124.045 45.015 ;
        RECT -123.265 41.655 -122.985 55.155 ;
        RECT -122.705 45.995 -122.425 55.435 ;
        RECT -122.145 45.015 -121.865 55.155 ;
        RECT -121.585 45.995 -121.305 55.435 ;
        RECT -122.205 43.815 -121.805 45.015 ;
        RECT -123.325 40.455 -122.925 41.655 ;
        RECT -121.025 38.295 -120.745 55.155 ;
        RECT -120.465 45.995 -120.185 55.435 ;
        RECT -119.905 45.015 -119.625 55.155 ;
        RECT -119.345 45.995 -119.065 55.435 ;
        RECT -119.965 43.815 -119.565 45.015 ;
        RECT -118.785 41.655 -118.505 55.155 ;
        RECT -118.225 45.995 -117.945 55.435 ;
        RECT -117.665 45.015 -117.385 55.155 ;
        RECT -117.105 45.995 -116.825 55.435 ;
        RECT -117.725 43.815 -117.325 45.015 ;
        RECT -118.845 40.455 -118.445 41.655 ;
        RECT -121.085 37.095 -120.685 38.295 ;
        RECT -125.565 33.735 -125.165 34.935 ;
        RECT -134.525 30.375 -134.125 31.575 ;
        RECT -152.445 27.015 -152.045 28.215 ;
        RECT -116.545 24.855 -116.265 55.155 ;
        RECT -115.985 45.995 -115.705 55.435 ;
        RECT -115.425 45.015 -115.145 55.155 ;
        RECT -114.865 45.995 -114.585 55.435 ;
        RECT -115.485 43.815 -115.085 45.015 ;
        RECT -114.305 41.655 -114.025 55.155 ;
        RECT -113.745 45.995 -113.465 55.435 ;
        RECT -113.185 45.015 -112.905 55.155 ;
        RECT -112.625 45.995 -112.345 55.435 ;
        RECT -113.245 43.815 -112.845 45.015 ;
        RECT -114.365 40.455 -113.965 41.655 ;
        RECT -112.065 38.295 -111.785 55.155 ;
        RECT -111.505 45.995 -111.225 55.435 ;
        RECT -110.945 45.015 -110.665 55.155 ;
        RECT -110.385 45.995 -110.105 55.435 ;
        RECT -111.005 43.815 -110.605 45.015 ;
        RECT -109.825 41.655 -109.545 55.155 ;
        RECT -109.265 45.995 -108.985 55.435 ;
        RECT -108.705 45.015 -108.425 55.155 ;
        RECT -108.145 45.995 -107.865 55.435 ;
        RECT -108.765 43.815 -108.365 45.015 ;
        RECT -109.885 40.455 -109.485 41.655 ;
        RECT -112.125 37.095 -111.725 38.295 ;
        RECT -107.585 34.935 -107.305 55.155 ;
        RECT -107.025 45.995 -106.745 55.435 ;
        RECT -106.465 45.015 -106.185 55.155 ;
        RECT -105.905 45.995 -105.625 55.435 ;
        RECT -106.525 43.815 -106.125 45.015 ;
        RECT -105.345 41.655 -105.065 55.155 ;
        RECT -104.785 45.995 -104.505 55.435 ;
        RECT -104.225 45.015 -103.945 55.155 ;
        RECT -103.665 45.995 -103.385 55.435 ;
        RECT -104.285 43.815 -103.885 45.015 ;
        RECT -105.405 40.455 -105.005 41.655 ;
        RECT -103.105 38.295 -102.825 55.155 ;
        RECT -102.545 45.995 -102.265 55.435 ;
        RECT -101.985 45.015 -101.705 55.155 ;
        RECT -101.425 45.995 -101.145 55.435 ;
        RECT -102.045 43.815 -101.645 45.015 ;
        RECT -100.865 41.655 -100.585 55.155 ;
        RECT -100.305 45.995 -100.025 55.435 ;
        RECT -99.745 45.015 -99.465 55.155 ;
        RECT -99.185 45.995 -98.905 55.435 ;
        RECT -99.805 43.815 -99.405 45.015 ;
        RECT -100.925 40.455 -100.525 41.655 ;
        RECT -103.165 37.095 -102.765 38.295 ;
        RECT -107.645 33.735 -107.245 34.935 ;
        RECT -98.625 31.575 -98.345 55.155 ;
        RECT -98.065 45.995 -97.785 55.435 ;
        RECT -97.505 45.015 -97.225 55.155 ;
        RECT -96.945 45.995 -96.665 55.435 ;
        RECT -97.565 43.815 -97.165 45.015 ;
        RECT -96.385 41.655 -96.105 55.155 ;
        RECT -95.825 45.995 -95.545 55.435 ;
        RECT -95.265 45.015 -94.985 55.155 ;
        RECT -94.705 45.995 -94.425 55.435 ;
        RECT -95.325 43.815 -94.925 45.015 ;
        RECT -96.445 40.455 -96.045 41.655 ;
        RECT -94.145 38.295 -93.865 55.155 ;
        RECT -93.585 45.995 -93.305 55.435 ;
        RECT -93.025 45.015 -92.745 55.155 ;
        RECT -92.465 45.995 -92.185 55.435 ;
        RECT -93.085 43.815 -92.685 45.015 ;
        RECT -91.905 41.655 -91.625 55.155 ;
        RECT -91.345 45.995 -91.065 55.435 ;
        RECT -90.785 45.015 -90.505 55.155 ;
        RECT -90.225 45.995 -89.945 55.435 ;
        RECT -90.845 43.815 -90.445 45.015 ;
        RECT -91.965 40.455 -91.565 41.655 ;
        RECT -94.205 37.095 -93.805 38.295 ;
        RECT -89.665 34.935 -89.385 55.155 ;
        RECT -89.105 45.995 -88.825 55.435 ;
        RECT -88.545 45.015 -88.265 55.155 ;
        RECT -87.985 45.995 -87.705 55.435 ;
        RECT -88.605 43.815 -88.205 45.015 ;
        RECT -87.425 41.655 -87.145 55.155 ;
        RECT -86.865 45.995 -86.585 55.435 ;
        RECT -86.305 45.015 -86.025 55.155 ;
        RECT -85.745 45.995 -85.465 55.435 ;
        RECT -86.365 43.815 -85.965 45.015 ;
        RECT -87.485 40.455 -87.085 41.655 ;
        RECT -85.185 38.295 -84.905 55.155 ;
        RECT -84.625 45.995 -84.345 55.435 ;
        RECT -84.065 45.015 -83.785 55.155 ;
        RECT -83.505 45.995 -83.225 55.435 ;
        RECT -84.125 43.815 -83.725 45.015 ;
        RECT -82.945 41.655 -82.665 55.155 ;
        RECT -82.385 45.995 -82.105 55.435 ;
        RECT -81.825 45.015 -81.545 55.155 ;
        RECT -81.265 45.995 -80.985 55.435 ;
        RECT -81.885 43.815 -81.485 45.015 ;
        RECT -83.005 40.455 -82.605 41.655 ;
        RECT -85.245 37.095 -84.845 38.295 ;
        RECT -89.725 33.735 -89.325 34.935 ;
        RECT -98.685 30.375 -98.285 31.575 ;
        RECT -80.705 28.215 -80.425 55.155 ;
        RECT -80.145 45.995 -79.865 55.435 ;
        RECT -79.585 45.015 -79.305 55.155 ;
        RECT -79.025 45.995 -78.745 55.435 ;
        RECT -79.645 43.815 -79.245 45.015 ;
        RECT -78.465 41.655 -78.185 55.155 ;
        RECT -77.905 45.995 -77.625 55.435 ;
        RECT -77.345 45.015 -77.065 55.155 ;
        RECT -76.785 45.995 -76.505 55.435 ;
        RECT -77.405 43.815 -77.005 45.015 ;
        RECT -78.525 40.455 -78.125 41.655 ;
        RECT -76.225 38.295 -75.945 55.155 ;
        RECT -75.665 45.995 -75.385 55.435 ;
        RECT -75.105 45.015 -74.825 55.155 ;
        RECT -74.545 45.995 -74.265 55.435 ;
        RECT -75.165 43.815 -74.765 45.015 ;
        RECT -73.985 41.655 -73.705 55.155 ;
        RECT -73.425 45.995 -73.145 55.435 ;
        RECT -72.865 45.015 -72.585 55.155 ;
        RECT -72.305 45.995 -72.025 55.435 ;
        RECT -72.925 43.815 -72.525 45.015 ;
        RECT -74.045 40.455 -73.645 41.655 ;
        RECT -76.285 37.095 -75.885 38.295 ;
        RECT -71.745 34.935 -71.465 55.155 ;
        RECT -71.185 45.995 -70.905 55.435 ;
        RECT -70.625 45.015 -70.345 55.155 ;
        RECT -70.065 45.995 -69.785 55.435 ;
        RECT -70.685 43.815 -70.285 45.015 ;
        RECT -69.505 41.655 -69.225 55.155 ;
        RECT -68.945 45.995 -68.665 55.435 ;
        RECT -68.385 45.015 -68.105 55.155 ;
        RECT -67.825 45.995 -67.545 55.435 ;
        RECT -68.445 43.815 -68.045 45.015 ;
        RECT -69.565 40.455 -69.165 41.655 ;
        RECT -67.265 38.295 -66.985 55.155 ;
        RECT -66.705 45.995 -66.425 55.435 ;
        RECT -66.145 45.015 -65.865 55.155 ;
        RECT -65.585 45.995 -65.305 55.435 ;
        RECT -66.205 43.815 -65.805 45.015 ;
        RECT -65.025 41.655 -64.745 55.155 ;
        RECT -64.465 45.995 -64.185 55.435 ;
        RECT -63.905 45.015 -63.625 55.155 ;
        RECT -63.345 45.995 -63.065 55.435 ;
        RECT -63.965 43.815 -63.565 45.015 ;
        RECT -65.085 40.455 -64.685 41.655 ;
        RECT -67.325 37.095 -66.925 38.295 ;
        RECT -71.805 33.735 -71.405 34.935 ;
        RECT -62.785 31.575 -62.505 55.155 ;
        RECT -62.225 45.995 -61.945 55.435 ;
        RECT -61.665 45.015 -61.385 55.155 ;
        RECT -61.105 45.995 -60.825 55.435 ;
        RECT -61.725 43.815 -61.325 45.015 ;
        RECT -60.545 41.655 -60.265 55.155 ;
        RECT -59.985 45.995 -59.705 55.435 ;
        RECT -59.425 45.015 -59.145 55.155 ;
        RECT -58.865 45.995 -58.585 55.435 ;
        RECT -59.485 43.815 -59.085 45.015 ;
        RECT -60.605 40.455 -60.205 41.655 ;
        RECT -58.305 38.295 -58.025 55.155 ;
        RECT -57.745 45.995 -57.465 55.435 ;
        RECT -57.185 45.015 -56.905 55.155 ;
        RECT -56.625 45.995 -56.345 55.435 ;
        RECT -57.245 43.815 -56.845 45.015 ;
        RECT -56.065 41.655 -55.785 55.155 ;
        RECT -55.505 45.995 -55.225 55.435 ;
        RECT -54.945 45.015 -54.665 55.155 ;
        RECT -54.385 45.995 -54.105 55.435 ;
        RECT -55.005 43.815 -54.605 45.015 ;
        RECT -56.125 40.455 -55.725 41.655 ;
        RECT -58.365 37.095 -57.965 38.295 ;
        RECT -53.825 34.935 -53.545 55.155 ;
        RECT -53.265 45.995 -52.985 55.435 ;
        RECT -52.705 45.015 -52.425 55.155 ;
        RECT -52.145 45.995 -51.865 55.435 ;
        RECT -52.765 43.815 -52.365 45.015 ;
        RECT -51.585 41.655 -51.305 55.155 ;
        RECT -51.025 45.995 -50.745 55.435 ;
        RECT -50.465 45.015 -50.185 55.155 ;
        RECT -49.905 45.995 -49.625 55.435 ;
        RECT -50.525 43.815 -50.125 45.015 ;
        RECT -51.645 40.455 -51.245 41.655 ;
        RECT -49.345 38.295 -49.065 55.155 ;
        RECT -48.785 45.995 -48.505 55.435 ;
        RECT -48.225 45.015 -47.945 55.155 ;
        RECT -47.665 45.995 -47.385 55.435 ;
        RECT -48.285 43.815 -47.885 45.015 ;
        RECT -47.105 41.655 -46.825 55.155 ;
        RECT -46.545 45.995 -46.265 55.435 ;
        RECT -45.985 45.015 -45.705 55.155 ;
        RECT -45.425 45.995 -45.145 55.435 ;
        RECT -46.045 43.815 -45.645 45.015 ;
        RECT -47.165 40.455 -46.765 41.655 ;
        RECT -49.405 37.095 -49.005 38.295 ;
        RECT -53.885 33.735 -53.485 34.935 ;
        RECT -62.845 30.375 -62.445 31.575 ;
        RECT -80.765 27.015 -80.365 28.215 ;
        RECT -116.605 23.655 -116.205 24.855 ;
        RECT -44.865 21.495 -44.585 55.155 ;
        RECT -44.305 45.995 -44.025 55.435 ;
        RECT -43.745 45.015 -43.465 55.155 ;
        RECT -43.185 45.995 -42.905 55.435 ;
        RECT -43.805 43.815 -43.405 45.015 ;
        RECT -42.625 41.655 -42.345 55.155 ;
        RECT -42.065 45.995 -41.785 55.435 ;
        RECT -41.505 45.015 -41.225 55.155 ;
        RECT -40.945 45.995 -40.665 55.435 ;
        RECT -41.565 43.815 -41.165 45.015 ;
        RECT -42.685 40.455 -42.285 41.655 ;
        RECT -40.385 38.295 -40.105 55.155 ;
        RECT -39.825 45.995 -39.545 55.435 ;
        RECT -39.265 45.015 -38.985 55.155 ;
        RECT -38.705 45.995 -38.425 55.435 ;
        RECT -39.325 43.815 -38.925 45.015 ;
        RECT -38.145 41.655 -37.865 55.155 ;
        RECT -37.585 45.995 -37.305 55.435 ;
        RECT -37.025 45.015 -36.745 55.155 ;
        RECT -36.465 45.995 -36.185 55.435 ;
        RECT -37.085 43.815 -36.685 45.015 ;
        RECT -38.205 40.455 -37.805 41.655 ;
        RECT -40.445 37.095 -40.045 38.295 ;
        RECT -35.905 34.935 -35.625 55.155 ;
        RECT -35.345 45.995 -35.065 55.435 ;
        RECT -34.785 45.015 -34.505 55.155 ;
        RECT -34.225 45.995 -33.945 55.435 ;
        RECT -34.845 43.815 -34.445 45.015 ;
        RECT -33.665 41.655 -33.385 55.155 ;
        RECT -33.105 45.995 -32.825 55.435 ;
        RECT -32.545 45.015 -32.265 55.155 ;
        RECT -31.985 45.995 -31.705 55.435 ;
        RECT -32.605 43.815 -32.205 45.015 ;
        RECT -33.725 40.455 -33.325 41.655 ;
        RECT -31.425 38.295 -31.145 55.155 ;
        RECT -30.865 45.995 -30.585 55.435 ;
        RECT -30.305 45.015 -30.025 55.155 ;
        RECT -29.745 45.995 -29.465 55.435 ;
        RECT -30.365 43.815 -29.965 45.015 ;
        RECT -29.185 41.655 -28.905 55.155 ;
        RECT -28.625 45.995 -28.345 55.435 ;
        RECT -28.065 45.015 -27.785 55.155 ;
        RECT -27.505 45.995 -27.225 55.435 ;
        RECT -28.125 43.815 -27.725 45.015 ;
        RECT -29.245 40.455 -28.845 41.655 ;
        RECT -31.485 37.095 -31.085 38.295 ;
        RECT -35.965 33.735 -35.565 34.935 ;
        RECT -26.945 31.575 -26.665 55.155 ;
        RECT -26.385 45.995 -26.105 55.435 ;
        RECT -25.825 45.015 -25.545 55.155 ;
        RECT -25.265 45.995 -24.985 55.435 ;
        RECT -25.885 43.815 -25.485 45.015 ;
        RECT -24.705 41.655 -24.425 55.155 ;
        RECT -24.145 45.995 -23.865 55.435 ;
        RECT -23.585 45.015 -23.305 55.155 ;
        RECT -23.025 45.995 -22.745 55.435 ;
        RECT -23.645 43.815 -23.245 45.015 ;
        RECT -24.765 40.455 -24.365 41.655 ;
        RECT -22.465 38.295 -22.185 55.155 ;
        RECT -21.905 45.995 -21.625 55.435 ;
        RECT -21.345 45.015 -21.065 55.155 ;
        RECT -20.785 45.995 -20.505 55.435 ;
        RECT -21.405 43.815 -21.005 45.015 ;
        RECT -20.225 41.655 -19.945 55.155 ;
        RECT -19.665 45.995 -19.385 55.435 ;
        RECT -19.105 45.015 -18.825 55.155 ;
        RECT -18.545 45.995 -18.265 55.435 ;
        RECT -19.165 43.815 -18.765 45.015 ;
        RECT -20.285 40.455 -19.885 41.655 ;
        RECT -22.525 37.095 -22.125 38.295 ;
        RECT -17.985 34.935 -17.705 55.155 ;
        RECT -17.425 45.995 -17.145 55.435 ;
        RECT -16.865 45.015 -16.585 55.155 ;
        RECT -16.305 45.995 -16.025 55.435 ;
        RECT -16.925 43.815 -16.525 45.015 ;
        RECT -15.745 41.655 -15.465 55.155 ;
        RECT -15.185 45.995 -14.905 55.435 ;
        RECT -14.625 45.015 -14.345 55.155 ;
        RECT -14.065 45.995 -13.785 55.435 ;
        RECT -14.685 43.815 -14.285 45.015 ;
        RECT -15.805 40.455 -15.405 41.655 ;
        RECT -13.505 38.295 -13.225 55.155 ;
        RECT -12.945 45.995 -12.665 55.435 ;
        RECT -12.385 45.015 -12.105 55.155 ;
        RECT -11.825 45.995 -11.545 55.435 ;
        RECT -12.445 43.815 -12.045 45.015 ;
        RECT -11.265 41.655 -10.985 55.155 ;
        RECT -10.705 45.995 -10.425 55.435 ;
        RECT -10.145 45.015 -9.865 55.155 ;
        RECT -9.585 45.995 -9.305 55.435 ;
        RECT -10.205 43.815 -9.805 45.015 ;
        RECT -11.325 40.455 -10.925 41.655 ;
        RECT -13.565 37.095 -13.165 38.295 ;
        RECT -18.045 33.735 -17.645 34.935 ;
        RECT -27.005 30.375 -26.605 31.575 ;
        RECT -9.025 28.215 -8.745 55.155 ;
        RECT -8.465 45.995 -8.185 55.435 ;
        RECT -7.905 45.015 -7.625 55.155 ;
        RECT -7.345 45.995 -7.065 55.435 ;
        RECT -7.965 43.815 -7.565 45.015 ;
        RECT -6.785 41.655 -6.505 55.155 ;
        RECT -6.225 45.995 -5.945 55.435 ;
        RECT -5.665 45.015 -5.385 55.155 ;
        RECT -5.105 45.995 -4.825 55.435 ;
        RECT -5.725 43.815 -5.325 45.015 ;
        RECT -6.845 40.455 -6.445 41.655 ;
        RECT -4.545 38.295 -4.265 55.155 ;
        RECT -3.985 45.995 -3.705 55.435 ;
        RECT -3.425 45.015 -3.145 55.155 ;
        RECT -2.865 45.995 -2.585 55.435 ;
        RECT -3.485 43.815 -3.085 45.015 ;
        RECT -2.305 41.655 -2.025 55.155 ;
        RECT -1.745 45.995 -1.465 55.435 ;
        RECT -1.185 45.015 -0.905 55.155 ;
        RECT -0.625 45.995 -0.345 55.435 ;
        RECT -1.245 43.815 -0.845 45.015 ;
        RECT -2.365 40.455 -1.965 41.655 ;
        RECT -4.605 37.095 -4.205 38.295 ;
        RECT -0.065 34.935 0.215 55.155 ;
        RECT 0.495 45.995 0.775 55.435 ;
        RECT 1.055 45.015 1.335 55.155 ;
        RECT 1.615 45.995 1.895 55.435 ;
        RECT 0.995 43.815 1.395 45.015 ;
        RECT 2.175 41.655 2.455 55.155 ;
        RECT 2.735 45.995 3.015 55.435 ;
        RECT 3.295 45.015 3.575 55.155 ;
        RECT 3.855 45.995 4.135 55.435 ;
        RECT 3.235 43.815 3.635 45.015 ;
        RECT 2.115 40.455 2.515 41.655 ;
        RECT 4.415 38.295 4.695 55.155 ;
        RECT 4.975 45.995 5.255 55.435 ;
        RECT 5.535 45.015 5.815 55.155 ;
        RECT 6.095 45.995 6.375 55.435 ;
        RECT 5.475 43.815 5.875 45.015 ;
        RECT 6.655 41.655 6.935 55.155 ;
        RECT 7.215 45.995 7.495 55.435 ;
        RECT 7.775 45.015 8.055 55.155 ;
        RECT 8.335 45.995 8.615 55.435 ;
        RECT 7.715 43.815 8.115 45.015 ;
        RECT 6.595 40.455 6.995 41.655 ;
        RECT 4.355 37.095 4.755 38.295 ;
        RECT -0.125 33.735 0.275 34.935 ;
        RECT 8.895 31.575 9.175 55.155 ;
        RECT 9.455 45.995 9.735 55.435 ;
        RECT 10.015 45.015 10.295 55.155 ;
        RECT 10.575 45.995 10.855 55.435 ;
        RECT 9.955 43.815 10.355 45.015 ;
        RECT 11.135 41.655 11.415 55.155 ;
        RECT 11.695 45.995 11.975 55.435 ;
        RECT 12.255 45.015 12.535 55.155 ;
        RECT 12.815 45.995 13.095 55.435 ;
        RECT 12.195 43.815 12.595 45.015 ;
        RECT 11.075 40.455 11.475 41.655 ;
        RECT 13.375 38.295 13.655 55.155 ;
        RECT 13.935 45.995 14.215 55.435 ;
        RECT 14.495 45.015 14.775 55.155 ;
        RECT 15.055 45.995 15.335 55.435 ;
        RECT 14.435 43.815 14.835 45.015 ;
        RECT 15.615 41.655 15.895 55.155 ;
        RECT 16.175 45.995 16.455 55.435 ;
        RECT 16.735 45.015 17.015 55.155 ;
        RECT 17.295 45.995 17.575 55.435 ;
        RECT 16.675 43.815 17.075 45.015 ;
        RECT 15.555 40.455 15.955 41.655 ;
        RECT 13.315 37.095 13.715 38.295 ;
        RECT 17.855 34.935 18.135 55.155 ;
        RECT 18.415 45.995 18.695 55.435 ;
        RECT 18.975 45.015 19.255 55.155 ;
        RECT 19.535 45.995 19.815 55.435 ;
        RECT 18.915 43.815 19.315 45.015 ;
        RECT 20.095 41.655 20.375 55.155 ;
        RECT 20.655 45.995 20.935 55.435 ;
        RECT 21.215 45.015 21.495 55.155 ;
        RECT 21.775 45.995 22.055 55.435 ;
        RECT 21.155 43.815 21.555 45.015 ;
        RECT 20.035 40.455 20.435 41.655 ;
        RECT 22.335 38.295 22.615 55.155 ;
        RECT 22.895 45.995 23.175 55.435 ;
        RECT 23.455 45.015 23.735 55.155 ;
        RECT 24.015 45.995 24.295 55.435 ;
        RECT 23.395 43.815 23.795 45.015 ;
        RECT 24.575 41.655 24.855 55.155 ;
        RECT 25.135 45.995 25.415 55.435 ;
        RECT 25.695 45.015 25.975 55.155 ;
        RECT 26.255 45.995 26.535 55.435 ;
        RECT 25.635 43.815 26.035 45.015 ;
        RECT 24.515 40.455 24.915 41.655 ;
        RECT 22.275 37.095 22.675 38.295 ;
        RECT 17.795 33.735 18.195 34.935 ;
        RECT 8.835 30.375 9.235 31.575 ;
        RECT -9.085 27.015 -8.685 28.215 ;
        RECT 26.815 24.855 27.095 55.155 ;
        RECT 27.375 45.995 27.655 55.435 ;
        RECT 27.935 45.015 28.215 55.155 ;
        RECT 28.495 45.995 28.775 55.435 ;
        RECT 27.875 43.815 28.275 45.015 ;
        RECT 29.055 41.655 29.335 55.155 ;
        RECT 29.615 45.995 29.895 55.435 ;
        RECT 30.175 45.015 30.455 55.155 ;
        RECT 30.735 45.995 31.015 55.435 ;
        RECT 30.115 43.815 30.515 45.015 ;
        RECT 28.995 40.455 29.395 41.655 ;
        RECT 31.295 38.295 31.575 55.155 ;
        RECT 31.855 45.995 32.135 55.435 ;
        RECT 32.415 45.015 32.695 55.155 ;
        RECT 32.975 45.995 33.255 55.435 ;
        RECT 32.355 43.815 32.755 45.015 ;
        RECT 33.535 41.655 33.815 55.155 ;
        RECT 34.095 45.995 34.375 55.435 ;
        RECT 34.655 45.015 34.935 55.155 ;
        RECT 35.215 45.995 35.495 55.435 ;
        RECT 34.595 43.815 34.995 45.015 ;
        RECT 33.475 40.455 33.875 41.655 ;
        RECT 31.235 37.095 31.635 38.295 ;
        RECT 35.775 34.935 36.055 55.155 ;
        RECT 36.335 45.995 36.615 55.435 ;
        RECT 36.895 45.015 37.175 55.155 ;
        RECT 37.455 45.995 37.735 55.435 ;
        RECT 36.835 43.815 37.235 45.015 ;
        RECT 38.015 41.655 38.295 55.155 ;
        RECT 38.575 45.995 38.855 55.435 ;
        RECT 39.135 45.015 39.415 55.155 ;
        RECT 39.695 45.995 39.975 55.435 ;
        RECT 39.075 43.815 39.475 45.015 ;
        RECT 37.955 40.455 38.355 41.655 ;
        RECT 40.255 38.295 40.535 55.155 ;
        RECT 40.815 45.995 41.095 55.435 ;
        RECT 41.375 45.015 41.655 55.155 ;
        RECT 41.935 45.995 42.215 55.435 ;
        RECT 41.315 43.815 41.715 45.015 ;
        RECT 42.495 41.655 42.775 55.155 ;
        RECT 43.055 45.995 43.335 55.435 ;
        RECT 43.615 45.015 43.895 55.155 ;
        RECT 44.175 45.995 44.455 55.435 ;
        RECT 43.555 43.815 43.955 45.015 ;
        RECT 42.435 40.455 42.835 41.655 ;
        RECT 40.195 37.095 40.595 38.295 ;
        RECT 35.715 33.735 36.115 34.935 ;
        RECT 44.735 31.575 45.015 55.155 ;
        RECT 45.295 45.995 45.575 55.435 ;
        RECT 45.855 45.015 46.135 55.155 ;
        RECT 46.415 45.995 46.695 55.435 ;
        RECT 45.795 43.815 46.195 45.015 ;
        RECT 46.975 41.655 47.255 55.155 ;
        RECT 47.535 45.995 47.815 55.435 ;
        RECT 48.095 45.015 48.375 55.155 ;
        RECT 48.655 45.995 48.935 55.435 ;
        RECT 48.035 43.815 48.435 45.015 ;
        RECT 46.915 40.455 47.315 41.655 ;
        RECT 49.215 38.295 49.495 55.155 ;
        RECT 49.775 45.995 50.055 55.435 ;
        RECT 50.335 45.015 50.615 55.155 ;
        RECT 50.895 45.995 51.175 55.435 ;
        RECT 50.275 43.815 50.675 45.015 ;
        RECT 51.455 41.655 51.735 55.155 ;
        RECT 52.015 45.995 52.295 55.435 ;
        RECT 52.575 45.015 52.855 55.155 ;
        RECT 53.135 45.995 53.415 55.435 ;
        RECT 52.515 43.815 52.915 45.015 ;
        RECT 51.395 40.455 51.795 41.655 ;
        RECT 49.155 37.095 49.555 38.295 ;
        RECT 53.695 34.935 53.975 55.155 ;
        RECT 54.255 45.995 54.535 55.435 ;
        RECT 54.815 45.015 55.095 55.155 ;
        RECT 55.375 45.995 55.655 55.435 ;
        RECT 54.755 43.815 55.155 45.015 ;
        RECT 55.935 41.655 56.215 55.155 ;
        RECT 56.495 45.995 56.775 55.435 ;
        RECT 57.055 45.015 57.335 55.155 ;
        RECT 57.615 45.995 57.895 55.435 ;
        RECT 56.995 43.815 57.395 45.015 ;
        RECT 55.875 40.455 56.275 41.655 ;
        RECT 58.175 38.295 58.455 55.155 ;
        RECT 58.735 45.995 59.015 55.435 ;
        RECT 59.295 45.015 59.575 55.155 ;
        RECT 59.855 45.995 60.135 55.435 ;
        RECT 59.235 43.815 59.635 45.015 ;
        RECT 60.415 41.655 60.695 55.155 ;
        RECT 60.975 45.995 61.255 55.435 ;
        RECT 61.535 45.015 61.815 55.155 ;
        RECT 62.095 45.995 62.375 55.435 ;
        RECT 61.475 43.815 61.875 45.015 ;
        RECT 60.355 40.455 60.755 41.655 ;
        RECT 58.115 37.095 58.515 38.295 ;
        RECT 53.635 33.735 54.035 34.935 ;
        RECT 44.675 30.375 45.075 31.575 ;
        RECT 62.655 28.215 62.935 55.155 ;
        RECT 63.215 45.995 63.495 55.435 ;
        RECT 63.775 45.015 64.055 55.155 ;
        RECT 64.335 45.995 64.615 55.435 ;
        RECT 63.715 43.815 64.115 45.015 ;
        RECT 64.895 41.655 65.175 55.155 ;
        RECT 65.455 45.995 65.735 55.435 ;
        RECT 66.015 45.015 66.295 55.155 ;
        RECT 66.575 45.995 66.855 55.435 ;
        RECT 65.955 43.815 66.355 45.015 ;
        RECT 64.835 40.455 65.235 41.655 ;
        RECT 67.135 38.295 67.415 55.155 ;
        RECT 67.695 45.995 67.975 55.435 ;
        RECT 68.255 45.015 68.535 55.155 ;
        RECT 68.815 45.995 69.095 55.435 ;
        RECT 68.195 43.815 68.595 45.015 ;
        RECT 69.375 41.655 69.655 55.155 ;
        RECT 69.935 45.995 70.215 55.435 ;
        RECT 70.495 45.015 70.775 55.155 ;
        RECT 71.055 45.995 71.335 55.435 ;
        RECT 70.435 43.815 70.835 45.015 ;
        RECT 69.315 40.455 69.715 41.655 ;
        RECT 67.075 37.095 67.475 38.295 ;
        RECT 71.615 34.935 71.895 55.155 ;
        RECT 72.175 45.995 72.455 55.435 ;
        RECT 72.735 45.015 73.015 55.155 ;
        RECT 73.295 45.995 73.575 55.435 ;
        RECT 72.675 43.815 73.075 45.015 ;
        RECT 73.855 41.655 74.135 55.155 ;
        RECT 74.415 45.995 74.695 55.435 ;
        RECT 74.975 45.015 75.255 55.155 ;
        RECT 75.535 45.995 75.815 55.435 ;
        RECT 74.915 43.815 75.315 45.015 ;
        RECT 73.795 40.455 74.195 41.655 ;
        RECT 76.095 38.295 76.375 55.155 ;
        RECT 76.655 45.995 76.935 55.435 ;
        RECT 77.215 45.015 77.495 55.155 ;
        RECT 77.775 45.995 78.055 55.435 ;
        RECT 77.155 43.815 77.555 45.015 ;
        RECT 78.335 41.655 78.615 55.155 ;
        RECT 78.895 45.995 79.175 55.435 ;
        RECT 79.455 45.015 79.735 55.155 ;
        RECT 80.015 45.995 80.295 55.435 ;
        RECT 79.395 43.815 79.795 45.015 ;
        RECT 78.275 40.455 78.675 41.655 ;
        RECT 76.035 37.095 76.435 38.295 ;
        RECT 71.555 33.735 71.955 34.935 ;
        RECT 80.575 31.575 80.855 55.155 ;
        RECT 81.135 45.995 81.415 55.435 ;
        RECT 81.695 45.015 81.975 55.155 ;
        RECT 82.255 45.995 82.535 55.435 ;
        RECT 81.635 43.815 82.035 45.015 ;
        RECT 82.815 41.655 83.095 55.155 ;
        RECT 83.375 45.995 83.655 55.435 ;
        RECT 83.935 45.015 84.215 55.155 ;
        RECT 84.495 45.995 84.775 55.435 ;
        RECT 83.875 43.815 84.275 45.015 ;
        RECT 82.755 40.455 83.155 41.655 ;
        RECT 85.055 38.295 85.335 55.155 ;
        RECT 85.615 45.995 85.895 55.435 ;
        RECT 86.175 45.015 86.455 55.155 ;
        RECT 86.735 45.995 87.015 55.435 ;
        RECT 86.115 43.815 86.515 45.015 ;
        RECT 87.295 41.655 87.575 55.155 ;
        RECT 87.855 45.995 88.135 55.435 ;
        RECT 88.415 45.015 88.695 55.155 ;
        RECT 88.975 45.995 89.255 55.435 ;
        RECT 88.355 43.815 88.755 45.015 ;
        RECT 87.235 40.455 87.635 41.655 ;
        RECT 84.995 37.095 85.395 38.295 ;
        RECT 89.535 34.935 89.815 55.155 ;
        RECT 90.095 45.995 90.375 55.435 ;
        RECT 90.655 45.015 90.935 55.155 ;
        RECT 91.215 45.995 91.495 55.435 ;
        RECT 90.595 43.815 90.995 45.015 ;
        RECT 91.775 41.655 92.055 55.155 ;
        RECT 92.335 45.995 92.615 55.435 ;
        RECT 92.895 45.015 93.175 55.155 ;
        RECT 93.455 45.995 93.735 55.435 ;
        RECT 92.835 43.815 93.235 45.015 ;
        RECT 91.715 40.455 92.115 41.655 ;
        RECT 94.015 38.295 94.295 55.155 ;
        RECT 94.575 45.995 94.855 55.435 ;
        RECT 95.135 45.015 95.415 55.155 ;
        RECT 95.695 45.995 95.975 55.435 ;
        RECT 95.075 43.815 95.475 45.015 ;
        RECT 96.255 41.655 96.535 55.155 ;
        RECT 96.815 45.995 97.095 55.435 ;
        RECT 97.375 45.015 97.655 55.155 ;
        RECT 97.935 45.995 98.215 55.435 ;
        RECT 98.495 45.405 98.775 54.995 ;
        RECT 99.055 45.995 99.335 55.435 ;
        RECT 99.615 45.405 99.895 54.995 ;
        RECT 100.175 45.405 100.455 55.435 ;
        RECT 97.315 43.815 97.715 45.015 ;
        RECT 98.495 45.005 100.455 45.405 ;
        RECT 96.195 40.455 96.595 41.655 ;
        RECT 93.955 37.095 94.355 38.295 ;
        RECT 89.475 33.735 89.875 34.935 ;
        RECT 80.515 30.375 80.915 31.575 ;
        RECT 62.595 27.015 62.995 28.215 ;
        RECT 26.755 23.655 27.155 24.855 ;
        RECT -44.925 20.295 -44.525 21.495 ;
        RECT -188.285 16.935 -187.885 18.135 ;
        RECT -189.405 13.575 -189.005 14.775 ;
        RECT 124.705 9.550 125.505 55.595 ;
        RECT 274.700 54.620 289.200 55.620 ;
        RECT 274.700 44.250 275.700 54.620 ;
        RECT 168.115 43.750 275.700 44.250 ;
        RECT 279.200 44.540 289.200 45.540 ;
        RECT 168.115 34.250 168.495 43.750 ;
        RECT 279.200 42.750 280.200 44.540 ;
        RECT 174.115 42.250 280.200 42.750 ;
        RECT 174.115 34.250 174.495 42.250 ;
        RECT 298.860 42.050 299.140 45.230 ;
        RECT 178.045 40.750 280.200 41.250 ;
        RECT 178.045 34.315 178.425 40.750 ;
        RECT 180.185 39.250 275.700 39.750 ;
        RECT 180.185 34.315 180.565 39.250 ;
        RECT 186.615 37.750 271.200 38.250 ;
        RECT 186.615 34.250 186.995 37.750 ;
        RECT 178.590 28.740 178.970 29.640 ;
        RECT 179.710 28.740 180.090 29.640 ;
        RECT 174.110 26.350 174.490 27.250 ;
        RECT 171.870 24.350 172.250 25.250 ;
        RECT 170.750 22.350 171.130 23.250 ;
        RECT 170.740 21.240 171.140 22.350 ;
        RECT 171.860 21.240 172.260 24.350 ;
        RECT 172.990 22.350 173.370 23.250 ;
        RECT 172.980 21.240 173.380 22.350 ;
        RECT 174.100 21.240 174.500 26.350 ;
        RECT 176.350 24.350 176.730 25.250 ;
        RECT 175.230 22.350 175.610 23.250 ;
        RECT 175.220 21.240 175.620 22.350 ;
        RECT 176.340 21.240 176.740 24.350 ;
        RECT 177.470 22.350 177.850 23.250 ;
        RECT 177.460 21.240 177.860 22.350 ;
        RECT 178.580 21.240 178.980 28.740 ;
        RECT 179.700 21.240 180.100 28.740 ;
        RECT 184.190 26.350 184.570 27.250 ;
        RECT 181.950 24.350 182.330 25.250 ;
        RECT 180.830 22.350 181.210 23.250 ;
        RECT 180.820 21.240 181.220 22.350 ;
        RECT 181.940 21.240 182.340 24.350 ;
        RECT 183.070 22.350 183.450 23.250 ;
        RECT 183.060 21.240 183.460 22.350 ;
        RECT 184.180 21.240 184.580 26.350 ;
        RECT 186.430 24.350 186.810 25.250 ;
        RECT 185.310 22.350 185.690 23.250 ;
        RECT 185.300 21.240 185.700 22.350 ;
        RECT 186.420 21.240 186.820 24.350 ;
        RECT 187.550 22.350 187.930 23.250 ;
        RECT 187.540 21.240 187.940 22.350 ;
        RECT 169.120 11.185 169.400 20.625 ;
        RECT 170.240 11.185 170.520 20.625 ;
        RECT 170.800 11.625 171.080 21.240 ;
        RECT 171.360 11.185 171.640 20.625 ;
        RECT 171.920 11.625 172.200 21.240 ;
        RECT 172.480 11.185 172.760 20.625 ;
        RECT 173.040 11.625 173.320 21.240 ;
        RECT 173.600 11.185 173.880 20.625 ;
        RECT 174.160 11.625 174.440 21.240 ;
        RECT 174.720 11.185 175.000 20.625 ;
        RECT 175.280 11.625 175.560 21.240 ;
        RECT 175.840 11.185 176.120 20.625 ;
        RECT 176.400 11.625 176.680 21.240 ;
        RECT 176.960 11.185 177.240 20.625 ;
        RECT 177.520 11.625 177.800 21.240 ;
        RECT 178.080 11.185 178.360 20.625 ;
        RECT 178.640 11.625 178.920 21.240 ;
        RECT 179.200 11.185 179.480 20.625 ;
        RECT 179.760 11.625 180.040 21.240 ;
        RECT 180.320 11.185 180.600 20.625 ;
        RECT 180.880 11.625 181.160 21.240 ;
        RECT 181.440 11.185 181.720 20.625 ;
        RECT 182.000 11.625 182.280 21.240 ;
        RECT 182.560 11.185 182.840 20.625 ;
        RECT 183.120 11.625 183.400 21.240 ;
        RECT 183.680 11.185 183.960 20.625 ;
        RECT 184.240 11.625 184.520 21.240 ;
        RECT 184.800 11.185 185.080 20.625 ;
        RECT 185.360 11.625 185.640 21.240 ;
        RECT 185.920 11.185 186.200 20.625 ;
        RECT 186.480 11.625 186.760 21.240 ;
        RECT 187.040 11.185 187.320 20.625 ;
        RECT 187.600 11.625 187.880 21.240 ;
        RECT 188.160 11.185 188.440 20.625 ;
        RECT 189.280 11.185 189.560 20.625 ;
        RECT 270.200 15.300 271.200 37.750 ;
        RECT 274.700 25.380 275.700 39.250 ;
        RECT 279.200 35.460 280.200 40.750 ;
        RECT 279.200 34.460 289.200 35.460 ;
        RECT 298.860 34.770 299.140 39.630 ;
        RECT 299.420 34.210 299.700 55.310 ;
        RECT 300.540 47.650 300.820 56.100 ;
        RECT 316.220 52.130 316.500 61.000 ;
        RECT 334.140 60.300 334.420 61.000 ;
        RECT 335.260 60.300 335.540 61.140 ;
        RECT 334.140 60.020 335.540 60.300 ;
        RECT 322.380 47.650 322.660 52.510 ;
        RECT 336.940 47.650 337.220 61.140 ;
        RECT 351.920 61.000 352.480 73.270 ;
        RECT 369.840 61.000 370.400 76.630 ;
        RECT 387.760 61.000 388.320 79.990 ;
        RECT 405.680 61.000 406.240 83.350 ;
        RECT 423.600 61.000 424.160 86.710 ;
        RECT 441.520 61.000 442.080 90.070 ;
        RECT 459.440 61.000 460.000 93.430 ;
        RECT 352.060 47.650 352.340 61.000 ;
        RECT 359.900 47.510 360.180 48.030 ;
        RECT 369.980 47.650 370.260 61.000 ;
        RECT 375.020 47.510 375.300 48.030 ;
        RECT 387.900 47.650 388.180 61.000 ;
        RECT 394.060 47.510 394.340 48.030 ;
        RECT 405.820 47.650 406.100 61.000 ;
        RECT 417.020 47.510 417.300 48.030 ;
        RECT 423.740 47.650 424.020 61.000 ;
        RECT 441.660 49.660 441.940 61.000 ;
        RECT 441.660 49.380 443.060 49.660 ;
        RECT 432.140 47.510 432.420 48.030 ;
        RECT 310.060 46.860 310.340 46.910 ;
        RECT 309.500 46.580 310.340 46.860 ;
        RECT 302.780 31.970 303.060 39.070 ;
        RECT 308.380 38.550 308.660 39.070 ;
        RECT 274.700 24.380 289.200 25.380 ;
        RECT 270.200 14.300 289.200 15.300 ;
        RECT 168.340 10.685 190.340 11.185 ;
        RECT 183.905 10.305 184.805 10.685 ;
        RECT 124.705 9.150 180.045 9.550 ;
        RECT 230.260 9.505 235.190 9.885 ;
        RECT 179.665 4.050 180.045 9.150 ;
        RECT 232.295 9.105 233.195 9.505 ;
        RECT 235.860 7.720 236.240 11.670 ;
        RECT 297.740 11.250 298.020 18.350 ;
        RECT 298.860 15.590 299.140 16.110 ;
        RECT 181.405 5.905 186.305 6.295 ;
        RECT 230.260 5.145 235.190 5.525 ;
        RECT 232.255 4.940 233.155 5.145 ;
        RECT 232.295 4.295 233.195 4.500 ;
        RECT 230.260 3.915 235.190 4.295 ;
        RECT 223.200 3.190 224.400 3.300 ;
        RECT 171.405 2.810 224.400 3.190 ;
        RECT 223.200 2.700 224.400 2.810 ;
        RECT 235.860 1.720 237.460 7.720 ;
        RECT 286.700 4.220 289.200 5.220 ;
        RECT 298.300 4.390 298.580 7.710 ;
        RECT 299.420 6.770 299.700 7.710 ;
        RECT 173.200 1.010 181.525 1.390 ;
        RECT 232.295 -0.065 233.195 0.335 ;
        RECT 230.260 -0.445 235.190 -0.065 ;
        RECT 173.200 -1.390 181.525 -1.010 ;
        RECT 235.860 -2.230 236.240 1.720 ;
        RECT 223.320 -2.810 224.520 -2.700 ;
        RECT 171.405 -3.190 224.520 -2.810 ;
        RECT 223.320 -3.300 224.520 -3.190 ;
        RECT 179.665 -9.150 180.045 -4.050 ;
        RECT 298.300 -4.100 298.580 -4.050 ;
        RECT 299.420 -4.100 299.700 -4.050 ;
        RECT 229.700 -5.485 235.700 -4.265 ;
        RECT 298.300 -4.380 299.700 -4.100 ;
        RECT 298.300 -4.430 298.580 -4.380 ;
        RECT 299.420 -4.430 299.700 -4.380 ;
        RECT 229.440 -5.865 235.960 -5.485 ;
        RECT 286.700 -5.860 289.200 -4.860 ;
        RECT 181.405 -6.300 186.305 -5.910 ;
        RECT 230.275 -8.550 230.655 -6.535 ;
        RECT 233.790 -8.550 234.170 -6.535 ;
        RECT 298.860 -7.230 299.140 -5.170 ;
        RECT 124.705 -9.550 180.045 -9.150 ;
        RECT 229.895 -9.450 230.655 -8.550 ;
        RECT 233.410 -9.450 234.170 -8.550 ;
        RECT -189.405 -14.775 -189.005 -13.575 ;
        RECT -332.765 -21.495 -332.365 -20.295 ;
        RECT -404.445 -24.855 -404.045 -23.655 ;
        RECT -440.285 -28.215 -439.885 -27.015 ;
        RECT -458.205 -31.575 -457.805 -30.375 ;
        RECT -467.165 -34.935 -466.765 -33.735 ;
        RECT -471.645 -38.295 -471.245 -37.095 ;
        RECT -473.885 -41.655 -473.485 -40.455 ;
        RECT -477.745 -45.405 -475.785 -45.005 ;
        RECT -475.005 -45.015 -474.605 -43.815 ;
        RECT -477.745 -55.435 -477.465 -45.405 ;
        RECT -477.185 -54.995 -476.905 -45.405 ;
        RECT -476.625 -55.435 -476.345 -45.995 ;
        RECT -476.065 -54.995 -475.785 -45.405 ;
        RECT -475.505 -55.435 -475.225 -45.995 ;
        RECT -474.945 -55.155 -474.665 -45.015 ;
        RECT -474.385 -55.435 -474.105 -45.995 ;
        RECT -473.825 -55.155 -473.545 -41.655 ;
        RECT -472.765 -45.015 -472.365 -43.815 ;
        RECT -473.265 -55.435 -472.985 -45.995 ;
        RECT -472.705 -55.155 -472.425 -45.015 ;
        RECT -472.145 -55.435 -471.865 -45.995 ;
        RECT -471.585 -55.155 -471.305 -38.295 ;
        RECT -469.405 -41.655 -469.005 -40.455 ;
        RECT -470.525 -45.015 -470.125 -43.815 ;
        RECT -471.025 -55.435 -470.745 -45.995 ;
        RECT -470.465 -55.155 -470.185 -45.015 ;
        RECT -469.905 -55.435 -469.625 -45.995 ;
        RECT -469.345 -55.155 -469.065 -41.655 ;
        RECT -468.285 -45.015 -467.885 -43.815 ;
        RECT -468.785 -55.435 -468.505 -45.995 ;
        RECT -468.225 -55.155 -467.945 -45.015 ;
        RECT -467.665 -55.435 -467.385 -45.995 ;
        RECT -467.105 -55.155 -466.825 -34.935 ;
        RECT -462.685 -38.295 -462.285 -37.095 ;
        RECT -464.925 -41.655 -464.525 -40.455 ;
        RECT -466.045 -45.015 -465.645 -43.815 ;
        RECT -466.545 -55.435 -466.265 -45.995 ;
        RECT -465.985 -55.155 -465.705 -45.015 ;
        RECT -465.425 -55.435 -465.145 -45.995 ;
        RECT -464.865 -55.155 -464.585 -41.655 ;
        RECT -463.805 -45.015 -463.405 -43.815 ;
        RECT -464.305 -55.435 -464.025 -45.995 ;
        RECT -463.745 -55.155 -463.465 -45.015 ;
        RECT -463.185 -55.435 -462.905 -45.995 ;
        RECT -462.625 -55.155 -462.345 -38.295 ;
        RECT -460.445 -41.655 -460.045 -40.455 ;
        RECT -461.565 -45.015 -461.165 -43.815 ;
        RECT -462.065 -55.435 -461.785 -45.995 ;
        RECT -461.505 -55.155 -461.225 -45.015 ;
        RECT -460.945 -55.435 -460.665 -45.995 ;
        RECT -460.385 -55.155 -460.105 -41.655 ;
        RECT -459.325 -45.015 -458.925 -43.815 ;
        RECT -459.825 -55.435 -459.545 -45.995 ;
        RECT -459.265 -55.155 -458.985 -45.015 ;
        RECT -458.705 -55.435 -458.425 -45.995 ;
        RECT -458.145 -55.155 -457.865 -31.575 ;
        RECT -449.245 -34.935 -448.845 -33.735 ;
        RECT -453.725 -38.295 -453.325 -37.095 ;
        RECT -455.965 -41.655 -455.565 -40.455 ;
        RECT -457.085 -45.015 -456.685 -43.815 ;
        RECT -457.585 -55.435 -457.305 -45.995 ;
        RECT -457.025 -55.155 -456.745 -45.015 ;
        RECT -456.465 -55.435 -456.185 -45.995 ;
        RECT -455.905 -55.155 -455.625 -41.655 ;
        RECT -454.845 -45.015 -454.445 -43.815 ;
        RECT -455.345 -55.435 -455.065 -45.995 ;
        RECT -454.785 -55.155 -454.505 -45.015 ;
        RECT -454.225 -55.435 -453.945 -45.995 ;
        RECT -453.665 -55.155 -453.385 -38.295 ;
        RECT -451.485 -41.655 -451.085 -40.455 ;
        RECT -452.605 -45.015 -452.205 -43.815 ;
        RECT -453.105 -55.435 -452.825 -45.995 ;
        RECT -452.545 -55.155 -452.265 -45.015 ;
        RECT -451.985 -55.435 -451.705 -45.995 ;
        RECT -451.425 -55.155 -451.145 -41.655 ;
        RECT -450.365 -45.015 -449.965 -43.815 ;
        RECT -450.865 -55.435 -450.585 -45.995 ;
        RECT -450.305 -55.155 -450.025 -45.015 ;
        RECT -449.745 -55.435 -449.465 -45.995 ;
        RECT -449.185 -55.155 -448.905 -34.935 ;
        RECT -444.765 -38.295 -444.365 -37.095 ;
        RECT -447.005 -41.655 -446.605 -40.455 ;
        RECT -448.125 -45.015 -447.725 -43.815 ;
        RECT -448.625 -55.435 -448.345 -45.995 ;
        RECT -448.065 -55.155 -447.785 -45.015 ;
        RECT -447.505 -55.435 -447.225 -45.995 ;
        RECT -446.945 -55.155 -446.665 -41.655 ;
        RECT -445.885 -45.015 -445.485 -43.815 ;
        RECT -446.385 -55.435 -446.105 -45.995 ;
        RECT -445.825 -55.155 -445.545 -45.015 ;
        RECT -445.265 -55.435 -444.985 -45.995 ;
        RECT -444.705 -55.155 -444.425 -38.295 ;
        RECT -442.525 -41.655 -442.125 -40.455 ;
        RECT -443.645 -45.015 -443.245 -43.815 ;
        RECT -444.145 -55.435 -443.865 -45.995 ;
        RECT -443.585 -55.155 -443.305 -45.015 ;
        RECT -443.025 -55.435 -442.745 -45.995 ;
        RECT -442.465 -55.155 -442.185 -41.655 ;
        RECT -441.405 -45.015 -441.005 -43.815 ;
        RECT -441.905 -55.435 -441.625 -45.995 ;
        RECT -441.345 -55.155 -441.065 -45.015 ;
        RECT -440.785 -55.435 -440.505 -45.995 ;
        RECT -440.225 -55.155 -439.945 -28.215 ;
        RECT -422.365 -31.575 -421.965 -30.375 ;
        RECT -431.325 -34.935 -430.925 -33.735 ;
        RECT -435.805 -38.295 -435.405 -37.095 ;
        RECT -438.045 -41.655 -437.645 -40.455 ;
        RECT -439.165 -45.015 -438.765 -43.815 ;
        RECT -439.665 -55.435 -439.385 -45.995 ;
        RECT -439.105 -55.155 -438.825 -45.015 ;
        RECT -438.545 -55.435 -438.265 -45.995 ;
        RECT -437.985 -55.155 -437.705 -41.655 ;
        RECT -436.925 -45.015 -436.525 -43.815 ;
        RECT -437.425 -55.435 -437.145 -45.995 ;
        RECT -436.865 -55.155 -436.585 -45.015 ;
        RECT -436.305 -55.435 -436.025 -45.995 ;
        RECT -435.745 -55.155 -435.465 -38.295 ;
        RECT -433.565 -41.655 -433.165 -40.455 ;
        RECT -434.685 -45.015 -434.285 -43.815 ;
        RECT -435.185 -55.435 -434.905 -45.995 ;
        RECT -434.625 -55.155 -434.345 -45.015 ;
        RECT -434.065 -55.435 -433.785 -45.995 ;
        RECT -433.505 -55.155 -433.225 -41.655 ;
        RECT -432.445 -45.015 -432.045 -43.815 ;
        RECT -432.945 -55.435 -432.665 -45.995 ;
        RECT -432.385 -55.155 -432.105 -45.015 ;
        RECT -431.825 -55.435 -431.545 -45.995 ;
        RECT -431.265 -55.155 -430.985 -34.935 ;
        RECT -426.845 -38.295 -426.445 -37.095 ;
        RECT -429.085 -41.655 -428.685 -40.455 ;
        RECT -430.205 -45.015 -429.805 -43.815 ;
        RECT -430.705 -55.435 -430.425 -45.995 ;
        RECT -430.145 -55.155 -429.865 -45.015 ;
        RECT -429.585 -55.435 -429.305 -45.995 ;
        RECT -429.025 -55.155 -428.745 -41.655 ;
        RECT -427.965 -45.015 -427.565 -43.815 ;
        RECT -428.465 -55.435 -428.185 -45.995 ;
        RECT -427.905 -55.155 -427.625 -45.015 ;
        RECT -427.345 -55.435 -427.065 -45.995 ;
        RECT -426.785 -55.155 -426.505 -38.295 ;
        RECT -424.605 -41.655 -424.205 -40.455 ;
        RECT -425.725 -45.015 -425.325 -43.815 ;
        RECT -426.225 -55.435 -425.945 -45.995 ;
        RECT -425.665 -55.155 -425.385 -45.015 ;
        RECT -425.105 -55.435 -424.825 -45.995 ;
        RECT -424.545 -55.155 -424.265 -41.655 ;
        RECT -423.485 -45.015 -423.085 -43.815 ;
        RECT -423.985 -55.435 -423.705 -45.995 ;
        RECT -423.425 -55.155 -423.145 -45.015 ;
        RECT -422.865 -55.435 -422.585 -45.995 ;
        RECT -422.305 -55.155 -422.025 -31.575 ;
        RECT -413.405 -34.935 -413.005 -33.735 ;
        RECT -417.885 -38.295 -417.485 -37.095 ;
        RECT -420.125 -41.655 -419.725 -40.455 ;
        RECT -421.245 -45.015 -420.845 -43.815 ;
        RECT -421.745 -55.435 -421.465 -45.995 ;
        RECT -421.185 -55.155 -420.905 -45.015 ;
        RECT -420.625 -55.435 -420.345 -45.995 ;
        RECT -420.065 -55.155 -419.785 -41.655 ;
        RECT -419.005 -45.015 -418.605 -43.815 ;
        RECT -419.505 -55.435 -419.225 -45.995 ;
        RECT -418.945 -55.155 -418.665 -45.015 ;
        RECT -418.385 -55.435 -418.105 -45.995 ;
        RECT -417.825 -55.155 -417.545 -38.295 ;
        RECT -415.645 -41.655 -415.245 -40.455 ;
        RECT -416.765 -45.015 -416.365 -43.815 ;
        RECT -417.265 -55.435 -416.985 -45.995 ;
        RECT -416.705 -55.155 -416.425 -45.015 ;
        RECT -416.145 -55.435 -415.865 -45.995 ;
        RECT -415.585 -55.155 -415.305 -41.655 ;
        RECT -414.525 -45.015 -414.125 -43.815 ;
        RECT -415.025 -55.435 -414.745 -45.995 ;
        RECT -414.465 -55.155 -414.185 -45.015 ;
        RECT -413.905 -55.435 -413.625 -45.995 ;
        RECT -413.345 -55.155 -413.065 -34.935 ;
        RECT -408.925 -38.295 -408.525 -37.095 ;
        RECT -411.165 -41.655 -410.765 -40.455 ;
        RECT -412.285 -45.015 -411.885 -43.815 ;
        RECT -412.785 -55.435 -412.505 -45.995 ;
        RECT -412.225 -55.155 -411.945 -45.015 ;
        RECT -411.665 -55.435 -411.385 -45.995 ;
        RECT -411.105 -55.155 -410.825 -41.655 ;
        RECT -410.045 -45.015 -409.645 -43.815 ;
        RECT -410.545 -55.435 -410.265 -45.995 ;
        RECT -409.985 -55.155 -409.705 -45.015 ;
        RECT -409.425 -55.435 -409.145 -45.995 ;
        RECT -408.865 -55.155 -408.585 -38.295 ;
        RECT -406.685 -41.655 -406.285 -40.455 ;
        RECT -407.805 -45.015 -407.405 -43.815 ;
        RECT -408.305 -55.435 -408.025 -45.995 ;
        RECT -407.745 -55.155 -407.465 -45.015 ;
        RECT -407.185 -55.435 -406.905 -45.995 ;
        RECT -406.625 -55.155 -406.345 -41.655 ;
        RECT -405.565 -45.015 -405.165 -43.815 ;
        RECT -406.065 -55.435 -405.785 -45.995 ;
        RECT -405.505 -55.155 -405.225 -45.015 ;
        RECT -404.945 -55.435 -404.665 -45.995 ;
        RECT -404.385 -55.155 -404.105 -24.855 ;
        RECT -368.605 -28.215 -368.205 -27.015 ;
        RECT -386.525 -31.575 -386.125 -30.375 ;
        RECT -395.485 -34.935 -395.085 -33.735 ;
        RECT -399.965 -38.295 -399.565 -37.095 ;
        RECT -402.205 -41.655 -401.805 -40.455 ;
        RECT -403.325 -45.015 -402.925 -43.815 ;
        RECT -403.825 -55.435 -403.545 -45.995 ;
        RECT -403.265 -55.155 -402.985 -45.015 ;
        RECT -402.705 -55.435 -402.425 -45.995 ;
        RECT -402.145 -55.155 -401.865 -41.655 ;
        RECT -401.085 -45.015 -400.685 -43.815 ;
        RECT -401.585 -55.435 -401.305 -45.995 ;
        RECT -401.025 -55.155 -400.745 -45.015 ;
        RECT -400.465 -55.435 -400.185 -45.995 ;
        RECT -399.905 -55.155 -399.625 -38.295 ;
        RECT -397.725 -41.655 -397.325 -40.455 ;
        RECT -398.845 -45.015 -398.445 -43.815 ;
        RECT -399.345 -55.435 -399.065 -45.995 ;
        RECT -398.785 -55.155 -398.505 -45.015 ;
        RECT -398.225 -55.435 -397.945 -45.995 ;
        RECT -397.665 -55.155 -397.385 -41.655 ;
        RECT -396.605 -45.015 -396.205 -43.815 ;
        RECT -397.105 -55.435 -396.825 -45.995 ;
        RECT -396.545 -55.155 -396.265 -45.015 ;
        RECT -395.985 -55.435 -395.705 -45.995 ;
        RECT -395.425 -55.155 -395.145 -34.935 ;
        RECT -391.005 -38.295 -390.605 -37.095 ;
        RECT -393.245 -41.655 -392.845 -40.455 ;
        RECT -394.365 -45.015 -393.965 -43.815 ;
        RECT -394.865 -55.435 -394.585 -45.995 ;
        RECT -394.305 -55.155 -394.025 -45.015 ;
        RECT -393.745 -55.435 -393.465 -45.995 ;
        RECT -393.185 -55.155 -392.905 -41.655 ;
        RECT -392.125 -45.015 -391.725 -43.815 ;
        RECT -392.625 -55.435 -392.345 -45.995 ;
        RECT -392.065 -55.155 -391.785 -45.015 ;
        RECT -391.505 -55.435 -391.225 -45.995 ;
        RECT -390.945 -55.155 -390.665 -38.295 ;
        RECT -388.765 -41.655 -388.365 -40.455 ;
        RECT -389.885 -45.015 -389.485 -43.815 ;
        RECT -390.385 -55.435 -390.105 -45.995 ;
        RECT -389.825 -55.155 -389.545 -45.015 ;
        RECT -389.265 -55.435 -388.985 -45.995 ;
        RECT -388.705 -55.155 -388.425 -41.655 ;
        RECT -387.645 -45.015 -387.245 -43.815 ;
        RECT -388.145 -55.435 -387.865 -45.995 ;
        RECT -387.585 -55.155 -387.305 -45.015 ;
        RECT -387.025 -55.435 -386.745 -45.995 ;
        RECT -386.465 -55.155 -386.185 -31.575 ;
        RECT -377.565 -34.935 -377.165 -33.735 ;
        RECT -382.045 -38.295 -381.645 -37.095 ;
        RECT -384.285 -41.655 -383.885 -40.455 ;
        RECT -385.405 -45.015 -385.005 -43.815 ;
        RECT -385.905 -55.435 -385.625 -45.995 ;
        RECT -385.345 -55.155 -385.065 -45.015 ;
        RECT -384.785 -55.435 -384.505 -45.995 ;
        RECT -384.225 -55.155 -383.945 -41.655 ;
        RECT -383.165 -45.015 -382.765 -43.815 ;
        RECT -383.665 -55.435 -383.385 -45.995 ;
        RECT -383.105 -55.155 -382.825 -45.015 ;
        RECT -382.545 -55.435 -382.265 -45.995 ;
        RECT -381.985 -55.155 -381.705 -38.295 ;
        RECT -379.805 -41.655 -379.405 -40.455 ;
        RECT -380.925 -45.015 -380.525 -43.815 ;
        RECT -381.425 -55.435 -381.145 -45.995 ;
        RECT -380.865 -55.155 -380.585 -45.015 ;
        RECT -380.305 -55.435 -380.025 -45.995 ;
        RECT -379.745 -55.155 -379.465 -41.655 ;
        RECT -378.685 -45.015 -378.285 -43.815 ;
        RECT -379.185 -55.435 -378.905 -45.995 ;
        RECT -378.625 -55.155 -378.345 -45.015 ;
        RECT -378.065 -55.435 -377.785 -45.995 ;
        RECT -377.505 -55.155 -377.225 -34.935 ;
        RECT -373.085 -38.295 -372.685 -37.095 ;
        RECT -375.325 -41.655 -374.925 -40.455 ;
        RECT -376.445 -45.015 -376.045 -43.815 ;
        RECT -376.945 -55.435 -376.665 -45.995 ;
        RECT -376.385 -55.155 -376.105 -45.015 ;
        RECT -375.825 -55.435 -375.545 -45.995 ;
        RECT -375.265 -55.155 -374.985 -41.655 ;
        RECT -374.205 -45.015 -373.805 -43.815 ;
        RECT -374.705 -55.435 -374.425 -45.995 ;
        RECT -374.145 -55.155 -373.865 -45.015 ;
        RECT -373.585 -55.435 -373.305 -45.995 ;
        RECT -373.025 -55.155 -372.745 -38.295 ;
        RECT -370.845 -41.655 -370.445 -40.455 ;
        RECT -371.965 -45.015 -371.565 -43.815 ;
        RECT -372.465 -55.435 -372.185 -45.995 ;
        RECT -371.905 -55.155 -371.625 -45.015 ;
        RECT -371.345 -55.435 -371.065 -45.995 ;
        RECT -370.785 -55.155 -370.505 -41.655 ;
        RECT -369.725 -45.015 -369.325 -43.815 ;
        RECT -370.225 -55.435 -369.945 -45.995 ;
        RECT -369.665 -55.155 -369.385 -45.015 ;
        RECT -369.105 -55.435 -368.825 -45.995 ;
        RECT -368.545 -55.155 -368.265 -28.215 ;
        RECT -350.685 -31.575 -350.285 -30.375 ;
        RECT -359.645 -34.935 -359.245 -33.735 ;
        RECT -364.125 -38.295 -363.725 -37.095 ;
        RECT -366.365 -41.655 -365.965 -40.455 ;
        RECT -367.485 -45.015 -367.085 -43.815 ;
        RECT -367.985 -55.435 -367.705 -45.995 ;
        RECT -367.425 -55.155 -367.145 -45.015 ;
        RECT -366.865 -55.435 -366.585 -45.995 ;
        RECT -366.305 -55.155 -366.025 -41.655 ;
        RECT -365.245 -45.015 -364.845 -43.815 ;
        RECT -365.745 -55.435 -365.465 -45.995 ;
        RECT -365.185 -55.155 -364.905 -45.015 ;
        RECT -364.625 -55.435 -364.345 -45.995 ;
        RECT -364.065 -55.155 -363.785 -38.295 ;
        RECT -361.885 -41.655 -361.485 -40.455 ;
        RECT -363.005 -45.015 -362.605 -43.815 ;
        RECT -363.505 -55.435 -363.225 -45.995 ;
        RECT -362.945 -55.155 -362.665 -45.015 ;
        RECT -362.385 -55.435 -362.105 -45.995 ;
        RECT -361.825 -55.155 -361.545 -41.655 ;
        RECT -360.765 -45.015 -360.365 -43.815 ;
        RECT -361.265 -55.435 -360.985 -45.995 ;
        RECT -360.705 -55.155 -360.425 -45.015 ;
        RECT -360.145 -55.435 -359.865 -45.995 ;
        RECT -359.585 -55.155 -359.305 -34.935 ;
        RECT -355.165 -38.295 -354.765 -37.095 ;
        RECT -357.405 -41.655 -357.005 -40.455 ;
        RECT -358.525 -45.015 -358.125 -43.815 ;
        RECT -359.025 -55.435 -358.745 -45.995 ;
        RECT -358.465 -55.155 -358.185 -45.015 ;
        RECT -357.905 -55.435 -357.625 -45.995 ;
        RECT -357.345 -55.155 -357.065 -41.655 ;
        RECT -356.285 -45.015 -355.885 -43.815 ;
        RECT -356.785 -55.435 -356.505 -45.995 ;
        RECT -356.225 -55.155 -355.945 -45.015 ;
        RECT -355.665 -55.435 -355.385 -45.995 ;
        RECT -355.105 -55.155 -354.825 -38.295 ;
        RECT -352.925 -41.655 -352.525 -40.455 ;
        RECT -354.045 -45.015 -353.645 -43.815 ;
        RECT -354.545 -55.435 -354.265 -45.995 ;
        RECT -353.985 -55.155 -353.705 -45.015 ;
        RECT -353.425 -55.435 -353.145 -45.995 ;
        RECT -352.865 -55.155 -352.585 -41.655 ;
        RECT -351.805 -45.015 -351.405 -43.815 ;
        RECT -352.305 -55.435 -352.025 -45.995 ;
        RECT -351.745 -55.155 -351.465 -45.015 ;
        RECT -351.185 -55.435 -350.905 -45.995 ;
        RECT -350.625 -55.155 -350.345 -31.575 ;
        RECT -341.725 -34.935 -341.325 -33.735 ;
        RECT -346.205 -38.295 -345.805 -37.095 ;
        RECT -348.445 -41.655 -348.045 -40.455 ;
        RECT -349.565 -45.015 -349.165 -43.815 ;
        RECT -350.065 -55.435 -349.785 -45.995 ;
        RECT -349.505 -55.155 -349.225 -45.015 ;
        RECT -348.945 -55.435 -348.665 -45.995 ;
        RECT -348.385 -55.155 -348.105 -41.655 ;
        RECT -347.325 -45.015 -346.925 -43.815 ;
        RECT -347.825 -55.435 -347.545 -45.995 ;
        RECT -347.265 -55.155 -346.985 -45.015 ;
        RECT -346.705 -55.435 -346.425 -45.995 ;
        RECT -346.145 -55.155 -345.865 -38.295 ;
        RECT -343.965 -41.655 -343.565 -40.455 ;
        RECT -345.085 -45.015 -344.685 -43.815 ;
        RECT -345.585 -55.435 -345.305 -45.995 ;
        RECT -345.025 -55.155 -344.745 -45.015 ;
        RECT -344.465 -55.435 -344.185 -45.995 ;
        RECT -343.905 -55.155 -343.625 -41.655 ;
        RECT -342.845 -45.015 -342.445 -43.815 ;
        RECT -343.345 -55.435 -343.065 -45.995 ;
        RECT -342.785 -55.155 -342.505 -45.015 ;
        RECT -342.225 -55.435 -341.945 -45.995 ;
        RECT -341.665 -55.155 -341.385 -34.935 ;
        RECT -337.245 -38.295 -336.845 -37.095 ;
        RECT -339.485 -41.655 -339.085 -40.455 ;
        RECT -340.605 -45.015 -340.205 -43.815 ;
        RECT -341.105 -55.435 -340.825 -45.995 ;
        RECT -340.545 -55.155 -340.265 -45.015 ;
        RECT -339.985 -55.435 -339.705 -45.995 ;
        RECT -339.425 -55.155 -339.145 -41.655 ;
        RECT -338.365 -45.015 -337.965 -43.815 ;
        RECT -338.865 -55.435 -338.585 -45.995 ;
        RECT -338.305 -55.155 -338.025 -45.015 ;
        RECT -337.745 -55.435 -337.465 -45.995 ;
        RECT -337.185 -55.155 -336.905 -38.295 ;
        RECT -335.005 -41.655 -334.605 -40.455 ;
        RECT -336.125 -45.015 -335.725 -43.815 ;
        RECT -336.625 -55.435 -336.345 -45.995 ;
        RECT -336.065 -55.155 -335.785 -45.015 ;
        RECT -335.505 -55.435 -335.225 -45.995 ;
        RECT -334.945 -55.155 -334.665 -41.655 ;
        RECT -333.885 -45.015 -333.485 -43.815 ;
        RECT -334.385 -55.435 -334.105 -45.995 ;
        RECT -333.825 -55.155 -333.545 -45.015 ;
        RECT -333.265 -55.435 -332.985 -45.995 ;
        RECT -332.705 -55.155 -332.425 -21.495 ;
        RECT -261.085 -24.855 -260.685 -23.655 ;
        RECT -296.925 -28.215 -296.525 -27.015 ;
        RECT -314.845 -31.575 -314.445 -30.375 ;
        RECT -323.805 -34.935 -323.405 -33.735 ;
        RECT -328.285 -38.295 -327.885 -37.095 ;
        RECT -330.525 -41.655 -330.125 -40.455 ;
        RECT -331.645 -45.015 -331.245 -43.815 ;
        RECT -332.145 -55.435 -331.865 -45.995 ;
        RECT -331.585 -55.155 -331.305 -45.015 ;
        RECT -331.025 -55.435 -330.745 -45.995 ;
        RECT -330.465 -55.155 -330.185 -41.655 ;
        RECT -329.405 -45.015 -329.005 -43.815 ;
        RECT -329.905 -55.435 -329.625 -45.995 ;
        RECT -329.345 -55.155 -329.065 -45.015 ;
        RECT -328.785 -55.435 -328.505 -45.995 ;
        RECT -328.225 -55.155 -327.945 -38.295 ;
        RECT -326.045 -41.655 -325.645 -40.455 ;
        RECT -327.165 -45.015 -326.765 -43.815 ;
        RECT -327.665 -55.435 -327.385 -45.995 ;
        RECT -327.105 -55.155 -326.825 -45.015 ;
        RECT -326.545 -55.435 -326.265 -45.995 ;
        RECT -325.985 -55.155 -325.705 -41.655 ;
        RECT -324.925 -45.015 -324.525 -43.815 ;
        RECT -325.425 -55.435 -325.145 -45.995 ;
        RECT -324.865 -55.155 -324.585 -45.015 ;
        RECT -324.305 -55.435 -324.025 -45.995 ;
        RECT -323.745 -55.155 -323.465 -34.935 ;
        RECT -319.325 -38.295 -318.925 -37.095 ;
        RECT -321.565 -41.655 -321.165 -40.455 ;
        RECT -322.685 -45.015 -322.285 -43.815 ;
        RECT -323.185 -55.435 -322.905 -45.995 ;
        RECT -322.625 -55.155 -322.345 -45.015 ;
        RECT -322.065 -55.435 -321.785 -45.995 ;
        RECT -321.505 -55.155 -321.225 -41.655 ;
        RECT -320.445 -45.015 -320.045 -43.815 ;
        RECT -320.945 -55.435 -320.665 -45.995 ;
        RECT -320.385 -55.155 -320.105 -45.015 ;
        RECT -319.825 -55.435 -319.545 -45.995 ;
        RECT -319.265 -55.155 -318.985 -38.295 ;
        RECT -317.085 -41.655 -316.685 -40.455 ;
        RECT -318.205 -45.015 -317.805 -43.815 ;
        RECT -318.705 -55.435 -318.425 -45.995 ;
        RECT -318.145 -55.155 -317.865 -45.015 ;
        RECT -317.585 -55.435 -317.305 -45.995 ;
        RECT -317.025 -55.155 -316.745 -41.655 ;
        RECT -315.965 -45.015 -315.565 -43.815 ;
        RECT -316.465 -55.435 -316.185 -45.995 ;
        RECT -315.905 -55.155 -315.625 -45.015 ;
        RECT -315.345 -55.435 -315.065 -45.995 ;
        RECT -314.785 -55.155 -314.505 -31.575 ;
        RECT -305.885 -34.935 -305.485 -33.735 ;
        RECT -310.365 -38.295 -309.965 -37.095 ;
        RECT -312.605 -41.655 -312.205 -40.455 ;
        RECT -313.725 -45.015 -313.325 -43.815 ;
        RECT -314.225 -55.435 -313.945 -45.995 ;
        RECT -313.665 -55.155 -313.385 -45.015 ;
        RECT -313.105 -55.435 -312.825 -45.995 ;
        RECT -312.545 -55.155 -312.265 -41.655 ;
        RECT -311.485 -45.015 -311.085 -43.815 ;
        RECT -311.985 -55.435 -311.705 -45.995 ;
        RECT -311.425 -55.155 -311.145 -45.015 ;
        RECT -310.865 -55.435 -310.585 -45.995 ;
        RECT -310.305 -55.155 -310.025 -38.295 ;
        RECT -308.125 -41.655 -307.725 -40.455 ;
        RECT -309.245 -45.015 -308.845 -43.815 ;
        RECT -309.745 -55.435 -309.465 -45.995 ;
        RECT -309.185 -55.155 -308.905 -45.015 ;
        RECT -308.625 -55.435 -308.345 -45.995 ;
        RECT -308.065 -55.155 -307.785 -41.655 ;
        RECT -307.005 -45.015 -306.605 -43.815 ;
        RECT -307.505 -55.435 -307.225 -45.995 ;
        RECT -306.945 -55.155 -306.665 -45.015 ;
        RECT -306.385 -55.435 -306.105 -45.995 ;
        RECT -305.825 -55.155 -305.545 -34.935 ;
        RECT -301.405 -38.295 -301.005 -37.095 ;
        RECT -303.645 -41.655 -303.245 -40.455 ;
        RECT -304.765 -45.015 -304.365 -43.815 ;
        RECT -305.265 -55.435 -304.985 -45.995 ;
        RECT -304.705 -55.155 -304.425 -45.015 ;
        RECT -304.145 -55.435 -303.865 -45.995 ;
        RECT -303.585 -55.155 -303.305 -41.655 ;
        RECT -302.525 -45.015 -302.125 -43.815 ;
        RECT -303.025 -55.435 -302.745 -45.995 ;
        RECT -302.465 -55.155 -302.185 -45.015 ;
        RECT -301.905 -55.435 -301.625 -45.995 ;
        RECT -301.345 -55.155 -301.065 -38.295 ;
        RECT -299.165 -41.655 -298.765 -40.455 ;
        RECT -300.285 -45.015 -299.885 -43.815 ;
        RECT -300.785 -55.435 -300.505 -45.995 ;
        RECT -300.225 -55.155 -299.945 -45.015 ;
        RECT -299.665 -55.435 -299.385 -45.995 ;
        RECT -299.105 -55.155 -298.825 -41.655 ;
        RECT -298.045 -45.015 -297.645 -43.815 ;
        RECT -298.545 -55.435 -298.265 -45.995 ;
        RECT -297.985 -55.155 -297.705 -45.015 ;
        RECT -297.425 -55.435 -297.145 -45.995 ;
        RECT -296.865 -55.155 -296.585 -28.215 ;
        RECT -279.005 -31.575 -278.605 -30.375 ;
        RECT -287.965 -34.935 -287.565 -33.735 ;
        RECT -292.445 -38.295 -292.045 -37.095 ;
        RECT -294.685 -41.655 -294.285 -40.455 ;
        RECT -295.805 -45.015 -295.405 -43.815 ;
        RECT -296.305 -55.435 -296.025 -45.995 ;
        RECT -295.745 -55.155 -295.465 -45.015 ;
        RECT -295.185 -55.435 -294.905 -45.995 ;
        RECT -294.625 -55.155 -294.345 -41.655 ;
        RECT -293.565 -45.015 -293.165 -43.815 ;
        RECT -294.065 -55.435 -293.785 -45.995 ;
        RECT -293.505 -55.155 -293.225 -45.015 ;
        RECT -292.945 -55.435 -292.665 -45.995 ;
        RECT -292.385 -55.155 -292.105 -38.295 ;
        RECT -290.205 -41.655 -289.805 -40.455 ;
        RECT -291.325 -45.015 -290.925 -43.815 ;
        RECT -291.825 -55.435 -291.545 -45.995 ;
        RECT -291.265 -55.155 -290.985 -45.015 ;
        RECT -290.705 -55.435 -290.425 -45.995 ;
        RECT -290.145 -55.155 -289.865 -41.655 ;
        RECT -289.085 -45.015 -288.685 -43.815 ;
        RECT -289.585 -55.435 -289.305 -45.995 ;
        RECT -289.025 -55.155 -288.745 -45.015 ;
        RECT -288.465 -55.435 -288.185 -45.995 ;
        RECT -287.905 -55.155 -287.625 -34.935 ;
        RECT -283.485 -38.295 -283.085 -37.095 ;
        RECT -285.725 -41.655 -285.325 -40.455 ;
        RECT -286.845 -45.015 -286.445 -43.815 ;
        RECT -287.345 -55.435 -287.065 -45.995 ;
        RECT -286.785 -55.155 -286.505 -45.015 ;
        RECT -286.225 -55.435 -285.945 -45.995 ;
        RECT -285.665 -55.155 -285.385 -41.655 ;
        RECT -284.605 -45.015 -284.205 -43.815 ;
        RECT -285.105 -55.435 -284.825 -45.995 ;
        RECT -284.545 -55.155 -284.265 -45.015 ;
        RECT -283.985 -55.435 -283.705 -45.995 ;
        RECT -283.425 -55.155 -283.145 -38.295 ;
        RECT -281.245 -41.655 -280.845 -40.455 ;
        RECT -282.365 -45.015 -281.965 -43.815 ;
        RECT -282.865 -55.435 -282.585 -45.995 ;
        RECT -282.305 -55.155 -282.025 -45.015 ;
        RECT -281.745 -55.435 -281.465 -45.995 ;
        RECT -281.185 -55.155 -280.905 -41.655 ;
        RECT -280.125 -45.015 -279.725 -43.815 ;
        RECT -280.625 -55.435 -280.345 -45.995 ;
        RECT -280.065 -55.155 -279.785 -45.015 ;
        RECT -279.505 -55.435 -279.225 -45.995 ;
        RECT -278.945 -55.155 -278.665 -31.575 ;
        RECT -270.045 -34.935 -269.645 -33.735 ;
        RECT -274.525 -38.295 -274.125 -37.095 ;
        RECT -276.765 -41.655 -276.365 -40.455 ;
        RECT -277.885 -45.015 -277.485 -43.815 ;
        RECT -278.385 -55.435 -278.105 -45.995 ;
        RECT -277.825 -55.155 -277.545 -45.015 ;
        RECT -277.265 -55.435 -276.985 -45.995 ;
        RECT -276.705 -55.155 -276.425 -41.655 ;
        RECT -275.645 -45.015 -275.245 -43.815 ;
        RECT -276.145 -55.435 -275.865 -45.995 ;
        RECT -275.585 -55.155 -275.305 -45.015 ;
        RECT -275.025 -55.435 -274.745 -45.995 ;
        RECT -274.465 -55.155 -274.185 -38.295 ;
        RECT -272.285 -41.655 -271.885 -40.455 ;
        RECT -273.405 -45.015 -273.005 -43.815 ;
        RECT -273.905 -55.435 -273.625 -45.995 ;
        RECT -273.345 -55.155 -273.065 -45.015 ;
        RECT -272.785 -55.435 -272.505 -45.995 ;
        RECT -272.225 -55.155 -271.945 -41.655 ;
        RECT -271.165 -45.015 -270.765 -43.815 ;
        RECT -271.665 -55.435 -271.385 -45.995 ;
        RECT -271.105 -55.155 -270.825 -45.015 ;
        RECT -270.545 -55.435 -270.265 -45.995 ;
        RECT -269.985 -55.155 -269.705 -34.935 ;
        RECT -265.565 -38.295 -265.165 -37.095 ;
        RECT -267.805 -41.655 -267.405 -40.455 ;
        RECT -268.925 -45.015 -268.525 -43.815 ;
        RECT -269.425 -55.435 -269.145 -45.995 ;
        RECT -268.865 -55.155 -268.585 -45.015 ;
        RECT -268.305 -55.435 -268.025 -45.995 ;
        RECT -267.745 -55.155 -267.465 -41.655 ;
        RECT -266.685 -45.015 -266.285 -43.815 ;
        RECT -267.185 -55.435 -266.905 -45.995 ;
        RECT -266.625 -55.155 -266.345 -45.015 ;
        RECT -266.065 -55.435 -265.785 -45.995 ;
        RECT -265.505 -55.155 -265.225 -38.295 ;
        RECT -263.325 -41.655 -262.925 -40.455 ;
        RECT -264.445 -45.015 -264.045 -43.815 ;
        RECT -264.945 -55.435 -264.665 -45.995 ;
        RECT -264.385 -55.155 -264.105 -45.015 ;
        RECT -263.825 -55.435 -263.545 -45.995 ;
        RECT -263.265 -55.155 -262.985 -41.655 ;
        RECT -262.205 -45.015 -261.805 -43.815 ;
        RECT -262.705 -55.435 -262.425 -45.995 ;
        RECT -262.145 -55.155 -261.865 -45.015 ;
        RECT -261.585 -55.435 -261.305 -45.995 ;
        RECT -261.025 -55.155 -260.745 -24.855 ;
        RECT -225.245 -28.215 -224.845 -27.015 ;
        RECT -243.165 -31.575 -242.765 -30.375 ;
        RECT -252.125 -34.935 -251.725 -33.735 ;
        RECT -256.605 -38.295 -256.205 -37.095 ;
        RECT -258.845 -41.655 -258.445 -40.455 ;
        RECT -259.965 -45.015 -259.565 -43.815 ;
        RECT -260.465 -55.435 -260.185 -45.995 ;
        RECT -259.905 -55.155 -259.625 -45.015 ;
        RECT -259.345 -55.435 -259.065 -45.995 ;
        RECT -258.785 -55.155 -258.505 -41.655 ;
        RECT -257.725 -45.015 -257.325 -43.815 ;
        RECT -258.225 -55.435 -257.945 -45.995 ;
        RECT -257.665 -55.155 -257.385 -45.015 ;
        RECT -257.105 -55.435 -256.825 -45.995 ;
        RECT -256.545 -55.155 -256.265 -38.295 ;
        RECT -254.365 -41.655 -253.965 -40.455 ;
        RECT -255.485 -45.015 -255.085 -43.815 ;
        RECT -255.985 -55.435 -255.705 -45.995 ;
        RECT -255.425 -55.155 -255.145 -45.015 ;
        RECT -254.865 -55.435 -254.585 -45.995 ;
        RECT -254.305 -55.155 -254.025 -41.655 ;
        RECT -253.245 -45.015 -252.845 -43.815 ;
        RECT -253.745 -55.435 -253.465 -45.995 ;
        RECT -253.185 -55.155 -252.905 -45.015 ;
        RECT -252.625 -55.435 -252.345 -45.995 ;
        RECT -252.065 -55.155 -251.785 -34.935 ;
        RECT -247.645 -38.295 -247.245 -37.095 ;
        RECT -249.885 -41.655 -249.485 -40.455 ;
        RECT -251.005 -45.015 -250.605 -43.815 ;
        RECT -251.505 -55.435 -251.225 -45.995 ;
        RECT -250.945 -55.155 -250.665 -45.015 ;
        RECT -250.385 -55.435 -250.105 -45.995 ;
        RECT -249.825 -55.155 -249.545 -41.655 ;
        RECT -248.765 -45.015 -248.365 -43.815 ;
        RECT -249.265 -55.435 -248.985 -45.995 ;
        RECT -248.705 -55.155 -248.425 -45.015 ;
        RECT -248.145 -55.435 -247.865 -45.995 ;
        RECT -247.585 -55.155 -247.305 -38.295 ;
        RECT -245.405 -41.655 -245.005 -40.455 ;
        RECT -246.525 -45.015 -246.125 -43.815 ;
        RECT -247.025 -55.435 -246.745 -45.995 ;
        RECT -246.465 -55.155 -246.185 -45.015 ;
        RECT -245.905 -55.435 -245.625 -45.995 ;
        RECT -245.345 -55.155 -245.065 -41.655 ;
        RECT -244.285 -45.015 -243.885 -43.815 ;
        RECT -244.785 -55.435 -244.505 -45.995 ;
        RECT -244.225 -55.155 -243.945 -45.015 ;
        RECT -243.665 -55.435 -243.385 -45.995 ;
        RECT -243.105 -55.155 -242.825 -31.575 ;
        RECT -234.205 -34.935 -233.805 -33.735 ;
        RECT -238.685 -38.295 -238.285 -37.095 ;
        RECT -240.925 -41.655 -240.525 -40.455 ;
        RECT -242.045 -45.015 -241.645 -43.815 ;
        RECT -242.545 -55.435 -242.265 -45.995 ;
        RECT -241.985 -55.155 -241.705 -45.015 ;
        RECT -241.425 -55.435 -241.145 -45.995 ;
        RECT -240.865 -55.155 -240.585 -41.655 ;
        RECT -239.805 -45.015 -239.405 -43.815 ;
        RECT -240.305 -55.435 -240.025 -45.995 ;
        RECT -239.745 -55.155 -239.465 -45.015 ;
        RECT -239.185 -55.435 -238.905 -45.995 ;
        RECT -238.625 -55.155 -238.345 -38.295 ;
        RECT -236.445 -41.655 -236.045 -40.455 ;
        RECT -237.565 -45.015 -237.165 -43.815 ;
        RECT -238.065 -55.435 -237.785 -45.995 ;
        RECT -237.505 -55.155 -237.225 -45.015 ;
        RECT -236.945 -55.435 -236.665 -45.995 ;
        RECT -236.385 -55.155 -236.105 -41.655 ;
        RECT -235.325 -45.015 -234.925 -43.815 ;
        RECT -235.825 -55.435 -235.545 -45.995 ;
        RECT -235.265 -55.155 -234.985 -45.015 ;
        RECT -234.705 -55.435 -234.425 -45.995 ;
        RECT -234.145 -55.155 -233.865 -34.935 ;
        RECT -229.725 -38.295 -229.325 -37.095 ;
        RECT -231.965 -41.655 -231.565 -40.455 ;
        RECT -233.085 -45.015 -232.685 -43.815 ;
        RECT -233.585 -55.435 -233.305 -45.995 ;
        RECT -233.025 -55.155 -232.745 -45.015 ;
        RECT -232.465 -55.435 -232.185 -45.995 ;
        RECT -231.905 -55.155 -231.625 -41.655 ;
        RECT -230.845 -45.015 -230.445 -43.815 ;
        RECT -231.345 -55.435 -231.065 -45.995 ;
        RECT -230.785 -55.155 -230.505 -45.015 ;
        RECT -230.225 -55.435 -229.945 -45.995 ;
        RECT -229.665 -55.155 -229.385 -38.295 ;
        RECT -227.485 -41.655 -227.085 -40.455 ;
        RECT -228.605 -45.015 -228.205 -43.815 ;
        RECT -229.105 -55.435 -228.825 -45.995 ;
        RECT -228.545 -55.155 -228.265 -45.015 ;
        RECT -227.985 -55.435 -227.705 -45.995 ;
        RECT -227.425 -55.155 -227.145 -41.655 ;
        RECT -226.365 -45.015 -225.965 -43.815 ;
        RECT -226.865 -55.435 -226.585 -45.995 ;
        RECT -226.305 -55.155 -226.025 -45.015 ;
        RECT -225.745 -55.435 -225.465 -45.995 ;
        RECT -225.185 -55.155 -224.905 -28.215 ;
        RECT -207.325 -31.575 -206.925 -30.375 ;
        RECT -216.285 -34.935 -215.885 -33.735 ;
        RECT -220.765 -38.295 -220.365 -37.095 ;
        RECT -223.005 -41.655 -222.605 -40.455 ;
        RECT -224.125 -45.015 -223.725 -43.815 ;
        RECT -224.625 -55.435 -224.345 -45.995 ;
        RECT -224.065 -55.155 -223.785 -45.015 ;
        RECT -223.505 -55.435 -223.225 -45.995 ;
        RECT -222.945 -55.155 -222.665 -41.655 ;
        RECT -221.885 -45.015 -221.485 -43.815 ;
        RECT -222.385 -55.435 -222.105 -45.995 ;
        RECT -221.825 -55.155 -221.545 -45.015 ;
        RECT -221.265 -55.435 -220.985 -45.995 ;
        RECT -220.705 -55.155 -220.425 -38.295 ;
        RECT -218.525 -41.655 -218.125 -40.455 ;
        RECT -219.645 -45.015 -219.245 -43.815 ;
        RECT -220.145 -55.435 -219.865 -45.995 ;
        RECT -219.585 -55.155 -219.305 -45.015 ;
        RECT -219.025 -55.435 -218.745 -45.995 ;
        RECT -218.465 -55.155 -218.185 -41.655 ;
        RECT -217.405 -45.015 -217.005 -43.815 ;
        RECT -217.905 -55.435 -217.625 -45.995 ;
        RECT -217.345 -55.155 -217.065 -45.015 ;
        RECT -216.785 -55.435 -216.505 -45.995 ;
        RECT -216.225 -55.155 -215.945 -34.935 ;
        RECT -211.805 -38.295 -211.405 -37.095 ;
        RECT -214.045 -41.655 -213.645 -40.455 ;
        RECT -215.165 -45.015 -214.765 -43.815 ;
        RECT -215.665 -55.435 -215.385 -45.995 ;
        RECT -215.105 -55.155 -214.825 -45.015 ;
        RECT -214.545 -55.435 -214.265 -45.995 ;
        RECT -213.985 -55.155 -213.705 -41.655 ;
        RECT -212.925 -45.015 -212.525 -43.815 ;
        RECT -213.425 -55.435 -213.145 -45.995 ;
        RECT -212.865 -55.155 -212.585 -45.015 ;
        RECT -212.305 -55.435 -212.025 -45.995 ;
        RECT -211.745 -55.155 -211.465 -38.295 ;
        RECT -209.565 -41.655 -209.165 -40.455 ;
        RECT -210.685 -45.015 -210.285 -43.815 ;
        RECT -211.185 -55.435 -210.905 -45.995 ;
        RECT -210.625 -55.155 -210.345 -45.015 ;
        RECT -210.065 -55.435 -209.785 -45.995 ;
        RECT -209.505 -55.155 -209.225 -41.655 ;
        RECT -208.445 -45.015 -208.045 -43.815 ;
        RECT -208.945 -55.435 -208.665 -45.995 ;
        RECT -208.385 -55.155 -208.105 -45.015 ;
        RECT -207.825 -55.435 -207.545 -45.995 ;
        RECT -207.265 -55.155 -206.985 -31.575 ;
        RECT -198.365 -34.935 -197.965 -33.735 ;
        RECT -202.845 -38.295 -202.445 -37.095 ;
        RECT -205.085 -41.655 -204.685 -40.455 ;
        RECT -206.205 -45.015 -205.805 -43.815 ;
        RECT -206.705 -55.435 -206.425 -45.995 ;
        RECT -206.145 -55.155 -205.865 -45.015 ;
        RECT -205.585 -55.435 -205.305 -45.995 ;
        RECT -205.025 -55.155 -204.745 -41.655 ;
        RECT -203.965 -45.015 -203.565 -43.815 ;
        RECT -204.465 -55.435 -204.185 -45.995 ;
        RECT -203.905 -55.155 -203.625 -45.015 ;
        RECT -203.345 -55.435 -203.065 -45.995 ;
        RECT -202.785 -55.155 -202.505 -38.295 ;
        RECT -200.605 -41.655 -200.205 -40.455 ;
        RECT -201.725 -45.015 -201.325 -43.815 ;
        RECT -202.225 -55.435 -201.945 -45.995 ;
        RECT -201.665 -55.155 -201.385 -45.015 ;
        RECT -201.105 -55.435 -200.825 -45.995 ;
        RECT -200.545 -55.155 -200.265 -41.655 ;
        RECT -199.485 -45.015 -199.085 -43.815 ;
        RECT -199.985 -55.435 -199.705 -45.995 ;
        RECT -199.425 -55.155 -199.145 -45.015 ;
        RECT -198.865 -55.435 -198.585 -45.995 ;
        RECT -198.305 -55.155 -198.025 -34.935 ;
        RECT -193.885 -38.295 -193.485 -37.095 ;
        RECT -196.125 -41.655 -195.725 -40.455 ;
        RECT -197.245 -45.015 -196.845 -43.815 ;
        RECT -197.745 -55.435 -197.465 -45.995 ;
        RECT -197.185 -55.155 -196.905 -45.015 ;
        RECT -196.625 -55.435 -196.345 -45.995 ;
        RECT -196.065 -55.155 -195.785 -41.655 ;
        RECT -195.005 -45.015 -194.605 -43.815 ;
        RECT -195.505 -55.435 -195.225 -45.995 ;
        RECT -194.945 -55.155 -194.665 -45.015 ;
        RECT -194.385 -55.435 -194.105 -45.995 ;
        RECT -193.825 -55.155 -193.545 -38.295 ;
        RECT -191.645 -41.655 -191.245 -40.455 ;
        RECT -192.765 -45.015 -192.365 -43.815 ;
        RECT -193.265 -55.435 -192.985 -45.995 ;
        RECT -192.705 -55.155 -192.425 -45.015 ;
        RECT -192.145 -55.435 -191.865 -45.995 ;
        RECT -191.585 -55.155 -191.305 -41.655 ;
        RECT -190.525 -45.015 -190.125 -43.815 ;
        RECT -191.025 -55.435 -190.745 -45.995 ;
        RECT -190.465 -55.155 -190.185 -45.015 ;
        RECT -189.905 -55.435 -189.625 -45.995 ;
        RECT -189.345 -55.155 -189.065 -14.775 ;
        RECT -188.285 -18.135 -187.885 -16.935 ;
        RECT -188.785 -55.435 -188.505 -45.995 ;
        RECT -188.225 -55.155 -187.945 -18.135 ;
        RECT -44.925 -21.495 -44.525 -20.295 ;
        RECT -116.605 -24.855 -116.205 -23.655 ;
        RECT -152.445 -28.215 -152.045 -27.015 ;
        RECT -170.365 -31.575 -169.965 -30.375 ;
        RECT -179.325 -34.935 -178.925 -33.735 ;
        RECT -183.805 -38.295 -183.405 -37.095 ;
        RECT -186.045 -41.655 -185.645 -40.455 ;
        RECT -187.165 -45.015 -186.765 -43.815 ;
        RECT -187.665 -55.435 -187.385 -45.995 ;
        RECT -187.105 -55.155 -186.825 -45.015 ;
        RECT -186.545 -55.435 -186.265 -45.995 ;
        RECT -185.985 -55.155 -185.705 -41.655 ;
        RECT -184.925 -45.015 -184.525 -43.815 ;
        RECT -185.425 -55.435 -185.145 -45.995 ;
        RECT -184.865 -55.155 -184.585 -45.015 ;
        RECT -184.305 -55.435 -184.025 -45.995 ;
        RECT -183.745 -55.155 -183.465 -38.295 ;
        RECT -181.565 -41.655 -181.165 -40.455 ;
        RECT -182.685 -45.015 -182.285 -43.815 ;
        RECT -183.185 -55.435 -182.905 -45.995 ;
        RECT -182.625 -55.155 -182.345 -45.015 ;
        RECT -182.065 -55.435 -181.785 -45.995 ;
        RECT -181.505 -55.155 -181.225 -41.655 ;
        RECT -180.445 -45.015 -180.045 -43.815 ;
        RECT -180.945 -55.435 -180.665 -45.995 ;
        RECT -180.385 -55.155 -180.105 -45.015 ;
        RECT -179.825 -55.435 -179.545 -45.995 ;
        RECT -179.265 -55.155 -178.985 -34.935 ;
        RECT -174.845 -38.295 -174.445 -37.095 ;
        RECT -177.085 -41.655 -176.685 -40.455 ;
        RECT -178.205 -45.015 -177.805 -43.815 ;
        RECT -178.705 -55.435 -178.425 -45.995 ;
        RECT -178.145 -55.155 -177.865 -45.015 ;
        RECT -177.585 -55.435 -177.305 -45.995 ;
        RECT -177.025 -55.155 -176.745 -41.655 ;
        RECT -175.965 -45.015 -175.565 -43.815 ;
        RECT -176.465 -55.435 -176.185 -45.995 ;
        RECT -175.905 -55.155 -175.625 -45.015 ;
        RECT -175.345 -55.435 -175.065 -45.995 ;
        RECT -174.785 -55.155 -174.505 -38.295 ;
        RECT -172.605 -41.655 -172.205 -40.455 ;
        RECT -173.725 -45.015 -173.325 -43.815 ;
        RECT -174.225 -55.435 -173.945 -45.995 ;
        RECT -173.665 -55.155 -173.385 -45.015 ;
        RECT -173.105 -55.435 -172.825 -45.995 ;
        RECT -172.545 -55.155 -172.265 -41.655 ;
        RECT -171.485 -45.015 -171.085 -43.815 ;
        RECT -171.985 -55.435 -171.705 -45.995 ;
        RECT -171.425 -55.155 -171.145 -45.015 ;
        RECT -170.865 -55.435 -170.585 -45.995 ;
        RECT -170.305 -55.155 -170.025 -31.575 ;
        RECT -161.405 -34.935 -161.005 -33.735 ;
        RECT -165.885 -38.295 -165.485 -37.095 ;
        RECT -168.125 -41.655 -167.725 -40.455 ;
        RECT -169.245 -45.015 -168.845 -43.815 ;
        RECT -169.745 -55.435 -169.465 -45.995 ;
        RECT -169.185 -55.155 -168.905 -45.015 ;
        RECT -168.625 -55.435 -168.345 -45.995 ;
        RECT -168.065 -55.155 -167.785 -41.655 ;
        RECT -167.005 -45.015 -166.605 -43.815 ;
        RECT -167.505 -55.435 -167.225 -45.995 ;
        RECT -166.945 -55.155 -166.665 -45.015 ;
        RECT -166.385 -55.435 -166.105 -45.995 ;
        RECT -165.825 -55.155 -165.545 -38.295 ;
        RECT -163.645 -41.655 -163.245 -40.455 ;
        RECT -164.765 -45.015 -164.365 -43.815 ;
        RECT -165.265 -55.435 -164.985 -45.995 ;
        RECT -164.705 -55.155 -164.425 -45.015 ;
        RECT -164.145 -55.435 -163.865 -45.995 ;
        RECT -163.585 -55.155 -163.305 -41.655 ;
        RECT -162.525 -45.015 -162.125 -43.815 ;
        RECT -163.025 -55.435 -162.745 -45.995 ;
        RECT -162.465 -55.155 -162.185 -45.015 ;
        RECT -161.905 -55.435 -161.625 -45.995 ;
        RECT -161.345 -55.155 -161.065 -34.935 ;
        RECT -156.925 -38.295 -156.525 -37.095 ;
        RECT -159.165 -41.655 -158.765 -40.455 ;
        RECT -160.285 -45.015 -159.885 -43.815 ;
        RECT -160.785 -55.435 -160.505 -45.995 ;
        RECT -160.225 -55.155 -159.945 -45.015 ;
        RECT -159.665 -55.435 -159.385 -45.995 ;
        RECT -159.105 -55.155 -158.825 -41.655 ;
        RECT -158.045 -45.015 -157.645 -43.815 ;
        RECT -158.545 -55.435 -158.265 -45.995 ;
        RECT -157.985 -55.155 -157.705 -45.015 ;
        RECT -157.425 -55.435 -157.145 -45.995 ;
        RECT -156.865 -55.155 -156.585 -38.295 ;
        RECT -154.685 -41.655 -154.285 -40.455 ;
        RECT -155.805 -45.015 -155.405 -43.815 ;
        RECT -156.305 -55.435 -156.025 -45.995 ;
        RECT -155.745 -55.155 -155.465 -45.015 ;
        RECT -155.185 -55.435 -154.905 -45.995 ;
        RECT -154.625 -55.155 -154.345 -41.655 ;
        RECT -153.565 -45.015 -153.165 -43.815 ;
        RECT -154.065 -55.435 -153.785 -45.995 ;
        RECT -153.505 -55.155 -153.225 -45.015 ;
        RECT -152.945 -55.435 -152.665 -45.995 ;
        RECT -152.385 -55.155 -152.105 -28.215 ;
        RECT -134.525 -31.575 -134.125 -30.375 ;
        RECT -143.485 -34.935 -143.085 -33.735 ;
        RECT -147.965 -38.295 -147.565 -37.095 ;
        RECT -150.205 -41.655 -149.805 -40.455 ;
        RECT -151.325 -45.015 -150.925 -43.815 ;
        RECT -151.825 -55.435 -151.545 -45.995 ;
        RECT -151.265 -55.155 -150.985 -45.015 ;
        RECT -150.705 -55.435 -150.425 -45.995 ;
        RECT -150.145 -55.155 -149.865 -41.655 ;
        RECT -149.085 -45.015 -148.685 -43.815 ;
        RECT -149.585 -55.435 -149.305 -45.995 ;
        RECT -149.025 -55.155 -148.745 -45.015 ;
        RECT -148.465 -55.435 -148.185 -45.995 ;
        RECT -147.905 -55.155 -147.625 -38.295 ;
        RECT -145.725 -41.655 -145.325 -40.455 ;
        RECT -146.845 -45.015 -146.445 -43.815 ;
        RECT -147.345 -55.435 -147.065 -45.995 ;
        RECT -146.785 -55.155 -146.505 -45.015 ;
        RECT -146.225 -55.435 -145.945 -45.995 ;
        RECT -145.665 -55.155 -145.385 -41.655 ;
        RECT -144.605 -45.015 -144.205 -43.815 ;
        RECT -145.105 -55.435 -144.825 -45.995 ;
        RECT -144.545 -55.155 -144.265 -45.015 ;
        RECT -143.985 -55.435 -143.705 -45.995 ;
        RECT -143.425 -55.155 -143.145 -34.935 ;
        RECT -139.005 -38.295 -138.605 -37.095 ;
        RECT -141.245 -41.655 -140.845 -40.455 ;
        RECT -142.365 -45.015 -141.965 -43.815 ;
        RECT -142.865 -55.435 -142.585 -45.995 ;
        RECT -142.305 -55.155 -142.025 -45.015 ;
        RECT -141.745 -55.435 -141.465 -45.995 ;
        RECT -141.185 -55.155 -140.905 -41.655 ;
        RECT -140.125 -45.015 -139.725 -43.815 ;
        RECT -140.625 -55.435 -140.345 -45.995 ;
        RECT -140.065 -55.155 -139.785 -45.015 ;
        RECT -139.505 -55.435 -139.225 -45.995 ;
        RECT -138.945 -55.155 -138.665 -38.295 ;
        RECT -136.765 -41.655 -136.365 -40.455 ;
        RECT -137.885 -45.015 -137.485 -43.815 ;
        RECT -138.385 -55.435 -138.105 -45.995 ;
        RECT -137.825 -55.155 -137.545 -45.015 ;
        RECT -137.265 -55.435 -136.985 -45.995 ;
        RECT -136.705 -55.155 -136.425 -41.655 ;
        RECT -135.645 -45.015 -135.245 -43.815 ;
        RECT -136.145 -55.435 -135.865 -45.995 ;
        RECT -135.585 -55.155 -135.305 -45.015 ;
        RECT -135.025 -55.435 -134.745 -45.995 ;
        RECT -134.465 -55.155 -134.185 -31.575 ;
        RECT -125.565 -34.935 -125.165 -33.735 ;
        RECT -130.045 -38.295 -129.645 -37.095 ;
        RECT -132.285 -41.655 -131.885 -40.455 ;
        RECT -133.405 -45.015 -133.005 -43.815 ;
        RECT -133.905 -55.435 -133.625 -45.995 ;
        RECT -133.345 -55.155 -133.065 -45.015 ;
        RECT -132.785 -55.435 -132.505 -45.995 ;
        RECT -132.225 -55.155 -131.945 -41.655 ;
        RECT -131.165 -45.015 -130.765 -43.815 ;
        RECT -131.665 -55.435 -131.385 -45.995 ;
        RECT -131.105 -55.155 -130.825 -45.015 ;
        RECT -130.545 -55.435 -130.265 -45.995 ;
        RECT -129.985 -55.155 -129.705 -38.295 ;
        RECT -127.805 -41.655 -127.405 -40.455 ;
        RECT -128.925 -45.015 -128.525 -43.815 ;
        RECT -129.425 -55.435 -129.145 -45.995 ;
        RECT -128.865 -55.155 -128.585 -45.015 ;
        RECT -128.305 -55.435 -128.025 -45.995 ;
        RECT -127.745 -55.155 -127.465 -41.655 ;
        RECT -126.685 -45.015 -126.285 -43.815 ;
        RECT -127.185 -55.435 -126.905 -45.995 ;
        RECT -126.625 -55.155 -126.345 -45.015 ;
        RECT -126.065 -55.435 -125.785 -45.995 ;
        RECT -125.505 -55.155 -125.225 -34.935 ;
        RECT -121.085 -38.295 -120.685 -37.095 ;
        RECT -123.325 -41.655 -122.925 -40.455 ;
        RECT -124.445 -45.015 -124.045 -43.815 ;
        RECT -124.945 -55.435 -124.665 -45.995 ;
        RECT -124.385 -55.155 -124.105 -45.015 ;
        RECT -123.825 -55.435 -123.545 -45.995 ;
        RECT -123.265 -55.155 -122.985 -41.655 ;
        RECT -122.205 -45.015 -121.805 -43.815 ;
        RECT -122.705 -55.435 -122.425 -45.995 ;
        RECT -122.145 -55.155 -121.865 -45.015 ;
        RECT -121.585 -55.435 -121.305 -45.995 ;
        RECT -121.025 -55.155 -120.745 -38.295 ;
        RECT -118.845 -41.655 -118.445 -40.455 ;
        RECT -119.965 -45.015 -119.565 -43.815 ;
        RECT -120.465 -55.435 -120.185 -45.995 ;
        RECT -119.905 -55.155 -119.625 -45.015 ;
        RECT -119.345 -55.435 -119.065 -45.995 ;
        RECT -118.785 -55.155 -118.505 -41.655 ;
        RECT -117.725 -45.015 -117.325 -43.815 ;
        RECT -118.225 -55.435 -117.945 -45.995 ;
        RECT -117.665 -55.155 -117.385 -45.015 ;
        RECT -117.105 -55.435 -116.825 -45.995 ;
        RECT -116.545 -55.155 -116.265 -24.855 ;
        RECT -80.765 -28.215 -80.365 -27.015 ;
        RECT -98.685 -31.575 -98.285 -30.375 ;
        RECT -107.645 -34.935 -107.245 -33.735 ;
        RECT -112.125 -38.295 -111.725 -37.095 ;
        RECT -114.365 -41.655 -113.965 -40.455 ;
        RECT -115.485 -45.015 -115.085 -43.815 ;
        RECT -115.985 -55.435 -115.705 -45.995 ;
        RECT -115.425 -55.155 -115.145 -45.015 ;
        RECT -114.865 -55.435 -114.585 -45.995 ;
        RECT -114.305 -55.155 -114.025 -41.655 ;
        RECT -113.245 -45.015 -112.845 -43.815 ;
        RECT -113.745 -55.435 -113.465 -45.995 ;
        RECT -113.185 -55.155 -112.905 -45.015 ;
        RECT -112.625 -55.435 -112.345 -45.995 ;
        RECT -112.065 -55.155 -111.785 -38.295 ;
        RECT -109.885 -41.655 -109.485 -40.455 ;
        RECT -111.005 -45.015 -110.605 -43.815 ;
        RECT -111.505 -55.435 -111.225 -45.995 ;
        RECT -110.945 -55.155 -110.665 -45.015 ;
        RECT -110.385 -55.435 -110.105 -45.995 ;
        RECT -109.825 -55.155 -109.545 -41.655 ;
        RECT -108.765 -45.015 -108.365 -43.815 ;
        RECT -109.265 -55.435 -108.985 -45.995 ;
        RECT -108.705 -55.155 -108.425 -45.015 ;
        RECT -108.145 -55.435 -107.865 -45.995 ;
        RECT -107.585 -55.155 -107.305 -34.935 ;
        RECT -103.165 -38.295 -102.765 -37.095 ;
        RECT -105.405 -41.655 -105.005 -40.455 ;
        RECT -106.525 -45.015 -106.125 -43.815 ;
        RECT -107.025 -55.435 -106.745 -45.995 ;
        RECT -106.465 -55.155 -106.185 -45.015 ;
        RECT -105.905 -55.435 -105.625 -45.995 ;
        RECT -105.345 -55.155 -105.065 -41.655 ;
        RECT -104.285 -45.015 -103.885 -43.815 ;
        RECT -104.785 -55.435 -104.505 -45.995 ;
        RECT -104.225 -55.155 -103.945 -45.015 ;
        RECT -103.665 -55.435 -103.385 -45.995 ;
        RECT -103.105 -55.155 -102.825 -38.295 ;
        RECT -100.925 -41.655 -100.525 -40.455 ;
        RECT -102.045 -45.015 -101.645 -43.815 ;
        RECT -102.545 -55.435 -102.265 -45.995 ;
        RECT -101.985 -55.155 -101.705 -45.015 ;
        RECT -101.425 -55.435 -101.145 -45.995 ;
        RECT -100.865 -55.155 -100.585 -41.655 ;
        RECT -99.805 -45.015 -99.405 -43.815 ;
        RECT -100.305 -55.435 -100.025 -45.995 ;
        RECT -99.745 -55.155 -99.465 -45.015 ;
        RECT -99.185 -55.435 -98.905 -45.995 ;
        RECT -98.625 -55.155 -98.345 -31.575 ;
        RECT -89.725 -34.935 -89.325 -33.735 ;
        RECT -94.205 -38.295 -93.805 -37.095 ;
        RECT -96.445 -41.655 -96.045 -40.455 ;
        RECT -97.565 -45.015 -97.165 -43.815 ;
        RECT -98.065 -55.435 -97.785 -45.995 ;
        RECT -97.505 -55.155 -97.225 -45.015 ;
        RECT -96.945 -55.435 -96.665 -45.995 ;
        RECT -96.385 -55.155 -96.105 -41.655 ;
        RECT -95.325 -45.015 -94.925 -43.815 ;
        RECT -95.825 -55.435 -95.545 -45.995 ;
        RECT -95.265 -55.155 -94.985 -45.015 ;
        RECT -94.705 -55.435 -94.425 -45.995 ;
        RECT -94.145 -55.155 -93.865 -38.295 ;
        RECT -91.965 -41.655 -91.565 -40.455 ;
        RECT -93.085 -45.015 -92.685 -43.815 ;
        RECT -93.585 -55.435 -93.305 -45.995 ;
        RECT -93.025 -55.155 -92.745 -45.015 ;
        RECT -92.465 -55.435 -92.185 -45.995 ;
        RECT -91.905 -55.155 -91.625 -41.655 ;
        RECT -90.845 -45.015 -90.445 -43.815 ;
        RECT -91.345 -55.435 -91.065 -45.995 ;
        RECT -90.785 -55.155 -90.505 -45.015 ;
        RECT -90.225 -55.435 -89.945 -45.995 ;
        RECT -89.665 -55.155 -89.385 -34.935 ;
        RECT -85.245 -38.295 -84.845 -37.095 ;
        RECT -87.485 -41.655 -87.085 -40.455 ;
        RECT -88.605 -45.015 -88.205 -43.815 ;
        RECT -89.105 -55.435 -88.825 -45.995 ;
        RECT -88.545 -55.155 -88.265 -45.015 ;
        RECT -87.985 -55.435 -87.705 -45.995 ;
        RECT -87.425 -55.155 -87.145 -41.655 ;
        RECT -86.365 -45.015 -85.965 -43.815 ;
        RECT -86.865 -55.435 -86.585 -45.995 ;
        RECT -86.305 -55.155 -86.025 -45.015 ;
        RECT -85.745 -55.435 -85.465 -45.995 ;
        RECT -85.185 -55.155 -84.905 -38.295 ;
        RECT -83.005 -41.655 -82.605 -40.455 ;
        RECT -84.125 -45.015 -83.725 -43.815 ;
        RECT -84.625 -55.435 -84.345 -45.995 ;
        RECT -84.065 -55.155 -83.785 -45.015 ;
        RECT -83.505 -55.435 -83.225 -45.995 ;
        RECT -82.945 -55.155 -82.665 -41.655 ;
        RECT -81.885 -45.015 -81.485 -43.815 ;
        RECT -82.385 -55.435 -82.105 -45.995 ;
        RECT -81.825 -55.155 -81.545 -45.015 ;
        RECT -81.265 -55.435 -80.985 -45.995 ;
        RECT -80.705 -55.155 -80.425 -28.215 ;
        RECT -62.845 -31.575 -62.445 -30.375 ;
        RECT -71.805 -34.935 -71.405 -33.735 ;
        RECT -76.285 -38.295 -75.885 -37.095 ;
        RECT -78.525 -41.655 -78.125 -40.455 ;
        RECT -79.645 -45.015 -79.245 -43.815 ;
        RECT -80.145 -55.435 -79.865 -45.995 ;
        RECT -79.585 -55.155 -79.305 -45.015 ;
        RECT -79.025 -55.435 -78.745 -45.995 ;
        RECT -78.465 -55.155 -78.185 -41.655 ;
        RECT -77.405 -45.015 -77.005 -43.815 ;
        RECT -77.905 -55.435 -77.625 -45.995 ;
        RECT -77.345 -55.155 -77.065 -45.015 ;
        RECT -76.785 -55.435 -76.505 -45.995 ;
        RECT -76.225 -55.155 -75.945 -38.295 ;
        RECT -74.045 -41.655 -73.645 -40.455 ;
        RECT -75.165 -45.015 -74.765 -43.815 ;
        RECT -75.665 -55.435 -75.385 -45.995 ;
        RECT -75.105 -55.155 -74.825 -45.015 ;
        RECT -74.545 -55.435 -74.265 -45.995 ;
        RECT -73.985 -55.155 -73.705 -41.655 ;
        RECT -72.925 -45.015 -72.525 -43.815 ;
        RECT -73.425 -55.435 -73.145 -45.995 ;
        RECT -72.865 -55.155 -72.585 -45.015 ;
        RECT -72.305 -55.435 -72.025 -45.995 ;
        RECT -71.745 -55.155 -71.465 -34.935 ;
        RECT -67.325 -38.295 -66.925 -37.095 ;
        RECT -69.565 -41.655 -69.165 -40.455 ;
        RECT -70.685 -45.015 -70.285 -43.815 ;
        RECT -71.185 -55.435 -70.905 -45.995 ;
        RECT -70.625 -55.155 -70.345 -45.015 ;
        RECT -70.065 -55.435 -69.785 -45.995 ;
        RECT -69.505 -55.155 -69.225 -41.655 ;
        RECT -68.445 -45.015 -68.045 -43.815 ;
        RECT -68.945 -55.435 -68.665 -45.995 ;
        RECT -68.385 -55.155 -68.105 -45.015 ;
        RECT -67.825 -55.435 -67.545 -45.995 ;
        RECT -67.265 -55.155 -66.985 -38.295 ;
        RECT -65.085 -41.655 -64.685 -40.455 ;
        RECT -66.205 -45.015 -65.805 -43.815 ;
        RECT -66.705 -55.435 -66.425 -45.995 ;
        RECT -66.145 -55.155 -65.865 -45.015 ;
        RECT -65.585 -55.435 -65.305 -45.995 ;
        RECT -65.025 -55.155 -64.745 -41.655 ;
        RECT -63.965 -45.015 -63.565 -43.815 ;
        RECT -64.465 -55.435 -64.185 -45.995 ;
        RECT -63.905 -55.155 -63.625 -45.015 ;
        RECT -63.345 -55.435 -63.065 -45.995 ;
        RECT -62.785 -55.155 -62.505 -31.575 ;
        RECT -53.885 -34.935 -53.485 -33.735 ;
        RECT -58.365 -38.295 -57.965 -37.095 ;
        RECT -60.605 -41.655 -60.205 -40.455 ;
        RECT -61.725 -45.015 -61.325 -43.815 ;
        RECT -62.225 -55.435 -61.945 -45.995 ;
        RECT -61.665 -55.155 -61.385 -45.015 ;
        RECT -61.105 -55.435 -60.825 -45.995 ;
        RECT -60.545 -55.155 -60.265 -41.655 ;
        RECT -59.485 -45.015 -59.085 -43.815 ;
        RECT -59.985 -55.435 -59.705 -45.995 ;
        RECT -59.425 -55.155 -59.145 -45.015 ;
        RECT -58.865 -55.435 -58.585 -45.995 ;
        RECT -58.305 -55.155 -58.025 -38.295 ;
        RECT -56.125 -41.655 -55.725 -40.455 ;
        RECT -57.245 -45.015 -56.845 -43.815 ;
        RECT -57.745 -55.435 -57.465 -45.995 ;
        RECT -57.185 -55.155 -56.905 -45.015 ;
        RECT -56.625 -55.435 -56.345 -45.995 ;
        RECT -56.065 -55.155 -55.785 -41.655 ;
        RECT -55.005 -45.015 -54.605 -43.815 ;
        RECT -55.505 -55.435 -55.225 -45.995 ;
        RECT -54.945 -55.155 -54.665 -45.015 ;
        RECT -54.385 -55.435 -54.105 -45.995 ;
        RECT -53.825 -55.155 -53.545 -34.935 ;
        RECT -49.405 -38.295 -49.005 -37.095 ;
        RECT -51.645 -41.655 -51.245 -40.455 ;
        RECT -52.765 -45.015 -52.365 -43.815 ;
        RECT -53.265 -55.435 -52.985 -45.995 ;
        RECT -52.705 -55.155 -52.425 -45.015 ;
        RECT -52.145 -55.435 -51.865 -45.995 ;
        RECT -51.585 -55.155 -51.305 -41.655 ;
        RECT -50.525 -45.015 -50.125 -43.815 ;
        RECT -51.025 -55.435 -50.745 -45.995 ;
        RECT -50.465 -55.155 -50.185 -45.015 ;
        RECT -49.905 -55.435 -49.625 -45.995 ;
        RECT -49.345 -55.155 -49.065 -38.295 ;
        RECT -47.165 -41.655 -46.765 -40.455 ;
        RECT -48.285 -45.015 -47.885 -43.815 ;
        RECT -48.785 -55.435 -48.505 -45.995 ;
        RECT -48.225 -55.155 -47.945 -45.015 ;
        RECT -47.665 -55.435 -47.385 -45.995 ;
        RECT -47.105 -55.155 -46.825 -41.655 ;
        RECT -46.045 -45.015 -45.645 -43.815 ;
        RECT -46.545 -55.435 -46.265 -45.995 ;
        RECT -45.985 -55.155 -45.705 -45.015 ;
        RECT -45.425 -55.435 -45.145 -45.995 ;
        RECT -44.865 -55.155 -44.585 -21.495 ;
        RECT 26.755 -24.855 27.155 -23.655 ;
        RECT -9.085 -28.215 -8.685 -27.015 ;
        RECT -27.005 -31.575 -26.605 -30.375 ;
        RECT -35.965 -34.935 -35.565 -33.735 ;
        RECT -40.445 -38.295 -40.045 -37.095 ;
        RECT -42.685 -41.655 -42.285 -40.455 ;
        RECT -43.805 -45.015 -43.405 -43.815 ;
        RECT -44.305 -55.435 -44.025 -45.995 ;
        RECT -43.745 -55.155 -43.465 -45.015 ;
        RECT -43.185 -55.435 -42.905 -45.995 ;
        RECT -42.625 -55.155 -42.345 -41.655 ;
        RECT -41.565 -45.015 -41.165 -43.815 ;
        RECT -42.065 -55.435 -41.785 -45.995 ;
        RECT -41.505 -55.155 -41.225 -45.015 ;
        RECT -40.945 -55.435 -40.665 -45.995 ;
        RECT -40.385 -55.155 -40.105 -38.295 ;
        RECT -38.205 -41.655 -37.805 -40.455 ;
        RECT -39.325 -45.015 -38.925 -43.815 ;
        RECT -39.825 -55.435 -39.545 -45.995 ;
        RECT -39.265 -55.155 -38.985 -45.015 ;
        RECT -38.705 -55.435 -38.425 -45.995 ;
        RECT -38.145 -55.155 -37.865 -41.655 ;
        RECT -37.085 -45.015 -36.685 -43.815 ;
        RECT -37.585 -55.435 -37.305 -45.995 ;
        RECT -37.025 -55.155 -36.745 -45.015 ;
        RECT -36.465 -55.435 -36.185 -45.995 ;
        RECT -35.905 -55.155 -35.625 -34.935 ;
        RECT -31.485 -38.295 -31.085 -37.095 ;
        RECT -33.725 -41.655 -33.325 -40.455 ;
        RECT -34.845 -45.015 -34.445 -43.815 ;
        RECT -35.345 -55.435 -35.065 -45.995 ;
        RECT -34.785 -55.155 -34.505 -45.015 ;
        RECT -34.225 -55.435 -33.945 -45.995 ;
        RECT -33.665 -55.155 -33.385 -41.655 ;
        RECT -32.605 -45.015 -32.205 -43.815 ;
        RECT -33.105 -55.435 -32.825 -45.995 ;
        RECT -32.545 -55.155 -32.265 -45.015 ;
        RECT -31.985 -55.435 -31.705 -45.995 ;
        RECT -31.425 -55.155 -31.145 -38.295 ;
        RECT -29.245 -41.655 -28.845 -40.455 ;
        RECT -30.365 -45.015 -29.965 -43.815 ;
        RECT -30.865 -55.435 -30.585 -45.995 ;
        RECT -30.305 -55.155 -30.025 -45.015 ;
        RECT -29.745 -55.435 -29.465 -45.995 ;
        RECT -29.185 -55.155 -28.905 -41.655 ;
        RECT -28.125 -45.015 -27.725 -43.815 ;
        RECT -28.625 -55.435 -28.345 -45.995 ;
        RECT -28.065 -55.155 -27.785 -45.015 ;
        RECT -27.505 -55.435 -27.225 -45.995 ;
        RECT -26.945 -55.155 -26.665 -31.575 ;
        RECT -18.045 -34.935 -17.645 -33.735 ;
        RECT -22.525 -38.295 -22.125 -37.095 ;
        RECT -24.765 -41.655 -24.365 -40.455 ;
        RECT -25.885 -45.015 -25.485 -43.815 ;
        RECT -26.385 -55.435 -26.105 -45.995 ;
        RECT -25.825 -55.155 -25.545 -45.015 ;
        RECT -25.265 -55.435 -24.985 -45.995 ;
        RECT -24.705 -55.155 -24.425 -41.655 ;
        RECT -23.645 -45.015 -23.245 -43.815 ;
        RECT -24.145 -55.435 -23.865 -45.995 ;
        RECT -23.585 -55.155 -23.305 -45.015 ;
        RECT -23.025 -55.435 -22.745 -45.995 ;
        RECT -22.465 -55.155 -22.185 -38.295 ;
        RECT -20.285 -41.655 -19.885 -40.455 ;
        RECT -21.405 -45.015 -21.005 -43.815 ;
        RECT -21.905 -55.435 -21.625 -45.995 ;
        RECT -21.345 -55.155 -21.065 -45.015 ;
        RECT -20.785 -55.435 -20.505 -45.995 ;
        RECT -20.225 -55.155 -19.945 -41.655 ;
        RECT -19.165 -45.015 -18.765 -43.815 ;
        RECT -19.665 -55.435 -19.385 -45.995 ;
        RECT -19.105 -55.155 -18.825 -45.015 ;
        RECT -18.545 -55.435 -18.265 -45.995 ;
        RECT -17.985 -55.155 -17.705 -34.935 ;
        RECT -13.565 -38.295 -13.165 -37.095 ;
        RECT -15.805 -41.655 -15.405 -40.455 ;
        RECT -16.925 -45.015 -16.525 -43.815 ;
        RECT -17.425 -55.435 -17.145 -45.995 ;
        RECT -16.865 -55.155 -16.585 -45.015 ;
        RECT -16.305 -55.435 -16.025 -45.995 ;
        RECT -15.745 -55.155 -15.465 -41.655 ;
        RECT -14.685 -45.015 -14.285 -43.815 ;
        RECT -15.185 -55.435 -14.905 -45.995 ;
        RECT -14.625 -55.155 -14.345 -45.015 ;
        RECT -14.065 -55.435 -13.785 -45.995 ;
        RECT -13.505 -55.155 -13.225 -38.295 ;
        RECT -11.325 -41.655 -10.925 -40.455 ;
        RECT -12.445 -45.015 -12.045 -43.815 ;
        RECT -12.945 -55.435 -12.665 -45.995 ;
        RECT -12.385 -55.155 -12.105 -45.015 ;
        RECT -11.825 -55.435 -11.545 -45.995 ;
        RECT -11.265 -55.155 -10.985 -41.655 ;
        RECT -10.205 -45.015 -9.805 -43.815 ;
        RECT -10.705 -55.435 -10.425 -45.995 ;
        RECT -10.145 -55.155 -9.865 -45.015 ;
        RECT -9.585 -55.435 -9.305 -45.995 ;
        RECT -9.025 -55.155 -8.745 -28.215 ;
        RECT 8.835 -31.575 9.235 -30.375 ;
        RECT -0.125 -34.935 0.275 -33.735 ;
        RECT -4.605 -38.295 -4.205 -37.095 ;
        RECT -6.845 -41.655 -6.445 -40.455 ;
        RECT -7.965 -45.015 -7.565 -43.815 ;
        RECT -8.465 -55.435 -8.185 -45.995 ;
        RECT -7.905 -55.155 -7.625 -45.015 ;
        RECT -7.345 -55.435 -7.065 -45.995 ;
        RECT -6.785 -55.155 -6.505 -41.655 ;
        RECT -5.725 -45.015 -5.325 -43.815 ;
        RECT -6.225 -55.435 -5.945 -45.995 ;
        RECT -5.665 -55.155 -5.385 -45.015 ;
        RECT -5.105 -55.435 -4.825 -45.995 ;
        RECT -4.545 -55.155 -4.265 -38.295 ;
        RECT -2.365 -41.655 -1.965 -40.455 ;
        RECT -3.485 -45.015 -3.085 -43.815 ;
        RECT -3.985 -55.435 -3.705 -45.995 ;
        RECT -3.425 -55.155 -3.145 -45.015 ;
        RECT -2.865 -55.435 -2.585 -45.995 ;
        RECT -2.305 -55.155 -2.025 -41.655 ;
        RECT -1.245 -45.015 -0.845 -43.815 ;
        RECT -1.745 -55.435 -1.465 -45.995 ;
        RECT -1.185 -55.155 -0.905 -45.015 ;
        RECT -0.625 -55.435 -0.345 -45.995 ;
        RECT -0.065 -55.155 0.215 -34.935 ;
        RECT 4.355 -38.295 4.755 -37.095 ;
        RECT 2.115 -41.655 2.515 -40.455 ;
        RECT 0.995 -45.015 1.395 -43.815 ;
        RECT 0.495 -55.435 0.775 -45.995 ;
        RECT 1.055 -55.155 1.335 -45.015 ;
        RECT 1.615 -55.435 1.895 -45.995 ;
        RECT 2.175 -55.155 2.455 -41.655 ;
        RECT 3.235 -45.015 3.635 -43.815 ;
        RECT 2.735 -55.435 3.015 -45.995 ;
        RECT 3.295 -55.155 3.575 -45.015 ;
        RECT 3.855 -55.435 4.135 -45.995 ;
        RECT 4.415 -55.155 4.695 -38.295 ;
        RECT 6.595 -41.655 6.995 -40.455 ;
        RECT 5.475 -45.015 5.875 -43.815 ;
        RECT 4.975 -55.435 5.255 -45.995 ;
        RECT 5.535 -55.155 5.815 -45.015 ;
        RECT 6.095 -55.435 6.375 -45.995 ;
        RECT 6.655 -55.155 6.935 -41.655 ;
        RECT 7.715 -45.015 8.115 -43.815 ;
        RECT 7.215 -55.435 7.495 -45.995 ;
        RECT 7.775 -55.155 8.055 -45.015 ;
        RECT 8.335 -55.435 8.615 -45.995 ;
        RECT 8.895 -55.155 9.175 -31.575 ;
        RECT 17.795 -34.935 18.195 -33.735 ;
        RECT 13.315 -38.295 13.715 -37.095 ;
        RECT 11.075 -41.655 11.475 -40.455 ;
        RECT 9.955 -45.015 10.355 -43.815 ;
        RECT 9.455 -55.435 9.735 -45.995 ;
        RECT 10.015 -55.155 10.295 -45.015 ;
        RECT 10.575 -55.435 10.855 -45.995 ;
        RECT 11.135 -55.155 11.415 -41.655 ;
        RECT 12.195 -45.015 12.595 -43.815 ;
        RECT 11.695 -55.435 11.975 -45.995 ;
        RECT 12.255 -55.155 12.535 -45.015 ;
        RECT 12.815 -55.435 13.095 -45.995 ;
        RECT 13.375 -55.155 13.655 -38.295 ;
        RECT 15.555 -41.655 15.955 -40.455 ;
        RECT 14.435 -45.015 14.835 -43.815 ;
        RECT 13.935 -55.435 14.215 -45.995 ;
        RECT 14.495 -55.155 14.775 -45.015 ;
        RECT 15.055 -55.435 15.335 -45.995 ;
        RECT 15.615 -55.155 15.895 -41.655 ;
        RECT 16.675 -45.015 17.075 -43.815 ;
        RECT 16.175 -55.435 16.455 -45.995 ;
        RECT 16.735 -55.155 17.015 -45.015 ;
        RECT 17.295 -55.435 17.575 -45.995 ;
        RECT 17.855 -55.155 18.135 -34.935 ;
        RECT 22.275 -38.295 22.675 -37.095 ;
        RECT 20.035 -41.655 20.435 -40.455 ;
        RECT 18.915 -45.015 19.315 -43.815 ;
        RECT 18.415 -55.435 18.695 -45.995 ;
        RECT 18.975 -55.155 19.255 -45.015 ;
        RECT 19.535 -55.435 19.815 -45.995 ;
        RECT 20.095 -55.155 20.375 -41.655 ;
        RECT 21.155 -45.015 21.555 -43.815 ;
        RECT 20.655 -55.435 20.935 -45.995 ;
        RECT 21.215 -55.155 21.495 -45.015 ;
        RECT 21.775 -55.435 22.055 -45.995 ;
        RECT 22.335 -55.155 22.615 -38.295 ;
        RECT 24.515 -41.655 24.915 -40.455 ;
        RECT 23.395 -45.015 23.795 -43.815 ;
        RECT 22.895 -55.435 23.175 -45.995 ;
        RECT 23.455 -55.155 23.735 -45.015 ;
        RECT 24.015 -55.435 24.295 -45.995 ;
        RECT 24.575 -55.155 24.855 -41.655 ;
        RECT 25.635 -45.015 26.035 -43.815 ;
        RECT 25.135 -55.435 25.415 -45.995 ;
        RECT 25.695 -55.155 25.975 -45.015 ;
        RECT 26.255 -55.435 26.535 -45.995 ;
        RECT 26.815 -55.155 27.095 -24.855 ;
        RECT 62.595 -28.215 62.995 -27.015 ;
        RECT 44.675 -31.575 45.075 -30.375 ;
        RECT 35.715 -34.935 36.115 -33.735 ;
        RECT 31.235 -38.295 31.635 -37.095 ;
        RECT 28.995 -41.655 29.395 -40.455 ;
        RECT 27.875 -45.015 28.275 -43.815 ;
        RECT 27.375 -55.435 27.655 -45.995 ;
        RECT 27.935 -55.155 28.215 -45.015 ;
        RECT 28.495 -55.435 28.775 -45.995 ;
        RECT 29.055 -55.155 29.335 -41.655 ;
        RECT 30.115 -45.015 30.515 -43.815 ;
        RECT 29.615 -55.435 29.895 -45.995 ;
        RECT 30.175 -55.155 30.455 -45.015 ;
        RECT 30.735 -55.435 31.015 -45.995 ;
        RECT 31.295 -55.155 31.575 -38.295 ;
        RECT 33.475 -41.655 33.875 -40.455 ;
        RECT 32.355 -45.015 32.755 -43.815 ;
        RECT 31.855 -55.435 32.135 -45.995 ;
        RECT 32.415 -55.155 32.695 -45.015 ;
        RECT 32.975 -55.435 33.255 -45.995 ;
        RECT 33.535 -55.155 33.815 -41.655 ;
        RECT 34.595 -45.015 34.995 -43.815 ;
        RECT 34.095 -55.435 34.375 -45.995 ;
        RECT 34.655 -55.155 34.935 -45.015 ;
        RECT 35.215 -55.435 35.495 -45.995 ;
        RECT 35.775 -55.155 36.055 -34.935 ;
        RECT 40.195 -38.295 40.595 -37.095 ;
        RECT 37.955 -41.655 38.355 -40.455 ;
        RECT 36.835 -45.015 37.235 -43.815 ;
        RECT 36.335 -55.435 36.615 -45.995 ;
        RECT 36.895 -55.155 37.175 -45.015 ;
        RECT 37.455 -55.435 37.735 -45.995 ;
        RECT 38.015 -55.155 38.295 -41.655 ;
        RECT 39.075 -45.015 39.475 -43.815 ;
        RECT 38.575 -55.435 38.855 -45.995 ;
        RECT 39.135 -55.155 39.415 -45.015 ;
        RECT 39.695 -55.435 39.975 -45.995 ;
        RECT 40.255 -55.155 40.535 -38.295 ;
        RECT 42.435 -41.655 42.835 -40.455 ;
        RECT 41.315 -45.015 41.715 -43.815 ;
        RECT 40.815 -55.435 41.095 -45.995 ;
        RECT 41.375 -55.155 41.655 -45.015 ;
        RECT 41.935 -55.435 42.215 -45.995 ;
        RECT 42.495 -55.155 42.775 -41.655 ;
        RECT 43.555 -45.015 43.955 -43.815 ;
        RECT 43.055 -55.435 43.335 -45.995 ;
        RECT 43.615 -55.155 43.895 -45.015 ;
        RECT 44.175 -55.435 44.455 -45.995 ;
        RECT 44.735 -55.155 45.015 -31.575 ;
        RECT 53.635 -34.935 54.035 -33.735 ;
        RECT 49.155 -38.295 49.555 -37.095 ;
        RECT 46.915 -41.655 47.315 -40.455 ;
        RECT 45.795 -45.015 46.195 -43.815 ;
        RECT 45.295 -55.435 45.575 -45.995 ;
        RECT 45.855 -55.155 46.135 -45.015 ;
        RECT 46.415 -55.435 46.695 -45.995 ;
        RECT 46.975 -55.155 47.255 -41.655 ;
        RECT 48.035 -45.015 48.435 -43.815 ;
        RECT 47.535 -55.435 47.815 -45.995 ;
        RECT 48.095 -55.155 48.375 -45.015 ;
        RECT 48.655 -55.435 48.935 -45.995 ;
        RECT 49.215 -55.155 49.495 -38.295 ;
        RECT 51.395 -41.655 51.795 -40.455 ;
        RECT 50.275 -45.015 50.675 -43.815 ;
        RECT 49.775 -55.435 50.055 -45.995 ;
        RECT 50.335 -55.155 50.615 -45.015 ;
        RECT 50.895 -55.435 51.175 -45.995 ;
        RECT 51.455 -55.155 51.735 -41.655 ;
        RECT 52.515 -45.015 52.915 -43.815 ;
        RECT 52.015 -55.435 52.295 -45.995 ;
        RECT 52.575 -55.155 52.855 -45.015 ;
        RECT 53.135 -55.435 53.415 -45.995 ;
        RECT 53.695 -55.155 53.975 -34.935 ;
        RECT 58.115 -38.295 58.515 -37.095 ;
        RECT 55.875 -41.655 56.275 -40.455 ;
        RECT 54.755 -45.015 55.155 -43.815 ;
        RECT 54.255 -55.435 54.535 -45.995 ;
        RECT 54.815 -55.155 55.095 -45.015 ;
        RECT 55.375 -55.435 55.655 -45.995 ;
        RECT 55.935 -55.155 56.215 -41.655 ;
        RECT 56.995 -45.015 57.395 -43.815 ;
        RECT 56.495 -55.435 56.775 -45.995 ;
        RECT 57.055 -55.155 57.335 -45.015 ;
        RECT 57.615 -55.435 57.895 -45.995 ;
        RECT 58.175 -55.155 58.455 -38.295 ;
        RECT 60.355 -41.655 60.755 -40.455 ;
        RECT 59.235 -45.015 59.635 -43.815 ;
        RECT 58.735 -55.435 59.015 -45.995 ;
        RECT 59.295 -55.155 59.575 -45.015 ;
        RECT 59.855 -55.435 60.135 -45.995 ;
        RECT 60.415 -55.155 60.695 -41.655 ;
        RECT 61.475 -45.015 61.875 -43.815 ;
        RECT 60.975 -55.435 61.255 -45.995 ;
        RECT 61.535 -55.155 61.815 -45.015 ;
        RECT 62.095 -55.435 62.375 -45.995 ;
        RECT 62.655 -55.155 62.935 -28.215 ;
        RECT 80.515 -31.575 80.915 -30.375 ;
        RECT 71.555 -34.935 71.955 -33.735 ;
        RECT 67.075 -38.295 67.475 -37.095 ;
        RECT 64.835 -41.655 65.235 -40.455 ;
        RECT 63.715 -45.015 64.115 -43.815 ;
        RECT 63.215 -55.435 63.495 -45.995 ;
        RECT 63.775 -55.155 64.055 -45.015 ;
        RECT 64.335 -55.435 64.615 -45.995 ;
        RECT 64.895 -55.155 65.175 -41.655 ;
        RECT 65.955 -45.015 66.355 -43.815 ;
        RECT 65.455 -55.435 65.735 -45.995 ;
        RECT 66.015 -55.155 66.295 -45.015 ;
        RECT 66.575 -55.435 66.855 -45.995 ;
        RECT 67.135 -55.155 67.415 -38.295 ;
        RECT 69.315 -41.655 69.715 -40.455 ;
        RECT 68.195 -45.015 68.595 -43.815 ;
        RECT 67.695 -55.435 67.975 -45.995 ;
        RECT 68.255 -55.155 68.535 -45.015 ;
        RECT 68.815 -55.435 69.095 -45.995 ;
        RECT 69.375 -55.155 69.655 -41.655 ;
        RECT 70.435 -45.015 70.835 -43.815 ;
        RECT 69.935 -55.435 70.215 -45.995 ;
        RECT 70.495 -55.155 70.775 -45.015 ;
        RECT 71.055 -55.435 71.335 -45.995 ;
        RECT 71.615 -55.155 71.895 -34.935 ;
        RECT 76.035 -38.295 76.435 -37.095 ;
        RECT 73.795 -41.655 74.195 -40.455 ;
        RECT 72.675 -45.015 73.075 -43.815 ;
        RECT 72.175 -55.435 72.455 -45.995 ;
        RECT 72.735 -55.155 73.015 -45.015 ;
        RECT 73.295 -55.435 73.575 -45.995 ;
        RECT 73.855 -55.155 74.135 -41.655 ;
        RECT 74.915 -45.015 75.315 -43.815 ;
        RECT 74.415 -55.435 74.695 -45.995 ;
        RECT 74.975 -55.155 75.255 -45.015 ;
        RECT 75.535 -55.435 75.815 -45.995 ;
        RECT 76.095 -55.155 76.375 -38.295 ;
        RECT 78.275 -41.655 78.675 -40.455 ;
        RECT 77.155 -45.015 77.555 -43.815 ;
        RECT 76.655 -55.435 76.935 -45.995 ;
        RECT 77.215 -55.155 77.495 -45.015 ;
        RECT 77.775 -55.435 78.055 -45.995 ;
        RECT 78.335 -55.155 78.615 -41.655 ;
        RECT 79.395 -45.015 79.795 -43.815 ;
        RECT 78.895 -55.435 79.175 -45.995 ;
        RECT 79.455 -55.155 79.735 -45.015 ;
        RECT 80.015 -55.435 80.295 -45.995 ;
        RECT 80.575 -55.155 80.855 -31.575 ;
        RECT 89.475 -34.935 89.875 -33.735 ;
        RECT 84.995 -38.295 85.395 -37.095 ;
        RECT 82.755 -41.655 83.155 -40.455 ;
        RECT 81.635 -45.015 82.035 -43.815 ;
        RECT 81.135 -55.435 81.415 -45.995 ;
        RECT 81.695 -55.155 81.975 -45.015 ;
        RECT 82.255 -55.435 82.535 -45.995 ;
        RECT 82.815 -55.155 83.095 -41.655 ;
        RECT 83.875 -45.015 84.275 -43.815 ;
        RECT 83.375 -55.435 83.655 -45.995 ;
        RECT 83.935 -55.155 84.215 -45.015 ;
        RECT 84.495 -55.435 84.775 -45.995 ;
        RECT 85.055 -55.155 85.335 -38.295 ;
        RECT 87.235 -41.655 87.635 -40.455 ;
        RECT 86.115 -45.015 86.515 -43.815 ;
        RECT 85.615 -55.435 85.895 -45.995 ;
        RECT 86.175 -55.155 86.455 -45.015 ;
        RECT 86.735 -55.435 87.015 -45.995 ;
        RECT 87.295 -55.155 87.575 -41.655 ;
        RECT 88.355 -45.015 88.755 -43.815 ;
        RECT 87.855 -55.435 88.135 -45.995 ;
        RECT 88.415 -55.155 88.695 -45.015 ;
        RECT 88.975 -55.435 89.255 -45.995 ;
        RECT 89.535 -55.155 89.815 -34.935 ;
        RECT 93.955 -38.295 94.355 -37.095 ;
        RECT 91.715 -41.655 92.115 -40.455 ;
        RECT 90.595 -45.015 90.995 -43.815 ;
        RECT 90.095 -55.435 90.375 -45.995 ;
        RECT 90.655 -55.155 90.935 -45.015 ;
        RECT 91.215 -55.435 91.495 -45.995 ;
        RECT 91.775 -55.155 92.055 -41.655 ;
        RECT 92.835 -45.015 93.235 -43.815 ;
        RECT 92.335 -55.435 92.615 -45.995 ;
        RECT 92.895 -55.155 93.175 -45.015 ;
        RECT 93.455 -55.435 93.735 -45.995 ;
        RECT 94.015 -55.155 94.295 -38.295 ;
        RECT 96.195 -41.655 96.595 -40.455 ;
        RECT 95.075 -45.015 95.475 -43.815 ;
        RECT 94.575 -55.435 94.855 -45.995 ;
        RECT 95.135 -55.155 95.415 -45.015 ;
        RECT 95.695 -55.435 95.975 -45.995 ;
        RECT 96.255 -55.155 96.535 -41.655 ;
        RECT 97.315 -45.015 97.715 -43.815 ;
        RECT 96.815 -55.435 97.095 -45.995 ;
        RECT 97.375 -55.155 97.655 -45.015 ;
        RECT 98.495 -45.405 100.455 -45.005 ;
        RECT 97.935 -55.435 98.215 -45.995 ;
        RECT 98.495 -54.995 98.775 -45.405 ;
        RECT 99.055 -55.435 99.335 -45.995 ;
        RECT 99.615 -54.995 99.895 -45.405 ;
        RECT 100.175 -55.435 100.455 -45.405 ;
        RECT -477.745 -55.595 100.455 -55.435 ;
        RECT 124.705 -55.595 125.505 -9.550 ;
        RECT 183.905 -10.685 184.805 -10.305 ;
        RECT 168.340 -11.185 190.340 -10.685 ;
        RECT 169.120 -20.625 169.400 -11.185 ;
        RECT 170.240 -20.625 170.520 -11.185 ;
        RECT 170.800 -21.240 171.080 -11.625 ;
        RECT 171.360 -20.625 171.640 -11.185 ;
        RECT 171.920 -21.240 172.200 -11.625 ;
        RECT 172.480 -20.625 172.760 -11.185 ;
        RECT 173.040 -21.240 173.320 -11.625 ;
        RECT 173.600 -20.625 173.880 -11.185 ;
        RECT 174.160 -21.240 174.440 -11.625 ;
        RECT 174.720 -20.625 175.000 -11.185 ;
        RECT 175.280 -21.240 175.560 -11.625 ;
        RECT 175.840 -20.625 176.120 -11.185 ;
        RECT 176.400 -21.240 176.680 -11.625 ;
        RECT 176.960 -20.625 177.240 -11.185 ;
        RECT 177.520 -21.240 177.800 -11.625 ;
        RECT 178.080 -20.625 178.360 -11.185 ;
        RECT 178.640 -21.240 178.920 -11.625 ;
        RECT 179.200 -20.625 179.480 -11.185 ;
        RECT 179.760 -21.240 180.040 -11.625 ;
        RECT 180.320 -20.625 180.600 -11.185 ;
        RECT 180.880 -21.240 181.160 -11.625 ;
        RECT 181.440 -20.625 181.720 -11.185 ;
        RECT 182.000 -21.240 182.280 -11.625 ;
        RECT 182.560 -20.625 182.840 -11.185 ;
        RECT 183.120 -21.240 183.400 -11.625 ;
        RECT 183.680 -20.625 183.960 -11.185 ;
        RECT 184.240 -21.240 184.520 -11.625 ;
        RECT 184.800 -20.625 185.080 -11.185 ;
        RECT 185.360 -21.240 185.640 -11.625 ;
        RECT 185.920 -20.625 186.200 -11.185 ;
        RECT 186.480 -21.240 186.760 -11.625 ;
        RECT 187.040 -20.625 187.320 -11.185 ;
        RECT 187.600 -21.240 187.880 -11.625 ;
        RECT 188.160 -20.625 188.440 -11.185 ;
        RECT 189.280 -20.625 189.560 -11.185 ;
        RECT 230.275 -11.465 230.655 -9.450 ;
        RECT 233.790 -11.465 234.170 -9.450 ;
        RECT 270.200 -15.940 289.200 -14.940 ;
        RECT 298.860 -15.630 299.140 -13.010 ;
        RECT 299.980 -15.070 300.260 27.310 ;
        RECT 302.780 25.670 303.060 26.190 ;
        RECT 302.780 18.950 303.060 19.470 ;
        RECT 302.220 7.190 302.500 7.710 ;
        RECT 301.660 2.850 301.940 3.790 ;
        RECT 303.340 0.940 303.620 30.670 ;
        RECT 306.140 12.140 306.420 12.190 ;
        RECT 306.140 11.860 308.100 12.140 ;
        RECT 306.140 11.810 306.420 11.860 ;
        RECT 305.580 7.190 305.860 7.710 ;
        RECT 303.900 6.630 304.180 7.150 ;
        RECT 307.260 6.770 307.540 11.070 ;
        RECT 307.820 10.740 308.100 11.860 ;
        RECT 308.380 11.110 308.660 11.630 ;
        RECT 307.820 10.460 308.660 10.740 ;
        RECT 308.380 5.090 308.660 10.460 ;
        RECT 303.900 4.390 304.180 4.910 ;
        RECT 306.140 3.830 306.420 4.350 ;
        RECT 303.340 0.660 304.180 0.940 ;
        RECT 300.540 -4.430 300.820 -2.930 ;
        RECT 170.740 -22.350 171.140 -21.240 ;
        RECT 170.750 -23.250 171.130 -22.350 ;
        RECT 171.860 -24.350 172.260 -21.240 ;
        RECT 172.980 -22.350 173.380 -21.240 ;
        RECT 172.990 -23.250 173.370 -22.350 ;
        RECT 171.870 -25.250 172.250 -24.350 ;
        RECT 174.100 -26.350 174.500 -21.240 ;
        RECT 175.220 -22.350 175.620 -21.240 ;
        RECT 175.230 -23.250 175.610 -22.350 ;
        RECT 176.340 -24.350 176.740 -21.240 ;
        RECT 177.460 -22.350 177.860 -21.240 ;
        RECT 177.470 -23.250 177.850 -22.350 ;
        RECT 176.350 -25.250 176.730 -24.350 ;
        RECT 174.110 -27.250 174.490 -26.350 ;
        RECT 178.580 -28.740 178.980 -21.240 ;
        RECT 179.700 -28.740 180.100 -21.240 ;
        RECT 180.820 -22.350 181.220 -21.240 ;
        RECT 180.830 -23.250 181.210 -22.350 ;
        RECT 181.940 -24.350 182.340 -21.240 ;
        RECT 183.060 -22.350 183.460 -21.240 ;
        RECT 183.070 -23.250 183.450 -22.350 ;
        RECT 181.950 -25.250 182.330 -24.350 ;
        RECT 184.180 -26.350 184.580 -21.240 ;
        RECT 185.300 -22.350 185.700 -21.240 ;
        RECT 185.310 -23.250 185.690 -22.350 ;
        RECT 186.420 -24.350 186.820 -21.240 ;
        RECT 187.540 -22.350 187.940 -21.240 ;
        RECT 187.550 -23.250 187.930 -22.350 ;
        RECT 186.430 -25.250 186.810 -24.350 ;
        RECT 184.190 -27.250 184.570 -26.350 ;
        RECT 178.590 -29.640 178.970 -28.740 ;
        RECT 179.710 -29.640 180.090 -28.740 ;
        RECT 168.115 -43.750 168.495 -34.250 ;
        RECT 174.115 -42.250 174.495 -34.250 ;
        RECT 178.045 -40.750 178.425 -34.315 ;
        RECT 180.185 -39.250 180.565 -34.315 ;
        RECT 186.615 -37.750 186.995 -34.250 ;
        RECT 270.200 -37.750 271.200 -15.940 ;
        RECT 300.540 -16.420 300.820 -16.370 ;
        RECT 300.540 -16.700 301.380 -16.420 ;
        RECT 300.540 -16.750 300.820 -16.700 ;
        RECT 298.300 -20.810 298.580 -20.290 ;
        RECT 186.615 -38.250 271.200 -37.750 ;
        RECT 274.700 -26.020 289.200 -25.020 ;
        RECT 298.860 -25.710 299.140 -23.090 ;
        RECT 274.700 -39.250 275.700 -26.020 ;
        RECT 299.420 -27.620 299.700 -27.570 ;
        RECT 299.420 -27.900 300.260 -27.620 ;
        RECT 299.420 -27.950 299.700 -27.900 ;
        RECT 180.185 -39.750 275.700 -39.250 ;
        RECT 279.200 -36.100 289.200 -35.100 ;
        RECT 299.980 -35.460 300.260 -27.900 ;
        RECT 300.540 -30.190 300.820 -19.730 ;
        RECT 301.100 -24.030 301.380 -16.700 ;
        RECT 302.780 -17.310 303.060 -15.810 ;
        RECT 303.900 -16.890 304.180 0.660 ;
        RECT 304.460 -20.250 304.740 0.430 ;
        RECT 305.020 -0.510 305.300 0.990 ;
        RECT 305.580 -8.350 305.860 -1.250 ;
        RECT 308.380 -8.490 308.660 -7.970 ;
        RECT 308.380 -11.940 308.660 -11.890 ;
        RECT 306.140 -12.220 308.660 -11.940 ;
        RECT 306.140 -15.070 306.420 -12.220 ;
        RECT 308.380 -12.270 308.660 -12.220 ;
        RECT 305.580 -15.770 305.860 -15.250 ;
        RECT 308.380 -15.300 308.660 -15.250 ;
        RECT 308.940 -15.300 309.220 9.950 ;
        RECT 309.500 3.740 309.780 46.580 ;
        RECT 310.060 46.530 310.340 46.580 ;
        RECT 310.620 42.940 310.900 42.990 ;
        RECT 312.300 42.940 312.580 42.990 ;
        RECT 310.620 42.660 312.580 42.940 ;
        RECT 310.620 42.610 310.900 42.660 ;
        RECT 312.300 42.610 312.580 42.660 ;
        RECT 310.620 34.770 310.900 41.870 ;
        RECT 312.860 35.940 313.140 42.430 ;
        RECT 315.100 42.380 315.380 42.430 ;
        RECT 317.340 42.380 317.620 42.430 ;
        RECT 315.100 42.100 317.620 42.380 ;
        RECT 314.540 41.350 314.820 41.870 ;
        RECT 315.100 35.940 315.380 42.100 ;
        RECT 317.340 42.050 317.620 42.100 ;
        RECT 312.860 35.660 313.700 35.940 ;
        RECT 310.620 15.500 310.900 15.550 ;
        RECT 312.860 15.500 313.140 15.550 ;
        RECT 310.620 15.220 313.140 15.500 ;
        RECT 310.060 8.780 310.340 10.510 ;
        RECT 310.620 9.570 310.900 15.220 ;
        RECT 312.860 15.170 313.140 15.220 ;
        RECT 312.300 11.020 312.580 11.630 ;
        RECT 311.180 10.740 312.580 11.020 ;
        RECT 311.180 10.460 313.140 10.740 ;
        RECT 311.180 8.780 311.460 8.830 ;
        RECT 312.860 8.780 313.140 10.460 ;
        RECT 310.060 8.500 310.900 8.780 ;
        RECT 310.620 7.330 310.900 8.500 ;
        RECT 311.180 8.500 313.140 8.780 ;
        RECT 311.180 8.450 311.460 8.500 ;
        RECT 310.060 6.630 310.340 7.150 ;
        RECT 312.860 6.070 313.140 6.590 ;
        RECT 311.180 3.970 311.460 5.470 ;
        RECT 310.060 3.740 310.340 3.790 ;
        RECT 309.500 3.460 310.340 3.740 ;
        RECT 308.380 -15.580 309.220 -15.300 ;
        RECT 308.380 -15.770 308.660 -15.580 ;
        RECT 306.700 -23.470 306.980 -19.730 ;
        RECT 308.380 -24.170 308.660 -23.650 ;
        RECT 301.660 -30.750 301.940 -27.570 ;
        RECT 300.540 -35.460 300.820 -35.410 ;
        RECT 299.980 -35.740 300.820 -35.460 ;
        RECT 300.540 -35.790 300.820 -35.740 ;
        RECT 301.660 -35.790 301.940 -32.050 ;
        RECT 303.900 -35.790 304.180 -30.930 ;
        RECT 279.200 -40.750 280.200 -36.100 ;
        RECT 178.045 -41.250 280.200 -40.750 ;
        RECT 305.580 -40.500 305.860 -40.450 ;
        RECT 305.580 -40.780 306.420 -40.500 ;
        RECT 305.580 -40.830 305.860 -40.780 ;
        RECT 174.115 -42.750 280.200 -42.250 ;
        RECT 168.115 -44.250 275.700 -43.750 ;
        RECT -483.245 -56.095 125.505 -55.595 ;
        RECT 274.700 -55.260 275.700 -44.250 ;
        RECT 279.200 -45.180 280.200 -42.750 ;
        RECT 298.860 -44.890 299.140 -44.370 ;
        RECT 279.200 -46.180 289.200 -45.180 ;
        RECT 300.540 -48.060 300.820 -46.610 ;
        RECT 298.300 -48.340 300.820 -48.060 ;
        RECT -483.245 -79.275 -482.495 -56.095 ;
        RECT -477.745 -56.255 100.455 -56.095 ;
        RECT -477.745 -66.285 -477.465 -56.255 ;
        RECT -477.185 -66.285 -476.905 -56.695 ;
        RECT -476.625 -65.695 -476.345 -56.255 ;
        RECT -476.065 -66.285 -475.785 -56.695 ;
        RECT -475.505 -65.695 -475.225 -56.255 ;
        RECT -477.745 -66.685 -475.785 -66.285 ;
        RECT -474.945 -66.675 -474.665 -56.535 ;
        RECT -474.385 -65.695 -474.105 -56.255 ;
        RECT -475.005 -67.875 -474.605 -66.675 ;
        RECT -473.825 -70.035 -473.545 -56.535 ;
        RECT -473.265 -65.695 -472.985 -56.255 ;
        RECT -472.705 -66.675 -472.425 -56.535 ;
        RECT -472.145 -65.695 -471.865 -56.255 ;
        RECT -472.765 -67.875 -472.365 -66.675 ;
        RECT -473.885 -71.235 -473.485 -70.035 ;
        RECT -471.585 -73.395 -471.305 -56.535 ;
        RECT -471.025 -65.695 -470.745 -56.255 ;
        RECT -470.465 -66.675 -470.185 -56.535 ;
        RECT -469.905 -65.695 -469.625 -56.255 ;
        RECT -470.525 -67.875 -470.125 -66.675 ;
        RECT -469.345 -70.035 -469.065 -56.535 ;
        RECT -468.785 -65.695 -468.505 -56.255 ;
        RECT -468.225 -66.675 -467.945 -56.535 ;
        RECT -467.665 -65.695 -467.385 -56.255 ;
        RECT -468.285 -67.875 -467.885 -66.675 ;
        RECT -469.405 -71.235 -469.005 -70.035 ;
        RECT -471.645 -74.595 -471.245 -73.395 ;
        RECT -467.105 -76.755 -466.825 -56.535 ;
        RECT -466.545 -65.695 -466.265 -56.255 ;
        RECT -465.985 -66.675 -465.705 -56.535 ;
        RECT -465.425 -65.695 -465.145 -56.255 ;
        RECT -466.045 -67.875 -465.645 -66.675 ;
        RECT -464.865 -70.035 -464.585 -56.535 ;
        RECT -464.305 -65.695 -464.025 -56.255 ;
        RECT -463.745 -66.675 -463.465 -56.535 ;
        RECT -463.185 -65.695 -462.905 -56.255 ;
        RECT -463.805 -67.875 -463.405 -66.675 ;
        RECT -464.925 -71.235 -464.525 -70.035 ;
        RECT -462.625 -73.395 -462.345 -56.535 ;
        RECT -462.065 -65.695 -461.785 -56.255 ;
        RECT -461.505 -66.675 -461.225 -56.535 ;
        RECT -460.945 -65.695 -460.665 -56.255 ;
        RECT -461.565 -67.875 -461.165 -66.675 ;
        RECT -460.385 -70.035 -460.105 -56.535 ;
        RECT -459.825 -65.695 -459.545 -56.255 ;
        RECT -459.265 -66.675 -458.985 -56.535 ;
        RECT -458.705 -65.695 -458.425 -56.255 ;
        RECT -459.325 -67.875 -458.925 -66.675 ;
        RECT -460.445 -71.235 -460.045 -70.035 ;
        RECT -462.685 -74.595 -462.285 -73.395 ;
        RECT -467.165 -77.955 -466.765 -76.755 ;
        RECT -484.745 -79.655 -482.495 -79.275 ;
        RECT -458.145 -80.115 -457.865 -56.535 ;
        RECT -457.585 -65.695 -457.305 -56.255 ;
        RECT -457.025 -66.675 -456.745 -56.535 ;
        RECT -456.465 -65.695 -456.185 -56.255 ;
        RECT -457.085 -67.875 -456.685 -66.675 ;
        RECT -455.905 -70.035 -455.625 -56.535 ;
        RECT -455.345 -65.695 -455.065 -56.255 ;
        RECT -454.785 -66.675 -454.505 -56.535 ;
        RECT -454.225 -65.695 -453.945 -56.255 ;
        RECT -454.845 -67.875 -454.445 -66.675 ;
        RECT -455.965 -71.235 -455.565 -70.035 ;
        RECT -453.665 -73.395 -453.385 -56.535 ;
        RECT -453.105 -65.695 -452.825 -56.255 ;
        RECT -452.545 -66.675 -452.265 -56.535 ;
        RECT -451.985 -65.695 -451.705 -56.255 ;
        RECT -452.605 -67.875 -452.205 -66.675 ;
        RECT -451.425 -70.035 -451.145 -56.535 ;
        RECT -450.865 -65.695 -450.585 -56.255 ;
        RECT -450.305 -66.675 -450.025 -56.535 ;
        RECT -449.745 -65.695 -449.465 -56.255 ;
        RECT -450.365 -67.875 -449.965 -66.675 ;
        RECT -451.485 -71.235 -451.085 -70.035 ;
        RECT -453.725 -74.595 -453.325 -73.395 ;
        RECT -449.185 -76.755 -448.905 -56.535 ;
        RECT -448.625 -65.695 -448.345 -56.255 ;
        RECT -448.065 -66.675 -447.785 -56.535 ;
        RECT -447.505 -65.695 -447.225 -56.255 ;
        RECT -448.125 -67.875 -447.725 -66.675 ;
        RECT -446.945 -70.035 -446.665 -56.535 ;
        RECT -446.385 -65.695 -446.105 -56.255 ;
        RECT -445.825 -66.675 -445.545 -56.535 ;
        RECT -445.265 -65.695 -444.985 -56.255 ;
        RECT -445.885 -67.875 -445.485 -66.675 ;
        RECT -447.005 -71.235 -446.605 -70.035 ;
        RECT -444.705 -73.395 -444.425 -56.535 ;
        RECT -444.145 -65.695 -443.865 -56.255 ;
        RECT -443.585 -66.675 -443.305 -56.535 ;
        RECT -443.025 -65.695 -442.745 -56.255 ;
        RECT -443.645 -67.875 -443.245 -66.675 ;
        RECT -442.465 -70.035 -442.185 -56.535 ;
        RECT -441.905 -65.695 -441.625 -56.255 ;
        RECT -441.345 -66.675 -441.065 -56.535 ;
        RECT -440.785 -65.695 -440.505 -56.255 ;
        RECT -441.405 -67.875 -441.005 -66.675 ;
        RECT -442.525 -71.235 -442.125 -70.035 ;
        RECT -444.765 -74.595 -444.365 -73.395 ;
        RECT -449.245 -77.955 -448.845 -76.755 ;
        RECT -486.955 -83.235 -486.555 -81.155 ;
        RECT -458.205 -81.315 -457.805 -80.115 ;
        RECT -497.595 -83.765 -495.515 -83.365 ;
        RECT -440.225 -83.475 -439.945 -56.535 ;
        RECT -439.665 -65.695 -439.385 -56.255 ;
        RECT -439.105 -66.675 -438.825 -56.535 ;
        RECT -438.545 -65.695 -438.265 -56.255 ;
        RECT -439.165 -67.875 -438.765 -66.675 ;
        RECT -437.985 -70.035 -437.705 -56.535 ;
        RECT -437.425 -65.695 -437.145 -56.255 ;
        RECT -436.865 -66.675 -436.585 -56.535 ;
        RECT -436.305 -65.695 -436.025 -56.255 ;
        RECT -436.925 -67.875 -436.525 -66.675 ;
        RECT -438.045 -71.235 -437.645 -70.035 ;
        RECT -435.745 -73.395 -435.465 -56.535 ;
        RECT -435.185 -65.695 -434.905 -56.255 ;
        RECT -434.625 -66.675 -434.345 -56.535 ;
        RECT -434.065 -65.695 -433.785 -56.255 ;
        RECT -434.685 -67.875 -434.285 -66.675 ;
        RECT -433.505 -70.035 -433.225 -56.535 ;
        RECT -432.945 -65.695 -432.665 -56.255 ;
        RECT -432.385 -66.675 -432.105 -56.535 ;
        RECT -431.825 -65.695 -431.545 -56.255 ;
        RECT -432.445 -67.875 -432.045 -66.675 ;
        RECT -433.565 -71.235 -433.165 -70.035 ;
        RECT -435.805 -74.595 -435.405 -73.395 ;
        RECT -431.265 -76.755 -430.985 -56.535 ;
        RECT -430.705 -65.695 -430.425 -56.255 ;
        RECT -430.145 -66.675 -429.865 -56.535 ;
        RECT -429.585 -65.695 -429.305 -56.255 ;
        RECT -430.205 -67.875 -429.805 -66.675 ;
        RECT -429.025 -70.035 -428.745 -56.535 ;
        RECT -428.465 -65.695 -428.185 -56.255 ;
        RECT -427.905 -66.675 -427.625 -56.535 ;
        RECT -427.345 -65.695 -427.065 -56.255 ;
        RECT -427.965 -67.875 -427.565 -66.675 ;
        RECT -429.085 -71.235 -428.685 -70.035 ;
        RECT -426.785 -73.395 -426.505 -56.535 ;
        RECT -426.225 -65.695 -425.945 -56.255 ;
        RECT -425.665 -66.675 -425.385 -56.535 ;
        RECT -425.105 -65.695 -424.825 -56.255 ;
        RECT -425.725 -67.875 -425.325 -66.675 ;
        RECT -424.545 -70.035 -424.265 -56.535 ;
        RECT -423.985 -65.695 -423.705 -56.255 ;
        RECT -423.425 -66.675 -423.145 -56.535 ;
        RECT -422.865 -65.695 -422.585 -56.255 ;
        RECT -423.485 -67.875 -423.085 -66.675 ;
        RECT -424.605 -71.235 -424.205 -70.035 ;
        RECT -426.845 -74.595 -426.445 -73.395 ;
        RECT -431.325 -77.955 -430.925 -76.755 ;
        RECT -422.305 -80.115 -422.025 -56.535 ;
        RECT -421.745 -65.695 -421.465 -56.255 ;
        RECT -421.185 -66.675 -420.905 -56.535 ;
        RECT -420.625 -65.695 -420.345 -56.255 ;
        RECT -421.245 -67.875 -420.845 -66.675 ;
        RECT -420.065 -70.035 -419.785 -56.535 ;
        RECT -419.505 -65.695 -419.225 -56.255 ;
        RECT -418.945 -66.675 -418.665 -56.535 ;
        RECT -418.385 -65.695 -418.105 -56.255 ;
        RECT -419.005 -67.875 -418.605 -66.675 ;
        RECT -420.125 -71.235 -419.725 -70.035 ;
        RECT -417.825 -73.395 -417.545 -56.535 ;
        RECT -417.265 -65.695 -416.985 -56.255 ;
        RECT -416.705 -66.675 -416.425 -56.535 ;
        RECT -416.145 -65.695 -415.865 -56.255 ;
        RECT -416.765 -67.875 -416.365 -66.675 ;
        RECT -415.585 -70.035 -415.305 -56.535 ;
        RECT -415.025 -65.695 -414.745 -56.255 ;
        RECT -414.465 -66.675 -414.185 -56.535 ;
        RECT -413.905 -65.695 -413.625 -56.255 ;
        RECT -414.525 -67.875 -414.125 -66.675 ;
        RECT -415.645 -71.235 -415.245 -70.035 ;
        RECT -417.885 -74.595 -417.485 -73.395 ;
        RECT -413.345 -76.755 -413.065 -56.535 ;
        RECT -412.785 -65.695 -412.505 -56.255 ;
        RECT -412.225 -66.675 -411.945 -56.535 ;
        RECT -411.665 -65.695 -411.385 -56.255 ;
        RECT -412.285 -67.875 -411.885 -66.675 ;
        RECT -411.105 -70.035 -410.825 -56.535 ;
        RECT -410.545 -65.695 -410.265 -56.255 ;
        RECT -409.985 -66.675 -409.705 -56.535 ;
        RECT -409.425 -65.695 -409.145 -56.255 ;
        RECT -410.045 -67.875 -409.645 -66.675 ;
        RECT -411.165 -71.235 -410.765 -70.035 ;
        RECT -408.865 -73.395 -408.585 -56.535 ;
        RECT -408.305 -65.695 -408.025 -56.255 ;
        RECT -407.745 -66.675 -407.465 -56.535 ;
        RECT -407.185 -65.695 -406.905 -56.255 ;
        RECT -407.805 -67.875 -407.405 -66.675 ;
        RECT -406.625 -70.035 -406.345 -56.535 ;
        RECT -406.065 -65.695 -405.785 -56.255 ;
        RECT -405.505 -66.675 -405.225 -56.535 ;
        RECT -404.945 -65.695 -404.665 -56.255 ;
        RECT -405.565 -67.875 -405.165 -66.675 ;
        RECT -406.685 -71.235 -406.285 -70.035 ;
        RECT -408.925 -74.595 -408.525 -73.395 ;
        RECT -413.405 -77.955 -413.005 -76.755 ;
        RECT -422.365 -81.315 -421.965 -80.115 ;
        RECT -492.330 -84.775 -490.235 -84.395 ;
        RECT -440.285 -84.675 -439.885 -83.475 ;
        RECT -490.615 -90.135 -490.235 -84.775 ;
        RECT -404.385 -86.835 -404.105 -56.535 ;
        RECT -403.825 -65.695 -403.545 -56.255 ;
        RECT -403.265 -66.675 -402.985 -56.535 ;
        RECT -402.705 -65.695 -402.425 -56.255 ;
        RECT -403.325 -67.875 -402.925 -66.675 ;
        RECT -402.145 -70.035 -401.865 -56.535 ;
        RECT -401.585 -65.695 -401.305 -56.255 ;
        RECT -401.025 -66.675 -400.745 -56.535 ;
        RECT -400.465 -65.695 -400.185 -56.255 ;
        RECT -401.085 -67.875 -400.685 -66.675 ;
        RECT -402.205 -71.235 -401.805 -70.035 ;
        RECT -399.905 -73.395 -399.625 -56.535 ;
        RECT -399.345 -65.695 -399.065 -56.255 ;
        RECT -398.785 -66.675 -398.505 -56.535 ;
        RECT -398.225 -65.695 -397.945 -56.255 ;
        RECT -398.845 -67.875 -398.445 -66.675 ;
        RECT -397.665 -70.035 -397.385 -56.535 ;
        RECT -397.105 -65.695 -396.825 -56.255 ;
        RECT -396.545 -66.675 -396.265 -56.535 ;
        RECT -395.985 -65.695 -395.705 -56.255 ;
        RECT -396.605 -67.875 -396.205 -66.675 ;
        RECT -397.725 -71.235 -397.325 -70.035 ;
        RECT -399.965 -74.595 -399.565 -73.395 ;
        RECT -395.425 -76.755 -395.145 -56.535 ;
        RECT -394.865 -65.695 -394.585 -56.255 ;
        RECT -394.305 -66.675 -394.025 -56.535 ;
        RECT -393.745 -65.695 -393.465 -56.255 ;
        RECT -394.365 -67.875 -393.965 -66.675 ;
        RECT -393.185 -70.035 -392.905 -56.535 ;
        RECT -392.625 -65.695 -392.345 -56.255 ;
        RECT -392.065 -66.675 -391.785 -56.535 ;
        RECT -391.505 -65.695 -391.225 -56.255 ;
        RECT -392.125 -67.875 -391.725 -66.675 ;
        RECT -393.245 -71.235 -392.845 -70.035 ;
        RECT -390.945 -73.395 -390.665 -56.535 ;
        RECT -390.385 -65.695 -390.105 -56.255 ;
        RECT -389.825 -66.675 -389.545 -56.535 ;
        RECT -389.265 -65.695 -388.985 -56.255 ;
        RECT -389.885 -67.875 -389.485 -66.675 ;
        RECT -388.705 -70.035 -388.425 -56.535 ;
        RECT -388.145 -65.695 -387.865 -56.255 ;
        RECT -387.585 -66.675 -387.305 -56.535 ;
        RECT -387.025 -65.695 -386.745 -56.255 ;
        RECT -387.645 -67.875 -387.245 -66.675 ;
        RECT -388.765 -71.235 -388.365 -70.035 ;
        RECT -391.005 -74.595 -390.605 -73.395 ;
        RECT -395.485 -77.955 -395.085 -76.755 ;
        RECT -386.465 -80.115 -386.185 -56.535 ;
        RECT -385.905 -65.695 -385.625 -56.255 ;
        RECT -385.345 -66.675 -385.065 -56.535 ;
        RECT -384.785 -65.695 -384.505 -56.255 ;
        RECT -385.405 -67.875 -385.005 -66.675 ;
        RECT -384.225 -70.035 -383.945 -56.535 ;
        RECT -383.665 -65.695 -383.385 -56.255 ;
        RECT -383.105 -66.675 -382.825 -56.535 ;
        RECT -382.545 -65.695 -382.265 -56.255 ;
        RECT -383.165 -67.875 -382.765 -66.675 ;
        RECT -384.285 -71.235 -383.885 -70.035 ;
        RECT -381.985 -73.395 -381.705 -56.535 ;
        RECT -381.425 -65.695 -381.145 -56.255 ;
        RECT -380.865 -66.675 -380.585 -56.535 ;
        RECT -380.305 -65.695 -380.025 -56.255 ;
        RECT -380.925 -67.875 -380.525 -66.675 ;
        RECT -379.745 -70.035 -379.465 -56.535 ;
        RECT -379.185 -65.695 -378.905 -56.255 ;
        RECT -378.625 -66.675 -378.345 -56.535 ;
        RECT -378.065 -65.695 -377.785 -56.255 ;
        RECT -378.685 -67.875 -378.285 -66.675 ;
        RECT -379.805 -71.235 -379.405 -70.035 ;
        RECT -382.045 -74.595 -381.645 -73.395 ;
        RECT -377.505 -76.755 -377.225 -56.535 ;
        RECT -376.945 -65.695 -376.665 -56.255 ;
        RECT -376.385 -66.675 -376.105 -56.535 ;
        RECT -375.825 -65.695 -375.545 -56.255 ;
        RECT -376.445 -67.875 -376.045 -66.675 ;
        RECT -375.265 -70.035 -374.985 -56.535 ;
        RECT -374.705 -65.695 -374.425 -56.255 ;
        RECT -374.145 -66.675 -373.865 -56.535 ;
        RECT -373.585 -65.695 -373.305 -56.255 ;
        RECT -374.205 -67.875 -373.805 -66.675 ;
        RECT -375.325 -71.235 -374.925 -70.035 ;
        RECT -373.025 -73.395 -372.745 -56.535 ;
        RECT -372.465 -65.695 -372.185 -56.255 ;
        RECT -371.905 -66.675 -371.625 -56.535 ;
        RECT -371.345 -65.695 -371.065 -56.255 ;
        RECT -371.965 -67.875 -371.565 -66.675 ;
        RECT -370.785 -70.035 -370.505 -56.535 ;
        RECT -370.225 -65.695 -369.945 -56.255 ;
        RECT -369.665 -66.675 -369.385 -56.535 ;
        RECT -369.105 -65.695 -368.825 -56.255 ;
        RECT -369.725 -67.875 -369.325 -66.675 ;
        RECT -370.845 -71.235 -370.445 -70.035 ;
        RECT -373.085 -74.595 -372.685 -73.395 ;
        RECT -377.565 -77.955 -377.165 -76.755 ;
        RECT -386.525 -81.315 -386.125 -80.115 ;
        RECT -368.545 -83.475 -368.265 -56.535 ;
        RECT -367.985 -65.695 -367.705 -56.255 ;
        RECT -367.425 -66.675 -367.145 -56.535 ;
        RECT -366.865 -65.695 -366.585 -56.255 ;
        RECT -367.485 -67.875 -367.085 -66.675 ;
        RECT -366.305 -70.035 -366.025 -56.535 ;
        RECT -365.745 -65.695 -365.465 -56.255 ;
        RECT -365.185 -66.675 -364.905 -56.535 ;
        RECT -364.625 -65.695 -364.345 -56.255 ;
        RECT -365.245 -67.875 -364.845 -66.675 ;
        RECT -366.365 -71.235 -365.965 -70.035 ;
        RECT -364.065 -73.395 -363.785 -56.535 ;
        RECT -363.505 -65.695 -363.225 -56.255 ;
        RECT -362.945 -66.675 -362.665 -56.535 ;
        RECT -362.385 -65.695 -362.105 -56.255 ;
        RECT -363.005 -67.875 -362.605 -66.675 ;
        RECT -361.825 -70.035 -361.545 -56.535 ;
        RECT -361.265 -65.695 -360.985 -56.255 ;
        RECT -360.705 -66.675 -360.425 -56.535 ;
        RECT -360.145 -65.695 -359.865 -56.255 ;
        RECT -360.765 -67.875 -360.365 -66.675 ;
        RECT -361.885 -71.235 -361.485 -70.035 ;
        RECT -364.125 -74.595 -363.725 -73.395 ;
        RECT -359.585 -76.755 -359.305 -56.535 ;
        RECT -359.025 -65.695 -358.745 -56.255 ;
        RECT -358.465 -66.675 -358.185 -56.535 ;
        RECT -357.905 -65.695 -357.625 -56.255 ;
        RECT -358.525 -67.875 -358.125 -66.675 ;
        RECT -357.345 -70.035 -357.065 -56.535 ;
        RECT -356.785 -65.695 -356.505 -56.255 ;
        RECT -356.225 -66.675 -355.945 -56.535 ;
        RECT -355.665 -65.695 -355.385 -56.255 ;
        RECT -356.285 -67.875 -355.885 -66.675 ;
        RECT -357.405 -71.235 -357.005 -70.035 ;
        RECT -355.105 -73.395 -354.825 -56.535 ;
        RECT -354.545 -65.695 -354.265 -56.255 ;
        RECT -353.985 -66.675 -353.705 -56.535 ;
        RECT -353.425 -65.695 -353.145 -56.255 ;
        RECT -354.045 -67.875 -353.645 -66.675 ;
        RECT -352.865 -70.035 -352.585 -56.535 ;
        RECT -352.305 -65.695 -352.025 -56.255 ;
        RECT -351.745 -66.675 -351.465 -56.535 ;
        RECT -351.185 -65.695 -350.905 -56.255 ;
        RECT -351.805 -67.875 -351.405 -66.675 ;
        RECT -352.925 -71.235 -352.525 -70.035 ;
        RECT -355.165 -74.595 -354.765 -73.395 ;
        RECT -359.645 -77.955 -359.245 -76.755 ;
        RECT -350.625 -80.115 -350.345 -56.535 ;
        RECT -350.065 -65.695 -349.785 -56.255 ;
        RECT -349.505 -66.675 -349.225 -56.535 ;
        RECT -348.945 -65.695 -348.665 -56.255 ;
        RECT -349.565 -67.875 -349.165 -66.675 ;
        RECT -348.385 -70.035 -348.105 -56.535 ;
        RECT -347.825 -65.695 -347.545 -56.255 ;
        RECT -347.265 -66.675 -346.985 -56.535 ;
        RECT -346.705 -65.695 -346.425 -56.255 ;
        RECT -347.325 -67.875 -346.925 -66.675 ;
        RECT -348.445 -71.235 -348.045 -70.035 ;
        RECT -346.145 -73.395 -345.865 -56.535 ;
        RECT -345.585 -65.695 -345.305 -56.255 ;
        RECT -345.025 -66.675 -344.745 -56.535 ;
        RECT -344.465 -65.695 -344.185 -56.255 ;
        RECT -345.085 -67.875 -344.685 -66.675 ;
        RECT -343.905 -70.035 -343.625 -56.535 ;
        RECT -343.345 -65.695 -343.065 -56.255 ;
        RECT -342.785 -66.675 -342.505 -56.535 ;
        RECT -342.225 -65.695 -341.945 -56.255 ;
        RECT -342.845 -67.875 -342.445 -66.675 ;
        RECT -343.965 -71.235 -343.565 -70.035 ;
        RECT -346.205 -74.595 -345.805 -73.395 ;
        RECT -341.665 -76.755 -341.385 -56.535 ;
        RECT -341.105 -65.695 -340.825 -56.255 ;
        RECT -340.545 -66.675 -340.265 -56.535 ;
        RECT -339.985 -65.695 -339.705 -56.255 ;
        RECT -340.605 -67.875 -340.205 -66.675 ;
        RECT -339.425 -70.035 -339.145 -56.535 ;
        RECT -338.865 -65.695 -338.585 -56.255 ;
        RECT -338.305 -66.675 -338.025 -56.535 ;
        RECT -337.745 -65.695 -337.465 -56.255 ;
        RECT -338.365 -67.875 -337.965 -66.675 ;
        RECT -339.485 -71.235 -339.085 -70.035 ;
        RECT -337.185 -73.395 -336.905 -56.535 ;
        RECT -336.625 -65.695 -336.345 -56.255 ;
        RECT -336.065 -66.675 -335.785 -56.535 ;
        RECT -335.505 -65.695 -335.225 -56.255 ;
        RECT -336.125 -67.875 -335.725 -66.675 ;
        RECT -334.945 -70.035 -334.665 -56.535 ;
        RECT -334.385 -65.695 -334.105 -56.255 ;
        RECT -333.825 -66.675 -333.545 -56.535 ;
        RECT -333.265 -65.695 -332.985 -56.255 ;
        RECT -333.885 -67.875 -333.485 -66.675 ;
        RECT -335.005 -71.235 -334.605 -70.035 ;
        RECT -337.245 -74.595 -336.845 -73.395 ;
        RECT -341.725 -77.955 -341.325 -76.755 ;
        RECT -350.685 -81.315 -350.285 -80.115 ;
        RECT -368.605 -84.675 -368.205 -83.475 ;
        RECT -404.445 -88.035 -404.045 -86.835 ;
        RECT -490.615 -90.515 -490.225 -90.135 ;
        RECT -332.705 -90.195 -332.425 -56.535 ;
        RECT -332.145 -65.695 -331.865 -56.255 ;
        RECT -331.585 -66.675 -331.305 -56.535 ;
        RECT -331.025 -65.695 -330.745 -56.255 ;
        RECT -331.645 -67.875 -331.245 -66.675 ;
        RECT -330.465 -70.035 -330.185 -56.535 ;
        RECT -329.905 -65.695 -329.625 -56.255 ;
        RECT -329.345 -66.675 -329.065 -56.535 ;
        RECT -328.785 -65.695 -328.505 -56.255 ;
        RECT -329.405 -67.875 -329.005 -66.675 ;
        RECT -330.525 -71.235 -330.125 -70.035 ;
        RECT -328.225 -73.395 -327.945 -56.535 ;
        RECT -327.665 -65.695 -327.385 -56.255 ;
        RECT -327.105 -66.675 -326.825 -56.535 ;
        RECT -326.545 -65.695 -326.265 -56.255 ;
        RECT -327.165 -67.875 -326.765 -66.675 ;
        RECT -325.985 -70.035 -325.705 -56.535 ;
        RECT -325.425 -65.695 -325.145 -56.255 ;
        RECT -324.865 -66.675 -324.585 -56.535 ;
        RECT -324.305 -65.695 -324.025 -56.255 ;
        RECT -324.925 -67.875 -324.525 -66.675 ;
        RECT -326.045 -71.235 -325.645 -70.035 ;
        RECT -328.285 -74.595 -327.885 -73.395 ;
        RECT -323.745 -76.755 -323.465 -56.535 ;
        RECT -323.185 -65.695 -322.905 -56.255 ;
        RECT -322.625 -66.675 -322.345 -56.535 ;
        RECT -322.065 -65.695 -321.785 -56.255 ;
        RECT -322.685 -67.875 -322.285 -66.675 ;
        RECT -321.505 -70.035 -321.225 -56.535 ;
        RECT -320.945 -65.695 -320.665 -56.255 ;
        RECT -320.385 -66.675 -320.105 -56.535 ;
        RECT -319.825 -65.695 -319.545 -56.255 ;
        RECT -320.445 -67.875 -320.045 -66.675 ;
        RECT -321.565 -71.235 -321.165 -70.035 ;
        RECT -319.265 -73.395 -318.985 -56.535 ;
        RECT -318.705 -65.695 -318.425 -56.255 ;
        RECT -318.145 -66.675 -317.865 -56.535 ;
        RECT -317.585 -65.695 -317.305 -56.255 ;
        RECT -318.205 -67.875 -317.805 -66.675 ;
        RECT -317.025 -70.035 -316.745 -56.535 ;
        RECT -316.465 -65.695 -316.185 -56.255 ;
        RECT -315.905 -66.675 -315.625 -56.535 ;
        RECT -315.345 -65.695 -315.065 -56.255 ;
        RECT -315.965 -67.875 -315.565 -66.675 ;
        RECT -317.085 -71.235 -316.685 -70.035 ;
        RECT -319.325 -74.595 -318.925 -73.395 ;
        RECT -323.805 -77.955 -323.405 -76.755 ;
        RECT -314.785 -80.115 -314.505 -56.535 ;
        RECT -314.225 -65.695 -313.945 -56.255 ;
        RECT -313.665 -66.675 -313.385 -56.535 ;
        RECT -313.105 -65.695 -312.825 -56.255 ;
        RECT -313.725 -67.875 -313.325 -66.675 ;
        RECT -312.545 -70.035 -312.265 -56.535 ;
        RECT -311.985 -65.695 -311.705 -56.255 ;
        RECT -311.425 -66.675 -311.145 -56.535 ;
        RECT -310.865 -65.695 -310.585 -56.255 ;
        RECT -311.485 -67.875 -311.085 -66.675 ;
        RECT -312.605 -71.235 -312.205 -70.035 ;
        RECT -310.305 -73.395 -310.025 -56.535 ;
        RECT -309.745 -65.695 -309.465 -56.255 ;
        RECT -309.185 -66.675 -308.905 -56.535 ;
        RECT -308.625 -65.695 -308.345 -56.255 ;
        RECT -309.245 -67.875 -308.845 -66.675 ;
        RECT -308.065 -70.035 -307.785 -56.535 ;
        RECT -307.505 -65.695 -307.225 -56.255 ;
        RECT -306.945 -66.675 -306.665 -56.535 ;
        RECT -306.385 -65.695 -306.105 -56.255 ;
        RECT -307.005 -67.875 -306.605 -66.675 ;
        RECT -308.125 -71.235 -307.725 -70.035 ;
        RECT -310.365 -74.595 -309.965 -73.395 ;
        RECT -305.825 -76.755 -305.545 -56.535 ;
        RECT -305.265 -65.695 -304.985 -56.255 ;
        RECT -304.705 -66.675 -304.425 -56.535 ;
        RECT -304.145 -65.695 -303.865 -56.255 ;
        RECT -304.765 -67.875 -304.365 -66.675 ;
        RECT -303.585 -70.035 -303.305 -56.535 ;
        RECT -303.025 -65.695 -302.745 -56.255 ;
        RECT -302.465 -66.675 -302.185 -56.535 ;
        RECT -301.905 -65.695 -301.625 -56.255 ;
        RECT -302.525 -67.875 -302.125 -66.675 ;
        RECT -303.645 -71.235 -303.245 -70.035 ;
        RECT -301.345 -73.395 -301.065 -56.535 ;
        RECT -300.785 -65.695 -300.505 -56.255 ;
        RECT -300.225 -66.675 -299.945 -56.535 ;
        RECT -299.665 -65.695 -299.385 -56.255 ;
        RECT -300.285 -67.875 -299.885 -66.675 ;
        RECT -299.105 -70.035 -298.825 -56.535 ;
        RECT -298.545 -65.695 -298.265 -56.255 ;
        RECT -297.985 -66.675 -297.705 -56.535 ;
        RECT -297.425 -65.695 -297.145 -56.255 ;
        RECT -298.045 -67.875 -297.645 -66.675 ;
        RECT -299.165 -71.235 -298.765 -70.035 ;
        RECT -301.405 -74.595 -301.005 -73.395 ;
        RECT -305.885 -77.955 -305.485 -76.755 ;
        RECT -314.845 -81.315 -314.445 -80.115 ;
        RECT -296.865 -83.475 -296.585 -56.535 ;
        RECT -296.305 -65.695 -296.025 -56.255 ;
        RECT -295.745 -66.675 -295.465 -56.535 ;
        RECT -295.185 -65.695 -294.905 -56.255 ;
        RECT -295.805 -67.875 -295.405 -66.675 ;
        RECT -294.625 -70.035 -294.345 -56.535 ;
        RECT -294.065 -65.695 -293.785 -56.255 ;
        RECT -293.505 -66.675 -293.225 -56.535 ;
        RECT -292.945 -65.695 -292.665 -56.255 ;
        RECT -293.565 -67.875 -293.165 -66.675 ;
        RECT -294.685 -71.235 -294.285 -70.035 ;
        RECT -292.385 -73.395 -292.105 -56.535 ;
        RECT -291.825 -65.695 -291.545 -56.255 ;
        RECT -291.265 -66.675 -290.985 -56.535 ;
        RECT -290.705 -65.695 -290.425 -56.255 ;
        RECT -291.325 -67.875 -290.925 -66.675 ;
        RECT -290.145 -70.035 -289.865 -56.535 ;
        RECT -289.585 -65.695 -289.305 -56.255 ;
        RECT -289.025 -66.675 -288.745 -56.535 ;
        RECT -288.465 -65.695 -288.185 -56.255 ;
        RECT -289.085 -67.875 -288.685 -66.675 ;
        RECT -290.205 -71.235 -289.805 -70.035 ;
        RECT -292.445 -74.595 -292.045 -73.395 ;
        RECT -287.905 -76.755 -287.625 -56.535 ;
        RECT -287.345 -65.695 -287.065 -56.255 ;
        RECT -286.785 -66.675 -286.505 -56.535 ;
        RECT -286.225 -65.695 -285.945 -56.255 ;
        RECT -286.845 -67.875 -286.445 -66.675 ;
        RECT -285.665 -70.035 -285.385 -56.535 ;
        RECT -285.105 -65.695 -284.825 -56.255 ;
        RECT -284.545 -66.675 -284.265 -56.535 ;
        RECT -283.985 -65.695 -283.705 -56.255 ;
        RECT -284.605 -67.875 -284.205 -66.675 ;
        RECT -285.725 -71.235 -285.325 -70.035 ;
        RECT -283.425 -73.395 -283.145 -56.535 ;
        RECT -282.865 -65.695 -282.585 -56.255 ;
        RECT -282.305 -66.675 -282.025 -56.535 ;
        RECT -281.745 -65.695 -281.465 -56.255 ;
        RECT -282.365 -67.875 -281.965 -66.675 ;
        RECT -281.185 -70.035 -280.905 -56.535 ;
        RECT -280.625 -65.695 -280.345 -56.255 ;
        RECT -280.065 -66.675 -279.785 -56.535 ;
        RECT -279.505 -65.695 -279.225 -56.255 ;
        RECT -280.125 -67.875 -279.725 -66.675 ;
        RECT -281.245 -71.235 -280.845 -70.035 ;
        RECT -283.485 -74.595 -283.085 -73.395 ;
        RECT -287.965 -77.955 -287.565 -76.755 ;
        RECT -278.945 -80.115 -278.665 -56.535 ;
        RECT -278.385 -65.695 -278.105 -56.255 ;
        RECT -277.825 -66.675 -277.545 -56.535 ;
        RECT -277.265 -65.695 -276.985 -56.255 ;
        RECT -277.885 -67.875 -277.485 -66.675 ;
        RECT -276.705 -70.035 -276.425 -56.535 ;
        RECT -276.145 -65.695 -275.865 -56.255 ;
        RECT -275.585 -66.675 -275.305 -56.535 ;
        RECT -275.025 -65.695 -274.745 -56.255 ;
        RECT -275.645 -67.875 -275.245 -66.675 ;
        RECT -276.765 -71.235 -276.365 -70.035 ;
        RECT -274.465 -73.395 -274.185 -56.535 ;
        RECT -273.905 -65.695 -273.625 -56.255 ;
        RECT -273.345 -66.675 -273.065 -56.535 ;
        RECT -272.785 -65.695 -272.505 -56.255 ;
        RECT -273.405 -67.875 -273.005 -66.675 ;
        RECT -272.225 -70.035 -271.945 -56.535 ;
        RECT -271.665 -65.695 -271.385 -56.255 ;
        RECT -271.105 -66.675 -270.825 -56.535 ;
        RECT -270.545 -65.695 -270.265 -56.255 ;
        RECT -271.165 -67.875 -270.765 -66.675 ;
        RECT -272.285 -71.235 -271.885 -70.035 ;
        RECT -274.525 -74.595 -274.125 -73.395 ;
        RECT -269.985 -76.755 -269.705 -56.535 ;
        RECT -269.425 -65.695 -269.145 -56.255 ;
        RECT -268.865 -66.675 -268.585 -56.535 ;
        RECT -268.305 -65.695 -268.025 -56.255 ;
        RECT -268.925 -67.875 -268.525 -66.675 ;
        RECT -267.745 -70.035 -267.465 -56.535 ;
        RECT -267.185 -65.695 -266.905 -56.255 ;
        RECT -266.625 -66.675 -266.345 -56.535 ;
        RECT -266.065 -65.695 -265.785 -56.255 ;
        RECT -266.685 -67.875 -266.285 -66.675 ;
        RECT -267.805 -71.235 -267.405 -70.035 ;
        RECT -265.505 -73.395 -265.225 -56.535 ;
        RECT -264.945 -65.695 -264.665 -56.255 ;
        RECT -264.385 -66.675 -264.105 -56.535 ;
        RECT -263.825 -65.695 -263.545 -56.255 ;
        RECT -264.445 -67.875 -264.045 -66.675 ;
        RECT -263.265 -70.035 -262.985 -56.535 ;
        RECT -262.705 -65.695 -262.425 -56.255 ;
        RECT -262.145 -66.675 -261.865 -56.535 ;
        RECT -261.585 -65.695 -261.305 -56.255 ;
        RECT -262.205 -67.875 -261.805 -66.675 ;
        RECT -263.325 -71.235 -262.925 -70.035 ;
        RECT -265.565 -74.595 -265.165 -73.395 ;
        RECT -270.045 -77.955 -269.645 -76.755 ;
        RECT -279.005 -81.315 -278.605 -80.115 ;
        RECT -296.925 -84.675 -296.525 -83.475 ;
        RECT -261.025 -86.835 -260.745 -56.535 ;
        RECT -260.465 -65.695 -260.185 -56.255 ;
        RECT -259.905 -66.675 -259.625 -56.535 ;
        RECT -259.345 -65.695 -259.065 -56.255 ;
        RECT -259.965 -67.875 -259.565 -66.675 ;
        RECT -258.785 -70.035 -258.505 -56.535 ;
        RECT -258.225 -65.695 -257.945 -56.255 ;
        RECT -257.665 -66.675 -257.385 -56.535 ;
        RECT -257.105 -65.695 -256.825 -56.255 ;
        RECT -257.725 -67.875 -257.325 -66.675 ;
        RECT -258.845 -71.235 -258.445 -70.035 ;
        RECT -256.545 -73.395 -256.265 -56.535 ;
        RECT -255.985 -65.695 -255.705 -56.255 ;
        RECT -255.425 -66.675 -255.145 -56.535 ;
        RECT -254.865 -65.695 -254.585 -56.255 ;
        RECT -255.485 -67.875 -255.085 -66.675 ;
        RECT -254.305 -70.035 -254.025 -56.535 ;
        RECT -253.745 -65.695 -253.465 -56.255 ;
        RECT -253.185 -66.675 -252.905 -56.535 ;
        RECT -252.625 -65.695 -252.345 -56.255 ;
        RECT -253.245 -67.875 -252.845 -66.675 ;
        RECT -254.365 -71.235 -253.965 -70.035 ;
        RECT -256.605 -74.595 -256.205 -73.395 ;
        RECT -252.065 -76.755 -251.785 -56.535 ;
        RECT -251.505 -65.695 -251.225 -56.255 ;
        RECT -250.945 -66.675 -250.665 -56.535 ;
        RECT -250.385 -65.695 -250.105 -56.255 ;
        RECT -251.005 -67.875 -250.605 -66.675 ;
        RECT -249.825 -70.035 -249.545 -56.535 ;
        RECT -249.265 -65.695 -248.985 -56.255 ;
        RECT -248.705 -66.675 -248.425 -56.535 ;
        RECT -248.145 -65.695 -247.865 -56.255 ;
        RECT -248.765 -67.875 -248.365 -66.675 ;
        RECT -249.885 -71.235 -249.485 -70.035 ;
        RECT -247.585 -73.395 -247.305 -56.535 ;
        RECT -247.025 -65.695 -246.745 -56.255 ;
        RECT -246.465 -66.675 -246.185 -56.535 ;
        RECT -245.905 -65.695 -245.625 -56.255 ;
        RECT -246.525 -67.875 -246.125 -66.675 ;
        RECT -245.345 -70.035 -245.065 -56.535 ;
        RECT -244.785 -65.695 -244.505 -56.255 ;
        RECT -244.225 -66.675 -243.945 -56.535 ;
        RECT -243.665 -65.695 -243.385 -56.255 ;
        RECT -244.285 -67.875 -243.885 -66.675 ;
        RECT -245.405 -71.235 -245.005 -70.035 ;
        RECT -247.645 -74.595 -247.245 -73.395 ;
        RECT -252.125 -77.955 -251.725 -76.755 ;
        RECT -243.105 -80.115 -242.825 -56.535 ;
        RECT -242.545 -65.695 -242.265 -56.255 ;
        RECT -241.985 -66.675 -241.705 -56.535 ;
        RECT -241.425 -65.695 -241.145 -56.255 ;
        RECT -242.045 -67.875 -241.645 -66.675 ;
        RECT -240.865 -70.035 -240.585 -56.535 ;
        RECT -240.305 -65.695 -240.025 -56.255 ;
        RECT -239.745 -66.675 -239.465 -56.535 ;
        RECT -239.185 -65.695 -238.905 -56.255 ;
        RECT -239.805 -67.875 -239.405 -66.675 ;
        RECT -240.925 -71.235 -240.525 -70.035 ;
        RECT -238.625 -73.395 -238.345 -56.535 ;
        RECT -238.065 -65.695 -237.785 -56.255 ;
        RECT -237.505 -66.675 -237.225 -56.535 ;
        RECT -236.945 -65.695 -236.665 -56.255 ;
        RECT -237.565 -67.875 -237.165 -66.675 ;
        RECT -236.385 -70.035 -236.105 -56.535 ;
        RECT -235.825 -65.695 -235.545 -56.255 ;
        RECT -235.265 -66.675 -234.985 -56.535 ;
        RECT -234.705 -65.695 -234.425 -56.255 ;
        RECT -235.325 -67.875 -234.925 -66.675 ;
        RECT -236.445 -71.235 -236.045 -70.035 ;
        RECT -238.685 -74.595 -238.285 -73.395 ;
        RECT -234.145 -76.755 -233.865 -56.535 ;
        RECT -233.585 -65.695 -233.305 -56.255 ;
        RECT -233.025 -66.675 -232.745 -56.535 ;
        RECT -232.465 -65.695 -232.185 -56.255 ;
        RECT -233.085 -67.875 -232.685 -66.675 ;
        RECT -231.905 -70.035 -231.625 -56.535 ;
        RECT -231.345 -65.695 -231.065 -56.255 ;
        RECT -230.785 -66.675 -230.505 -56.535 ;
        RECT -230.225 -65.695 -229.945 -56.255 ;
        RECT -230.845 -67.875 -230.445 -66.675 ;
        RECT -231.965 -71.235 -231.565 -70.035 ;
        RECT -229.665 -73.395 -229.385 -56.535 ;
        RECT -229.105 -65.695 -228.825 -56.255 ;
        RECT -228.545 -66.675 -228.265 -56.535 ;
        RECT -227.985 -65.695 -227.705 -56.255 ;
        RECT -228.605 -67.875 -228.205 -66.675 ;
        RECT -227.425 -70.035 -227.145 -56.535 ;
        RECT -226.865 -65.695 -226.585 -56.255 ;
        RECT -226.305 -66.675 -226.025 -56.535 ;
        RECT -225.745 -65.695 -225.465 -56.255 ;
        RECT -226.365 -67.875 -225.965 -66.675 ;
        RECT -227.485 -71.235 -227.085 -70.035 ;
        RECT -229.725 -74.595 -229.325 -73.395 ;
        RECT -234.205 -77.955 -233.805 -76.755 ;
        RECT -243.165 -81.315 -242.765 -80.115 ;
        RECT -225.185 -83.475 -224.905 -56.535 ;
        RECT -224.625 -65.695 -224.345 -56.255 ;
        RECT -224.065 -66.675 -223.785 -56.535 ;
        RECT -223.505 -65.695 -223.225 -56.255 ;
        RECT -224.125 -67.875 -223.725 -66.675 ;
        RECT -222.945 -70.035 -222.665 -56.535 ;
        RECT -222.385 -65.695 -222.105 -56.255 ;
        RECT -221.825 -66.675 -221.545 -56.535 ;
        RECT -221.265 -65.695 -220.985 -56.255 ;
        RECT -221.885 -67.875 -221.485 -66.675 ;
        RECT -223.005 -71.235 -222.605 -70.035 ;
        RECT -220.705 -73.395 -220.425 -56.535 ;
        RECT -220.145 -65.695 -219.865 -56.255 ;
        RECT -219.585 -66.675 -219.305 -56.535 ;
        RECT -219.025 -65.695 -218.745 -56.255 ;
        RECT -219.645 -67.875 -219.245 -66.675 ;
        RECT -218.465 -70.035 -218.185 -56.535 ;
        RECT -217.905 -65.695 -217.625 -56.255 ;
        RECT -217.345 -66.675 -217.065 -56.535 ;
        RECT -216.785 -65.695 -216.505 -56.255 ;
        RECT -217.405 -67.875 -217.005 -66.675 ;
        RECT -218.525 -71.235 -218.125 -70.035 ;
        RECT -220.765 -74.595 -220.365 -73.395 ;
        RECT -216.225 -76.755 -215.945 -56.535 ;
        RECT -215.665 -65.695 -215.385 -56.255 ;
        RECT -215.105 -66.675 -214.825 -56.535 ;
        RECT -214.545 -65.695 -214.265 -56.255 ;
        RECT -215.165 -67.875 -214.765 -66.675 ;
        RECT -213.985 -70.035 -213.705 -56.535 ;
        RECT -213.425 -65.695 -213.145 -56.255 ;
        RECT -212.865 -66.675 -212.585 -56.535 ;
        RECT -212.305 -65.695 -212.025 -56.255 ;
        RECT -212.925 -67.875 -212.525 -66.675 ;
        RECT -214.045 -71.235 -213.645 -70.035 ;
        RECT -211.745 -73.395 -211.465 -56.535 ;
        RECT -211.185 -65.695 -210.905 -56.255 ;
        RECT -210.625 -66.675 -210.345 -56.535 ;
        RECT -210.065 -65.695 -209.785 -56.255 ;
        RECT -210.685 -67.875 -210.285 -66.675 ;
        RECT -209.505 -70.035 -209.225 -56.535 ;
        RECT -208.945 -65.695 -208.665 -56.255 ;
        RECT -208.385 -66.675 -208.105 -56.535 ;
        RECT -207.825 -65.695 -207.545 -56.255 ;
        RECT -208.445 -67.875 -208.045 -66.675 ;
        RECT -209.565 -71.235 -209.165 -70.035 ;
        RECT -211.805 -74.595 -211.405 -73.395 ;
        RECT -216.285 -77.955 -215.885 -76.755 ;
        RECT -207.265 -80.115 -206.985 -56.535 ;
        RECT -206.705 -65.695 -206.425 -56.255 ;
        RECT -206.145 -66.675 -205.865 -56.535 ;
        RECT -205.585 -65.695 -205.305 -56.255 ;
        RECT -206.205 -67.875 -205.805 -66.675 ;
        RECT -205.025 -70.035 -204.745 -56.535 ;
        RECT -204.465 -65.695 -204.185 -56.255 ;
        RECT -203.905 -66.675 -203.625 -56.535 ;
        RECT -203.345 -65.695 -203.065 -56.255 ;
        RECT -203.965 -67.875 -203.565 -66.675 ;
        RECT -205.085 -71.235 -204.685 -70.035 ;
        RECT -202.785 -73.395 -202.505 -56.535 ;
        RECT -202.225 -65.695 -201.945 -56.255 ;
        RECT -201.665 -66.675 -201.385 -56.535 ;
        RECT -201.105 -65.695 -200.825 -56.255 ;
        RECT -201.725 -67.875 -201.325 -66.675 ;
        RECT -200.545 -70.035 -200.265 -56.535 ;
        RECT -199.985 -65.695 -199.705 -56.255 ;
        RECT -199.425 -66.675 -199.145 -56.535 ;
        RECT -198.865 -65.695 -198.585 -56.255 ;
        RECT -199.485 -67.875 -199.085 -66.675 ;
        RECT -200.605 -71.235 -200.205 -70.035 ;
        RECT -202.845 -74.595 -202.445 -73.395 ;
        RECT -198.305 -76.755 -198.025 -56.535 ;
        RECT -197.745 -65.695 -197.465 -56.255 ;
        RECT -197.185 -66.675 -196.905 -56.535 ;
        RECT -196.625 -65.695 -196.345 -56.255 ;
        RECT -197.245 -67.875 -196.845 -66.675 ;
        RECT -196.065 -70.035 -195.785 -56.535 ;
        RECT -195.505 -65.695 -195.225 -56.255 ;
        RECT -194.945 -66.675 -194.665 -56.535 ;
        RECT -194.385 -65.695 -194.105 -56.255 ;
        RECT -195.005 -67.875 -194.605 -66.675 ;
        RECT -196.125 -71.235 -195.725 -70.035 ;
        RECT -193.825 -73.395 -193.545 -56.535 ;
        RECT -193.265 -65.695 -192.985 -56.255 ;
        RECT -192.705 -66.675 -192.425 -56.535 ;
        RECT -192.145 -65.695 -191.865 -56.255 ;
        RECT -192.765 -67.875 -192.365 -66.675 ;
        RECT -191.585 -70.035 -191.305 -56.535 ;
        RECT -191.025 -65.695 -190.745 -56.255 ;
        RECT -190.465 -66.675 -190.185 -56.535 ;
        RECT -189.905 -65.695 -189.625 -56.255 ;
        RECT -190.525 -67.875 -190.125 -66.675 ;
        RECT -191.645 -71.235 -191.245 -70.035 ;
        RECT -193.885 -74.595 -193.485 -73.395 ;
        RECT -198.365 -77.955 -197.965 -76.755 ;
        RECT -207.325 -81.315 -206.925 -80.115 ;
        RECT -225.245 -84.675 -224.845 -83.475 ;
        RECT -261.085 -88.035 -260.685 -86.835 ;
        RECT -490.615 -95.450 -490.235 -90.515 ;
        RECT -332.765 -91.395 -332.365 -90.195 ;
        RECT -493.475 -95.830 -488.545 -95.450 ;
        RECT -189.345 -96.915 -189.065 -56.535 ;
        RECT -188.785 -65.695 -188.505 -56.255 ;
        RECT -188.225 -93.555 -187.945 -56.535 ;
        RECT -187.665 -65.695 -187.385 -56.255 ;
        RECT -187.105 -66.675 -186.825 -56.535 ;
        RECT -186.545 -65.695 -186.265 -56.255 ;
        RECT -187.165 -67.875 -186.765 -66.675 ;
        RECT -185.985 -70.035 -185.705 -56.535 ;
        RECT -185.425 -65.695 -185.145 -56.255 ;
        RECT -184.865 -66.675 -184.585 -56.535 ;
        RECT -184.305 -65.695 -184.025 -56.255 ;
        RECT -184.925 -67.875 -184.525 -66.675 ;
        RECT -186.045 -71.235 -185.645 -70.035 ;
        RECT -183.745 -73.395 -183.465 -56.535 ;
        RECT -183.185 -65.695 -182.905 -56.255 ;
        RECT -182.625 -66.675 -182.345 -56.535 ;
        RECT -182.065 -65.695 -181.785 -56.255 ;
        RECT -182.685 -67.875 -182.285 -66.675 ;
        RECT -181.505 -70.035 -181.225 -56.535 ;
        RECT -180.945 -65.695 -180.665 -56.255 ;
        RECT -180.385 -66.675 -180.105 -56.535 ;
        RECT -179.825 -65.695 -179.545 -56.255 ;
        RECT -180.445 -67.875 -180.045 -66.675 ;
        RECT -181.565 -71.235 -181.165 -70.035 ;
        RECT -183.805 -74.595 -183.405 -73.395 ;
        RECT -179.265 -76.755 -178.985 -56.535 ;
        RECT -178.705 -65.695 -178.425 -56.255 ;
        RECT -178.145 -66.675 -177.865 -56.535 ;
        RECT -177.585 -65.695 -177.305 -56.255 ;
        RECT -178.205 -67.875 -177.805 -66.675 ;
        RECT -177.025 -70.035 -176.745 -56.535 ;
        RECT -176.465 -65.695 -176.185 -56.255 ;
        RECT -175.905 -66.675 -175.625 -56.535 ;
        RECT -175.345 -65.695 -175.065 -56.255 ;
        RECT -175.965 -67.875 -175.565 -66.675 ;
        RECT -177.085 -71.235 -176.685 -70.035 ;
        RECT -174.785 -73.395 -174.505 -56.535 ;
        RECT -174.225 -65.695 -173.945 -56.255 ;
        RECT -173.665 -66.675 -173.385 -56.535 ;
        RECT -173.105 -65.695 -172.825 -56.255 ;
        RECT -173.725 -67.875 -173.325 -66.675 ;
        RECT -172.545 -70.035 -172.265 -56.535 ;
        RECT -171.985 -65.695 -171.705 -56.255 ;
        RECT -171.425 -66.675 -171.145 -56.535 ;
        RECT -170.865 -65.695 -170.585 -56.255 ;
        RECT -171.485 -67.875 -171.085 -66.675 ;
        RECT -172.605 -71.235 -172.205 -70.035 ;
        RECT -174.845 -74.595 -174.445 -73.395 ;
        RECT -179.325 -77.955 -178.925 -76.755 ;
        RECT -170.305 -80.115 -170.025 -56.535 ;
        RECT -169.745 -65.695 -169.465 -56.255 ;
        RECT -169.185 -66.675 -168.905 -56.535 ;
        RECT -168.625 -65.695 -168.345 -56.255 ;
        RECT -169.245 -67.875 -168.845 -66.675 ;
        RECT -168.065 -70.035 -167.785 -56.535 ;
        RECT -167.505 -65.695 -167.225 -56.255 ;
        RECT -166.945 -66.675 -166.665 -56.535 ;
        RECT -166.385 -65.695 -166.105 -56.255 ;
        RECT -167.005 -67.875 -166.605 -66.675 ;
        RECT -168.125 -71.235 -167.725 -70.035 ;
        RECT -165.825 -73.395 -165.545 -56.535 ;
        RECT -165.265 -65.695 -164.985 -56.255 ;
        RECT -164.705 -66.675 -164.425 -56.535 ;
        RECT -164.145 -65.695 -163.865 -56.255 ;
        RECT -164.765 -67.875 -164.365 -66.675 ;
        RECT -163.585 -70.035 -163.305 -56.535 ;
        RECT -163.025 -65.695 -162.745 -56.255 ;
        RECT -162.465 -66.675 -162.185 -56.535 ;
        RECT -161.905 -65.695 -161.625 -56.255 ;
        RECT -162.525 -67.875 -162.125 -66.675 ;
        RECT -163.645 -71.235 -163.245 -70.035 ;
        RECT -165.885 -74.595 -165.485 -73.395 ;
        RECT -161.345 -76.755 -161.065 -56.535 ;
        RECT -160.785 -65.695 -160.505 -56.255 ;
        RECT -160.225 -66.675 -159.945 -56.535 ;
        RECT -159.665 -65.695 -159.385 -56.255 ;
        RECT -160.285 -67.875 -159.885 -66.675 ;
        RECT -159.105 -70.035 -158.825 -56.535 ;
        RECT -158.545 -65.695 -158.265 -56.255 ;
        RECT -157.985 -66.675 -157.705 -56.535 ;
        RECT -157.425 -65.695 -157.145 -56.255 ;
        RECT -158.045 -67.875 -157.645 -66.675 ;
        RECT -159.165 -71.235 -158.765 -70.035 ;
        RECT -156.865 -73.395 -156.585 -56.535 ;
        RECT -156.305 -65.695 -156.025 -56.255 ;
        RECT -155.745 -66.675 -155.465 -56.535 ;
        RECT -155.185 -65.695 -154.905 -56.255 ;
        RECT -155.805 -67.875 -155.405 -66.675 ;
        RECT -154.625 -70.035 -154.345 -56.535 ;
        RECT -154.065 -65.695 -153.785 -56.255 ;
        RECT -153.505 -66.675 -153.225 -56.535 ;
        RECT -152.945 -65.695 -152.665 -56.255 ;
        RECT -153.565 -67.875 -153.165 -66.675 ;
        RECT -154.685 -71.235 -154.285 -70.035 ;
        RECT -156.925 -74.595 -156.525 -73.395 ;
        RECT -161.405 -77.955 -161.005 -76.755 ;
        RECT -170.365 -81.315 -169.965 -80.115 ;
        RECT -152.385 -83.475 -152.105 -56.535 ;
        RECT -151.825 -65.695 -151.545 -56.255 ;
        RECT -151.265 -66.675 -150.985 -56.535 ;
        RECT -150.705 -65.695 -150.425 -56.255 ;
        RECT -151.325 -67.875 -150.925 -66.675 ;
        RECT -150.145 -70.035 -149.865 -56.535 ;
        RECT -149.585 -65.695 -149.305 -56.255 ;
        RECT -149.025 -66.675 -148.745 -56.535 ;
        RECT -148.465 -65.695 -148.185 -56.255 ;
        RECT -149.085 -67.875 -148.685 -66.675 ;
        RECT -150.205 -71.235 -149.805 -70.035 ;
        RECT -147.905 -73.395 -147.625 -56.535 ;
        RECT -147.345 -65.695 -147.065 -56.255 ;
        RECT -146.785 -66.675 -146.505 -56.535 ;
        RECT -146.225 -65.695 -145.945 -56.255 ;
        RECT -146.845 -67.875 -146.445 -66.675 ;
        RECT -145.665 -70.035 -145.385 -56.535 ;
        RECT -145.105 -65.695 -144.825 -56.255 ;
        RECT -144.545 -66.675 -144.265 -56.535 ;
        RECT -143.985 -65.695 -143.705 -56.255 ;
        RECT -144.605 -67.875 -144.205 -66.675 ;
        RECT -145.725 -71.235 -145.325 -70.035 ;
        RECT -147.965 -74.595 -147.565 -73.395 ;
        RECT -143.425 -76.755 -143.145 -56.535 ;
        RECT -142.865 -65.695 -142.585 -56.255 ;
        RECT -142.305 -66.675 -142.025 -56.535 ;
        RECT -141.745 -65.695 -141.465 -56.255 ;
        RECT -142.365 -67.875 -141.965 -66.675 ;
        RECT -141.185 -70.035 -140.905 -56.535 ;
        RECT -140.625 -65.695 -140.345 -56.255 ;
        RECT -140.065 -66.675 -139.785 -56.535 ;
        RECT -139.505 -65.695 -139.225 -56.255 ;
        RECT -140.125 -67.875 -139.725 -66.675 ;
        RECT -141.245 -71.235 -140.845 -70.035 ;
        RECT -138.945 -73.395 -138.665 -56.535 ;
        RECT -138.385 -65.695 -138.105 -56.255 ;
        RECT -137.825 -66.675 -137.545 -56.535 ;
        RECT -137.265 -65.695 -136.985 -56.255 ;
        RECT -137.885 -67.875 -137.485 -66.675 ;
        RECT -136.705 -70.035 -136.425 -56.535 ;
        RECT -136.145 -65.695 -135.865 -56.255 ;
        RECT -135.585 -66.675 -135.305 -56.535 ;
        RECT -135.025 -65.695 -134.745 -56.255 ;
        RECT -135.645 -67.875 -135.245 -66.675 ;
        RECT -136.765 -71.235 -136.365 -70.035 ;
        RECT -139.005 -74.595 -138.605 -73.395 ;
        RECT -143.485 -77.955 -143.085 -76.755 ;
        RECT -134.465 -80.115 -134.185 -56.535 ;
        RECT -133.905 -65.695 -133.625 -56.255 ;
        RECT -133.345 -66.675 -133.065 -56.535 ;
        RECT -132.785 -65.695 -132.505 -56.255 ;
        RECT -133.405 -67.875 -133.005 -66.675 ;
        RECT -132.225 -70.035 -131.945 -56.535 ;
        RECT -131.665 -65.695 -131.385 -56.255 ;
        RECT -131.105 -66.675 -130.825 -56.535 ;
        RECT -130.545 -65.695 -130.265 -56.255 ;
        RECT -131.165 -67.875 -130.765 -66.675 ;
        RECT -132.285 -71.235 -131.885 -70.035 ;
        RECT -129.985 -73.395 -129.705 -56.535 ;
        RECT -129.425 -65.695 -129.145 -56.255 ;
        RECT -128.865 -66.675 -128.585 -56.535 ;
        RECT -128.305 -65.695 -128.025 -56.255 ;
        RECT -128.925 -67.875 -128.525 -66.675 ;
        RECT -127.745 -70.035 -127.465 -56.535 ;
        RECT -127.185 -65.695 -126.905 -56.255 ;
        RECT -126.625 -66.675 -126.345 -56.535 ;
        RECT -126.065 -65.695 -125.785 -56.255 ;
        RECT -126.685 -67.875 -126.285 -66.675 ;
        RECT -127.805 -71.235 -127.405 -70.035 ;
        RECT -130.045 -74.595 -129.645 -73.395 ;
        RECT -125.505 -76.755 -125.225 -56.535 ;
        RECT -124.945 -65.695 -124.665 -56.255 ;
        RECT -124.385 -66.675 -124.105 -56.535 ;
        RECT -123.825 -65.695 -123.545 -56.255 ;
        RECT -124.445 -67.875 -124.045 -66.675 ;
        RECT -123.265 -70.035 -122.985 -56.535 ;
        RECT -122.705 -65.695 -122.425 -56.255 ;
        RECT -122.145 -66.675 -121.865 -56.535 ;
        RECT -121.585 -65.695 -121.305 -56.255 ;
        RECT -122.205 -67.875 -121.805 -66.675 ;
        RECT -123.325 -71.235 -122.925 -70.035 ;
        RECT -121.025 -73.395 -120.745 -56.535 ;
        RECT -120.465 -65.695 -120.185 -56.255 ;
        RECT -119.905 -66.675 -119.625 -56.535 ;
        RECT -119.345 -65.695 -119.065 -56.255 ;
        RECT -119.965 -67.875 -119.565 -66.675 ;
        RECT -118.785 -70.035 -118.505 -56.535 ;
        RECT -118.225 -65.695 -117.945 -56.255 ;
        RECT -117.665 -66.675 -117.385 -56.535 ;
        RECT -117.105 -65.695 -116.825 -56.255 ;
        RECT -117.725 -67.875 -117.325 -66.675 ;
        RECT -118.845 -71.235 -118.445 -70.035 ;
        RECT -121.085 -74.595 -120.685 -73.395 ;
        RECT -125.565 -77.955 -125.165 -76.755 ;
        RECT -134.525 -81.315 -134.125 -80.115 ;
        RECT -152.445 -84.675 -152.045 -83.475 ;
        RECT -116.545 -86.835 -116.265 -56.535 ;
        RECT -115.985 -65.695 -115.705 -56.255 ;
        RECT -115.425 -66.675 -115.145 -56.535 ;
        RECT -114.865 -65.695 -114.585 -56.255 ;
        RECT -115.485 -67.875 -115.085 -66.675 ;
        RECT -114.305 -70.035 -114.025 -56.535 ;
        RECT -113.745 -65.695 -113.465 -56.255 ;
        RECT -113.185 -66.675 -112.905 -56.535 ;
        RECT -112.625 -65.695 -112.345 -56.255 ;
        RECT -113.245 -67.875 -112.845 -66.675 ;
        RECT -114.365 -71.235 -113.965 -70.035 ;
        RECT -112.065 -73.395 -111.785 -56.535 ;
        RECT -111.505 -65.695 -111.225 -56.255 ;
        RECT -110.945 -66.675 -110.665 -56.535 ;
        RECT -110.385 -65.695 -110.105 -56.255 ;
        RECT -111.005 -67.875 -110.605 -66.675 ;
        RECT -109.825 -70.035 -109.545 -56.535 ;
        RECT -109.265 -65.695 -108.985 -56.255 ;
        RECT -108.705 -66.675 -108.425 -56.535 ;
        RECT -108.145 -65.695 -107.865 -56.255 ;
        RECT -108.765 -67.875 -108.365 -66.675 ;
        RECT -109.885 -71.235 -109.485 -70.035 ;
        RECT -112.125 -74.595 -111.725 -73.395 ;
        RECT -107.585 -76.755 -107.305 -56.535 ;
        RECT -107.025 -65.695 -106.745 -56.255 ;
        RECT -106.465 -66.675 -106.185 -56.535 ;
        RECT -105.905 -65.695 -105.625 -56.255 ;
        RECT -106.525 -67.875 -106.125 -66.675 ;
        RECT -105.345 -70.035 -105.065 -56.535 ;
        RECT -104.785 -65.695 -104.505 -56.255 ;
        RECT -104.225 -66.675 -103.945 -56.535 ;
        RECT -103.665 -65.695 -103.385 -56.255 ;
        RECT -104.285 -67.875 -103.885 -66.675 ;
        RECT -105.405 -71.235 -105.005 -70.035 ;
        RECT -103.105 -73.395 -102.825 -56.535 ;
        RECT -102.545 -65.695 -102.265 -56.255 ;
        RECT -101.985 -66.675 -101.705 -56.535 ;
        RECT -101.425 -65.695 -101.145 -56.255 ;
        RECT -102.045 -67.875 -101.645 -66.675 ;
        RECT -100.865 -70.035 -100.585 -56.535 ;
        RECT -100.305 -65.695 -100.025 -56.255 ;
        RECT -99.745 -66.675 -99.465 -56.535 ;
        RECT -99.185 -65.695 -98.905 -56.255 ;
        RECT -99.805 -67.875 -99.405 -66.675 ;
        RECT -100.925 -71.235 -100.525 -70.035 ;
        RECT -103.165 -74.595 -102.765 -73.395 ;
        RECT -107.645 -77.955 -107.245 -76.755 ;
        RECT -98.625 -80.115 -98.345 -56.535 ;
        RECT -98.065 -65.695 -97.785 -56.255 ;
        RECT -97.505 -66.675 -97.225 -56.535 ;
        RECT -96.945 -65.695 -96.665 -56.255 ;
        RECT -97.565 -67.875 -97.165 -66.675 ;
        RECT -96.385 -70.035 -96.105 -56.535 ;
        RECT -95.825 -65.695 -95.545 -56.255 ;
        RECT -95.265 -66.675 -94.985 -56.535 ;
        RECT -94.705 -65.695 -94.425 -56.255 ;
        RECT -95.325 -67.875 -94.925 -66.675 ;
        RECT -96.445 -71.235 -96.045 -70.035 ;
        RECT -94.145 -73.395 -93.865 -56.535 ;
        RECT -93.585 -65.695 -93.305 -56.255 ;
        RECT -93.025 -66.675 -92.745 -56.535 ;
        RECT -92.465 -65.695 -92.185 -56.255 ;
        RECT -93.085 -67.875 -92.685 -66.675 ;
        RECT -91.905 -70.035 -91.625 -56.535 ;
        RECT -91.345 -65.695 -91.065 -56.255 ;
        RECT -90.785 -66.675 -90.505 -56.535 ;
        RECT -90.225 -65.695 -89.945 -56.255 ;
        RECT -90.845 -67.875 -90.445 -66.675 ;
        RECT -91.965 -71.235 -91.565 -70.035 ;
        RECT -94.205 -74.595 -93.805 -73.395 ;
        RECT -89.665 -76.755 -89.385 -56.535 ;
        RECT -89.105 -65.695 -88.825 -56.255 ;
        RECT -88.545 -66.675 -88.265 -56.535 ;
        RECT -87.985 -65.695 -87.705 -56.255 ;
        RECT -88.605 -67.875 -88.205 -66.675 ;
        RECT -87.425 -70.035 -87.145 -56.535 ;
        RECT -86.865 -65.695 -86.585 -56.255 ;
        RECT -86.305 -66.675 -86.025 -56.535 ;
        RECT -85.745 -65.695 -85.465 -56.255 ;
        RECT -86.365 -67.875 -85.965 -66.675 ;
        RECT -87.485 -71.235 -87.085 -70.035 ;
        RECT -85.185 -73.395 -84.905 -56.535 ;
        RECT -84.625 -65.695 -84.345 -56.255 ;
        RECT -84.065 -66.675 -83.785 -56.535 ;
        RECT -83.505 -65.695 -83.225 -56.255 ;
        RECT -84.125 -67.875 -83.725 -66.675 ;
        RECT -82.945 -70.035 -82.665 -56.535 ;
        RECT -82.385 -65.695 -82.105 -56.255 ;
        RECT -81.825 -66.675 -81.545 -56.535 ;
        RECT -81.265 -65.695 -80.985 -56.255 ;
        RECT -81.885 -67.875 -81.485 -66.675 ;
        RECT -83.005 -71.235 -82.605 -70.035 ;
        RECT -85.245 -74.595 -84.845 -73.395 ;
        RECT -89.725 -77.955 -89.325 -76.755 ;
        RECT -98.685 -81.315 -98.285 -80.115 ;
        RECT -80.705 -83.475 -80.425 -56.535 ;
        RECT -80.145 -65.695 -79.865 -56.255 ;
        RECT -79.585 -66.675 -79.305 -56.535 ;
        RECT -79.025 -65.695 -78.745 -56.255 ;
        RECT -79.645 -67.875 -79.245 -66.675 ;
        RECT -78.465 -70.035 -78.185 -56.535 ;
        RECT -77.905 -65.695 -77.625 -56.255 ;
        RECT -77.345 -66.675 -77.065 -56.535 ;
        RECT -76.785 -65.695 -76.505 -56.255 ;
        RECT -77.405 -67.875 -77.005 -66.675 ;
        RECT -78.525 -71.235 -78.125 -70.035 ;
        RECT -76.225 -73.395 -75.945 -56.535 ;
        RECT -75.665 -65.695 -75.385 -56.255 ;
        RECT -75.105 -66.675 -74.825 -56.535 ;
        RECT -74.545 -65.695 -74.265 -56.255 ;
        RECT -75.165 -67.875 -74.765 -66.675 ;
        RECT -73.985 -70.035 -73.705 -56.535 ;
        RECT -73.425 -65.695 -73.145 -56.255 ;
        RECT -72.865 -66.675 -72.585 -56.535 ;
        RECT -72.305 -65.695 -72.025 -56.255 ;
        RECT -72.925 -67.875 -72.525 -66.675 ;
        RECT -74.045 -71.235 -73.645 -70.035 ;
        RECT -76.285 -74.595 -75.885 -73.395 ;
        RECT -71.745 -76.755 -71.465 -56.535 ;
        RECT -71.185 -65.695 -70.905 -56.255 ;
        RECT -70.625 -66.675 -70.345 -56.535 ;
        RECT -70.065 -65.695 -69.785 -56.255 ;
        RECT -70.685 -67.875 -70.285 -66.675 ;
        RECT -69.505 -70.035 -69.225 -56.535 ;
        RECT -68.945 -65.695 -68.665 -56.255 ;
        RECT -68.385 -66.675 -68.105 -56.535 ;
        RECT -67.825 -65.695 -67.545 -56.255 ;
        RECT -68.445 -67.875 -68.045 -66.675 ;
        RECT -69.565 -71.235 -69.165 -70.035 ;
        RECT -67.265 -73.395 -66.985 -56.535 ;
        RECT -66.705 -65.695 -66.425 -56.255 ;
        RECT -66.145 -66.675 -65.865 -56.535 ;
        RECT -65.585 -65.695 -65.305 -56.255 ;
        RECT -66.205 -67.875 -65.805 -66.675 ;
        RECT -65.025 -70.035 -64.745 -56.535 ;
        RECT -64.465 -65.695 -64.185 -56.255 ;
        RECT -63.905 -66.675 -63.625 -56.535 ;
        RECT -63.345 -65.695 -63.065 -56.255 ;
        RECT -63.965 -67.875 -63.565 -66.675 ;
        RECT -65.085 -71.235 -64.685 -70.035 ;
        RECT -67.325 -74.595 -66.925 -73.395 ;
        RECT -71.805 -77.955 -71.405 -76.755 ;
        RECT -62.785 -80.115 -62.505 -56.535 ;
        RECT -62.225 -65.695 -61.945 -56.255 ;
        RECT -61.665 -66.675 -61.385 -56.535 ;
        RECT -61.105 -65.695 -60.825 -56.255 ;
        RECT -61.725 -67.875 -61.325 -66.675 ;
        RECT -60.545 -70.035 -60.265 -56.535 ;
        RECT -59.985 -65.695 -59.705 -56.255 ;
        RECT -59.425 -66.675 -59.145 -56.535 ;
        RECT -58.865 -65.695 -58.585 -56.255 ;
        RECT -59.485 -67.875 -59.085 -66.675 ;
        RECT -60.605 -71.235 -60.205 -70.035 ;
        RECT -58.305 -73.395 -58.025 -56.535 ;
        RECT -57.745 -65.695 -57.465 -56.255 ;
        RECT -57.185 -66.675 -56.905 -56.535 ;
        RECT -56.625 -65.695 -56.345 -56.255 ;
        RECT -57.245 -67.875 -56.845 -66.675 ;
        RECT -56.065 -70.035 -55.785 -56.535 ;
        RECT -55.505 -65.695 -55.225 -56.255 ;
        RECT -54.945 -66.675 -54.665 -56.535 ;
        RECT -54.385 -65.695 -54.105 -56.255 ;
        RECT -55.005 -67.875 -54.605 -66.675 ;
        RECT -56.125 -71.235 -55.725 -70.035 ;
        RECT -58.365 -74.595 -57.965 -73.395 ;
        RECT -53.825 -76.755 -53.545 -56.535 ;
        RECT -53.265 -65.695 -52.985 -56.255 ;
        RECT -52.705 -66.675 -52.425 -56.535 ;
        RECT -52.145 -65.695 -51.865 -56.255 ;
        RECT -52.765 -67.875 -52.365 -66.675 ;
        RECT -51.585 -70.035 -51.305 -56.535 ;
        RECT -51.025 -65.695 -50.745 -56.255 ;
        RECT -50.465 -66.675 -50.185 -56.535 ;
        RECT -49.905 -65.695 -49.625 -56.255 ;
        RECT -50.525 -67.875 -50.125 -66.675 ;
        RECT -51.645 -71.235 -51.245 -70.035 ;
        RECT -49.345 -73.395 -49.065 -56.535 ;
        RECT -48.785 -65.695 -48.505 -56.255 ;
        RECT -48.225 -66.675 -47.945 -56.535 ;
        RECT -47.665 -65.695 -47.385 -56.255 ;
        RECT -48.285 -67.875 -47.885 -66.675 ;
        RECT -47.105 -70.035 -46.825 -56.535 ;
        RECT -46.545 -65.695 -46.265 -56.255 ;
        RECT -45.985 -66.675 -45.705 -56.535 ;
        RECT -45.425 -65.695 -45.145 -56.255 ;
        RECT -46.045 -67.875 -45.645 -66.675 ;
        RECT -47.165 -71.235 -46.765 -70.035 ;
        RECT -49.405 -74.595 -49.005 -73.395 ;
        RECT -53.885 -77.955 -53.485 -76.755 ;
        RECT -62.845 -81.315 -62.445 -80.115 ;
        RECT -80.765 -84.675 -80.365 -83.475 ;
        RECT -116.605 -88.035 -116.205 -86.835 ;
        RECT -44.865 -90.195 -44.585 -56.535 ;
        RECT -44.305 -65.695 -44.025 -56.255 ;
        RECT -43.745 -66.675 -43.465 -56.535 ;
        RECT -43.185 -65.695 -42.905 -56.255 ;
        RECT -43.805 -67.875 -43.405 -66.675 ;
        RECT -42.625 -70.035 -42.345 -56.535 ;
        RECT -42.065 -65.695 -41.785 -56.255 ;
        RECT -41.505 -66.675 -41.225 -56.535 ;
        RECT -40.945 -65.695 -40.665 -56.255 ;
        RECT -41.565 -67.875 -41.165 -66.675 ;
        RECT -42.685 -71.235 -42.285 -70.035 ;
        RECT -40.385 -73.395 -40.105 -56.535 ;
        RECT -39.825 -65.695 -39.545 -56.255 ;
        RECT -39.265 -66.675 -38.985 -56.535 ;
        RECT -38.705 -65.695 -38.425 -56.255 ;
        RECT -39.325 -67.875 -38.925 -66.675 ;
        RECT -38.145 -70.035 -37.865 -56.535 ;
        RECT -37.585 -65.695 -37.305 -56.255 ;
        RECT -37.025 -66.675 -36.745 -56.535 ;
        RECT -36.465 -65.695 -36.185 -56.255 ;
        RECT -37.085 -67.875 -36.685 -66.675 ;
        RECT -38.205 -71.235 -37.805 -70.035 ;
        RECT -40.445 -74.595 -40.045 -73.395 ;
        RECT -35.905 -76.755 -35.625 -56.535 ;
        RECT -35.345 -65.695 -35.065 -56.255 ;
        RECT -34.785 -66.675 -34.505 -56.535 ;
        RECT -34.225 -65.695 -33.945 -56.255 ;
        RECT -34.845 -67.875 -34.445 -66.675 ;
        RECT -33.665 -70.035 -33.385 -56.535 ;
        RECT -33.105 -65.695 -32.825 -56.255 ;
        RECT -32.545 -66.675 -32.265 -56.535 ;
        RECT -31.985 -65.695 -31.705 -56.255 ;
        RECT -32.605 -67.875 -32.205 -66.675 ;
        RECT -33.725 -71.235 -33.325 -70.035 ;
        RECT -31.425 -73.395 -31.145 -56.535 ;
        RECT -30.865 -65.695 -30.585 -56.255 ;
        RECT -30.305 -66.675 -30.025 -56.535 ;
        RECT -29.745 -65.695 -29.465 -56.255 ;
        RECT -30.365 -67.875 -29.965 -66.675 ;
        RECT -29.185 -70.035 -28.905 -56.535 ;
        RECT -28.625 -65.695 -28.345 -56.255 ;
        RECT -28.065 -66.675 -27.785 -56.535 ;
        RECT -27.505 -65.695 -27.225 -56.255 ;
        RECT -28.125 -67.875 -27.725 -66.675 ;
        RECT -29.245 -71.235 -28.845 -70.035 ;
        RECT -31.485 -74.595 -31.085 -73.395 ;
        RECT -35.965 -77.955 -35.565 -76.755 ;
        RECT -26.945 -80.115 -26.665 -56.535 ;
        RECT -26.385 -65.695 -26.105 -56.255 ;
        RECT -25.825 -66.675 -25.545 -56.535 ;
        RECT -25.265 -65.695 -24.985 -56.255 ;
        RECT -25.885 -67.875 -25.485 -66.675 ;
        RECT -24.705 -70.035 -24.425 -56.535 ;
        RECT -24.145 -65.695 -23.865 -56.255 ;
        RECT -23.585 -66.675 -23.305 -56.535 ;
        RECT -23.025 -65.695 -22.745 -56.255 ;
        RECT -23.645 -67.875 -23.245 -66.675 ;
        RECT -24.765 -71.235 -24.365 -70.035 ;
        RECT -22.465 -73.395 -22.185 -56.535 ;
        RECT -21.905 -65.695 -21.625 -56.255 ;
        RECT -21.345 -66.675 -21.065 -56.535 ;
        RECT -20.785 -65.695 -20.505 -56.255 ;
        RECT -21.405 -67.875 -21.005 -66.675 ;
        RECT -20.225 -70.035 -19.945 -56.535 ;
        RECT -19.665 -65.695 -19.385 -56.255 ;
        RECT -19.105 -66.675 -18.825 -56.535 ;
        RECT -18.545 -65.695 -18.265 -56.255 ;
        RECT -19.165 -67.875 -18.765 -66.675 ;
        RECT -20.285 -71.235 -19.885 -70.035 ;
        RECT -22.525 -74.595 -22.125 -73.395 ;
        RECT -17.985 -76.755 -17.705 -56.535 ;
        RECT -17.425 -65.695 -17.145 -56.255 ;
        RECT -16.865 -66.675 -16.585 -56.535 ;
        RECT -16.305 -65.695 -16.025 -56.255 ;
        RECT -16.925 -67.875 -16.525 -66.675 ;
        RECT -15.745 -70.035 -15.465 -56.535 ;
        RECT -15.185 -65.695 -14.905 -56.255 ;
        RECT -14.625 -66.675 -14.345 -56.535 ;
        RECT -14.065 -65.695 -13.785 -56.255 ;
        RECT -14.685 -67.875 -14.285 -66.675 ;
        RECT -15.805 -71.235 -15.405 -70.035 ;
        RECT -13.505 -73.395 -13.225 -56.535 ;
        RECT -12.945 -65.695 -12.665 -56.255 ;
        RECT -12.385 -66.675 -12.105 -56.535 ;
        RECT -11.825 -65.695 -11.545 -56.255 ;
        RECT -12.445 -67.875 -12.045 -66.675 ;
        RECT -11.265 -70.035 -10.985 -56.535 ;
        RECT -10.705 -65.695 -10.425 -56.255 ;
        RECT -10.145 -66.675 -9.865 -56.535 ;
        RECT -9.585 -65.695 -9.305 -56.255 ;
        RECT -10.205 -67.875 -9.805 -66.675 ;
        RECT -11.325 -71.235 -10.925 -70.035 ;
        RECT -13.565 -74.595 -13.165 -73.395 ;
        RECT -18.045 -77.955 -17.645 -76.755 ;
        RECT -27.005 -81.315 -26.605 -80.115 ;
        RECT -9.025 -83.475 -8.745 -56.535 ;
        RECT -8.465 -65.695 -8.185 -56.255 ;
        RECT -7.905 -66.675 -7.625 -56.535 ;
        RECT -7.345 -65.695 -7.065 -56.255 ;
        RECT -7.965 -67.875 -7.565 -66.675 ;
        RECT -6.785 -70.035 -6.505 -56.535 ;
        RECT -6.225 -65.695 -5.945 -56.255 ;
        RECT -5.665 -66.675 -5.385 -56.535 ;
        RECT -5.105 -65.695 -4.825 -56.255 ;
        RECT -5.725 -67.875 -5.325 -66.675 ;
        RECT -6.845 -71.235 -6.445 -70.035 ;
        RECT -4.545 -73.395 -4.265 -56.535 ;
        RECT -3.985 -65.695 -3.705 -56.255 ;
        RECT -3.425 -66.675 -3.145 -56.535 ;
        RECT -2.865 -65.695 -2.585 -56.255 ;
        RECT -3.485 -67.875 -3.085 -66.675 ;
        RECT -2.305 -70.035 -2.025 -56.535 ;
        RECT -1.745 -65.695 -1.465 -56.255 ;
        RECT -1.185 -66.675 -0.905 -56.535 ;
        RECT -0.625 -65.695 -0.345 -56.255 ;
        RECT -1.245 -67.875 -0.845 -66.675 ;
        RECT -2.365 -71.235 -1.965 -70.035 ;
        RECT -4.605 -74.595 -4.205 -73.395 ;
        RECT -0.065 -76.755 0.215 -56.535 ;
        RECT 0.495 -65.695 0.775 -56.255 ;
        RECT 1.055 -66.675 1.335 -56.535 ;
        RECT 1.615 -65.695 1.895 -56.255 ;
        RECT 0.995 -67.875 1.395 -66.675 ;
        RECT 2.175 -70.035 2.455 -56.535 ;
        RECT 2.735 -65.695 3.015 -56.255 ;
        RECT 3.295 -66.675 3.575 -56.535 ;
        RECT 3.855 -65.695 4.135 -56.255 ;
        RECT 3.235 -67.875 3.635 -66.675 ;
        RECT 2.115 -71.235 2.515 -70.035 ;
        RECT 4.415 -73.395 4.695 -56.535 ;
        RECT 4.975 -65.695 5.255 -56.255 ;
        RECT 5.535 -66.675 5.815 -56.535 ;
        RECT 6.095 -65.695 6.375 -56.255 ;
        RECT 5.475 -67.875 5.875 -66.675 ;
        RECT 6.655 -70.035 6.935 -56.535 ;
        RECT 7.215 -65.695 7.495 -56.255 ;
        RECT 7.775 -66.675 8.055 -56.535 ;
        RECT 8.335 -65.695 8.615 -56.255 ;
        RECT 7.715 -67.875 8.115 -66.675 ;
        RECT 6.595 -71.235 6.995 -70.035 ;
        RECT 4.355 -74.595 4.755 -73.395 ;
        RECT -0.125 -77.955 0.275 -76.755 ;
        RECT 8.895 -80.115 9.175 -56.535 ;
        RECT 9.455 -65.695 9.735 -56.255 ;
        RECT 10.015 -66.675 10.295 -56.535 ;
        RECT 10.575 -65.695 10.855 -56.255 ;
        RECT 9.955 -67.875 10.355 -66.675 ;
        RECT 11.135 -70.035 11.415 -56.535 ;
        RECT 11.695 -65.695 11.975 -56.255 ;
        RECT 12.255 -66.675 12.535 -56.535 ;
        RECT 12.815 -65.695 13.095 -56.255 ;
        RECT 12.195 -67.875 12.595 -66.675 ;
        RECT 11.075 -71.235 11.475 -70.035 ;
        RECT 13.375 -73.395 13.655 -56.535 ;
        RECT 13.935 -65.695 14.215 -56.255 ;
        RECT 14.495 -66.675 14.775 -56.535 ;
        RECT 15.055 -65.695 15.335 -56.255 ;
        RECT 14.435 -67.875 14.835 -66.675 ;
        RECT 15.615 -70.035 15.895 -56.535 ;
        RECT 16.175 -65.695 16.455 -56.255 ;
        RECT 16.735 -66.675 17.015 -56.535 ;
        RECT 17.295 -65.695 17.575 -56.255 ;
        RECT 16.675 -67.875 17.075 -66.675 ;
        RECT 15.555 -71.235 15.955 -70.035 ;
        RECT 13.315 -74.595 13.715 -73.395 ;
        RECT 17.855 -76.755 18.135 -56.535 ;
        RECT 18.415 -65.695 18.695 -56.255 ;
        RECT 18.975 -66.675 19.255 -56.535 ;
        RECT 19.535 -65.695 19.815 -56.255 ;
        RECT 18.915 -67.875 19.315 -66.675 ;
        RECT 20.095 -70.035 20.375 -56.535 ;
        RECT 20.655 -65.695 20.935 -56.255 ;
        RECT 21.215 -66.675 21.495 -56.535 ;
        RECT 21.775 -65.695 22.055 -56.255 ;
        RECT 21.155 -67.875 21.555 -66.675 ;
        RECT 20.035 -71.235 20.435 -70.035 ;
        RECT 22.335 -73.395 22.615 -56.535 ;
        RECT 22.895 -65.695 23.175 -56.255 ;
        RECT 23.455 -66.675 23.735 -56.535 ;
        RECT 24.015 -65.695 24.295 -56.255 ;
        RECT 23.395 -67.875 23.795 -66.675 ;
        RECT 24.575 -70.035 24.855 -56.535 ;
        RECT 25.135 -65.695 25.415 -56.255 ;
        RECT 25.695 -66.675 25.975 -56.535 ;
        RECT 26.255 -65.695 26.535 -56.255 ;
        RECT 25.635 -67.875 26.035 -66.675 ;
        RECT 24.515 -71.235 24.915 -70.035 ;
        RECT 22.275 -74.595 22.675 -73.395 ;
        RECT 17.795 -77.955 18.195 -76.755 ;
        RECT 8.835 -81.315 9.235 -80.115 ;
        RECT -9.085 -84.675 -8.685 -83.475 ;
        RECT 26.815 -86.835 27.095 -56.535 ;
        RECT 27.375 -65.695 27.655 -56.255 ;
        RECT 27.935 -66.675 28.215 -56.535 ;
        RECT 28.495 -65.695 28.775 -56.255 ;
        RECT 27.875 -67.875 28.275 -66.675 ;
        RECT 29.055 -70.035 29.335 -56.535 ;
        RECT 29.615 -65.695 29.895 -56.255 ;
        RECT 30.175 -66.675 30.455 -56.535 ;
        RECT 30.735 -65.695 31.015 -56.255 ;
        RECT 30.115 -67.875 30.515 -66.675 ;
        RECT 28.995 -71.235 29.395 -70.035 ;
        RECT 31.295 -73.395 31.575 -56.535 ;
        RECT 31.855 -65.695 32.135 -56.255 ;
        RECT 32.415 -66.675 32.695 -56.535 ;
        RECT 32.975 -65.695 33.255 -56.255 ;
        RECT 32.355 -67.875 32.755 -66.675 ;
        RECT 33.535 -70.035 33.815 -56.535 ;
        RECT 34.095 -65.695 34.375 -56.255 ;
        RECT 34.655 -66.675 34.935 -56.535 ;
        RECT 35.215 -65.695 35.495 -56.255 ;
        RECT 34.595 -67.875 34.995 -66.675 ;
        RECT 33.475 -71.235 33.875 -70.035 ;
        RECT 31.235 -74.595 31.635 -73.395 ;
        RECT 35.775 -76.755 36.055 -56.535 ;
        RECT 36.335 -65.695 36.615 -56.255 ;
        RECT 36.895 -66.675 37.175 -56.535 ;
        RECT 37.455 -65.695 37.735 -56.255 ;
        RECT 36.835 -67.875 37.235 -66.675 ;
        RECT 38.015 -70.035 38.295 -56.535 ;
        RECT 38.575 -65.695 38.855 -56.255 ;
        RECT 39.135 -66.675 39.415 -56.535 ;
        RECT 39.695 -65.695 39.975 -56.255 ;
        RECT 39.075 -67.875 39.475 -66.675 ;
        RECT 37.955 -71.235 38.355 -70.035 ;
        RECT 40.255 -73.395 40.535 -56.535 ;
        RECT 40.815 -65.695 41.095 -56.255 ;
        RECT 41.375 -66.675 41.655 -56.535 ;
        RECT 41.935 -65.695 42.215 -56.255 ;
        RECT 41.315 -67.875 41.715 -66.675 ;
        RECT 42.495 -70.035 42.775 -56.535 ;
        RECT 43.055 -65.695 43.335 -56.255 ;
        RECT 43.615 -66.675 43.895 -56.535 ;
        RECT 44.175 -65.695 44.455 -56.255 ;
        RECT 43.555 -67.875 43.955 -66.675 ;
        RECT 42.435 -71.235 42.835 -70.035 ;
        RECT 40.195 -74.595 40.595 -73.395 ;
        RECT 35.715 -77.955 36.115 -76.755 ;
        RECT 44.735 -80.115 45.015 -56.535 ;
        RECT 45.295 -65.695 45.575 -56.255 ;
        RECT 45.855 -66.675 46.135 -56.535 ;
        RECT 46.415 -65.695 46.695 -56.255 ;
        RECT 45.795 -67.875 46.195 -66.675 ;
        RECT 46.975 -70.035 47.255 -56.535 ;
        RECT 47.535 -65.695 47.815 -56.255 ;
        RECT 48.095 -66.675 48.375 -56.535 ;
        RECT 48.655 -65.695 48.935 -56.255 ;
        RECT 48.035 -67.875 48.435 -66.675 ;
        RECT 46.915 -71.235 47.315 -70.035 ;
        RECT 49.215 -73.395 49.495 -56.535 ;
        RECT 49.775 -65.695 50.055 -56.255 ;
        RECT 50.335 -66.675 50.615 -56.535 ;
        RECT 50.895 -65.695 51.175 -56.255 ;
        RECT 50.275 -67.875 50.675 -66.675 ;
        RECT 51.455 -70.035 51.735 -56.535 ;
        RECT 52.015 -65.695 52.295 -56.255 ;
        RECT 52.575 -66.675 52.855 -56.535 ;
        RECT 53.135 -65.695 53.415 -56.255 ;
        RECT 52.515 -67.875 52.915 -66.675 ;
        RECT 51.395 -71.235 51.795 -70.035 ;
        RECT 49.155 -74.595 49.555 -73.395 ;
        RECT 53.695 -76.755 53.975 -56.535 ;
        RECT 54.255 -65.695 54.535 -56.255 ;
        RECT 54.815 -66.675 55.095 -56.535 ;
        RECT 55.375 -65.695 55.655 -56.255 ;
        RECT 54.755 -67.875 55.155 -66.675 ;
        RECT 55.935 -70.035 56.215 -56.535 ;
        RECT 56.495 -65.695 56.775 -56.255 ;
        RECT 57.055 -66.675 57.335 -56.535 ;
        RECT 57.615 -65.695 57.895 -56.255 ;
        RECT 56.995 -67.875 57.395 -66.675 ;
        RECT 55.875 -71.235 56.275 -70.035 ;
        RECT 58.175 -73.395 58.455 -56.535 ;
        RECT 58.735 -65.695 59.015 -56.255 ;
        RECT 59.295 -66.675 59.575 -56.535 ;
        RECT 59.855 -65.695 60.135 -56.255 ;
        RECT 59.235 -67.875 59.635 -66.675 ;
        RECT 60.415 -70.035 60.695 -56.535 ;
        RECT 60.975 -65.695 61.255 -56.255 ;
        RECT 61.535 -66.675 61.815 -56.535 ;
        RECT 62.095 -65.695 62.375 -56.255 ;
        RECT 61.475 -67.875 61.875 -66.675 ;
        RECT 60.355 -71.235 60.755 -70.035 ;
        RECT 58.115 -74.595 58.515 -73.395 ;
        RECT 53.635 -77.955 54.035 -76.755 ;
        RECT 44.675 -81.315 45.075 -80.115 ;
        RECT 62.655 -83.475 62.935 -56.535 ;
        RECT 63.215 -65.695 63.495 -56.255 ;
        RECT 63.775 -66.675 64.055 -56.535 ;
        RECT 64.335 -65.695 64.615 -56.255 ;
        RECT 63.715 -67.875 64.115 -66.675 ;
        RECT 64.895 -70.035 65.175 -56.535 ;
        RECT 65.455 -65.695 65.735 -56.255 ;
        RECT 66.015 -66.675 66.295 -56.535 ;
        RECT 66.575 -65.695 66.855 -56.255 ;
        RECT 65.955 -67.875 66.355 -66.675 ;
        RECT 64.835 -71.235 65.235 -70.035 ;
        RECT 67.135 -73.395 67.415 -56.535 ;
        RECT 67.695 -65.695 67.975 -56.255 ;
        RECT 68.255 -66.675 68.535 -56.535 ;
        RECT 68.815 -65.695 69.095 -56.255 ;
        RECT 68.195 -67.875 68.595 -66.675 ;
        RECT 69.375 -70.035 69.655 -56.535 ;
        RECT 69.935 -65.695 70.215 -56.255 ;
        RECT 70.495 -66.675 70.775 -56.535 ;
        RECT 71.055 -65.695 71.335 -56.255 ;
        RECT 70.435 -67.875 70.835 -66.675 ;
        RECT 69.315 -71.235 69.715 -70.035 ;
        RECT 67.075 -74.595 67.475 -73.395 ;
        RECT 71.615 -76.755 71.895 -56.535 ;
        RECT 72.175 -65.695 72.455 -56.255 ;
        RECT 72.735 -66.675 73.015 -56.535 ;
        RECT 73.295 -65.695 73.575 -56.255 ;
        RECT 72.675 -67.875 73.075 -66.675 ;
        RECT 73.855 -70.035 74.135 -56.535 ;
        RECT 74.415 -65.695 74.695 -56.255 ;
        RECT 74.975 -66.675 75.255 -56.535 ;
        RECT 75.535 -65.695 75.815 -56.255 ;
        RECT 74.915 -67.875 75.315 -66.675 ;
        RECT 73.795 -71.235 74.195 -70.035 ;
        RECT 76.095 -73.395 76.375 -56.535 ;
        RECT 76.655 -65.695 76.935 -56.255 ;
        RECT 77.215 -66.675 77.495 -56.535 ;
        RECT 77.775 -65.695 78.055 -56.255 ;
        RECT 77.155 -67.875 77.555 -66.675 ;
        RECT 78.335 -70.035 78.615 -56.535 ;
        RECT 78.895 -65.695 79.175 -56.255 ;
        RECT 79.455 -66.675 79.735 -56.535 ;
        RECT 80.015 -65.695 80.295 -56.255 ;
        RECT 79.395 -67.875 79.795 -66.675 ;
        RECT 78.275 -71.235 78.675 -70.035 ;
        RECT 76.035 -74.595 76.435 -73.395 ;
        RECT 71.555 -77.955 71.955 -76.755 ;
        RECT 80.575 -80.115 80.855 -56.535 ;
        RECT 81.135 -65.695 81.415 -56.255 ;
        RECT 81.695 -66.675 81.975 -56.535 ;
        RECT 82.255 -65.695 82.535 -56.255 ;
        RECT 81.635 -67.875 82.035 -66.675 ;
        RECT 82.815 -70.035 83.095 -56.535 ;
        RECT 83.375 -65.695 83.655 -56.255 ;
        RECT 83.935 -66.675 84.215 -56.535 ;
        RECT 84.495 -65.695 84.775 -56.255 ;
        RECT 83.875 -67.875 84.275 -66.675 ;
        RECT 82.755 -71.235 83.155 -70.035 ;
        RECT 85.055 -73.395 85.335 -56.535 ;
        RECT 85.615 -65.695 85.895 -56.255 ;
        RECT 86.175 -66.675 86.455 -56.535 ;
        RECT 86.735 -65.695 87.015 -56.255 ;
        RECT 86.115 -67.875 86.515 -66.675 ;
        RECT 87.295 -70.035 87.575 -56.535 ;
        RECT 87.855 -65.695 88.135 -56.255 ;
        RECT 88.415 -66.675 88.695 -56.535 ;
        RECT 88.975 -65.695 89.255 -56.255 ;
        RECT 88.355 -67.875 88.755 -66.675 ;
        RECT 87.235 -71.235 87.635 -70.035 ;
        RECT 84.995 -74.595 85.395 -73.395 ;
        RECT 89.535 -76.755 89.815 -56.535 ;
        RECT 90.095 -65.695 90.375 -56.255 ;
        RECT 90.655 -66.675 90.935 -56.535 ;
        RECT 91.215 -65.695 91.495 -56.255 ;
        RECT 90.595 -67.875 90.995 -66.675 ;
        RECT 91.775 -70.035 92.055 -56.535 ;
        RECT 92.335 -65.695 92.615 -56.255 ;
        RECT 92.895 -66.675 93.175 -56.535 ;
        RECT 93.455 -65.695 93.735 -56.255 ;
        RECT 92.835 -67.875 93.235 -66.675 ;
        RECT 91.715 -71.235 92.115 -70.035 ;
        RECT 94.015 -73.395 94.295 -56.535 ;
        RECT 94.575 -65.695 94.855 -56.255 ;
        RECT 95.135 -66.675 95.415 -56.535 ;
        RECT 95.695 -65.695 95.975 -56.255 ;
        RECT 95.075 -67.875 95.475 -66.675 ;
        RECT 96.255 -70.035 96.535 -56.535 ;
        RECT 96.815 -65.695 97.095 -56.255 ;
        RECT 97.375 -66.675 97.655 -56.535 ;
        RECT 97.935 -65.695 98.215 -56.255 ;
        RECT 98.495 -66.285 98.775 -56.695 ;
        RECT 99.055 -65.695 99.335 -56.255 ;
        RECT 99.615 -66.285 99.895 -56.695 ;
        RECT 100.175 -66.285 100.455 -56.255 ;
        RECT 274.700 -56.260 289.200 -55.260 ;
        RECT 298.300 -61.000 298.580 -48.340 ;
        RECT 306.140 -55.950 306.420 -40.780 ;
        RECT 308.940 -43.630 309.220 -20.290 ;
        RECT 309.500 -31.870 309.780 -16.370 ;
        RECT 310.060 -39.150 310.340 3.460 ;
        RECT 312.300 2.850 312.580 3.790 ;
        RECT 311.740 -4.570 312.020 -4.050 ;
        RECT 312.300 -24.590 312.580 -23.650 ;
        RECT 312.860 -29.070 313.140 -15.250 ;
        RECT 313.420 -20.670 313.700 35.660 ;
        RECT 314.540 35.660 315.380 35.940 ;
        RECT 313.980 18.950 314.260 19.470 ;
        RECT 313.980 5.090 314.260 11.630 ;
        RECT 313.980 -25.290 314.260 -24.770 ;
        RECT 313.420 -30.750 313.700 -26.450 ;
        RECT 314.540 -28.740 314.820 35.660 ;
        RECT 317.340 31.180 317.620 31.230 ;
        RECT 318.460 31.180 318.740 39.070 ;
        RECT 317.340 30.900 318.740 31.180 ;
        RECT 317.340 26.140 317.620 30.900 ;
        RECT 317.900 26.790 318.180 27.310 ;
        RECT 319.020 27.260 319.300 46.910 ;
        RECT 346.460 46.860 346.740 46.910 ;
        RECT 354.860 46.860 355.140 46.910 ;
        RECT 344.220 46.580 346.740 46.860 ;
        RECT 334.140 43.170 334.420 44.110 ;
        RECT 340.860 44.060 341.140 44.110 ;
        RECT 342.540 44.060 342.820 44.110 ;
        RECT 340.860 43.780 342.820 44.060 ;
        RECT 340.860 43.730 341.140 43.780 ;
        RECT 342.540 43.730 342.820 43.780 ;
        RECT 344.220 43.590 344.500 46.580 ;
        RECT 346.460 46.530 346.740 46.580 ;
        RECT 352.060 46.580 355.140 46.860 ;
        RECT 352.060 44.060 352.340 46.580 ;
        RECT 354.860 46.530 355.140 46.580 ;
        RECT 384.540 45.740 384.820 46.910 ;
        RECT 389.020 45.740 389.300 45.790 ;
        RECT 384.540 45.460 389.300 45.740 ;
        RECT 349.820 43.780 352.340 44.060 ;
        RECT 349.820 43.170 350.100 43.780 ;
        RECT 352.060 43.730 352.340 43.780 ;
        RECT 353.740 43.590 354.020 44.110 ;
        RECT 376.140 43.590 376.420 44.110 ;
        RECT 384.540 44.060 384.820 45.460 ;
        RECT 389.020 45.410 389.300 45.460 ;
        RECT 405.820 45.410 406.100 46.910 ;
        RECT 408.060 45.270 408.340 45.790 ;
        RECT 383.420 43.780 384.820 44.060 ;
        RECT 392.380 44.060 392.660 44.110 ;
        RECT 392.380 43.780 397.140 44.060 ;
        RECT 319.580 41.910 319.860 42.430 ;
        RECT 338.060 42.380 338.340 42.430 ;
        RECT 338.060 42.100 338.900 42.380 ;
        RECT 338.060 42.050 338.340 42.100 ;
        RECT 321.820 35.330 322.100 39.070 ;
        RECT 320.140 31.180 320.420 31.230 ;
        RECT 320.140 30.900 322.100 31.180 ;
        RECT 320.140 30.850 320.420 30.900 ;
        RECT 321.260 27.260 321.540 27.310 ;
        RECT 319.020 26.980 321.540 27.260 ;
        RECT 321.260 26.930 321.540 26.980 ;
        RECT 320.700 26.140 320.980 26.190 ;
        RECT 317.340 25.860 318.180 26.140 ;
        RECT 316.780 19.420 317.060 19.470 ;
        RECT 317.900 19.420 318.180 25.860 ;
        RECT 316.780 19.140 318.180 19.420 ;
        RECT 319.020 25.860 320.980 26.140 ;
        RECT 316.780 17.970 317.060 19.140 ;
        RECT 316.780 6.210 317.060 7.710 ;
        RECT 318.460 7.330 318.740 11.630 ;
        RECT 317.900 3.970 318.180 6.590 ;
        RECT 319.020 4.300 319.300 25.860 ;
        RECT 320.700 25.810 320.980 25.860 ;
        RECT 321.820 24.130 322.100 30.900 ;
        RECT 332.460 30.060 332.740 30.110 ;
        RECT 333.020 30.060 333.300 37.950 ;
        RECT 332.460 29.780 333.300 30.060 ;
        RECT 331.340 26.230 331.620 26.750 ;
        RECT 332.460 19.650 332.740 29.780 ;
        RECT 333.020 26.930 333.300 28.430 ;
        RECT 320.140 10.740 320.420 14.990 ;
        RECT 320.700 13.910 320.980 14.430 ;
        RECT 321.260 12.700 321.540 14.430 ;
        RECT 321.260 12.420 322.660 12.700 ;
        RECT 321.260 11.110 321.540 11.630 ;
        RECT 320.140 10.460 322.100 10.740 ;
        RECT 319.580 7.190 319.860 7.710 ;
        RECT 321.820 6.770 322.100 10.460 ;
        RECT 322.380 6.770 322.660 12.420 ;
        RECT 323.500 11.810 323.780 19.470 ;
        RECT 324.060 18.950 324.340 19.470 ;
        RECT 325.180 15.170 325.460 19.470 ;
        RECT 326.300 15.730 326.580 19.470 ;
        RECT 326.860 14.470 327.140 14.990 ;
        RECT 325.180 12.370 325.460 14.430 ;
        RECT 325.740 12.370 326.020 14.430 ;
        RECT 324.620 12.140 324.900 12.190 ;
        RECT 324.060 11.860 324.900 12.140 ;
        RECT 324.060 10.740 324.340 11.860 ;
        RECT 324.620 11.810 324.900 11.860 ;
        RECT 327.420 11.670 327.700 12.190 ;
        RECT 325.740 11.110 326.020 11.630 ;
        RECT 323.500 10.460 324.340 10.740 ;
        RECT 323.500 7.330 323.780 10.460 ;
        RECT 321.820 4.390 322.100 4.910 ;
        RECT 326.300 4.530 326.580 11.630 ;
        RECT 327.420 6.540 327.700 6.590 ;
        RECT 326.860 6.260 327.700 6.540 ;
        RECT 326.860 4.530 327.140 6.260 ;
        RECT 327.420 6.070 327.700 6.260 ;
        RECT 329.100 4.860 329.380 18.350 ;
        RECT 329.660 7.750 329.940 8.270 ;
        RECT 329.660 4.860 329.940 4.910 ;
        RECT 329.100 4.580 329.940 4.860 ;
        RECT 318.460 4.020 319.300 4.300 ;
        RECT 318.460 3.180 318.740 4.020 ;
        RECT 313.980 -29.020 314.820 -28.740 ;
        RECT 315.100 2.900 318.740 3.180 ;
        RECT 315.100 -28.740 315.380 2.900 ;
        RECT 316.220 -3.310 316.500 -0.690 ;
        RECT 317.340 -3.310 317.620 -0.130 ;
        RECT 318.460 -3.310 318.740 -0.690 ;
        RECT 319.020 -1.860 319.300 3.230 ;
        RECT 321.260 3.180 321.540 3.230 ;
        RECT 319.580 2.900 321.540 3.180 ;
        RECT 319.580 -0.650 319.860 2.900 ;
        RECT 321.260 2.850 321.540 2.900 ;
        RECT 324.620 3.180 324.900 3.230 ;
        RECT 324.620 2.900 325.460 3.180 ;
        RECT 324.620 2.710 324.900 2.900 ;
        RECT 319.020 -2.140 319.860 -1.860 ;
        RECT 319.020 -4.010 319.300 -3.490 ;
        RECT 319.580 -4.100 319.860 -2.140 ;
        RECT 320.140 -3.310 320.420 -1.250 ;
        RECT 320.700 -2.190 320.980 -1.250 ;
        RECT 321.820 -4.010 322.100 -3.490 ;
        RECT 320.700 -4.100 320.980 -4.050 ;
        RECT 319.580 -4.380 320.980 -4.100 ;
        RECT 320.700 -4.430 320.980 -4.380 ;
        RECT 321.260 -6.340 321.540 -4.610 ;
        RECT 323.500 -4.990 323.780 -1.250 ;
        RECT 325.180 -2.980 325.460 2.900 ;
        RECT 329.100 -0.510 329.380 4.580 ;
        RECT 329.660 4.530 329.940 4.580 ;
        RECT 331.900 4.530 332.180 7.150 ;
        RECT 330.780 3.270 331.060 3.790 ;
        RECT 331.340 -1.630 331.620 -0.130 ;
        RECT 325.740 -2.980 326.020 -2.930 ;
        RECT 325.180 -3.260 326.020 -2.980 ;
        RECT 325.740 -3.450 326.020 -3.260 ;
        RECT 328.540 -3.450 328.820 -2.930 ;
        RECT 324.060 -4.100 324.340 -4.050 ;
        RECT 324.620 -4.100 324.900 -3.490 ;
        RECT 324.060 -4.380 324.900 -4.100 ;
        RECT 324.060 -4.430 324.340 -4.380 ;
        RECT 326.300 -4.990 326.580 -4.050 ;
        RECT 321.260 -6.620 323.780 -6.340 ;
        RECT 321.820 -16.190 322.100 -7.970 ;
        RECT 323.500 -8.350 323.780 -6.620 ;
        RECT 330.780 -15.630 331.060 -4.610 ;
        RECT 323.500 -15.860 323.780 -15.810 ;
        RECT 323.500 -16.140 324.340 -15.860 ;
        RECT 323.500 -16.190 323.780 -16.140 ;
        RECT 321.820 -17.450 322.100 -16.930 ;
        RECT 319.020 -19.130 319.300 -18.610 ;
        RECT 323.500 -18.660 323.780 -18.610 ;
        RECT 322.380 -18.940 323.780 -18.660 ;
        RECT 321.820 -19.690 322.100 -19.170 ;
        RECT 322.380 -22.020 322.660 -18.940 ;
        RECT 323.500 -18.990 323.780 -18.940 ;
        RECT 321.260 -22.300 322.660 -22.020 ;
        RECT 319.580 -23.610 319.860 -23.090 ;
        RECT 321.260 -23.470 321.540 -22.300 ;
        RECT 319.020 -27.530 319.300 -27.010 ;
        RECT 316.780 -27.620 317.060 -27.570 ;
        RECT 318.460 -27.620 318.740 -27.570 ;
        RECT 316.780 -27.900 318.740 -27.620 ;
        RECT 316.780 -27.950 317.060 -27.900 ;
        RECT 318.460 -28.090 318.740 -27.900 ;
        RECT 315.100 -29.020 318.740 -28.740 ;
        RECT 312.860 -31.540 313.140 -31.490 ;
        RECT 313.980 -31.540 314.260 -29.020 ;
        RECT 310.620 -31.820 314.260 -31.540 ;
        RECT 310.620 -39.380 310.900 -31.820 ;
        RECT 312.860 -31.870 313.140 -31.820 ;
        RECT 314.540 -38.260 314.820 -29.810 ;
        RECT 317.340 -30.890 317.620 -30.370 ;
        RECT 315.100 -34.670 315.380 -31.490 ;
        RECT 317.900 -34.670 318.180 -32.610 ;
        RECT 317.900 -38.260 318.180 -38.210 ;
        RECT 314.540 -38.540 318.180 -38.260 ;
        RECT 317.900 -38.590 318.180 -38.540 ;
        RECT 312.860 -39.290 313.140 -38.770 ;
        RECT 310.620 -39.660 311.460 -39.380 ;
        RECT 310.620 -39.710 310.900 -39.660 ;
        RECT 311.180 -43.300 311.460 -39.660 ;
        RECT 312.300 -40.500 312.580 -40.450 ;
        RECT 312.300 -40.780 313.140 -40.500 ;
        RECT 312.300 -40.830 312.580 -40.780 ;
        RECT 312.300 -43.300 312.580 -43.250 ;
        RECT 311.180 -43.580 312.580 -43.300 ;
        RECT 312.300 -43.630 312.580 -43.580 ;
        RECT 312.300 -47.220 312.580 -47.170 ;
        RECT 312.860 -47.220 313.140 -40.780 ;
        RECT 315.100 -44.190 315.380 -43.250 ;
        RECT 317.340 -43.630 317.620 -39.330 ;
        RECT 312.300 -47.500 313.140 -47.220 ;
        RECT 318.460 -47.220 318.740 -29.020 ;
        RECT 319.020 -30.420 319.300 -30.370 ;
        RECT 319.580 -30.420 319.860 -26.450 ;
        RECT 319.020 -30.700 319.860 -30.420 ;
        RECT 319.020 -30.750 319.300 -30.700 ;
        RECT 320.140 -32.660 320.420 -24.770 ;
        RECT 322.380 -26.830 322.660 -24.770 ;
        RECT 321.260 -30.420 321.540 -27.570 ;
        RECT 322.940 -30.420 323.220 -19.730 ;
        RECT 324.060 -19.780 324.340 -16.140 ;
        RECT 324.620 -16.420 324.900 -16.370 ;
        RECT 324.620 -16.700 325.460 -16.420 ;
        RECT 324.620 -16.750 324.900 -16.700 ;
        RECT 324.620 -19.780 324.900 -19.730 ;
        RECT 324.060 -20.060 324.900 -19.780 ;
        RECT 324.620 -20.670 324.900 -20.060 ;
        RECT 325.180 -20.110 325.460 -16.700 ;
        RECT 326.860 -20.340 327.140 -16.930 ;
        RECT 327.980 -20.340 328.260 -20.290 ;
        RECT 326.860 -20.620 328.260 -20.340 ;
        RECT 327.980 -20.810 328.260 -20.620 ;
        RECT 325.180 -27.530 325.460 -27.010 ;
        RECT 324.060 -28.090 324.340 -27.570 ;
        RECT 321.260 -30.700 323.220 -30.420 ;
        RECT 320.700 -31.450 320.980 -30.930 ;
        RECT 321.260 -32.660 321.540 -32.610 ;
        RECT 320.140 -32.940 321.540 -32.660 ;
        RECT 321.260 -34.670 321.540 -32.940 ;
        RECT 322.380 -34.670 322.660 -32.050 ;
        RECT 322.940 -34.900 323.220 -30.700 ;
        RECT 327.980 -32.010 328.260 -31.490 ;
        RECT 323.500 -34.900 323.780 -34.850 ;
        RECT 322.940 -35.180 323.780 -34.900 ;
        RECT 319.020 -35.460 319.300 -35.410 ;
        RECT 320.140 -35.460 320.420 -35.410 ;
        RECT 321.820 -35.460 322.100 -35.410 ;
        RECT 319.020 -35.740 320.420 -35.460 ;
        RECT 319.020 -35.790 319.300 -35.740 ;
        RECT 319.020 -43.630 319.300 -36.530 ;
        RECT 319.580 -38.590 319.860 -35.740 ;
        RECT 320.140 -35.790 320.420 -35.740 ;
        RECT 320.700 -35.740 322.100 -35.460 ;
        RECT 320.700 -39.150 320.980 -35.740 ;
        RECT 321.820 -35.930 322.100 -35.740 ;
        RECT 323.500 -35.790 323.780 -35.180 ;
        RECT 325.180 -36.490 325.460 -35.970 ;
        RECT 322.940 -39.290 323.220 -38.770 ;
        RECT 326.300 -40.270 326.580 -32.050 ;
        RECT 329.100 -32.430 329.380 -15.810 ;
        RECT 330.780 -16.980 331.060 -16.930 ;
        RECT 331.900 -16.980 332.180 -15.810 ;
        RECT 330.780 -17.260 332.180 -16.980 ;
        RECT 330.780 -20.110 331.060 -17.260 ;
        RECT 327.980 -39.710 328.260 -38.210 ;
        RECT 330.220 -39.380 330.500 -39.330 ;
        RECT 330.780 -39.380 331.060 -31.490 ;
        RECT 331.340 -31.870 331.620 -28.130 ;
        RECT 331.900 -35.790 332.180 -32.050 ;
        RECT 330.220 -39.660 331.060 -39.380 ;
        RECT 332.460 -39.380 332.740 -39.330 ;
        RECT 333.020 -39.380 333.300 -35.970 ;
        RECT 332.460 -39.660 333.300 -39.380 ;
        RECT 330.220 -39.710 330.500 -39.660 ;
        RECT 332.460 -39.710 332.740 -39.660 ;
        RECT 331.900 -42.510 332.180 -39.890 ;
        RECT 333.580 -45.540 333.860 41.870 ;
        RECT 336.940 39.580 337.220 39.630 ;
        RECT 338.060 39.580 338.340 39.630 ;
        RECT 336.940 39.300 338.340 39.580 ;
        RECT 336.940 39.250 337.220 39.300 ;
        RECT 338.060 38.690 338.340 39.300 ;
        RECT 338.620 39.020 338.900 42.100 ;
        RECT 339.180 39.810 339.460 41.870 ;
        RECT 339.180 39.020 339.460 39.070 ;
        RECT 338.620 38.740 339.460 39.020 ;
        RECT 339.180 38.550 339.460 38.740 ;
        RECT 339.740 35.940 340.020 37.950 ;
        RECT 337.500 32.300 337.780 35.710 ;
        RECT 338.060 35.190 338.340 35.710 ;
        RECT 338.620 35.660 340.020 35.940 ;
        RECT 338.620 35.330 338.900 35.660 ;
        RECT 340.860 32.300 341.140 34.590 ;
        RECT 337.500 32.020 341.140 32.300 ;
        RECT 335.820 31.460 337.780 31.740 ;
        RECT 335.260 28.610 335.540 30.670 ;
        RECT 334.140 27.820 334.420 27.870 ;
        RECT 335.820 27.820 336.100 31.460 ;
        RECT 337.500 30.850 337.780 31.460 ;
        RECT 336.380 30.150 336.660 30.670 ;
        RECT 337.500 27.910 337.780 28.430 ;
        RECT 334.140 27.540 336.100 27.820 ;
        RECT 334.140 27.490 334.420 27.540 ;
        RECT 334.700 26.930 334.980 27.540 ;
        RECT 338.620 25.580 338.900 30.110 ;
        RECT 335.260 25.300 338.900 25.580 ;
        RECT 334.140 23.570 334.420 24.510 ;
        RECT 335.260 24.130 335.540 25.300 ;
        RECT 334.140 22.310 334.420 22.830 ;
        RECT 337.500 22.310 337.780 22.830 ;
        RECT 339.180 22.780 339.460 32.020 ;
        RECT 341.420 31.740 341.700 39.070 ;
        RECT 339.740 31.460 341.700 31.740 ;
        RECT 339.740 30.850 340.020 31.460 ;
        RECT 341.420 31.410 341.700 31.460 ;
        RECT 340.300 27.260 340.580 27.310 ;
        RECT 341.980 27.260 342.260 35.710 ;
        RECT 343.660 31.970 343.940 37.950 ;
        RECT 350.380 35.940 350.660 41.870 ;
        RECT 350.380 35.660 352.900 35.940 ;
        RECT 345.340 34.630 345.620 35.150 ;
        RECT 349.260 31.970 349.540 35.150 ;
        RECT 349.820 31.410 350.100 34.590 ;
        RECT 343.660 27.820 343.940 30.110 ;
        RECT 343.660 27.540 345.060 27.820 ;
        RECT 340.300 26.980 342.260 27.260 ;
        RECT 342.540 27.260 342.820 27.310 ;
        RECT 342.540 26.980 343.940 27.260 ;
        RECT 340.300 26.930 340.580 26.980 ;
        RECT 342.540 26.930 342.820 26.980 ;
        RECT 343.660 24.130 343.940 26.980 ;
        RECT 344.220 22.870 344.500 23.390 ;
        RECT 339.740 22.780 340.020 22.830 ;
        RECT 339.180 22.500 340.020 22.780 ;
        RECT 339.740 22.450 340.020 22.500 ;
        RECT 341.420 15.500 341.700 15.550 ;
        RECT 340.300 15.220 341.700 15.500 ;
        RECT 340.300 7.890 340.580 15.220 ;
        RECT 341.420 15.170 341.700 15.220 ;
        RECT 342.540 10.740 342.820 20.030 ;
        RECT 343.100 15.170 343.380 15.690 ;
        RECT 343.100 13.910 343.380 14.430 ;
        RECT 341.420 7.890 341.700 10.510 ;
        RECT 342.540 10.460 343.940 10.740 ;
        RECT 339.180 6.210 339.460 7.150 ;
        RECT 343.660 -1.630 343.940 10.460 ;
        RECT 344.220 8.450 344.500 15.550 ;
        RECT 344.780 11.810 345.060 27.540 ;
        RECT 346.460 20.210 346.740 23.390 ;
        RECT 347.580 23.010 347.860 27.310 ;
        RECT 348.140 22.870 348.420 23.390 ;
        RECT 344.780 6.770 345.060 8.270 ;
        RECT 345.340 7.100 345.620 14.990 ;
        RECT 349.260 14.940 349.540 23.390 ;
        RECT 350.940 20.210 351.220 22.270 ;
        RECT 349.260 14.660 350.660 14.940 ;
        RECT 349.260 14.610 349.540 14.660 ;
        RECT 346.460 11.110 346.740 11.630 ;
        RECT 345.900 7.100 346.180 7.150 ;
        RECT 345.340 6.820 346.180 7.100 ;
        RECT 335.260 -8.910 335.540 -4.050 ;
        RECT 336.940 -4.430 337.220 -3.490 ;
        RECT 335.260 -23.470 335.540 -15.810 ;
        RECT 338.620 -32.660 338.900 -4.050 ;
        RECT 339.180 -7.230 339.460 -2.930 ;
        RECT 345.340 -7.790 345.620 6.820 ;
        RECT 345.900 6.770 346.180 6.820 ;
        RECT 346.460 2.850 346.740 3.790 ;
        RECT 348.700 3.740 348.980 3.790 ;
        RECT 347.020 3.460 348.980 3.740 ;
        RECT 346.460 0.940 346.740 0.990 ;
        RECT 347.020 0.940 347.300 3.460 ;
        RECT 348.700 3.410 348.980 3.460 ;
        RECT 346.460 0.660 347.300 0.940 ;
        RECT 347.580 0.940 347.860 0.990 ;
        RECT 348.140 0.940 348.420 2.670 ;
        RECT 347.580 0.660 348.420 0.940 ;
        RECT 346.460 0.610 346.740 0.660 ;
        RECT 347.580 0.470 347.860 0.660 ;
        RECT 349.260 -3.310 349.540 -0.130 ;
        RECT 350.380 -0.180 350.660 14.660 ;
        RECT 350.940 2.710 351.220 3.230 ;
        RECT 350.940 -0.180 351.220 -0.130 ;
        RECT 350.380 -0.460 351.220 -0.180 ;
        RECT 350.940 -0.510 351.220 -0.460 ;
        RECT 346.460 -4.010 346.740 -3.490 ;
        RECT 345.900 -10.820 346.180 -4.050 ;
        RECT 347.020 -4.570 347.300 -4.050 ;
        RECT 347.580 -10.820 347.860 -10.770 ;
        RECT 345.900 -11.100 347.860 -10.820 ;
        RECT 347.580 -11.150 347.860 -11.100 ;
        RECT 349.260 -12.270 349.540 -4.610 ;
        RECT 349.820 -6.670 350.100 -1.250 ;
        RECT 350.380 -1.770 350.660 -1.250 ;
        RECT 351.500 -3.870 351.780 0.430 ;
        RECT 350.940 -4.570 351.220 -4.050 ;
        RECT 350.380 -15.300 350.660 -15.250 ;
        RECT 352.060 -15.300 352.340 -11.330 ;
        RECT 350.380 -15.580 352.340 -15.300 ;
        RECT 350.380 -15.630 350.660 -15.580 ;
        RECT 352.060 -16.190 352.340 -15.580 ;
        RECT 346.460 -18.660 346.740 -16.930 ;
        RECT 346.460 -18.940 347.300 -18.660 ;
        RECT 346.460 -18.990 346.740 -18.940 ;
        RECT 338.620 -32.940 339.460 -32.660 ;
        RECT 337.500 -34.340 337.780 -34.290 ;
        RECT 338.620 -34.340 338.900 -33.730 ;
        RECT 337.500 -34.620 338.900 -34.340 ;
        RECT 337.500 -34.810 337.780 -34.620 ;
        RECT 336.940 -37.050 337.220 -36.530 ;
        RECT 338.620 -42.510 338.900 -36.530 ;
        RECT 339.180 -39.380 339.460 -32.940 ;
        RECT 342.540 -33.130 342.820 -32.610 ;
        RECT 343.660 -33.780 343.940 -24.770 ;
        RECT 345.340 -25.290 345.620 -24.770 ;
        RECT 346.460 -31.870 346.740 -27.010 ;
        RECT 342.540 -34.060 343.940 -33.780 ;
        RECT 339.180 -39.660 340.020 -39.380 ;
        RECT 334.700 -43.770 334.980 -43.250 ;
        RECT 338.620 -43.860 338.900 -43.810 ;
        RECT 339.180 -43.860 339.460 -40.450 ;
        RECT 339.740 -43.300 340.020 -39.660 ;
        RECT 342.540 -43.070 342.820 -34.060 ;
        RECT 344.780 -40.830 345.060 -32.610 ;
        RECT 347.020 -40.270 347.300 -18.940 ;
        RECT 352.620 -22.580 352.900 35.660 ;
        RECT 355.420 35.330 355.700 42.990 ;
        RECT 358.780 42.940 359.060 42.990 ;
        RECT 358.780 42.660 361.300 42.940 ;
        RECT 358.780 42.610 359.060 42.660 ;
        RECT 361.020 39.810 361.300 42.660 ;
        RECT 360.460 35.890 360.740 39.070 ;
        RECT 361.580 37.990 361.860 38.510 ;
        RECT 363.260 36.220 363.540 39.070 ;
        RECT 365.500 38.550 365.780 39.070 ;
        RECT 364.940 37.990 365.220 38.510 ;
        RECT 363.820 36.220 364.100 36.270 ;
        RECT 363.260 35.940 364.100 36.220 ;
        RECT 363.820 35.890 364.100 35.940 ;
        RECT 364.380 35.940 364.660 37.950 ;
        RECT 354.860 28.380 355.140 28.430 ;
        RECT 356.540 28.380 356.820 35.710 ;
        RECT 364.380 35.660 365.220 35.940 ;
        RECT 360.460 30.290 360.740 35.150 ;
        RECT 354.860 28.100 356.820 28.380 ;
        RECT 354.860 28.050 355.140 28.100 ;
        RECT 357.660 26.790 357.940 27.310 ;
        RECT 361.580 26.930 361.860 35.150 ;
        RECT 362.140 21.890 362.420 30.670 ;
        RECT 362.700 28.380 362.980 35.150 ;
        RECT 364.380 34.630 364.660 35.150 ;
        RECT 363.260 34.070 363.540 34.590 ;
        RECT 363.260 30.710 363.540 31.230 ;
        RECT 363.260 28.380 363.540 28.430 ;
        RECT 362.700 28.100 364.660 28.380 ;
        RECT 363.260 28.050 363.540 28.100 ;
        RECT 364.380 20.540 364.660 28.100 ;
        RECT 364.940 28.050 365.220 35.660 ;
        RECT 366.060 34.770 366.340 37.950 ;
        RECT 369.980 35.330 370.260 43.550 ;
        RECT 373.900 38.690 374.180 41.870 ;
        RECT 377.820 39.810 378.100 41.870 ;
        RECT 378.940 41.490 379.220 42.430 ;
        RECT 381.740 42.380 382.020 42.430 ;
        RECT 383.420 42.380 383.700 43.780 ;
        RECT 392.380 43.730 392.660 43.780 ;
        RECT 383.980 42.940 384.260 42.990 ;
        RECT 383.980 42.660 385.380 42.940 ;
        RECT 383.980 42.610 384.260 42.660 ;
        RECT 381.740 42.100 383.700 42.380 ;
        RECT 381.740 35.940 382.020 42.100 ;
        RECT 385.100 40.140 385.380 42.660 ;
        RECT 385.660 41.490 385.940 42.990 ;
        RECT 386.220 40.140 386.500 40.190 ;
        RECT 385.100 39.860 386.500 40.140 ;
        RECT 386.220 39.810 386.500 39.860 ;
        RECT 366.620 31.180 366.900 31.230 ;
        RECT 366.620 30.900 369.700 31.180 ;
        RECT 366.620 30.850 366.900 30.900 ;
        RECT 369.420 28.050 369.700 30.900 ;
        RECT 369.980 26.930 370.260 30.110 ;
        RECT 377.820 27.260 378.100 35.710 ;
        RECT 381.740 35.660 382.580 35.940 ;
        RECT 381.740 30.150 382.020 30.670 ;
        RECT 378.940 27.260 379.220 27.310 ;
        RECT 377.820 26.980 379.220 27.260 ;
        RECT 378.940 26.930 379.220 26.980 ;
        RECT 369.980 22.220 370.260 22.270 ;
        RECT 369.980 21.940 370.820 22.220 ;
        RECT 369.980 21.890 370.260 21.940 ;
        RECT 365.500 20.540 365.780 20.590 ;
        RECT 362.700 20.260 365.780 20.540 ;
        RECT 357.100 11.250 357.380 14.430 ;
        RECT 359.340 10.690 359.620 11.630 ;
        RECT 355.980 3.410 356.260 10.510 ;
        RECT 358.780 3.740 359.060 3.790 ;
        RECT 358.780 3.460 359.620 3.740 ;
        RECT 358.780 3.410 359.060 3.460 ;
        RECT 353.740 -11.710 354.020 -1.250 ;
        RECT 356.540 -4.990 356.820 0.990 ;
        RECT 359.340 0.380 359.620 3.460 ;
        RECT 362.140 0.380 362.420 0.430 ;
        RECT 359.340 0.100 362.420 0.380 ;
        RECT 362.140 0.050 362.420 0.100 ;
        RECT 358.220 -1.300 358.500 -0.690 ;
        RECT 361.580 -0.740 361.860 -0.690 ;
        RECT 361.580 -1.020 362.420 -0.740 ;
        RECT 361.580 -1.070 361.860 -1.020 ;
        RECT 358.780 -1.300 359.060 -1.250 ;
        RECT 358.220 -1.580 359.060 -1.300 ;
        RECT 358.780 -1.630 359.060 -1.580 ;
        RECT 362.140 -3.310 362.420 -1.020 ;
        RECT 361.580 -4.100 361.860 -4.050 ;
        RECT 359.900 -4.380 361.860 -4.100 ;
        RECT 353.180 -16.190 353.460 -11.890 ;
        RECT 359.900 -15.630 360.180 -4.380 ;
        RECT 361.580 -4.430 361.860 -4.380 ;
        RECT 362.700 -4.430 362.980 20.260 ;
        RECT 365.500 20.210 365.780 20.260 ;
        RECT 367.180 19.090 367.460 20.030 ;
        RECT 369.420 18.530 369.700 19.470 ;
        RECT 368.860 18.300 369.140 18.350 ;
        RECT 366.620 18.020 369.140 18.300 ;
        RECT 363.260 10.690 363.540 15.550 ;
        RECT 363.820 10.740 364.100 15.550 ;
        RECT 366.620 15.170 366.900 18.020 ;
        RECT 368.860 17.970 369.140 18.020 ;
        RECT 367.180 11.020 367.460 12.190 ;
        RECT 368.860 12.140 369.140 12.190 ;
        RECT 370.540 12.140 370.820 21.940 ;
        RECT 368.860 11.860 370.820 12.140 ;
        RECT 368.860 11.810 369.140 11.860 ;
        RECT 370.540 11.810 370.820 11.860 ;
        RECT 367.180 10.740 368.580 11.020 ;
        RECT 363.820 10.460 364.660 10.740 ;
        RECT 367.180 10.690 367.460 10.740 ;
        RECT 363.820 -0.510 364.100 0.430 ;
        RECT 363.260 -1.210 363.540 -0.690 ;
        RECT 360.460 -13.060 360.740 -5.170 ;
        RECT 361.020 -12.270 361.300 -8.530 ;
        RECT 361.580 -10.260 361.860 -5.730 ;
        RECT 363.820 -6.110 364.100 -5.170 ;
        RECT 364.380 -5.550 364.660 10.460 ;
        RECT 368.300 7.330 368.580 10.740 ;
        RECT 369.980 4.530 370.260 10.510 ;
        RECT 364.940 -8.020 365.220 -7.970 ;
        RECT 363.820 -8.300 365.220 -8.020 ;
        RECT 362.140 -9.050 362.420 -8.530 ;
        RECT 363.260 -9.050 363.540 -8.530 ;
        RECT 362.700 -9.610 362.980 -9.090 ;
        RECT 361.580 -10.540 362.420 -10.260 ;
        RECT 360.460 -13.340 361.300 -13.060 ;
        RECT 360.460 -16.890 360.740 -16.370 ;
        RECT 350.940 -22.860 352.900 -22.580 ;
        RECT 349.820 -26.970 350.100 -26.450 ;
        RECT 349.260 -27.530 349.540 -27.010 ;
        RECT 350.380 -34.340 350.660 -34.290 ;
        RECT 349.820 -34.620 350.660 -34.340 ;
        RECT 349.820 -35.230 350.100 -34.620 ;
        RECT 350.380 -34.670 350.660 -34.620 ;
        RECT 348.140 -36.020 348.420 -35.410 ;
        RECT 349.260 -36.020 349.540 -35.970 ;
        RECT 348.140 -36.300 349.540 -36.020 ;
        RECT 347.580 -38.260 347.860 -38.210 ;
        RECT 348.140 -38.260 348.420 -36.300 ;
        RECT 349.260 -36.350 349.540 -36.300 ;
        RECT 350.940 -37.140 351.220 -22.860 ;
        RECT 351.500 -24.730 351.780 -24.210 ;
        RECT 353.180 -24.730 353.460 -16.930 ;
        RECT 359.340 -17.450 359.620 -16.930 ;
        RECT 361.020 -20.110 361.300 -13.340 ;
        RECT 359.340 -23.610 359.620 -23.090 ;
        RECT 356.540 -23.700 356.820 -23.650 ;
        RECT 354.300 -23.980 356.820 -23.700 ;
        RECT 353.740 -25.290 354.020 -24.770 ;
        RECT 354.300 -26.970 354.580 -23.980 ;
        RECT 356.540 -24.030 356.820 -23.980 ;
        RECT 353.740 -27.950 354.020 -27.010 ;
        RECT 358.220 -27.060 358.500 -23.650 ;
        RECT 361.580 -24.170 361.860 -23.650 ;
        RECT 362.140 -24.260 362.420 -10.540 ;
        RECT 363.260 -10.820 363.540 -10.770 ;
        RECT 363.820 -10.820 364.100 -8.300 ;
        RECT 364.940 -8.350 365.220 -8.300 ;
        RECT 362.700 -11.100 364.100 -10.820 ;
        RECT 362.700 -15.070 362.980 -11.100 ;
        RECT 363.260 -11.150 363.540 -11.100 ;
        RECT 366.620 -11.290 366.900 -10.770 ;
        RECT 363.260 -24.030 363.540 -14.690 ;
        RECT 363.820 -16.330 364.100 -15.810 ;
        RECT 365.500 -20.250 365.780 -19.730 ;
        RECT 366.060 -24.030 366.340 -11.330 ;
        RECT 367.180 -15.860 367.460 2.670 ;
        RECT 367.740 -8.350 368.020 0.430 ;
        RECT 370.540 0.380 370.820 0.430 ;
        RECT 371.100 0.380 371.380 7.710 ;
        RECT 371.660 2.290 371.940 11.630 ;
        RECT 377.820 11.250 378.100 14.430 ;
        RECT 381.180 12.370 381.460 27.310 ;
        RECT 382.300 20.540 382.580 35.660 ;
        RECT 386.220 35.330 386.500 38.510 ;
        RECT 384.540 32.860 384.820 35.150 ;
        RECT 381.740 20.260 382.580 20.540 ;
        RECT 383.420 32.580 384.820 32.860 ;
        RECT 381.740 15.500 382.020 20.260 ;
        RECT 383.420 19.650 383.700 32.580 ;
        RECT 385.100 30.710 385.380 31.230 ;
        RECT 383.980 23.340 384.260 30.670 ;
        RECT 385.660 30.620 385.940 35.150 ;
        RECT 386.780 30.850 387.060 42.990 ;
        RECT 387.900 42.940 388.180 42.990 ;
        RECT 389.020 42.940 389.300 42.990 ;
        RECT 387.900 42.660 388.740 42.940 ;
        RECT 387.900 42.610 388.180 42.660 ;
        RECT 387.340 41.910 387.620 42.430 ;
        RECT 388.460 39.580 388.740 42.660 ;
        RECT 389.020 42.660 389.860 42.940 ;
        RECT 389.020 42.610 389.300 42.660 ;
        RECT 389.020 39.580 389.300 39.630 ;
        RECT 388.460 39.300 389.300 39.580 ;
        RECT 387.900 38.550 388.180 39.070 ;
        RECT 388.460 35.940 388.740 39.300 ;
        RECT 389.020 39.250 389.300 39.300 ;
        RECT 387.900 35.660 388.740 35.940 ;
        RECT 387.900 35.330 388.180 35.660 ;
        RECT 386.220 30.620 386.500 30.670 ;
        RECT 385.660 30.340 386.500 30.620 ;
        RECT 386.220 30.150 386.500 30.340 ;
        RECT 384.540 29.590 384.820 30.110 ;
        RECT 387.900 30.060 388.180 30.110 ;
        RECT 387.340 29.780 388.180 30.060 ;
        RECT 385.660 23.340 385.940 23.390 ;
        RECT 383.980 23.060 385.940 23.340 ;
        RECT 385.660 22.450 385.940 23.060 ;
        RECT 386.780 22.870 387.060 23.390 ;
        RECT 387.340 23.340 387.620 29.780 ;
        RECT 387.900 29.730 388.180 29.780 ;
        RECT 389.020 28.380 389.300 28.430 ;
        RECT 389.580 28.380 389.860 42.660 ;
        RECT 391.820 41.910 392.100 42.430 ;
        RECT 390.700 37.990 390.980 38.510 ;
        RECT 391.260 35.940 391.540 37.950 ;
        RECT 391.260 35.660 393.220 35.940 ;
        RECT 391.260 35.100 391.540 35.150 ;
        RECT 391.260 34.820 392.660 35.100 ;
        RECT 391.260 34.770 391.540 34.820 ;
        RECT 389.020 28.100 389.860 28.380 ;
        RECT 392.380 33.980 392.660 34.820 ;
        RECT 392.940 34.770 393.220 35.660 ;
        RECT 394.060 33.980 394.340 42.990 ;
        RECT 396.860 42.610 397.140 43.780 ;
        RECT 408.620 43.500 408.900 43.550 ;
        RECT 408.060 43.220 408.900 43.500 ;
        RECT 404.700 38.550 404.980 39.070 ;
        RECT 392.380 33.700 394.340 33.980 ;
        RECT 404.700 35.940 404.980 36.270 ;
        RECT 408.060 35.940 408.340 43.220 ;
        RECT 408.620 43.170 408.900 43.220 ;
        RECT 404.700 35.660 408.340 35.940 ;
        RECT 389.020 28.050 389.300 28.100 ;
        RECT 390.700 27.260 390.980 27.310 ;
        RECT 391.820 27.260 392.100 27.310 ;
        RECT 390.700 26.980 392.100 27.260 ;
        RECT 390.700 26.930 390.980 26.980 ;
        RECT 391.820 26.930 392.100 26.980 ;
        RECT 389.580 23.340 389.860 23.390 ;
        RECT 390.140 23.340 390.420 23.390 ;
        RECT 387.340 23.060 388.180 23.340 ;
        RECT 386.220 21.100 386.500 22.270 ;
        RECT 384.540 20.820 386.500 21.100 ;
        RECT 382.300 18.950 382.580 19.470 ;
        RECT 381.740 15.220 382.580 15.500 ;
        RECT 381.740 13.910 382.020 14.430 ;
        RECT 382.300 6.540 382.580 15.220 ;
        RECT 382.860 14.050 383.140 19.470 ;
        RECT 383.980 19.420 384.260 19.470 ;
        RECT 384.540 19.420 384.820 20.820 ;
        RECT 385.100 19.980 385.380 20.030 ;
        RECT 387.340 19.980 387.620 22.270 ;
        RECT 385.100 19.700 387.620 19.980 ;
        RECT 385.100 19.650 385.380 19.700 ;
        RECT 383.980 19.140 384.820 19.420 ;
        RECT 383.420 18.390 383.700 18.910 ;
        RECT 383.980 17.970 384.260 19.140 ;
        RECT 387.900 19.090 388.180 23.060 ;
        RECT 389.580 23.060 390.420 23.340 ;
        RECT 389.580 23.010 389.860 23.060 ;
        RECT 390.140 23.010 390.420 23.060 ;
        RECT 390.700 20.540 390.980 22.270 ;
        RECT 390.700 20.260 392.100 20.540 ;
        RECT 389.580 18.950 389.860 19.470 ;
        RECT 391.820 19.090 392.100 20.260 ;
        RECT 392.380 19.090 392.660 33.700 ;
        RECT 393.500 32.300 393.780 32.350 ;
        RECT 392.940 32.020 393.780 32.300 ;
        RECT 391.260 14.380 391.540 14.430 ;
        RECT 390.140 14.100 391.540 14.380 ;
        RECT 382.860 11.020 383.140 11.630 ;
        RECT 386.220 11.250 386.500 12.750 ;
        RECT 388.460 12.230 388.740 12.750 ;
        RECT 389.580 11.580 389.860 11.630 ;
        RECT 390.140 11.580 390.420 14.100 ;
        RECT 391.260 14.050 391.540 14.100 ;
        RECT 392.380 12.700 392.660 12.750 ;
        RECT 392.940 12.700 393.220 32.020 ;
        RECT 393.500 31.970 393.780 32.020 ;
        RECT 392.380 12.420 393.220 12.700 ;
        RECT 392.380 11.810 392.660 12.420 ;
        RECT 389.020 11.300 390.420 11.580 ;
        RECT 383.980 11.020 384.260 11.070 ;
        RECT 382.860 10.740 384.260 11.020 ;
        RECT 382.860 6.770 383.140 10.740 ;
        RECT 383.980 10.690 384.260 10.740 ;
        RECT 386.780 6.540 387.060 6.590 ;
        RECT 381.740 6.260 382.580 6.540 ;
        RECT 386.220 6.260 387.060 6.540 ;
        RECT 373.900 2.150 374.180 2.670 ;
        RECT 370.540 0.100 371.380 0.380 ;
        RECT 370.540 0.050 370.820 0.100 ;
        RECT 368.300 -0.650 368.580 -0.130 ;
        RECT 369.420 -1.210 369.700 -0.690 ;
        RECT 371.100 -0.740 371.380 -0.690 ;
        RECT 369.980 -1.020 371.380 -0.740 ;
        RECT 369.980 -3.310 370.260 -1.020 ;
        RECT 371.100 -1.070 371.380 -1.020 ;
        RECT 368.300 -12.270 368.580 -9.090 ;
        RECT 369.420 -12.830 369.700 -3.490 ;
        RECT 370.540 -5.220 370.820 -5.170 ;
        RECT 370.540 -5.500 371.940 -5.220 ;
        RECT 370.540 -5.550 370.820 -5.500 ;
        RECT 371.100 -11.850 371.380 -11.330 ;
        RECT 371.660 -15.300 371.940 -5.500 ;
        RECT 372.220 -12.270 372.500 -0.690 ;
        RECT 368.300 -15.580 371.940 -15.300 ;
        RECT 367.180 -16.140 368.020 -15.860 ;
        RECT 362.700 -24.260 362.980 -24.210 ;
        RECT 362.140 -24.540 362.980 -24.260 ;
        RECT 362.700 -24.590 362.980 -24.540 ;
        RECT 367.180 -24.590 367.460 -16.930 ;
        RECT 367.740 -22.860 368.020 -16.140 ;
        RECT 368.300 -20.110 368.580 -15.580 ;
        RECT 371.660 -15.630 371.940 -15.580 ;
        RECT 370.540 -19.780 370.820 -16.370 ;
        RECT 372.220 -18.990 372.500 -15.810 ;
        RECT 372.780 -19.550 373.060 -16.370 ;
        RECT 371.660 -19.780 371.940 -19.730 ;
        RECT 370.540 -20.060 371.940 -19.780 ;
        RECT 371.660 -20.250 371.940 -20.060 ;
        RECT 367.740 -23.140 371.940 -22.860 ;
        RECT 358.780 -25.290 359.060 -24.770 ;
        RECT 358.220 -27.340 359.620 -27.060 ;
        RECT 358.220 -27.390 358.500 -27.340 ;
        RECT 355.420 -27.620 355.700 -27.570 ;
        RECT 355.420 -27.900 356.820 -27.620 ;
        RECT 355.420 -28.090 355.700 -27.900 ;
        RECT 354.860 -28.650 355.140 -28.130 ;
        RECT 352.060 -28.740 352.340 -28.690 ;
        RECT 352.060 -29.020 352.900 -28.740 ;
        RECT 352.060 -29.070 352.340 -29.020 ;
        RECT 352.060 -35.790 352.340 -30.370 ;
        RECT 352.620 -34.340 352.900 -29.020 ;
        RECT 356.540 -30.420 356.820 -27.900 ;
        RECT 356.540 -30.700 357.940 -30.420 ;
        RECT 356.540 -30.890 356.820 -30.700 ;
        RECT 353.180 -34.340 353.460 -34.290 ;
        RECT 352.620 -34.620 353.460 -34.340 ;
        RECT 352.620 -34.810 352.900 -34.620 ;
        RECT 353.180 -34.670 353.460 -34.620 ;
        RECT 357.660 -34.670 357.940 -30.700 ;
        RECT 354.300 -35.790 354.580 -34.850 ;
        RECT 355.420 -35.460 355.700 -35.410 ;
        RECT 355.420 -35.740 356.820 -35.460 ;
        RECT 355.420 -35.930 355.700 -35.740 ;
        RECT 352.620 -36.490 352.900 -35.970 ;
        RECT 350.940 -37.420 352.900 -37.140 ;
        RECT 347.580 -38.540 348.420 -38.260 ;
        RECT 347.580 -38.590 347.860 -38.540 ;
        RECT 343.100 -42.650 343.380 -42.130 ;
        RECT 344.220 -43.210 344.500 -42.690 ;
        RECT 349.820 -43.210 350.100 -42.690 ;
        RECT 340.300 -43.300 340.580 -43.250 ;
        RECT 339.740 -43.580 340.580 -43.300 ;
        RECT 340.300 -43.630 340.580 -43.580 ;
        RECT 344.780 -43.770 345.060 -43.250 ;
        RECT 348.700 -43.770 348.980 -43.250 ;
        RECT 338.620 -44.140 339.460 -43.860 ;
        RECT 338.620 -44.190 338.900 -44.140 ;
        RECT 347.020 -44.330 347.300 -43.810 ;
        RECT 333.580 -45.820 336.100 -45.540 ;
        RECT 333.580 -46.990 333.860 -45.820 ;
        RECT 319.020 -47.220 319.300 -47.170 ;
        RECT 318.460 -47.500 319.300 -47.220 ;
        RECT 312.300 -47.550 312.580 -47.500 ;
        RECT 319.020 -47.550 319.300 -47.500 ;
        RECT 316.220 -61.000 316.500 -47.730 ;
        RECT 322.380 -48.670 322.660 -47.730 ;
        RECT 334.140 -61.000 334.420 -46.610 ;
        RECT 335.820 -47.550 336.100 -45.820 ;
        RECT 340.860 -47.130 341.140 -46.610 ;
        RECT 352.060 -61.000 352.340 -46.610 ;
        RECT 352.620 -46.660 352.900 -37.420 ;
        RECT 356.540 -38.260 356.820 -35.740 ;
        RECT 358.780 -35.930 359.060 -35.410 ;
        RECT 359.340 -35.790 359.620 -27.340 ;
        RECT 359.900 -27.950 360.180 -24.770 ;
        RECT 364.940 -27.950 365.220 -27.010 ;
        RECT 365.500 -34.110 365.780 -24.770 ;
        RECT 366.620 -32.430 366.900 -27.570 ;
        RECT 371.100 -30.890 371.380 -30.370 ;
        RECT 369.420 -32.660 369.700 -32.610 ;
        RECT 368.860 -32.940 369.700 -32.660 ;
        RECT 363.260 -35.230 363.540 -34.290 ;
        RECT 358.220 -36.580 358.500 -35.970 ;
        RECT 361.020 -36.580 361.300 -36.530 ;
        RECT 362.700 -36.580 362.980 -36.530 ;
        RECT 358.220 -36.860 359.620 -36.580 ;
        RECT 357.100 -38.260 357.380 -38.210 ;
        RECT 356.540 -38.540 357.380 -38.260 ;
        RECT 357.100 -38.590 357.380 -38.540 ;
        RECT 356.540 -39.940 356.820 -39.890 ;
        RECT 354.860 -40.220 356.820 -39.940 ;
        RECT 354.860 -43.070 355.140 -40.220 ;
        RECT 356.540 -40.270 356.820 -40.220 ;
        RECT 359.340 -40.830 359.620 -36.860 ;
        RECT 361.020 -36.860 362.980 -36.580 ;
        RECT 361.020 -36.910 361.300 -36.860 ;
        RECT 362.700 -36.910 362.980 -36.860 ;
        RECT 364.940 -38.590 365.220 -34.850 ;
        RECT 367.180 -34.900 367.460 -34.850 ;
        RECT 366.620 -35.180 367.460 -34.900 ;
        RECT 366.620 -35.790 366.900 -35.180 ;
        RECT 367.180 -35.230 367.460 -35.180 ;
        RECT 368.860 -35.790 369.140 -32.940 ;
        RECT 369.420 -32.990 369.700 -32.940 ;
        RECT 369.420 -39.710 369.700 -38.210 ;
        RECT 369.980 -39.380 370.260 -34.850 ;
        RECT 371.660 -35.230 371.940 -23.140 ;
        RECT 372.220 -32.570 372.500 -20.290 ;
        RECT 375.580 -22.860 375.860 -7.970 ;
        RECT 376.140 -15.070 376.420 -3.490 ;
        RECT 377.260 -9.610 377.540 -9.090 ;
        RECT 379.500 -12.410 379.780 -11.890 ;
        RECT 377.820 -15.210 378.100 -14.690 ;
        RECT 378.940 -16.980 379.220 -16.370 ;
        RECT 377.820 -17.260 379.220 -16.980 ;
        RECT 376.700 -19.550 376.980 -18.610 ;
        RECT 376.140 -20.810 376.420 -20.290 ;
        RECT 374.460 -23.140 375.860 -22.860 ;
        RECT 372.780 -24.170 373.060 -23.650 ;
        RECT 374.460 -24.030 374.740 -23.140 ;
        RECT 377.820 -26.830 378.100 -17.260 ;
        RECT 380.060 -22.860 380.340 -11.330 ;
        RECT 381.180 -12.970 381.460 -12.450 ;
        RECT 380.620 -16.330 380.900 -15.810 ;
        RECT 380.060 -23.140 380.900 -22.860 ;
        RECT 380.620 -24.030 380.900 -23.140 ;
        RECT 376.140 -30.750 376.420 -27.010 ;
        RECT 373.900 -34.670 374.180 -32.050 ;
        RECT 377.820 -34.340 378.100 -34.290 ;
        RECT 376.700 -34.620 378.100 -34.340 ;
        RECT 372.780 -35.930 373.060 -35.410 ;
        RECT 372.220 -38.260 372.500 -38.210 ;
        RECT 372.220 -38.540 373.060 -38.260 ;
        RECT 372.220 -38.590 372.500 -38.540 ;
        RECT 372.220 -39.380 372.500 -39.330 ;
        RECT 369.980 -39.660 372.500 -39.380 ;
        RECT 372.220 -39.710 372.500 -39.660 ;
        RECT 357.660 -42.510 357.940 -41.570 ;
        RECT 369.980 -43.630 370.260 -40.450 ;
        RECT 372.780 -43.630 373.060 -38.540 ;
        RECT 376.700 -43.070 376.980 -34.620 ;
        RECT 377.820 -34.810 378.100 -34.620 ;
        RECT 381.740 -34.670 382.020 6.260 ;
        RECT 382.300 -0.510 382.580 2.670 ;
        RECT 382.860 -1.300 383.140 -1.250 ;
        RECT 384.540 -1.300 384.820 -1.250 ;
        RECT 382.860 -1.580 384.820 -1.300 ;
        RECT 382.860 -1.630 383.140 -1.580 ;
        RECT 384.540 -1.770 384.820 -1.580 ;
        RECT 383.980 -4.430 384.260 -3.910 ;
        RECT 386.220 -4.430 386.500 6.260 ;
        RECT 386.780 6.210 387.060 6.260 ;
        RECT 386.780 2.290 387.060 3.790 ;
        RECT 382.300 -8.910 382.580 -5.170 ;
        RECT 383.420 -13.950 383.700 -11.890 ;
        RECT 383.980 -11.940 384.260 -5.170 ;
        RECT 384.540 -11.940 384.820 -11.890 ;
        RECT 383.980 -12.220 384.820 -11.940 ;
        RECT 384.540 -12.270 384.820 -12.220 ;
        RECT 382.300 -16.420 382.580 -16.370 ;
        RECT 382.300 -16.700 383.140 -16.420 ;
        RECT 382.300 -16.890 382.580 -16.700 ;
        RECT 382.860 -19.550 383.140 -16.700 ;
        RECT 383.980 -26.270 384.260 -13.010 ;
        RECT 385.100 -14.510 385.380 -7.970 ;
        RECT 387.340 -8.350 387.620 -0.690 ;
        RECT 387.900 -3.540 388.180 -1.250 ;
        RECT 388.460 -2.190 388.740 4.350 ;
        RECT 388.460 -3.540 388.740 -3.490 ;
        RECT 387.900 -3.820 388.740 -3.540 ;
        RECT 388.460 -3.870 388.740 -3.820 ;
        RECT 387.900 -8.350 388.180 -4.610 ;
        RECT 384.540 -16.190 384.820 -14.690 ;
        RECT 385.100 -20.250 385.380 -17.490 ;
        RECT 385.660 -26.830 385.940 -20.290 ;
        RECT 386.780 -27.390 387.060 -24.770 ;
        RECT 383.980 -30.190 384.260 -28.130 ;
        RECT 380.060 -35.370 380.340 -34.850 ;
        RECT 382.300 -35.790 382.580 -34.850 ;
        RECT 380.060 -43.630 380.340 -38.210 ;
        RECT 382.300 -42.510 382.580 -36.530 ;
        RECT 383.980 -40.970 384.260 -35.970 ;
        RECT 385.100 -38.590 385.380 -32.610 ;
        RECT 386.220 -36.350 386.500 -27.570 ;
        RECT 386.780 -30.420 387.060 -30.370 ;
        RECT 387.340 -30.420 387.620 -24.770 ;
        RECT 387.900 -30.190 388.180 -24.770 ;
        RECT 386.780 -30.700 387.620 -30.420 ;
        RECT 386.780 -30.750 387.060 -30.700 ;
        RECT 386.780 -34.340 387.060 -32.610 ;
        RECT 389.020 -34.340 389.300 11.300 ;
        RECT 389.580 11.110 389.860 11.300 ;
        RECT 391.820 7.890 392.100 11.630 ;
        RECT 393.500 11.250 393.780 27.310 ;
        RECT 396.300 15.030 396.580 15.550 ;
        RECT 400.220 15.500 400.500 16.670 ;
        RECT 401.900 16.060 402.180 16.110 ;
        RECT 401.900 15.780 403.860 16.060 ;
        RECT 401.900 15.730 402.180 15.780 ;
        RECT 400.220 15.220 401.060 15.500 ;
        RECT 400.220 15.170 400.500 15.220 ;
        RECT 399.100 14.470 399.380 14.990 ;
        RECT 397.420 13.910 397.700 14.430 ;
        RECT 400.780 12.700 401.060 15.220 ;
        RECT 401.340 13.260 401.620 14.430 ;
        RECT 401.900 14.380 402.180 14.430 ;
        RECT 401.900 14.100 403.300 14.380 ;
        RECT 401.900 13.910 402.180 14.100 ;
        RECT 401.340 12.980 402.740 13.260 ;
        RECT 400.780 12.420 402.180 12.700 ;
        RECT 401.340 7.330 401.620 11.070 ;
        RECT 401.900 7.330 402.180 12.420 ;
        RECT 402.460 10.690 402.740 12.980 ;
        RECT 403.020 11.020 403.300 14.100 ;
        RECT 403.580 11.810 403.860 15.780 ;
        RECT 404.140 14.940 404.420 19.470 ;
        RECT 404.700 16.290 404.980 35.660 ;
        RECT 410.300 34.540 410.580 34.590 ;
        RECT 411.980 34.540 412.260 46.910 ;
        RECT 412.540 35.890 412.820 41.870 ;
        RECT 410.300 34.260 412.260 34.540 ;
        RECT 408.620 30.290 408.900 34.030 ;
        RECT 409.180 31.410 409.460 32.350 ;
        RECT 409.180 26.700 409.460 26.750 ;
        RECT 410.300 26.700 410.580 34.260 ;
        RECT 411.420 31.740 411.700 31.790 ;
        RECT 413.100 31.740 413.380 45.790 ;
        RECT 422.060 43.730 422.340 46.350 ;
        RECT 426.540 45.830 426.820 46.350 ;
        RECT 415.340 38.130 415.620 42.990 ;
        RECT 416.460 41.490 416.740 42.990 ;
        RECT 417.580 41.910 417.860 42.430 ;
        RECT 417.020 34.770 417.300 39.070 ;
        RECT 418.700 38.460 418.980 42.990 ;
        RECT 419.820 38.690 420.100 42.990 ;
        RECT 417.580 38.180 418.980 38.460 ;
        RECT 415.340 33.980 415.620 34.030 ;
        RECT 411.420 31.460 413.380 31.740 ;
        RECT 413.660 33.700 415.620 33.980 ;
        RECT 411.420 31.410 411.700 31.460 ;
        RECT 411.420 26.790 411.700 27.310 ;
        RECT 409.180 26.420 410.580 26.700 ;
        RECT 407.500 19.650 407.780 21.710 ;
        RECT 404.140 14.660 405.540 14.940 ;
        RECT 404.140 12.370 404.420 13.310 ;
        RECT 405.260 12.700 405.540 14.660 ;
        RECT 406.940 12.930 407.220 15.550 ;
        RECT 405.820 12.700 406.100 12.750 ;
        RECT 405.260 12.420 406.100 12.700 ;
        RECT 405.820 12.370 406.100 12.420 ;
        RECT 403.020 10.740 404.420 11.020 ;
        RECT 403.580 7.330 403.860 8.270 ;
        RECT 404.140 7.330 404.420 10.740 ;
        RECT 407.500 10.130 407.780 11.630 ;
        RECT 409.180 9.900 409.460 26.420 ;
        RECT 409.740 11.020 410.020 11.070 ;
        RECT 409.740 10.740 410.580 11.020 ;
        RECT 409.740 10.690 410.020 10.740 ;
        RECT 410.300 10.130 410.580 10.740 ;
        RECT 409.180 9.620 410.020 9.900 ;
        RECT 406.940 7.190 407.220 7.710 ;
        RECT 391.260 6.070 391.540 6.590 ;
        RECT 392.380 3.410 392.660 7.150 ;
        RECT 407.500 6.630 407.780 7.150 ;
        RECT 396.300 6.070 396.580 6.590 ;
        RECT 403.020 6.070 403.300 6.590 ;
        RECT 397.980 4.860 398.260 4.910 ;
        RECT 397.980 4.580 398.820 4.860 ;
        RECT 397.980 4.530 398.260 4.580 ;
        RECT 394.620 3.740 394.900 3.790 ;
        RECT 392.940 3.460 394.900 3.740 ;
        RECT 391.820 0.610 392.100 3.230 ;
        RECT 392.940 0.050 393.220 3.460 ;
        RECT 394.620 3.270 394.900 3.460 ;
        RECT 396.860 -0.180 397.140 -0.130 ;
        RECT 396.300 -0.460 397.140 -0.180 ;
        RECT 395.740 -0.740 396.020 -0.690 ;
        RECT 394.620 -1.020 396.020 -0.740 ;
        RECT 390.140 -4.990 390.420 -1.250 ;
        RECT 394.620 -4.570 394.900 -1.020 ;
        RECT 395.740 -1.070 396.020 -1.020 ;
        RECT 389.580 -7.930 389.860 -7.410 ;
        RECT 391.260 -8.910 391.540 -5.730 ;
        RECT 390.140 -21.230 390.420 -15.810 ;
        RECT 390.700 -16.750 390.980 -11.890 ;
        RECT 391.820 -12.500 392.100 -7.970 ;
        RECT 396.300 -8.350 396.580 -0.460 ;
        RECT 396.860 -0.510 397.140 -0.460 ;
        RECT 395.740 -9.140 396.020 -8.530 ;
        RECT 396.300 -9.140 396.580 -9.090 ;
        RECT 395.740 -9.420 396.580 -9.140 ;
        RECT 396.300 -9.610 396.580 -9.420 ;
        RECT 396.300 -11.380 396.580 -11.330 ;
        RECT 396.860 -11.380 397.140 -1.250 ;
        RECT 397.980 -4.100 398.260 3.790 ;
        RECT 398.540 0.050 398.820 4.580 ;
        RECT 400.220 4.300 400.500 4.350 ;
        RECT 400.220 4.020 401.620 4.300 ;
        RECT 400.220 3.830 400.500 4.020 ;
        RECT 401.340 0.050 401.620 4.020 ;
        RECT 406.380 3.410 406.660 6.590 ;
        RECT 409.180 1.170 409.460 7.710 ;
        RECT 399.660 -0.650 399.940 -0.130 ;
        RECT 400.780 -4.100 401.060 -4.050 ;
        RECT 397.980 -4.380 401.060 -4.100 ;
        RECT 402.460 -4.100 402.740 -0.690 ;
        RECT 404.700 -2.980 404.980 -1.250 ;
        RECT 404.700 -3.260 406.660 -2.980 ;
        RECT 404.700 -3.310 404.980 -3.260 ;
        RECT 403.580 -4.100 403.860 -4.050 ;
        RECT 402.460 -4.380 403.860 -4.100 ;
        RECT 396.300 -11.660 397.140 -11.380 ;
        RECT 396.300 -11.710 396.580 -11.660 ;
        RECT 397.420 -11.940 397.700 -4.610 ;
        RECT 400.780 -4.660 401.060 -4.380 ;
        RECT 400.780 -4.940 401.620 -4.660 ;
        RECT 399.660 -8.350 399.940 -6.850 ;
        RECT 401.340 -8.350 401.620 -4.940 ;
        RECT 401.900 -5.220 402.180 -5.170 ;
        RECT 401.900 -5.500 402.740 -5.220 ;
        RECT 401.900 -5.550 402.180 -5.500 ;
        RECT 398.540 -11.940 398.820 -11.890 ;
        RECT 397.420 -12.220 398.820 -11.940 ;
        RECT 398.540 -12.270 398.820 -12.220 ;
        RECT 391.260 -12.780 392.100 -12.500 ;
        RECT 390.700 -21.230 390.980 -20.290 ;
        RECT 391.260 -20.670 391.540 -12.780 ;
        RECT 392.380 -12.970 392.660 -12.450 ;
        RECT 400.780 -13.390 401.060 -11.890 ;
        RECT 392.940 -16.330 393.220 -15.810 ;
        RECT 391.820 -18.990 392.100 -16.930 ;
        RECT 391.820 -20.250 392.100 -19.730 ;
        RECT 392.380 -19.780 392.660 -16.930 ;
        RECT 395.740 -17.540 396.020 -14.130 ;
        RECT 397.980 -17.310 398.260 -14.690 ;
        RECT 401.900 -16.190 402.180 -6.290 ;
        RECT 395.740 -17.820 396.580 -17.540 ;
        RECT 394.620 -19.780 394.900 -19.730 ;
        RECT 392.380 -20.060 394.900 -19.780 ;
        RECT 394.620 -20.110 394.900 -20.060 ;
        RECT 390.700 -24.170 390.980 -23.650 ;
        RECT 389.580 -31.870 389.860 -24.210 ;
        RECT 392.380 -25.290 392.660 -24.770 ;
        RECT 395.180 -27.390 395.460 -20.850 ;
        RECT 395.740 -24.590 396.020 -20.850 ;
        RECT 395.740 -26.500 396.020 -26.450 ;
        RECT 396.300 -26.500 396.580 -17.820 ;
        RECT 401.900 -21.790 402.180 -20.290 ;
        RECT 402.460 -21.230 402.740 -5.500 ;
        RECT 403.580 -6.670 403.860 -4.380 ;
        RECT 406.380 -4.430 406.660 -3.260 ;
        RECT 403.580 -11.710 403.860 -7.410 ;
        RECT 404.140 -9.050 404.420 -8.530 ;
        RECT 403.580 -14.180 403.860 -14.130 ;
        RECT 403.580 -14.460 404.420 -14.180 ;
        RECT 403.580 -14.510 403.860 -14.460 ;
        RECT 404.140 -16.190 404.420 -14.460 ;
        RECT 403.020 -16.890 403.300 -16.370 ;
        RECT 404.700 -16.750 404.980 -7.970 ;
        RECT 406.380 -17.870 406.660 -9.090 ;
        RECT 406.940 -12.270 407.220 -7.970 ;
        RECT 407.500 -16.420 407.780 -1.810 ;
        RECT 408.620 -2.980 408.900 -0.130 ;
        RECT 409.180 -2.190 409.460 -1.250 ;
        RECT 409.180 -2.980 409.460 -2.930 ;
        RECT 408.620 -3.260 409.460 -2.980 ;
        RECT 409.180 -3.310 409.460 -3.260 ;
        RECT 408.620 -9.050 408.900 -8.530 ;
        RECT 408.620 -16.420 408.900 -16.370 ;
        RECT 407.500 -16.700 408.900 -16.420 ;
        RECT 408.620 -16.890 408.900 -16.700 ;
        RECT 403.580 -22.860 403.860 -19.170 ;
        RECT 409.740 -22.860 410.020 9.620 ;
        RECT 410.300 7.100 410.580 7.150 ;
        RECT 411.420 7.100 411.700 7.710 ;
        RECT 410.300 6.820 411.700 7.100 ;
        RECT 410.300 6.770 410.580 6.820 ;
        RECT 411.980 6.540 412.260 31.460 ;
        RECT 413.660 30.850 413.940 33.700 ;
        RECT 415.340 33.650 415.620 33.700 ;
        RECT 415.900 30.850 416.180 32.350 ;
        RECT 417.580 30.290 417.860 38.180 ;
        RECT 420.940 37.900 421.220 42.990 ;
        RECT 418.140 37.620 421.220 37.900 ;
        RECT 418.140 33.650 418.420 37.620 ;
        RECT 422.060 34.770 422.340 35.710 ;
        RECT 415.340 26.370 415.620 27.310 ;
        RECT 417.020 26.790 417.300 27.310 ;
        RECT 420.380 26.790 420.660 27.310 ;
        RECT 418.140 22.450 418.420 26.750 ;
        RECT 421.500 26.370 421.780 27.310 ;
        RECT 423.180 26.930 423.460 42.990 ;
        RECT 424.860 26.930 425.140 41.870 ;
        RECT 427.100 41.490 427.380 45.790 ;
        RECT 427.100 39.110 427.380 39.630 ;
        RECT 427.100 31.830 427.380 32.350 ;
        RECT 422.060 26.700 422.340 26.750 ;
        RECT 422.060 26.420 422.900 26.700 ;
        RECT 422.060 26.370 422.340 26.420 ;
        RECT 419.820 23.340 420.100 23.390 ;
        RECT 422.060 23.340 422.340 23.390 ;
        RECT 419.260 23.060 422.340 23.340 ;
        RECT 418.700 21.330 418.980 22.270 ;
        RECT 416.460 20.540 416.740 20.590 ;
        RECT 419.260 20.540 419.540 23.060 ;
        RECT 419.820 23.010 420.100 23.060 ;
        RECT 422.060 23.010 422.340 23.060 ;
        RECT 416.460 20.260 419.540 20.540 ;
        RECT 416.460 20.210 416.740 20.260 ;
        RECT 411.420 6.260 412.260 6.540 ;
        RECT 410.860 -14.510 411.140 -13.010 ;
        RECT 410.860 -20.810 411.140 -20.290 ;
        RECT 410.300 -21.790 410.580 -20.850 ;
        RECT 403.580 -23.140 407.220 -22.860 ;
        RECT 395.740 -26.780 396.580 -26.500 ;
        RECT 395.740 -26.830 396.020 -26.780 ;
        RECT 396.860 -28.090 397.140 -27.570 ;
        RECT 399.660 -29.070 399.940 -23.650 ;
        RECT 401.900 -26.500 402.180 -26.450 ;
        RECT 402.460 -26.500 402.740 -23.650 ;
        RECT 401.900 -26.780 402.740 -26.500 ;
        RECT 401.900 -26.830 402.180 -26.780 ;
        RECT 405.820 -27.390 406.100 -23.140 ;
        RECT 406.940 -23.470 407.220 -23.140 ;
        RECT 409.180 -23.140 410.020 -22.860 ;
        RECT 400.220 -27.620 400.500 -27.570 ;
        RECT 402.460 -27.620 402.740 -27.570 ;
        RECT 403.580 -27.620 403.860 -27.570 ;
        RECT 405.260 -27.620 405.540 -27.570 ;
        RECT 400.220 -27.900 402.180 -27.620 ;
        RECT 400.220 -28.090 400.500 -27.900 ;
        RECT 389.580 -34.340 389.860 -34.290 ;
        RECT 386.780 -34.620 387.620 -34.340 ;
        RECT 386.780 -34.670 387.060 -34.620 ;
        RECT 387.340 -38.260 387.620 -34.620 ;
        RECT 389.020 -34.620 389.860 -34.340 ;
        RECT 389.020 -35.230 389.300 -34.620 ;
        RECT 389.580 -34.670 389.860 -34.620 ;
        RECT 387.900 -37.050 388.180 -36.530 ;
        RECT 390.140 -36.910 390.420 -32.050 ;
        RECT 387.900 -38.260 388.180 -38.210 ;
        RECT 387.340 -38.540 388.180 -38.260 ;
        RECT 387.900 -38.590 388.180 -38.540 ;
        RECT 386.220 -42.650 386.500 -42.130 ;
        RECT 381.180 -43.210 381.460 -42.690 ;
        RECT 390.700 -42.740 390.980 -35.410 ;
        RECT 391.260 -39.150 391.540 -35.410 ;
        RECT 389.020 -43.020 390.980 -42.740 ;
        RECT 400.780 -39.380 401.060 -39.330 ;
        RECT 401.340 -39.380 401.620 -28.690 ;
        RECT 401.900 -31.870 402.180 -27.900 ;
        RECT 402.460 -27.900 403.300 -27.620 ;
        RECT 402.460 -27.950 402.740 -27.900 ;
        RECT 403.020 -31.540 403.300 -27.900 ;
        RECT 403.580 -27.900 405.540 -27.620 ;
        RECT 403.580 -27.950 403.860 -27.900 ;
        RECT 405.260 -27.950 405.540 -27.900 ;
        RECT 403.580 -31.540 403.860 -31.490 ;
        RECT 403.020 -31.820 403.860 -31.540 ;
        RECT 403.580 -31.870 403.860 -31.820 ;
        RECT 405.260 -32.570 405.540 -32.050 ;
        RECT 400.780 -39.660 401.620 -39.380 ;
        RECT 352.620 -46.940 355.140 -46.660 ;
        RECT 352.620 -46.990 352.900 -46.940 ;
        RECT 354.860 -47.550 355.140 -46.940 ;
        RECT 359.900 -47.130 360.180 -46.610 ;
        RECT 376.140 -47.550 376.420 -44.370 ;
        RECT 369.980 -61.000 370.260 -47.730 ;
        RECT 381.740 -48.250 382.020 -47.730 ;
        RECT 387.900 -61.000 388.180 -46.610 ;
        RECT 389.020 -46.990 389.300 -43.020 ;
        RECT 397.420 -43.770 397.700 -43.250 ;
        RECT 400.780 -43.630 401.060 -39.660 ;
        RECT 403.020 -39.710 403.300 -32.610 ;
        RECT 402.460 -42.650 402.740 -40.450 ;
        RECT 409.180 -42.180 409.460 -23.140 ;
        RECT 411.420 -35.790 411.700 6.260 ;
        RECT 412.540 -1.210 412.820 -0.690 ;
        RECT 411.980 -1.770 412.260 -1.250 ;
        RECT 411.980 -8.910 412.260 -4.050 ;
        RECT 414.220 -7.460 414.500 -7.410 ;
        RECT 415.340 -7.460 415.620 19.470 ;
        RECT 422.620 18.530 422.900 26.420 ;
        RECT 427.100 23.010 427.380 23.950 ;
        RECT 423.740 20.540 424.020 22.270 ;
        RECT 428.220 21.660 428.500 46.910 ;
        RECT 428.780 31.410 429.060 43.550 ;
        RECT 431.580 35.890 431.860 39.070 ;
        RECT 434.940 38.690 435.220 40.190 ;
        RECT 436.060 38.690 436.340 43.550 ;
        RECT 437.180 39.580 437.460 39.630 ;
        RECT 439.420 39.580 439.700 39.630 ;
        RECT 437.180 39.300 439.700 39.580 ;
        RECT 437.180 39.250 437.460 39.300 ;
        RECT 439.420 39.250 439.700 39.300 ;
        RECT 439.980 39.250 440.260 42.990 ;
        RECT 442.780 39.250 443.060 49.380 ;
        RECT 443.900 45.740 444.180 46.910 ;
        RECT 446.140 45.740 446.420 45.790 ;
        RECT 443.900 45.460 446.420 45.740 ;
        RECT 441.100 38.550 441.380 39.070 ;
        RECT 437.740 37.990 438.020 38.510 ;
        RECT 433.820 35.190 434.100 35.710 ;
        RECT 431.580 30.290 431.860 31.230 ;
        RECT 427.100 21.380 428.500 21.660 ;
        RECT 427.100 20.540 427.380 21.380 ;
        RECT 423.740 20.260 427.380 20.540 ;
        RECT 427.100 20.210 427.380 20.260 ;
        RECT 425.980 18.390 426.260 18.910 ;
        RECT 427.660 18.530 427.940 20.590 ;
        RECT 417.020 -5.220 417.300 18.350 ;
        RECT 428.780 17.740 429.060 23.390 ;
        RECT 429.340 22.220 429.620 22.270 ;
        RECT 429.340 21.940 430.180 22.220 ;
        RECT 429.340 21.890 429.620 21.940 ;
        RECT 429.900 20.210 430.180 21.940 ;
        RECT 432.140 21.750 432.420 22.270 ;
        RECT 434.380 21.330 434.660 30.110 ;
        RECT 437.740 30.060 438.020 35.710 ;
        RECT 438.300 30.060 438.580 30.110 ;
        RECT 437.740 29.780 438.580 30.060 ;
        RECT 438.300 29.590 438.580 29.780 ;
        RECT 438.860 26.930 439.140 37.950 ;
        RECT 442.220 37.430 442.500 37.950 ;
        RECT 434.940 21.750 435.220 22.270 ;
        RECT 435.500 21.100 435.780 26.190 ;
        RECT 438.860 24.460 439.140 24.510 ;
        RECT 434.940 20.820 435.780 21.100 ;
        RECT 436.060 24.180 439.140 24.460 ;
        RECT 434.940 20.210 435.220 20.820 ;
        RECT 432.700 19.510 432.980 20.030 ;
        RECT 431.580 18.530 431.860 19.470 ;
        RECT 425.420 17.460 429.060 17.740 ;
        RECT 419.820 14.050 420.100 15.550 ;
        RECT 423.740 15.030 424.020 15.550 ;
        RECT 422.620 10.690 422.900 14.430 ;
        RECT 423.180 6.630 423.460 7.150 ;
        RECT 418.140 -0.740 418.420 -0.690 ;
        RECT 418.140 -1.020 418.980 -0.740 ;
        RECT 418.140 -1.070 418.420 -1.020 ;
        RECT 417.580 -5.220 417.860 -5.170 ;
        RECT 417.020 -5.500 417.860 -5.220 ;
        RECT 417.580 -5.550 417.860 -5.500 ;
        RECT 414.220 -7.740 415.620 -7.460 ;
        RECT 414.220 -7.930 414.500 -7.740 ;
        RECT 411.980 -11.850 412.260 -11.330 ;
        RECT 417.020 -11.850 417.300 -11.330 ;
        RECT 412.540 -12.830 412.820 -11.890 ;
        RECT 415.340 -16.190 415.620 -12.450 ;
        RECT 417.020 -15.630 417.300 -14.690 ;
        RECT 414.780 -16.890 415.060 -16.370 ;
        RECT 411.980 -20.250 412.260 -19.730 ;
        RECT 418.140 -20.810 418.420 -3.490 ;
        RECT 418.700 -20.110 418.980 -1.020 ;
        RECT 419.820 -7.790 420.100 -4.050 ;
        RECT 423.740 -4.570 424.020 -4.050 ;
        RECT 424.860 -4.100 425.140 -0.690 ;
        RECT 424.300 -4.380 425.140 -4.100 ;
        RECT 424.300 -5.780 424.580 -4.380 ;
        RECT 424.860 -4.430 425.140 -4.380 ;
        RECT 423.180 -6.060 424.580 -5.780 ;
        RECT 422.620 -8.490 422.900 -7.970 ;
        RECT 419.260 -18.660 419.540 -12.450 ;
        RECT 421.500 -15.300 421.780 -15.250 ;
        RECT 421.500 -15.580 422.340 -15.300 ;
        RECT 421.500 -15.630 421.780 -15.580 ;
        RECT 420.940 -16.330 421.220 -15.810 ;
        RECT 419.260 -18.940 420.100 -18.660 ;
        RECT 419.820 -20.110 420.100 -18.940 ;
        RECT 412.540 -24.030 412.820 -20.850 ;
        RECT 421.500 -21.370 421.780 -20.850 ;
        RECT 422.060 -22.860 422.340 -15.580 ;
        RECT 422.620 -15.860 422.900 -15.810 ;
        RECT 423.180 -15.860 423.460 -6.060 ;
        RECT 424.300 -11.710 424.580 -7.970 ;
        RECT 425.420 -11.940 425.700 17.460 ;
        RECT 426.540 14.380 426.820 14.430 ;
        RECT 426.540 14.100 427.940 14.380 ;
        RECT 426.540 14.050 426.820 14.100 ;
        RECT 426.540 12.230 426.820 12.750 ;
        RECT 427.660 7.100 427.940 14.100 ;
        RECT 428.220 12.370 428.500 14.430 ;
        RECT 429.900 13.910 430.180 14.430 ;
        RECT 432.700 12.370 432.980 13.310 ;
        RECT 433.820 12.140 434.100 15.550 ;
        RECT 434.380 14.940 434.660 19.470 ;
        RECT 435.500 19.090 435.780 20.030 ;
        RECT 436.060 18.300 436.340 24.180 ;
        RECT 438.860 24.130 439.140 24.180 ;
        RECT 435.500 18.020 436.340 18.300 ;
        RECT 435.500 15.730 435.780 18.020 ;
        RECT 436.060 15.030 436.340 15.550 ;
        RECT 434.940 14.940 435.220 14.990 ;
        RECT 434.380 14.660 435.220 14.940 ;
        RECT 434.380 12.140 434.660 12.190 ;
        RECT 433.820 11.860 434.660 12.140 ;
        RECT 434.380 11.810 434.660 11.860 ;
        RECT 427.660 6.820 429.060 7.100 ;
        RECT 427.100 6.540 427.380 6.590 ;
        RECT 427.100 6.260 428.500 6.540 ;
        RECT 427.100 6.070 427.380 6.260 ;
        RECT 426.540 4.390 426.820 4.910 ;
        RECT 428.220 3.410 428.500 6.260 ;
        RECT 428.780 -2.980 429.060 6.820 ;
        RECT 432.140 3.830 432.420 4.350 ;
        RECT 429.340 3.180 429.620 3.230 ;
        RECT 431.580 3.180 431.860 3.790 ;
        RECT 429.340 2.900 431.860 3.180 ;
        RECT 429.340 2.850 429.620 2.900 ;
        RECT 428.780 -3.260 429.620 -2.980 ;
        RECT 427.100 -8.020 427.380 -7.970 ;
        RECT 425.980 -8.300 427.380 -8.020 ;
        RECT 425.980 -11.150 426.260 -8.300 ;
        RECT 427.100 -8.490 427.380 -8.300 ;
        RECT 428.780 -11.150 429.060 -8.530 ;
        RECT 429.340 -11.710 429.620 -3.260 ;
        RECT 425.420 -12.220 426.260 -11.940 ;
        RECT 422.620 -16.140 423.460 -15.860 ;
        RECT 422.620 -16.190 422.900 -16.140 ;
        RECT 423.180 -20.900 423.460 -16.140 ;
        RECT 418.140 -23.610 418.420 -23.090 ;
        RECT 421.500 -23.140 422.340 -22.860 ;
        RECT 422.620 -21.180 423.460 -20.900 ;
        RECT 418.700 -24.170 418.980 -23.650 ;
        RECT 420.380 -23.700 420.660 -23.650 ;
        RECT 419.820 -23.980 420.660 -23.700 ;
        RECT 413.100 -27.950 413.380 -25.330 ;
        RECT 415.340 -29.300 415.620 -24.770 ;
        RECT 418.140 -24.820 418.420 -24.210 ;
        RECT 419.820 -24.820 420.100 -23.980 ;
        RECT 420.380 -24.030 420.660 -23.980 ;
        RECT 421.500 -24.030 421.780 -23.140 ;
        RECT 418.140 -25.100 420.100 -24.820 ;
        RECT 418.140 -26.830 418.420 -25.100 ;
        RECT 420.380 -25.150 420.660 -24.630 ;
        RECT 421.500 -24.820 421.780 -24.770 ;
        RECT 421.500 -25.100 422.340 -24.820 ;
        RECT 421.500 -25.150 421.780 -25.100 ;
        RECT 422.060 -27.060 422.340 -25.100 ;
        RECT 421.500 -27.340 422.340 -27.060 ;
        RECT 419.820 -29.300 420.100 -28.130 ;
        RECT 414.780 -29.580 415.620 -29.300 ;
        RECT 414.780 -40.970 415.060 -29.580 ;
        RECT 415.340 -29.630 415.620 -29.580 ;
        RECT 418.700 -29.580 420.100 -29.300 ;
        RECT 418.700 -34.670 418.980 -29.580 ;
        RECT 419.820 -29.630 420.100 -29.580 ;
        RECT 421.500 -31.870 421.780 -27.340 ;
        RECT 422.060 -27.530 422.340 -27.340 ;
        RECT 422.060 -32.570 422.340 -32.050 ;
        RECT 422.620 -36.910 422.900 -21.180 ;
        RECT 423.740 -21.460 424.020 -15.810 ;
        RECT 425.420 -19.690 425.700 -19.170 ;
        RECT 423.180 -21.740 424.020 -21.460 ;
        RECT 423.180 -26.830 423.460 -21.740 ;
        RECT 423.740 -22.860 424.020 -22.530 ;
        RECT 425.980 -22.860 426.260 -12.220 ;
        RECT 430.460 -12.270 430.740 -9.090 ;
        RECT 431.580 -10.590 431.860 2.900 ;
        RECT 432.700 -6.670 432.980 10.510 ;
        RECT 433.820 7.890 434.100 11.070 ;
        RECT 434.380 7.660 434.660 7.710 ;
        RECT 434.940 7.660 435.220 14.660 ;
        RECT 435.500 11.250 435.780 14.990 ;
        RECT 436.620 9.340 436.900 23.390 ;
        RECT 440.540 22.870 440.820 23.390 ;
        RECT 437.180 19.510 437.460 20.030 ;
        RECT 438.860 19.090 439.140 21.710 ;
        RECT 439.420 16.290 439.700 22.270 ;
        RECT 442.220 19.650 442.500 22.270 ;
        RECT 437.740 14.470 438.020 14.990 ;
        RECT 438.860 11.250 439.140 13.310 ;
        RECT 437.180 10.460 437.460 10.510 ;
        RECT 437.180 10.180 439.700 10.460 ;
        RECT 437.180 10.130 437.460 10.180 ;
        RECT 434.380 7.380 435.220 7.660 ;
        RECT 436.060 9.060 436.900 9.340 ;
        RECT 434.380 3.410 434.660 7.380 ;
        RECT 435.500 3.970 435.780 6.590 ;
        RECT 436.060 4.860 436.340 9.060 ;
        RECT 436.620 5.980 436.900 8.270 ;
        RECT 439.420 7.330 439.700 10.180 ;
        RECT 437.740 7.100 438.020 7.150 ;
        RECT 437.740 6.820 438.580 7.100 ;
        RECT 437.740 6.770 438.020 6.820 ;
        RECT 436.620 5.700 438.020 5.980 ;
        RECT 436.620 4.860 436.900 4.910 ;
        RECT 436.060 4.580 436.900 4.860 ;
        RECT 433.260 1.500 433.540 3.230 ;
        RECT 433.260 1.220 435.220 1.500 ;
        RECT 434.940 0.610 435.220 1.220 ;
        RECT 435.500 -3.310 435.780 1.550 ;
        RECT 436.060 -1.070 436.340 4.580 ;
        RECT 436.620 4.530 436.900 4.580 ;
        RECT 437.180 0.610 437.460 2.670 ;
        RECT 436.620 -7.230 436.900 0.430 ;
        RECT 437.740 0.380 438.020 5.700 ;
        RECT 438.300 1.500 438.580 6.820 ;
        RECT 439.980 3.410 440.260 14.990 ;
        RECT 442.220 14.470 442.500 14.990 ;
        RECT 442.780 10.740 443.060 36.270 ;
        RECT 443.340 30.850 443.620 42.990 ;
        RECT 443.340 23.900 443.620 23.950 ;
        RECT 443.900 23.900 444.180 45.460 ;
        RECT 446.140 45.410 446.420 45.460 ;
        RECT 444.460 41.910 444.740 42.430 ;
        RECT 445.580 38.690 445.860 43.550 ;
        RECT 446.140 40.140 446.420 41.870 ;
        RECT 446.140 39.860 446.980 40.140 ;
        RECT 446.700 39.580 446.980 39.860 ;
        RECT 446.700 39.300 448.100 39.580 ;
        RECT 443.340 23.620 444.180 23.900 ;
        RECT 443.340 23.570 443.620 23.620 ;
        RECT 446.140 21.750 446.420 37.950 ;
        RECT 447.820 35.100 448.100 39.300 ;
        RECT 448.380 35.890 448.660 42.430 ;
        RECT 457.340 38.690 457.620 41.870 ;
        RECT 459.580 40.140 459.860 61.000 ;
        RECT 459.020 39.860 459.860 40.140 ;
        RECT 448.940 35.100 449.220 35.150 ;
        RECT 447.820 34.820 449.220 35.100 ;
        RECT 448.940 34.770 449.220 34.820 ;
        RECT 452.300 35.100 452.580 35.150 ;
        RECT 452.300 34.820 453.140 35.100 ;
        RECT 452.300 34.770 452.580 34.820 ;
        RECT 449.500 20.210 449.780 31.230 ;
        RECT 452.860 30.060 453.140 34.820 ;
        RECT 455.100 30.710 455.380 31.230 ;
        RECT 453.980 30.060 454.260 30.110 ;
        RECT 452.860 29.780 454.260 30.060 ;
        RECT 453.980 29.590 454.260 29.780 ;
        RECT 455.660 27.820 455.940 34.590 ;
        RECT 459.020 31.970 459.300 39.860 ;
        RECT 457.900 28.050 458.180 31.230 ;
        RECT 458.460 29.170 458.740 31.790 ;
        RECT 455.100 27.540 455.940 27.820 ;
        RECT 454.540 25.670 454.820 26.190 ;
        RECT 446.140 10.740 446.420 14.430 ;
        RECT 447.260 10.740 447.540 11.070 ;
        RECT 442.780 10.460 443.620 10.740 ;
        RECT 442.220 6.540 442.500 7.710 ;
        RECT 443.340 6.540 443.620 10.460 ;
        RECT 446.140 10.460 447.540 10.740 ;
        RECT 442.220 6.260 444.180 6.540 ;
        RECT 438.300 1.220 439.700 1.500 ;
        RECT 439.420 0.940 439.700 1.220 ;
        RECT 441.100 0.940 441.380 0.990 ;
        RECT 442.780 0.940 443.060 2.670 ;
        RECT 439.420 0.660 440.820 0.940 ;
        RECT 439.420 0.610 439.700 0.660 ;
        RECT 438.300 0.380 438.580 0.430 ;
        RECT 437.740 0.100 438.580 0.380 ;
        RECT 438.300 0.050 438.580 0.100 ;
        RECT 440.540 -0.180 440.820 0.660 ;
        RECT 441.100 0.660 443.060 0.940 ;
        RECT 441.100 0.610 441.380 0.660 ;
        RECT 442.220 -0.180 442.500 -0.130 ;
        RECT 440.540 -0.460 442.500 -0.180 ;
        RECT 437.180 -6.340 437.460 -4.050 ;
        RECT 440.540 -4.430 440.820 -0.460 ;
        RECT 442.220 -0.510 442.500 -0.460 ;
        RECT 437.180 -6.620 438.580 -6.340 ;
        RECT 437.180 -6.670 437.460 -6.620 ;
        RECT 438.300 -7.930 438.580 -6.620 ;
        RECT 441.100 -12.410 441.380 -11.890 ;
        RECT 432.700 -18.660 432.980 -18.610 ;
        RECT 432.140 -18.940 432.980 -18.660 ;
        RECT 423.740 -23.140 424.580 -22.860 ;
        RECT 425.980 -23.140 426.820 -22.860 ;
        RECT 424.300 -23.470 424.580 -23.140 ;
        RECT 424.300 -27.620 424.580 -27.010 ;
        RECT 425.980 -27.530 426.260 -27.010 ;
        RECT 424.300 -27.900 425.700 -27.620 ;
        RECT 425.420 -28.180 425.700 -27.900 ;
        RECT 425.420 -28.460 426.260 -28.180 ;
        RECT 424.860 -28.740 425.140 -28.690 ;
        RECT 424.860 -29.020 425.700 -28.740 ;
        RECT 424.860 -29.070 425.140 -29.020 ;
        RECT 423.180 -31.870 423.460 -30.930 ;
        RECT 423.740 -36.020 424.020 -31.490 ;
        RECT 424.860 -31.540 425.140 -31.490 ;
        RECT 423.180 -36.300 424.020 -36.020 ;
        RECT 424.300 -31.820 425.140 -31.540 ;
        RECT 418.140 -38.730 418.420 -38.210 ;
        RECT 423.180 -38.590 423.460 -36.300 ;
        RECT 424.300 -37.700 424.580 -31.820 ;
        RECT 424.860 -31.870 425.140 -31.820 ;
        RECT 425.420 -31.870 425.700 -29.020 ;
        RECT 425.980 -32.660 426.260 -28.460 ;
        RECT 426.540 -31.870 426.820 -23.140 ;
        RECT 431.580 -23.470 431.860 -19.730 ;
        RECT 432.140 -20.110 432.420 -18.940 ;
        RECT 432.700 -18.990 432.980 -18.940 ;
        RECT 433.820 -19.780 434.100 -19.730 ;
        RECT 432.700 -20.060 434.100 -19.780 ;
        RECT 427.660 -28.180 427.940 -27.010 ;
        RECT 427.660 -28.460 429.060 -28.180 ;
        RECT 427.660 -28.510 427.940 -28.460 ;
        RECT 428.780 -32.010 429.060 -28.460 ;
        RECT 431.580 -28.510 431.860 -27.570 ;
        RECT 430.460 -31.450 430.740 -30.930 ;
        RECT 432.140 -32.570 432.420 -32.050 ;
        RECT 427.660 -32.660 427.940 -32.610 ;
        RECT 425.980 -32.940 427.940 -32.660 ;
        RECT 427.660 -33.130 427.940 -32.940 ;
        RECT 423.740 -37.980 424.580 -37.700 ;
        RECT 406.380 -42.460 409.460 -42.180 ;
        RECT 406.380 -43.070 406.660 -42.460 ;
        RECT 409.180 -42.510 409.460 -42.460 ;
        RECT 417.580 -42.180 417.860 -42.130 ;
        RECT 418.700 -42.180 418.980 -39.890 ;
        RECT 423.740 -40.270 424.020 -37.980 ;
        RECT 428.220 -39.380 428.500 -32.610 ;
        RECT 424.860 -39.660 428.500 -39.380 ;
        RECT 417.580 -42.460 418.980 -42.180 ;
        RECT 417.580 -42.510 417.860 -42.460 ;
        RECT 418.700 -43.070 418.980 -42.460 ;
        RECT 421.500 -43.770 421.780 -43.250 ;
        RECT 423.740 -43.860 424.020 -43.250 ;
        RECT 424.860 -43.860 425.140 -39.660 ;
        RECT 431.020 -39.710 431.300 -32.610 ;
        RECT 432.700 -33.220 432.980 -20.060 ;
        RECT 433.820 -20.110 434.100 -20.060 ;
        RECT 436.620 -20.110 436.900 -19.590 ;
        RECT 432.140 -33.500 432.980 -33.220 ;
        RECT 423.740 -44.140 425.140 -43.860 ;
        RECT 398.540 -47.130 398.820 -46.610 ;
        RECT 389.580 -47.690 389.860 -47.170 ;
        RECT 392.940 -47.690 393.220 -47.170 ;
        RECT 405.820 -61.000 406.100 -46.610 ;
        RECT 406.940 -47.220 407.220 -44.370 ;
        RECT 417.020 -47.130 417.300 -46.610 ;
        RECT 411.980 -47.220 412.260 -47.170 ;
        RECT 406.940 -47.500 412.260 -47.220 ;
        RECT 411.980 -47.550 412.260 -47.500 ;
        RECT 419.260 -47.550 419.540 -44.370 ;
        RECT 427.100 -46.430 427.380 -40.450 ;
        RECT 431.580 -44.190 431.860 -39.330 ;
        RECT 432.140 -43.630 432.420 -33.500 ;
        RECT 432.700 -33.690 432.980 -33.500 ;
        RECT 432.700 -35.370 432.980 -34.850 ;
        RECT 433.260 -36.350 433.540 -21.410 ;
        RECT 435.500 -23.610 435.780 -23.090 ;
        RECT 435.500 -27.620 435.780 -27.570 ;
        RECT 436.620 -27.620 436.900 -20.850 ;
        RECT 437.180 -23.470 437.460 -18.610 ;
        RECT 438.300 -24.730 438.580 -24.210 ;
        RECT 439.980 -24.260 440.260 -24.210 ;
        RECT 438.860 -24.540 440.260 -24.260 ;
        RECT 438.860 -25.940 439.140 -24.540 ;
        RECT 439.980 -24.590 440.260 -24.540 ;
        RECT 437.180 -26.220 439.140 -25.940 ;
        RECT 437.180 -26.830 437.460 -26.220 ;
        RECT 438.860 -27.620 439.140 -27.570 ;
        RECT 435.500 -27.900 436.340 -27.620 ;
        RECT 436.620 -27.900 439.140 -27.620 ;
        RECT 435.500 -28.090 435.780 -27.900 ;
        RECT 434.380 -30.750 434.660 -28.130 ;
        RECT 436.060 -28.740 436.340 -27.900 ;
        RECT 438.860 -27.950 439.140 -27.900 ;
        RECT 436.060 -29.020 438.580 -28.740 ;
        RECT 437.180 -31.450 437.460 -30.930 ;
        RECT 438.300 -31.310 438.580 -29.020 ;
        RECT 435.500 -38.590 435.780 -35.410 ;
        RECT 436.060 -39.150 436.340 -31.490 ;
        RECT 438.860 -31.540 439.140 -31.490 ;
        RECT 438.860 -31.820 439.700 -31.540 ;
        RECT 438.860 -31.870 439.140 -31.820 ;
        RECT 439.420 -32.430 439.700 -31.820 ;
        RECT 439.980 -32.010 440.260 -31.490 ;
        RECT 442.220 -31.540 442.500 -31.490 ;
        RECT 442.780 -31.540 443.060 -7.970 ;
        RECT 443.340 -12.270 443.620 -7.410 ;
        RECT 443.900 -22.860 444.180 6.260 ;
        RECT 446.140 -1.070 446.420 10.460 ;
        RECT 447.820 7.330 448.100 20.030 ;
        RECT 454.540 3.270 454.820 3.790 ;
        RECT 455.100 2.620 455.380 27.540 ;
        RECT 456.220 27.260 456.500 27.310 ;
        RECT 455.660 26.980 456.500 27.260 ;
        RECT 455.660 23.010 455.940 26.980 ;
        RECT 456.220 26.930 456.500 26.980 ;
        RECT 456.220 26.140 456.500 26.190 ;
        RECT 456.220 25.860 457.620 26.140 ;
        RECT 456.220 25.810 456.500 25.860 ;
        RECT 457.340 23.010 457.620 25.860 ;
        RECT 457.340 19.090 457.620 22.270 ;
        RECT 457.340 15.170 457.620 16.670 ;
        RECT 459.020 15.500 459.300 27.310 ;
        RECT 459.580 23.010 459.860 39.070 ;
        RECT 460.140 30.620 460.420 30.670 ;
        RECT 460.140 30.340 460.980 30.620 ;
        RECT 460.140 30.290 460.420 30.340 ;
        RECT 460.140 20.210 460.420 29.550 ;
        RECT 459.580 15.500 459.860 15.550 ;
        RECT 459.020 15.220 459.860 15.500 ;
        RECT 456.780 2.620 457.060 3.230 ;
        RECT 454.540 2.340 457.060 2.620 ;
        RECT 445.020 -8.350 445.300 -6.850 ;
        RECT 442.220 -31.820 443.060 -31.540 ;
        RECT 443.340 -23.140 444.180 -22.860 ;
        RECT 440.540 -32.570 440.820 -32.050 ;
        RECT 437.180 -35.930 437.460 -32.610 ;
        RECT 442.220 -33.550 442.500 -31.820 ;
        RECT 436.060 -42.180 436.340 -42.130 ;
        RECT 436.620 -42.180 436.900 -38.210 ;
        RECT 439.420 -38.820 439.700 -35.410 ;
        RECT 437.180 -39.100 439.700 -38.820 ;
        RECT 437.180 -39.710 437.460 -39.100 ;
        RECT 438.860 -40.410 439.140 -39.890 ;
        RECT 436.060 -42.460 436.900 -42.180 ;
        RECT 438.860 -42.180 439.140 -42.130 ;
        RECT 439.420 -42.180 439.700 -39.100 ;
        RECT 442.780 -39.380 443.060 -39.330 ;
        RECT 438.860 -42.460 439.700 -42.180 ;
        RECT 441.660 -39.660 443.060 -39.380 ;
        RECT 436.060 -42.510 436.340 -42.460 ;
        RECT 438.860 -42.510 439.140 -42.460 ;
        RECT 441.660 -42.510 441.940 -39.660 ;
        RECT 442.780 -39.710 443.060 -39.660 ;
        RECT 443.340 -42.180 443.620 -23.140 ;
        RECT 443.900 -36.350 444.180 -24.770 ;
        RECT 445.020 -32.010 445.300 -31.490 ;
        RECT 444.460 -34.670 444.740 -32.050 ;
        RECT 445.020 -35.230 445.300 -32.610 ;
        RECT 445.580 -36.910 445.860 -24.210 ;
        RECT 446.140 -34.670 446.420 -10.770 ;
        RECT 448.380 -16.190 448.660 -10.210 ;
        RECT 447.260 -26.830 447.540 -23.650 ;
        RECT 448.380 -34.810 448.660 -34.290 ;
        RECT 446.700 -36.350 446.980 -35.410 ;
        RECT 449.500 -38.590 449.780 -16.930 ;
        RECT 452.300 -19.130 452.580 -18.610 ;
        RECT 450.060 -34.670 450.340 -28.130 ;
        RECT 451.180 -35.790 451.460 -34.290 ;
        RECT 453.420 -39.150 453.700 -19.730 ;
        RECT 447.820 -40.500 448.100 -40.450 ;
        RECT 445.580 -40.780 448.100 -40.500 ;
        RECT 443.900 -42.180 444.180 -42.130 ;
        RECT 442.220 -42.460 444.180 -42.180 ;
        RECT 441.100 -43.300 441.380 -43.250 ;
        RECT 442.220 -43.300 442.500 -42.460 ;
        RECT 443.900 -42.510 444.180 -42.460 ;
        RECT 441.100 -43.580 442.500 -43.300 ;
        RECT 441.100 -43.630 441.380 -43.580 ;
        RECT 423.740 -61.000 424.020 -46.610 ;
        RECT 436.060 -47.130 436.340 -46.610 ;
        RECT 432.140 -47.690 432.420 -47.170 ;
        RECT 441.660 -60.380 443.620 -60.100 ;
        RECT 441.660 -61.000 441.940 -60.380 ;
        RECT 298.160 -63.190 298.720 -61.000 ;
        RECT 144.850 -63.590 298.720 -63.190 ;
        RECT 120.925 -63.715 121.925 -63.665 ;
        RECT 120.925 -64.115 143.995 -63.715 ;
        RECT 120.925 -64.165 121.925 -64.115 ;
        RECT 298.160 -65.000 298.720 -63.590 ;
        RECT 97.315 -67.875 97.715 -66.675 ;
        RECT 98.495 -66.685 100.455 -66.285 ;
        RECT 316.080 -66.550 316.640 -61.000 ;
        RECT 144.850 -66.950 316.640 -66.550 ;
        RECT 120.925 -67.075 121.925 -67.025 ;
        RECT 120.925 -67.475 143.995 -67.075 ;
        RECT 120.925 -67.525 121.925 -67.475 ;
        RECT 334.000 -69.910 334.560 -61.000 ;
        RECT 96.195 -71.235 96.595 -70.035 ;
        RECT 144.850 -70.310 334.560 -69.910 ;
        RECT 120.925 -70.435 121.925 -70.385 ;
        RECT 120.925 -70.835 143.995 -70.435 ;
        RECT 120.925 -70.885 121.925 -70.835 ;
        RECT 351.920 -73.270 352.480 -61.000 ;
        RECT 93.955 -74.595 94.355 -73.395 ;
        RECT 144.850 -73.670 352.480 -73.270 ;
        RECT 120.925 -73.795 121.925 -73.745 ;
        RECT 120.925 -74.195 143.995 -73.795 ;
        RECT 120.925 -74.245 121.925 -74.195 ;
        RECT 369.840 -76.630 370.400 -61.000 ;
        RECT 89.475 -77.955 89.875 -76.755 ;
        RECT 144.850 -77.030 370.400 -76.630 ;
        RECT 120.925 -77.155 121.925 -77.105 ;
        RECT 120.925 -77.555 143.995 -77.155 ;
        RECT 120.925 -77.605 121.925 -77.555 ;
        RECT 387.760 -79.990 388.320 -61.000 ;
        RECT 80.515 -81.315 80.915 -80.115 ;
        RECT 144.850 -80.390 388.320 -79.990 ;
        RECT 120.925 -80.515 121.925 -80.465 ;
        RECT 120.925 -80.915 143.995 -80.515 ;
        RECT 120.925 -80.965 121.925 -80.915 ;
        RECT 405.680 -83.350 406.240 -61.000 ;
        RECT 62.595 -84.675 62.995 -83.475 ;
        RECT 144.850 -83.750 406.240 -83.350 ;
        RECT 120.925 -83.875 121.925 -83.825 ;
        RECT 120.925 -84.275 143.995 -83.875 ;
        RECT 120.925 -84.325 121.925 -84.275 ;
        RECT 423.600 -86.710 424.160 -61.000 ;
        RECT 26.755 -88.035 27.155 -86.835 ;
        RECT 144.850 -87.110 424.160 -86.710 ;
        RECT 120.925 -87.235 121.925 -87.185 ;
        RECT 120.925 -87.635 143.995 -87.235 ;
        RECT 120.925 -87.685 121.925 -87.635 ;
        RECT 441.520 -90.070 442.080 -61.000 ;
        RECT 443.340 -61.220 443.620 -60.380 ;
        RECT 445.580 -61.220 445.860 -40.780 ;
        RECT 447.820 -40.830 448.100 -40.780 ;
        RECT 450.060 -42.180 450.340 -42.130 ;
        RECT 454.540 -42.180 454.820 2.340 ;
        RECT 457.340 -0.650 457.620 -0.130 ;
        RECT 459.580 -1.070 459.860 15.220 ;
        RECT 460.140 10.740 460.420 11.070 ;
        RECT 460.700 10.740 460.980 30.340 ;
        RECT 460.140 10.460 460.980 10.740 ;
        RECT 457.340 -8.020 457.620 -4.050 ;
        RECT 460.140 -4.430 460.420 10.460 ;
        RECT 455.100 -8.300 457.620 -8.020 ;
        RECT 455.100 -22.860 455.380 -8.300 ;
        RECT 456.780 -9.140 457.060 -9.090 ;
        RECT 456.220 -9.420 457.060 -9.140 ;
        RECT 456.220 -17.310 456.500 -9.420 ;
        RECT 456.780 -9.470 457.060 -9.420 ;
        RECT 460.700 -9.610 460.980 -9.090 ;
        RECT 456.220 -19.780 456.500 -19.730 ;
        RECT 458.460 -19.780 458.740 -19.170 ;
        RECT 456.220 -20.060 458.740 -19.780 ;
        RECT 456.220 -20.250 456.500 -20.060 ;
        RECT 455.100 -23.140 457.620 -22.860 ;
        RECT 459.020 -22.910 459.300 -19.730 ;
        RECT 457.340 -26.830 457.620 -23.140 ;
        RECT 456.780 -30.420 457.060 -30.370 ;
        RECT 456.220 -30.700 457.060 -30.420 ;
        RECT 455.100 -34.810 455.380 -34.290 ;
        RECT 455.100 -41.620 455.380 -35.970 ;
        RECT 455.100 -41.900 455.940 -41.620 ;
        RECT 450.060 -42.460 454.820 -42.180 ;
        RECT 450.060 -42.510 450.340 -42.460 ;
        RECT 454.540 -42.740 454.820 -42.460 ;
        RECT 455.100 -42.740 455.380 -42.690 ;
        RECT 454.540 -43.020 455.380 -42.740 ;
        RECT 455.100 -43.070 455.380 -43.020 ;
        RECT 454.540 -44.330 454.820 -43.810 ;
        RECT 455.660 -44.980 455.940 -41.900 ;
        RECT 453.980 -45.260 455.940 -44.980 ;
        RECT 453.980 -46.990 454.260 -45.260 ;
        RECT 456.220 -47.780 456.500 -30.700 ;
        RECT 456.780 -30.750 457.060 -30.700 ;
        RECT 459.580 -30.750 459.860 -19.730 ;
        RECT 456.780 -35.460 457.060 -32.050 ;
        RECT 457.340 -35.460 457.620 -35.410 ;
        RECT 456.780 -35.740 457.620 -35.460 ;
        RECT 457.340 -35.790 457.620 -35.740 ;
        RECT 457.340 -39.150 457.620 -37.650 ;
        RECT 456.780 -47.780 457.060 -47.730 ;
        RECT 456.220 -48.060 457.060 -47.780 ;
        RECT 457.900 -47.780 458.180 -36.530 ;
        RECT 458.460 -42.510 458.740 -30.930 ;
        RECT 460.140 -36.350 460.420 -28.130 ;
        RECT 460.700 -33.130 460.980 -32.610 ;
        RECT 458.460 -47.780 458.740 -47.730 ;
        RECT 457.900 -48.060 458.740 -47.780 ;
        RECT 456.780 -48.110 457.060 -48.060 ;
        RECT 458.460 -48.110 458.740 -48.060 ;
        RECT 459.580 -61.000 459.860 -46.050 ;
        RECT 443.340 -61.500 445.860 -61.220 ;
        RECT -44.925 -91.395 -44.525 -90.195 ;
        RECT 144.850 -90.470 442.080 -90.070 ;
        RECT 120.925 -90.595 121.925 -90.545 ;
        RECT 120.925 -90.995 143.995 -90.595 ;
        RECT 120.925 -91.045 121.925 -90.995 ;
        RECT 459.440 -93.430 460.000 -61.000 ;
        RECT -188.285 -94.755 -187.885 -93.555 ;
        RECT 144.850 -93.830 460.000 -93.430 ;
        RECT 120.925 -93.955 121.925 -93.905 ;
        RECT 120.925 -94.355 143.995 -93.955 ;
        RECT 120.925 -94.405 121.925 -94.355 ;
        RECT -491.830 -105.625 -491.430 -97.075 ;
        RECT -189.405 -98.115 -189.005 -96.915 ;
        RECT 120.925 -97.315 121.925 -97.265 ;
        RECT 120.925 -97.715 143.995 -97.315 ;
        RECT 120.925 -97.765 121.925 -97.715 ;
        RECT 468.200 -105.525 469.200 105.525 ;
        RECT -492.150 -106.425 -491.110 -105.625 ;
        RECT 466.700 -106.525 469.200 -105.525 ;
      LAYER Via2 ;
        RECT -492.030 105.885 -491.230 106.165 ;
        RECT 467.250 106.165 467.530 106.445 ;
        RECT 467.810 106.165 468.090 106.445 ;
        RECT 468.370 106.165 468.650 106.445 ;
        RECT 467.250 105.605 467.530 105.885 ;
        RECT 467.810 105.605 468.090 105.885 ;
        RECT 468.370 105.605 468.650 105.885 ;
        RECT -189.345 97.675 -189.065 97.955 ;
        RECT -189.345 97.075 -189.065 97.355 ;
        RECT 121.025 97.375 121.825 97.655 ;
        RECT -332.705 90.955 -332.425 91.235 ;
        RECT -332.705 90.355 -332.425 90.635 ;
        RECT -404.385 87.595 -404.105 87.875 ;
        RECT -404.385 86.995 -404.105 87.275 ;
        RECT -440.225 84.235 -439.945 84.515 ;
        RECT -497.475 83.425 -495.635 83.705 ;
        RECT -440.225 83.635 -439.945 83.915 ;
        RECT -486.895 81.275 -486.615 83.115 ;
        RECT -458.145 80.875 -457.865 81.155 ;
        RECT -458.145 80.275 -457.865 80.555 ;
        RECT -467.105 77.515 -466.825 77.795 ;
        RECT -467.105 76.915 -466.825 77.195 ;
        RECT -471.585 74.155 -471.305 74.435 ;
        RECT -471.585 73.555 -471.305 73.835 ;
        RECT -473.825 70.795 -473.545 71.075 ;
        RECT -473.825 70.195 -473.545 70.475 ;
        RECT -474.945 67.435 -474.665 67.715 ;
        RECT -474.945 66.835 -474.665 67.115 ;
        RECT -472.705 67.435 -472.425 67.715 ;
        RECT -472.705 66.835 -472.425 67.115 ;
        RECT -469.345 70.795 -469.065 71.075 ;
        RECT -469.345 70.195 -469.065 70.475 ;
        RECT -470.465 67.435 -470.185 67.715 ;
        RECT -470.465 66.835 -470.185 67.115 ;
        RECT -468.225 67.435 -467.945 67.715 ;
        RECT -468.225 66.835 -467.945 67.115 ;
        RECT -462.625 74.155 -462.345 74.435 ;
        RECT -462.625 73.555 -462.345 73.835 ;
        RECT -464.865 70.795 -464.585 71.075 ;
        RECT -464.865 70.195 -464.585 70.475 ;
        RECT -465.985 67.435 -465.705 67.715 ;
        RECT -465.985 66.835 -465.705 67.115 ;
        RECT -463.745 67.435 -463.465 67.715 ;
        RECT -463.745 66.835 -463.465 67.115 ;
        RECT -460.385 70.795 -460.105 71.075 ;
        RECT -460.385 70.195 -460.105 70.475 ;
        RECT -461.505 67.435 -461.225 67.715 ;
        RECT -461.505 66.835 -461.225 67.115 ;
        RECT -459.265 67.435 -458.985 67.715 ;
        RECT -459.265 66.835 -458.985 67.115 ;
        RECT -449.185 77.515 -448.905 77.795 ;
        RECT -449.185 76.915 -448.905 77.195 ;
        RECT -453.665 74.155 -453.385 74.435 ;
        RECT -453.665 73.555 -453.385 73.835 ;
        RECT -455.905 70.795 -455.625 71.075 ;
        RECT -455.905 70.195 -455.625 70.475 ;
        RECT -457.025 67.435 -456.745 67.715 ;
        RECT -457.025 66.835 -456.745 67.115 ;
        RECT -454.785 67.435 -454.505 67.715 ;
        RECT -454.785 66.835 -454.505 67.115 ;
        RECT -451.425 70.795 -451.145 71.075 ;
        RECT -451.425 70.195 -451.145 70.475 ;
        RECT -452.545 67.435 -452.265 67.715 ;
        RECT -452.545 66.835 -452.265 67.115 ;
        RECT -450.305 67.435 -450.025 67.715 ;
        RECT -450.305 66.835 -450.025 67.115 ;
        RECT -444.705 74.155 -444.425 74.435 ;
        RECT -444.705 73.555 -444.425 73.835 ;
        RECT -446.945 70.795 -446.665 71.075 ;
        RECT -446.945 70.195 -446.665 70.475 ;
        RECT -448.065 67.435 -447.785 67.715 ;
        RECT -448.065 66.835 -447.785 67.115 ;
        RECT -445.825 67.435 -445.545 67.715 ;
        RECT -445.825 66.835 -445.545 67.115 ;
        RECT -442.465 70.795 -442.185 71.075 ;
        RECT -442.465 70.195 -442.185 70.475 ;
        RECT -443.585 67.435 -443.305 67.715 ;
        RECT -443.585 66.835 -443.305 67.115 ;
        RECT -441.345 67.435 -441.065 67.715 ;
        RECT -441.345 66.835 -441.065 67.115 ;
        RECT -422.305 80.875 -422.025 81.155 ;
        RECT -422.305 80.275 -422.025 80.555 ;
        RECT -431.265 77.515 -430.985 77.795 ;
        RECT -431.265 76.915 -430.985 77.195 ;
        RECT -435.745 74.155 -435.465 74.435 ;
        RECT -435.745 73.555 -435.465 73.835 ;
        RECT -437.985 70.795 -437.705 71.075 ;
        RECT -437.985 70.195 -437.705 70.475 ;
        RECT -439.105 67.435 -438.825 67.715 ;
        RECT -439.105 66.835 -438.825 67.115 ;
        RECT -436.865 67.435 -436.585 67.715 ;
        RECT -436.865 66.835 -436.585 67.115 ;
        RECT -433.505 70.795 -433.225 71.075 ;
        RECT -433.505 70.195 -433.225 70.475 ;
        RECT -434.625 67.435 -434.345 67.715 ;
        RECT -434.625 66.835 -434.345 67.115 ;
        RECT -432.385 67.435 -432.105 67.715 ;
        RECT -432.385 66.835 -432.105 67.115 ;
        RECT -426.785 74.155 -426.505 74.435 ;
        RECT -426.785 73.555 -426.505 73.835 ;
        RECT -429.025 70.795 -428.745 71.075 ;
        RECT -429.025 70.195 -428.745 70.475 ;
        RECT -430.145 67.435 -429.865 67.715 ;
        RECT -430.145 66.835 -429.865 67.115 ;
        RECT -427.905 67.435 -427.625 67.715 ;
        RECT -427.905 66.835 -427.625 67.115 ;
        RECT -424.545 70.795 -424.265 71.075 ;
        RECT -424.545 70.195 -424.265 70.475 ;
        RECT -425.665 67.435 -425.385 67.715 ;
        RECT -425.665 66.835 -425.385 67.115 ;
        RECT -423.425 67.435 -423.145 67.715 ;
        RECT -423.425 66.835 -423.145 67.115 ;
        RECT -413.345 77.515 -413.065 77.795 ;
        RECT -413.345 76.915 -413.065 77.195 ;
        RECT -417.825 74.155 -417.545 74.435 ;
        RECT -417.825 73.555 -417.545 73.835 ;
        RECT -420.065 70.795 -419.785 71.075 ;
        RECT -420.065 70.195 -419.785 70.475 ;
        RECT -421.185 67.435 -420.905 67.715 ;
        RECT -421.185 66.835 -420.905 67.115 ;
        RECT -418.945 67.435 -418.665 67.715 ;
        RECT -418.945 66.835 -418.665 67.115 ;
        RECT -415.585 70.795 -415.305 71.075 ;
        RECT -415.585 70.195 -415.305 70.475 ;
        RECT -416.705 67.435 -416.425 67.715 ;
        RECT -416.705 66.835 -416.425 67.115 ;
        RECT -414.465 67.435 -414.185 67.715 ;
        RECT -414.465 66.835 -414.185 67.115 ;
        RECT -408.865 74.155 -408.585 74.435 ;
        RECT -408.865 73.555 -408.585 73.835 ;
        RECT -411.105 70.795 -410.825 71.075 ;
        RECT -411.105 70.195 -410.825 70.475 ;
        RECT -412.225 67.435 -411.945 67.715 ;
        RECT -412.225 66.835 -411.945 67.115 ;
        RECT -409.985 67.435 -409.705 67.715 ;
        RECT -409.985 66.835 -409.705 67.115 ;
        RECT -406.625 70.795 -406.345 71.075 ;
        RECT -406.625 70.195 -406.345 70.475 ;
        RECT -407.745 67.435 -407.465 67.715 ;
        RECT -407.745 66.835 -407.465 67.115 ;
        RECT -405.505 67.435 -405.225 67.715 ;
        RECT -405.505 66.835 -405.225 67.115 ;
        RECT -368.545 84.235 -368.265 84.515 ;
        RECT -368.545 83.635 -368.265 83.915 ;
        RECT -386.465 80.875 -386.185 81.155 ;
        RECT -386.465 80.275 -386.185 80.555 ;
        RECT -395.425 77.515 -395.145 77.795 ;
        RECT -395.425 76.915 -395.145 77.195 ;
        RECT -399.905 74.155 -399.625 74.435 ;
        RECT -399.905 73.555 -399.625 73.835 ;
        RECT -402.145 70.795 -401.865 71.075 ;
        RECT -402.145 70.195 -401.865 70.475 ;
        RECT -403.265 67.435 -402.985 67.715 ;
        RECT -403.265 66.835 -402.985 67.115 ;
        RECT -401.025 67.435 -400.745 67.715 ;
        RECT -401.025 66.835 -400.745 67.115 ;
        RECT -397.665 70.795 -397.385 71.075 ;
        RECT -397.665 70.195 -397.385 70.475 ;
        RECT -398.785 67.435 -398.505 67.715 ;
        RECT -398.785 66.835 -398.505 67.115 ;
        RECT -396.545 67.435 -396.265 67.715 ;
        RECT -396.545 66.835 -396.265 67.115 ;
        RECT -390.945 74.155 -390.665 74.435 ;
        RECT -390.945 73.555 -390.665 73.835 ;
        RECT -393.185 70.795 -392.905 71.075 ;
        RECT -393.185 70.195 -392.905 70.475 ;
        RECT -394.305 67.435 -394.025 67.715 ;
        RECT -394.305 66.835 -394.025 67.115 ;
        RECT -392.065 67.435 -391.785 67.715 ;
        RECT -392.065 66.835 -391.785 67.115 ;
        RECT -388.705 70.795 -388.425 71.075 ;
        RECT -388.705 70.195 -388.425 70.475 ;
        RECT -389.825 67.435 -389.545 67.715 ;
        RECT -389.825 66.835 -389.545 67.115 ;
        RECT -387.585 67.435 -387.305 67.715 ;
        RECT -387.585 66.835 -387.305 67.115 ;
        RECT -377.505 77.515 -377.225 77.795 ;
        RECT -377.505 76.915 -377.225 77.195 ;
        RECT -381.985 74.155 -381.705 74.435 ;
        RECT -381.985 73.555 -381.705 73.835 ;
        RECT -384.225 70.795 -383.945 71.075 ;
        RECT -384.225 70.195 -383.945 70.475 ;
        RECT -385.345 67.435 -385.065 67.715 ;
        RECT -385.345 66.835 -385.065 67.115 ;
        RECT -383.105 67.435 -382.825 67.715 ;
        RECT -383.105 66.835 -382.825 67.115 ;
        RECT -379.745 70.795 -379.465 71.075 ;
        RECT -379.745 70.195 -379.465 70.475 ;
        RECT -380.865 67.435 -380.585 67.715 ;
        RECT -380.865 66.835 -380.585 67.115 ;
        RECT -378.625 67.435 -378.345 67.715 ;
        RECT -378.625 66.835 -378.345 67.115 ;
        RECT -373.025 74.155 -372.745 74.435 ;
        RECT -373.025 73.555 -372.745 73.835 ;
        RECT -375.265 70.795 -374.985 71.075 ;
        RECT -375.265 70.195 -374.985 70.475 ;
        RECT -376.385 67.435 -376.105 67.715 ;
        RECT -376.385 66.835 -376.105 67.115 ;
        RECT -374.145 67.435 -373.865 67.715 ;
        RECT -374.145 66.835 -373.865 67.115 ;
        RECT -370.785 70.795 -370.505 71.075 ;
        RECT -370.785 70.195 -370.505 70.475 ;
        RECT -371.905 67.435 -371.625 67.715 ;
        RECT -371.905 66.835 -371.625 67.115 ;
        RECT -369.665 67.435 -369.385 67.715 ;
        RECT -369.665 66.835 -369.385 67.115 ;
        RECT -350.625 80.875 -350.345 81.155 ;
        RECT -350.625 80.275 -350.345 80.555 ;
        RECT -359.585 77.515 -359.305 77.795 ;
        RECT -359.585 76.915 -359.305 77.195 ;
        RECT -364.065 74.155 -363.785 74.435 ;
        RECT -364.065 73.555 -363.785 73.835 ;
        RECT -366.305 70.795 -366.025 71.075 ;
        RECT -366.305 70.195 -366.025 70.475 ;
        RECT -367.425 67.435 -367.145 67.715 ;
        RECT -367.425 66.835 -367.145 67.115 ;
        RECT -365.185 67.435 -364.905 67.715 ;
        RECT -365.185 66.835 -364.905 67.115 ;
        RECT -361.825 70.795 -361.545 71.075 ;
        RECT -361.825 70.195 -361.545 70.475 ;
        RECT -362.945 67.435 -362.665 67.715 ;
        RECT -362.945 66.835 -362.665 67.115 ;
        RECT -360.705 67.435 -360.425 67.715 ;
        RECT -360.705 66.835 -360.425 67.115 ;
        RECT -355.105 74.155 -354.825 74.435 ;
        RECT -355.105 73.555 -354.825 73.835 ;
        RECT -357.345 70.795 -357.065 71.075 ;
        RECT -357.345 70.195 -357.065 70.475 ;
        RECT -358.465 67.435 -358.185 67.715 ;
        RECT -358.465 66.835 -358.185 67.115 ;
        RECT -356.225 67.435 -355.945 67.715 ;
        RECT -356.225 66.835 -355.945 67.115 ;
        RECT -352.865 70.795 -352.585 71.075 ;
        RECT -352.865 70.195 -352.585 70.475 ;
        RECT -353.985 67.435 -353.705 67.715 ;
        RECT -353.985 66.835 -353.705 67.115 ;
        RECT -351.745 67.435 -351.465 67.715 ;
        RECT -351.745 66.835 -351.465 67.115 ;
        RECT -341.665 77.515 -341.385 77.795 ;
        RECT -341.665 76.915 -341.385 77.195 ;
        RECT -346.145 74.155 -345.865 74.435 ;
        RECT -346.145 73.555 -345.865 73.835 ;
        RECT -348.385 70.795 -348.105 71.075 ;
        RECT -348.385 70.195 -348.105 70.475 ;
        RECT -349.505 67.435 -349.225 67.715 ;
        RECT -349.505 66.835 -349.225 67.115 ;
        RECT -347.265 67.435 -346.985 67.715 ;
        RECT -347.265 66.835 -346.985 67.115 ;
        RECT -343.905 70.795 -343.625 71.075 ;
        RECT -343.905 70.195 -343.625 70.475 ;
        RECT -345.025 67.435 -344.745 67.715 ;
        RECT -345.025 66.835 -344.745 67.115 ;
        RECT -342.785 67.435 -342.505 67.715 ;
        RECT -342.785 66.835 -342.505 67.115 ;
        RECT -337.185 74.155 -336.905 74.435 ;
        RECT -337.185 73.555 -336.905 73.835 ;
        RECT -339.425 70.795 -339.145 71.075 ;
        RECT -339.425 70.195 -339.145 70.475 ;
        RECT -340.545 67.435 -340.265 67.715 ;
        RECT -340.545 66.835 -340.265 67.115 ;
        RECT -338.305 67.435 -338.025 67.715 ;
        RECT -338.305 66.835 -338.025 67.115 ;
        RECT -334.945 70.795 -334.665 71.075 ;
        RECT -334.945 70.195 -334.665 70.475 ;
        RECT -336.065 67.435 -335.785 67.715 ;
        RECT -336.065 66.835 -335.785 67.115 ;
        RECT -333.825 67.435 -333.545 67.715 ;
        RECT -333.825 66.835 -333.545 67.115 ;
        RECT -261.025 87.595 -260.745 87.875 ;
        RECT -261.025 86.995 -260.745 87.275 ;
        RECT -296.865 84.235 -296.585 84.515 ;
        RECT -296.865 83.635 -296.585 83.915 ;
        RECT -314.785 80.875 -314.505 81.155 ;
        RECT -314.785 80.275 -314.505 80.555 ;
        RECT -323.745 77.515 -323.465 77.795 ;
        RECT -323.745 76.915 -323.465 77.195 ;
        RECT -328.225 74.155 -327.945 74.435 ;
        RECT -328.225 73.555 -327.945 73.835 ;
        RECT -330.465 70.795 -330.185 71.075 ;
        RECT -330.465 70.195 -330.185 70.475 ;
        RECT -331.585 67.435 -331.305 67.715 ;
        RECT -331.585 66.835 -331.305 67.115 ;
        RECT -329.345 67.435 -329.065 67.715 ;
        RECT -329.345 66.835 -329.065 67.115 ;
        RECT -325.985 70.795 -325.705 71.075 ;
        RECT -325.985 70.195 -325.705 70.475 ;
        RECT -327.105 67.435 -326.825 67.715 ;
        RECT -327.105 66.835 -326.825 67.115 ;
        RECT -324.865 67.435 -324.585 67.715 ;
        RECT -324.865 66.835 -324.585 67.115 ;
        RECT -319.265 74.155 -318.985 74.435 ;
        RECT -319.265 73.555 -318.985 73.835 ;
        RECT -321.505 70.795 -321.225 71.075 ;
        RECT -321.505 70.195 -321.225 70.475 ;
        RECT -322.625 67.435 -322.345 67.715 ;
        RECT -322.625 66.835 -322.345 67.115 ;
        RECT -320.385 67.435 -320.105 67.715 ;
        RECT -320.385 66.835 -320.105 67.115 ;
        RECT -317.025 70.795 -316.745 71.075 ;
        RECT -317.025 70.195 -316.745 70.475 ;
        RECT -318.145 67.435 -317.865 67.715 ;
        RECT -318.145 66.835 -317.865 67.115 ;
        RECT -315.905 67.435 -315.625 67.715 ;
        RECT -315.905 66.835 -315.625 67.115 ;
        RECT -305.825 77.515 -305.545 77.795 ;
        RECT -305.825 76.915 -305.545 77.195 ;
        RECT -310.305 74.155 -310.025 74.435 ;
        RECT -310.305 73.555 -310.025 73.835 ;
        RECT -312.545 70.795 -312.265 71.075 ;
        RECT -312.545 70.195 -312.265 70.475 ;
        RECT -313.665 67.435 -313.385 67.715 ;
        RECT -313.665 66.835 -313.385 67.115 ;
        RECT -311.425 67.435 -311.145 67.715 ;
        RECT -311.425 66.835 -311.145 67.115 ;
        RECT -308.065 70.795 -307.785 71.075 ;
        RECT -308.065 70.195 -307.785 70.475 ;
        RECT -309.185 67.435 -308.905 67.715 ;
        RECT -309.185 66.835 -308.905 67.115 ;
        RECT -306.945 67.435 -306.665 67.715 ;
        RECT -306.945 66.835 -306.665 67.115 ;
        RECT -301.345 74.155 -301.065 74.435 ;
        RECT -301.345 73.555 -301.065 73.835 ;
        RECT -303.585 70.795 -303.305 71.075 ;
        RECT -303.585 70.195 -303.305 70.475 ;
        RECT -304.705 67.435 -304.425 67.715 ;
        RECT -304.705 66.835 -304.425 67.115 ;
        RECT -302.465 67.435 -302.185 67.715 ;
        RECT -302.465 66.835 -302.185 67.115 ;
        RECT -299.105 70.795 -298.825 71.075 ;
        RECT -299.105 70.195 -298.825 70.475 ;
        RECT -300.225 67.435 -299.945 67.715 ;
        RECT -300.225 66.835 -299.945 67.115 ;
        RECT -297.985 67.435 -297.705 67.715 ;
        RECT -297.985 66.835 -297.705 67.115 ;
        RECT -278.945 80.875 -278.665 81.155 ;
        RECT -278.945 80.275 -278.665 80.555 ;
        RECT -287.905 77.515 -287.625 77.795 ;
        RECT -287.905 76.915 -287.625 77.195 ;
        RECT -292.385 74.155 -292.105 74.435 ;
        RECT -292.385 73.555 -292.105 73.835 ;
        RECT -294.625 70.795 -294.345 71.075 ;
        RECT -294.625 70.195 -294.345 70.475 ;
        RECT -295.745 67.435 -295.465 67.715 ;
        RECT -295.745 66.835 -295.465 67.115 ;
        RECT -293.505 67.435 -293.225 67.715 ;
        RECT -293.505 66.835 -293.225 67.115 ;
        RECT -290.145 70.795 -289.865 71.075 ;
        RECT -290.145 70.195 -289.865 70.475 ;
        RECT -291.265 67.435 -290.985 67.715 ;
        RECT -291.265 66.835 -290.985 67.115 ;
        RECT -289.025 67.435 -288.745 67.715 ;
        RECT -289.025 66.835 -288.745 67.115 ;
        RECT -283.425 74.155 -283.145 74.435 ;
        RECT -283.425 73.555 -283.145 73.835 ;
        RECT -285.665 70.795 -285.385 71.075 ;
        RECT -285.665 70.195 -285.385 70.475 ;
        RECT -286.785 67.435 -286.505 67.715 ;
        RECT -286.785 66.835 -286.505 67.115 ;
        RECT -284.545 67.435 -284.265 67.715 ;
        RECT -284.545 66.835 -284.265 67.115 ;
        RECT -281.185 70.795 -280.905 71.075 ;
        RECT -281.185 70.195 -280.905 70.475 ;
        RECT -282.305 67.435 -282.025 67.715 ;
        RECT -282.305 66.835 -282.025 67.115 ;
        RECT -280.065 67.435 -279.785 67.715 ;
        RECT -280.065 66.835 -279.785 67.115 ;
        RECT -269.985 77.515 -269.705 77.795 ;
        RECT -269.985 76.915 -269.705 77.195 ;
        RECT -274.465 74.155 -274.185 74.435 ;
        RECT -274.465 73.555 -274.185 73.835 ;
        RECT -276.705 70.795 -276.425 71.075 ;
        RECT -276.705 70.195 -276.425 70.475 ;
        RECT -277.825 67.435 -277.545 67.715 ;
        RECT -277.825 66.835 -277.545 67.115 ;
        RECT -275.585 67.435 -275.305 67.715 ;
        RECT -275.585 66.835 -275.305 67.115 ;
        RECT -272.225 70.795 -271.945 71.075 ;
        RECT -272.225 70.195 -271.945 70.475 ;
        RECT -273.345 67.435 -273.065 67.715 ;
        RECT -273.345 66.835 -273.065 67.115 ;
        RECT -271.105 67.435 -270.825 67.715 ;
        RECT -271.105 66.835 -270.825 67.115 ;
        RECT -265.505 74.155 -265.225 74.435 ;
        RECT -265.505 73.555 -265.225 73.835 ;
        RECT -267.745 70.795 -267.465 71.075 ;
        RECT -267.745 70.195 -267.465 70.475 ;
        RECT -268.865 67.435 -268.585 67.715 ;
        RECT -268.865 66.835 -268.585 67.115 ;
        RECT -266.625 67.435 -266.345 67.715 ;
        RECT -266.625 66.835 -266.345 67.115 ;
        RECT -263.265 70.795 -262.985 71.075 ;
        RECT -263.265 70.195 -262.985 70.475 ;
        RECT -264.385 67.435 -264.105 67.715 ;
        RECT -264.385 66.835 -264.105 67.115 ;
        RECT -262.145 67.435 -261.865 67.715 ;
        RECT -262.145 66.835 -261.865 67.115 ;
        RECT -225.185 84.235 -224.905 84.515 ;
        RECT -225.185 83.635 -224.905 83.915 ;
        RECT -243.105 80.875 -242.825 81.155 ;
        RECT -243.105 80.275 -242.825 80.555 ;
        RECT -252.065 77.515 -251.785 77.795 ;
        RECT -252.065 76.915 -251.785 77.195 ;
        RECT -256.545 74.155 -256.265 74.435 ;
        RECT -256.545 73.555 -256.265 73.835 ;
        RECT -258.785 70.795 -258.505 71.075 ;
        RECT -258.785 70.195 -258.505 70.475 ;
        RECT -259.905 67.435 -259.625 67.715 ;
        RECT -259.905 66.835 -259.625 67.115 ;
        RECT -257.665 67.435 -257.385 67.715 ;
        RECT -257.665 66.835 -257.385 67.115 ;
        RECT -254.305 70.795 -254.025 71.075 ;
        RECT -254.305 70.195 -254.025 70.475 ;
        RECT -255.425 67.435 -255.145 67.715 ;
        RECT -255.425 66.835 -255.145 67.115 ;
        RECT -253.185 67.435 -252.905 67.715 ;
        RECT -253.185 66.835 -252.905 67.115 ;
        RECT -247.585 74.155 -247.305 74.435 ;
        RECT -247.585 73.555 -247.305 73.835 ;
        RECT -249.825 70.795 -249.545 71.075 ;
        RECT -249.825 70.195 -249.545 70.475 ;
        RECT -250.945 67.435 -250.665 67.715 ;
        RECT -250.945 66.835 -250.665 67.115 ;
        RECT -248.705 67.435 -248.425 67.715 ;
        RECT -248.705 66.835 -248.425 67.115 ;
        RECT -245.345 70.795 -245.065 71.075 ;
        RECT -245.345 70.195 -245.065 70.475 ;
        RECT -246.465 67.435 -246.185 67.715 ;
        RECT -246.465 66.835 -246.185 67.115 ;
        RECT -244.225 67.435 -243.945 67.715 ;
        RECT -244.225 66.835 -243.945 67.115 ;
        RECT -234.145 77.515 -233.865 77.795 ;
        RECT -234.145 76.915 -233.865 77.195 ;
        RECT -238.625 74.155 -238.345 74.435 ;
        RECT -238.625 73.555 -238.345 73.835 ;
        RECT -240.865 70.795 -240.585 71.075 ;
        RECT -240.865 70.195 -240.585 70.475 ;
        RECT -241.985 67.435 -241.705 67.715 ;
        RECT -241.985 66.835 -241.705 67.115 ;
        RECT -239.745 67.435 -239.465 67.715 ;
        RECT -239.745 66.835 -239.465 67.115 ;
        RECT -236.385 70.795 -236.105 71.075 ;
        RECT -236.385 70.195 -236.105 70.475 ;
        RECT -237.505 67.435 -237.225 67.715 ;
        RECT -237.505 66.835 -237.225 67.115 ;
        RECT -235.265 67.435 -234.985 67.715 ;
        RECT -235.265 66.835 -234.985 67.115 ;
        RECT -229.665 74.155 -229.385 74.435 ;
        RECT -229.665 73.555 -229.385 73.835 ;
        RECT -231.905 70.795 -231.625 71.075 ;
        RECT -231.905 70.195 -231.625 70.475 ;
        RECT -233.025 67.435 -232.745 67.715 ;
        RECT -233.025 66.835 -232.745 67.115 ;
        RECT -230.785 67.435 -230.505 67.715 ;
        RECT -230.785 66.835 -230.505 67.115 ;
        RECT -227.425 70.795 -227.145 71.075 ;
        RECT -227.425 70.195 -227.145 70.475 ;
        RECT -228.545 67.435 -228.265 67.715 ;
        RECT -228.545 66.835 -228.265 67.115 ;
        RECT -226.305 67.435 -226.025 67.715 ;
        RECT -226.305 66.835 -226.025 67.115 ;
        RECT -207.265 80.875 -206.985 81.155 ;
        RECT -207.265 80.275 -206.985 80.555 ;
        RECT -216.225 77.515 -215.945 77.795 ;
        RECT -216.225 76.915 -215.945 77.195 ;
        RECT -220.705 74.155 -220.425 74.435 ;
        RECT -220.705 73.555 -220.425 73.835 ;
        RECT -222.945 70.795 -222.665 71.075 ;
        RECT -222.945 70.195 -222.665 70.475 ;
        RECT -224.065 67.435 -223.785 67.715 ;
        RECT -224.065 66.835 -223.785 67.115 ;
        RECT -221.825 67.435 -221.545 67.715 ;
        RECT -221.825 66.835 -221.545 67.115 ;
        RECT -218.465 70.795 -218.185 71.075 ;
        RECT -218.465 70.195 -218.185 70.475 ;
        RECT -219.585 67.435 -219.305 67.715 ;
        RECT -219.585 66.835 -219.305 67.115 ;
        RECT -217.345 67.435 -217.065 67.715 ;
        RECT -217.345 66.835 -217.065 67.115 ;
        RECT -211.745 74.155 -211.465 74.435 ;
        RECT -211.745 73.555 -211.465 73.835 ;
        RECT -213.985 70.795 -213.705 71.075 ;
        RECT -213.985 70.195 -213.705 70.475 ;
        RECT -215.105 67.435 -214.825 67.715 ;
        RECT -215.105 66.835 -214.825 67.115 ;
        RECT -212.865 67.435 -212.585 67.715 ;
        RECT -212.865 66.835 -212.585 67.115 ;
        RECT -209.505 70.795 -209.225 71.075 ;
        RECT -209.505 70.195 -209.225 70.475 ;
        RECT -210.625 67.435 -210.345 67.715 ;
        RECT -210.625 66.835 -210.345 67.115 ;
        RECT -208.385 67.435 -208.105 67.715 ;
        RECT -208.385 66.835 -208.105 67.115 ;
        RECT -198.305 77.515 -198.025 77.795 ;
        RECT -198.305 76.915 -198.025 77.195 ;
        RECT -202.785 74.155 -202.505 74.435 ;
        RECT -202.785 73.555 -202.505 73.835 ;
        RECT -205.025 70.795 -204.745 71.075 ;
        RECT -205.025 70.195 -204.745 70.475 ;
        RECT -206.145 67.435 -205.865 67.715 ;
        RECT -206.145 66.835 -205.865 67.115 ;
        RECT -203.905 67.435 -203.625 67.715 ;
        RECT -203.905 66.835 -203.625 67.115 ;
        RECT -200.545 70.795 -200.265 71.075 ;
        RECT -200.545 70.195 -200.265 70.475 ;
        RECT -201.665 67.435 -201.385 67.715 ;
        RECT -201.665 66.835 -201.385 67.115 ;
        RECT -199.425 67.435 -199.145 67.715 ;
        RECT -199.425 66.835 -199.145 67.115 ;
        RECT -193.825 74.155 -193.545 74.435 ;
        RECT -193.825 73.555 -193.545 73.835 ;
        RECT -196.065 70.795 -195.785 71.075 ;
        RECT -196.065 70.195 -195.785 70.475 ;
        RECT -197.185 67.435 -196.905 67.715 ;
        RECT -197.185 66.835 -196.905 67.115 ;
        RECT -194.945 67.435 -194.665 67.715 ;
        RECT -194.945 66.835 -194.665 67.115 ;
        RECT -191.585 70.795 -191.305 71.075 ;
        RECT -191.585 70.195 -191.305 70.475 ;
        RECT -192.705 67.435 -192.425 67.715 ;
        RECT -192.705 66.835 -192.425 67.115 ;
        RECT -190.465 67.435 -190.185 67.715 ;
        RECT -190.465 66.835 -190.185 67.115 ;
        RECT -188.225 94.315 -187.945 94.595 ;
        RECT -188.225 93.715 -187.945 93.995 ;
        RECT 121.025 94.015 121.825 94.295 ;
        RECT -44.865 90.955 -44.585 91.235 ;
        RECT -44.865 90.355 -44.585 90.635 ;
        RECT 121.025 90.655 121.825 90.935 ;
        RECT -116.545 87.595 -116.265 87.875 ;
        RECT -116.545 86.995 -116.265 87.275 ;
        RECT -152.385 84.235 -152.105 84.515 ;
        RECT -152.385 83.635 -152.105 83.915 ;
        RECT -170.305 80.875 -170.025 81.155 ;
        RECT -170.305 80.275 -170.025 80.555 ;
        RECT -179.265 77.515 -178.985 77.795 ;
        RECT -179.265 76.915 -178.985 77.195 ;
        RECT -183.745 74.155 -183.465 74.435 ;
        RECT -183.745 73.555 -183.465 73.835 ;
        RECT -185.985 70.795 -185.705 71.075 ;
        RECT -185.985 70.195 -185.705 70.475 ;
        RECT -187.105 67.435 -186.825 67.715 ;
        RECT -187.105 66.835 -186.825 67.115 ;
        RECT -184.865 67.435 -184.585 67.715 ;
        RECT -184.865 66.835 -184.585 67.115 ;
        RECT -181.505 70.795 -181.225 71.075 ;
        RECT -181.505 70.195 -181.225 70.475 ;
        RECT -182.625 67.435 -182.345 67.715 ;
        RECT -182.625 66.835 -182.345 67.115 ;
        RECT -180.385 67.435 -180.105 67.715 ;
        RECT -180.385 66.835 -180.105 67.115 ;
        RECT -174.785 74.155 -174.505 74.435 ;
        RECT -174.785 73.555 -174.505 73.835 ;
        RECT -177.025 70.795 -176.745 71.075 ;
        RECT -177.025 70.195 -176.745 70.475 ;
        RECT -178.145 67.435 -177.865 67.715 ;
        RECT -178.145 66.835 -177.865 67.115 ;
        RECT -175.905 67.435 -175.625 67.715 ;
        RECT -175.905 66.835 -175.625 67.115 ;
        RECT -172.545 70.795 -172.265 71.075 ;
        RECT -172.545 70.195 -172.265 70.475 ;
        RECT -173.665 67.435 -173.385 67.715 ;
        RECT -173.665 66.835 -173.385 67.115 ;
        RECT -171.425 67.435 -171.145 67.715 ;
        RECT -171.425 66.835 -171.145 67.115 ;
        RECT -161.345 77.515 -161.065 77.795 ;
        RECT -161.345 76.915 -161.065 77.195 ;
        RECT -165.825 74.155 -165.545 74.435 ;
        RECT -165.825 73.555 -165.545 73.835 ;
        RECT -168.065 70.795 -167.785 71.075 ;
        RECT -168.065 70.195 -167.785 70.475 ;
        RECT -169.185 67.435 -168.905 67.715 ;
        RECT -169.185 66.835 -168.905 67.115 ;
        RECT -166.945 67.435 -166.665 67.715 ;
        RECT -166.945 66.835 -166.665 67.115 ;
        RECT -163.585 70.795 -163.305 71.075 ;
        RECT -163.585 70.195 -163.305 70.475 ;
        RECT -164.705 67.435 -164.425 67.715 ;
        RECT -164.705 66.835 -164.425 67.115 ;
        RECT -162.465 67.435 -162.185 67.715 ;
        RECT -162.465 66.835 -162.185 67.115 ;
        RECT -156.865 74.155 -156.585 74.435 ;
        RECT -156.865 73.555 -156.585 73.835 ;
        RECT -159.105 70.795 -158.825 71.075 ;
        RECT -159.105 70.195 -158.825 70.475 ;
        RECT -160.225 67.435 -159.945 67.715 ;
        RECT -160.225 66.835 -159.945 67.115 ;
        RECT -157.985 67.435 -157.705 67.715 ;
        RECT -157.985 66.835 -157.705 67.115 ;
        RECT -154.625 70.795 -154.345 71.075 ;
        RECT -154.625 70.195 -154.345 70.475 ;
        RECT -155.745 67.435 -155.465 67.715 ;
        RECT -155.745 66.835 -155.465 67.115 ;
        RECT -153.505 67.435 -153.225 67.715 ;
        RECT -153.505 66.835 -153.225 67.115 ;
        RECT -134.465 80.875 -134.185 81.155 ;
        RECT -134.465 80.275 -134.185 80.555 ;
        RECT -143.425 77.515 -143.145 77.795 ;
        RECT -143.425 76.915 -143.145 77.195 ;
        RECT -147.905 74.155 -147.625 74.435 ;
        RECT -147.905 73.555 -147.625 73.835 ;
        RECT -150.145 70.795 -149.865 71.075 ;
        RECT -150.145 70.195 -149.865 70.475 ;
        RECT -151.265 67.435 -150.985 67.715 ;
        RECT -151.265 66.835 -150.985 67.115 ;
        RECT -149.025 67.435 -148.745 67.715 ;
        RECT -149.025 66.835 -148.745 67.115 ;
        RECT -145.665 70.795 -145.385 71.075 ;
        RECT -145.665 70.195 -145.385 70.475 ;
        RECT -146.785 67.435 -146.505 67.715 ;
        RECT -146.785 66.835 -146.505 67.115 ;
        RECT -144.545 67.435 -144.265 67.715 ;
        RECT -144.545 66.835 -144.265 67.115 ;
        RECT -138.945 74.155 -138.665 74.435 ;
        RECT -138.945 73.555 -138.665 73.835 ;
        RECT -141.185 70.795 -140.905 71.075 ;
        RECT -141.185 70.195 -140.905 70.475 ;
        RECT -142.305 67.435 -142.025 67.715 ;
        RECT -142.305 66.835 -142.025 67.115 ;
        RECT -140.065 67.435 -139.785 67.715 ;
        RECT -140.065 66.835 -139.785 67.115 ;
        RECT -136.705 70.795 -136.425 71.075 ;
        RECT -136.705 70.195 -136.425 70.475 ;
        RECT -137.825 67.435 -137.545 67.715 ;
        RECT -137.825 66.835 -137.545 67.115 ;
        RECT -135.585 67.435 -135.305 67.715 ;
        RECT -135.585 66.835 -135.305 67.115 ;
        RECT -125.505 77.515 -125.225 77.795 ;
        RECT -125.505 76.915 -125.225 77.195 ;
        RECT -129.985 74.155 -129.705 74.435 ;
        RECT -129.985 73.555 -129.705 73.835 ;
        RECT -132.225 70.795 -131.945 71.075 ;
        RECT -132.225 70.195 -131.945 70.475 ;
        RECT -133.345 67.435 -133.065 67.715 ;
        RECT -133.345 66.835 -133.065 67.115 ;
        RECT -131.105 67.435 -130.825 67.715 ;
        RECT -131.105 66.835 -130.825 67.115 ;
        RECT -127.745 70.795 -127.465 71.075 ;
        RECT -127.745 70.195 -127.465 70.475 ;
        RECT -128.865 67.435 -128.585 67.715 ;
        RECT -128.865 66.835 -128.585 67.115 ;
        RECT -126.625 67.435 -126.345 67.715 ;
        RECT -126.625 66.835 -126.345 67.115 ;
        RECT -121.025 74.155 -120.745 74.435 ;
        RECT -121.025 73.555 -120.745 73.835 ;
        RECT -123.265 70.795 -122.985 71.075 ;
        RECT -123.265 70.195 -122.985 70.475 ;
        RECT -124.385 67.435 -124.105 67.715 ;
        RECT -124.385 66.835 -124.105 67.115 ;
        RECT -122.145 67.435 -121.865 67.715 ;
        RECT -122.145 66.835 -121.865 67.115 ;
        RECT -118.785 70.795 -118.505 71.075 ;
        RECT -118.785 70.195 -118.505 70.475 ;
        RECT -119.905 67.435 -119.625 67.715 ;
        RECT -119.905 66.835 -119.625 67.115 ;
        RECT -117.665 67.435 -117.385 67.715 ;
        RECT -117.665 66.835 -117.385 67.115 ;
        RECT -80.705 84.235 -80.425 84.515 ;
        RECT -80.705 83.635 -80.425 83.915 ;
        RECT -98.625 80.875 -98.345 81.155 ;
        RECT -98.625 80.275 -98.345 80.555 ;
        RECT -107.585 77.515 -107.305 77.795 ;
        RECT -107.585 76.915 -107.305 77.195 ;
        RECT -112.065 74.155 -111.785 74.435 ;
        RECT -112.065 73.555 -111.785 73.835 ;
        RECT -114.305 70.795 -114.025 71.075 ;
        RECT -114.305 70.195 -114.025 70.475 ;
        RECT -115.425 67.435 -115.145 67.715 ;
        RECT -115.425 66.835 -115.145 67.115 ;
        RECT -113.185 67.435 -112.905 67.715 ;
        RECT -113.185 66.835 -112.905 67.115 ;
        RECT -109.825 70.795 -109.545 71.075 ;
        RECT -109.825 70.195 -109.545 70.475 ;
        RECT -110.945 67.435 -110.665 67.715 ;
        RECT -110.945 66.835 -110.665 67.115 ;
        RECT -108.705 67.435 -108.425 67.715 ;
        RECT -108.705 66.835 -108.425 67.115 ;
        RECT -103.105 74.155 -102.825 74.435 ;
        RECT -103.105 73.555 -102.825 73.835 ;
        RECT -105.345 70.795 -105.065 71.075 ;
        RECT -105.345 70.195 -105.065 70.475 ;
        RECT -106.465 67.435 -106.185 67.715 ;
        RECT -106.465 66.835 -106.185 67.115 ;
        RECT -104.225 67.435 -103.945 67.715 ;
        RECT -104.225 66.835 -103.945 67.115 ;
        RECT -100.865 70.795 -100.585 71.075 ;
        RECT -100.865 70.195 -100.585 70.475 ;
        RECT -101.985 67.435 -101.705 67.715 ;
        RECT -101.985 66.835 -101.705 67.115 ;
        RECT -99.745 67.435 -99.465 67.715 ;
        RECT -99.745 66.835 -99.465 67.115 ;
        RECT -89.665 77.515 -89.385 77.795 ;
        RECT -89.665 76.915 -89.385 77.195 ;
        RECT -94.145 74.155 -93.865 74.435 ;
        RECT -94.145 73.555 -93.865 73.835 ;
        RECT -96.385 70.795 -96.105 71.075 ;
        RECT -96.385 70.195 -96.105 70.475 ;
        RECT -97.505 67.435 -97.225 67.715 ;
        RECT -97.505 66.835 -97.225 67.115 ;
        RECT -95.265 67.435 -94.985 67.715 ;
        RECT -95.265 66.835 -94.985 67.115 ;
        RECT -91.905 70.795 -91.625 71.075 ;
        RECT -91.905 70.195 -91.625 70.475 ;
        RECT -93.025 67.435 -92.745 67.715 ;
        RECT -93.025 66.835 -92.745 67.115 ;
        RECT -90.785 67.435 -90.505 67.715 ;
        RECT -90.785 66.835 -90.505 67.115 ;
        RECT -85.185 74.155 -84.905 74.435 ;
        RECT -85.185 73.555 -84.905 73.835 ;
        RECT -87.425 70.795 -87.145 71.075 ;
        RECT -87.425 70.195 -87.145 70.475 ;
        RECT -88.545 67.435 -88.265 67.715 ;
        RECT -88.545 66.835 -88.265 67.115 ;
        RECT -86.305 67.435 -86.025 67.715 ;
        RECT -86.305 66.835 -86.025 67.115 ;
        RECT -82.945 70.795 -82.665 71.075 ;
        RECT -82.945 70.195 -82.665 70.475 ;
        RECT -84.065 67.435 -83.785 67.715 ;
        RECT -84.065 66.835 -83.785 67.115 ;
        RECT -81.825 67.435 -81.545 67.715 ;
        RECT -81.825 66.835 -81.545 67.115 ;
        RECT -62.785 80.875 -62.505 81.155 ;
        RECT -62.785 80.275 -62.505 80.555 ;
        RECT -71.745 77.515 -71.465 77.795 ;
        RECT -71.745 76.915 -71.465 77.195 ;
        RECT -76.225 74.155 -75.945 74.435 ;
        RECT -76.225 73.555 -75.945 73.835 ;
        RECT -78.465 70.795 -78.185 71.075 ;
        RECT -78.465 70.195 -78.185 70.475 ;
        RECT -79.585 67.435 -79.305 67.715 ;
        RECT -79.585 66.835 -79.305 67.115 ;
        RECT -77.345 67.435 -77.065 67.715 ;
        RECT -77.345 66.835 -77.065 67.115 ;
        RECT -73.985 70.795 -73.705 71.075 ;
        RECT -73.985 70.195 -73.705 70.475 ;
        RECT -75.105 67.435 -74.825 67.715 ;
        RECT -75.105 66.835 -74.825 67.115 ;
        RECT -72.865 67.435 -72.585 67.715 ;
        RECT -72.865 66.835 -72.585 67.115 ;
        RECT -67.265 74.155 -66.985 74.435 ;
        RECT -67.265 73.555 -66.985 73.835 ;
        RECT -69.505 70.795 -69.225 71.075 ;
        RECT -69.505 70.195 -69.225 70.475 ;
        RECT -70.625 67.435 -70.345 67.715 ;
        RECT -70.625 66.835 -70.345 67.115 ;
        RECT -68.385 67.435 -68.105 67.715 ;
        RECT -68.385 66.835 -68.105 67.115 ;
        RECT -65.025 70.795 -64.745 71.075 ;
        RECT -65.025 70.195 -64.745 70.475 ;
        RECT -66.145 67.435 -65.865 67.715 ;
        RECT -66.145 66.835 -65.865 67.115 ;
        RECT -63.905 67.435 -63.625 67.715 ;
        RECT -63.905 66.835 -63.625 67.115 ;
        RECT -53.825 77.515 -53.545 77.795 ;
        RECT -53.825 76.915 -53.545 77.195 ;
        RECT -58.305 74.155 -58.025 74.435 ;
        RECT -58.305 73.555 -58.025 73.835 ;
        RECT -60.545 70.795 -60.265 71.075 ;
        RECT -60.545 70.195 -60.265 70.475 ;
        RECT -61.665 67.435 -61.385 67.715 ;
        RECT -61.665 66.835 -61.385 67.115 ;
        RECT -59.425 67.435 -59.145 67.715 ;
        RECT -59.425 66.835 -59.145 67.115 ;
        RECT -56.065 70.795 -55.785 71.075 ;
        RECT -56.065 70.195 -55.785 70.475 ;
        RECT -57.185 67.435 -56.905 67.715 ;
        RECT -57.185 66.835 -56.905 67.115 ;
        RECT -54.945 67.435 -54.665 67.715 ;
        RECT -54.945 66.835 -54.665 67.115 ;
        RECT -49.345 74.155 -49.065 74.435 ;
        RECT -49.345 73.555 -49.065 73.835 ;
        RECT -51.585 70.795 -51.305 71.075 ;
        RECT -51.585 70.195 -51.305 70.475 ;
        RECT -52.705 67.435 -52.425 67.715 ;
        RECT -52.705 66.835 -52.425 67.115 ;
        RECT -50.465 67.435 -50.185 67.715 ;
        RECT -50.465 66.835 -50.185 67.115 ;
        RECT -47.105 70.795 -46.825 71.075 ;
        RECT -47.105 70.195 -46.825 70.475 ;
        RECT -48.225 67.435 -47.945 67.715 ;
        RECT -48.225 66.835 -47.945 67.115 ;
        RECT -45.985 67.435 -45.705 67.715 ;
        RECT -45.985 66.835 -45.705 67.115 ;
        RECT 26.815 87.595 27.095 87.875 ;
        RECT 26.815 86.995 27.095 87.275 ;
        RECT 121.025 87.295 121.825 87.575 ;
        RECT -9.025 84.235 -8.745 84.515 ;
        RECT -9.025 83.635 -8.745 83.915 ;
        RECT -26.945 80.875 -26.665 81.155 ;
        RECT -26.945 80.275 -26.665 80.555 ;
        RECT -35.905 77.515 -35.625 77.795 ;
        RECT -35.905 76.915 -35.625 77.195 ;
        RECT -40.385 74.155 -40.105 74.435 ;
        RECT -40.385 73.555 -40.105 73.835 ;
        RECT -42.625 70.795 -42.345 71.075 ;
        RECT -42.625 70.195 -42.345 70.475 ;
        RECT -43.745 67.435 -43.465 67.715 ;
        RECT -43.745 66.835 -43.465 67.115 ;
        RECT -41.505 67.435 -41.225 67.715 ;
        RECT -41.505 66.835 -41.225 67.115 ;
        RECT -38.145 70.795 -37.865 71.075 ;
        RECT -38.145 70.195 -37.865 70.475 ;
        RECT -39.265 67.435 -38.985 67.715 ;
        RECT -39.265 66.835 -38.985 67.115 ;
        RECT -37.025 67.435 -36.745 67.715 ;
        RECT -37.025 66.835 -36.745 67.115 ;
        RECT -31.425 74.155 -31.145 74.435 ;
        RECT -31.425 73.555 -31.145 73.835 ;
        RECT -33.665 70.795 -33.385 71.075 ;
        RECT -33.665 70.195 -33.385 70.475 ;
        RECT -34.785 67.435 -34.505 67.715 ;
        RECT -34.785 66.835 -34.505 67.115 ;
        RECT -32.545 67.435 -32.265 67.715 ;
        RECT -32.545 66.835 -32.265 67.115 ;
        RECT -29.185 70.795 -28.905 71.075 ;
        RECT -29.185 70.195 -28.905 70.475 ;
        RECT -30.305 67.435 -30.025 67.715 ;
        RECT -30.305 66.835 -30.025 67.115 ;
        RECT -28.065 67.435 -27.785 67.715 ;
        RECT -28.065 66.835 -27.785 67.115 ;
        RECT -17.985 77.515 -17.705 77.795 ;
        RECT -17.985 76.915 -17.705 77.195 ;
        RECT -22.465 74.155 -22.185 74.435 ;
        RECT -22.465 73.555 -22.185 73.835 ;
        RECT -24.705 70.795 -24.425 71.075 ;
        RECT -24.705 70.195 -24.425 70.475 ;
        RECT -25.825 67.435 -25.545 67.715 ;
        RECT -25.825 66.835 -25.545 67.115 ;
        RECT -23.585 67.435 -23.305 67.715 ;
        RECT -23.585 66.835 -23.305 67.115 ;
        RECT -20.225 70.795 -19.945 71.075 ;
        RECT -20.225 70.195 -19.945 70.475 ;
        RECT -21.345 67.435 -21.065 67.715 ;
        RECT -21.345 66.835 -21.065 67.115 ;
        RECT -19.105 67.435 -18.825 67.715 ;
        RECT -19.105 66.835 -18.825 67.115 ;
        RECT -13.505 74.155 -13.225 74.435 ;
        RECT -13.505 73.555 -13.225 73.835 ;
        RECT -15.745 70.795 -15.465 71.075 ;
        RECT -15.745 70.195 -15.465 70.475 ;
        RECT -16.865 67.435 -16.585 67.715 ;
        RECT -16.865 66.835 -16.585 67.115 ;
        RECT -14.625 67.435 -14.345 67.715 ;
        RECT -14.625 66.835 -14.345 67.115 ;
        RECT -11.265 70.795 -10.985 71.075 ;
        RECT -11.265 70.195 -10.985 70.475 ;
        RECT -12.385 67.435 -12.105 67.715 ;
        RECT -12.385 66.835 -12.105 67.115 ;
        RECT -10.145 67.435 -9.865 67.715 ;
        RECT -10.145 66.835 -9.865 67.115 ;
        RECT 8.895 80.875 9.175 81.155 ;
        RECT 8.895 80.275 9.175 80.555 ;
        RECT -0.065 77.515 0.215 77.795 ;
        RECT -0.065 76.915 0.215 77.195 ;
        RECT -4.545 74.155 -4.265 74.435 ;
        RECT -4.545 73.555 -4.265 73.835 ;
        RECT -6.785 70.795 -6.505 71.075 ;
        RECT -6.785 70.195 -6.505 70.475 ;
        RECT -7.905 67.435 -7.625 67.715 ;
        RECT -7.905 66.835 -7.625 67.115 ;
        RECT -5.665 67.435 -5.385 67.715 ;
        RECT -5.665 66.835 -5.385 67.115 ;
        RECT -2.305 70.795 -2.025 71.075 ;
        RECT -2.305 70.195 -2.025 70.475 ;
        RECT -3.425 67.435 -3.145 67.715 ;
        RECT -3.425 66.835 -3.145 67.115 ;
        RECT -1.185 67.435 -0.905 67.715 ;
        RECT -1.185 66.835 -0.905 67.115 ;
        RECT 4.415 74.155 4.695 74.435 ;
        RECT 4.415 73.555 4.695 73.835 ;
        RECT 2.175 70.795 2.455 71.075 ;
        RECT 2.175 70.195 2.455 70.475 ;
        RECT 1.055 67.435 1.335 67.715 ;
        RECT 1.055 66.835 1.335 67.115 ;
        RECT 3.295 67.435 3.575 67.715 ;
        RECT 3.295 66.835 3.575 67.115 ;
        RECT 6.655 70.795 6.935 71.075 ;
        RECT 6.655 70.195 6.935 70.475 ;
        RECT 5.535 67.435 5.815 67.715 ;
        RECT 5.535 66.835 5.815 67.115 ;
        RECT 7.775 67.435 8.055 67.715 ;
        RECT 7.775 66.835 8.055 67.115 ;
        RECT 17.855 77.515 18.135 77.795 ;
        RECT 17.855 76.915 18.135 77.195 ;
        RECT 13.375 74.155 13.655 74.435 ;
        RECT 13.375 73.555 13.655 73.835 ;
        RECT 11.135 70.795 11.415 71.075 ;
        RECT 11.135 70.195 11.415 70.475 ;
        RECT 10.015 67.435 10.295 67.715 ;
        RECT 10.015 66.835 10.295 67.115 ;
        RECT 12.255 67.435 12.535 67.715 ;
        RECT 12.255 66.835 12.535 67.115 ;
        RECT 15.615 70.795 15.895 71.075 ;
        RECT 15.615 70.195 15.895 70.475 ;
        RECT 14.495 67.435 14.775 67.715 ;
        RECT 14.495 66.835 14.775 67.115 ;
        RECT 16.735 67.435 17.015 67.715 ;
        RECT 16.735 66.835 17.015 67.115 ;
        RECT 22.335 74.155 22.615 74.435 ;
        RECT 22.335 73.555 22.615 73.835 ;
        RECT 20.095 70.795 20.375 71.075 ;
        RECT 20.095 70.195 20.375 70.475 ;
        RECT 18.975 67.435 19.255 67.715 ;
        RECT 18.975 66.835 19.255 67.115 ;
        RECT 21.215 67.435 21.495 67.715 ;
        RECT 21.215 66.835 21.495 67.115 ;
        RECT 24.575 70.795 24.855 71.075 ;
        RECT 24.575 70.195 24.855 70.475 ;
        RECT 23.455 67.435 23.735 67.715 ;
        RECT 23.455 66.835 23.735 67.115 ;
        RECT 25.695 67.435 25.975 67.715 ;
        RECT 25.695 66.835 25.975 67.115 ;
        RECT 62.655 84.235 62.935 84.515 ;
        RECT 62.655 83.635 62.935 83.915 ;
        RECT 121.025 83.935 121.825 84.215 ;
        RECT 44.735 80.875 45.015 81.155 ;
        RECT 44.735 80.275 45.015 80.555 ;
        RECT 35.775 77.515 36.055 77.795 ;
        RECT 35.775 76.915 36.055 77.195 ;
        RECT 31.295 74.155 31.575 74.435 ;
        RECT 31.295 73.555 31.575 73.835 ;
        RECT 29.055 70.795 29.335 71.075 ;
        RECT 29.055 70.195 29.335 70.475 ;
        RECT 27.935 67.435 28.215 67.715 ;
        RECT 27.935 66.835 28.215 67.115 ;
        RECT 30.175 67.435 30.455 67.715 ;
        RECT 30.175 66.835 30.455 67.115 ;
        RECT 33.535 70.795 33.815 71.075 ;
        RECT 33.535 70.195 33.815 70.475 ;
        RECT 32.415 67.435 32.695 67.715 ;
        RECT 32.415 66.835 32.695 67.115 ;
        RECT 34.655 67.435 34.935 67.715 ;
        RECT 34.655 66.835 34.935 67.115 ;
        RECT 40.255 74.155 40.535 74.435 ;
        RECT 40.255 73.555 40.535 73.835 ;
        RECT 38.015 70.795 38.295 71.075 ;
        RECT 38.015 70.195 38.295 70.475 ;
        RECT 36.895 67.435 37.175 67.715 ;
        RECT 36.895 66.835 37.175 67.115 ;
        RECT 39.135 67.435 39.415 67.715 ;
        RECT 39.135 66.835 39.415 67.115 ;
        RECT 42.495 70.795 42.775 71.075 ;
        RECT 42.495 70.195 42.775 70.475 ;
        RECT 41.375 67.435 41.655 67.715 ;
        RECT 41.375 66.835 41.655 67.115 ;
        RECT 43.615 67.435 43.895 67.715 ;
        RECT 43.615 66.835 43.895 67.115 ;
        RECT 53.695 77.515 53.975 77.795 ;
        RECT 53.695 76.915 53.975 77.195 ;
        RECT 49.215 74.155 49.495 74.435 ;
        RECT 49.215 73.555 49.495 73.835 ;
        RECT 46.975 70.795 47.255 71.075 ;
        RECT 46.975 70.195 47.255 70.475 ;
        RECT 45.855 67.435 46.135 67.715 ;
        RECT 45.855 66.835 46.135 67.115 ;
        RECT 48.095 67.435 48.375 67.715 ;
        RECT 48.095 66.835 48.375 67.115 ;
        RECT 51.455 70.795 51.735 71.075 ;
        RECT 51.455 70.195 51.735 70.475 ;
        RECT 50.335 67.435 50.615 67.715 ;
        RECT 50.335 66.835 50.615 67.115 ;
        RECT 52.575 67.435 52.855 67.715 ;
        RECT 52.575 66.835 52.855 67.115 ;
        RECT 58.175 74.155 58.455 74.435 ;
        RECT 58.175 73.555 58.455 73.835 ;
        RECT 55.935 70.795 56.215 71.075 ;
        RECT 55.935 70.195 56.215 70.475 ;
        RECT 54.815 67.435 55.095 67.715 ;
        RECT 54.815 66.835 55.095 67.115 ;
        RECT 57.055 67.435 57.335 67.715 ;
        RECT 57.055 66.835 57.335 67.115 ;
        RECT 60.415 70.795 60.695 71.075 ;
        RECT 60.415 70.195 60.695 70.475 ;
        RECT 59.295 67.435 59.575 67.715 ;
        RECT 59.295 66.835 59.575 67.115 ;
        RECT 61.535 67.435 61.815 67.715 ;
        RECT 61.535 66.835 61.815 67.115 ;
        RECT 80.575 80.875 80.855 81.155 ;
        RECT 80.575 80.275 80.855 80.555 ;
        RECT 121.025 80.575 121.825 80.855 ;
        RECT 71.615 77.515 71.895 77.795 ;
        RECT 71.615 76.915 71.895 77.195 ;
        RECT 67.135 74.155 67.415 74.435 ;
        RECT 67.135 73.555 67.415 73.835 ;
        RECT 64.895 70.795 65.175 71.075 ;
        RECT 64.895 70.195 65.175 70.475 ;
        RECT 63.775 67.435 64.055 67.715 ;
        RECT 63.775 66.835 64.055 67.115 ;
        RECT 66.015 67.435 66.295 67.715 ;
        RECT 66.015 66.835 66.295 67.115 ;
        RECT 69.375 70.795 69.655 71.075 ;
        RECT 69.375 70.195 69.655 70.475 ;
        RECT 68.255 67.435 68.535 67.715 ;
        RECT 68.255 66.835 68.535 67.115 ;
        RECT 70.495 67.435 70.775 67.715 ;
        RECT 70.495 66.835 70.775 67.115 ;
        RECT 76.095 74.155 76.375 74.435 ;
        RECT 76.095 73.555 76.375 73.835 ;
        RECT 73.855 70.795 74.135 71.075 ;
        RECT 73.855 70.195 74.135 70.475 ;
        RECT 72.735 67.435 73.015 67.715 ;
        RECT 72.735 66.835 73.015 67.115 ;
        RECT 74.975 67.435 75.255 67.715 ;
        RECT 74.975 66.835 75.255 67.115 ;
        RECT 78.335 70.795 78.615 71.075 ;
        RECT 78.335 70.195 78.615 70.475 ;
        RECT 77.215 67.435 77.495 67.715 ;
        RECT 77.215 66.835 77.495 67.115 ;
        RECT 79.455 67.435 79.735 67.715 ;
        RECT 79.455 66.835 79.735 67.115 ;
        RECT 89.535 77.515 89.815 77.795 ;
        RECT 89.535 76.915 89.815 77.195 ;
        RECT 121.025 77.215 121.825 77.495 ;
        RECT 85.055 74.155 85.335 74.435 ;
        RECT 85.055 73.555 85.335 73.835 ;
        RECT 82.815 70.795 83.095 71.075 ;
        RECT 82.815 70.195 83.095 70.475 ;
        RECT 81.695 67.435 81.975 67.715 ;
        RECT 81.695 66.835 81.975 67.115 ;
        RECT 83.935 67.435 84.215 67.715 ;
        RECT 83.935 66.835 84.215 67.115 ;
        RECT 87.295 70.795 87.575 71.075 ;
        RECT 87.295 70.195 87.575 70.475 ;
        RECT 86.175 67.435 86.455 67.715 ;
        RECT 86.175 66.835 86.455 67.115 ;
        RECT 88.415 67.435 88.695 67.715 ;
        RECT 88.415 66.835 88.695 67.115 ;
        RECT 94.015 74.155 94.295 74.435 ;
        RECT 94.015 73.555 94.295 73.835 ;
        RECT 121.025 73.855 121.825 74.135 ;
        RECT 91.775 70.795 92.055 71.075 ;
        RECT 91.775 70.195 92.055 70.475 ;
        RECT 90.655 67.435 90.935 67.715 ;
        RECT 90.655 66.835 90.935 67.115 ;
        RECT 92.895 67.435 93.175 67.715 ;
        RECT 92.895 66.835 93.175 67.115 ;
        RECT 96.255 70.795 96.535 71.075 ;
        RECT 96.255 70.195 96.535 70.475 ;
        RECT 121.025 70.495 121.825 70.775 ;
        RECT 95.135 67.435 95.415 67.715 ;
        RECT 95.135 66.835 95.415 67.115 ;
        RECT 97.375 67.435 97.655 67.715 ;
        RECT 97.375 66.835 97.655 67.115 ;
        RECT 121.025 67.135 121.825 67.415 ;
        RECT 121.025 63.775 121.825 64.055 ;
        RECT -474.945 44.575 -474.665 44.855 ;
        RECT -474.945 43.975 -474.665 44.255 ;
        RECT -472.705 44.575 -472.425 44.855 ;
        RECT -472.705 43.975 -472.425 44.255 ;
        RECT -473.825 41.215 -473.545 41.495 ;
        RECT -473.825 40.615 -473.545 40.895 ;
        RECT -470.465 44.575 -470.185 44.855 ;
        RECT -470.465 43.975 -470.185 44.255 ;
        RECT -468.225 44.575 -467.945 44.855 ;
        RECT -468.225 43.975 -467.945 44.255 ;
        RECT -469.345 41.215 -469.065 41.495 ;
        RECT -469.345 40.615 -469.065 40.895 ;
        RECT -471.585 37.855 -471.305 38.135 ;
        RECT -471.585 37.255 -471.305 37.535 ;
        RECT -465.985 44.575 -465.705 44.855 ;
        RECT -465.985 43.975 -465.705 44.255 ;
        RECT -463.745 44.575 -463.465 44.855 ;
        RECT -463.745 43.975 -463.465 44.255 ;
        RECT -464.865 41.215 -464.585 41.495 ;
        RECT -464.865 40.615 -464.585 40.895 ;
        RECT -461.505 44.575 -461.225 44.855 ;
        RECT -461.505 43.975 -461.225 44.255 ;
        RECT -459.265 44.575 -458.985 44.855 ;
        RECT -459.265 43.975 -458.985 44.255 ;
        RECT -460.385 41.215 -460.105 41.495 ;
        RECT -460.385 40.615 -460.105 40.895 ;
        RECT -462.625 37.855 -462.345 38.135 ;
        RECT -462.625 37.255 -462.345 37.535 ;
        RECT -467.105 34.495 -466.825 34.775 ;
        RECT -467.105 33.895 -466.825 34.175 ;
        RECT -457.025 44.575 -456.745 44.855 ;
        RECT -457.025 43.975 -456.745 44.255 ;
        RECT -454.785 44.575 -454.505 44.855 ;
        RECT -454.785 43.975 -454.505 44.255 ;
        RECT -455.905 41.215 -455.625 41.495 ;
        RECT -455.905 40.615 -455.625 40.895 ;
        RECT -452.545 44.575 -452.265 44.855 ;
        RECT -452.545 43.975 -452.265 44.255 ;
        RECT -450.305 44.575 -450.025 44.855 ;
        RECT -450.305 43.975 -450.025 44.255 ;
        RECT -451.425 41.215 -451.145 41.495 ;
        RECT -451.425 40.615 -451.145 40.895 ;
        RECT -453.665 37.855 -453.385 38.135 ;
        RECT -453.665 37.255 -453.385 37.535 ;
        RECT -448.065 44.575 -447.785 44.855 ;
        RECT -448.065 43.975 -447.785 44.255 ;
        RECT -445.825 44.575 -445.545 44.855 ;
        RECT -445.825 43.975 -445.545 44.255 ;
        RECT -446.945 41.215 -446.665 41.495 ;
        RECT -446.945 40.615 -446.665 40.895 ;
        RECT -443.585 44.575 -443.305 44.855 ;
        RECT -443.585 43.975 -443.305 44.255 ;
        RECT -441.345 44.575 -441.065 44.855 ;
        RECT -441.345 43.975 -441.065 44.255 ;
        RECT -442.465 41.215 -442.185 41.495 ;
        RECT -442.465 40.615 -442.185 40.895 ;
        RECT -444.705 37.855 -444.425 38.135 ;
        RECT -444.705 37.255 -444.425 37.535 ;
        RECT -449.185 34.495 -448.905 34.775 ;
        RECT -449.185 33.895 -448.905 34.175 ;
        RECT -458.145 31.135 -457.865 31.415 ;
        RECT -458.145 30.535 -457.865 30.815 ;
        RECT -439.105 44.575 -438.825 44.855 ;
        RECT -439.105 43.975 -438.825 44.255 ;
        RECT -436.865 44.575 -436.585 44.855 ;
        RECT -436.865 43.975 -436.585 44.255 ;
        RECT -437.985 41.215 -437.705 41.495 ;
        RECT -437.985 40.615 -437.705 40.895 ;
        RECT -434.625 44.575 -434.345 44.855 ;
        RECT -434.625 43.975 -434.345 44.255 ;
        RECT -432.385 44.575 -432.105 44.855 ;
        RECT -432.385 43.975 -432.105 44.255 ;
        RECT -433.505 41.215 -433.225 41.495 ;
        RECT -433.505 40.615 -433.225 40.895 ;
        RECT -435.745 37.855 -435.465 38.135 ;
        RECT -435.745 37.255 -435.465 37.535 ;
        RECT -430.145 44.575 -429.865 44.855 ;
        RECT -430.145 43.975 -429.865 44.255 ;
        RECT -427.905 44.575 -427.625 44.855 ;
        RECT -427.905 43.975 -427.625 44.255 ;
        RECT -429.025 41.215 -428.745 41.495 ;
        RECT -429.025 40.615 -428.745 40.895 ;
        RECT -425.665 44.575 -425.385 44.855 ;
        RECT -425.665 43.975 -425.385 44.255 ;
        RECT -423.425 44.575 -423.145 44.855 ;
        RECT -423.425 43.975 -423.145 44.255 ;
        RECT -424.545 41.215 -424.265 41.495 ;
        RECT -424.545 40.615 -424.265 40.895 ;
        RECT -426.785 37.855 -426.505 38.135 ;
        RECT -426.785 37.255 -426.505 37.535 ;
        RECT -431.265 34.495 -430.985 34.775 ;
        RECT -431.265 33.895 -430.985 34.175 ;
        RECT -421.185 44.575 -420.905 44.855 ;
        RECT -421.185 43.975 -420.905 44.255 ;
        RECT -418.945 44.575 -418.665 44.855 ;
        RECT -418.945 43.975 -418.665 44.255 ;
        RECT -420.065 41.215 -419.785 41.495 ;
        RECT -420.065 40.615 -419.785 40.895 ;
        RECT -416.705 44.575 -416.425 44.855 ;
        RECT -416.705 43.975 -416.425 44.255 ;
        RECT -414.465 44.575 -414.185 44.855 ;
        RECT -414.465 43.975 -414.185 44.255 ;
        RECT -415.585 41.215 -415.305 41.495 ;
        RECT -415.585 40.615 -415.305 40.895 ;
        RECT -417.825 37.855 -417.545 38.135 ;
        RECT -417.825 37.255 -417.545 37.535 ;
        RECT -412.225 44.575 -411.945 44.855 ;
        RECT -412.225 43.975 -411.945 44.255 ;
        RECT -409.985 44.575 -409.705 44.855 ;
        RECT -409.985 43.975 -409.705 44.255 ;
        RECT -411.105 41.215 -410.825 41.495 ;
        RECT -411.105 40.615 -410.825 40.895 ;
        RECT -407.745 44.575 -407.465 44.855 ;
        RECT -407.745 43.975 -407.465 44.255 ;
        RECT -405.505 44.575 -405.225 44.855 ;
        RECT -405.505 43.975 -405.225 44.255 ;
        RECT -406.625 41.215 -406.345 41.495 ;
        RECT -406.625 40.615 -406.345 40.895 ;
        RECT -408.865 37.855 -408.585 38.135 ;
        RECT -408.865 37.255 -408.585 37.535 ;
        RECT -413.345 34.495 -413.065 34.775 ;
        RECT -413.345 33.895 -413.065 34.175 ;
        RECT -422.305 31.135 -422.025 31.415 ;
        RECT -422.305 30.535 -422.025 30.815 ;
        RECT -440.225 27.775 -439.945 28.055 ;
        RECT -440.225 27.175 -439.945 27.455 ;
        RECT -403.265 44.575 -402.985 44.855 ;
        RECT -403.265 43.975 -402.985 44.255 ;
        RECT -401.025 44.575 -400.745 44.855 ;
        RECT -401.025 43.975 -400.745 44.255 ;
        RECT -402.145 41.215 -401.865 41.495 ;
        RECT -402.145 40.615 -401.865 40.895 ;
        RECT -398.785 44.575 -398.505 44.855 ;
        RECT -398.785 43.975 -398.505 44.255 ;
        RECT -396.545 44.575 -396.265 44.855 ;
        RECT -396.545 43.975 -396.265 44.255 ;
        RECT -397.665 41.215 -397.385 41.495 ;
        RECT -397.665 40.615 -397.385 40.895 ;
        RECT -399.905 37.855 -399.625 38.135 ;
        RECT -399.905 37.255 -399.625 37.535 ;
        RECT -394.305 44.575 -394.025 44.855 ;
        RECT -394.305 43.975 -394.025 44.255 ;
        RECT -392.065 44.575 -391.785 44.855 ;
        RECT -392.065 43.975 -391.785 44.255 ;
        RECT -393.185 41.215 -392.905 41.495 ;
        RECT -393.185 40.615 -392.905 40.895 ;
        RECT -389.825 44.575 -389.545 44.855 ;
        RECT -389.825 43.975 -389.545 44.255 ;
        RECT -387.585 44.575 -387.305 44.855 ;
        RECT -387.585 43.975 -387.305 44.255 ;
        RECT -388.705 41.215 -388.425 41.495 ;
        RECT -388.705 40.615 -388.425 40.895 ;
        RECT -390.945 37.855 -390.665 38.135 ;
        RECT -390.945 37.255 -390.665 37.535 ;
        RECT -395.425 34.495 -395.145 34.775 ;
        RECT -395.425 33.895 -395.145 34.175 ;
        RECT -385.345 44.575 -385.065 44.855 ;
        RECT -385.345 43.975 -385.065 44.255 ;
        RECT -383.105 44.575 -382.825 44.855 ;
        RECT -383.105 43.975 -382.825 44.255 ;
        RECT -384.225 41.215 -383.945 41.495 ;
        RECT -384.225 40.615 -383.945 40.895 ;
        RECT -380.865 44.575 -380.585 44.855 ;
        RECT -380.865 43.975 -380.585 44.255 ;
        RECT -378.625 44.575 -378.345 44.855 ;
        RECT -378.625 43.975 -378.345 44.255 ;
        RECT -379.745 41.215 -379.465 41.495 ;
        RECT -379.745 40.615 -379.465 40.895 ;
        RECT -381.985 37.855 -381.705 38.135 ;
        RECT -381.985 37.255 -381.705 37.535 ;
        RECT -376.385 44.575 -376.105 44.855 ;
        RECT -376.385 43.975 -376.105 44.255 ;
        RECT -374.145 44.575 -373.865 44.855 ;
        RECT -374.145 43.975 -373.865 44.255 ;
        RECT -375.265 41.215 -374.985 41.495 ;
        RECT -375.265 40.615 -374.985 40.895 ;
        RECT -371.905 44.575 -371.625 44.855 ;
        RECT -371.905 43.975 -371.625 44.255 ;
        RECT -369.665 44.575 -369.385 44.855 ;
        RECT -369.665 43.975 -369.385 44.255 ;
        RECT -370.785 41.215 -370.505 41.495 ;
        RECT -370.785 40.615 -370.505 40.895 ;
        RECT -373.025 37.855 -372.745 38.135 ;
        RECT -373.025 37.255 -372.745 37.535 ;
        RECT -377.505 34.495 -377.225 34.775 ;
        RECT -377.505 33.895 -377.225 34.175 ;
        RECT -386.465 31.135 -386.185 31.415 ;
        RECT -386.465 30.535 -386.185 30.815 ;
        RECT -367.425 44.575 -367.145 44.855 ;
        RECT -367.425 43.975 -367.145 44.255 ;
        RECT -365.185 44.575 -364.905 44.855 ;
        RECT -365.185 43.975 -364.905 44.255 ;
        RECT -366.305 41.215 -366.025 41.495 ;
        RECT -366.305 40.615 -366.025 40.895 ;
        RECT -362.945 44.575 -362.665 44.855 ;
        RECT -362.945 43.975 -362.665 44.255 ;
        RECT -360.705 44.575 -360.425 44.855 ;
        RECT -360.705 43.975 -360.425 44.255 ;
        RECT -361.825 41.215 -361.545 41.495 ;
        RECT -361.825 40.615 -361.545 40.895 ;
        RECT -364.065 37.855 -363.785 38.135 ;
        RECT -364.065 37.255 -363.785 37.535 ;
        RECT -358.465 44.575 -358.185 44.855 ;
        RECT -358.465 43.975 -358.185 44.255 ;
        RECT -356.225 44.575 -355.945 44.855 ;
        RECT -356.225 43.975 -355.945 44.255 ;
        RECT -357.345 41.215 -357.065 41.495 ;
        RECT -357.345 40.615 -357.065 40.895 ;
        RECT -353.985 44.575 -353.705 44.855 ;
        RECT -353.985 43.975 -353.705 44.255 ;
        RECT -351.745 44.575 -351.465 44.855 ;
        RECT -351.745 43.975 -351.465 44.255 ;
        RECT -352.865 41.215 -352.585 41.495 ;
        RECT -352.865 40.615 -352.585 40.895 ;
        RECT -355.105 37.855 -354.825 38.135 ;
        RECT -355.105 37.255 -354.825 37.535 ;
        RECT -359.585 34.495 -359.305 34.775 ;
        RECT -359.585 33.895 -359.305 34.175 ;
        RECT -349.505 44.575 -349.225 44.855 ;
        RECT -349.505 43.975 -349.225 44.255 ;
        RECT -347.265 44.575 -346.985 44.855 ;
        RECT -347.265 43.975 -346.985 44.255 ;
        RECT -348.385 41.215 -348.105 41.495 ;
        RECT -348.385 40.615 -348.105 40.895 ;
        RECT -345.025 44.575 -344.745 44.855 ;
        RECT -345.025 43.975 -344.745 44.255 ;
        RECT -342.785 44.575 -342.505 44.855 ;
        RECT -342.785 43.975 -342.505 44.255 ;
        RECT -343.905 41.215 -343.625 41.495 ;
        RECT -343.905 40.615 -343.625 40.895 ;
        RECT -346.145 37.855 -345.865 38.135 ;
        RECT -346.145 37.255 -345.865 37.535 ;
        RECT -340.545 44.575 -340.265 44.855 ;
        RECT -340.545 43.975 -340.265 44.255 ;
        RECT -338.305 44.575 -338.025 44.855 ;
        RECT -338.305 43.975 -338.025 44.255 ;
        RECT -339.425 41.215 -339.145 41.495 ;
        RECT -339.425 40.615 -339.145 40.895 ;
        RECT -336.065 44.575 -335.785 44.855 ;
        RECT -336.065 43.975 -335.785 44.255 ;
        RECT -333.825 44.575 -333.545 44.855 ;
        RECT -333.825 43.975 -333.545 44.255 ;
        RECT -334.945 41.215 -334.665 41.495 ;
        RECT -334.945 40.615 -334.665 40.895 ;
        RECT -337.185 37.855 -336.905 38.135 ;
        RECT -337.185 37.255 -336.905 37.535 ;
        RECT -341.665 34.495 -341.385 34.775 ;
        RECT -341.665 33.895 -341.385 34.175 ;
        RECT -350.625 31.135 -350.345 31.415 ;
        RECT -350.625 30.535 -350.345 30.815 ;
        RECT -368.545 27.775 -368.265 28.055 ;
        RECT -368.545 27.175 -368.265 27.455 ;
        RECT -404.385 24.415 -404.105 24.695 ;
        RECT -404.385 23.815 -404.105 24.095 ;
        RECT -331.585 44.575 -331.305 44.855 ;
        RECT -331.585 43.975 -331.305 44.255 ;
        RECT -329.345 44.575 -329.065 44.855 ;
        RECT -329.345 43.975 -329.065 44.255 ;
        RECT -330.465 41.215 -330.185 41.495 ;
        RECT -330.465 40.615 -330.185 40.895 ;
        RECT -327.105 44.575 -326.825 44.855 ;
        RECT -327.105 43.975 -326.825 44.255 ;
        RECT -324.865 44.575 -324.585 44.855 ;
        RECT -324.865 43.975 -324.585 44.255 ;
        RECT -325.985 41.215 -325.705 41.495 ;
        RECT -325.985 40.615 -325.705 40.895 ;
        RECT -328.225 37.855 -327.945 38.135 ;
        RECT -328.225 37.255 -327.945 37.535 ;
        RECT -322.625 44.575 -322.345 44.855 ;
        RECT -322.625 43.975 -322.345 44.255 ;
        RECT -320.385 44.575 -320.105 44.855 ;
        RECT -320.385 43.975 -320.105 44.255 ;
        RECT -321.505 41.215 -321.225 41.495 ;
        RECT -321.505 40.615 -321.225 40.895 ;
        RECT -318.145 44.575 -317.865 44.855 ;
        RECT -318.145 43.975 -317.865 44.255 ;
        RECT -315.905 44.575 -315.625 44.855 ;
        RECT -315.905 43.975 -315.625 44.255 ;
        RECT -317.025 41.215 -316.745 41.495 ;
        RECT -317.025 40.615 -316.745 40.895 ;
        RECT -319.265 37.855 -318.985 38.135 ;
        RECT -319.265 37.255 -318.985 37.535 ;
        RECT -323.745 34.495 -323.465 34.775 ;
        RECT -323.745 33.895 -323.465 34.175 ;
        RECT -313.665 44.575 -313.385 44.855 ;
        RECT -313.665 43.975 -313.385 44.255 ;
        RECT -311.425 44.575 -311.145 44.855 ;
        RECT -311.425 43.975 -311.145 44.255 ;
        RECT -312.545 41.215 -312.265 41.495 ;
        RECT -312.545 40.615 -312.265 40.895 ;
        RECT -309.185 44.575 -308.905 44.855 ;
        RECT -309.185 43.975 -308.905 44.255 ;
        RECT -306.945 44.575 -306.665 44.855 ;
        RECT -306.945 43.975 -306.665 44.255 ;
        RECT -308.065 41.215 -307.785 41.495 ;
        RECT -308.065 40.615 -307.785 40.895 ;
        RECT -310.305 37.855 -310.025 38.135 ;
        RECT -310.305 37.255 -310.025 37.535 ;
        RECT -304.705 44.575 -304.425 44.855 ;
        RECT -304.705 43.975 -304.425 44.255 ;
        RECT -302.465 44.575 -302.185 44.855 ;
        RECT -302.465 43.975 -302.185 44.255 ;
        RECT -303.585 41.215 -303.305 41.495 ;
        RECT -303.585 40.615 -303.305 40.895 ;
        RECT -300.225 44.575 -299.945 44.855 ;
        RECT -300.225 43.975 -299.945 44.255 ;
        RECT -297.985 44.575 -297.705 44.855 ;
        RECT -297.985 43.975 -297.705 44.255 ;
        RECT -299.105 41.215 -298.825 41.495 ;
        RECT -299.105 40.615 -298.825 40.895 ;
        RECT -301.345 37.855 -301.065 38.135 ;
        RECT -301.345 37.255 -301.065 37.535 ;
        RECT -305.825 34.495 -305.545 34.775 ;
        RECT -305.825 33.895 -305.545 34.175 ;
        RECT -314.785 31.135 -314.505 31.415 ;
        RECT -314.785 30.535 -314.505 30.815 ;
        RECT -295.745 44.575 -295.465 44.855 ;
        RECT -295.745 43.975 -295.465 44.255 ;
        RECT -293.505 44.575 -293.225 44.855 ;
        RECT -293.505 43.975 -293.225 44.255 ;
        RECT -294.625 41.215 -294.345 41.495 ;
        RECT -294.625 40.615 -294.345 40.895 ;
        RECT -291.265 44.575 -290.985 44.855 ;
        RECT -291.265 43.975 -290.985 44.255 ;
        RECT -289.025 44.575 -288.745 44.855 ;
        RECT -289.025 43.975 -288.745 44.255 ;
        RECT -290.145 41.215 -289.865 41.495 ;
        RECT -290.145 40.615 -289.865 40.895 ;
        RECT -292.385 37.855 -292.105 38.135 ;
        RECT -292.385 37.255 -292.105 37.535 ;
        RECT -286.785 44.575 -286.505 44.855 ;
        RECT -286.785 43.975 -286.505 44.255 ;
        RECT -284.545 44.575 -284.265 44.855 ;
        RECT -284.545 43.975 -284.265 44.255 ;
        RECT -285.665 41.215 -285.385 41.495 ;
        RECT -285.665 40.615 -285.385 40.895 ;
        RECT -282.305 44.575 -282.025 44.855 ;
        RECT -282.305 43.975 -282.025 44.255 ;
        RECT -280.065 44.575 -279.785 44.855 ;
        RECT -280.065 43.975 -279.785 44.255 ;
        RECT -281.185 41.215 -280.905 41.495 ;
        RECT -281.185 40.615 -280.905 40.895 ;
        RECT -283.425 37.855 -283.145 38.135 ;
        RECT -283.425 37.255 -283.145 37.535 ;
        RECT -287.905 34.495 -287.625 34.775 ;
        RECT -287.905 33.895 -287.625 34.175 ;
        RECT -277.825 44.575 -277.545 44.855 ;
        RECT -277.825 43.975 -277.545 44.255 ;
        RECT -275.585 44.575 -275.305 44.855 ;
        RECT -275.585 43.975 -275.305 44.255 ;
        RECT -276.705 41.215 -276.425 41.495 ;
        RECT -276.705 40.615 -276.425 40.895 ;
        RECT -273.345 44.575 -273.065 44.855 ;
        RECT -273.345 43.975 -273.065 44.255 ;
        RECT -271.105 44.575 -270.825 44.855 ;
        RECT -271.105 43.975 -270.825 44.255 ;
        RECT -272.225 41.215 -271.945 41.495 ;
        RECT -272.225 40.615 -271.945 40.895 ;
        RECT -274.465 37.855 -274.185 38.135 ;
        RECT -274.465 37.255 -274.185 37.535 ;
        RECT -268.865 44.575 -268.585 44.855 ;
        RECT -268.865 43.975 -268.585 44.255 ;
        RECT -266.625 44.575 -266.345 44.855 ;
        RECT -266.625 43.975 -266.345 44.255 ;
        RECT -267.745 41.215 -267.465 41.495 ;
        RECT -267.745 40.615 -267.465 40.895 ;
        RECT -264.385 44.575 -264.105 44.855 ;
        RECT -264.385 43.975 -264.105 44.255 ;
        RECT -262.145 44.575 -261.865 44.855 ;
        RECT -262.145 43.975 -261.865 44.255 ;
        RECT -263.265 41.215 -262.985 41.495 ;
        RECT -263.265 40.615 -262.985 40.895 ;
        RECT -265.505 37.855 -265.225 38.135 ;
        RECT -265.505 37.255 -265.225 37.535 ;
        RECT -269.985 34.495 -269.705 34.775 ;
        RECT -269.985 33.895 -269.705 34.175 ;
        RECT -278.945 31.135 -278.665 31.415 ;
        RECT -278.945 30.535 -278.665 30.815 ;
        RECT -296.865 27.775 -296.585 28.055 ;
        RECT -296.865 27.175 -296.585 27.455 ;
        RECT -259.905 44.575 -259.625 44.855 ;
        RECT -259.905 43.975 -259.625 44.255 ;
        RECT -257.665 44.575 -257.385 44.855 ;
        RECT -257.665 43.975 -257.385 44.255 ;
        RECT -258.785 41.215 -258.505 41.495 ;
        RECT -258.785 40.615 -258.505 40.895 ;
        RECT -255.425 44.575 -255.145 44.855 ;
        RECT -255.425 43.975 -255.145 44.255 ;
        RECT -253.185 44.575 -252.905 44.855 ;
        RECT -253.185 43.975 -252.905 44.255 ;
        RECT -254.305 41.215 -254.025 41.495 ;
        RECT -254.305 40.615 -254.025 40.895 ;
        RECT -256.545 37.855 -256.265 38.135 ;
        RECT -256.545 37.255 -256.265 37.535 ;
        RECT -250.945 44.575 -250.665 44.855 ;
        RECT -250.945 43.975 -250.665 44.255 ;
        RECT -248.705 44.575 -248.425 44.855 ;
        RECT -248.705 43.975 -248.425 44.255 ;
        RECT -249.825 41.215 -249.545 41.495 ;
        RECT -249.825 40.615 -249.545 40.895 ;
        RECT -246.465 44.575 -246.185 44.855 ;
        RECT -246.465 43.975 -246.185 44.255 ;
        RECT -244.225 44.575 -243.945 44.855 ;
        RECT -244.225 43.975 -243.945 44.255 ;
        RECT -245.345 41.215 -245.065 41.495 ;
        RECT -245.345 40.615 -245.065 40.895 ;
        RECT -247.585 37.855 -247.305 38.135 ;
        RECT -247.585 37.255 -247.305 37.535 ;
        RECT -252.065 34.495 -251.785 34.775 ;
        RECT -252.065 33.895 -251.785 34.175 ;
        RECT -241.985 44.575 -241.705 44.855 ;
        RECT -241.985 43.975 -241.705 44.255 ;
        RECT -239.745 44.575 -239.465 44.855 ;
        RECT -239.745 43.975 -239.465 44.255 ;
        RECT -240.865 41.215 -240.585 41.495 ;
        RECT -240.865 40.615 -240.585 40.895 ;
        RECT -237.505 44.575 -237.225 44.855 ;
        RECT -237.505 43.975 -237.225 44.255 ;
        RECT -235.265 44.575 -234.985 44.855 ;
        RECT -235.265 43.975 -234.985 44.255 ;
        RECT -236.385 41.215 -236.105 41.495 ;
        RECT -236.385 40.615 -236.105 40.895 ;
        RECT -238.625 37.855 -238.345 38.135 ;
        RECT -238.625 37.255 -238.345 37.535 ;
        RECT -233.025 44.575 -232.745 44.855 ;
        RECT -233.025 43.975 -232.745 44.255 ;
        RECT -230.785 44.575 -230.505 44.855 ;
        RECT -230.785 43.975 -230.505 44.255 ;
        RECT -231.905 41.215 -231.625 41.495 ;
        RECT -231.905 40.615 -231.625 40.895 ;
        RECT -228.545 44.575 -228.265 44.855 ;
        RECT -228.545 43.975 -228.265 44.255 ;
        RECT -226.305 44.575 -226.025 44.855 ;
        RECT -226.305 43.975 -226.025 44.255 ;
        RECT -227.425 41.215 -227.145 41.495 ;
        RECT -227.425 40.615 -227.145 40.895 ;
        RECT -229.665 37.855 -229.385 38.135 ;
        RECT -229.665 37.255 -229.385 37.535 ;
        RECT -234.145 34.495 -233.865 34.775 ;
        RECT -234.145 33.895 -233.865 34.175 ;
        RECT -243.105 31.135 -242.825 31.415 ;
        RECT -243.105 30.535 -242.825 30.815 ;
        RECT -224.065 44.575 -223.785 44.855 ;
        RECT -224.065 43.975 -223.785 44.255 ;
        RECT -221.825 44.575 -221.545 44.855 ;
        RECT -221.825 43.975 -221.545 44.255 ;
        RECT -222.945 41.215 -222.665 41.495 ;
        RECT -222.945 40.615 -222.665 40.895 ;
        RECT -219.585 44.575 -219.305 44.855 ;
        RECT -219.585 43.975 -219.305 44.255 ;
        RECT -217.345 44.575 -217.065 44.855 ;
        RECT -217.345 43.975 -217.065 44.255 ;
        RECT -218.465 41.215 -218.185 41.495 ;
        RECT -218.465 40.615 -218.185 40.895 ;
        RECT -220.705 37.855 -220.425 38.135 ;
        RECT -220.705 37.255 -220.425 37.535 ;
        RECT -215.105 44.575 -214.825 44.855 ;
        RECT -215.105 43.975 -214.825 44.255 ;
        RECT -212.865 44.575 -212.585 44.855 ;
        RECT -212.865 43.975 -212.585 44.255 ;
        RECT -213.985 41.215 -213.705 41.495 ;
        RECT -213.985 40.615 -213.705 40.895 ;
        RECT -210.625 44.575 -210.345 44.855 ;
        RECT -210.625 43.975 -210.345 44.255 ;
        RECT -208.385 44.575 -208.105 44.855 ;
        RECT -208.385 43.975 -208.105 44.255 ;
        RECT -209.505 41.215 -209.225 41.495 ;
        RECT -209.505 40.615 -209.225 40.895 ;
        RECT -211.745 37.855 -211.465 38.135 ;
        RECT -211.745 37.255 -211.465 37.535 ;
        RECT -216.225 34.495 -215.945 34.775 ;
        RECT -216.225 33.895 -215.945 34.175 ;
        RECT -206.145 44.575 -205.865 44.855 ;
        RECT -206.145 43.975 -205.865 44.255 ;
        RECT -203.905 44.575 -203.625 44.855 ;
        RECT -203.905 43.975 -203.625 44.255 ;
        RECT -205.025 41.215 -204.745 41.495 ;
        RECT -205.025 40.615 -204.745 40.895 ;
        RECT -201.665 44.575 -201.385 44.855 ;
        RECT -201.665 43.975 -201.385 44.255 ;
        RECT -199.425 44.575 -199.145 44.855 ;
        RECT -199.425 43.975 -199.145 44.255 ;
        RECT -200.545 41.215 -200.265 41.495 ;
        RECT -200.545 40.615 -200.265 40.895 ;
        RECT -202.785 37.855 -202.505 38.135 ;
        RECT -202.785 37.255 -202.505 37.535 ;
        RECT -197.185 44.575 -196.905 44.855 ;
        RECT -197.185 43.975 -196.905 44.255 ;
        RECT -194.945 44.575 -194.665 44.855 ;
        RECT -194.945 43.975 -194.665 44.255 ;
        RECT -196.065 41.215 -195.785 41.495 ;
        RECT -196.065 40.615 -195.785 40.895 ;
        RECT -192.705 44.575 -192.425 44.855 ;
        RECT -192.705 43.975 -192.425 44.255 ;
        RECT -190.465 44.575 -190.185 44.855 ;
        RECT -190.465 43.975 -190.185 44.255 ;
        RECT -191.585 41.215 -191.305 41.495 ;
        RECT -191.585 40.615 -191.305 40.895 ;
        RECT -193.825 37.855 -193.545 38.135 ;
        RECT -193.825 37.255 -193.545 37.535 ;
        RECT -198.305 34.495 -198.025 34.775 ;
        RECT -198.305 33.895 -198.025 34.175 ;
        RECT -207.265 31.135 -206.985 31.415 ;
        RECT -207.265 30.535 -206.985 30.815 ;
        RECT -225.185 27.775 -224.905 28.055 ;
        RECT -225.185 27.175 -224.905 27.455 ;
        RECT -261.025 24.415 -260.745 24.695 ;
        RECT -261.025 23.815 -260.745 24.095 ;
        RECT -332.705 21.055 -332.425 21.335 ;
        RECT -332.705 20.455 -332.425 20.735 ;
        RECT -187.105 44.575 -186.825 44.855 ;
        RECT -187.105 43.975 -186.825 44.255 ;
        RECT -184.865 44.575 -184.585 44.855 ;
        RECT -184.865 43.975 -184.585 44.255 ;
        RECT -185.985 41.215 -185.705 41.495 ;
        RECT -185.985 40.615 -185.705 40.895 ;
        RECT -182.625 44.575 -182.345 44.855 ;
        RECT -182.625 43.975 -182.345 44.255 ;
        RECT -180.385 44.575 -180.105 44.855 ;
        RECT -180.385 43.975 -180.105 44.255 ;
        RECT -181.505 41.215 -181.225 41.495 ;
        RECT -181.505 40.615 -181.225 40.895 ;
        RECT -183.745 37.855 -183.465 38.135 ;
        RECT -183.745 37.255 -183.465 37.535 ;
        RECT -178.145 44.575 -177.865 44.855 ;
        RECT -178.145 43.975 -177.865 44.255 ;
        RECT -175.905 44.575 -175.625 44.855 ;
        RECT -175.905 43.975 -175.625 44.255 ;
        RECT -177.025 41.215 -176.745 41.495 ;
        RECT -177.025 40.615 -176.745 40.895 ;
        RECT -173.665 44.575 -173.385 44.855 ;
        RECT -173.665 43.975 -173.385 44.255 ;
        RECT -171.425 44.575 -171.145 44.855 ;
        RECT -171.425 43.975 -171.145 44.255 ;
        RECT -172.545 41.215 -172.265 41.495 ;
        RECT -172.545 40.615 -172.265 40.895 ;
        RECT -174.785 37.855 -174.505 38.135 ;
        RECT -174.785 37.255 -174.505 37.535 ;
        RECT -179.265 34.495 -178.985 34.775 ;
        RECT -179.265 33.895 -178.985 34.175 ;
        RECT -169.185 44.575 -168.905 44.855 ;
        RECT -169.185 43.975 -168.905 44.255 ;
        RECT -166.945 44.575 -166.665 44.855 ;
        RECT -166.945 43.975 -166.665 44.255 ;
        RECT -168.065 41.215 -167.785 41.495 ;
        RECT -168.065 40.615 -167.785 40.895 ;
        RECT -164.705 44.575 -164.425 44.855 ;
        RECT -164.705 43.975 -164.425 44.255 ;
        RECT -162.465 44.575 -162.185 44.855 ;
        RECT -162.465 43.975 -162.185 44.255 ;
        RECT -163.585 41.215 -163.305 41.495 ;
        RECT -163.585 40.615 -163.305 40.895 ;
        RECT -165.825 37.855 -165.545 38.135 ;
        RECT -165.825 37.255 -165.545 37.535 ;
        RECT -160.225 44.575 -159.945 44.855 ;
        RECT -160.225 43.975 -159.945 44.255 ;
        RECT -157.985 44.575 -157.705 44.855 ;
        RECT -157.985 43.975 -157.705 44.255 ;
        RECT -159.105 41.215 -158.825 41.495 ;
        RECT -159.105 40.615 -158.825 40.895 ;
        RECT -155.745 44.575 -155.465 44.855 ;
        RECT -155.745 43.975 -155.465 44.255 ;
        RECT -153.505 44.575 -153.225 44.855 ;
        RECT -153.505 43.975 -153.225 44.255 ;
        RECT -154.625 41.215 -154.345 41.495 ;
        RECT -154.625 40.615 -154.345 40.895 ;
        RECT -156.865 37.855 -156.585 38.135 ;
        RECT -156.865 37.255 -156.585 37.535 ;
        RECT -161.345 34.495 -161.065 34.775 ;
        RECT -161.345 33.895 -161.065 34.175 ;
        RECT -170.305 31.135 -170.025 31.415 ;
        RECT -170.305 30.535 -170.025 30.815 ;
        RECT -151.265 44.575 -150.985 44.855 ;
        RECT -151.265 43.975 -150.985 44.255 ;
        RECT -149.025 44.575 -148.745 44.855 ;
        RECT -149.025 43.975 -148.745 44.255 ;
        RECT -150.145 41.215 -149.865 41.495 ;
        RECT -150.145 40.615 -149.865 40.895 ;
        RECT -146.785 44.575 -146.505 44.855 ;
        RECT -146.785 43.975 -146.505 44.255 ;
        RECT -144.545 44.575 -144.265 44.855 ;
        RECT -144.545 43.975 -144.265 44.255 ;
        RECT -145.665 41.215 -145.385 41.495 ;
        RECT -145.665 40.615 -145.385 40.895 ;
        RECT -147.905 37.855 -147.625 38.135 ;
        RECT -147.905 37.255 -147.625 37.535 ;
        RECT -142.305 44.575 -142.025 44.855 ;
        RECT -142.305 43.975 -142.025 44.255 ;
        RECT -140.065 44.575 -139.785 44.855 ;
        RECT -140.065 43.975 -139.785 44.255 ;
        RECT -141.185 41.215 -140.905 41.495 ;
        RECT -141.185 40.615 -140.905 40.895 ;
        RECT -137.825 44.575 -137.545 44.855 ;
        RECT -137.825 43.975 -137.545 44.255 ;
        RECT -135.585 44.575 -135.305 44.855 ;
        RECT -135.585 43.975 -135.305 44.255 ;
        RECT -136.705 41.215 -136.425 41.495 ;
        RECT -136.705 40.615 -136.425 40.895 ;
        RECT -138.945 37.855 -138.665 38.135 ;
        RECT -138.945 37.255 -138.665 37.535 ;
        RECT -143.425 34.495 -143.145 34.775 ;
        RECT -143.425 33.895 -143.145 34.175 ;
        RECT -133.345 44.575 -133.065 44.855 ;
        RECT -133.345 43.975 -133.065 44.255 ;
        RECT -131.105 44.575 -130.825 44.855 ;
        RECT -131.105 43.975 -130.825 44.255 ;
        RECT -132.225 41.215 -131.945 41.495 ;
        RECT -132.225 40.615 -131.945 40.895 ;
        RECT -128.865 44.575 -128.585 44.855 ;
        RECT -128.865 43.975 -128.585 44.255 ;
        RECT -126.625 44.575 -126.345 44.855 ;
        RECT -126.625 43.975 -126.345 44.255 ;
        RECT -127.745 41.215 -127.465 41.495 ;
        RECT -127.745 40.615 -127.465 40.895 ;
        RECT -129.985 37.855 -129.705 38.135 ;
        RECT -129.985 37.255 -129.705 37.535 ;
        RECT -124.385 44.575 -124.105 44.855 ;
        RECT -124.385 43.975 -124.105 44.255 ;
        RECT -122.145 44.575 -121.865 44.855 ;
        RECT -122.145 43.975 -121.865 44.255 ;
        RECT -123.265 41.215 -122.985 41.495 ;
        RECT -123.265 40.615 -122.985 40.895 ;
        RECT -119.905 44.575 -119.625 44.855 ;
        RECT -119.905 43.975 -119.625 44.255 ;
        RECT -117.665 44.575 -117.385 44.855 ;
        RECT -117.665 43.975 -117.385 44.255 ;
        RECT -118.785 41.215 -118.505 41.495 ;
        RECT -118.785 40.615 -118.505 40.895 ;
        RECT -121.025 37.855 -120.745 38.135 ;
        RECT -121.025 37.255 -120.745 37.535 ;
        RECT -125.505 34.495 -125.225 34.775 ;
        RECT -125.505 33.895 -125.225 34.175 ;
        RECT -134.465 31.135 -134.185 31.415 ;
        RECT -134.465 30.535 -134.185 30.815 ;
        RECT -152.385 27.775 -152.105 28.055 ;
        RECT -152.385 27.175 -152.105 27.455 ;
        RECT -115.425 44.575 -115.145 44.855 ;
        RECT -115.425 43.975 -115.145 44.255 ;
        RECT -113.185 44.575 -112.905 44.855 ;
        RECT -113.185 43.975 -112.905 44.255 ;
        RECT -114.305 41.215 -114.025 41.495 ;
        RECT -114.305 40.615 -114.025 40.895 ;
        RECT -110.945 44.575 -110.665 44.855 ;
        RECT -110.945 43.975 -110.665 44.255 ;
        RECT -108.705 44.575 -108.425 44.855 ;
        RECT -108.705 43.975 -108.425 44.255 ;
        RECT -109.825 41.215 -109.545 41.495 ;
        RECT -109.825 40.615 -109.545 40.895 ;
        RECT -112.065 37.855 -111.785 38.135 ;
        RECT -112.065 37.255 -111.785 37.535 ;
        RECT -106.465 44.575 -106.185 44.855 ;
        RECT -106.465 43.975 -106.185 44.255 ;
        RECT -104.225 44.575 -103.945 44.855 ;
        RECT -104.225 43.975 -103.945 44.255 ;
        RECT -105.345 41.215 -105.065 41.495 ;
        RECT -105.345 40.615 -105.065 40.895 ;
        RECT -101.985 44.575 -101.705 44.855 ;
        RECT -101.985 43.975 -101.705 44.255 ;
        RECT -99.745 44.575 -99.465 44.855 ;
        RECT -99.745 43.975 -99.465 44.255 ;
        RECT -100.865 41.215 -100.585 41.495 ;
        RECT -100.865 40.615 -100.585 40.895 ;
        RECT -103.105 37.855 -102.825 38.135 ;
        RECT -103.105 37.255 -102.825 37.535 ;
        RECT -107.585 34.495 -107.305 34.775 ;
        RECT -107.585 33.895 -107.305 34.175 ;
        RECT -97.505 44.575 -97.225 44.855 ;
        RECT -97.505 43.975 -97.225 44.255 ;
        RECT -95.265 44.575 -94.985 44.855 ;
        RECT -95.265 43.975 -94.985 44.255 ;
        RECT -96.385 41.215 -96.105 41.495 ;
        RECT -96.385 40.615 -96.105 40.895 ;
        RECT -93.025 44.575 -92.745 44.855 ;
        RECT -93.025 43.975 -92.745 44.255 ;
        RECT -90.785 44.575 -90.505 44.855 ;
        RECT -90.785 43.975 -90.505 44.255 ;
        RECT -91.905 41.215 -91.625 41.495 ;
        RECT -91.905 40.615 -91.625 40.895 ;
        RECT -94.145 37.855 -93.865 38.135 ;
        RECT -94.145 37.255 -93.865 37.535 ;
        RECT -88.545 44.575 -88.265 44.855 ;
        RECT -88.545 43.975 -88.265 44.255 ;
        RECT -86.305 44.575 -86.025 44.855 ;
        RECT -86.305 43.975 -86.025 44.255 ;
        RECT -87.425 41.215 -87.145 41.495 ;
        RECT -87.425 40.615 -87.145 40.895 ;
        RECT -84.065 44.575 -83.785 44.855 ;
        RECT -84.065 43.975 -83.785 44.255 ;
        RECT -81.825 44.575 -81.545 44.855 ;
        RECT -81.825 43.975 -81.545 44.255 ;
        RECT -82.945 41.215 -82.665 41.495 ;
        RECT -82.945 40.615 -82.665 40.895 ;
        RECT -85.185 37.855 -84.905 38.135 ;
        RECT -85.185 37.255 -84.905 37.535 ;
        RECT -89.665 34.495 -89.385 34.775 ;
        RECT -89.665 33.895 -89.385 34.175 ;
        RECT -98.625 31.135 -98.345 31.415 ;
        RECT -98.625 30.535 -98.345 30.815 ;
        RECT -79.585 44.575 -79.305 44.855 ;
        RECT -79.585 43.975 -79.305 44.255 ;
        RECT -77.345 44.575 -77.065 44.855 ;
        RECT -77.345 43.975 -77.065 44.255 ;
        RECT -78.465 41.215 -78.185 41.495 ;
        RECT -78.465 40.615 -78.185 40.895 ;
        RECT -75.105 44.575 -74.825 44.855 ;
        RECT -75.105 43.975 -74.825 44.255 ;
        RECT -72.865 44.575 -72.585 44.855 ;
        RECT -72.865 43.975 -72.585 44.255 ;
        RECT -73.985 41.215 -73.705 41.495 ;
        RECT -73.985 40.615 -73.705 40.895 ;
        RECT -76.225 37.855 -75.945 38.135 ;
        RECT -76.225 37.255 -75.945 37.535 ;
        RECT -70.625 44.575 -70.345 44.855 ;
        RECT -70.625 43.975 -70.345 44.255 ;
        RECT -68.385 44.575 -68.105 44.855 ;
        RECT -68.385 43.975 -68.105 44.255 ;
        RECT -69.505 41.215 -69.225 41.495 ;
        RECT -69.505 40.615 -69.225 40.895 ;
        RECT -66.145 44.575 -65.865 44.855 ;
        RECT -66.145 43.975 -65.865 44.255 ;
        RECT -63.905 44.575 -63.625 44.855 ;
        RECT -63.905 43.975 -63.625 44.255 ;
        RECT -65.025 41.215 -64.745 41.495 ;
        RECT -65.025 40.615 -64.745 40.895 ;
        RECT -67.265 37.855 -66.985 38.135 ;
        RECT -67.265 37.255 -66.985 37.535 ;
        RECT -71.745 34.495 -71.465 34.775 ;
        RECT -71.745 33.895 -71.465 34.175 ;
        RECT -61.665 44.575 -61.385 44.855 ;
        RECT -61.665 43.975 -61.385 44.255 ;
        RECT -59.425 44.575 -59.145 44.855 ;
        RECT -59.425 43.975 -59.145 44.255 ;
        RECT -60.545 41.215 -60.265 41.495 ;
        RECT -60.545 40.615 -60.265 40.895 ;
        RECT -57.185 44.575 -56.905 44.855 ;
        RECT -57.185 43.975 -56.905 44.255 ;
        RECT -54.945 44.575 -54.665 44.855 ;
        RECT -54.945 43.975 -54.665 44.255 ;
        RECT -56.065 41.215 -55.785 41.495 ;
        RECT -56.065 40.615 -55.785 40.895 ;
        RECT -58.305 37.855 -58.025 38.135 ;
        RECT -58.305 37.255 -58.025 37.535 ;
        RECT -52.705 44.575 -52.425 44.855 ;
        RECT -52.705 43.975 -52.425 44.255 ;
        RECT -50.465 44.575 -50.185 44.855 ;
        RECT -50.465 43.975 -50.185 44.255 ;
        RECT -51.585 41.215 -51.305 41.495 ;
        RECT -51.585 40.615 -51.305 40.895 ;
        RECT -48.225 44.575 -47.945 44.855 ;
        RECT -48.225 43.975 -47.945 44.255 ;
        RECT -45.985 44.575 -45.705 44.855 ;
        RECT -45.985 43.975 -45.705 44.255 ;
        RECT -47.105 41.215 -46.825 41.495 ;
        RECT -47.105 40.615 -46.825 40.895 ;
        RECT -49.345 37.855 -49.065 38.135 ;
        RECT -49.345 37.255 -49.065 37.535 ;
        RECT -53.825 34.495 -53.545 34.775 ;
        RECT -53.825 33.895 -53.545 34.175 ;
        RECT -62.785 31.135 -62.505 31.415 ;
        RECT -62.785 30.535 -62.505 30.815 ;
        RECT -80.705 27.775 -80.425 28.055 ;
        RECT -80.705 27.175 -80.425 27.455 ;
        RECT -116.545 24.415 -116.265 24.695 ;
        RECT -116.545 23.815 -116.265 24.095 ;
        RECT -43.745 44.575 -43.465 44.855 ;
        RECT -43.745 43.975 -43.465 44.255 ;
        RECT -41.505 44.575 -41.225 44.855 ;
        RECT -41.505 43.975 -41.225 44.255 ;
        RECT -42.625 41.215 -42.345 41.495 ;
        RECT -42.625 40.615 -42.345 40.895 ;
        RECT -39.265 44.575 -38.985 44.855 ;
        RECT -39.265 43.975 -38.985 44.255 ;
        RECT -37.025 44.575 -36.745 44.855 ;
        RECT -37.025 43.975 -36.745 44.255 ;
        RECT -38.145 41.215 -37.865 41.495 ;
        RECT -38.145 40.615 -37.865 40.895 ;
        RECT -40.385 37.855 -40.105 38.135 ;
        RECT -40.385 37.255 -40.105 37.535 ;
        RECT -34.785 44.575 -34.505 44.855 ;
        RECT -34.785 43.975 -34.505 44.255 ;
        RECT -32.545 44.575 -32.265 44.855 ;
        RECT -32.545 43.975 -32.265 44.255 ;
        RECT -33.665 41.215 -33.385 41.495 ;
        RECT -33.665 40.615 -33.385 40.895 ;
        RECT -30.305 44.575 -30.025 44.855 ;
        RECT -30.305 43.975 -30.025 44.255 ;
        RECT -28.065 44.575 -27.785 44.855 ;
        RECT -28.065 43.975 -27.785 44.255 ;
        RECT -29.185 41.215 -28.905 41.495 ;
        RECT -29.185 40.615 -28.905 40.895 ;
        RECT -31.425 37.855 -31.145 38.135 ;
        RECT -31.425 37.255 -31.145 37.535 ;
        RECT -35.905 34.495 -35.625 34.775 ;
        RECT -35.905 33.895 -35.625 34.175 ;
        RECT -25.825 44.575 -25.545 44.855 ;
        RECT -25.825 43.975 -25.545 44.255 ;
        RECT -23.585 44.575 -23.305 44.855 ;
        RECT -23.585 43.975 -23.305 44.255 ;
        RECT -24.705 41.215 -24.425 41.495 ;
        RECT -24.705 40.615 -24.425 40.895 ;
        RECT -21.345 44.575 -21.065 44.855 ;
        RECT -21.345 43.975 -21.065 44.255 ;
        RECT -19.105 44.575 -18.825 44.855 ;
        RECT -19.105 43.975 -18.825 44.255 ;
        RECT -20.225 41.215 -19.945 41.495 ;
        RECT -20.225 40.615 -19.945 40.895 ;
        RECT -22.465 37.855 -22.185 38.135 ;
        RECT -22.465 37.255 -22.185 37.535 ;
        RECT -16.865 44.575 -16.585 44.855 ;
        RECT -16.865 43.975 -16.585 44.255 ;
        RECT -14.625 44.575 -14.345 44.855 ;
        RECT -14.625 43.975 -14.345 44.255 ;
        RECT -15.745 41.215 -15.465 41.495 ;
        RECT -15.745 40.615 -15.465 40.895 ;
        RECT -12.385 44.575 -12.105 44.855 ;
        RECT -12.385 43.975 -12.105 44.255 ;
        RECT -10.145 44.575 -9.865 44.855 ;
        RECT -10.145 43.975 -9.865 44.255 ;
        RECT -11.265 41.215 -10.985 41.495 ;
        RECT -11.265 40.615 -10.985 40.895 ;
        RECT -13.505 37.855 -13.225 38.135 ;
        RECT -13.505 37.255 -13.225 37.535 ;
        RECT -17.985 34.495 -17.705 34.775 ;
        RECT -17.985 33.895 -17.705 34.175 ;
        RECT -26.945 31.135 -26.665 31.415 ;
        RECT -26.945 30.535 -26.665 30.815 ;
        RECT -7.905 44.575 -7.625 44.855 ;
        RECT -7.905 43.975 -7.625 44.255 ;
        RECT -5.665 44.575 -5.385 44.855 ;
        RECT -5.665 43.975 -5.385 44.255 ;
        RECT -6.785 41.215 -6.505 41.495 ;
        RECT -6.785 40.615 -6.505 40.895 ;
        RECT -3.425 44.575 -3.145 44.855 ;
        RECT -3.425 43.975 -3.145 44.255 ;
        RECT -1.185 44.575 -0.905 44.855 ;
        RECT -1.185 43.975 -0.905 44.255 ;
        RECT -2.305 41.215 -2.025 41.495 ;
        RECT -2.305 40.615 -2.025 40.895 ;
        RECT -4.545 37.855 -4.265 38.135 ;
        RECT -4.545 37.255 -4.265 37.535 ;
        RECT 1.055 44.575 1.335 44.855 ;
        RECT 1.055 43.975 1.335 44.255 ;
        RECT 3.295 44.575 3.575 44.855 ;
        RECT 3.295 43.975 3.575 44.255 ;
        RECT 2.175 41.215 2.455 41.495 ;
        RECT 2.175 40.615 2.455 40.895 ;
        RECT 5.535 44.575 5.815 44.855 ;
        RECT 5.535 43.975 5.815 44.255 ;
        RECT 7.775 44.575 8.055 44.855 ;
        RECT 7.775 43.975 8.055 44.255 ;
        RECT 6.655 41.215 6.935 41.495 ;
        RECT 6.655 40.615 6.935 40.895 ;
        RECT 4.415 37.855 4.695 38.135 ;
        RECT 4.415 37.255 4.695 37.535 ;
        RECT -0.065 34.495 0.215 34.775 ;
        RECT -0.065 33.895 0.215 34.175 ;
        RECT 10.015 44.575 10.295 44.855 ;
        RECT 10.015 43.975 10.295 44.255 ;
        RECT 12.255 44.575 12.535 44.855 ;
        RECT 12.255 43.975 12.535 44.255 ;
        RECT 11.135 41.215 11.415 41.495 ;
        RECT 11.135 40.615 11.415 40.895 ;
        RECT 14.495 44.575 14.775 44.855 ;
        RECT 14.495 43.975 14.775 44.255 ;
        RECT 16.735 44.575 17.015 44.855 ;
        RECT 16.735 43.975 17.015 44.255 ;
        RECT 15.615 41.215 15.895 41.495 ;
        RECT 15.615 40.615 15.895 40.895 ;
        RECT 13.375 37.855 13.655 38.135 ;
        RECT 13.375 37.255 13.655 37.535 ;
        RECT 18.975 44.575 19.255 44.855 ;
        RECT 18.975 43.975 19.255 44.255 ;
        RECT 21.215 44.575 21.495 44.855 ;
        RECT 21.215 43.975 21.495 44.255 ;
        RECT 20.095 41.215 20.375 41.495 ;
        RECT 20.095 40.615 20.375 40.895 ;
        RECT 23.455 44.575 23.735 44.855 ;
        RECT 23.455 43.975 23.735 44.255 ;
        RECT 25.695 44.575 25.975 44.855 ;
        RECT 25.695 43.975 25.975 44.255 ;
        RECT 24.575 41.215 24.855 41.495 ;
        RECT 24.575 40.615 24.855 40.895 ;
        RECT 22.335 37.855 22.615 38.135 ;
        RECT 22.335 37.255 22.615 37.535 ;
        RECT 17.855 34.495 18.135 34.775 ;
        RECT 17.855 33.895 18.135 34.175 ;
        RECT 8.895 31.135 9.175 31.415 ;
        RECT 8.895 30.535 9.175 30.815 ;
        RECT -9.025 27.775 -8.745 28.055 ;
        RECT -9.025 27.175 -8.745 27.455 ;
        RECT 27.935 44.575 28.215 44.855 ;
        RECT 27.935 43.975 28.215 44.255 ;
        RECT 30.175 44.575 30.455 44.855 ;
        RECT 30.175 43.975 30.455 44.255 ;
        RECT 29.055 41.215 29.335 41.495 ;
        RECT 29.055 40.615 29.335 40.895 ;
        RECT 32.415 44.575 32.695 44.855 ;
        RECT 32.415 43.975 32.695 44.255 ;
        RECT 34.655 44.575 34.935 44.855 ;
        RECT 34.655 43.975 34.935 44.255 ;
        RECT 33.535 41.215 33.815 41.495 ;
        RECT 33.535 40.615 33.815 40.895 ;
        RECT 31.295 37.855 31.575 38.135 ;
        RECT 31.295 37.255 31.575 37.535 ;
        RECT 36.895 44.575 37.175 44.855 ;
        RECT 36.895 43.975 37.175 44.255 ;
        RECT 39.135 44.575 39.415 44.855 ;
        RECT 39.135 43.975 39.415 44.255 ;
        RECT 38.015 41.215 38.295 41.495 ;
        RECT 38.015 40.615 38.295 40.895 ;
        RECT 41.375 44.575 41.655 44.855 ;
        RECT 41.375 43.975 41.655 44.255 ;
        RECT 43.615 44.575 43.895 44.855 ;
        RECT 43.615 43.975 43.895 44.255 ;
        RECT 42.495 41.215 42.775 41.495 ;
        RECT 42.495 40.615 42.775 40.895 ;
        RECT 40.255 37.855 40.535 38.135 ;
        RECT 40.255 37.255 40.535 37.535 ;
        RECT 35.775 34.495 36.055 34.775 ;
        RECT 35.775 33.895 36.055 34.175 ;
        RECT 45.855 44.575 46.135 44.855 ;
        RECT 45.855 43.975 46.135 44.255 ;
        RECT 48.095 44.575 48.375 44.855 ;
        RECT 48.095 43.975 48.375 44.255 ;
        RECT 46.975 41.215 47.255 41.495 ;
        RECT 46.975 40.615 47.255 40.895 ;
        RECT 50.335 44.575 50.615 44.855 ;
        RECT 50.335 43.975 50.615 44.255 ;
        RECT 52.575 44.575 52.855 44.855 ;
        RECT 52.575 43.975 52.855 44.255 ;
        RECT 51.455 41.215 51.735 41.495 ;
        RECT 51.455 40.615 51.735 40.895 ;
        RECT 49.215 37.855 49.495 38.135 ;
        RECT 49.215 37.255 49.495 37.535 ;
        RECT 54.815 44.575 55.095 44.855 ;
        RECT 54.815 43.975 55.095 44.255 ;
        RECT 57.055 44.575 57.335 44.855 ;
        RECT 57.055 43.975 57.335 44.255 ;
        RECT 55.935 41.215 56.215 41.495 ;
        RECT 55.935 40.615 56.215 40.895 ;
        RECT 59.295 44.575 59.575 44.855 ;
        RECT 59.295 43.975 59.575 44.255 ;
        RECT 61.535 44.575 61.815 44.855 ;
        RECT 61.535 43.975 61.815 44.255 ;
        RECT 60.415 41.215 60.695 41.495 ;
        RECT 60.415 40.615 60.695 40.895 ;
        RECT 58.175 37.855 58.455 38.135 ;
        RECT 58.175 37.255 58.455 37.535 ;
        RECT 53.695 34.495 53.975 34.775 ;
        RECT 53.695 33.895 53.975 34.175 ;
        RECT 44.735 31.135 45.015 31.415 ;
        RECT 44.735 30.535 45.015 30.815 ;
        RECT 63.775 44.575 64.055 44.855 ;
        RECT 63.775 43.975 64.055 44.255 ;
        RECT 66.015 44.575 66.295 44.855 ;
        RECT 66.015 43.975 66.295 44.255 ;
        RECT 64.895 41.215 65.175 41.495 ;
        RECT 64.895 40.615 65.175 40.895 ;
        RECT 68.255 44.575 68.535 44.855 ;
        RECT 68.255 43.975 68.535 44.255 ;
        RECT 70.495 44.575 70.775 44.855 ;
        RECT 70.495 43.975 70.775 44.255 ;
        RECT 69.375 41.215 69.655 41.495 ;
        RECT 69.375 40.615 69.655 40.895 ;
        RECT 67.135 37.855 67.415 38.135 ;
        RECT 67.135 37.255 67.415 37.535 ;
        RECT 72.735 44.575 73.015 44.855 ;
        RECT 72.735 43.975 73.015 44.255 ;
        RECT 74.975 44.575 75.255 44.855 ;
        RECT 74.975 43.975 75.255 44.255 ;
        RECT 73.855 41.215 74.135 41.495 ;
        RECT 73.855 40.615 74.135 40.895 ;
        RECT 77.215 44.575 77.495 44.855 ;
        RECT 77.215 43.975 77.495 44.255 ;
        RECT 79.455 44.575 79.735 44.855 ;
        RECT 79.455 43.975 79.735 44.255 ;
        RECT 78.335 41.215 78.615 41.495 ;
        RECT 78.335 40.615 78.615 40.895 ;
        RECT 76.095 37.855 76.375 38.135 ;
        RECT 76.095 37.255 76.375 37.535 ;
        RECT 71.615 34.495 71.895 34.775 ;
        RECT 71.615 33.895 71.895 34.175 ;
        RECT 81.695 44.575 81.975 44.855 ;
        RECT 81.695 43.975 81.975 44.255 ;
        RECT 83.935 44.575 84.215 44.855 ;
        RECT 83.935 43.975 84.215 44.255 ;
        RECT 82.815 41.215 83.095 41.495 ;
        RECT 82.815 40.615 83.095 40.895 ;
        RECT 86.175 44.575 86.455 44.855 ;
        RECT 86.175 43.975 86.455 44.255 ;
        RECT 88.415 44.575 88.695 44.855 ;
        RECT 88.415 43.975 88.695 44.255 ;
        RECT 87.295 41.215 87.575 41.495 ;
        RECT 87.295 40.615 87.575 40.895 ;
        RECT 85.055 37.855 85.335 38.135 ;
        RECT 85.055 37.255 85.335 37.535 ;
        RECT 90.655 44.575 90.935 44.855 ;
        RECT 90.655 43.975 90.935 44.255 ;
        RECT 92.895 44.575 93.175 44.855 ;
        RECT 92.895 43.975 93.175 44.255 ;
        RECT 91.775 41.215 92.055 41.495 ;
        RECT 91.775 40.615 92.055 40.895 ;
        RECT 95.135 44.575 95.415 44.855 ;
        RECT 95.135 43.975 95.415 44.255 ;
        RECT 97.375 44.575 97.655 44.855 ;
        RECT 97.375 43.975 97.655 44.255 ;
        RECT 96.255 41.215 96.535 41.495 ;
        RECT 96.255 40.615 96.535 40.895 ;
        RECT 94.015 37.855 94.295 38.135 ;
        RECT 94.015 37.255 94.295 37.535 ;
        RECT 89.535 34.495 89.815 34.775 ;
        RECT 89.535 33.895 89.815 34.175 ;
        RECT 80.575 31.135 80.855 31.415 ;
        RECT 80.575 30.535 80.855 30.815 ;
        RECT 62.655 27.775 62.935 28.055 ;
        RECT 62.655 27.175 62.935 27.455 ;
        RECT 26.815 24.415 27.095 24.695 ;
        RECT 26.815 23.815 27.095 24.095 ;
        RECT -44.865 21.055 -44.585 21.335 ;
        RECT -44.865 20.455 -44.585 20.735 ;
        RECT -188.225 17.695 -187.945 17.975 ;
        RECT -188.225 17.095 -187.945 17.375 ;
        RECT -189.345 14.335 -189.065 14.615 ;
        RECT -189.345 13.735 -189.065 14.015 ;
        RECT 287.250 55.260 287.530 55.540 ;
        RECT 287.810 55.260 288.090 55.540 ;
        RECT 288.370 55.260 288.650 55.540 ;
        RECT 287.250 54.700 287.530 54.980 ;
        RECT 287.810 54.700 288.090 54.980 ;
        RECT 288.370 54.700 288.650 54.980 ;
        RECT 299.420 54.980 299.700 55.260 ;
        RECT 287.250 45.180 287.530 45.460 ;
        RECT 287.810 45.180 288.090 45.460 ;
        RECT 288.370 45.180 288.650 45.460 ;
        RECT 287.250 44.620 287.530 44.900 ;
        RECT 287.810 44.620 288.090 44.900 ;
        RECT 288.370 44.620 288.650 44.900 ;
        RECT 298.860 44.900 299.140 45.180 ;
        RECT 287.250 35.100 287.530 35.380 ;
        RECT 287.810 35.100 288.090 35.380 ;
        RECT 288.370 35.100 288.650 35.380 ;
        RECT 287.250 34.540 287.530 34.820 ;
        RECT 287.810 34.540 288.090 34.820 ;
        RECT 288.370 34.540 288.650 34.820 ;
        RECT 298.860 34.820 299.140 35.100 ;
        RECT 316.220 52.180 316.500 52.460 ;
        RECT 322.380 52.180 322.660 52.460 ;
        RECT 352.060 47.700 352.340 47.980 ;
        RECT 359.900 47.700 360.180 47.980 ;
        RECT 369.980 47.700 370.260 47.980 ;
        RECT 375.020 47.700 375.300 47.980 ;
        RECT 387.900 47.700 388.180 47.980 ;
        RECT 394.060 47.700 394.340 47.980 ;
        RECT 405.820 47.700 406.100 47.980 ;
        RECT 417.020 47.700 417.300 47.980 ;
        RECT 423.740 47.700 424.020 47.980 ;
        RECT 432.140 47.700 432.420 47.980 ;
        RECT 309.500 42.100 309.780 42.380 ;
        RECT 302.780 38.740 303.060 39.020 ;
        RECT 308.380 38.740 308.660 39.020 ;
        RECT 287.250 25.020 287.530 25.300 ;
        RECT 287.810 25.020 288.090 25.300 ;
        RECT 288.370 25.020 288.650 25.300 ;
        RECT 287.250 24.460 287.530 24.740 ;
        RECT 287.810 24.460 288.090 24.740 ;
        RECT 288.370 24.460 288.650 24.740 ;
        RECT 287.250 14.940 287.530 15.220 ;
        RECT 287.810 14.940 288.090 15.220 ;
        RECT 288.370 14.940 288.650 15.220 ;
        RECT 287.250 14.380 287.530 14.660 ;
        RECT 287.810 14.380 288.090 14.660 ;
        RECT 288.370 14.380 288.650 14.660 ;
        RECT 298.860 15.780 299.140 16.060 ;
        RECT 297.740 11.300 298.020 11.580 ;
        RECT 236.000 5.040 237.320 7.400 ;
        RECT 236.000 2.040 237.320 4.400 ;
        RECT 287.250 4.860 287.530 5.140 ;
        RECT 287.810 4.860 288.090 5.140 ;
        RECT 288.370 4.860 288.650 5.140 ;
        RECT 287.250 4.300 287.530 4.580 ;
        RECT 287.810 4.300 288.090 4.580 ;
        RECT 288.370 4.300 288.650 4.580 ;
        RECT 299.420 7.380 299.700 7.660 ;
        RECT 298.300 4.580 298.580 4.860 ;
        RECT 230.020 -5.725 232.380 -4.405 ;
        RECT 233.020 -5.725 235.380 -4.405 ;
        RECT 299.420 -4.380 299.700 -4.100 ;
        RECT 287.250 -5.220 287.530 -4.940 ;
        RECT 287.810 -5.220 288.090 -4.940 ;
        RECT 288.370 -5.220 288.650 -4.940 ;
        RECT 287.250 -5.780 287.530 -5.500 ;
        RECT 287.810 -5.780 288.090 -5.500 ;
        RECT 288.370 -5.780 288.650 -5.500 ;
        RECT 298.860 -5.500 299.140 -5.220 ;
        RECT -189.345 -14.015 -189.065 -13.735 ;
        RECT -189.345 -14.615 -189.065 -14.335 ;
        RECT -332.705 -20.735 -332.425 -20.455 ;
        RECT -332.705 -21.335 -332.425 -21.055 ;
        RECT -404.385 -24.095 -404.105 -23.815 ;
        RECT -404.385 -24.695 -404.105 -24.415 ;
        RECT -440.225 -27.455 -439.945 -27.175 ;
        RECT -440.225 -28.055 -439.945 -27.775 ;
        RECT -458.145 -30.815 -457.865 -30.535 ;
        RECT -458.145 -31.415 -457.865 -31.135 ;
        RECT -467.105 -34.175 -466.825 -33.895 ;
        RECT -467.105 -34.775 -466.825 -34.495 ;
        RECT -471.585 -37.535 -471.305 -37.255 ;
        RECT -471.585 -38.135 -471.305 -37.855 ;
        RECT -473.825 -40.895 -473.545 -40.615 ;
        RECT -473.825 -41.495 -473.545 -41.215 ;
        RECT -474.945 -44.255 -474.665 -43.975 ;
        RECT -474.945 -44.855 -474.665 -44.575 ;
        RECT -472.705 -44.255 -472.425 -43.975 ;
        RECT -472.705 -44.855 -472.425 -44.575 ;
        RECT -469.345 -40.895 -469.065 -40.615 ;
        RECT -469.345 -41.495 -469.065 -41.215 ;
        RECT -470.465 -44.255 -470.185 -43.975 ;
        RECT -470.465 -44.855 -470.185 -44.575 ;
        RECT -468.225 -44.255 -467.945 -43.975 ;
        RECT -468.225 -44.855 -467.945 -44.575 ;
        RECT -462.625 -37.535 -462.345 -37.255 ;
        RECT -462.625 -38.135 -462.345 -37.855 ;
        RECT -464.865 -40.895 -464.585 -40.615 ;
        RECT -464.865 -41.495 -464.585 -41.215 ;
        RECT -465.985 -44.255 -465.705 -43.975 ;
        RECT -465.985 -44.855 -465.705 -44.575 ;
        RECT -463.745 -44.255 -463.465 -43.975 ;
        RECT -463.745 -44.855 -463.465 -44.575 ;
        RECT -460.385 -40.895 -460.105 -40.615 ;
        RECT -460.385 -41.495 -460.105 -41.215 ;
        RECT -461.505 -44.255 -461.225 -43.975 ;
        RECT -461.505 -44.855 -461.225 -44.575 ;
        RECT -459.265 -44.255 -458.985 -43.975 ;
        RECT -459.265 -44.855 -458.985 -44.575 ;
        RECT -449.185 -34.175 -448.905 -33.895 ;
        RECT -449.185 -34.775 -448.905 -34.495 ;
        RECT -453.665 -37.535 -453.385 -37.255 ;
        RECT -453.665 -38.135 -453.385 -37.855 ;
        RECT -455.905 -40.895 -455.625 -40.615 ;
        RECT -455.905 -41.495 -455.625 -41.215 ;
        RECT -457.025 -44.255 -456.745 -43.975 ;
        RECT -457.025 -44.855 -456.745 -44.575 ;
        RECT -454.785 -44.255 -454.505 -43.975 ;
        RECT -454.785 -44.855 -454.505 -44.575 ;
        RECT -451.425 -40.895 -451.145 -40.615 ;
        RECT -451.425 -41.495 -451.145 -41.215 ;
        RECT -452.545 -44.255 -452.265 -43.975 ;
        RECT -452.545 -44.855 -452.265 -44.575 ;
        RECT -450.305 -44.255 -450.025 -43.975 ;
        RECT -450.305 -44.855 -450.025 -44.575 ;
        RECT -444.705 -37.535 -444.425 -37.255 ;
        RECT -444.705 -38.135 -444.425 -37.855 ;
        RECT -446.945 -40.895 -446.665 -40.615 ;
        RECT -446.945 -41.495 -446.665 -41.215 ;
        RECT -448.065 -44.255 -447.785 -43.975 ;
        RECT -448.065 -44.855 -447.785 -44.575 ;
        RECT -445.825 -44.255 -445.545 -43.975 ;
        RECT -445.825 -44.855 -445.545 -44.575 ;
        RECT -442.465 -40.895 -442.185 -40.615 ;
        RECT -442.465 -41.495 -442.185 -41.215 ;
        RECT -443.585 -44.255 -443.305 -43.975 ;
        RECT -443.585 -44.855 -443.305 -44.575 ;
        RECT -441.345 -44.255 -441.065 -43.975 ;
        RECT -441.345 -44.855 -441.065 -44.575 ;
        RECT -422.305 -30.815 -422.025 -30.535 ;
        RECT -422.305 -31.415 -422.025 -31.135 ;
        RECT -431.265 -34.175 -430.985 -33.895 ;
        RECT -431.265 -34.775 -430.985 -34.495 ;
        RECT -435.745 -37.535 -435.465 -37.255 ;
        RECT -435.745 -38.135 -435.465 -37.855 ;
        RECT -437.985 -40.895 -437.705 -40.615 ;
        RECT -437.985 -41.495 -437.705 -41.215 ;
        RECT -439.105 -44.255 -438.825 -43.975 ;
        RECT -439.105 -44.855 -438.825 -44.575 ;
        RECT -436.865 -44.255 -436.585 -43.975 ;
        RECT -436.865 -44.855 -436.585 -44.575 ;
        RECT -433.505 -40.895 -433.225 -40.615 ;
        RECT -433.505 -41.495 -433.225 -41.215 ;
        RECT -434.625 -44.255 -434.345 -43.975 ;
        RECT -434.625 -44.855 -434.345 -44.575 ;
        RECT -432.385 -44.255 -432.105 -43.975 ;
        RECT -432.385 -44.855 -432.105 -44.575 ;
        RECT -426.785 -37.535 -426.505 -37.255 ;
        RECT -426.785 -38.135 -426.505 -37.855 ;
        RECT -429.025 -40.895 -428.745 -40.615 ;
        RECT -429.025 -41.495 -428.745 -41.215 ;
        RECT -430.145 -44.255 -429.865 -43.975 ;
        RECT -430.145 -44.855 -429.865 -44.575 ;
        RECT -427.905 -44.255 -427.625 -43.975 ;
        RECT -427.905 -44.855 -427.625 -44.575 ;
        RECT -424.545 -40.895 -424.265 -40.615 ;
        RECT -424.545 -41.495 -424.265 -41.215 ;
        RECT -425.665 -44.255 -425.385 -43.975 ;
        RECT -425.665 -44.855 -425.385 -44.575 ;
        RECT -423.425 -44.255 -423.145 -43.975 ;
        RECT -423.425 -44.855 -423.145 -44.575 ;
        RECT -413.345 -34.175 -413.065 -33.895 ;
        RECT -413.345 -34.775 -413.065 -34.495 ;
        RECT -417.825 -37.535 -417.545 -37.255 ;
        RECT -417.825 -38.135 -417.545 -37.855 ;
        RECT -420.065 -40.895 -419.785 -40.615 ;
        RECT -420.065 -41.495 -419.785 -41.215 ;
        RECT -421.185 -44.255 -420.905 -43.975 ;
        RECT -421.185 -44.855 -420.905 -44.575 ;
        RECT -418.945 -44.255 -418.665 -43.975 ;
        RECT -418.945 -44.855 -418.665 -44.575 ;
        RECT -415.585 -40.895 -415.305 -40.615 ;
        RECT -415.585 -41.495 -415.305 -41.215 ;
        RECT -416.705 -44.255 -416.425 -43.975 ;
        RECT -416.705 -44.855 -416.425 -44.575 ;
        RECT -414.465 -44.255 -414.185 -43.975 ;
        RECT -414.465 -44.855 -414.185 -44.575 ;
        RECT -408.865 -37.535 -408.585 -37.255 ;
        RECT -408.865 -38.135 -408.585 -37.855 ;
        RECT -411.105 -40.895 -410.825 -40.615 ;
        RECT -411.105 -41.495 -410.825 -41.215 ;
        RECT -412.225 -44.255 -411.945 -43.975 ;
        RECT -412.225 -44.855 -411.945 -44.575 ;
        RECT -409.985 -44.255 -409.705 -43.975 ;
        RECT -409.985 -44.855 -409.705 -44.575 ;
        RECT -406.625 -40.895 -406.345 -40.615 ;
        RECT -406.625 -41.495 -406.345 -41.215 ;
        RECT -407.745 -44.255 -407.465 -43.975 ;
        RECT -407.745 -44.855 -407.465 -44.575 ;
        RECT -405.505 -44.255 -405.225 -43.975 ;
        RECT -405.505 -44.855 -405.225 -44.575 ;
        RECT -368.545 -27.455 -368.265 -27.175 ;
        RECT -368.545 -28.055 -368.265 -27.775 ;
        RECT -386.465 -30.815 -386.185 -30.535 ;
        RECT -386.465 -31.415 -386.185 -31.135 ;
        RECT -395.425 -34.175 -395.145 -33.895 ;
        RECT -395.425 -34.775 -395.145 -34.495 ;
        RECT -399.905 -37.535 -399.625 -37.255 ;
        RECT -399.905 -38.135 -399.625 -37.855 ;
        RECT -402.145 -40.895 -401.865 -40.615 ;
        RECT -402.145 -41.495 -401.865 -41.215 ;
        RECT -403.265 -44.255 -402.985 -43.975 ;
        RECT -403.265 -44.855 -402.985 -44.575 ;
        RECT -401.025 -44.255 -400.745 -43.975 ;
        RECT -401.025 -44.855 -400.745 -44.575 ;
        RECT -397.665 -40.895 -397.385 -40.615 ;
        RECT -397.665 -41.495 -397.385 -41.215 ;
        RECT -398.785 -44.255 -398.505 -43.975 ;
        RECT -398.785 -44.855 -398.505 -44.575 ;
        RECT -396.545 -44.255 -396.265 -43.975 ;
        RECT -396.545 -44.855 -396.265 -44.575 ;
        RECT -390.945 -37.535 -390.665 -37.255 ;
        RECT -390.945 -38.135 -390.665 -37.855 ;
        RECT -393.185 -40.895 -392.905 -40.615 ;
        RECT -393.185 -41.495 -392.905 -41.215 ;
        RECT -394.305 -44.255 -394.025 -43.975 ;
        RECT -394.305 -44.855 -394.025 -44.575 ;
        RECT -392.065 -44.255 -391.785 -43.975 ;
        RECT -392.065 -44.855 -391.785 -44.575 ;
        RECT -388.705 -40.895 -388.425 -40.615 ;
        RECT -388.705 -41.495 -388.425 -41.215 ;
        RECT -389.825 -44.255 -389.545 -43.975 ;
        RECT -389.825 -44.855 -389.545 -44.575 ;
        RECT -387.585 -44.255 -387.305 -43.975 ;
        RECT -387.585 -44.855 -387.305 -44.575 ;
        RECT -377.505 -34.175 -377.225 -33.895 ;
        RECT -377.505 -34.775 -377.225 -34.495 ;
        RECT -381.985 -37.535 -381.705 -37.255 ;
        RECT -381.985 -38.135 -381.705 -37.855 ;
        RECT -384.225 -40.895 -383.945 -40.615 ;
        RECT -384.225 -41.495 -383.945 -41.215 ;
        RECT -385.345 -44.255 -385.065 -43.975 ;
        RECT -385.345 -44.855 -385.065 -44.575 ;
        RECT -383.105 -44.255 -382.825 -43.975 ;
        RECT -383.105 -44.855 -382.825 -44.575 ;
        RECT -379.745 -40.895 -379.465 -40.615 ;
        RECT -379.745 -41.495 -379.465 -41.215 ;
        RECT -380.865 -44.255 -380.585 -43.975 ;
        RECT -380.865 -44.855 -380.585 -44.575 ;
        RECT -378.625 -44.255 -378.345 -43.975 ;
        RECT -378.625 -44.855 -378.345 -44.575 ;
        RECT -373.025 -37.535 -372.745 -37.255 ;
        RECT -373.025 -38.135 -372.745 -37.855 ;
        RECT -375.265 -40.895 -374.985 -40.615 ;
        RECT -375.265 -41.495 -374.985 -41.215 ;
        RECT -376.385 -44.255 -376.105 -43.975 ;
        RECT -376.385 -44.855 -376.105 -44.575 ;
        RECT -374.145 -44.255 -373.865 -43.975 ;
        RECT -374.145 -44.855 -373.865 -44.575 ;
        RECT -370.785 -40.895 -370.505 -40.615 ;
        RECT -370.785 -41.495 -370.505 -41.215 ;
        RECT -371.905 -44.255 -371.625 -43.975 ;
        RECT -371.905 -44.855 -371.625 -44.575 ;
        RECT -369.665 -44.255 -369.385 -43.975 ;
        RECT -369.665 -44.855 -369.385 -44.575 ;
        RECT -350.625 -30.815 -350.345 -30.535 ;
        RECT -350.625 -31.415 -350.345 -31.135 ;
        RECT -359.585 -34.175 -359.305 -33.895 ;
        RECT -359.585 -34.775 -359.305 -34.495 ;
        RECT -364.065 -37.535 -363.785 -37.255 ;
        RECT -364.065 -38.135 -363.785 -37.855 ;
        RECT -366.305 -40.895 -366.025 -40.615 ;
        RECT -366.305 -41.495 -366.025 -41.215 ;
        RECT -367.425 -44.255 -367.145 -43.975 ;
        RECT -367.425 -44.855 -367.145 -44.575 ;
        RECT -365.185 -44.255 -364.905 -43.975 ;
        RECT -365.185 -44.855 -364.905 -44.575 ;
        RECT -361.825 -40.895 -361.545 -40.615 ;
        RECT -361.825 -41.495 -361.545 -41.215 ;
        RECT -362.945 -44.255 -362.665 -43.975 ;
        RECT -362.945 -44.855 -362.665 -44.575 ;
        RECT -360.705 -44.255 -360.425 -43.975 ;
        RECT -360.705 -44.855 -360.425 -44.575 ;
        RECT -355.105 -37.535 -354.825 -37.255 ;
        RECT -355.105 -38.135 -354.825 -37.855 ;
        RECT -357.345 -40.895 -357.065 -40.615 ;
        RECT -357.345 -41.495 -357.065 -41.215 ;
        RECT -358.465 -44.255 -358.185 -43.975 ;
        RECT -358.465 -44.855 -358.185 -44.575 ;
        RECT -356.225 -44.255 -355.945 -43.975 ;
        RECT -356.225 -44.855 -355.945 -44.575 ;
        RECT -352.865 -40.895 -352.585 -40.615 ;
        RECT -352.865 -41.495 -352.585 -41.215 ;
        RECT -353.985 -44.255 -353.705 -43.975 ;
        RECT -353.985 -44.855 -353.705 -44.575 ;
        RECT -351.745 -44.255 -351.465 -43.975 ;
        RECT -351.745 -44.855 -351.465 -44.575 ;
        RECT -341.665 -34.175 -341.385 -33.895 ;
        RECT -341.665 -34.775 -341.385 -34.495 ;
        RECT -346.145 -37.535 -345.865 -37.255 ;
        RECT -346.145 -38.135 -345.865 -37.855 ;
        RECT -348.385 -40.895 -348.105 -40.615 ;
        RECT -348.385 -41.495 -348.105 -41.215 ;
        RECT -349.505 -44.255 -349.225 -43.975 ;
        RECT -349.505 -44.855 -349.225 -44.575 ;
        RECT -347.265 -44.255 -346.985 -43.975 ;
        RECT -347.265 -44.855 -346.985 -44.575 ;
        RECT -343.905 -40.895 -343.625 -40.615 ;
        RECT -343.905 -41.495 -343.625 -41.215 ;
        RECT -345.025 -44.255 -344.745 -43.975 ;
        RECT -345.025 -44.855 -344.745 -44.575 ;
        RECT -342.785 -44.255 -342.505 -43.975 ;
        RECT -342.785 -44.855 -342.505 -44.575 ;
        RECT -337.185 -37.535 -336.905 -37.255 ;
        RECT -337.185 -38.135 -336.905 -37.855 ;
        RECT -339.425 -40.895 -339.145 -40.615 ;
        RECT -339.425 -41.495 -339.145 -41.215 ;
        RECT -340.545 -44.255 -340.265 -43.975 ;
        RECT -340.545 -44.855 -340.265 -44.575 ;
        RECT -338.305 -44.255 -338.025 -43.975 ;
        RECT -338.305 -44.855 -338.025 -44.575 ;
        RECT -334.945 -40.895 -334.665 -40.615 ;
        RECT -334.945 -41.495 -334.665 -41.215 ;
        RECT -336.065 -44.255 -335.785 -43.975 ;
        RECT -336.065 -44.855 -335.785 -44.575 ;
        RECT -333.825 -44.255 -333.545 -43.975 ;
        RECT -333.825 -44.855 -333.545 -44.575 ;
        RECT -261.025 -24.095 -260.745 -23.815 ;
        RECT -261.025 -24.695 -260.745 -24.415 ;
        RECT -296.865 -27.455 -296.585 -27.175 ;
        RECT -296.865 -28.055 -296.585 -27.775 ;
        RECT -314.785 -30.815 -314.505 -30.535 ;
        RECT -314.785 -31.415 -314.505 -31.135 ;
        RECT -323.745 -34.175 -323.465 -33.895 ;
        RECT -323.745 -34.775 -323.465 -34.495 ;
        RECT -328.225 -37.535 -327.945 -37.255 ;
        RECT -328.225 -38.135 -327.945 -37.855 ;
        RECT -330.465 -40.895 -330.185 -40.615 ;
        RECT -330.465 -41.495 -330.185 -41.215 ;
        RECT -331.585 -44.255 -331.305 -43.975 ;
        RECT -331.585 -44.855 -331.305 -44.575 ;
        RECT -329.345 -44.255 -329.065 -43.975 ;
        RECT -329.345 -44.855 -329.065 -44.575 ;
        RECT -325.985 -40.895 -325.705 -40.615 ;
        RECT -325.985 -41.495 -325.705 -41.215 ;
        RECT -327.105 -44.255 -326.825 -43.975 ;
        RECT -327.105 -44.855 -326.825 -44.575 ;
        RECT -324.865 -44.255 -324.585 -43.975 ;
        RECT -324.865 -44.855 -324.585 -44.575 ;
        RECT -319.265 -37.535 -318.985 -37.255 ;
        RECT -319.265 -38.135 -318.985 -37.855 ;
        RECT -321.505 -40.895 -321.225 -40.615 ;
        RECT -321.505 -41.495 -321.225 -41.215 ;
        RECT -322.625 -44.255 -322.345 -43.975 ;
        RECT -322.625 -44.855 -322.345 -44.575 ;
        RECT -320.385 -44.255 -320.105 -43.975 ;
        RECT -320.385 -44.855 -320.105 -44.575 ;
        RECT -317.025 -40.895 -316.745 -40.615 ;
        RECT -317.025 -41.495 -316.745 -41.215 ;
        RECT -318.145 -44.255 -317.865 -43.975 ;
        RECT -318.145 -44.855 -317.865 -44.575 ;
        RECT -315.905 -44.255 -315.625 -43.975 ;
        RECT -315.905 -44.855 -315.625 -44.575 ;
        RECT -305.825 -34.175 -305.545 -33.895 ;
        RECT -305.825 -34.775 -305.545 -34.495 ;
        RECT -310.305 -37.535 -310.025 -37.255 ;
        RECT -310.305 -38.135 -310.025 -37.855 ;
        RECT -312.545 -40.895 -312.265 -40.615 ;
        RECT -312.545 -41.495 -312.265 -41.215 ;
        RECT -313.665 -44.255 -313.385 -43.975 ;
        RECT -313.665 -44.855 -313.385 -44.575 ;
        RECT -311.425 -44.255 -311.145 -43.975 ;
        RECT -311.425 -44.855 -311.145 -44.575 ;
        RECT -308.065 -40.895 -307.785 -40.615 ;
        RECT -308.065 -41.495 -307.785 -41.215 ;
        RECT -309.185 -44.255 -308.905 -43.975 ;
        RECT -309.185 -44.855 -308.905 -44.575 ;
        RECT -306.945 -44.255 -306.665 -43.975 ;
        RECT -306.945 -44.855 -306.665 -44.575 ;
        RECT -301.345 -37.535 -301.065 -37.255 ;
        RECT -301.345 -38.135 -301.065 -37.855 ;
        RECT -303.585 -40.895 -303.305 -40.615 ;
        RECT -303.585 -41.495 -303.305 -41.215 ;
        RECT -304.705 -44.255 -304.425 -43.975 ;
        RECT -304.705 -44.855 -304.425 -44.575 ;
        RECT -302.465 -44.255 -302.185 -43.975 ;
        RECT -302.465 -44.855 -302.185 -44.575 ;
        RECT -299.105 -40.895 -298.825 -40.615 ;
        RECT -299.105 -41.495 -298.825 -41.215 ;
        RECT -300.225 -44.255 -299.945 -43.975 ;
        RECT -300.225 -44.855 -299.945 -44.575 ;
        RECT -297.985 -44.255 -297.705 -43.975 ;
        RECT -297.985 -44.855 -297.705 -44.575 ;
        RECT -278.945 -30.815 -278.665 -30.535 ;
        RECT -278.945 -31.415 -278.665 -31.135 ;
        RECT -287.905 -34.175 -287.625 -33.895 ;
        RECT -287.905 -34.775 -287.625 -34.495 ;
        RECT -292.385 -37.535 -292.105 -37.255 ;
        RECT -292.385 -38.135 -292.105 -37.855 ;
        RECT -294.625 -40.895 -294.345 -40.615 ;
        RECT -294.625 -41.495 -294.345 -41.215 ;
        RECT -295.745 -44.255 -295.465 -43.975 ;
        RECT -295.745 -44.855 -295.465 -44.575 ;
        RECT -293.505 -44.255 -293.225 -43.975 ;
        RECT -293.505 -44.855 -293.225 -44.575 ;
        RECT -290.145 -40.895 -289.865 -40.615 ;
        RECT -290.145 -41.495 -289.865 -41.215 ;
        RECT -291.265 -44.255 -290.985 -43.975 ;
        RECT -291.265 -44.855 -290.985 -44.575 ;
        RECT -289.025 -44.255 -288.745 -43.975 ;
        RECT -289.025 -44.855 -288.745 -44.575 ;
        RECT -283.425 -37.535 -283.145 -37.255 ;
        RECT -283.425 -38.135 -283.145 -37.855 ;
        RECT -285.665 -40.895 -285.385 -40.615 ;
        RECT -285.665 -41.495 -285.385 -41.215 ;
        RECT -286.785 -44.255 -286.505 -43.975 ;
        RECT -286.785 -44.855 -286.505 -44.575 ;
        RECT -284.545 -44.255 -284.265 -43.975 ;
        RECT -284.545 -44.855 -284.265 -44.575 ;
        RECT -281.185 -40.895 -280.905 -40.615 ;
        RECT -281.185 -41.495 -280.905 -41.215 ;
        RECT -282.305 -44.255 -282.025 -43.975 ;
        RECT -282.305 -44.855 -282.025 -44.575 ;
        RECT -280.065 -44.255 -279.785 -43.975 ;
        RECT -280.065 -44.855 -279.785 -44.575 ;
        RECT -269.985 -34.175 -269.705 -33.895 ;
        RECT -269.985 -34.775 -269.705 -34.495 ;
        RECT -274.465 -37.535 -274.185 -37.255 ;
        RECT -274.465 -38.135 -274.185 -37.855 ;
        RECT -276.705 -40.895 -276.425 -40.615 ;
        RECT -276.705 -41.495 -276.425 -41.215 ;
        RECT -277.825 -44.255 -277.545 -43.975 ;
        RECT -277.825 -44.855 -277.545 -44.575 ;
        RECT -275.585 -44.255 -275.305 -43.975 ;
        RECT -275.585 -44.855 -275.305 -44.575 ;
        RECT -272.225 -40.895 -271.945 -40.615 ;
        RECT -272.225 -41.495 -271.945 -41.215 ;
        RECT -273.345 -44.255 -273.065 -43.975 ;
        RECT -273.345 -44.855 -273.065 -44.575 ;
        RECT -271.105 -44.255 -270.825 -43.975 ;
        RECT -271.105 -44.855 -270.825 -44.575 ;
        RECT -265.505 -37.535 -265.225 -37.255 ;
        RECT -265.505 -38.135 -265.225 -37.855 ;
        RECT -267.745 -40.895 -267.465 -40.615 ;
        RECT -267.745 -41.495 -267.465 -41.215 ;
        RECT -268.865 -44.255 -268.585 -43.975 ;
        RECT -268.865 -44.855 -268.585 -44.575 ;
        RECT -266.625 -44.255 -266.345 -43.975 ;
        RECT -266.625 -44.855 -266.345 -44.575 ;
        RECT -263.265 -40.895 -262.985 -40.615 ;
        RECT -263.265 -41.495 -262.985 -41.215 ;
        RECT -264.385 -44.255 -264.105 -43.975 ;
        RECT -264.385 -44.855 -264.105 -44.575 ;
        RECT -262.145 -44.255 -261.865 -43.975 ;
        RECT -262.145 -44.855 -261.865 -44.575 ;
        RECT -225.185 -27.455 -224.905 -27.175 ;
        RECT -225.185 -28.055 -224.905 -27.775 ;
        RECT -243.105 -30.815 -242.825 -30.535 ;
        RECT -243.105 -31.415 -242.825 -31.135 ;
        RECT -252.065 -34.175 -251.785 -33.895 ;
        RECT -252.065 -34.775 -251.785 -34.495 ;
        RECT -256.545 -37.535 -256.265 -37.255 ;
        RECT -256.545 -38.135 -256.265 -37.855 ;
        RECT -258.785 -40.895 -258.505 -40.615 ;
        RECT -258.785 -41.495 -258.505 -41.215 ;
        RECT -259.905 -44.255 -259.625 -43.975 ;
        RECT -259.905 -44.855 -259.625 -44.575 ;
        RECT -257.665 -44.255 -257.385 -43.975 ;
        RECT -257.665 -44.855 -257.385 -44.575 ;
        RECT -254.305 -40.895 -254.025 -40.615 ;
        RECT -254.305 -41.495 -254.025 -41.215 ;
        RECT -255.425 -44.255 -255.145 -43.975 ;
        RECT -255.425 -44.855 -255.145 -44.575 ;
        RECT -253.185 -44.255 -252.905 -43.975 ;
        RECT -253.185 -44.855 -252.905 -44.575 ;
        RECT -247.585 -37.535 -247.305 -37.255 ;
        RECT -247.585 -38.135 -247.305 -37.855 ;
        RECT -249.825 -40.895 -249.545 -40.615 ;
        RECT -249.825 -41.495 -249.545 -41.215 ;
        RECT -250.945 -44.255 -250.665 -43.975 ;
        RECT -250.945 -44.855 -250.665 -44.575 ;
        RECT -248.705 -44.255 -248.425 -43.975 ;
        RECT -248.705 -44.855 -248.425 -44.575 ;
        RECT -245.345 -40.895 -245.065 -40.615 ;
        RECT -245.345 -41.495 -245.065 -41.215 ;
        RECT -246.465 -44.255 -246.185 -43.975 ;
        RECT -246.465 -44.855 -246.185 -44.575 ;
        RECT -244.225 -44.255 -243.945 -43.975 ;
        RECT -244.225 -44.855 -243.945 -44.575 ;
        RECT -234.145 -34.175 -233.865 -33.895 ;
        RECT -234.145 -34.775 -233.865 -34.495 ;
        RECT -238.625 -37.535 -238.345 -37.255 ;
        RECT -238.625 -38.135 -238.345 -37.855 ;
        RECT -240.865 -40.895 -240.585 -40.615 ;
        RECT -240.865 -41.495 -240.585 -41.215 ;
        RECT -241.985 -44.255 -241.705 -43.975 ;
        RECT -241.985 -44.855 -241.705 -44.575 ;
        RECT -239.745 -44.255 -239.465 -43.975 ;
        RECT -239.745 -44.855 -239.465 -44.575 ;
        RECT -236.385 -40.895 -236.105 -40.615 ;
        RECT -236.385 -41.495 -236.105 -41.215 ;
        RECT -237.505 -44.255 -237.225 -43.975 ;
        RECT -237.505 -44.855 -237.225 -44.575 ;
        RECT -235.265 -44.255 -234.985 -43.975 ;
        RECT -235.265 -44.855 -234.985 -44.575 ;
        RECT -229.665 -37.535 -229.385 -37.255 ;
        RECT -229.665 -38.135 -229.385 -37.855 ;
        RECT -231.905 -40.895 -231.625 -40.615 ;
        RECT -231.905 -41.495 -231.625 -41.215 ;
        RECT -233.025 -44.255 -232.745 -43.975 ;
        RECT -233.025 -44.855 -232.745 -44.575 ;
        RECT -230.785 -44.255 -230.505 -43.975 ;
        RECT -230.785 -44.855 -230.505 -44.575 ;
        RECT -227.425 -40.895 -227.145 -40.615 ;
        RECT -227.425 -41.495 -227.145 -41.215 ;
        RECT -228.545 -44.255 -228.265 -43.975 ;
        RECT -228.545 -44.855 -228.265 -44.575 ;
        RECT -226.305 -44.255 -226.025 -43.975 ;
        RECT -226.305 -44.855 -226.025 -44.575 ;
        RECT -207.265 -30.815 -206.985 -30.535 ;
        RECT -207.265 -31.415 -206.985 -31.135 ;
        RECT -216.225 -34.175 -215.945 -33.895 ;
        RECT -216.225 -34.775 -215.945 -34.495 ;
        RECT -220.705 -37.535 -220.425 -37.255 ;
        RECT -220.705 -38.135 -220.425 -37.855 ;
        RECT -222.945 -40.895 -222.665 -40.615 ;
        RECT -222.945 -41.495 -222.665 -41.215 ;
        RECT -224.065 -44.255 -223.785 -43.975 ;
        RECT -224.065 -44.855 -223.785 -44.575 ;
        RECT -221.825 -44.255 -221.545 -43.975 ;
        RECT -221.825 -44.855 -221.545 -44.575 ;
        RECT -218.465 -40.895 -218.185 -40.615 ;
        RECT -218.465 -41.495 -218.185 -41.215 ;
        RECT -219.585 -44.255 -219.305 -43.975 ;
        RECT -219.585 -44.855 -219.305 -44.575 ;
        RECT -217.345 -44.255 -217.065 -43.975 ;
        RECT -217.345 -44.855 -217.065 -44.575 ;
        RECT -211.745 -37.535 -211.465 -37.255 ;
        RECT -211.745 -38.135 -211.465 -37.855 ;
        RECT -213.985 -40.895 -213.705 -40.615 ;
        RECT -213.985 -41.495 -213.705 -41.215 ;
        RECT -215.105 -44.255 -214.825 -43.975 ;
        RECT -215.105 -44.855 -214.825 -44.575 ;
        RECT -212.865 -44.255 -212.585 -43.975 ;
        RECT -212.865 -44.855 -212.585 -44.575 ;
        RECT -209.505 -40.895 -209.225 -40.615 ;
        RECT -209.505 -41.495 -209.225 -41.215 ;
        RECT -210.625 -44.255 -210.345 -43.975 ;
        RECT -210.625 -44.855 -210.345 -44.575 ;
        RECT -208.385 -44.255 -208.105 -43.975 ;
        RECT -208.385 -44.855 -208.105 -44.575 ;
        RECT -198.305 -34.175 -198.025 -33.895 ;
        RECT -198.305 -34.775 -198.025 -34.495 ;
        RECT -202.785 -37.535 -202.505 -37.255 ;
        RECT -202.785 -38.135 -202.505 -37.855 ;
        RECT -205.025 -40.895 -204.745 -40.615 ;
        RECT -205.025 -41.495 -204.745 -41.215 ;
        RECT -206.145 -44.255 -205.865 -43.975 ;
        RECT -206.145 -44.855 -205.865 -44.575 ;
        RECT -203.905 -44.255 -203.625 -43.975 ;
        RECT -203.905 -44.855 -203.625 -44.575 ;
        RECT -200.545 -40.895 -200.265 -40.615 ;
        RECT -200.545 -41.495 -200.265 -41.215 ;
        RECT -201.665 -44.255 -201.385 -43.975 ;
        RECT -201.665 -44.855 -201.385 -44.575 ;
        RECT -199.425 -44.255 -199.145 -43.975 ;
        RECT -199.425 -44.855 -199.145 -44.575 ;
        RECT -193.825 -37.535 -193.545 -37.255 ;
        RECT -193.825 -38.135 -193.545 -37.855 ;
        RECT -196.065 -40.895 -195.785 -40.615 ;
        RECT -196.065 -41.495 -195.785 -41.215 ;
        RECT -197.185 -44.255 -196.905 -43.975 ;
        RECT -197.185 -44.855 -196.905 -44.575 ;
        RECT -194.945 -44.255 -194.665 -43.975 ;
        RECT -194.945 -44.855 -194.665 -44.575 ;
        RECT -191.585 -40.895 -191.305 -40.615 ;
        RECT -191.585 -41.495 -191.305 -41.215 ;
        RECT -192.705 -44.255 -192.425 -43.975 ;
        RECT -192.705 -44.855 -192.425 -44.575 ;
        RECT -190.465 -44.255 -190.185 -43.975 ;
        RECT -190.465 -44.855 -190.185 -44.575 ;
        RECT -188.225 -17.375 -187.945 -17.095 ;
        RECT -188.225 -17.975 -187.945 -17.695 ;
        RECT -44.865 -20.735 -44.585 -20.455 ;
        RECT -44.865 -21.335 -44.585 -21.055 ;
        RECT -116.545 -24.095 -116.265 -23.815 ;
        RECT -116.545 -24.695 -116.265 -24.415 ;
        RECT -152.385 -27.455 -152.105 -27.175 ;
        RECT -152.385 -28.055 -152.105 -27.775 ;
        RECT -170.305 -30.815 -170.025 -30.535 ;
        RECT -170.305 -31.415 -170.025 -31.135 ;
        RECT -179.265 -34.175 -178.985 -33.895 ;
        RECT -179.265 -34.775 -178.985 -34.495 ;
        RECT -183.745 -37.535 -183.465 -37.255 ;
        RECT -183.745 -38.135 -183.465 -37.855 ;
        RECT -185.985 -40.895 -185.705 -40.615 ;
        RECT -185.985 -41.495 -185.705 -41.215 ;
        RECT -187.105 -44.255 -186.825 -43.975 ;
        RECT -187.105 -44.855 -186.825 -44.575 ;
        RECT -184.865 -44.255 -184.585 -43.975 ;
        RECT -184.865 -44.855 -184.585 -44.575 ;
        RECT -181.505 -40.895 -181.225 -40.615 ;
        RECT -181.505 -41.495 -181.225 -41.215 ;
        RECT -182.625 -44.255 -182.345 -43.975 ;
        RECT -182.625 -44.855 -182.345 -44.575 ;
        RECT -180.385 -44.255 -180.105 -43.975 ;
        RECT -180.385 -44.855 -180.105 -44.575 ;
        RECT -174.785 -37.535 -174.505 -37.255 ;
        RECT -174.785 -38.135 -174.505 -37.855 ;
        RECT -177.025 -40.895 -176.745 -40.615 ;
        RECT -177.025 -41.495 -176.745 -41.215 ;
        RECT -178.145 -44.255 -177.865 -43.975 ;
        RECT -178.145 -44.855 -177.865 -44.575 ;
        RECT -175.905 -44.255 -175.625 -43.975 ;
        RECT -175.905 -44.855 -175.625 -44.575 ;
        RECT -172.545 -40.895 -172.265 -40.615 ;
        RECT -172.545 -41.495 -172.265 -41.215 ;
        RECT -173.665 -44.255 -173.385 -43.975 ;
        RECT -173.665 -44.855 -173.385 -44.575 ;
        RECT -171.425 -44.255 -171.145 -43.975 ;
        RECT -171.425 -44.855 -171.145 -44.575 ;
        RECT -161.345 -34.175 -161.065 -33.895 ;
        RECT -161.345 -34.775 -161.065 -34.495 ;
        RECT -165.825 -37.535 -165.545 -37.255 ;
        RECT -165.825 -38.135 -165.545 -37.855 ;
        RECT -168.065 -40.895 -167.785 -40.615 ;
        RECT -168.065 -41.495 -167.785 -41.215 ;
        RECT -169.185 -44.255 -168.905 -43.975 ;
        RECT -169.185 -44.855 -168.905 -44.575 ;
        RECT -166.945 -44.255 -166.665 -43.975 ;
        RECT -166.945 -44.855 -166.665 -44.575 ;
        RECT -163.585 -40.895 -163.305 -40.615 ;
        RECT -163.585 -41.495 -163.305 -41.215 ;
        RECT -164.705 -44.255 -164.425 -43.975 ;
        RECT -164.705 -44.855 -164.425 -44.575 ;
        RECT -162.465 -44.255 -162.185 -43.975 ;
        RECT -162.465 -44.855 -162.185 -44.575 ;
        RECT -156.865 -37.535 -156.585 -37.255 ;
        RECT -156.865 -38.135 -156.585 -37.855 ;
        RECT -159.105 -40.895 -158.825 -40.615 ;
        RECT -159.105 -41.495 -158.825 -41.215 ;
        RECT -160.225 -44.255 -159.945 -43.975 ;
        RECT -160.225 -44.855 -159.945 -44.575 ;
        RECT -157.985 -44.255 -157.705 -43.975 ;
        RECT -157.985 -44.855 -157.705 -44.575 ;
        RECT -154.625 -40.895 -154.345 -40.615 ;
        RECT -154.625 -41.495 -154.345 -41.215 ;
        RECT -155.745 -44.255 -155.465 -43.975 ;
        RECT -155.745 -44.855 -155.465 -44.575 ;
        RECT -153.505 -44.255 -153.225 -43.975 ;
        RECT -153.505 -44.855 -153.225 -44.575 ;
        RECT -134.465 -30.815 -134.185 -30.535 ;
        RECT -134.465 -31.415 -134.185 -31.135 ;
        RECT -143.425 -34.175 -143.145 -33.895 ;
        RECT -143.425 -34.775 -143.145 -34.495 ;
        RECT -147.905 -37.535 -147.625 -37.255 ;
        RECT -147.905 -38.135 -147.625 -37.855 ;
        RECT -150.145 -40.895 -149.865 -40.615 ;
        RECT -150.145 -41.495 -149.865 -41.215 ;
        RECT -151.265 -44.255 -150.985 -43.975 ;
        RECT -151.265 -44.855 -150.985 -44.575 ;
        RECT -149.025 -44.255 -148.745 -43.975 ;
        RECT -149.025 -44.855 -148.745 -44.575 ;
        RECT -145.665 -40.895 -145.385 -40.615 ;
        RECT -145.665 -41.495 -145.385 -41.215 ;
        RECT -146.785 -44.255 -146.505 -43.975 ;
        RECT -146.785 -44.855 -146.505 -44.575 ;
        RECT -144.545 -44.255 -144.265 -43.975 ;
        RECT -144.545 -44.855 -144.265 -44.575 ;
        RECT -138.945 -37.535 -138.665 -37.255 ;
        RECT -138.945 -38.135 -138.665 -37.855 ;
        RECT -141.185 -40.895 -140.905 -40.615 ;
        RECT -141.185 -41.495 -140.905 -41.215 ;
        RECT -142.305 -44.255 -142.025 -43.975 ;
        RECT -142.305 -44.855 -142.025 -44.575 ;
        RECT -140.065 -44.255 -139.785 -43.975 ;
        RECT -140.065 -44.855 -139.785 -44.575 ;
        RECT -136.705 -40.895 -136.425 -40.615 ;
        RECT -136.705 -41.495 -136.425 -41.215 ;
        RECT -137.825 -44.255 -137.545 -43.975 ;
        RECT -137.825 -44.855 -137.545 -44.575 ;
        RECT -135.585 -44.255 -135.305 -43.975 ;
        RECT -135.585 -44.855 -135.305 -44.575 ;
        RECT -125.505 -34.175 -125.225 -33.895 ;
        RECT -125.505 -34.775 -125.225 -34.495 ;
        RECT -129.985 -37.535 -129.705 -37.255 ;
        RECT -129.985 -38.135 -129.705 -37.855 ;
        RECT -132.225 -40.895 -131.945 -40.615 ;
        RECT -132.225 -41.495 -131.945 -41.215 ;
        RECT -133.345 -44.255 -133.065 -43.975 ;
        RECT -133.345 -44.855 -133.065 -44.575 ;
        RECT -131.105 -44.255 -130.825 -43.975 ;
        RECT -131.105 -44.855 -130.825 -44.575 ;
        RECT -127.745 -40.895 -127.465 -40.615 ;
        RECT -127.745 -41.495 -127.465 -41.215 ;
        RECT -128.865 -44.255 -128.585 -43.975 ;
        RECT -128.865 -44.855 -128.585 -44.575 ;
        RECT -126.625 -44.255 -126.345 -43.975 ;
        RECT -126.625 -44.855 -126.345 -44.575 ;
        RECT -121.025 -37.535 -120.745 -37.255 ;
        RECT -121.025 -38.135 -120.745 -37.855 ;
        RECT -123.265 -40.895 -122.985 -40.615 ;
        RECT -123.265 -41.495 -122.985 -41.215 ;
        RECT -124.385 -44.255 -124.105 -43.975 ;
        RECT -124.385 -44.855 -124.105 -44.575 ;
        RECT -122.145 -44.255 -121.865 -43.975 ;
        RECT -122.145 -44.855 -121.865 -44.575 ;
        RECT -118.785 -40.895 -118.505 -40.615 ;
        RECT -118.785 -41.495 -118.505 -41.215 ;
        RECT -119.905 -44.255 -119.625 -43.975 ;
        RECT -119.905 -44.855 -119.625 -44.575 ;
        RECT -117.665 -44.255 -117.385 -43.975 ;
        RECT -117.665 -44.855 -117.385 -44.575 ;
        RECT -80.705 -27.455 -80.425 -27.175 ;
        RECT -80.705 -28.055 -80.425 -27.775 ;
        RECT -98.625 -30.815 -98.345 -30.535 ;
        RECT -98.625 -31.415 -98.345 -31.135 ;
        RECT -107.585 -34.175 -107.305 -33.895 ;
        RECT -107.585 -34.775 -107.305 -34.495 ;
        RECT -112.065 -37.535 -111.785 -37.255 ;
        RECT -112.065 -38.135 -111.785 -37.855 ;
        RECT -114.305 -40.895 -114.025 -40.615 ;
        RECT -114.305 -41.495 -114.025 -41.215 ;
        RECT -115.425 -44.255 -115.145 -43.975 ;
        RECT -115.425 -44.855 -115.145 -44.575 ;
        RECT -113.185 -44.255 -112.905 -43.975 ;
        RECT -113.185 -44.855 -112.905 -44.575 ;
        RECT -109.825 -40.895 -109.545 -40.615 ;
        RECT -109.825 -41.495 -109.545 -41.215 ;
        RECT -110.945 -44.255 -110.665 -43.975 ;
        RECT -110.945 -44.855 -110.665 -44.575 ;
        RECT -108.705 -44.255 -108.425 -43.975 ;
        RECT -108.705 -44.855 -108.425 -44.575 ;
        RECT -103.105 -37.535 -102.825 -37.255 ;
        RECT -103.105 -38.135 -102.825 -37.855 ;
        RECT -105.345 -40.895 -105.065 -40.615 ;
        RECT -105.345 -41.495 -105.065 -41.215 ;
        RECT -106.465 -44.255 -106.185 -43.975 ;
        RECT -106.465 -44.855 -106.185 -44.575 ;
        RECT -104.225 -44.255 -103.945 -43.975 ;
        RECT -104.225 -44.855 -103.945 -44.575 ;
        RECT -100.865 -40.895 -100.585 -40.615 ;
        RECT -100.865 -41.495 -100.585 -41.215 ;
        RECT -101.985 -44.255 -101.705 -43.975 ;
        RECT -101.985 -44.855 -101.705 -44.575 ;
        RECT -99.745 -44.255 -99.465 -43.975 ;
        RECT -99.745 -44.855 -99.465 -44.575 ;
        RECT -89.665 -34.175 -89.385 -33.895 ;
        RECT -89.665 -34.775 -89.385 -34.495 ;
        RECT -94.145 -37.535 -93.865 -37.255 ;
        RECT -94.145 -38.135 -93.865 -37.855 ;
        RECT -96.385 -40.895 -96.105 -40.615 ;
        RECT -96.385 -41.495 -96.105 -41.215 ;
        RECT -97.505 -44.255 -97.225 -43.975 ;
        RECT -97.505 -44.855 -97.225 -44.575 ;
        RECT -95.265 -44.255 -94.985 -43.975 ;
        RECT -95.265 -44.855 -94.985 -44.575 ;
        RECT -91.905 -40.895 -91.625 -40.615 ;
        RECT -91.905 -41.495 -91.625 -41.215 ;
        RECT -93.025 -44.255 -92.745 -43.975 ;
        RECT -93.025 -44.855 -92.745 -44.575 ;
        RECT -90.785 -44.255 -90.505 -43.975 ;
        RECT -90.785 -44.855 -90.505 -44.575 ;
        RECT -85.185 -37.535 -84.905 -37.255 ;
        RECT -85.185 -38.135 -84.905 -37.855 ;
        RECT -87.425 -40.895 -87.145 -40.615 ;
        RECT -87.425 -41.495 -87.145 -41.215 ;
        RECT -88.545 -44.255 -88.265 -43.975 ;
        RECT -88.545 -44.855 -88.265 -44.575 ;
        RECT -86.305 -44.255 -86.025 -43.975 ;
        RECT -86.305 -44.855 -86.025 -44.575 ;
        RECT -82.945 -40.895 -82.665 -40.615 ;
        RECT -82.945 -41.495 -82.665 -41.215 ;
        RECT -84.065 -44.255 -83.785 -43.975 ;
        RECT -84.065 -44.855 -83.785 -44.575 ;
        RECT -81.825 -44.255 -81.545 -43.975 ;
        RECT -81.825 -44.855 -81.545 -44.575 ;
        RECT -62.785 -30.815 -62.505 -30.535 ;
        RECT -62.785 -31.415 -62.505 -31.135 ;
        RECT -71.745 -34.175 -71.465 -33.895 ;
        RECT -71.745 -34.775 -71.465 -34.495 ;
        RECT -76.225 -37.535 -75.945 -37.255 ;
        RECT -76.225 -38.135 -75.945 -37.855 ;
        RECT -78.465 -40.895 -78.185 -40.615 ;
        RECT -78.465 -41.495 -78.185 -41.215 ;
        RECT -79.585 -44.255 -79.305 -43.975 ;
        RECT -79.585 -44.855 -79.305 -44.575 ;
        RECT -77.345 -44.255 -77.065 -43.975 ;
        RECT -77.345 -44.855 -77.065 -44.575 ;
        RECT -73.985 -40.895 -73.705 -40.615 ;
        RECT -73.985 -41.495 -73.705 -41.215 ;
        RECT -75.105 -44.255 -74.825 -43.975 ;
        RECT -75.105 -44.855 -74.825 -44.575 ;
        RECT -72.865 -44.255 -72.585 -43.975 ;
        RECT -72.865 -44.855 -72.585 -44.575 ;
        RECT -67.265 -37.535 -66.985 -37.255 ;
        RECT -67.265 -38.135 -66.985 -37.855 ;
        RECT -69.505 -40.895 -69.225 -40.615 ;
        RECT -69.505 -41.495 -69.225 -41.215 ;
        RECT -70.625 -44.255 -70.345 -43.975 ;
        RECT -70.625 -44.855 -70.345 -44.575 ;
        RECT -68.385 -44.255 -68.105 -43.975 ;
        RECT -68.385 -44.855 -68.105 -44.575 ;
        RECT -65.025 -40.895 -64.745 -40.615 ;
        RECT -65.025 -41.495 -64.745 -41.215 ;
        RECT -66.145 -44.255 -65.865 -43.975 ;
        RECT -66.145 -44.855 -65.865 -44.575 ;
        RECT -63.905 -44.255 -63.625 -43.975 ;
        RECT -63.905 -44.855 -63.625 -44.575 ;
        RECT -53.825 -34.175 -53.545 -33.895 ;
        RECT -53.825 -34.775 -53.545 -34.495 ;
        RECT -58.305 -37.535 -58.025 -37.255 ;
        RECT -58.305 -38.135 -58.025 -37.855 ;
        RECT -60.545 -40.895 -60.265 -40.615 ;
        RECT -60.545 -41.495 -60.265 -41.215 ;
        RECT -61.665 -44.255 -61.385 -43.975 ;
        RECT -61.665 -44.855 -61.385 -44.575 ;
        RECT -59.425 -44.255 -59.145 -43.975 ;
        RECT -59.425 -44.855 -59.145 -44.575 ;
        RECT -56.065 -40.895 -55.785 -40.615 ;
        RECT -56.065 -41.495 -55.785 -41.215 ;
        RECT -57.185 -44.255 -56.905 -43.975 ;
        RECT -57.185 -44.855 -56.905 -44.575 ;
        RECT -54.945 -44.255 -54.665 -43.975 ;
        RECT -54.945 -44.855 -54.665 -44.575 ;
        RECT -49.345 -37.535 -49.065 -37.255 ;
        RECT -49.345 -38.135 -49.065 -37.855 ;
        RECT -51.585 -40.895 -51.305 -40.615 ;
        RECT -51.585 -41.495 -51.305 -41.215 ;
        RECT -52.705 -44.255 -52.425 -43.975 ;
        RECT -52.705 -44.855 -52.425 -44.575 ;
        RECT -50.465 -44.255 -50.185 -43.975 ;
        RECT -50.465 -44.855 -50.185 -44.575 ;
        RECT -47.105 -40.895 -46.825 -40.615 ;
        RECT -47.105 -41.495 -46.825 -41.215 ;
        RECT -48.225 -44.255 -47.945 -43.975 ;
        RECT -48.225 -44.855 -47.945 -44.575 ;
        RECT -45.985 -44.255 -45.705 -43.975 ;
        RECT -45.985 -44.855 -45.705 -44.575 ;
        RECT 26.815 -24.095 27.095 -23.815 ;
        RECT 26.815 -24.695 27.095 -24.415 ;
        RECT -9.025 -27.455 -8.745 -27.175 ;
        RECT -9.025 -28.055 -8.745 -27.775 ;
        RECT -26.945 -30.815 -26.665 -30.535 ;
        RECT -26.945 -31.415 -26.665 -31.135 ;
        RECT -35.905 -34.175 -35.625 -33.895 ;
        RECT -35.905 -34.775 -35.625 -34.495 ;
        RECT -40.385 -37.535 -40.105 -37.255 ;
        RECT -40.385 -38.135 -40.105 -37.855 ;
        RECT -42.625 -40.895 -42.345 -40.615 ;
        RECT -42.625 -41.495 -42.345 -41.215 ;
        RECT -43.745 -44.255 -43.465 -43.975 ;
        RECT -43.745 -44.855 -43.465 -44.575 ;
        RECT -41.505 -44.255 -41.225 -43.975 ;
        RECT -41.505 -44.855 -41.225 -44.575 ;
        RECT -38.145 -40.895 -37.865 -40.615 ;
        RECT -38.145 -41.495 -37.865 -41.215 ;
        RECT -39.265 -44.255 -38.985 -43.975 ;
        RECT -39.265 -44.855 -38.985 -44.575 ;
        RECT -37.025 -44.255 -36.745 -43.975 ;
        RECT -37.025 -44.855 -36.745 -44.575 ;
        RECT -31.425 -37.535 -31.145 -37.255 ;
        RECT -31.425 -38.135 -31.145 -37.855 ;
        RECT -33.665 -40.895 -33.385 -40.615 ;
        RECT -33.665 -41.495 -33.385 -41.215 ;
        RECT -34.785 -44.255 -34.505 -43.975 ;
        RECT -34.785 -44.855 -34.505 -44.575 ;
        RECT -32.545 -44.255 -32.265 -43.975 ;
        RECT -32.545 -44.855 -32.265 -44.575 ;
        RECT -29.185 -40.895 -28.905 -40.615 ;
        RECT -29.185 -41.495 -28.905 -41.215 ;
        RECT -30.305 -44.255 -30.025 -43.975 ;
        RECT -30.305 -44.855 -30.025 -44.575 ;
        RECT -28.065 -44.255 -27.785 -43.975 ;
        RECT -28.065 -44.855 -27.785 -44.575 ;
        RECT -17.985 -34.175 -17.705 -33.895 ;
        RECT -17.985 -34.775 -17.705 -34.495 ;
        RECT -22.465 -37.535 -22.185 -37.255 ;
        RECT -22.465 -38.135 -22.185 -37.855 ;
        RECT -24.705 -40.895 -24.425 -40.615 ;
        RECT -24.705 -41.495 -24.425 -41.215 ;
        RECT -25.825 -44.255 -25.545 -43.975 ;
        RECT -25.825 -44.855 -25.545 -44.575 ;
        RECT -23.585 -44.255 -23.305 -43.975 ;
        RECT -23.585 -44.855 -23.305 -44.575 ;
        RECT -20.225 -40.895 -19.945 -40.615 ;
        RECT -20.225 -41.495 -19.945 -41.215 ;
        RECT -21.345 -44.255 -21.065 -43.975 ;
        RECT -21.345 -44.855 -21.065 -44.575 ;
        RECT -19.105 -44.255 -18.825 -43.975 ;
        RECT -19.105 -44.855 -18.825 -44.575 ;
        RECT -13.505 -37.535 -13.225 -37.255 ;
        RECT -13.505 -38.135 -13.225 -37.855 ;
        RECT -15.745 -40.895 -15.465 -40.615 ;
        RECT -15.745 -41.495 -15.465 -41.215 ;
        RECT -16.865 -44.255 -16.585 -43.975 ;
        RECT -16.865 -44.855 -16.585 -44.575 ;
        RECT -14.625 -44.255 -14.345 -43.975 ;
        RECT -14.625 -44.855 -14.345 -44.575 ;
        RECT -11.265 -40.895 -10.985 -40.615 ;
        RECT -11.265 -41.495 -10.985 -41.215 ;
        RECT -12.385 -44.255 -12.105 -43.975 ;
        RECT -12.385 -44.855 -12.105 -44.575 ;
        RECT -10.145 -44.255 -9.865 -43.975 ;
        RECT -10.145 -44.855 -9.865 -44.575 ;
        RECT 8.895 -30.815 9.175 -30.535 ;
        RECT 8.895 -31.415 9.175 -31.135 ;
        RECT -0.065 -34.175 0.215 -33.895 ;
        RECT -0.065 -34.775 0.215 -34.495 ;
        RECT -4.545 -37.535 -4.265 -37.255 ;
        RECT -4.545 -38.135 -4.265 -37.855 ;
        RECT -6.785 -40.895 -6.505 -40.615 ;
        RECT -6.785 -41.495 -6.505 -41.215 ;
        RECT -7.905 -44.255 -7.625 -43.975 ;
        RECT -7.905 -44.855 -7.625 -44.575 ;
        RECT -5.665 -44.255 -5.385 -43.975 ;
        RECT -5.665 -44.855 -5.385 -44.575 ;
        RECT -2.305 -40.895 -2.025 -40.615 ;
        RECT -2.305 -41.495 -2.025 -41.215 ;
        RECT -3.425 -44.255 -3.145 -43.975 ;
        RECT -3.425 -44.855 -3.145 -44.575 ;
        RECT -1.185 -44.255 -0.905 -43.975 ;
        RECT -1.185 -44.855 -0.905 -44.575 ;
        RECT 4.415 -37.535 4.695 -37.255 ;
        RECT 4.415 -38.135 4.695 -37.855 ;
        RECT 2.175 -40.895 2.455 -40.615 ;
        RECT 2.175 -41.495 2.455 -41.215 ;
        RECT 1.055 -44.255 1.335 -43.975 ;
        RECT 1.055 -44.855 1.335 -44.575 ;
        RECT 3.295 -44.255 3.575 -43.975 ;
        RECT 3.295 -44.855 3.575 -44.575 ;
        RECT 6.655 -40.895 6.935 -40.615 ;
        RECT 6.655 -41.495 6.935 -41.215 ;
        RECT 5.535 -44.255 5.815 -43.975 ;
        RECT 5.535 -44.855 5.815 -44.575 ;
        RECT 7.775 -44.255 8.055 -43.975 ;
        RECT 7.775 -44.855 8.055 -44.575 ;
        RECT 17.855 -34.175 18.135 -33.895 ;
        RECT 17.855 -34.775 18.135 -34.495 ;
        RECT 13.375 -37.535 13.655 -37.255 ;
        RECT 13.375 -38.135 13.655 -37.855 ;
        RECT 11.135 -40.895 11.415 -40.615 ;
        RECT 11.135 -41.495 11.415 -41.215 ;
        RECT 10.015 -44.255 10.295 -43.975 ;
        RECT 10.015 -44.855 10.295 -44.575 ;
        RECT 12.255 -44.255 12.535 -43.975 ;
        RECT 12.255 -44.855 12.535 -44.575 ;
        RECT 15.615 -40.895 15.895 -40.615 ;
        RECT 15.615 -41.495 15.895 -41.215 ;
        RECT 14.495 -44.255 14.775 -43.975 ;
        RECT 14.495 -44.855 14.775 -44.575 ;
        RECT 16.735 -44.255 17.015 -43.975 ;
        RECT 16.735 -44.855 17.015 -44.575 ;
        RECT 22.335 -37.535 22.615 -37.255 ;
        RECT 22.335 -38.135 22.615 -37.855 ;
        RECT 20.095 -40.895 20.375 -40.615 ;
        RECT 20.095 -41.495 20.375 -41.215 ;
        RECT 18.975 -44.255 19.255 -43.975 ;
        RECT 18.975 -44.855 19.255 -44.575 ;
        RECT 21.215 -44.255 21.495 -43.975 ;
        RECT 21.215 -44.855 21.495 -44.575 ;
        RECT 24.575 -40.895 24.855 -40.615 ;
        RECT 24.575 -41.495 24.855 -41.215 ;
        RECT 23.455 -44.255 23.735 -43.975 ;
        RECT 23.455 -44.855 23.735 -44.575 ;
        RECT 25.695 -44.255 25.975 -43.975 ;
        RECT 25.695 -44.855 25.975 -44.575 ;
        RECT 62.655 -27.455 62.935 -27.175 ;
        RECT 62.655 -28.055 62.935 -27.775 ;
        RECT 44.735 -30.815 45.015 -30.535 ;
        RECT 44.735 -31.415 45.015 -31.135 ;
        RECT 35.775 -34.175 36.055 -33.895 ;
        RECT 35.775 -34.775 36.055 -34.495 ;
        RECT 31.295 -37.535 31.575 -37.255 ;
        RECT 31.295 -38.135 31.575 -37.855 ;
        RECT 29.055 -40.895 29.335 -40.615 ;
        RECT 29.055 -41.495 29.335 -41.215 ;
        RECT 27.935 -44.255 28.215 -43.975 ;
        RECT 27.935 -44.855 28.215 -44.575 ;
        RECT 30.175 -44.255 30.455 -43.975 ;
        RECT 30.175 -44.855 30.455 -44.575 ;
        RECT 33.535 -40.895 33.815 -40.615 ;
        RECT 33.535 -41.495 33.815 -41.215 ;
        RECT 32.415 -44.255 32.695 -43.975 ;
        RECT 32.415 -44.855 32.695 -44.575 ;
        RECT 34.655 -44.255 34.935 -43.975 ;
        RECT 34.655 -44.855 34.935 -44.575 ;
        RECT 40.255 -37.535 40.535 -37.255 ;
        RECT 40.255 -38.135 40.535 -37.855 ;
        RECT 38.015 -40.895 38.295 -40.615 ;
        RECT 38.015 -41.495 38.295 -41.215 ;
        RECT 36.895 -44.255 37.175 -43.975 ;
        RECT 36.895 -44.855 37.175 -44.575 ;
        RECT 39.135 -44.255 39.415 -43.975 ;
        RECT 39.135 -44.855 39.415 -44.575 ;
        RECT 42.495 -40.895 42.775 -40.615 ;
        RECT 42.495 -41.495 42.775 -41.215 ;
        RECT 41.375 -44.255 41.655 -43.975 ;
        RECT 41.375 -44.855 41.655 -44.575 ;
        RECT 43.615 -44.255 43.895 -43.975 ;
        RECT 43.615 -44.855 43.895 -44.575 ;
        RECT 53.695 -34.175 53.975 -33.895 ;
        RECT 53.695 -34.775 53.975 -34.495 ;
        RECT 49.215 -37.535 49.495 -37.255 ;
        RECT 49.215 -38.135 49.495 -37.855 ;
        RECT 46.975 -40.895 47.255 -40.615 ;
        RECT 46.975 -41.495 47.255 -41.215 ;
        RECT 45.855 -44.255 46.135 -43.975 ;
        RECT 45.855 -44.855 46.135 -44.575 ;
        RECT 48.095 -44.255 48.375 -43.975 ;
        RECT 48.095 -44.855 48.375 -44.575 ;
        RECT 51.455 -40.895 51.735 -40.615 ;
        RECT 51.455 -41.495 51.735 -41.215 ;
        RECT 50.335 -44.255 50.615 -43.975 ;
        RECT 50.335 -44.855 50.615 -44.575 ;
        RECT 52.575 -44.255 52.855 -43.975 ;
        RECT 52.575 -44.855 52.855 -44.575 ;
        RECT 58.175 -37.535 58.455 -37.255 ;
        RECT 58.175 -38.135 58.455 -37.855 ;
        RECT 55.935 -40.895 56.215 -40.615 ;
        RECT 55.935 -41.495 56.215 -41.215 ;
        RECT 54.815 -44.255 55.095 -43.975 ;
        RECT 54.815 -44.855 55.095 -44.575 ;
        RECT 57.055 -44.255 57.335 -43.975 ;
        RECT 57.055 -44.855 57.335 -44.575 ;
        RECT 60.415 -40.895 60.695 -40.615 ;
        RECT 60.415 -41.495 60.695 -41.215 ;
        RECT 59.295 -44.255 59.575 -43.975 ;
        RECT 59.295 -44.855 59.575 -44.575 ;
        RECT 61.535 -44.255 61.815 -43.975 ;
        RECT 61.535 -44.855 61.815 -44.575 ;
        RECT 80.575 -30.815 80.855 -30.535 ;
        RECT 80.575 -31.415 80.855 -31.135 ;
        RECT 71.615 -34.175 71.895 -33.895 ;
        RECT 71.615 -34.775 71.895 -34.495 ;
        RECT 67.135 -37.535 67.415 -37.255 ;
        RECT 67.135 -38.135 67.415 -37.855 ;
        RECT 64.895 -40.895 65.175 -40.615 ;
        RECT 64.895 -41.495 65.175 -41.215 ;
        RECT 63.775 -44.255 64.055 -43.975 ;
        RECT 63.775 -44.855 64.055 -44.575 ;
        RECT 66.015 -44.255 66.295 -43.975 ;
        RECT 66.015 -44.855 66.295 -44.575 ;
        RECT 69.375 -40.895 69.655 -40.615 ;
        RECT 69.375 -41.495 69.655 -41.215 ;
        RECT 68.255 -44.255 68.535 -43.975 ;
        RECT 68.255 -44.855 68.535 -44.575 ;
        RECT 70.495 -44.255 70.775 -43.975 ;
        RECT 70.495 -44.855 70.775 -44.575 ;
        RECT 76.095 -37.535 76.375 -37.255 ;
        RECT 76.095 -38.135 76.375 -37.855 ;
        RECT 73.855 -40.895 74.135 -40.615 ;
        RECT 73.855 -41.495 74.135 -41.215 ;
        RECT 72.735 -44.255 73.015 -43.975 ;
        RECT 72.735 -44.855 73.015 -44.575 ;
        RECT 74.975 -44.255 75.255 -43.975 ;
        RECT 74.975 -44.855 75.255 -44.575 ;
        RECT 78.335 -40.895 78.615 -40.615 ;
        RECT 78.335 -41.495 78.615 -41.215 ;
        RECT 77.215 -44.255 77.495 -43.975 ;
        RECT 77.215 -44.855 77.495 -44.575 ;
        RECT 79.455 -44.255 79.735 -43.975 ;
        RECT 79.455 -44.855 79.735 -44.575 ;
        RECT 89.535 -34.175 89.815 -33.895 ;
        RECT 89.535 -34.775 89.815 -34.495 ;
        RECT 85.055 -37.535 85.335 -37.255 ;
        RECT 85.055 -38.135 85.335 -37.855 ;
        RECT 82.815 -40.895 83.095 -40.615 ;
        RECT 82.815 -41.495 83.095 -41.215 ;
        RECT 81.695 -44.255 81.975 -43.975 ;
        RECT 81.695 -44.855 81.975 -44.575 ;
        RECT 83.935 -44.255 84.215 -43.975 ;
        RECT 83.935 -44.855 84.215 -44.575 ;
        RECT 87.295 -40.895 87.575 -40.615 ;
        RECT 87.295 -41.495 87.575 -41.215 ;
        RECT 86.175 -44.255 86.455 -43.975 ;
        RECT 86.175 -44.855 86.455 -44.575 ;
        RECT 88.415 -44.255 88.695 -43.975 ;
        RECT 88.415 -44.855 88.695 -44.575 ;
        RECT 94.015 -37.535 94.295 -37.255 ;
        RECT 94.015 -38.135 94.295 -37.855 ;
        RECT 91.775 -40.895 92.055 -40.615 ;
        RECT 91.775 -41.495 92.055 -41.215 ;
        RECT 90.655 -44.255 90.935 -43.975 ;
        RECT 90.655 -44.855 90.935 -44.575 ;
        RECT 92.895 -44.255 93.175 -43.975 ;
        RECT 92.895 -44.855 93.175 -44.575 ;
        RECT 96.255 -40.895 96.535 -40.615 ;
        RECT 96.255 -41.495 96.535 -41.215 ;
        RECT 95.135 -44.255 95.415 -43.975 ;
        RECT 95.135 -44.855 95.415 -44.575 ;
        RECT 97.375 -44.255 97.655 -43.975 ;
        RECT 97.375 -44.855 97.655 -44.575 ;
        RECT 287.250 -15.300 287.530 -15.020 ;
        RECT 287.810 -15.300 288.090 -15.020 ;
        RECT 288.370 -15.300 288.650 -15.020 ;
        RECT 287.250 -15.860 287.530 -15.580 ;
        RECT 287.810 -15.860 288.090 -15.580 ;
        RECT 288.370 -15.860 288.650 -15.580 ;
        RECT 302.780 25.860 303.060 26.140 ;
        RECT 302.780 19.140 303.060 19.420 ;
        RECT 302.220 7.380 302.500 7.660 ;
        RECT 301.660 3.460 301.940 3.740 ;
        RECT 305.580 7.380 305.860 7.660 ;
        RECT 303.900 6.820 304.180 7.100 ;
        RECT 308.380 11.300 308.660 11.580 ;
        RECT 307.260 6.820 307.540 7.100 ;
        RECT 308.380 5.140 308.660 5.420 ;
        RECT 308.940 9.620 309.220 9.900 ;
        RECT 303.900 4.580 304.180 4.860 ;
        RECT 306.140 4.020 306.420 4.300 ;
        RECT 300.540 -3.260 300.820 -2.980 ;
        RECT 298.860 -15.580 299.140 -15.300 ;
        RECT 298.300 -20.620 298.580 -20.340 ;
        RECT 287.250 -25.380 287.530 -25.100 ;
        RECT 287.810 -25.380 288.090 -25.100 ;
        RECT 288.370 -25.380 288.650 -25.100 ;
        RECT 287.250 -25.940 287.530 -25.660 ;
        RECT 287.810 -25.940 288.090 -25.660 ;
        RECT 288.370 -25.940 288.650 -25.660 ;
        RECT 298.860 -25.660 299.140 -25.380 ;
        RECT 305.020 0.660 305.300 0.940 ;
        RECT 303.900 -16.700 304.180 -16.420 ;
        RECT 304.460 -4.380 304.740 -4.100 ;
        RECT 302.780 -17.260 303.060 -16.980 ;
        RECT 305.580 -8.300 305.860 -8.020 ;
        RECT 308.380 -8.300 308.660 -8.020 ;
        RECT 305.580 -15.580 305.860 -15.300 ;
        RECT 310.620 41.540 310.900 41.820 ;
        RECT 314.540 41.540 314.820 41.820 ;
        RECT 312.300 11.300 312.580 11.580 ;
        RECT 310.620 9.620 310.900 9.900 ;
        RECT 310.620 7.380 310.900 7.660 ;
        RECT 310.060 6.820 310.340 7.100 ;
        RECT 312.860 6.260 313.140 6.540 ;
        RECT 311.180 5.140 311.460 5.420 ;
        RECT 310.060 3.460 310.340 3.740 ;
        RECT 309.500 -16.700 309.780 -16.420 ;
        RECT 304.460 -20.060 304.740 -19.780 ;
        RECT 306.700 -23.420 306.980 -23.140 ;
        RECT 308.940 -20.620 309.220 -20.340 ;
        RECT 301.100 -23.980 301.380 -23.700 ;
        RECT 308.380 -23.980 308.660 -23.700 ;
        RECT 300.540 -30.140 300.820 -29.860 ;
        RECT 301.660 -30.700 301.940 -30.420 ;
        RECT 299.980 -31.820 300.260 -31.540 ;
        RECT 287.250 -35.460 287.530 -35.180 ;
        RECT 287.810 -35.460 288.090 -35.180 ;
        RECT 288.370 -35.460 288.650 -35.180 ;
        RECT 303.900 -31.260 304.180 -30.980 ;
        RECT 287.250 -36.020 287.530 -35.740 ;
        RECT 287.810 -36.020 288.090 -35.740 ;
        RECT 288.370 -36.020 288.650 -35.740 ;
        RECT 301.660 -35.740 301.940 -35.460 ;
        RECT 308.940 -36.300 309.220 -36.020 ;
        RECT 298.860 -44.700 299.140 -44.420 ;
        RECT 287.250 -45.540 287.530 -45.260 ;
        RECT 287.810 -45.540 288.090 -45.260 ;
        RECT 288.370 -45.540 288.650 -45.260 ;
        RECT 287.250 -46.100 287.530 -45.820 ;
        RECT 287.810 -46.100 288.090 -45.820 ;
        RECT 288.370 -46.100 288.650 -45.820 ;
        RECT 287.250 -55.620 287.530 -55.340 ;
        RECT 287.810 -55.620 288.090 -55.340 ;
        RECT 288.370 -55.620 288.650 -55.340 ;
        RECT -474.945 -67.115 -474.665 -66.835 ;
        RECT -474.945 -67.715 -474.665 -67.435 ;
        RECT -472.705 -67.115 -472.425 -66.835 ;
        RECT -472.705 -67.715 -472.425 -67.435 ;
        RECT -473.825 -70.475 -473.545 -70.195 ;
        RECT -473.825 -71.075 -473.545 -70.795 ;
        RECT -470.465 -67.115 -470.185 -66.835 ;
        RECT -470.465 -67.715 -470.185 -67.435 ;
        RECT -468.225 -67.115 -467.945 -66.835 ;
        RECT -468.225 -67.715 -467.945 -67.435 ;
        RECT -469.345 -70.475 -469.065 -70.195 ;
        RECT -469.345 -71.075 -469.065 -70.795 ;
        RECT -471.585 -73.835 -471.305 -73.555 ;
        RECT -471.585 -74.435 -471.305 -74.155 ;
        RECT -465.985 -67.115 -465.705 -66.835 ;
        RECT -465.985 -67.715 -465.705 -67.435 ;
        RECT -463.745 -67.115 -463.465 -66.835 ;
        RECT -463.745 -67.715 -463.465 -67.435 ;
        RECT -464.865 -70.475 -464.585 -70.195 ;
        RECT -464.865 -71.075 -464.585 -70.795 ;
        RECT -461.505 -67.115 -461.225 -66.835 ;
        RECT -461.505 -67.715 -461.225 -67.435 ;
        RECT -459.265 -67.115 -458.985 -66.835 ;
        RECT -459.265 -67.715 -458.985 -67.435 ;
        RECT -460.385 -70.475 -460.105 -70.195 ;
        RECT -460.385 -71.075 -460.105 -70.795 ;
        RECT -462.625 -73.835 -462.345 -73.555 ;
        RECT -462.625 -74.435 -462.345 -74.155 ;
        RECT -467.105 -77.195 -466.825 -76.915 ;
        RECT -467.105 -77.795 -466.825 -77.515 ;
        RECT -457.025 -67.115 -456.745 -66.835 ;
        RECT -457.025 -67.715 -456.745 -67.435 ;
        RECT -454.785 -67.115 -454.505 -66.835 ;
        RECT -454.785 -67.715 -454.505 -67.435 ;
        RECT -455.905 -70.475 -455.625 -70.195 ;
        RECT -455.905 -71.075 -455.625 -70.795 ;
        RECT -452.545 -67.115 -452.265 -66.835 ;
        RECT -452.545 -67.715 -452.265 -67.435 ;
        RECT -450.305 -67.115 -450.025 -66.835 ;
        RECT -450.305 -67.715 -450.025 -67.435 ;
        RECT -451.425 -70.475 -451.145 -70.195 ;
        RECT -451.425 -71.075 -451.145 -70.795 ;
        RECT -453.665 -73.835 -453.385 -73.555 ;
        RECT -453.665 -74.435 -453.385 -74.155 ;
        RECT -448.065 -67.115 -447.785 -66.835 ;
        RECT -448.065 -67.715 -447.785 -67.435 ;
        RECT -445.825 -67.115 -445.545 -66.835 ;
        RECT -445.825 -67.715 -445.545 -67.435 ;
        RECT -446.945 -70.475 -446.665 -70.195 ;
        RECT -446.945 -71.075 -446.665 -70.795 ;
        RECT -443.585 -67.115 -443.305 -66.835 ;
        RECT -443.585 -67.715 -443.305 -67.435 ;
        RECT -441.345 -67.115 -441.065 -66.835 ;
        RECT -441.345 -67.715 -441.065 -67.435 ;
        RECT -442.465 -70.475 -442.185 -70.195 ;
        RECT -442.465 -71.075 -442.185 -70.795 ;
        RECT -444.705 -73.835 -444.425 -73.555 ;
        RECT -444.705 -74.435 -444.425 -74.155 ;
        RECT -449.185 -77.195 -448.905 -76.915 ;
        RECT -449.185 -77.795 -448.905 -77.515 ;
        RECT -458.145 -80.555 -457.865 -80.275 ;
        RECT -458.145 -81.155 -457.865 -80.875 ;
        RECT -486.895 -83.115 -486.615 -81.275 ;
        RECT -497.475 -83.705 -495.635 -83.425 ;
        RECT -439.105 -67.115 -438.825 -66.835 ;
        RECT -439.105 -67.715 -438.825 -67.435 ;
        RECT -436.865 -67.115 -436.585 -66.835 ;
        RECT -436.865 -67.715 -436.585 -67.435 ;
        RECT -437.985 -70.475 -437.705 -70.195 ;
        RECT -437.985 -71.075 -437.705 -70.795 ;
        RECT -434.625 -67.115 -434.345 -66.835 ;
        RECT -434.625 -67.715 -434.345 -67.435 ;
        RECT -432.385 -67.115 -432.105 -66.835 ;
        RECT -432.385 -67.715 -432.105 -67.435 ;
        RECT -433.505 -70.475 -433.225 -70.195 ;
        RECT -433.505 -71.075 -433.225 -70.795 ;
        RECT -435.745 -73.835 -435.465 -73.555 ;
        RECT -435.745 -74.435 -435.465 -74.155 ;
        RECT -430.145 -67.115 -429.865 -66.835 ;
        RECT -430.145 -67.715 -429.865 -67.435 ;
        RECT -427.905 -67.115 -427.625 -66.835 ;
        RECT -427.905 -67.715 -427.625 -67.435 ;
        RECT -429.025 -70.475 -428.745 -70.195 ;
        RECT -429.025 -71.075 -428.745 -70.795 ;
        RECT -425.665 -67.115 -425.385 -66.835 ;
        RECT -425.665 -67.715 -425.385 -67.435 ;
        RECT -423.425 -67.115 -423.145 -66.835 ;
        RECT -423.425 -67.715 -423.145 -67.435 ;
        RECT -424.545 -70.475 -424.265 -70.195 ;
        RECT -424.545 -71.075 -424.265 -70.795 ;
        RECT -426.785 -73.835 -426.505 -73.555 ;
        RECT -426.785 -74.435 -426.505 -74.155 ;
        RECT -431.265 -77.195 -430.985 -76.915 ;
        RECT -431.265 -77.795 -430.985 -77.515 ;
        RECT -421.185 -67.115 -420.905 -66.835 ;
        RECT -421.185 -67.715 -420.905 -67.435 ;
        RECT -418.945 -67.115 -418.665 -66.835 ;
        RECT -418.945 -67.715 -418.665 -67.435 ;
        RECT -420.065 -70.475 -419.785 -70.195 ;
        RECT -420.065 -71.075 -419.785 -70.795 ;
        RECT -416.705 -67.115 -416.425 -66.835 ;
        RECT -416.705 -67.715 -416.425 -67.435 ;
        RECT -414.465 -67.115 -414.185 -66.835 ;
        RECT -414.465 -67.715 -414.185 -67.435 ;
        RECT -415.585 -70.475 -415.305 -70.195 ;
        RECT -415.585 -71.075 -415.305 -70.795 ;
        RECT -417.825 -73.835 -417.545 -73.555 ;
        RECT -417.825 -74.435 -417.545 -74.155 ;
        RECT -412.225 -67.115 -411.945 -66.835 ;
        RECT -412.225 -67.715 -411.945 -67.435 ;
        RECT -409.985 -67.115 -409.705 -66.835 ;
        RECT -409.985 -67.715 -409.705 -67.435 ;
        RECT -411.105 -70.475 -410.825 -70.195 ;
        RECT -411.105 -71.075 -410.825 -70.795 ;
        RECT -407.745 -67.115 -407.465 -66.835 ;
        RECT -407.745 -67.715 -407.465 -67.435 ;
        RECT -405.505 -67.115 -405.225 -66.835 ;
        RECT -405.505 -67.715 -405.225 -67.435 ;
        RECT -406.625 -70.475 -406.345 -70.195 ;
        RECT -406.625 -71.075 -406.345 -70.795 ;
        RECT -408.865 -73.835 -408.585 -73.555 ;
        RECT -408.865 -74.435 -408.585 -74.155 ;
        RECT -413.345 -77.195 -413.065 -76.915 ;
        RECT -413.345 -77.795 -413.065 -77.515 ;
        RECT -422.305 -80.555 -422.025 -80.275 ;
        RECT -422.305 -81.155 -422.025 -80.875 ;
        RECT -440.225 -83.915 -439.945 -83.635 ;
        RECT -440.225 -84.515 -439.945 -84.235 ;
        RECT -403.265 -67.115 -402.985 -66.835 ;
        RECT -403.265 -67.715 -402.985 -67.435 ;
        RECT -401.025 -67.115 -400.745 -66.835 ;
        RECT -401.025 -67.715 -400.745 -67.435 ;
        RECT -402.145 -70.475 -401.865 -70.195 ;
        RECT -402.145 -71.075 -401.865 -70.795 ;
        RECT -398.785 -67.115 -398.505 -66.835 ;
        RECT -398.785 -67.715 -398.505 -67.435 ;
        RECT -396.545 -67.115 -396.265 -66.835 ;
        RECT -396.545 -67.715 -396.265 -67.435 ;
        RECT -397.665 -70.475 -397.385 -70.195 ;
        RECT -397.665 -71.075 -397.385 -70.795 ;
        RECT -399.905 -73.835 -399.625 -73.555 ;
        RECT -399.905 -74.435 -399.625 -74.155 ;
        RECT -394.305 -67.115 -394.025 -66.835 ;
        RECT -394.305 -67.715 -394.025 -67.435 ;
        RECT -392.065 -67.115 -391.785 -66.835 ;
        RECT -392.065 -67.715 -391.785 -67.435 ;
        RECT -393.185 -70.475 -392.905 -70.195 ;
        RECT -393.185 -71.075 -392.905 -70.795 ;
        RECT -389.825 -67.115 -389.545 -66.835 ;
        RECT -389.825 -67.715 -389.545 -67.435 ;
        RECT -387.585 -67.115 -387.305 -66.835 ;
        RECT -387.585 -67.715 -387.305 -67.435 ;
        RECT -388.705 -70.475 -388.425 -70.195 ;
        RECT -388.705 -71.075 -388.425 -70.795 ;
        RECT -390.945 -73.835 -390.665 -73.555 ;
        RECT -390.945 -74.435 -390.665 -74.155 ;
        RECT -395.425 -77.195 -395.145 -76.915 ;
        RECT -395.425 -77.795 -395.145 -77.515 ;
        RECT -385.345 -67.115 -385.065 -66.835 ;
        RECT -385.345 -67.715 -385.065 -67.435 ;
        RECT -383.105 -67.115 -382.825 -66.835 ;
        RECT -383.105 -67.715 -382.825 -67.435 ;
        RECT -384.225 -70.475 -383.945 -70.195 ;
        RECT -384.225 -71.075 -383.945 -70.795 ;
        RECT -380.865 -67.115 -380.585 -66.835 ;
        RECT -380.865 -67.715 -380.585 -67.435 ;
        RECT -378.625 -67.115 -378.345 -66.835 ;
        RECT -378.625 -67.715 -378.345 -67.435 ;
        RECT -379.745 -70.475 -379.465 -70.195 ;
        RECT -379.745 -71.075 -379.465 -70.795 ;
        RECT -381.985 -73.835 -381.705 -73.555 ;
        RECT -381.985 -74.435 -381.705 -74.155 ;
        RECT -376.385 -67.115 -376.105 -66.835 ;
        RECT -376.385 -67.715 -376.105 -67.435 ;
        RECT -374.145 -67.115 -373.865 -66.835 ;
        RECT -374.145 -67.715 -373.865 -67.435 ;
        RECT -375.265 -70.475 -374.985 -70.195 ;
        RECT -375.265 -71.075 -374.985 -70.795 ;
        RECT -371.905 -67.115 -371.625 -66.835 ;
        RECT -371.905 -67.715 -371.625 -67.435 ;
        RECT -369.665 -67.115 -369.385 -66.835 ;
        RECT -369.665 -67.715 -369.385 -67.435 ;
        RECT -370.785 -70.475 -370.505 -70.195 ;
        RECT -370.785 -71.075 -370.505 -70.795 ;
        RECT -373.025 -73.835 -372.745 -73.555 ;
        RECT -373.025 -74.435 -372.745 -74.155 ;
        RECT -377.505 -77.195 -377.225 -76.915 ;
        RECT -377.505 -77.795 -377.225 -77.515 ;
        RECT -386.465 -80.555 -386.185 -80.275 ;
        RECT -386.465 -81.155 -386.185 -80.875 ;
        RECT -367.425 -67.115 -367.145 -66.835 ;
        RECT -367.425 -67.715 -367.145 -67.435 ;
        RECT -365.185 -67.115 -364.905 -66.835 ;
        RECT -365.185 -67.715 -364.905 -67.435 ;
        RECT -366.305 -70.475 -366.025 -70.195 ;
        RECT -366.305 -71.075 -366.025 -70.795 ;
        RECT -362.945 -67.115 -362.665 -66.835 ;
        RECT -362.945 -67.715 -362.665 -67.435 ;
        RECT -360.705 -67.115 -360.425 -66.835 ;
        RECT -360.705 -67.715 -360.425 -67.435 ;
        RECT -361.825 -70.475 -361.545 -70.195 ;
        RECT -361.825 -71.075 -361.545 -70.795 ;
        RECT -364.065 -73.835 -363.785 -73.555 ;
        RECT -364.065 -74.435 -363.785 -74.155 ;
        RECT -358.465 -67.115 -358.185 -66.835 ;
        RECT -358.465 -67.715 -358.185 -67.435 ;
        RECT -356.225 -67.115 -355.945 -66.835 ;
        RECT -356.225 -67.715 -355.945 -67.435 ;
        RECT -357.345 -70.475 -357.065 -70.195 ;
        RECT -357.345 -71.075 -357.065 -70.795 ;
        RECT -353.985 -67.115 -353.705 -66.835 ;
        RECT -353.985 -67.715 -353.705 -67.435 ;
        RECT -351.745 -67.115 -351.465 -66.835 ;
        RECT -351.745 -67.715 -351.465 -67.435 ;
        RECT -352.865 -70.475 -352.585 -70.195 ;
        RECT -352.865 -71.075 -352.585 -70.795 ;
        RECT -355.105 -73.835 -354.825 -73.555 ;
        RECT -355.105 -74.435 -354.825 -74.155 ;
        RECT -359.585 -77.195 -359.305 -76.915 ;
        RECT -359.585 -77.795 -359.305 -77.515 ;
        RECT -349.505 -67.115 -349.225 -66.835 ;
        RECT -349.505 -67.715 -349.225 -67.435 ;
        RECT -347.265 -67.115 -346.985 -66.835 ;
        RECT -347.265 -67.715 -346.985 -67.435 ;
        RECT -348.385 -70.475 -348.105 -70.195 ;
        RECT -348.385 -71.075 -348.105 -70.795 ;
        RECT -345.025 -67.115 -344.745 -66.835 ;
        RECT -345.025 -67.715 -344.745 -67.435 ;
        RECT -342.785 -67.115 -342.505 -66.835 ;
        RECT -342.785 -67.715 -342.505 -67.435 ;
        RECT -343.905 -70.475 -343.625 -70.195 ;
        RECT -343.905 -71.075 -343.625 -70.795 ;
        RECT -346.145 -73.835 -345.865 -73.555 ;
        RECT -346.145 -74.435 -345.865 -74.155 ;
        RECT -340.545 -67.115 -340.265 -66.835 ;
        RECT -340.545 -67.715 -340.265 -67.435 ;
        RECT -338.305 -67.115 -338.025 -66.835 ;
        RECT -338.305 -67.715 -338.025 -67.435 ;
        RECT -339.425 -70.475 -339.145 -70.195 ;
        RECT -339.425 -71.075 -339.145 -70.795 ;
        RECT -336.065 -67.115 -335.785 -66.835 ;
        RECT -336.065 -67.715 -335.785 -67.435 ;
        RECT -333.825 -67.115 -333.545 -66.835 ;
        RECT -333.825 -67.715 -333.545 -67.435 ;
        RECT -334.945 -70.475 -334.665 -70.195 ;
        RECT -334.945 -71.075 -334.665 -70.795 ;
        RECT -337.185 -73.835 -336.905 -73.555 ;
        RECT -337.185 -74.435 -336.905 -74.155 ;
        RECT -341.665 -77.195 -341.385 -76.915 ;
        RECT -341.665 -77.795 -341.385 -77.515 ;
        RECT -350.625 -80.555 -350.345 -80.275 ;
        RECT -350.625 -81.155 -350.345 -80.875 ;
        RECT -368.545 -83.915 -368.265 -83.635 ;
        RECT -368.545 -84.515 -368.265 -84.235 ;
        RECT -404.385 -87.275 -404.105 -86.995 ;
        RECT -404.385 -87.875 -404.105 -87.595 ;
        RECT -331.585 -67.115 -331.305 -66.835 ;
        RECT -331.585 -67.715 -331.305 -67.435 ;
        RECT -329.345 -67.115 -329.065 -66.835 ;
        RECT -329.345 -67.715 -329.065 -67.435 ;
        RECT -330.465 -70.475 -330.185 -70.195 ;
        RECT -330.465 -71.075 -330.185 -70.795 ;
        RECT -327.105 -67.115 -326.825 -66.835 ;
        RECT -327.105 -67.715 -326.825 -67.435 ;
        RECT -324.865 -67.115 -324.585 -66.835 ;
        RECT -324.865 -67.715 -324.585 -67.435 ;
        RECT -325.985 -70.475 -325.705 -70.195 ;
        RECT -325.985 -71.075 -325.705 -70.795 ;
        RECT -328.225 -73.835 -327.945 -73.555 ;
        RECT -328.225 -74.435 -327.945 -74.155 ;
        RECT -322.625 -67.115 -322.345 -66.835 ;
        RECT -322.625 -67.715 -322.345 -67.435 ;
        RECT -320.385 -67.115 -320.105 -66.835 ;
        RECT -320.385 -67.715 -320.105 -67.435 ;
        RECT -321.505 -70.475 -321.225 -70.195 ;
        RECT -321.505 -71.075 -321.225 -70.795 ;
        RECT -318.145 -67.115 -317.865 -66.835 ;
        RECT -318.145 -67.715 -317.865 -67.435 ;
        RECT -315.905 -67.115 -315.625 -66.835 ;
        RECT -315.905 -67.715 -315.625 -67.435 ;
        RECT -317.025 -70.475 -316.745 -70.195 ;
        RECT -317.025 -71.075 -316.745 -70.795 ;
        RECT -319.265 -73.835 -318.985 -73.555 ;
        RECT -319.265 -74.435 -318.985 -74.155 ;
        RECT -323.745 -77.195 -323.465 -76.915 ;
        RECT -323.745 -77.795 -323.465 -77.515 ;
        RECT -313.665 -67.115 -313.385 -66.835 ;
        RECT -313.665 -67.715 -313.385 -67.435 ;
        RECT -311.425 -67.115 -311.145 -66.835 ;
        RECT -311.425 -67.715 -311.145 -67.435 ;
        RECT -312.545 -70.475 -312.265 -70.195 ;
        RECT -312.545 -71.075 -312.265 -70.795 ;
        RECT -309.185 -67.115 -308.905 -66.835 ;
        RECT -309.185 -67.715 -308.905 -67.435 ;
        RECT -306.945 -67.115 -306.665 -66.835 ;
        RECT -306.945 -67.715 -306.665 -67.435 ;
        RECT -308.065 -70.475 -307.785 -70.195 ;
        RECT -308.065 -71.075 -307.785 -70.795 ;
        RECT -310.305 -73.835 -310.025 -73.555 ;
        RECT -310.305 -74.435 -310.025 -74.155 ;
        RECT -304.705 -67.115 -304.425 -66.835 ;
        RECT -304.705 -67.715 -304.425 -67.435 ;
        RECT -302.465 -67.115 -302.185 -66.835 ;
        RECT -302.465 -67.715 -302.185 -67.435 ;
        RECT -303.585 -70.475 -303.305 -70.195 ;
        RECT -303.585 -71.075 -303.305 -70.795 ;
        RECT -300.225 -67.115 -299.945 -66.835 ;
        RECT -300.225 -67.715 -299.945 -67.435 ;
        RECT -297.985 -67.115 -297.705 -66.835 ;
        RECT -297.985 -67.715 -297.705 -67.435 ;
        RECT -299.105 -70.475 -298.825 -70.195 ;
        RECT -299.105 -71.075 -298.825 -70.795 ;
        RECT -301.345 -73.835 -301.065 -73.555 ;
        RECT -301.345 -74.435 -301.065 -74.155 ;
        RECT -305.825 -77.195 -305.545 -76.915 ;
        RECT -305.825 -77.795 -305.545 -77.515 ;
        RECT -314.785 -80.555 -314.505 -80.275 ;
        RECT -314.785 -81.155 -314.505 -80.875 ;
        RECT -295.745 -67.115 -295.465 -66.835 ;
        RECT -295.745 -67.715 -295.465 -67.435 ;
        RECT -293.505 -67.115 -293.225 -66.835 ;
        RECT -293.505 -67.715 -293.225 -67.435 ;
        RECT -294.625 -70.475 -294.345 -70.195 ;
        RECT -294.625 -71.075 -294.345 -70.795 ;
        RECT -291.265 -67.115 -290.985 -66.835 ;
        RECT -291.265 -67.715 -290.985 -67.435 ;
        RECT -289.025 -67.115 -288.745 -66.835 ;
        RECT -289.025 -67.715 -288.745 -67.435 ;
        RECT -290.145 -70.475 -289.865 -70.195 ;
        RECT -290.145 -71.075 -289.865 -70.795 ;
        RECT -292.385 -73.835 -292.105 -73.555 ;
        RECT -292.385 -74.435 -292.105 -74.155 ;
        RECT -286.785 -67.115 -286.505 -66.835 ;
        RECT -286.785 -67.715 -286.505 -67.435 ;
        RECT -284.545 -67.115 -284.265 -66.835 ;
        RECT -284.545 -67.715 -284.265 -67.435 ;
        RECT -285.665 -70.475 -285.385 -70.195 ;
        RECT -285.665 -71.075 -285.385 -70.795 ;
        RECT -282.305 -67.115 -282.025 -66.835 ;
        RECT -282.305 -67.715 -282.025 -67.435 ;
        RECT -280.065 -67.115 -279.785 -66.835 ;
        RECT -280.065 -67.715 -279.785 -67.435 ;
        RECT -281.185 -70.475 -280.905 -70.195 ;
        RECT -281.185 -71.075 -280.905 -70.795 ;
        RECT -283.425 -73.835 -283.145 -73.555 ;
        RECT -283.425 -74.435 -283.145 -74.155 ;
        RECT -287.905 -77.195 -287.625 -76.915 ;
        RECT -287.905 -77.795 -287.625 -77.515 ;
        RECT -277.825 -67.115 -277.545 -66.835 ;
        RECT -277.825 -67.715 -277.545 -67.435 ;
        RECT -275.585 -67.115 -275.305 -66.835 ;
        RECT -275.585 -67.715 -275.305 -67.435 ;
        RECT -276.705 -70.475 -276.425 -70.195 ;
        RECT -276.705 -71.075 -276.425 -70.795 ;
        RECT -273.345 -67.115 -273.065 -66.835 ;
        RECT -273.345 -67.715 -273.065 -67.435 ;
        RECT -271.105 -67.115 -270.825 -66.835 ;
        RECT -271.105 -67.715 -270.825 -67.435 ;
        RECT -272.225 -70.475 -271.945 -70.195 ;
        RECT -272.225 -71.075 -271.945 -70.795 ;
        RECT -274.465 -73.835 -274.185 -73.555 ;
        RECT -274.465 -74.435 -274.185 -74.155 ;
        RECT -268.865 -67.115 -268.585 -66.835 ;
        RECT -268.865 -67.715 -268.585 -67.435 ;
        RECT -266.625 -67.115 -266.345 -66.835 ;
        RECT -266.625 -67.715 -266.345 -67.435 ;
        RECT -267.745 -70.475 -267.465 -70.195 ;
        RECT -267.745 -71.075 -267.465 -70.795 ;
        RECT -264.385 -67.115 -264.105 -66.835 ;
        RECT -264.385 -67.715 -264.105 -67.435 ;
        RECT -262.145 -67.115 -261.865 -66.835 ;
        RECT -262.145 -67.715 -261.865 -67.435 ;
        RECT -263.265 -70.475 -262.985 -70.195 ;
        RECT -263.265 -71.075 -262.985 -70.795 ;
        RECT -265.505 -73.835 -265.225 -73.555 ;
        RECT -265.505 -74.435 -265.225 -74.155 ;
        RECT -269.985 -77.195 -269.705 -76.915 ;
        RECT -269.985 -77.795 -269.705 -77.515 ;
        RECT -278.945 -80.555 -278.665 -80.275 ;
        RECT -278.945 -81.155 -278.665 -80.875 ;
        RECT -296.865 -83.915 -296.585 -83.635 ;
        RECT -296.865 -84.515 -296.585 -84.235 ;
        RECT -259.905 -67.115 -259.625 -66.835 ;
        RECT -259.905 -67.715 -259.625 -67.435 ;
        RECT -257.665 -67.115 -257.385 -66.835 ;
        RECT -257.665 -67.715 -257.385 -67.435 ;
        RECT -258.785 -70.475 -258.505 -70.195 ;
        RECT -258.785 -71.075 -258.505 -70.795 ;
        RECT -255.425 -67.115 -255.145 -66.835 ;
        RECT -255.425 -67.715 -255.145 -67.435 ;
        RECT -253.185 -67.115 -252.905 -66.835 ;
        RECT -253.185 -67.715 -252.905 -67.435 ;
        RECT -254.305 -70.475 -254.025 -70.195 ;
        RECT -254.305 -71.075 -254.025 -70.795 ;
        RECT -256.545 -73.835 -256.265 -73.555 ;
        RECT -256.545 -74.435 -256.265 -74.155 ;
        RECT -250.945 -67.115 -250.665 -66.835 ;
        RECT -250.945 -67.715 -250.665 -67.435 ;
        RECT -248.705 -67.115 -248.425 -66.835 ;
        RECT -248.705 -67.715 -248.425 -67.435 ;
        RECT -249.825 -70.475 -249.545 -70.195 ;
        RECT -249.825 -71.075 -249.545 -70.795 ;
        RECT -246.465 -67.115 -246.185 -66.835 ;
        RECT -246.465 -67.715 -246.185 -67.435 ;
        RECT -244.225 -67.115 -243.945 -66.835 ;
        RECT -244.225 -67.715 -243.945 -67.435 ;
        RECT -245.345 -70.475 -245.065 -70.195 ;
        RECT -245.345 -71.075 -245.065 -70.795 ;
        RECT -247.585 -73.835 -247.305 -73.555 ;
        RECT -247.585 -74.435 -247.305 -74.155 ;
        RECT -252.065 -77.195 -251.785 -76.915 ;
        RECT -252.065 -77.795 -251.785 -77.515 ;
        RECT -241.985 -67.115 -241.705 -66.835 ;
        RECT -241.985 -67.715 -241.705 -67.435 ;
        RECT -239.745 -67.115 -239.465 -66.835 ;
        RECT -239.745 -67.715 -239.465 -67.435 ;
        RECT -240.865 -70.475 -240.585 -70.195 ;
        RECT -240.865 -71.075 -240.585 -70.795 ;
        RECT -237.505 -67.115 -237.225 -66.835 ;
        RECT -237.505 -67.715 -237.225 -67.435 ;
        RECT -235.265 -67.115 -234.985 -66.835 ;
        RECT -235.265 -67.715 -234.985 -67.435 ;
        RECT -236.385 -70.475 -236.105 -70.195 ;
        RECT -236.385 -71.075 -236.105 -70.795 ;
        RECT -238.625 -73.835 -238.345 -73.555 ;
        RECT -238.625 -74.435 -238.345 -74.155 ;
        RECT -233.025 -67.115 -232.745 -66.835 ;
        RECT -233.025 -67.715 -232.745 -67.435 ;
        RECT -230.785 -67.115 -230.505 -66.835 ;
        RECT -230.785 -67.715 -230.505 -67.435 ;
        RECT -231.905 -70.475 -231.625 -70.195 ;
        RECT -231.905 -71.075 -231.625 -70.795 ;
        RECT -228.545 -67.115 -228.265 -66.835 ;
        RECT -228.545 -67.715 -228.265 -67.435 ;
        RECT -226.305 -67.115 -226.025 -66.835 ;
        RECT -226.305 -67.715 -226.025 -67.435 ;
        RECT -227.425 -70.475 -227.145 -70.195 ;
        RECT -227.425 -71.075 -227.145 -70.795 ;
        RECT -229.665 -73.835 -229.385 -73.555 ;
        RECT -229.665 -74.435 -229.385 -74.155 ;
        RECT -234.145 -77.195 -233.865 -76.915 ;
        RECT -234.145 -77.795 -233.865 -77.515 ;
        RECT -243.105 -80.555 -242.825 -80.275 ;
        RECT -243.105 -81.155 -242.825 -80.875 ;
        RECT -224.065 -67.115 -223.785 -66.835 ;
        RECT -224.065 -67.715 -223.785 -67.435 ;
        RECT -221.825 -67.115 -221.545 -66.835 ;
        RECT -221.825 -67.715 -221.545 -67.435 ;
        RECT -222.945 -70.475 -222.665 -70.195 ;
        RECT -222.945 -71.075 -222.665 -70.795 ;
        RECT -219.585 -67.115 -219.305 -66.835 ;
        RECT -219.585 -67.715 -219.305 -67.435 ;
        RECT -217.345 -67.115 -217.065 -66.835 ;
        RECT -217.345 -67.715 -217.065 -67.435 ;
        RECT -218.465 -70.475 -218.185 -70.195 ;
        RECT -218.465 -71.075 -218.185 -70.795 ;
        RECT -220.705 -73.835 -220.425 -73.555 ;
        RECT -220.705 -74.435 -220.425 -74.155 ;
        RECT -215.105 -67.115 -214.825 -66.835 ;
        RECT -215.105 -67.715 -214.825 -67.435 ;
        RECT -212.865 -67.115 -212.585 -66.835 ;
        RECT -212.865 -67.715 -212.585 -67.435 ;
        RECT -213.985 -70.475 -213.705 -70.195 ;
        RECT -213.985 -71.075 -213.705 -70.795 ;
        RECT -210.625 -67.115 -210.345 -66.835 ;
        RECT -210.625 -67.715 -210.345 -67.435 ;
        RECT -208.385 -67.115 -208.105 -66.835 ;
        RECT -208.385 -67.715 -208.105 -67.435 ;
        RECT -209.505 -70.475 -209.225 -70.195 ;
        RECT -209.505 -71.075 -209.225 -70.795 ;
        RECT -211.745 -73.835 -211.465 -73.555 ;
        RECT -211.745 -74.435 -211.465 -74.155 ;
        RECT -216.225 -77.195 -215.945 -76.915 ;
        RECT -216.225 -77.795 -215.945 -77.515 ;
        RECT -206.145 -67.115 -205.865 -66.835 ;
        RECT -206.145 -67.715 -205.865 -67.435 ;
        RECT -203.905 -67.115 -203.625 -66.835 ;
        RECT -203.905 -67.715 -203.625 -67.435 ;
        RECT -205.025 -70.475 -204.745 -70.195 ;
        RECT -205.025 -71.075 -204.745 -70.795 ;
        RECT -201.665 -67.115 -201.385 -66.835 ;
        RECT -201.665 -67.715 -201.385 -67.435 ;
        RECT -199.425 -67.115 -199.145 -66.835 ;
        RECT -199.425 -67.715 -199.145 -67.435 ;
        RECT -200.545 -70.475 -200.265 -70.195 ;
        RECT -200.545 -71.075 -200.265 -70.795 ;
        RECT -202.785 -73.835 -202.505 -73.555 ;
        RECT -202.785 -74.435 -202.505 -74.155 ;
        RECT -197.185 -67.115 -196.905 -66.835 ;
        RECT -197.185 -67.715 -196.905 -67.435 ;
        RECT -194.945 -67.115 -194.665 -66.835 ;
        RECT -194.945 -67.715 -194.665 -67.435 ;
        RECT -196.065 -70.475 -195.785 -70.195 ;
        RECT -196.065 -71.075 -195.785 -70.795 ;
        RECT -192.705 -67.115 -192.425 -66.835 ;
        RECT -192.705 -67.715 -192.425 -67.435 ;
        RECT -190.465 -67.115 -190.185 -66.835 ;
        RECT -190.465 -67.715 -190.185 -67.435 ;
        RECT -191.585 -70.475 -191.305 -70.195 ;
        RECT -191.585 -71.075 -191.305 -70.795 ;
        RECT -193.825 -73.835 -193.545 -73.555 ;
        RECT -193.825 -74.435 -193.545 -74.155 ;
        RECT -198.305 -77.195 -198.025 -76.915 ;
        RECT -198.305 -77.795 -198.025 -77.515 ;
        RECT -207.265 -80.555 -206.985 -80.275 ;
        RECT -207.265 -81.155 -206.985 -80.875 ;
        RECT -225.185 -83.915 -224.905 -83.635 ;
        RECT -225.185 -84.515 -224.905 -84.235 ;
        RECT -261.025 -87.275 -260.745 -86.995 ;
        RECT -261.025 -87.875 -260.745 -87.595 ;
        RECT -332.705 -90.635 -332.425 -90.355 ;
        RECT -332.705 -91.235 -332.425 -90.955 ;
        RECT -187.105 -67.115 -186.825 -66.835 ;
        RECT -187.105 -67.715 -186.825 -67.435 ;
        RECT -184.865 -67.115 -184.585 -66.835 ;
        RECT -184.865 -67.715 -184.585 -67.435 ;
        RECT -185.985 -70.475 -185.705 -70.195 ;
        RECT -185.985 -71.075 -185.705 -70.795 ;
        RECT -182.625 -67.115 -182.345 -66.835 ;
        RECT -182.625 -67.715 -182.345 -67.435 ;
        RECT -180.385 -67.115 -180.105 -66.835 ;
        RECT -180.385 -67.715 -180.105 -67.435 ;
        RECT -181.505 -70.475 -181.225 -70.195 ;
        RECT -181.505 -71.075 -181.225 -70.795 ;
        RECT -183.745 -73.835 -183.465 -73.555 ;
        RECT -183.745 -74.435 -183.465 -74.155 ;
        RECT -178.145 -67.115 -177.865 -66.835 ;
        RECT -178.145 -67.715 -177.865 -67.435 ;
        RECT -175.905 -67.115 -175.625 -66.835 ;
        RECT -175.905 -67.715 -175.625 -67.435 ;
        RECT -177.025 -70.475 -176.745 -70.195 ;
        RECT -177.025 -71.075 -176.745 -70.795 ;
        RECT -173.665 -67.115 -173.385 -66.835 ;
        RECT -173.665 -67.715 -173.385 -67.435 ;
        RECT -171.425 -67.115 -171.145 -66.835 ;
        RECT -171.425 -67.715 -171.145 -67.435 ;
        RECT -172.545 -70.475 -172.265 -70.195 ;
        RECT -172.545 -71.075 -172.265 -70.795 ;
        RECT -174.785 -73.835 -174.505 -73.555 ;
        RECT -174.785 -74.435 -174.505 -74.155 ;
        RECT -179.265 -77.195 -178.985 -76.915 ;
        RECT -179.265 -77.795 -178.985 -77.515 ;
        RECT -169.185 -67.115 -168.905 -66.835 ;
        RECT -169.185 -67.715 -168.905 -67.435 ;
        RECT -166.945 -67.115 -166.665 -66.835 ;
        RECT -166.945 -67.715 -166.665 -67.435 ;
        RECT -168.065 -70.475 -167.785 -70.195 ;
        RECT -168.065 -71.075 -167.785 -70.795 ;
        RECT -164.705 -67.115 -164.425 -66.835 ;
        RECT -164.705 -67.715 -164.425 -67.435 ;
        RECT -162.465 -67.115 -162.185 -66.835 ;
        RECT -162.465 -67.715 -162.185 -67.435 ;
        RECT -163.585 -70.475 -163.305 -70.195 ;
        RECT -163.585 -71.075 -163.305 -70.795 ;
        RECT -165.825 -73.835 -165.545 -73.555 ;
        RECT -165.825 -74.435 -165.545 -74.155 ;
        RECT -160.225 -67.115 -159.945 -66.835 ;
        RECT -160.225 -67.715 -159.945 -67.435 ;
        RECT -157.985 -67.115 -157.705 -66.835 ;
        RECT -157.985 -67.715 -157.705 -67.435 ;
        RECT -159.105 -70.475 -158.825 -70.195 ;
        RECT -159.105 -71.075 -158.825 -70.795 ;
        RECT -155.745 -67.115 -155.465 -66.835 ;
        RECT -155.745 -67.715 -155.465 -67.435 ;
        RECT -153.505 -67.115 -153.225 -66.835 ;
        RECT -153.505 -67.715 -153.225 -67.435 ;
        RECT -154.625 -70.475 -154.345 -70.195 ;
        RECT -154.625 -71.075 -154.345 -70.795 ;
        RECT -156.865 -73.835 -156.585 -73.555 ;
        RECT -156.865 -74.435 -156.585 -74.155 ;
        RECT -161.345 -77.195 -161.065 -76.915 ;
        RECT -161.345 -77.795 -161.065 -77.515 ;
        RECT -170.305 -80.555 -170.025 -80.275 ;
        RECT -170.305 -81.155 -170.025 -80.875 ;
        RECT -151.265 -67.115 -150.985 -66.835 ;
        RECT -151.265 -67.715 -150.985 -67.435 ;
        RECT -149.025 -67.115 -148.745 -66.835 ;
        RECT -149.025 -67.715 -148.745 -67.435 ;
        RECT -150.145 -70.475 -149.865 -70.195 ;
        RECT -150.145 -71.075 -149.865 -70.795 ;
        RECT -146.785 -67.115 -146.505 -66.835 ;
        RECT -146.785 -67.715 -146.505 -67.435 ;
        RECT -144.545 -67.115 -144.265 -66.835 ;
        RECT -144.545 -67.715 -144.265 -67.435 ;
        RECT -145.665 -70.475 -145.385 -70.195 ;
        RECT -145.665 -71.075 -145.385 -70.795 ;
        RECT -147.905 -73.835 -147.625 -73.555 ;
        RECT -147.905 -74.435 -147.625 -74.155 ;
        RECT -142.305 -67.115 -142.025 -66.835 ;
        RECT -142.305 -67.715 -142.025 -67.435 ;
        RECT -140.065 -67.115 -139.785 -66.835 ;
        RECT -140.065 -67.715 -139.785 -67.435 ;
        RECT -141.185 -70.475 -140.905 -70.195 ;
        RECT -141.185 -71.075 -140.905 -70.795 ;
        RECT -137.825 -67.115 -137.545 -66.835 ;
        RECT -137.825 -67.715 -137.545 -67.435 ;
        RECT -135.585 -67.115 -135.305 -66.835 ;
        RECT -135.585 -67.715 -135.305 -67.435 ;
        RECT -136.705 -70.475 -136.425 -70.195 ;
        RECT -136.705 -71.075 -136.425 -70.795 ;
        RECT -138.945 -73.835 -138.665 -73.555 ;
        RECT -138.945 -74.435 -138.665 -74.155 ;
        RECT -143.425 -77.195 -143.145 -76.915 ;
        RECT -143.425 -77.795 -143.145 -77.515 ;
        RECT -133.345 -67.115 -133.065 -66.835 ;
        RECT -133.345 -67.715 -133.065 -67.435 ;
        RECT -131.105 -67.115 -130.825 -66.835 ;
        RECT -131.105 -67.715 -130.825 -67.435 ;
        RECT -132.225 -70.475 -131.945 -70.195 ;
        RECT -132.225 -71.075 -131.945 -70.795 ;
        RECT -128.865 -67.115 -128.585 -66.835 ;
        RECT -128.865 -67.715 -128.585 -67.435 ;
        RECT -126.625 -67.115 -126.345 -66.835 ;
        RECT -126.625 -67.715 -126.345 -67.435 ;
        RECT -127.745 -70.475 -127.465 -70.195 ;
        RECT -127.745 -71.075 -127.465 -70.795 ;
        RECT -129.985 -73.835 -129.705 -73.555 ;
        RECT -129.985 -74.435 -129.705 -74.155 ;
        RECT -124.385 -67.115 -124.105 -66.835 ;
        RECT -124.385 -67.715 -124.105 -67.435 ;
        RECT -122.145 -67.115 -121.865 -66.835 ;
        RECT -122.145 -67.715 -121.865 -67.435 ;
        RECT -123.265 -70.475 -122.985 -70.195 ;
        RECT -123.265 -71.075 -122.985 -70.795 ;
        RECT -119.905 -67.115 -119.625 -66.835 ;
        RECT -119.905 -67.715 -119.625 -67.435 ;
        RECT -117.665 -67.115 -117.385 -66.835 ;
        RECT -117.665 -67.715 -117.385 -67.435 ;
        RECT -118.785 -70.475 -118.505 -70.195 ;
        RECT -118.785 -71.075 -118.505 -70.795 ;
        RECT -121.025 -73.835 -120.745 -73.555 ;
        RECT -121.025 -74.435 -120.745 -74.155 ;
        RECT -125.505 -77.195 -125.225 -76.915 ;
        RECT -125.505 -77.795 -125.225 -77.515 ;
        RECT -134.465 -80.555 -134.185 -80.275 ;
        RECT -134.465 -81.155 -134.185 -80.875 ;
        RECT -152.385 -83.915 -152.105 -83.635 ;
        RECT -152.385 -84.515 -152.105 -84.235 ;
        RECT -115.425 -67.115 -115.145 -66.835 ;
        RECT -115.425 -67.715 -115.145 -67.435 ;
        RECT -113.185 -67.115 -112.905 -66.835 ;
        RECT -113.185 -67.715 -112.905 -67.435 ;
        RECT -114.305 -70.475 -114.025 -70.195 ;
        RECT -114.305 -71.075 -114.025 -70.795 ;
        RECT -110.945 -67.115 -110.665 -66.835 ;
        RECT -110.945 -67.715 -110.665 -67.435 ;
        RECT -108.705 -67.115 -108.425 -66.835 ;
        RECT -108.705 -67.715 -108.425 -67.435 ;
        RECT -109.825 -70.475 -109.545 -70.195 ;
        RECT -109.825 -71.075 -109.545 -70.795 ;
        RECT -112.065 -73.835 -111.785 -73.555 ;
        RECT -112.065 -74.435 -111.785 -74.155 ;
        RECT -106.465 -67.115 -106.185 -66.835 ;
        RECT -106.465 -67.715 -106.185 -67.435 ;
        RECT -104.225 -67.115 -103.945 -66.835 ;
        RECT -104.225 -67.715 -103.945 -67.435 ;
        RECT -105.345 -70.475 -105.065 -70.195 ;
        RECT -105.345 -71.075 -105.065 -70.795 ;
        RECT -101.985 -67.115 -101.705 -66.835 ;
        RECT -101.985 -67.715 -101.705 -67.435 ;
        RECT -99.745 -67.115 -99.465 -66.835 ;
        RECT -99.745 -67.715 -99.465 -67.435 ;
        RECT -100.865 -70.475 -100.585 -70.195 ;
        RECT -100.865 -71.075 -100.585 -70.795 ;
        RECT -103.105 -73.835 -102.825 -73.555 ;
        RECT -103.105 -74.435 -102.825 -74.155 ;
        RECT -107.585 -77.195 -107.305 -76.915 ;
        RECT -107.585 -77.795 -107.305 -77.515 ;
        RECT -97.505 -67.115 -97.225 -66.835 ;
        RECT -97.505 -67.715 -97.225 -67.435 ;
        RECT -95.265 -67.115 -94.985 -66.835 ;
        RECT -95.265 -67.715 -94.985 -67.435 ;
        RECT -96.385 -70.475 -96.105 -70.195 ;
        RECT -96.385 -71.075 -96.105 -70.795 ;
        RECT -93.025 -67.115 -92.745 -66.835 ;
        RECT -93.025 -67.715 -92.745 -67.435 ;
        RECT -90.785 -67.115 -90.505 -66.835 ;
        RECT -90.785 -67.715 -90.505 -67.435 ;
        RECT -91.905 -70.475 -91.625 -70.195 ;
        RECT -91.905 -71.075 -91.625 -70.795 ;
        RECT -94.145 -73.835 -93.865 -73.555 ;
        RECT -94.145 -74.435 -93.865 -74.155 ;
        RECT -88.545 -67.115 -88.265 -66.835 ;
        RECT -88.545 -67.715 -88.265 -67.435 ;
        RECT -86.305 -67.115 -86.025 -66.835 ;
        RECT -86.305 -67.715 -86.025 -67.435 ;
        RECT -87.425 -70.475 -87.145 -70.195 ;
        RECT -87.425 -71.075 -87.145 -70.795 ;
        RECT -84.065 -67.115 -83.785 -66.835 ;
        RECT -84.065 -67.715 -83.785 -67.435 ;
        RECT -81.825 -67.115 -81.545 -66.835 ;
        RECT -81.825 -67.715 -81.545 -67.435 ;
        RECT -82.945 -70.475 -82.665 -70.195 ;
        RECT -82.945 -71.075 -82.665 -70.795 ;
        RECT -85.185 -73.835 -84.905 -73.555 ;
        RECT -85.185 -74.435 -84.905 -74.155 ;
        RECT -89.665 -77.195 -89.385 -76.915 ;
        RECT -89.665 -77.795 -89.385 -77.515 ;
        RECT -98.625 -80.555 -98.345 -80.275 ;
        RECT -98.625 -81.155 -98.345 -80.875 ;
        RECT -79.585 -67.115 -79.305 -66.835 ;
        RECT -79.585 -67.715 -79.305 -67.435 ;
        RECT -77.345 -67.115 -77.065 -66.835 ;
        RECT -77.345 -67.715 -77.065 -67.435 ;
        RECT -78.465 -70.475 -78.185 -70.195 ;
        RECT -78.465 -71.075 -78.185 -70.795 ;
        RECT -75.105 -67.115 -74.825 -66.835 ;
        RECT -75.105 -67.715 -74.825 -67.435 ;
        RECT -72.865 -67.115 -72.585 -66.835 ;
        RECT -72.865 -67.715 -72.585 -67.435 ;
        RECT -73.985 -70.475 -73.705 -70.195 ;
        RECT -73.985 -71.075 -73.705 -70.795 ;
        RECT -76.225 -73.835 -75.945 -73.555 ;
        RECT -76.225 -74.435 -75.945 -74.155 ;
        RECT -70.625 -67.115 -70.345 -66.835 ;
        RECT -70.625 -67.715 -70.345 -67.435 ;
        RECT -68.385 -67.115 -68.105 -66.835 ;
        RECT -68.385 -67.715 -68.105 -67.435 ;
        RECT -69.505 -70.475 -69.225 -70.195 ;
        RECT -69.505 -71.075 -69.225 -70.795 ;
        RECT -66.145 -67.115 -65.865 -66.835 ;
        RECT -66.145 -67.715 -65.865 -67.435 ;
        RECT -63.905 -67.115 -63.625 -66.835 ;
        RECT -63.905 -67.715 -63.625 -67.435 ;
        RECT -65.025 -70.475 -64.745 -70.195 ;
        RECT -65.025 -71.075 -64.745 -70.795 ;
        RECT -67.265 -73.835 -66.985 -73.555 ;
        RECT -67.265 -74.435 -66.985 -74.155 ;
        RECT -71.745 -77.195 -71.465 -76.915 ;
        RECT -71.745 -77.795 -71.465 -77.515 ;
        RECT -61.665 -67.115 -61.385 -66.835 ;
        RECT -61.665 -67.715 -61.385 -67.435 ;
        RECT -59.425 -67.115 -59.145 -66.835 ;
        RECT -59.425 -67.715 -59.145 -67.435 ;
        RECT -60.545 -70.475 -60.265 -70.195 ;
        RECT -60.545 -71.075 -60.265 -70.795 ;
        RECT -57.185 -67.115 -56.905 -66.835 ;
        RECT -57.185 -67.715 -56.905 -67.435 ;
        RECT -54.945 -67.115 -54.665 -66.835 ;
        RECT -54.945 -67.715 -54.665 -67.435 ;
        RECT -56.065 -70.475 -55.785 -70.195 ;
        RECT -56.065 -71.075 -55.785 -70.795 ;
        RECT -58.305 -73.835 -58.025 -73.555 ;
        RECT -58.305 -74.435 -58.025 -74.155 ;
        RECT -52.705 -67.115 -52.425 -66.835 ;
        RECT -52.705 -67.715 -52.425 -67.435 ;
        RECT -50.465 -67.115 -50.185 -66.835 ;
        RECT -50.465 -67.715 -50.185 -67.435 ;
        RECT -51.585 -70.475 -51.305 -70.195 ;
        RECT -51.585 -71.075 -51.305 -70.795 ;
        RECT -48.225 -67.115 -47.945 -66.835 ;
        RECT -48.225 -67.715 -47.945 -67.435 ;
        RECT -45.985 -67.115 -45.705 -66.835 ;
        RECT -45.985 -67.715 -45.705 -67.435 ;
        RECT -47.105 -70.475 -46.825 -70.195 ;
        RECT -47.105 -71.075 -46.825 -70.795 ;
        RECT -49.345 -73.835 -49.065 -73.555 ;
        RECT -49.345 -74.435 -49.065 -74.155 ;
        RECT -53.825 -77.195 -53.545 -76.915 ;
        RECT -53.825 -77.795 -53.545 -77.515 ;
        RECT -62.785 -80.555 -62.505 -80.275 ;
        RECT -62.785 -81.155 -62.505 -80.875 ;
        RECT -80.705 -83.915 -80.425 -83.635 ;
        RECT -80.705 -84.515 -80.425 -84.235 ;
        RECT -116.545 -87.275 -116.265 -86.995 ;
        RECT -116.545 -87.875 -116.265 -87.595 ;
        RECT -43.745 -67.115 -43.465 -66.835 ;
        RECT -43.745 -67.715 -43.465 -67.435 ;
        RECT -41.505 -67.115 -41.225 -66.835 ;
        RECT -41.505 -67.715 -41.225 -67.435 ;
        RECT -42.625 -70.475 -42.345 -70.195 ;
        RECT -42.625 -71.075 -42.345 -70.795 ;
        RECT -39.265 -67.115 -38.985 -66.835 ;
        RECT -39.265 -67.715 -38.985 -67.435 ;
        RECT -37.025 -67.115 -36.745 -66.835 ;
        RECT -37.025 -67.715 -36.745 -67.435 ;
        RECT -38.145 -70.475 -37.865 -70.195 ;
        RECT -38.145 -71.075 -37.865 -70.795 ;
        RECT -40.385 -73.835 -40.105 -73.555 ;
        RECT -40.385 -74.435 -40.105 -74.155 ;
        RECT -34.785 -67.115 -34.505 -66.835 ;
        RECT -34.785 -67.715 -34.505 -67.435 ;
        RECT -32.545 -67.115 -32.265 -66.835 ;
        RECT -32.545 -67.715 -32.265 -67.435 ;
        RECT -33.665 -70.475 -33.385 -70.195 ;
        RECT -33.665 -71.075 -33.385 -70.795 ;
        RECT -30.305 -67.115 -30.025 -66.835 ;
        RECT -30.305 -67.715 -30.025 -67.435 ;
        RECT -28.065 -67.115 -27.785 -66.835 ;
        RECT -28.065 -67.715 -27.785 -67.435 ;
        RECT -29.185 -70.475 -28.905 -70.195 ;
        RECT -29.185 -71.075 -28.905 -70.795 ;
        RECT -31.425 -73.835 -31.145 -73.555 ;
        RECT -31.425 -74.435 -31.145 -74.155 ;
        RECT -35.905 -77.195 -35.625 -76.915 ;
        RECT -35.905 -77.795 -35.625 -77.515 ;
        RECT -25.825 -67.115 -25.545 -66.835 ;
        RECT -25.825 -67.715 -25.545 -67.435 ;
        RECT -23.585 -67.115 -23.305 -66.835 ;
        RECT -23.585 -67.715 -23.305 -67.435 ;
        RECT -24.705 -70.475 -24.425 -70.195 ;
        RECT -24.705 -71.075 -24.425 -70.795 ;
        RECT -21.345 -67.115 -21.065 -66.835 ;
        RECT -21.345 -67.715 -21.065 -67.435 ;
        RECT -19.105 -67.115 -18.825 -66.835 ;
        RECT -19.105 -67.715 -18.825 -67.435 ;
        RECT -20.225 -70.475 -19.945 -70.195 ;
        RECT -20.225 -71.075 -19.945 -70.795 ;
        RECT -22.465 -73.835 -22.185 -73.555 ;
        RECT -22.465 -74.435 -22.185 -74.155 ;
        RECT -16.865 -67.115 -16.585 -66.835 ;
        RECT -16.865 -67.715 -16.585 -67.435 ;
        RECT -14.625 -67.115 -14.345 -66.835 ;
        RECT -14.625 -67.715 -14.345 -67.435 ;
        RECT -15.745 -70.475 -15.465 -70.195 ;
        RECT -15.745 -71.075 -15.465 -70.795 ;
        RECT -12.385 -67.115 -12.105 -66.835 ;
        RECT -12.385 -67.715 -12.105 -67.435 ;
        RECT -10.145 -67.115 -9.865 -66.835 ;
        RECT -10.145 -67.715 -9.865 -67.435 ;
        RECT -11.265 -70.475 -10.985 -70.195 ;
        RECT -11.265 -71.075 -10.985 -70.795 ;
        RECT -13.505 -73.835 -13.225 -73.555 ;
        RECT -13.505 -74.435 -13.225 -74.155 ;
        RECT -17.985 -77.195 -17.705 -76.915 ;
        RECT -17.985 -77.795 -17.705 -77.515 ;
        RECT -26.945 -80.555 -26.665 -80.275 ;
        RECT -26.945 -81.155 -26.665 -80.875 ;
        RECT -7.905 -67.115 -7.625 -66.835 ;
        RECT -7.905 -67.715 -7.625 -67.435 ;
        RECT -5.665 -67.115 -5.385 -66.835 ;
        RECT -5.665 -67.715 -5.385 -67.435 ;
        RECT -6.785 -70.475 -6.505 -70.195 ;
        RECT -6.785 -71.075 -6.505 -70.795 ;
        RECT -3.425 -67.115 -3.145 -66.835 ;
        RECT -3.425 -67.715 -3.145 -67.435 ;
        RECT -1.185 -67.115 -0.905 -66.835 ;
        RECT -1.185 -67.715 -0.905 -67.435 ;
        RECT -2.305 -70.475 -2.025 -70.195 ;
        RECT -2.305 -71.075 -2.025 -70.795 ;
        RECT -4.545 -73.835 -4.265 -73.555 ;
        RECT -4.545 -74.435 -4.265 -74.155 ;
        RECT 1.055 -67.115 1.335 -66.835 ;
        RECT 1.055 -67.715 1.335 -67.435 ;
        RECT 3.295 -67.115 3.575 -66.835 ;
        RECT 3.295 -67.715 3.575 -67.435 ;
        RECT 2.175 -70.475 2.455 -70.195 ;
        RECT 2.175 -71.075 2.455 -70.795 ;
        RECT 5.535 -67.115 5.815 -66.835 ;
        RECT 5.535 -67.715 5.815 -67.435 ;
        RECT 7.775 -67.115 8.055 -66.835 ;
        RECT 7.775 -67.715 8.055 -67.435 ;
        RECT 6.655 -70.475 6.935 -70.195 ;
        RECT 6.655 -71.075 6.935 -70.795 ;
        RECT 4.415 -73.835 4.695 -73.555 ;
        RECT 4.415 -74.435 4.695 -74.155 ;
        RECT -0.065 -77.195 0.215 -76.915 ;
        RECT -0.065 -77.795 0.215 -77.515 ;
        RECT 10.015 -67.115 10.295 -66.835 ;
        RECT 10.015 -67.715 10.295 -67.435 ;
        RECT 12.255 -67.115 12.535 -66.835 ;
        RECT 12.255 -67.715 12.535 -67.435 ;
        RECT 11.135 -70.475 11.415 -70.195 ;
        RECT 11.135 -71.075 11.415 -70.795 ;
        RECT 14.495 -67.115 14.775 -66.835 ;
        RECT 14.495 -67.715 14.775 -67.435 ;
        RECT 16.735 -67.115 17.015 -66.835 ;
        RECT 16.735 -67.715 17.015 -67.435 ;
        RECT 15.615 -70.475 15.895 -70.195 ;
        RECT 15.615 -71.075 15.895 -70.795 ;
        RECT 13.375 -73.835 13.655 -73.555 ;
        RECT 13.375 -74.435 13.655 -74.155 ;
        RECT 18.975 -67.115 19.255 -66.835 ;
        RECT 18.975 -67.715 19.255 -67.435 ;
        RECT 21.215 -67.115 21.495 -66.835 ;
        RECT 21.215 -67.715 21.495 -67.435 ;
        RECT 20.095 -70.475 20.375 -70.195 ;
        RECT 20.095 -71.075 20.375 -70.795 ;
        RECT 23.455 -67.115 23.735 -66.835 ;
        RECT 23.455 -67.715 23.735 -67.435 ;
        RECT 25.695 -67.115 25.975 -66.835 ;
        RECT 25.695 -67.715 25.975 -67.435 ;
        RECT 24.575 -70.475 24.855 -70.195 ;
        RECT 24.575 -71.075 24.855 -70.795 ;
        RECT 22.335 -73.835 22.615 -73.555 ;
        RECT 22.335 -74.435 22.615 -74.155 ;
        RECT 17.855 -77.195 18.135 -76.915 ;
        RECT 17.855 -77.795 18.135 -77.515 ;
        RECT 8.895 -80.555 9.175 -80.275 ;
        RECT 8.895 -81.155 9.175 -80.875 ;
        RECT -9.025 -83.915 -8.745 -83.635 ;
        RECT -9.025 -84.515 -8.745 -84.235 ;
        RECT 27.935 -67.115 28.215 -66.835 ;
        RECT 27.935 -67.715 28.215 -67.435 ;
        RECT 30.175 -67.115 30.455 -66.835 ;
        RECT 30.175 -67.715 30.455 -67.435 ;
        RECT 29.055 -70.475 29.335 -70.195 ;
        RECT 29.055 -71.075 29.335 -70.795 ;
        RECT 32.415 -67.115 32.695 -66.835 ;
        RECT 32.415 -67.715 32.695 -67.435 ;
        RECT 34.655 -67.115 34.935 -66.835 ;
        RECT 34.655 -67.715 34.935 -67.435 ;
        RECT 33.535 -70.475 33.815 -70.195 ;
        RECT 33.535 -71.075 33.815 -70.795 ;
        RECT 31.295 -73.835 31.575 -73.555 ;
        RECT 31.295 -74.435 31.575 -74.155 ;
        RECT 36.895 -67.115 37.175 -66.835 ;
        RECT 36.895 -67.715 37.175 -67.435 ;
        RECT 39.135 -67.115 39.415 -66.835 ;
        RECT 39.135 -67.715 39.415 -67.435 ;
        RECT 38.015 -70.475 38.295 -70.195 ;
        RECT 38.015 -71.075 38.295 -70.795 ;
        RECT 41.375 -67.115 41.655 -66.835 ;
        RECT 41.375 -67.715 41.655 -67.435 ;
        RECT 43.615 -67.115 43.895 -66.835 ;
        RECT 43.615 -67.715 43.895 -67.435 ;
        RECT 42.495 -70.475 42.775 -70.195 ;
        RECT 42.495 -71.075 42.775 -70.795 ;
        RECT 40.255 -73.835 40.535 -73.555 ;
        RECT 40.255 -74.435 40.535 -74.155 ;
        RECT 35.775 -77.195 36.055 -76.915 ;
        RECT 35.775 -77.795 36.055 -77.515 ;
        RECT 45.855 -67.115 46.135 -66.835 ;
        RECT 45.855 -67.715 46.135 -67.435 ;
        RECT 48.095 -67.115 48.375 -66.835 ;
        RECT 48.095 -67.715 48.375 -67.435 ;
        RECT 46.975 -70.475 47.255 -70.195 ;
        RECT 46.975 -71.075 47.255 -70.795 ;
        RECT 50.335 -67.115 50.615 -66.835 ;
        RECT 50.335 -67.715 50.615 -67.435 ;
        RECT 52.575 -67.115 52.855 -66.835 ;
        RECT 52.575 -67.715 52.855 -67.435 ;
        RECT 51.455 -70.475 51.735 -70.195 ;
        RECT 51.455 -71.075 51.735 -70.795 ;
        RECT 49.215 -73.835 49.495 -73.555 ;
        RECT 49.215 -74.435 49.495 -74.155 ;
        RECT 54.815 -67.115 55.095 -66.835 ;
        RECT 54.815 -67.715 55.095 -67.435 ;
        RECT 57.055 -67.115 57.335 -66.835 ;
        RECT 57.055 -67.715 57.335 -67.435 ;
        RECT 55.935 -70.475 56.215 -70.195 ;
        RECT 55.935 -71.075 56.215 -70.795 ;
        RECT 59.295 -67.115 59.575 -66.835 ;
        RECT 59.295 -67.715 59.575 -67.435 ;
        RECT 61.535 -67.115 61.815 -66.835 ;
        RECT 61.535 -67.715 61.815 -67.435 ;
        RECT 60.415 -70.475 60.695 -70.195 ;
        RECT 60.415 -71.075 60.695 -70.795 ;
        RECT 58.175 -73.835 58.455 -73.555 ;
        RECT 58.175 -74.435 58.455 -74.155 ;
        RECT 53.695 -77.195 53.975 -76.915 ;
        RECT 53.695 -77.795 53.975 -77.515 ;
        RECT 44.735 -80.555 45.015 -80.275 ;
        RECT 44.735 -81.155 45.015 -80.875 ;
        RECT 63.775 -67.115 64.055 -66.835 ;
        RECT 63.775 -67.715 64.055 -67.435 ;
        RECT 66.015 -67.115 66.295 -66.835 ;
        RECT 66.015 -67.715 66.295 -67.435 ;
        RECT 64.895 -70.475 65.175 -70.195 ;
        RECT 64.895 -71.075 65.175 -70.795 ;
        RECT 68.255 -67.115 68.535 -66.835 ;
        RECT 68.255 -67.715 68.535 -67.435 ;
        RECT 70.495 -67.115 70.775 -66.835 ;
        RECT 70.495 -67.715 70.775 -67.435 ;
        RECT 69.375 -70.475 69.655 -70.195 ;
        RECT 69.375 -71.075 69.655 -70.795 ;
        RECT 67.135 -73.835 67.415 -73.555 ;
        RECT 67.135 -74.435 67.415 -74.155 ;
        RECT 72.735 -67.115 73.015 -66.835 ;
        RECT 72.735 -67.715 73.015 -67.435 ;
        RECT 74.975 -67.115 75.255 -66.835 ;
        RECT 74.975 -67.715 75.255 -67.435 ;
        RECT 73.855 -70.475 74.135 -70.195 ;
        RECT 73.855 -71.075 74.135 -70.795 ;
        RECT 77.215 -67.115 77.495 -66.835 ;
        RECT 77.215 -67.715 77.495 -67.435 ;
        RECT 79.455 -67.115 79.735 -66.835 ;
        RECT 79.455 -67.715 79.735 -67.435 ;
        RECT 78.335 -70.475 78.615 -70.195 ;
        RECT 78.335 -71.075 78.615 -70.795 ;
        RECT 76.095 -73.835 76.375 -73.555 ;
        RECT 76.095 -74.435 76.375 -74.155 ;
        RECT 71.615 -77.195 71.895 -76.915 ;
        RECT 71.615 -77.795 71.895 -77.515 ;
        RECT 81.695 -67.115 81.975 -66.835 ;
        RECT 81.695 -67.715 81.975 -67.435 ;
        RECT 83.935 -67.115 84.215 -66.835 ;
        RECT 83.935 -67.715 84.215 -67.435 ;
        RECT 82.815 -70.475 83.095 -70.195 ;
        RECT 82.815 -71.075 83.095 -70.795 ;
        RECT 86.175 -67.115 86.455 -66.835 ;
        RECT 86.175 -67.715 86.455 -67.435 ;
        RECT 88.415 -67.115 88.695 -66.835 ;
        RECT 88.415 -67.715 88.695 -67.435 ;
        RECT 87.295 -70.475 87.575 -70.195 ;
        RECT 87.295 -71.075 87.575 -70.795 ;
        RECT 85.055 -73.835 85.335 -73.555 ;
        RECT 85.055 -74.435 85.335 -74.155 ;
        RECT 90.655 -67.115 90.935 -66.835 ;
        RECT 90.655 -67.715 90.935 -67.435 ;
        RECT 92.895 -67.115 93.175 -66.835 ;
        RECT 92.895 -67.715 93.175 -67.435 ;
        RECT 91.775 -70.475 92.055 -70.195 ;
        RECT 91.775 -71.075 92.055 -70.795 ;
        RECT 95.135 -67.115 95.415 -66.835 ;
        RECT 95.135 -67.715 95.415 -67.435 ;
        RECT 287.250 -56.180 287.530 -55.900 ;
        RECT 287.810 -56.180 288.090 -55.900 ;
        RECT 288.370 -56.180 288.650 -55.900 ;
        RECT 312.300 2.900 312.580 3.180 ;
        RECT 311.740 -4.380 312.020 -4.100 ;
        RECT 312.860 -15.580 313.140 -15.300 ;
        RECT 312.300 -23.980 312.580 -23.700 ;
        RECT 313.980 19.140 314.260 19.420 ;
        RECT 313.980 5.140 314.260 5.420 ;
        RECT 313.420 -20.620 313.700 -20.340 ;
        RECT 313.980 -25.100 314.260 -24.820 ;
        RECT 312.860 -29.020 313.140 -28.740 ;
        RECT 317.900 26.980 318.180 27.260 ;
        RECT 334.140 43.780 334.420 44.060 ;
        RECT 344.220 43.780 344.500 44.060 ;
        RECT 353.740 43.780 354.020 44.060 ;
        RECT 405.820 45.460 406.100 45.740 ;
        RECT 408.060 45.460 408.340 45.740 ;
        RECT 376.140 43.780 376.420 44.060 ;
        RECT 319.580 42.100 319.860 42.380 ;
        RECT 321.820 35.380 322.100 35.660 ;
        RECT 316.780 18.020 317.060 18.300 ;
        RECT 318.460 11.300 318.740 11.580 ;
        RECT 316.780 6.260 317.060 6.540 ;
        RECT 331.340 26.420 331.620 26.700 ;
        RECT 321.820 24.180 322.100 24.460 ;
        RECT 333.020 28.100 333.300 28.380 ;
        RECT 332.460 19.700 332.740 19.980 ;
        RECT 320.700 14.100 320.980 14.380 ;
        RECT 321.260 11.300 321.540 11.580 ;
        RECT 319.580 7.380 319.860 7.660 ;
        RECT 321.820 6.820 322.100 7.100 ;
        RECT 324.060 19.140 324.340 19.420 ;
        RECT 329.100 18.020 329.380 18.300 ;
        RECT 325.180 15.220 325.460 15.500 ;
        RECT 326.860 14.660 327.140 14.940 ;
        RECT 325.180 14.100 325.460 14.380 ;
        RECT 325.740 12.420 326.020 12.700 ;
        RECT 324.620 11.860 324.900 12.140 ;
        RECT 327.420 11.860 327.700 12.140 ;
        RECT 325.740 11.300 326.020 11.580 ;
        RECT 322.380 7.940 322.660 8.220 ;
        RECT 321.820 4.580 322.100 4.860 ;
        RECT 326.300 4.580 326.580 4.860 ;
        RECT 327.420 6.260 327.700 6.540 ;
        RECT 326.860 5.140 327.140 5.420 ;
        RECT 329.660 7.940 329.940 8.220 ;
        RECT 316.220 -1.020 316.500 -0.740 ;
        RECT 318.460 -1.020 318.740 -0.740 ;
        RECT 319.580 -0.460 319.860 -0.180 ;
        RECT 319.020 -3.820 319.300 -3.540 ;
        RECT 320.700 -2.140 320.980 -1.860 ;
        RECT 323.500 -2.140 323.780 -1.860 ;
        RECT 320.140 -3.260 320.420 -2.980 ;
        RECT 321.820 -3.820 322.100 -3.540 ;
        RECT 331.900 4.580 332.180 4.860 ;
        RECT 330.780 3.460 331.060 3.740 ;
        RECT 331.340 -1.580 331.620 -1.300 ;
        RECT 325.740 -3.260 326.020 -2.980 ;
        RECT 328.540 -3.260 328.820 -2.980 ;
        RECT 323.500 -4.940 323.780 -4.660 ;
        RECT 326.300 -4.940 326.580 -4.660 ;
        RECT 330.780 -4.940 331.060 -4.660 ;
        RECT 330.780 -15.580 331.060 -15.300 ;
        RECT 321.820 -16.140 322.100 -15.860 ;
        RECT 321.820 -17.260 322.100 -16.980 ;
        RECT 319.020 -18.940 319.300 -18.660 ;
        RECT 321.820 -19.500 322.100 -19.220 ;
        RECT 319.580 -23.420 319.860 -23.140 ;
        RECT 319.020 -27.340 319.300 -27.060 ;
        RECT 318.460 -27.900 318.740 -27.620 ;
        RECT 310.060 -39.100 310.340 -38.820 ;
        RECT 314.540 -30.140 314.820 -29.860 ;
        RECT 317.340 -30.700 317.620 -30.420 ;
        RECT 315.100 -32.940 315.380 -32.660 ;
        RECT 317.900 -34.620 318.180 -34.340 ;
        RECT 312.860 -39.100 313.140 -38.820 ;
        RECT 317.340 -39.660 317.620 -39.380 ;
        RECT 315.100 -44.140 315.380 -43.860 ;
        RECT 322.380 -25.100 322.660 -24.820 ;
        RECT 329.100 -16.140 329.380 -15.860 ;
        RECT 325.180 -19.500 325.460 -19.220 ;
        RECT 324.620 -20.620 324.900 -20.340 ;
        RECT 327.980 -20.620 328.260 -20.340 ;
        RECT 325.180 -27.340 325.460 -27.060 ;
        RECT 324.060 -27.900 324.340 -27.620 ;
        RECT 320.700 -31.260 320.980 -30.980 ;
        RECT 321.260 -34.620 321.540 -34.340 ;
        RECT 327.980 -31.820 328.260 -31.540 ;
        RECT 326.300 -32.380 326.580 -32.100 ;
        RECT 323.500 -35.180 323.780 -34.900 ;
        RECT 319.020 -36.860 319.300 -36.580 ;
        RECT 321.820 -35.740 322.100 -35.460 ;
        RECT 325.180 -36.300 325.460 -36.020 ;
        RECT 322.940 -39.100 323.220 -38.820 ;
        RECT 330.780 -20.060 331.060 -19.780 ;
        RECT 331.340 -28.460 331.620 -28.180 ;
        RECT 329.100 -32.380 329.380 -32.100 ;
        RECT 330.780 -31.820 331.060 -31.540 ;
        RECT 326.300 -39.660 326.580 -39.380 ;
        RECT 327.980 -38.540 328.260 -38.260 ;
        RECT 331.900 -32.380 332.180 -32.100 ;
        RECT 333.020 -36.300 333.300 -36.020 ;
        RECT 331.900 -40.220 332.180 -39.940 ;
        RECT 338.060 39.300 338.340 39.580 ;
        RECT 339.180 39.860 339.460 40.140 ;
        RECT 339.180 38.740 339.460 39.020 ;
        RECT 338.060 35.380 338.340 35.660 ;
        RECT 341.420 34.820 341.700 35.100 ;
        RECT 335.260 30.340 335.540 30.620 ;
        RECT 335.260 28.660 335.540 28.940 ;
        RECT 336.380 30.340 336.660 30.620 ;
        RECT 337.500 28.100 337.780 28.380 ;
        RECT 334.700 26.980 334.980 27.260 ;
        RECT 334.140 24.180 334.420 24.460 ;
        RECT 334.140 22.500 334.420 22.780 ;
        RECT 337.500 22.500 337.780 22.780 ;
        RECT 341.980 35.380 342.260 35.660 ;
        RECT 343.660 34.820 343.940 35.100 ;
        RECT 345.340 34.820 345.620 35.100 ;
        RECT 349.260 34.820 349.540 35.100 ;
        RECT 343.660 32.020 343.940 32.300 ;
        RECT 349.820 34.260 350.100 34.540 ;
        RECT 343.660 28.100 343.940 28.380 ;
        RECT 344.220 23.060 344.500 23.340 ;
        RECT 339.740 22.500 340.020 22.780 ;
        RECT 342.540 19.700 342.820 19.980 ;
        RECT 343.100 15.220 343.380 15.500 ;
        RECT 343.100 14.100 343.380 14.380 ;
        RECT 341.420 7.940 341.700 8.220 ;
        RECT 339.180 6.260 339.460 6.540 ;
        RECT 347.580 26.980 347.860 27.260 ;
        RECT 348.140 23.060 348.420 23.340 ;
        RECT 346.460 22.500 346.740 22.780 ;
        RECT 346.460 20.260 346.740 20.540 ;
        RECT 344.780 11.860 345.060 12.140 ;
        RECT 345.340 14.660 345.620 14.940 ;
        RECT 344.780 7.940 345.060 8.220 ;
        RECT 350.940 20.260 351.220 20.540 ;
        RECT 346.460 11.300 346.740 11.580 ;
        RECT 339.180 -3.260 339.460 -2.980 ;
        RECT 335.260 -4.380 335.540 -4.100 ;
        RECT 336.940 -4.380 337.220 -4.100 ;
        RECT 335.260 -23.420 335.540 -23.140 ;
        RECT 346.460 2.900 346.740 3.180 ;
        RECT 350.940 2.900 351.220 3.180 ;
        RECT 351.500 0.100 351.780 0.380 ;
        RECT 346.460 -3.820 346.740 -3.540 ;
        RECT 345.340 -7.740 345.620 -7.460 ;
        RECT 347.020 -4.380 347.300 -4.100 ;
        RECT 345.900 -8.860 346.180 -8.580 ;
        RECT 349.260 -4.940 349.540 -4.660 ;
        RECT 350.380 -1.580 350.660 -1.300 ;
        RECT 350.940 -4.380 351.220 -4.100 ;
        RECT 349.820 -6.620 350.100 -6.340 ;
        RECT 338.620 -34.060 338.900 -33.780 ;
        RECT 336.940 -36.860 337.220 -36.580 ;
        RECT 342.540 -32.940 342.820 -32.660 ;
        RECT 345.340 -25.100 345.620 -24.820 ;
        RECT 346.460 -27.340 346.740 -27.060 ;
        RECT 344.780 -32.940 345.060 -32.660 ;
        RECT 342.540 -35.180 342.820 -34.900 ;
        RECT 338.620 -42.460 338.900 -42.180 ;
        RECT 339.180 -40.780 339.460 -40.500 ;
        RECT 334.700 -43.580 334.980 -43.300 ;
        RECT 339.740 -41.900 340.020 -41.620 ;
        RECT 360.460 38.740 360.740 39.020 ;
        RECT 363.260 38.740 363.540 39.020 ;
        RECT 361.580 38.180 361.860 38.460 ;
        RECT 365.500 38.740 365.780 39.020 ;
        RECT 364.940 38.180 365.220 38.460 ;
        RECT 355.420 35.380 355.700 35.660 ;
        RECT 356.540 35.380 356.820 35.660 ;
        RECT 360.460 34.820 360.740 35.100 ;
        RECT 360.460 30.900 360.740 31.180 ;
        RECT 357.660 26.980 357.940 27.260 ;
        RECT 361.580 26.980 361.860 27.260 ;
        RECT 364.380 34.820 364.660 35.100 ;
        RECT 363.260 34.260 363.540 34.540 ;
        RECT 363.260 30.900 363.540 31.180 ;
        RECT 373.900 41.540 374.180 41.820 ;
        RECT 378.940 41.540 379.220 41.820 ;
        RECT 377.820 39.860 378.100 40.140 ;
        RECT 373.900 38.740 374.180 39.020 ;
        RECT 385.660 41.540 385.940 41.820 ;
        RECT 386.220 38.180 386.500 38.460 ;
        RECT 369.980 35.380 370.260 35.660 ;
        RECT 377.820 35.380 378.100 35.660 ;
        RECT 366.060 34.820 366.340 35.100 ;
        RECT 364.940 30.900 365.220 31.180 ;
        RECT 362.140 21.940 362.420 22.220 ;
        RECT 369.980 29.780 370.260 30.060 ;
        RECT 381.740 30.340 382.020 30.620 ;
        RECT 357.100 14.100 357.380 14.380 ;
        RECT 359.340 10.740 359.620 11.020 ;
        RECT 355.980 10.180 356.260 10.460 ;
        RECT 356.540 0.660 356.820 0.940 ;
        RECT 358.780 -1.580 359.060 -1.300 ;
        RECT 367.180 19.140 367.460 19.420 ;
        RECT 369.420 18.580 369.700 18.860 ;
        RECT 363.260 10.740 363.540 11.020 ;
        RECT 363.820 15.220 364.100 15.500 ;
        RECT 363.820 0.100 364.100 0.380 ;
        RECT 369.980 10.180 370.260 10.460 ;
        RECT 364.380 -0.460 364.660 -0.180 ;
        RECT 363.260 -1.020 363.540 -0.740 ;
        RECT 362.700 -1.580 362.980 -1.300 ;
        RECT 356.540 -4.940 356.820 -4.660 ;
        RECT 353.740 -6.620 354.020 -6.340 ;
        RECT 353.740 -11.660 354.020 -11.380 ;
        RECT 360.460 -5.500 360.740 -5.220 ;
        RECT 361.580 -6.060 361.860 -5.780 ;
        RECT 361.020 -8.860 361.300 -8.580 ;
        RECT 364.380 -5.500 364.660 -5.220 ;
        RECT 367.180 2.340 367.460 2.620 ;
        RECT 363.820 -6.060 364.100 -5.780 ;
        RECT 362.140 -8.860 362.420 -8.580 ;
        RECT 363.260 -8.860 363.540 -8.580 ;
        RECT 362.700 -9.420 362.980 -9.140 ;
        RECT 361.020 -12.220 361.300 -11.940 ;
        RECT 353.180 -16.140 353.460 -15.860 ;
        RECT 360.460 -16.700 360.740 -16.420 ;
        RECT 359.340 -17.260 359.620 -16.980 ;
        RECT 361.020 -20.060 361.300 -19.780 ;
        RECT 353.180 -20.620 353.460 -20.340 ;
        RECT 349.820 -26.780 350.100 -26.500 ;
        RECT 349.260 -27.340 349.540 -27.060 ;
        RECT 350.380 -34.620 350.660 -34.340 ;
        RECT 348.140 -35.740 348.420 -35.460 ;
        RECT 351.500 -24.540 351.780 -24.260 ;
        RECT 359.340 -23.420 359.620 -23.140 ;
        RECT 353.180 -24.540 353.460 -24.260 ;
        RECT 353.740 -25.100 354.020 -24.820 ;
        RECT 358.220 -23.980 358.500 -23.700 ;
        RECT 354.300 -26.780 354.580 -26.500 ;
        RECT 353.740 -27.340 354.020 -27.060 ;
        RECT 361.580 -23.980 361.860 -23.700 ;
        RECT 366.620 -11.100 366.900 -10.820 ;
        RECT 366.060 -11.660 366.340 -11.380 ;
        RECT 366.060 -14.460 366.340 -14.180 ;
        RECT 363.260 -15.020 363.540 -14.740 ;
        RECT 363.820 -16.140 364.100 -15.860 ;
        RECT 365.500 -20.060 365.780 -19.780 ;
        RECT 367.740 0.100 368.020 0.380 ;
        RECT 385.100 30.900 385.380 31.180 ;
        RECT 383.980 30.340 384.260 30.620 ;
        RECT 387.340 42.100 387.620 42.380 ;
        RECT 387.900 38.740 388.180 39.020 ;
        RECT 386.780 30.900 387.060 31.180 ;
        RECT 391.820 42.100 392.100 42.380 ;
        RECT 390.700 38.180 390.980 38.460 ;
        RECT 389.580 34.820 389.860 35.100 ;
        RECT 386.220 30.340 386.500 30.620 ;
        RECT 384.540 29.780 384.820 30.060 ;
        RECT 386.780 23.060 387.060 23.340 ;
        RECT 404.700 38.740 404.980 39.020 ;
        RECT 391.820 26.980 392.100 27.260 ;
        RECT 385.660 22.500 385.940 22.780 ;
        RECT 383.420 19.700 383.700 19.980 ;
        RECT 387.340 21.380 387.620 21.660 ;
        RECT 382.300 19.140 382.580 19.420 ;
        RECT 381.740 14.100 382.020 14.380 ;
        RECT 381.180 12.420 381.460 12.700 ;
        RECT 377.820 11.300 378.100 11.580 ;
        RECT 387.900 19.140 388.180 19.420 ;
        RECT 383.420 18.580 383.700 18.860 ;
        RECT 389.580 19.140 389.860 19.420 ;
        RECT 392.380 19.140 392.660 19.420 ;
        RECT 393.500 32.020 393.780 32.300 ;
        RECT 383.980 18.020 384.260 18.300 ;
        RECT 382.860 14.100 383.140 14.380 ;
        RECT 386.220 12.420 386.500 12.700 ;
        RECT 382.860 11.300 383.140 11.580 ;
        RECT 388.460 12.420 388.740 12.700 ;
        RECT 393.500 26.980 393.780 27.260 ;
        RECT 404.140 19.140 404.420 19.420 ;
        RECT 400.220 16.340 400.500 16.620 ;
        RECT 393.500 15.220 393.780 15.500 ;
        RECT 392.380 11.860 392.660 12.140 ;
        RECT 371.660 2.340 371.940 2.620 ;
        RECT 373.900 2.340 374.180 2.620 ;
        RECT 368.300 -0.460 368.580 -0.180 ;
        RECT 369.420 -1.020 369.700 -0.740 ;
        RECT 372.220 -1.020 372.500 -0.740 ;
        RECT 369.420 -8.860 369.700 -8.580 ;
        RECT 368.300 -9.420 368.580 -9.140 ;
        RECT 371.100 -11.660 371.380 -11.380 ;
        RECT 369.420 -12.780 369.700 -12.500 ;
        RECT 376.140 -3.820 376.420 -3.540 ;
        RECT 372.220 -9.420 372.500 -9.140 ;
        RECT 366.060 -23.980 366.340 -23.700 ;
        RECT 367.180 -17.260 367.460 -16.980 ;
        RECT 367.180 -20.620 367.460 -20.340 ;
        RECT 370.540 -16.700 370.820 -16.420 ;
        RECT 372.220 -18.940 372.500 -18.660 ;
        RECT 372.780 -16.700 373.060 -16.420 ;
        RECT 377.260 -9.420 377.540 -9.140 ;
        RECT 380.060 -11.660 380.340 -11.380 ;
        RECT 379.500 -12.220 379.780 -11.940 ;
        RECT 376.140 -13.900 376.420 -13.620 ;
        RECT 381.180 -12.780 381.460 -12.500 ;
        RECT 380.060 -13.340 380.340 -13.060 ;
        RECT 377.820 -15.020 378.100 -14.740 ;
        RECT 378.940 -16.700 379.220 -16.420 ;
        RECT 375.580 -17.260 375.860 -16.980 ;
        RECT 371.660 -20.060 371.940 -19.780 ;
        RECT 358.780 -25.100 359.060 -24.820 ;
        RECT 354.860 -28.460 355.140 -28.180 ;
        RECT 352.060 -30.700 352.340 -30.420 ;
        RECT 354.300 -35.180 354.580 -34.900 ;
        RECT 359.900 -27.900 360.180 -27.620 ;
        RECT 364.940 -27.900 365.220 -27.620 ;
        RECT 371.100 -30.700 371.380 -30.420 ;
        RECT 366.620 -32.380 366.900 -32.100 ;
        RECT 365.500 -34.060 365.780 -33.780 ;
        RECT 359.340 -35.180 359.620 -34.900 ;
        RECT 352.620 -36.300 352.900 -36.020 ;
        RECT 347.020 -40.220 347.300 -39.940 ;
        RECT 343.100 -42.460 343.380 -42.180 ;
        RECT 344.220 -43.020 344.500 -42.740 ;
        RECT 349.820 -43.020 350.100 -42.740 ;
        RECT 344.780 -43.580 345.060 -43.300 ;
        RECT 348.700 -43.580 348.980 -43.300 ;
        RECT 347.020 -44.140 347.300 -43.860 ;
        RECT 334.140 -46.940 334.420 -46.660 ;
        RECT 306.140 -55.900 306.420 -55.620 ;
        RECT 316.220 -48.060 316.500 -47.780 ;
        RECT 322.380 -48.060 322.660 -47.780 ;
        RECT 340.860 -46.940 341.140 -46.660 ;
        RECT 352.060 -46.940 352.340 -46.660 ;
        RECT 358.780 -35.740 359.060 -35.460 ;
        RECT 363.260 -34.620 363.540 -34.340 ;
        RECT 367.180 -35.180 367.460 -34.900 ;
        RECT 364.940 -38.540 365.220 -38.260 ;
        RECT 369.420 -38.540 369.700 -38.260 ;
        RECT 376.700 -18.940 376.980 -18.660 ;
        RECT 376.140 -20.620 376.420 -20.340 ;
        RECT 372.780 -23.980 373.060 -23.700 ;
        RECT 380.620 -16.140 380.900 -15.860 ;
        RECT 376.140 -27.340 376.420 -27.060 ;
        RECT 376.140 -30.700 376.420 -30.420 ;
        RECT 372.220 -32.380 372.500 -32.100 ;
        RECT 373.900 -32.940 374.180 -32.660 ;
        RECT 373.900 -34.620 374.180 -34.340 ;
        RECT 377.820 -34.620 378.100 -34.340 ;
        RECT 371.660 -35.180 371.940 -34.900 ;
        RECT 372.780 -35.740 373.060 -35.460 ;
        RECT 359.340 -40.780 359.620 -40.500 ;
        RECT 369.980 -40.780 370.260 -40.500 ;
        RECT 357.660 -41.900 357.940 -41.620 ;
        RECT 354.860 -43.020 355.140 -42.740 ;
        RECT 382.300 2.340 382.580 2.620 ;
        RECT 386.780 2.340 387.060 2.620 ;
        RECT 386.220 -0.460 386.500 -0.180 ;
        RECT 384.540 -1.580 384.820 -1.300 ;
        RECT 383.980 -4.380 384.260 -4.100 ;
        RECT 382.300 -7.180 382.580 -6.900 ;
        RECT 387.900 -1.580 388.180 -1.300 ;
        RECT 388.460 -2.140 388.740 -1.860 ;
        RECT 396.300 15.220 396.580 15.500 ;
        RECT 399.100 14.660 399.380 14.940 ;
        RECT 397.420 14.100 397.700 14.380 ;
        RECT 401.340 10.740 401.620 11.020 ;
        RECT 402.460 10.740 402.740 11.020 ;
        RECT 422.060 46.020 422.340 46.300 ;
        RECT 413.100 45.460 413.380 45.740 ;
        RECT 412.540 41.540 412.820 41.820 ;
        RECT 412.540 35.940 412.820 36.220 ;
        RECT 408.620 33.700 408.900 33.980 ;
        RECT 409.180 32.020 409.460 32.300 ;
        RECT 408.620 30.340 408.900 30.620 ;
        RECT 426.540 46.020 426.820 46.300 ;
        RECT 418.700 42.660 418.980 42.940 ;
        RECT 417.580 42.100 417.860 42.380 ;
        RECT 416.460 41.540 416.740 41.820 ;
        RECT 415.340 38.180 415.620 38.460 ;
        RECT 417.020 38.740 417.300 39.020 ;
        RECT 419.820 38.740 420.100 39.020 ;
        RECT 411.420 26.980 411.700 27.260 ;
        RECT 407.500 21.380 407.780 21.660 ;
        RECT 407.500 19.700 407.780 19.980 ;
        RECT 404.700 16.340 404.980 16.620 ;
        RECT 404.140 12.980 404.420 13.260 ;
        RECT 406.940 12.980 407.220 13.260 ;
        RECT 403.580 7.380 403.860 7.660 ;
        RECT 407.500 10.180 407.780 10.460 ;
        RECT 410.300 10.180 410.580 10.460 ;
        RECT 406.940 7.380 407.220 7.660 ;
        RECT 391.260 6.260 391.540 6.540 ;
        RECT 407.500 6.820 407.780 7.100 ;
        RECT 396.300 6.260 396.580 6.540 ;
        RECT 403.020 6.260 403.300 6.540 ;
        RECT 406.380 6.260 406.660 6.540 ;
        RECT 392.380 4.020 392.660 4.300 ;
        RECT 394.620 3.460 394.900 3.740 ;
        RECT 389.020 2.900 389.300 3.180 ;
        RECT 387.340 -8.300 387.620 -8.020 ;
        RECT 387.900 -4.940 388.180 -4.660 ;
        RECT 385.100 -8.860 385.380 -8.580 ;
        RECT 383.420 -13.900 383.700 -13.620 ;
        RECT 385.100 -14.460 385.380 -14.180 ;
        RECT 384.540 -15.020 384.820 -14.740 ;
        RECT 384.540 -16.140 384.820 -15.860 ;
        RECT 385.100 -17.820 385.380 -17.540 ;
        RECT 385.100 -20.060 385.380 -19.780 ;
        RECT 383.980 -26.220 384.260 -25.940 ;
        RECT 385.660 -26.780 385.940 -26.500 ;
        RECT 386.780 -25.660 387.060 -25.380 ;
        RECT 386.780 -27.340 387.060 -27.060 ;
        RECT 383.980 -30.140 384.260 -29.860 ;
        RECT 381.740 -34.620 382.020 -34.340 ;
        RECT 380.060 -35.180 380.340 -34.900 ;
        RECT 382.300 -35.180 382.580 -34.900 ;
        RECT 382.300 -36.860 382.580 -36.580 ;
        RECT 380.060 -38.540 380.340 -38.260 ;
        RECT 387.900 -25.100 388.180 -24.820 ;
        RECT 387.900 -30.140 388.180 -29.860 ;
        RECT 386.780 -32.940 387.060 -32.660 ;
        RECT 391.820 0.660 392.100 0.940 ;
        RECT 397.980 3.460 398.260 3.740 ;
        RECT 390.140 -2.140 390.420 -1.860 ;
        RECT 394.620 -4.380 394.900 -4.100 ;
        RECT 390.140 -4.940 390.420 -4.660 ;
        RECT 391.260 -6.060 391.540 -5.780 ;
        RECT 389.580 -7.740 389.860 -7.460 ;
        RECT 391.820 -8.300 392.100 -8.020 ;
        RECT 390.700 -12.220 390.980 -11.940 ;
        RECT 390.140 -16.140 390.420 -15.860 ;
        RECT 396.300 -8.300 396.580 -8.020 ;
        RECT 396.860 -1.580 397.140 -1.300 ;
        RECT 398.540 0.100 398.820 0.380 ;
        RECT 409.180 1.220 409.460 1.500 ;
        RECT 399.660 -0.460 399.940 -0.180 ;
        RECT 408.620 -0.460 408.900 -0.180 ;
        RECT 407.500 -2.140 407.780 -1.860 ;
        RECT 396.860 -6.060 397.140 -5.780 ;
        RECT 395.740 -8.860 396.020 -8.580 ;
        RECT 396.300 -9.420 396.580 -9.140 ;
        RECT 397.420 -5.500 397.700 -5.220 ;
        RECT 399.660 -7.180 399.940 -6.900 ;
        RECT 401.900 -6.620 402.180 -6.340 ;
        RECT 392.380 -12.780 392.660 -12.500 ;
        RECT 400.780 -13.340 401.060 -13.060 ;
        RECT 395.740 -14.460 396.020 -14.180 ;
        RECT 392.940 -16.140 393.220 -15.860 ;
        RECT 391.820 -18.940 392.100 -18.660 ;
        RECT 391.820 -20.060 392.100 -19.780 ;
        RECT 401.900 -14.460 402.180 -14.180 ;
        RECT 397.980 -15.020 398.260 -14.740 ;
        RECT 397.980 -17.260 398.260 -16.980 ;
        RECT 391.260 -20.620 391.540 -20.340 ;
        RECT 390.700 -21.180 390.980 -20.900 ;
        RECT 395.180 -21.180 395.460 -20.900 ;
        RECT 390.700 -23.980 390.980 -23.700 ;
        RECT 389.580 -24.540 389.860 -24.260 ;
        RECT 392.380 -25.100 392.660 -24.820 ;
        RECT 395.740 -24.540 396.020 -24.260 ;
        RECT 403.580 -6.620 403.860 -6.340 ;
        RECT 404.700 -8.300 404.980 -8.020 ;
        RECT 404.140 -8.860 404.420 -8.580 ;
        RECT 404.700 -11.660 404.980 -11.380 ;
        RECT 403.020 -16.700 403.300 -16.420 ;
        RECT 406.940 -12.220 407.220 -11.940 ;
        RECT 409.180 -2.140 409.460 -1.860 ;
        RECT 408.620 -8.860 408.900 -8.580 ;
        RECT 407.500 -16.140 407.780 -15.860 ;
        RECT 408.620 -16.700 408.900 -16.420 ;
        RECT 406.380 -17.820 406.660 -17.540 ;
        RECT 403.580 -20.060 403.860 -19.780 ;
        RECT 401.900 -21.740 402.180 -21.460 ;
        RECT 415.900 32.020 416.180 32.300 ;
        RECT 423.180 42.660 423.460 42.940 ;
        RECT 423.180 38.180 423.460 38.460 ;
        RECT 422.060 35.380 422.340 35.660 ;
        RECT 418.140 33.700 418.420 33.980 ;
        RECT 415.340 26.980 415.620 27.260 ;
        RECT 417.020 26.980 417.300 27.260 ;
        RECT 420.380 26.980 420.660 27.260 ;
        RECT 418.140 26.420 418.420 26.700 ;
        RECT 427.100 41.540 427.380 41.820 ;
        RECT 424.860 39.860 425.140 40.140 ;
        RECT 427.100 39.300 427.380 39.580 ;
        RECT 428.220 38.740 428.500 39.020 ;
        RECT 427.100 32.020 427.380 32.300 ;
        RECT 421.500 26.420 421.780 26.700 ;
        RECT 418.140 22.500 418.420 22.780 ;
        RECT 418.700 21.380 418.980 21.660 ;
        RECT 410.860 -14.460 411.140 -14.180 ;
        RECT 410.860 -20.620 411.140 -20.340 ;
        RECT 410.300 -21.740 410.580 -21.460 ;
        RECT 396.860 -27.900 397.140 -27.620 ;
        RECT 406.940 -23.420 407.220 -23.140 ;
        RECT 399.660 -29.020 399.940 -28.740 ;
        RECT 401.340 -29.020 401.620 -28.740 ;
        RECT 385.100 -38.540 385.380 -38.260 ;
        RECT 389.020 -35.180 389.300 -34.900 ;
        RECT 387.900 -36.860 388.180 -36.580 ;
        RECT 390.140 -36.860 390.420 -36.580 ;
        RECT 390.700 -35.740 390.980 -35.460 ;
        RECT 383.980 -40.780 384.260 -40.500 ;
        RECT 386.220 -42.460 386.500 -42.180 ;
        RECT 391.260 -39.100 391.540 -38.820 ;
        RECT 381.180 -43.020 381.460 -42.740 ;
        RECT 403.020 -28.460 403.300 -28.180 ;
        RECT 405.260 -32.380 405.540 -32.100 ;
        RECT 359.900 -46.940 360.180 -46.660 ;
        RECT 387.900 -46.940 388.180 -46.660 ;
        RECT 369.980 -48.060 370.260 -47.780 ;
        RECT 381.740 -48.060 382.020 -47.780 ;
        RECT 397.420 -43.580 397.700 -43.300 ;
        RECT 402.460 -40.780 402.740 -40.500 ;
        RECT 412.540 -1.020 412.820 -0.740 ;
        RECT 411.980 -1.580 412.260 -1.300 ;
        RECT 411.980 -4.380 412.260 -4.100 ;
        RECT 427.100 23.060 427.380 23.340 ;
        RECT 436.060 43.220 436.340 43.500 ;
        RECT 434.940 39.860 435.220 40.140 ;
        RECT 442.780 39.300 443.060 39.580 ;
        RECT 441.100 38.740 441.380 39.020 ;
        RECT 437.740 38.180 438.020 38.460 ;
        RECT 431.580 35.940 431.860 36.220 ;
        RECT 438.860 37.620 439.140 37.900 ;
        RECT 433.820 35.380 434.100 35.660 ;
        RECT 428.780 31.460 429.060 31.740 ;
        RECT 431.580 30.340 431.860 30.620 ;
        RECT 438.300 29.780 438.580 30.060 ;
        RECT 434.380 26.980 434.660 27.260 ;
        RECT 428.780 23.060 429.060 23.340 ;
        RECT 427.660 20.260 427.940 20.540 ;
        RECT 422.620 18.580 422.900 18.860 ;
        RECT 425.980 18.580 426.260 18.860 ;
        RECT 432.140 21.940 432.420 22.220 ;
        RECT 442.220 37.620 442.500 37.900 ;
        RECT 442.780 35.940 443.060 36.220 ;
        RECT 435.500 25.860 435.780 26.140 ;
        RECT 434.940 21.940 435.220 22.220 ;
        RECT 434.380 21.380 434.660 21.660 ;
        RECT 432.700 19.700 432.980 19.980 ;
        RECT 435.500 19.700 435.780 19.980 ;
        RECT 431.580 19.140 431.860 19.420 ;
        RECT 417.020 15.220 417.300 15.500 ;
        RECT 419.820 15.220 420.100 15.500 ;
        RECT 423.740 15.220 424.020 15.500 ;
        RECT 422.620 10.740 422.900 11.020 ;
        RECT 423.180 6.820 423.460 7.100 ;
        RECT 411.980 -8.860 412.260 -8.580 ;
        RECT 411.980 -11.660 412.260 -11.380 ;
        RECT 417.020 -11.660 417.300 -11.380 ;
        RECT 412.540 -12.220 412.820 -11.940 ;
        RECT 415.340 -12.780 415.620 -12.500 ;
        RECT 417.020 -15.580 417.300 -15.300 ;
        RECT 414.780 -16.700 415.060 -16.420 ;
        RECT 411.980 -20.060 412.260 -19.780 ;
        RECT 424.860 -1.020 425.140 -0.740 ;
        RECT 423.740 -4.380 424.020 -4.100 ;
        RECT 419.820 -6.620 420.100 -6.340 ;
        RECT 422.620 -8.300 422.900 -8.020 ;
        RECT 418.700 -9.420 418.980 -9.140 ;
        RECT 419.260 -12.780 419.540 -12.500 ;
        RECT 420.940 -16.140 421.220 -15.860 ;
        RECT 418.700 -19.500 418.980 -19.220 ;
        RECT 418.140 -20.620 418.420 -20.340 ;
        RECT 421.500 -21.180 421.780 -20.900 ;
        RECT 424.300 -11.660 424.580 -11.380 ;
        RECT 433.820 15.220 434.100 15.500 ;
        RECT 426.540 12.420 426.820 12.700 ;
        RECT 429.900 14.100 430.180 14.380 ;
        RECT 428.220 12.420 428.500 12.700 ;
        RECT 432.700 12.980 432.980 13.260 ;
        RECT 436.620 23.060 436.900 23.340 ;
        RECT 436.060 15.220 436.340 15.500 ;
        RECT 434.940 14.100 435.220 14.380 ;
        RECT 433.820 10.740 434.100 11.020 ;
        RECT 432.700 10.180 432.980 10.460 ;
        RECT 426.540 4.580 426.820 4.860 ;
        RECT 428.220 4.020 428.500 4.300 ;
        RECT 432.140 4.020 432.420 4.300 ;
        RECT 427.100 -8.300 427.380 -8.020 ;
        RECT 428.780 -11.100 429.060 -10.820 ;
        RECT 429.340 -11.660 429.620 -11.380 ;
        RECT 433.820 7.940 434.100 8.220 ;
        RECT 435.500 14.660 435.780 14.940 ;
        RECT 440.540 23.060 440.820 23.340 ;
        RECT 438.860 21.380 439.140 21.660 ;
        RECT 437.180 19.700 437.460 19.980 ;
        RECT 442.220 19.700 442.500 19.980 ;
        RECT 439.420 16.340 439.700 16.620 ;
        RECT 437.740 14.660 438.020 14.940 ;
        RECT 439.980 14.660 440.260 14.940 ;
        RECT 438.860 12.980 439.140 13.260 ;
        RECT 436.620 7.940 436.900 8.220 ;
        RECT 435.500 1.220 435.780 1.500 ;
        RECT 435.500 -0.460 435.780 -0.180 ;
        RECT 437.180 0.660 437.460 0.940 ;
        RECT 432.700 -6.620 432.980 -6.340 ;
        RECT 442.220 14.660 442.500 14.940 ;
        RECT 443.340 30.900 443.620 31.180 ;
        RECT 444.460 42.100 444.740 42.380 ;
        RECT 445.580 38.740 445.860 39.020 ;
        RECT 457.340 41.540 457.620 41.820 ;
        RECT 448.380 35.940 448.660 36.220 ;
        RECT 446.140 29.780 446.420 30.060 ;
        RECT 446.140 21.940 446.420 22.220 ;
        RECT 455.100 30.900 455.380 31.180 ;
        RECT 459.020 32.020 459.300 32.300 ;
        RECT 458.460 31.460 458.740 31.740 ;
        RECT 455.660 30.340 455.940 30.620 ;
        RECT 453.980 29.780 454.260 30.060 ;
        RECT 457.900 30.900 458.180 31.180 ;
        RECT 458.460 29.220 458.740 29.500 ;
        RECT 459.580 29.780 459.860 30.060 ;
        RECT 454.540 25.860 454.820 26.140 ;
        RECT 449.500 20.260 449.780 20.540 ;
        RECT 447.820 19.700 448.100 19.980 ;
        RECT 446.140 6.820 446.420 7.100 ;
        RECT 442.780 2.340 443.060 2.620 ;
        RECT 436.620 -7.180 436.900 -6.900 ;
        RECT 438.300 -7.740 438.580 -7.460 ;
        RECT 443.340 -7.740 443.620 -7.460 ;
        RECT 431.580 -10.540 431.860 -10.260 ;
        RECT 418.140 -23.420 418.420 -23.140 ;
        RECT 423.740 -16.140 424.020 -15.860 ;
        RECT 412.540 -23.980 412.820 -23.700 ;
        RECT 418.700 -23.980 418.980 -23.700 ;
        RECT 418.140 -24.540 418.420 -24.260 ;
        RECT 413.100 -25.660 413.380 -25.380 ;
        RECT 413.100 -27.900 413.380 -27.620 ;
        RECT 420.380 -25.100 420.660 -24.820 ;
        RECT 422.060 -27.340 422.340 -27.060 ;
        RECT 411.420 -35.740 411.700 -35.460 ;
        RECT 415.340 -29.580 415.620 -29.300 ;
        RECT 419.820 -29.580 420.100 -29.300 ;
        RECT 422.060 -32.380 422.340 -32.100 ;
        RECT 425.420 -19.500 425.700 -19.220 ;
        RECT 430.460 -12.220 430.740 -11.940 ;
        RECT 441.100 -12.220 441.380 -11.940 ;
        RECT 425.980 -27.340 426.260 -27.060 ;
        RECT 423.180 -31.260 423.460 -30.980 ;
        RECT 423.740 -35.180 424.020 -34.900 ;
        RECT 422.620 -36.860 422.900 -36.580 ;
        RECT 424.860 -31.820 425.140 -31.540 ;
        RECT 418.140 -38.540 418.420 -38.260 ;
        RECT 437.180 -18.940 437.460 -18.660 ;
        RECT 432.140 -20.060 432.420 -19.780 ;
        RECT 431.580 -23.420 431.860 -23.140 ;
        RECT 426.540 -31.820 426.820 -31.540 ;
        RECT 431.580 -28.460 431.860 -28.180 ;
        RECT 430.460 -31.260 430.740 -30.980 ;
        RECT 428.780 -31.820 429.060 -31.540 ;
        RECT 432.140 -32.380 432.420 -32.100 ;
        RECT 427.660 -32.940 427.940 -32.660 ;
        RECT 423.180 -38.540 423.460 -38.260 ;
        RECT 414.780 -40.780 415.060 -40.500 ;
        RECT 418.700 -40.220 418.980 -39.940 ;
        RECT 402.460 -42.460 402.740 -42.180 ;
        RECT 423.740 -40.220 424.020 -39.940 ;
        RECT 431.020 -32.940 431.300 -32.660 ;
        RECT 436.620 -20.060 436.900 -19.780 ;
        RECT 436.620 -21.180 436.900 -20.900 ;
        RECT 432.700 -33.500 432.980 -33.220 ;
        RECT 431.020 -39.660 431.300 -39.380 ;
        RECT 421.500 -43.580 421.780 -43.300 ;
        RECT 398.540 -46.940 398.820 -46.660 ;
        RECT 405.820 -46.940 406.100 -46.660 ;
        RECT 389.580 -47.500 389.860 -47.220 ;
        RECT 392.940 -47.500 393.220 -47.220 ;
        RECT 417.020 -46.940 417.300 -46.660 ;
        RECT 433.260 -21.740 433.540 -21.460 ;
        RECT 432.700 -35.180 432.980 -34.900 ;
        RECT 435.500 -23.420 435.780 -23.140 ;
        RECT 438.300 -24.540 438.580 -24.260 ;
        RECT 434.380 -30.700 434.660 -30.420 ;
        RECT 437.180 -31.260 437.460 -30.980 ;
        RECT 435.500 -35.740 435.780 -35.460 ;
        RECT 439.980 -31.820 440.260 -31.540 ;
        RECT 443.340 -11.100 443.620 -10.820 ;
        RECT 454.540 3.460 454.820 3.740 ;
        RECT 455.660 23.060 455.940 23.340 ;
        RECT 457.340 21.940 457.620 22.220 ;
        RECT 457.340 16.340 457.620 16.620 ;
        RECT 460.140 29.220 460.420 29.500 ;
        RECT 445.020 -7.180 445.300 -6.900 ;
        RECT 448.380 -10.540 448.660 -10.260 ;
        RECT 446.140 -11.100 446.420 -10.820 ;
        RECT 440.540 -32.380 440.820 -32.100 ;
        RECT 437.180 -32.940 437.460 -32.660 ;
        RECT 442.220 -33.500 442.500 -33.220 ;
        RECT 437.180 -35.740 437.460 -35.460 ;
        RECT 436.620 -38.540 436.900 -38.260 ;
        RECT 438.860 -40.220 439.140 -39.940 ;
        RECT 445.020 -31.820 445.300 -31.540 ;
        RECT 444.460 -32.380 444.740 -32.100 ;
        RECT 445.020 -32.940 445.300 -32.660 ;
        RECT 443.900 -36.300 444.180 -36.020 ;
        RECT 449.500 -17.260 449.780 -16.980 ;
        RECT 447.260 -26.780 447.540 -26.500 ;
        RECT 452.300 -18.940 452.580 -18.660 ;
        RECT 453.420 -20.060 453.700 -19.780 ;
        RECT 449.500 -32.380 449.780 -32.100 ;
        RECT 446.140 -34.620 446.420 -34.340 ;
        RECT 448.380 -34.620 448.660 -34.340 ;
        RECT 446.700 -36.300 446.980 -36.020 ;
        RECT 445.580 -36.860 445.860 -36.580 ;
        RECT 450.060 -28.460 450.340 -28.180 ;
        RECT 451.180 -34.620 451.460 -34.340 ;
        RECT 449.500 -38.540 449.780 -38.260 ;
        RECT 453.420 -39.100 453.700 -38.820 ;
        RECT 432.140 -43.580 432.420 -43.300 ;
        RECT 431.580 -44.140 431.860 -43.860 ;
        RECT 427.100 -46.380 427.380 -46.100 ;
        RECT 419.260 -47.500 419.540 -47.220 ;
        RECT 423.740 -46.940 424.020 -46.660 ;
        RECT 436.060 -46.940 436.340 -46.660 ;
        RECT 432.140 -47.500 432.420 -47.220 ;
        RECT 121.025 -64.055 121.825 -63.775 ;
        RECT 97.375 -67.115 97.655 -66.835 ;
        RECT 97.375 -67.715 97.655 -67.435 ;
        RECT 121.025 -67.415 121.825 -67.135 ;
        RECT 96.255 -70.475 96.535 -70.195 ;
        RECT 96.255 -71.075 96.535 -70.795 ;
        RECT 121.025 -70.775 121.825 -70.495 ;
        RECT 94.015 -73.835 94.295 -73.555 ;
        RECT 94.015 -74.435 94.295 -74.155 ;
        RECT 121.025 -74.135 121.825 -73.855 ;
        RECT 89.535 -77.195 89.815 -76.915 ;
        RECT 89.535 -77.795 89.815 -77.515 ;
        RECT 121.025 -77.495 121.825 -77.215 ;
        RECT 80.575 -80.555 80.855 -80.275 ;
        RECT 80.575 -81.155 80.855 -80.875 ;
        RECT 121.025 -80.855 121.825 -80.575 ;
        RECT 62.655 -83.915 62.935 -83.635 ;
        RECT 62.655 -84.515 62.935 -84.235 ;
        RECT 121.025 -84.215 121.825 -83.935 ;
        RECT 26.815 -87.275 27.095 -86.995 ;
        RECT 26.815 -87.875 27.095 -87.595 ;
        RECT 121.025 -87.575 121.825 -87.295 ;
        RECT 457.340 -0.460 457.620 -0.180 ;
        RECT 459.580 -1.020 459.860 -0.740 ;
        RECT 455.100 -11.660 455.380 -11.380 ;
        RECT 460.700 -9.420 460.980 -9.140 ;
        RECT 456.220 -17.260 456.500 -16.980 ;
        RECT 468.280 -19.500 468.560 -19.220 ;
        RECT 468.840 -19.500 469.120 -19.220 ;
        RECT 459.020 -20.060 459.300 -19.780 ;
        RECT 456.780 -30.700 457.060 -30.420 ;
        RECT 455.100 -34.620 455.380 -34.340 ;
        RECT 455.100 -36.300 455.380 -36.020 ;
        RECT 454.540 -44.140 454.820 -43.860 ;
        RECT 468.280 -20.060 468.560 -19.780 ;
        RECT 468.840 -20.060 469.120 -19.780 ;
        RECT 468.280 -20.620 468.560 -20.340 ;
        RECT 468.840 -20.620 469.120 -20.340 ;
        RECT 459.580 -30.700 459.860 -30.420 ;
        RECT 460.140 -29.020 460.420 -28.740 ;
        RECT 458.460 -31.260 458.740 -30.980 ;
        RECT 456.780 -32.380 457.060 -32.100 ;
        RECT 457.900 -36.860 458.180 -36.580 ;
        RECT 457.340 -37.980 457.620 -37.700 ;
        RECT 460.700 -32.940 460.980 -32.660 ;
        RECT 460.140 -36.300 460.420 -36.020 ;
        RECT 459.580 -46.380 459.860 -46.100 ;
        RECT -44.865 -90.635 -44.585 -90.355 ;
        RECT -44.865 -91.235 -44.585 -90.955 ;
        RECT 121.025 -90.935 121.825 -90.655 ;
        RECT -188.225 -93.995 -187.945 -93.715 ;
        RECT -188.225 -94.595 -187.945 -94.315 ;
        RECT 121.025 -94.295 121.825 -94.015 ;
        RECT -189.345 -97.355 -189.065 -97.075 ;
        RECT -189.345 -97.955 -189.065 -97.675 ;
        RECT 121.025 -97.655 121.825 -97.375 ;
        RECT -492.030 -106.165 -491.230 -105.885 ;
        RECT 467.250 -105.885 467.530 -105.605 ;
        RECT 467.810 -105.885 468.090 -105.605 ;
        RECT 468.370 -105.885 468.650 -105.605 ;
        RECT 467.250 -106.445 467.530 -106.165 ;
        RECT 467.810 -106.445 468.090 -106.165 ;
        RECT 468.370 -106.445 468.650 -106.165 ;
      LAYER Metal3 ;
        RECT 135.505 106.425 469.200 106.525 ;
        RECT -492.150 105.625 469.200 106.425 ;
        RECT 135.505 105.525 469.200 105.625 ;
        RECT -189.405 96.915 -189.005 98.115 ;
        RECT 120.925 97.265 121.925 97.765 ;
        RECT -188.285 93.555 -187.885 94.755 ;
        RECT 115.555 93.955 116.755 94.355 ;
        RECT -332.765 90.195 -332.365 91.395 ;
        RECT -44.925 90.195 -44.525 91.395 ;
        RECT 113.755 90.595 114.955 90.995 ;
        RECT -404.445 86.835 -404.045 88.035 ;
        RECT -261.085 86.835 -260.685 88.035 ;
        RECT -116.605 86.835 -116.205 88.035 ;
        RECT 26.755 86.835 27.155 88.035 ;
        RECT 111.955 87.235 113.155 87.635 ;
        RECT -497.595 83.365 -495.515 83.765 ;
        RECT -440.285 83.475 -439.885 84.675 ;
        RECT -368.605 83.475 -368.205 84.675 ;
        RECT -296.925 83.475 -296.525 84.675 ;
        RECT -225.245 83.475 -224.845 84.675 ;
        RECT -152.445 83.475 -152.045 84.675 ;
        RECT -80.765 83.475 -80.365 84.675 ;
        RECT -9.085 83.475 -8.685 84.675 ;
        RECT 62.595 83.475 62.995 84.675 ;
        RECT 110.155 83.875 111.355 84.275 ;
        RECT -486.955 81.155 -486.555 83.235 ;
        RECT -458.205 80.115 -457.805 81.315 ;
        RECT -422.365 80.115 -421.965 81.315 ;
        RECT -386.525 80.115 -386.125 81.315 ;
        RECT -350.685 80.115 -350.285 81.315 ;
        RECT -314.845 80.115 -314.445 81.315 ;
        RECT -279.005 80.115 -278.605 81.315 ;
        RECT -243.165 80.115 -242.765 81.315 ;
        RECT -207.325 80.115 -206.925 81.315 ;
        RECT -170.365 80.115 -169.965 81.315 ;
        RECT -134.525 80.115 -134.125 81.315 ;
        RECT -98.685 80.115 -98.285 81.315 ;
        RECT -62.845 80.115 -62.445 81.315 ;
        RECT -27.005 80.115 -26.605 81.315 ;
        RECT 8.835 80.115 9.235 81.315 ;
        RECT 44.675 80.115 45.075 81.315 ;
        RECT 80.515 80.115 80.915 81.315 ;
        RECT 108.355 80.515 109.555 80.915 ;
        RECT -467.165 76.755 -466.765 77.955 ;
        RECT -449.245 76.755 -448.845 77.955 ;
        RECT -431.325 76.755 -430.925 77.955 ;
        RECT -413.405 76.755 -413.005 77.955 ;
        RECT -395.485 76.755 -395.085 77.955 ;
        RECT -377.565 76.755 -377.165 77.955 ;
        RECT -359.645 76.755 -359.245 77.955 ;
        RECT -341.725 76.755 -341.325 77.955 ;
        RECT -323.805 76.755 -323.405 77.955 ;
        RECT -305.885 76.755 -305.485 77.955 ;
        RECT -287.965 76.755 -287.565 77.955 ;
        RECT -270.045 76.755 -269.645 77.955 ;
        RECT -252.125 76.755 -251.725 77.955 ;
        RECT -234.205 76.755 -233.805 77.955 ;
        RECT -216.285 76.755 -215.885 77.955 ;
        RECT -198.365 76.755 -197.965 77.955 ;
        RECT -179.325 76.755 -178.925 77.955 ;
        RECT -161.405 76.755 -161.005 77.955 ;
        RECT -143.485 76.755 -143.085 77.955 ;
        RECT -125.565 76.755 -125.165 77.955 ;
        RECT -107.645 76.755 -107.245 77.955 ;
        RECT -89.725 76.755 -89.325 77.955 ;
        RECT -71.805 76.755 -71.405 77.955 ;
        RECT -53.885 76.755 -53.485 77.955 ;
        RECT -35.965 76.755 -35.565 77.955 ;
        RECT -18.045 76.755 -17.645 77.955 ;
        RECT -0.125 76.755 0.275 77.955 ;
        RECT 17.795 76.755 18.195 77.955 ;
        RECT 35.715 76.755 36.115 77.955 ;
        RECT 53.635 76.755 54.035 77.955 ;
        RECT 71.555 76.755 71.955 77.955 ;
        RECT 89.475 76.755 89.875 77.955 ;
        RECT 106.555 77.155 107.755 77.555 ;
        RECT -471.645 73.395 -471.245 74.595 ;
        RECT -462.685 73.395 -462.285 74.595 ;
        RECT -453.725 73.395 -453.325 74.595 ;
        RECT -444.765 73.395 -444.365 74.595 ;
        RECT -435.805 73.395 -435.405 74.595 ;
        RECT -426.845 73.395 -426.445 74.595 ;
        RECT -417.885 73.395 -417.485 74.595 ;
        RECT -408.925 73.395 -408.525 74.595 ;
        RECT -399.965 73.395 -399.565 74.595 ;
        RECT -391.005 73.395 -390.605 74.595 ;
        RECT -382.045 73.395 -381.645 74.595 ;
        RECT -373.085 73.395 -372.685 74.595 ;
        RECT -364.125 73.395 -363.725 74.595 ;
        RECT -355.165 73.395 -354.765 74.595 ;
        RECT -346.205 73.395 -345.805 74.595 ;
        RECT -337.245 73.395 -336.845 74.595 ;
        RECT -328.285 73.395 -327.885 74.595 ;
        RECT -319.325 73.395 -318.925 74.595 ;
        RECT -310.365 73.395 -309.965 74.595 ;
        RECT -301.405 73.395 -301.005 74.595 ;
        RECT -292.445 73.395 -292.045 74.595 ;
        RECT -283.485 73.395 -283.085 74.595 ;
        RECT -274.525 73.395 -274.125 74.595 ;
        RECT -265.565 73.395 -265.165 74.595 ;
        RECT -256.605 73.395 -256.205 74.595 ;
        RECT -247.645 73.395 -247.245 74.595 ;
        RECT -238.685 73.395 -238.285 74.595 ;
        RECT -229.725 73.395 -229.325 74.595 ;
        RECT -220.765 73.395 -220.365 74.595 ;
        RECT -211.805 73.395 -211.405 74.595 ;
        RECT -202.845 73.395 -202.445 74.595 ;
        RECT -193.885 73.395 -193.485 74.595 ;
        RECT -183.805 73.395 -183.405 74.595 ;
        RECT -174.845 73.395 -174.445 74.595 ;
        RECT -165.885 73.395 -165.485 74.595 ;
        RECT -156.925 73.395 -156.525 74.595 ;
        RECT -147.965 73.395 -147.565 74.595 ;
        RECT -139.005 73.395 -138.605 74.595 ;
        RECT -130.045 73.395 -129.645 74.595 ;
        RECT -121.085 73.395 -120.685 74.595 ;
        RECT -112.125 73.395 -111.725 74.595 ;
        RECT -103.165 73.395 -102.765 74.595 ;
        RECT -94.205 73.395 -93.805 74.595 ;
        RECT -85.245 73.395 -84.845 74.595 ;
        RECT -76.285 73.395 -75.885 74.595 ;
        RECT -67.325 73.395 -66.925 74.595 ;
        RECT -58.365 73.395 -57.965 74.595 ;
        RECT -49.405 73.395 -49.005 74.595 ;
        RECT -40.445 73.395 -40.045 74.595 ;
        RECT -31.485 73.395 -31.085 74.595 ;
        RECT -22.525 73.395 -22.125 74.595 ;
        RECT -13.565 73.395 -13.165 74.595 ;
        RECT -4.605 73.395 -4.205 74.595 ;
        RECT 4.355 73.395 4.755 74.595 ;
        RECT 13.315 73.395 13.715 74.595 ;
        RECT 22.275 73.395 22.675 74.595 ;
        RECT 31.235 73.395 31.635 74.595 ;
        RECT 40.195 73.395 40.595 74.595 ;
        RECT 49.155 73.395 49.555 74.595 ;
        RECT 58.115 73.395 58.515 74.595 ;
        RECT 67.075 73.395 67.475 74.595 ;
        RECT 76.035 73.395 76.435 74.595 ;
        RECT 84.995 73.395 85.395 74.595 ;
        RECT 93.955 73.395 94.355 74.595 ;
        RECT 104.755 73.795 105.955 74.195 ;
        RECT -473.885 70.035 -473.485 71.235 ;
        RECT -469.405 70.035 -469.005 71.235 ;
        RECT -464.925 70.035 -464.525 71.235 ;
        RECT -460.445 70.035 -460.045 71.235 ;
        RECT -455.965 70.035 -455.565 71.235 ;
        RECT -451.485 70.035 -451.085 71.235 ;
        RECT -447.005 70.035 -446.605 71.235 ;
        RECT -442.525 70.035 -442.125 71.235 ;
        RECT -438.045 70.035 -437.645 71.235 ;
        RECT -433.565 70.035 -433.165 71.235 ;
        RECT -429.085 70.035 -428.685 71.235 ;
        RECT -424.605 70.035 -424.205 71.235 ;
        RECT -420.125 70.035 -419.725 71.235 ;
        RECT -415.645 70.035 -415.245 71.235 ;
        RECT -411.165 70.035 -410.765 71.235 ;
        RECT -406.685 70.035 -406.285 71.235 ;
        RECT -402.205 70.035 -401.805 71.235 ;
        RECT -397.725 70.035 -397.325 71.235 ;
        RECT -393.245 70.035 -392.845 71.235 ;
        RECT -388.765 70.035 -388.365 71.235 ;
        RECT -384.285 70.035 -383.885 71.235 ;
        RECT -379.805 70.035 -379.405 71.235 ;
        RECT -375.325 70.035 -374.925 71.235 ;
        RECT -370.845 70.035 -370.445 71.235 ;
        RECT -366.365 70.035 -365.965 71.235 ;
        RECT -361.885 70.035 -361.485 71.235 ;
        RECT -357.405 70.035 -357.005 71.235 ;
        RECT -352.925 70.035 -352.525 71.235 ;
        RECT -348.445 70.035 -348.045 71.235 ;
        RECT -343.965 70.035 -343.565 71.235 ;
        RECT -339.485 70.035 -339.085 71.235 ;
        RECT -335.005 70.035 -334.605 71.235 ;
        RECT -330.525 70.035 -330.125 71.235 ;
        RECT -326.045 70.035 -325.645 71.235 ;
        RECT -321.565 70.035 -321.165 71.235 ;
        RECT -317.085 70.035 -316.685 71.235 ;
        RECT -312.605 70.035 -312.205 71.235 ;
        RECT -308.125 70.035 -307.725 71.235 ;
        RECT -303.645 70.035 -303.245 71.235 ;
        RECT -299.165 70.035 -298.765 71.235 ;
        RECT -294.685 70.035 -294.285 71.235 ;
        RECT -290.205 70.035 -289.805 71.235 ;
        RECT -285.725 70.035 -285.325 71.235 ;
        RECT -281.245 70.035 -280.845 71.235 ;
        RECT -276.765 70.035 -276.365 71.235 ;
        RECT -272.285 70.035 -271.885 71.235 ;
        RECT -267.805 70.035 -267.405 71.235 ;
        RECT -263.325 70.035 -262.925 71.235 ;
        RECT -258.845 70.035 -258.445 71.235 ;
        RECT -254.365 70.035 -253.965 71.235 ;
        RECT -249.885 70.035 -249.485 71.235 ;
        RECT -245.405 70.035 -245.005 71.235 ;
        RECT -240.925 70.035 -240.525 71.235 ;
        RECT -236.445 70.035 -236.045 71.235 ;
        RECT -231.965 70.035 -231.565 71.235 ;
        RECT -227.485 70.035 -227.085 71.235 ;
        RECT -223.005 70.035 -222.605 71.235 ;
        RECT -218.525 70.035 -218.125 71.235 ;
        RECT -214.045 70.035 -213.645 71.235 ;
        RECT -209.565 70.035 -209.165 71.235 ;
        RECT -205.085 70.035 -204.685 71.235 ;
        RECT -200.605 70.035 -200.205 71.235 ;
        RECT -196.125 70.035 -195.725 71.235 ;
        RECT -191.645 70.035 -191.245 71.235 ;
        RECT -186.045 70.035 -185.645 71.235 ;
        RECT -181.565 70.035 -181.165 71.235 ;
        RECT -177.085 70.035 -176.685 71.235 ;
        RECT -172.605 70.035 -172.205 71.235 ;
        RECT -168.125 70.035 -167.725 71.235 ;
        RECT -163.645 70.035 -163.245 71.235 ;
        RECT -159.165 70.035 -158.765 71.235 ;
        RECT -154.685 70.035 -154.285 71.235 ;
        RECT -150.205 70.035 -149.805 71.235 ;
        RECT -145.725 70.035 -145.325 71.235 ;
        RECT -141.245 70.035 -140.845 71.235 ;
        RECT -136.765 70.035 -136.365 71.235 ;
        RECT -132.285 70.035 -131.885 71.235 ;
        RECT -127.805 70.035 -127.405 71.235 ;
        RECT -123.325 70.035 -122.925 71.235 ;
        RECT -118.845 70.035 -118.445 71.235 ;
        RECT -114.365 70.035 -113.965 71.235 ;
        RECT -109.885 70.035 -109.485 71.235 ;
        RECT -105.405 70.035 -105.005 71.235 ;
        RECT -100.925 70.035 -100.525 71.235 ;
        RECT -96.445 70.035 -96.045 71.235 ;
        RECT -91.965 70.035 -91.565 71.235 ;
        RECT -87.485 70.035 -87.085 71.235 ;
        RECT -83.005 70.035 -82.605 71.235 ;
        RECT -78.525 70.035 -78.125 71.235 ;
        RECT -74.045 70.035 -73.645 71.235 ;
        RECT -69.565 70.035 -69.165 71.235 ;
        RECT -65.085 70.035 -64.685 71.235 ;
        RECT -60.605 70.035 -60.205 71.235 ;
        RECT -56.125 70.035 -55.725 71.235 ;
        RECT -51.645 70.035 -51.245 71.235 ;
        RECT -47.165 70.035 -46.765 71.235 ;
        RECT -42.685 70.035 -42.285 71.235 ;
        RECT -38.205 70.035 -37.805 71.235 ;
        RECT -33.725 70.035 -33.325 71.235 ;
        RECT -29.245 70.035 -28.845 71.235 ;
        RECT -24.765 70.035 -24.365 71.235 ;
        RECT -20.285 70.035 -19.885 71.235 ;
        RECT -15.805 70.035 -15.405 71.235 ;
        RECT -11.325 70.035 -10.925 71.235 ;
        RECT -6.845 70.035 -6.445 71.235 ;
        RECT -2.365 70.035 -1.965 71.235 ;
        RECT 2.115 70.035 2.515 71.235 ;
        RECT 6.595 70.035 6.995 71.235 ;
        RECT 11.075 70.035 11.475 71.235 ;
        RECT 15.555 70.035 15.955 71.235 ;
        RECT 20.035 70.035 20.435 71.235 ;
        RECT 24.515 70.035 24.915 71.235 ;
        RECT 28.995 70.035 29.395 71.235 ;
        RECT 33.475 70.035 33.875 71.235 ;
        RECT 37.955 70.035 38.355 71.235 ;
        RECT 42.435 70.035 42.835 71.235 ;
        RECT 46.915 70.035 47.315 71.235 ;
        RECT 51.395 70.035 51.795 71.235 ;
        RECT 55.875 70.035 56.275 71.235 ;
        RECT 60.355 70.035 60.755 71.235 ;
        RECT 64.835 70.035 65.235 71.235 ;
        RECT 69.315 70.035 69.715 71.235 ;
        RECT 73.795 70.035 74.195 71.235 ;
        RECT 78.275 70.035 78.675 71.235 ;
        RECT 82.755 70.035 83.155 71.235 ;
        RECT 87.235 70.035 87.635 71.235 ;
        RECT 91.715 70.035 92.115 71.235 ;
        RECT 96.195 70.035 96.595 71.235 ;
        RECT 102.955 70.435 104.155 70.835 ;
        RECT -475.005 66.675 -474.605 67.875 ;
        RECT -472.765 66.675 -472.365 67.875 ;
        RECT -470.525 66.675 -470.125 67.875 ;
        RECT -468.285 66.675 -467.885 67.875 ;
        RECT -466.045 66.675 -465.645 67.875 ;
        RECT -463.805 66.675 -463.405 67.875 ;
        RECT -461.565 66.675 -461.165 67.875 ;
        RECT -459.325 66.675 -458.925 67.875 ;
        RECT -457.085 66.675 -456.685 67.875 ;
        RECT -454.845 66.675 -454.445 67.875 ;
        RECT -452.605 66.675 -452.205 67.875 ;
        RECT -450.365 66.675 -449.965 67.875 ;
        RECT -448.125 66.675 -447.725 67.875 ;
        RECT -445.885 66.675 -445.485 67.875 ;
        RECT -443.645 66.675 -443.245 67.875 ;
        RECT -441.405 66.675 -441.005 67.875 ;
        RECT -439.165 66.675 -438.765 67.875 ;
        RECT -436.925 66.675 -436.525 67.875 ;
        RECT -434.685 66.675 -434.285 67.875 ;
        RECT -432.445 66.675 -432.045 67.875 ;
        RECT -430.205 66.675 -429.805 67.875 ;
        RECT -427.965 66.675 -427.565 67.875 ;
        RECT -425.725 66.675 -425.325 67.875 ;
        RECT -423.485 66.675 -423.085 67.875 ;
        RECT -421.245 66.675 -420.845 67.875 ;
        RECT -419.005 66.675 -418.605 67.875 ;
        RECT -416.765 66.675 -416.365 67.875 ;
        RECT -414.525 66.675 -414.125 67.875 ;
        RECT -412.285 66.675 -411.885 67.875 ;
        RECT -410.045 66.675 -409.645 67.875 ;
        RECT -407.805 66.675 -407.405 67.875 ;
        RECT -405.565 66.675 -405.165 67.875 ;
        RECT -403.325 66.675 -402.925 67.875 ;
        RECT -401.085 66.675 -400.685 67.875 ;
        RECT -398.845 66.675 -398.445 67.875 ;
        RECT -396.605 66.675 -396.205 67.875 ;
        RECT -394.365 66.675 -393.965 67.875 ;
        RECT -392.125 66.675 -391.725 67.875 ;
        RECT -389.885 66.675 -389.485 67.875 ;
        RECT -387.645 66.675 -387.245 67.875 ;
        RECT -385.405 66.675 -385.005 67.875 ;
        RECT -383.165 66.675 -382.765 67.875 ;
        RECT -380.925 66.675 -380.525 67.875 ;
        RECT -378.685 66.675 -378.285 67.875 ;
        RECT -376.445 66.675 -376.045 67.875 ;
        RECT -374.205 66.675 -373.805 67.875 ;
        RECT -371.965 66.675 -371.565 67.875 ;
        RECT -369.725 66.675 -369.325 67.875 ;
        RECT -367.485 66.675 -367.085 67.875 ;
        RECT -365.245 66.675 -364.845 67.875 ;
        RECT -363.005 66.675 -362.605 67.875 ;
        RECT -360.765 66.675 -360.365 67.875 ;
        RECT -358.525 66.675 -358.125 67.875 ;
        RECT -356.285 66.675 -355.885 67.875 ;
        RECT -354.045 66.675 -353.645 67.875 ;
        RECT -351.805 66.675 -351.405 67.875 ;
        RECT -349.565 66.675 -349.165 67.875 ;
        RECT -347.325 66.675 -346.925 67.875 ;
        RECT -345.085 66.675 -344.685 67.875 ;
        RECT -342.845 66.675 -342.445 67.875 ;
        RECT -340.605 66.675 -340.205 67.875 ;
        RECT -338.365 66.675 -337.965 67.875 ;
        RECT -336.125 66.675 -335.725 67.875 ;
        RECT -333.885 66.675 -333.485 67.875 ;
        RECT -331.645 66.675 -331.245 67.875 ;
        RECT -329.405 66.675 -329.005 67.875 ;
        RECT -327.165 66.675 -326.765 67.875 ;
        RECT -324.925 66.675 -324.525 67.875 ;
        RECT -322.685 66.675 -322.285 67.875 ;
        RECT -320.445 66.675 -320.045 67.875 ;
        RECT -318.205 66.675 -317.805 67.875 ;
        RECT -315.965 66.675 -315.565 67.875 ;
        RECT -313.725 66.675 -313.325 67.875 ;
        RECT -311.485 66.675 -311.085 67.875 ;
        RECT -309.245 66.675 -308.845 67.875 ;
        RECT -307.005 66.675 -306.605 67.875 ;
        RECT -304.765 66.675 -304.365 67.875 ;
        RECT -302.525 66.675 -302.125 67.875 ;
        RECT -300.285 66.675 -299.885 67.875 ;
        RECT -298.045 66.675 -297.645 67.875 ;
        RECT -295.805 66.675 -295.405 67.875 ;
        RECT -293.565 66.675 -293.165 67.875 ;
        RECT -291.325 66.675 -290.925 67.875 ;
        RECT -289.085 66.675 -288.685 67.875 ;
        RECT -286.845 66.675 -286.445 67.875 ;
        RECT -284.605 66.675 -284.205 67.875 ;
        RECT -282.365 66.675 -281.965 67.875 ;
        RECT -280.125 66.675 -279.725 67.875 ;
        RECT -277.885 66.675 -277.485 67.875 ;
        RECT -275.645 66.675 -275.245 67.875 ;
        RECT -273.405 66.675 -273.005 67.875 ;
        RECT -271.165 66.675 -270.765 67.875 ;
        RECT -268.925 66.675 -268.525 67.875 ;
        RECT -266.685 66.675 -266.285 67.875 ;
        RECT -264.445 66.675 -264.045 67.875 ;
        RECT -262.205 66.675 -261.805 67.875 ;
        RECT -259.965 66.675 -259.565 67.875 ;
        RECT -257.725 66.675 -257.325 67.875 ;
        RECT -255.485 66.675 -255.085 67.875 ;
        RECT -253.245 66.675 -252.845 67.875 ;
        RECT -251.005 66.675 -250.605 67.875 ;
        RECT -248.765 66.675 -248.365 67.875 ;
        RECT -246.525 66.675 -246.125 67.875 ;
        RECT -244.285 66.675 -243.885 67.875 ;
        RECT -242.045 66.675 -241.645 67.875 ;
        RECT -239.805 66.675 -239.405 67.875 ;
        RECT -237.565 66.675 -237.165 67.875 ;
        RECT -235.325 66.675 -234.925 67.875 ;
        RECT -233.085 66.675 -232.685 67.875 ;
        RECT -230.845 66.675 -230.445 67.875 ;
        RECT -228.605 66.675 -228.205 67.875 ;
        RECT -226.365 66.675 -225.965 67.875 ;
        RECT -224.125 66.675 -223.725 67.875 ;
        RECT -221.885 66.675 -221.485 67.875 ;
        RECT -219.645 66.675 -219.245 67.875 ;
        RECT -217.405 66.675 -217.005 67.875 ;
        RECT -215.165 66.675 -214.765 67.875 ;
        RECT -212.925 66.675 -212.525 67.875 ;
        RECT -210.685 66.675 -210.285 67.875 ;
        RECT -208.445 66.675 -208.045 67.875 ;
        RECT -206.205 66.675 -205.805 67.875 ;
        RECT -203.965 66.675 -203.565 67.875 ;
        RECT -201.725 66.675 -201.325 67.875 ;
        RECT -199.485 66.675 -199.085 67.875 ;
        RECT -197.245 66.675 -196.845 67.875 ;
        RECT -195.005 66.675 -194.605 67.875 ;
        RECT -192.765 66.675 -192.365 67.875 ;
        RECT -190.525 66.675 -190.125 67.875 ;
        RECT -187.165 66.675 -186.765 67.875 ;
        RECT -184.925 66.675 -184.525 67.875 ;
        RECT -182.685 66.675 -182.285 67.875 ;
        RECT -180.445 66.675 -180.045 67.875 ;
        RECT -178.205 66.675 -177.805 67.875 ;
        RECT -175.965 66.675 -175.565 67.875 ;
        RECT -173.725 66.675 -173.325 67.875 ;
        RECT -171.485 66.675 -171.085 67.875 ;
        RECT -169.245 66.675 -168.845 67.875 ;
        RECT -167.005 66.675 -166.605 67.875 ;
        RECT -164.765 66.675 -164.365 67.875 ;
        RECT -162.525 66.675 -162.125 67.875 ;
        RECT -160.285 66.675 -159.885 67.875 ;
        RECT -158.045 66.675 -157.645 67.875 ;
        RECT -155.805 66.675 -155.405 67.875 ;
        RECT -153.565 66.675 -153.165 67.875 ;
        RECT -151.325 66.675 -150.925 67.875 ;
        RECT -149.085 66.675 -148.685 67.875 ;
        RECT -146.845 66.675 -146.445 67.875 ;
        RECT -144.605 66.675 -144.205 67.875 ;
        RECT -142.365 66.675 -141.965 67.875 ;
        RECT -140.125 66.675 -139.725 67.875 ;
        RECT -137.885 66.675 -137.485 67.875 ;
        RECT -135.645 66.675 -135.245 67.875 ;
        RECT -133.405 66.675 -133.005 67.875 ;
        RECT -131.165 66.675 -130.765 67.875 ;
        RECT -128.925 66.675 -128.525 67.875 ;
        RECT -126.685 66.675 -126.285 67.875 ;
        RECT -124.445 66.675 -124.045 67.875 ;
        RECT -122.205 66.675 -121.805 67.875 ;
        RECT -119.965 66.675 -119.565 67.875 ;
        RECT -117.725 66.675 -117.325 67.875 ;
        RECT -115.485 66.675 -115.085 67.875 ;
        RECT -113.245 66.675 -112.845 67.875 ;
        RECT -111.005 66.675 -110.605 67.875 ;
        RECT -108.765 66.675 -108.365 67.875 ;
        RECT -106.525 66.675 -106.125 67.875 ;
        RECT -104.285 66.675 -103.885 67.875 ;
        RECT -102.045 66.675 -101.645 67.875 ;
        RECT -99.805 66.675 -99.405 67.875 ;
        RECT -97.565 66.675 -97.165 67.875 ;
        RECT -95.325 66.675 -94.925 67.875 ;
        RECT -93.085 66.675 -92.685 67.875 ;
        RECT -90.845 66.675 -90.445 67.875 ;
        RECT -88.605 66.675 -88.205 67.875 ;
        RECT -86.365 66.675 -85.965 67.875 ;
        RECT -84.125 66.675 -83.725 67.875 ;
        RECT -81.885 66.675 -81.485 67.875 ;
        RECT -79.645 66.675 -79.245 67.875 ;
        RECT -77.405 66.675 -77.005 67.875 ;
        RECT -75.165 66.675 -74.765 67.875 ;
        RECT -72.925 66.675 -72.525 67.875 ;
        RECT -70.685 66.675 -70.285 67.875 ;
        RECT -68.445 66.675 -68.045 67.875 ;
        RECT -66.205 66.675 -65.805 67.875 ;
        RECT -63.965 66.675 -63.565 67.875 ;
        RECT -61.725 66.675 -61.325 67.875 ;
        RECT -59.485 66.675 -59.085 67.875 ;
        RECT -57.245 66.675 -56.845 67.875 ;
        RECT -55.005 66.675 -54.605 67.875 ;
        RECT -52.765 66.675 -52.365 67.875 ;
        RECT -50.525 66.675 -50.125 67.875 ;
        RECT -48.285 66.675 -47.885 67.875 ;
        RECT -46.045 66.675 -45.645 67.875 ;
        RECT -43.805 66.675 -43.405 67.875 ;
        RECT -41.565 66.675 -41.165 67.875 ;
        RECT -39.325 66.675 -38.925 67.875 ;
        RECT -37.085 66.675 -36.685 67.875 ;
        RECT -34.845 66.675 -34.445 67.875 ;
        RECT -32.605 66.675 -32.205 67.875 ;
        RECT -30.365 66.675 -29.965 67.875 ;
        RECT -28.125 66.675 -27.725 67.875 ;
        RECT -25.885 66.675 -25.485 67.875 ;
        RECT -23.645 66.675 -23.245 67.875 ;
        RECT -21.405 66.675 -21.005 67.875 ;
        RECT -19.165 66.675 -18.765 67.875 ;
        RECT -16.925 66.675 -16.525 67.875 ;
        RECT -14.685 66.675 -14.285 67.875 ;
        RECT -12.445 66.675 -12.045 67.875 ;
        RECT -10.205 66.675 -9.805 67.875 ;
        RECT -7.965 66.675 -7.565 67.875 ;
        RECT -5.725 66.675 -5.325 67.875 ;
        RECT -3.485 66.675 -3.085 67.875 ;
        RECT -1.245 66.675 -0.845 67.875 ;
        RECT 0.995 66.675 1.395 67.875 ;
        RECT 3.235 66.675 3.635 67.875 ;
        RECT 5.475 66.675 5.875 67.875 ;
        RECT 7.715 66.675 8.115 67.875 ;
        RECT 9.955 66.675 10.355 67.875 ;
        RECT 12.195 66.675 12.595 67.875 ;
        RECT 14.435 66.675 14.835 67.875 ;
        RECT 16.675 66.675 17.075 67.875 ;
        RECT 18.915 66.675 19.315 67.875 ;
        RECT 21.155 66.675 21.555 67.875 ;
        RECT 23.395 66.675 23.795 67.875 ;
        RECT 25.635 66.675 26.035 67.875 ;
        RECT 27.875 66.675 28.275 67.875 ;
        RECT 30.115 66.675 30.515 67.875 ;
        RECT 32.355 66.675 32.755 67.875 ;
        RECT 34.595 66.675 34.995 67.875 ;
        RECT 36.835 66.675 37.235 67.875 ;
        RECT 39.075 66.675 39.475 67.875 ;
        RECT 41.315 66.675 41.715 67.875 ;
        RECT 43.555 66.675 43.955 67.875 ;
        RECT 45.795 66.675 46.195 67.875 ;
        RECT 48.035 66.675 48.435 67.875 ;
        RECT 50.275 66.675 50.675 67.875 ;
        RECT 52.515 66.675 52.915 67.875 ;
        RECT 54.755 66.675 55.155 67.875 ;
        RECT 56.995 66.675 57.395 67.875 ;
        RECT 59.235 66.675 59.635 67.875 ;
        RECT 61.475 66.675 61.875 67.875 ;
        RECT 63.715 66.675 64.115 67.875 ;
        RECT 65.955 66.675 66.355 67.875 ;
        RECT 68.195 66.675 68.595 67.875 ;
        RECT 70.435 66.675 70.835 67.875 ;
        RECT 72.675 66.675 73.075 67.875 ;
        RECT 74.915 66.675 75.315 67.875 ;
        RECT 77.155 66.675 77.555 67.875 ;
        RECT 79.395 66.675 79.795 67.875 ;
        RECT 81.635 66.675 82.035 67.875 ;
        RECT 83.875 66.675 84.275 67.875 ;
        RECT 86.115 66.675 86.515 67.875 ;
        RECT 88.355 66.675 88.755 67.875 ;
        RECT 90.595 66.675 90.995 67.875 ;
        RECT 92.835 66.675 93.235 67.875 ;
        RECT 95.075 66.675 95.475 67.875 ;
        RECT 97.315 66.675 97.715 67.875 ;
        RECT 101.155 67.075 102.355 67.475 ;
        RECT -475.005 43.815 -474.605 45.015 ;
        RECT -472.765 43.815 -472.365 45.015 ;
        RECT -470.525 43.815 -470.125 45.015 ;
        RECT -468.285 43.815 -467.885 45.015 ;
        RECT -466.045 43.815 -465.645 45.015 ;
        RECT -463.805 43.815 -463.405 45.015 ;
        RECT -461.565 43.815 -461.165 45.015 ;
        RECT -459.325 43.815 -458.925 45.015 ;
        RECT -457.085 43.815 -456.685 45.015 ;
        RECT -454.845 43.815 -454.445 45.015 ;
        RECT -452.605 43.815 -452.205 45.015 ;
        RECT -450.365 43.815 -449.965 45.015 ;
        RECT -448.125 43.815 -447.725 45.015 ;
        RECT -445.885 43.815 -445.485 45.015 ;
        RECT -443.645 43.815 -443.245 45.015 ;
        RECT -441.405 43.815 -441.005 45.015 ;
        RECT -439.165 43.815 -438.765 45.015 ;
        RECT -436.925 43.815 -436.525 45.015 ;
        RECT -434.685 43.815 -434.285 45.015 ;
        RECT -432.445 43.815 -432.045 45.015 ;
        RECT -430.205 43.815 -429.805 45.015 ;
        RECT -427.965 43.815 -427.565 45.015 ;
        RECT -425.725 43.815 -425.325 45.015 ;
        RECT -423.485 43.815 -423.085 45.015 ;
        RECT -421.245 43.815 -420.845 45.015 ;
        RECT -419.005 43.815 -418.605 45.015 ;
        RECT -416.765 43.815 -416.365 45.015 ;
        RECT -414.525 43.815 -414.125 45.015 ;
        RECT -412.285 43.815 -411.885 45.015 ;
        RECT -410.045 43.815 -409.645 45.015 ;
        RECT -407.805 43.815 -407.405 45.015 ;
        RECT -405.565 43.815 -405.165 45.015 ;
        RECT -403.325 43.815 -402.925 45.015 ;
        RECT -401.085 43.815 -400.685 45.015 ;
        RECT -398.845 43.815 -398.445 45.015 ;
        RECT -396.605 43.815 -396.205 45.015 ;
        RECT -394.365 43.815 -393.965 45.015 ;
        RECT -392.125 43.815 -391.725 45.015 ;
        RECT -389.885 43.815 -389.485 45.015 ;
        RECT -387.645 43.815 -387.245 45.015 ;
        RECT -385.405 43.815 -385.005 45.015 ;
        RECT -383.165 43.815 -382.765 45.015 ;
        RECT -380.925 43.815 -380.525 45.015 ;
        RECT -378.685 43.815 -378.285 45.015 ;
        RECT -376.445 43.815 -376.045 45.015 ;
        RECT -374.205 43.815 -373.805 45.015 ;
        RECT -371.965 43.815 -371.565 45.015 ;
        RECT -369.725 43.815 -369.325 45.015 ;
        RECT -367.485 43.815 -367.085 45.015 ;
        RECT -365.245 43.815 -364.845 45.015 ;
        RECT -363.005 43.815 -362.605 45.015 ;
        RECT -360.765 43.815 -360.365 45.015 ;
        RECT -358.525 43.815 -358.125 45.015 ;
        RECT -356.285 43.815 -355.885 45.015 ;
        RECT -354.045 43.815 -353.645 45.015 ;
        RECT -351.805 43.815 -351.405 45.015 ;
        RECT -349.565 43.815 -349.165 45.015 ;
        RECT -347.325 43.815 -346.925 45.015 ;
        RECT -345.085 43.815 -344.685 45.015 ;
        RECT -342.845 43.815 -342.445 45.015 ;
        RECT -340.605 43.815 -340.205 45.015 ;
        RECT -338.365 43.815 -337.965 45.015 ;
        RECT -336.125 43.815 -335.725 45.015 ;
        RECT -333.885 43.815 -333.485 45.015 ;
        RECT -331.645 43.815 -331.245 45.015 ;
        RECT -329.405 43.815 -329.005 45.015 ;
        RECT -327.165 43.815 -326.765 45.015 ;
        RECT -324.925 43.815 -324.525 45.015 ;
        RECT -322.685 43.815 -322.285 45.015 ;
        RECT -320.445 43.815 -320.045 45.015 ;
        RECT -318.205 43.815 -317.805 45.015 ;
        RECT -315.965 43.815 -315.565 45.015 ;
        RECT -313.725 43.815 -313.325 45.015 ;
        RECT -311.485 43.815 -311.085 45.015 ;
        RECT -309.245 43.815 -308.845 45.015 ;
        RECT -307.005 43.815 -306.605 45.015 ;
        RECT -304.765 43.815 -304.365 45.015 ;
        RECT -302.525 43.815 -302.125 45.015 ;
        RECT -300.285 43.815 -299.885 45.015 ;
        RECT -298.045 43.815 -297.645 45.015 ;
        RECT -295.805 43.815 -295.405 45.015 ;
        RECT -293.565 43.815 -293.165 45.015 ;
        RECT -291.325 43.815 -290.925 45.015 ;
        RECT -289.085 43.815 -288.685 45.015 ;
        RECT -286.845 43.815 -286.445 45.015 ;
        RECT -284.605 43.815 -284.205 45.015 ;
        RECT -282.365 43.815 -281.965 45.015 ;
        RECT -280.125 43.815 -279.725 45.015 ;
        RECT -277.885 43.815 -277.485 45.015 ;
        RECT -275.645 43.815 -275.245 45.015 ;
        RECT -273.405 43.815 -273.005 45.015 ;
        RECT -271.165 43.815 -270.765 45.015 ;
        RECT -268.925 43.815 -268.525 45.015 ;
        RECT -266.685 43.815 -266.285 45.015 ;
        RECT -264.445 43.815 -264.045 45.015 ;
        RECT -262.205 43.815 -261.805 45.015 ;
        RECT -259.965 43.815 -259.565 45.015 ;
        RECT -257.725 43.815 -257.325 45.015 ;
        RECT -255.485 43.815 -255.085 45.015 ;
        RECT -253.245 43.815 -252.845 45.015 ;
        RECT -251.005 43.815 -250.605 45.015 ;
        RECT -248.765 43.815 -248.365 45.015 ;
        RECT -246.525 43.815 -246.125 45.015 ;
        RECT -244.285 43.815 -243.885 45.015 ;
        RECT -242.045 43.815 -241.645 45.015 ;
        RECT -239.805 43.815 -239.405 45.015 ;
        RECT -237.565 43.815 -237.165 45.015 ;
        RECT -235.325 43.815 -234.925 45.015 ;
        RECT -233.085 43.815 -232.685 45.015 ;
        RECT -230.845 43.815 -230.445 45.015 ;
        RECT -228.605 43.815 -228.205 45.015 ;
        RECT -226.365 43.815 -225.965 45.015 ;
        RECT -224.125 43.815 -223.725 45.015 ;
        RECT -221.885 43.815 -221.485 45.015 ;
        RECT -219.645 43.815 -219.245 45.015 ;
        RECT -217.405 43.815 -217.005 45.015 ;
        RECT -215.165 43.815 -214.765 45.015 ;
        RECT -212.925 43.815 -212.525 45.015 ;
        RECT -210.685 43.815 -210.285 45.015 ;
        RECT -208.445 43.815 -208.045 45.015 ;
        RECT -206.205 43.815 -205.805 45.015 ;
        RECT -203.965 43.815 -203.565 45.015 ;
        RECT -201.725 43.815 -201.325 45.015 ;
        RECT -199.485 43.815 -199.085 45.015 ;
        RECT -197.245 43.815 -196.845 45.015 ;
        RECT -195.005 43.815 -194.605 45.015 ;
        RECT -192.765 43.815 -192.365 45.015 ;
        RECT -190.525 43.815 -190.125 45.015 ;
        RECT -187.165 43.815 -186.765 45.015 ;
        RECT -184.925 43.815 -184.525 45.015 ;
        RECT -182.685 43.815 -182.285 45.015 ;
        RECT -180.445 43.815 -180.045 45.015 ;
        RECT -178.205 43.815 -177.805 45.015 ;
        RECT -175.965 43.815 -175.565 45.015 ;
        RECT -173.725 43.815 -173.325 45.015 ;
        RECT -171.485 43.815 -171.085 45.015 ;
        RECT -169.245 43.815 -168.845 45.015 ;
        RECT -167.005 43.815 -166.605 45.015 ;
        RECT -164.765 43.815 -164.365 45.015 ;
        RECT -162.525 43.815 -162.125 45.015 ;
        RECT -160.285 43.815 -159.885 45.015 ;
        RECT -158.045 43.815 -157.645 45.015 ;
        RECT -155.805 43.815 -155.405 45.015 ;
        RECT -153.565 43.815 -153.165 45.015 ;
        RECT -151.325 43.815 -150.925 45.015 ;
        RECT -149.085 43.815 -148.685 45.015 ;
        RECT -146.845 43.815 -146.445 45.015 ;
        RECT -144.605 43.815 -144.205 45.015 ;
        RECT -142.365 43.815 -141.965 45.015 ;
        RECT -140.125 43.815 -139.725 45.015 ;
        RECT -137.885 43.815 -137.485 45.015 ;
        RECT -135.645 43.815 -135.245 45.015 ;
        RECT -133.405 43.815 -133.005 45.015 ;
        RECT -131.165 43.815 -130.765 45.015 ;
        RECT -128.925 43.815 -128.525 45.015 ;
        RECT -126.685 43.815 -126.285 45.015 ;
        RECT -124.445 43.815 -124.045 45.015 ;
        RECT -122.205 43.815 -121.805 45.015 ;
        RECT -119.965 43.815 -119.565 45.015 ;
        RECT -117.725 43.815 -117.325 45.015 ;
        RECT -115.485 43.815 -115.085 45.015 ;
        RECT -113.245 43.815 -112.845 45.015 ;
        RECT -111.005 43.815 -110.605 45.015 ;
        RECT -108.765 43.815 -108.365 45.015 ;
        RECT -106.525 43.815 -106.125 45.015 ;
        RECT -104.285 43.815 -103.885 45.015 ;
        RECT -102.045 43.815 -101.645 45.015 ;
        RECT -99.805 43.815 -99.405 45.015 ;
        RECT -97.565 43.815 -97.165 45.015 ;
        RECT -95.325 43.815 -94.925 45.015 ;
        RECT -93.085 43.815 -92.685 45.015 ;
        RECT -90.845 43.815 -90.445 45.015 ;
        RECT -88.605 43.815 -88.205 45.015 ;
        RECT -86.365 43.815 -85.965 45.015 ;
        RECT -84.125 43.815 -83.725 45.015 ;
        RECT -81.885 43.815 -81.485 45.015 ;
        RECT -79.645 43.815 -79.245 45.015 ;
        RECT -77.405 43.815 -77.005 45.015 ;
        RECT -75.165 43.815 -74.765 45.015 ;
        RECT -72.925 43.815 -72.525 45.015 ;
        RECT -70.685 43.815 -70.285 45.015 ;
        RECT -68.445 43.815 -68.045 45.015 ;
        RECT -66.205 43.815 -65.805 45.015 ;
        RECT -63.965 43.815 -63.565 45.015 ;
        RECT -61.725 43.815 -61.325 45.015 ;
        RECT -59.485 43.815 -59.085 45.015 ;
        RECT -57.245 43.815 -56.845 45.015 ;
        RECT -55.005 43.815 -54.605 45.015 ;
        RECT -52.765 43.815 -52.365 45.015 ;
        RECT -50.525 43.815 -50.125 45.015 ;
        RECT -48.285 43.815 -47.885 45.015 ;
        RECT -46.045 43.815 -45.645 45.015 ;
        RECT -43.805 43.815 -43.405 45.015 ;
        RECT -41.565 43.815 -41.165 45.015 ;
        RECT -39.325 43.815 -38.925 45.015 ;
        RECT -37.085 43.815 -36.685 45.015 ;
        RECT -34.845 43.815 -34.445 45.015 ;
        RECT -32.605 43.815 -32.205 45.015 ;
        RECT -30.365 43.815 -29.965 45.015 ;
        RECT -28.125 43.815 -27.725 45.015 ;
        RECT -25.885 43.815 -25.485 45.015 ;
        RECT -23.645 43.815 -23.245 45.015 ;
        RECT -21.405 43.815 -21.005 45.015 ;
        RECT -19.165 43.815 -18.765 45.015 ;
        RECT -16.925 43.815 -16.525 45.015 ;
        RECT -14.685 43.815 -14.285 45.015 ;
        RECT -12.445 43.815 -12.045 45.015 ;
        RECT -10.205 43.815 -9.805 45.015 ;
        RECT -7.965 43.815 -7.565 45.015 ;
        RECT -5.725 43.815 -5.325 45.015 ;
        RECT -3.485 43.815 -3.085 45.015 ;
        RECT -1.245 43.815 -0.845 45.015 ;
        RECT 0.995 43.815 1.395 45.015 ;
        RECT 3.235 43.815 3.635 45.015 ;
        RECT 5.475 43.815 5.875 45.015 ;
        RECT 7.715 43.815 8.115 45.015 ;
        RECT 9.955 43.815 10.355 45.015 ;
        RECT 12.195 43.815 12.595 45.015 ;
        RECT 14.435 43.815 14.835 45.015 ;
        RECT 16.675 43.815 17.075 45.015 ;
        RECT 18.915 43.815 19.315 45.015 ;
        RECT 21.155 43.815 21.555 45.015 ;
        RECT 23.395 43.815 23.795 45.015 ;
        RECT 25.635 43.815 26.035 45.015 ;
        RECT 27.875 43.815 28.275 45.015 ;
        RECT 30.115 43.815 30.515 45.015 ;
        RECT 32.355 43.815 32.755 45.015 ;
        RECT 34.595 43.815 34.995 45.015 ;
        RECT 36.835 43.815 37.235 45.015 ;
        RECT 39.075 43.815 39.475 45.015 ;
        RECT 41.315 43.815 41.715 45.015 ;
        RECT 43.555 43.815 43.955 45.015 ;
        RECT 45.795 43.815 46.195 45.015 ;
        RECT 48.035 43.815 48.435 45.015 ;
        RECT 50.275 43.815 50.675 45.015 ;
        RECT 52.515 43.815 52.915 45.015 ;
        RECT 54.755 43.815 55.155 45.015 ;
        RECT 56.995 43.815 57.395 45.015 ;
        RECT 59.235 43.815 59.635 45.015 ;
        RECT 61.475 43.815 61.875 45.015 ;
        RECT 63.715 43.815 64.115 45.015 ;
        RECT 65.955 43.815 66.355 45.015 ;
        RECT 68.195 43.815 68.595 45.015 ;
        RECT 70.435 43.815 70.835 45.015 ;
        RECT 72.675 43.815 73.075 45.015 ;
        RECT 74.915 43.815 75.315 45.015 ;
        RECT 77.155 43.815 77.555 45.015 ;
        RECT 79.395 43.815 79.795 45.015 ;
        RECT 81.635 43.815 82.035 45.015 ;
        RECT 83.875 43.815 84.275 45.015 ;
        RECT 86.115 43.815 86.515 45.015 ;
        RECT 88.355 43.815 88.755 45.015 ;
        RECT 90.595 43.815 90.995 45.015 ;
        RECT 92.835 43.815 93.235 45.015 ;
        RECT 95.075 43.815 95.475 45.015 ;
        RECT 97.315 43.815 97.715 45.015 ;
        RECT 101.505 44.615 102.005 67.075 ;
        RECT 101.155 44.215 102.355 44.615 ;
        RECT -473.885 40.455 -473.485 41.655 ;
        RECT -469.405 40.455 -469.005 41.655 ;
        RECT -464.925 40.455 -464.525 41.655 ;
        RECT -460.445 40.455 -460.045 41.655 ;
        RECT -455.965 40.455 -455.565 41.655 ;
        RECT -451.485 40.455 -451.085 41.655 ;
        RECT -447.005 40.455 -446.605 41.655 ;
        RECT -442.525 40.455 -442.125 41.655 ;
        RECT -438.045 40.455 -437.645 41.655 ;
        RECT -433.565 40.455 -433.165 41.655 ;
        RECT -429.085 40.455 -428.685 41.655 ;
        RECT -424.605 40.455 -424.205 41.655 ;
        RECT -420.125 40.455 -419.725 41.655 ;
        RECT -415.645 40.455 -415.245 41.655 ;
        RECT -411.165 40.455 -410.765 41.655 ;
        RECT -406.685 40.455 -406.285 41.655 ;
        RECT -402.205 40.455 -401.805 41.655 ;
        RECT -397.725 40.455 -397.325 41.655 ;
        RECT -393.245 40.455 -392.845 41.655 ;
        RECT -388.765 40.455 -388.365 41.655 ;
        RECT -384.285 40.455 -383.885 41.655 ;
        RECT -379.805 40.455 -379.405 41.655 ;
        RECT -375.325 40.455 -374.925 41.655 ;
        RECT -370.845 40.455 -370.445 41.655 ;
        RECT -366.365 40.455 -365.965 41.655 ;
        RECT -361.885 40.455 -361.485 41.655 ;
        RECT -357.405 40.455 -357.005 41.655 ;
        RECT -352.925 40.455 -352.525 41.655 ;
        RECT -348.445 40.455 -348.045 41.655 ;
        RECT -343.965 40.455 -343.565 41.655 ;
        RECT -339.485 40.455 -339.085 41.655 ;
        RECT -335.005 40.455 -334.605 41.655 ;
        RECT -330.525 40.455 -330.125 41.655 ;
        RECT -326.045 40.455 -325.645 41.655 ;
        RECT -321.565 40.455 -321.165 41.655 ;
        RECT -317.085 40.455 -316.685 41.655 ;
        RECT -312.605 40.455 -312.205 41.655 ;
        RECT -308.125 40.455 -307.725 41.655 ;
        RECT -303.645 40.455 -303.245 41.655 ;
        RECT -299.165 40.455 -298.765 41.655 ;
        RECT -294.685 40.455 -294.285 41.655 ;
        RECT -290.205 40.455 -289.805 41.655 ;
        RECT -285.725 40.455 -285.325 41.655 ;
        RECT -281.245 40.455 -280.845 41.655 ;
        RECT -276.765 40.455 -276.365 41.655 ;
        RECT -272.285 40.455 -271.885 41.655 ;
        RECT -267.805 40.455 -267.405 41.655 ;
        RECT -263.325 40.455 -262.925 41.655 ;
        RECT -258.845 40.455 -258.445 41.655 ;
        RECT -254.365 40.455 -253.965 41.655 ;
        RECT -249.885 40.455 -249.485 41.655 ;
        RECT -245.405 40.455 -245.005 41.655 ;
        RECT -240.925 40.455 -240.525 41.655 ;
        RECT -236.445 40.455 -236.045 41.655 ;
        RECT -231.965 40.455 -231.565 41.655 ;
        RECT -227.485 40.455 -227.085 41.655 ;
        RECT -223.005 40.455 -222.605 41.655 ;
        RECT -218.525 40.455 -218.125 41.655 ;
        RECT -214.045 40.455 -213.645 41.655 ;
        RECT -209.565 40.455 -209.165 41.655 ;
        RECT -205.085 40.455 -204.685 41.655 ;
        RECT -200.605 40.455 -200.205 41.655 ;
        RECT -196.125 40.455 -195.725 41.655 ;
        RECT -191.645 40.455 -191.245 41.655 ;
        RECT -186.045 40.455 -185.645 41.655 ;
        RECT -181.565 40.455 -181.165 41.655 ;
        RECT -177.085 40.455 -176.685 41.655 ;
        RECT -172.605 40.455 -172.205 41.655 ;
        RECT -168.125 40.455 -167.725 41.655 ;
        RECT -163.645 40.455 -163.245 41.655 ;
        RECT -159.165 40.455 -158.765 41.655 ;
        RECT -154.685 40.455 -154.285 41.655 ;
        RECT -150.205 40.455 -149.805 41.655 ;
        RECT -145.725 40.455 -145.325 41.655 ;
        RECT -141.245 40.455 -140.845 41.655 ;
        RECT -136.765 40.455 -136.365 41.655 ;
        RECT -132.285 40.455 -131.885 41.655 ;
        RECT -127.805 40.455 -127.405 41.655 ;
        RECT -123.325 40.455 -122.925 41.655 ;
        RECT -118.845 40.455 -118.445 41.655 ;
        RECT -114.365 40.455 -113.965 41.655 ;
        RECT -109.885 40.455 -109.485 41.655 ;
        RECT -105.405 40.455 -105.005 41.655 ;
        RECT -100.925 40.455 -100.525 41.655 ;
        RECT -96.445 40.455 -96.045 41.655 ;
        RECT -91.965 40.455 -91.565 41.655 ;
        RECT -87.485 40.455 -87.085 41.655 ;
        RECT -83.005 40.455 -82.605 41.655 ;
        RECT -78.525 40.455 -78.125 41.655 ;
        RECT -74.045 40.455 -73.645 41.655 ;
        RECT -69.565 40.455 -69.165 41.655 ;
        RECT -65.085 40.455 -64.685 41.655 ;
        RECT -60.605 40.455 -60.205 41.655 ;
        RECT -56.125 40.455 -55.725 41.655 ;
        RECT -51.645 40.455 -51.245 41.655 ;
        RECT -47.165 40.455 -46.765 41.655 ;
        RECT -42.685 40.455 -42.285 41.655 ;
        RECT -38.205 40.455 -37.805 41.655 ;
        RECT -33.725 40.455 -33.325 41.655 ;
        RECT -29.245 40.455 -28.845 41.655 ;
        RECT -24.765 40.455 -24.365 41.655 ;
        RECT -20.285 40.455 -19.885 41.655 ;
        RECT -15.805 40.455 -15.405 41.655 ;
        RECT -11.325 40.455 -10.925 41.655 ;
        RECT -6.845 40.455 -6.445 41.655 ;
        RECT -2.365 40.455 -1.965 41.655 ;
        RECT 2.115 40.455 2.515 41.655 ;
        RECT 6.595 40.455 6.995 41.655 ;
        RECT 11.075 40.455 11.475 41.655 ;
        RECT 15.555 40.455 15.955 41.655 ;
        RECT 20.035 40.455 20.435 41.655 ;
        RECT 24.515 40.455 24.915 41.655 ;
        RECT 28.995 40.455 29.395 41.655 ;
        RECT 33.475 40.455 33.875 41.655 ;
        RECT 37.955 40.455 38.355 41.655 ;
        RECT 42.435 40.455 42.835 41.655 ;
        RECT 46.915 40.455 47.315 41.655 ;
        RECT 51.395 40.455 51.795 41.655 ;
        RECT 55.875 40.455 56.275 41.655 ;
        RECT 60.355 40.455 60.755 41.655 ;
        RECT 64.835 40.455 65.235 41.655 ;
        RECT 69.315 40.455 69.715 41.655 ;
        RECT 73.795 40.455 74.195 41.655 ;
        RECT 78.275 40.455 78.675 41.655 ;
        RECT 82.755 40.455 83.155 41.655 ;
        RECT 87.235 40.455 87.635 41.655 ;
        RECT 91.715 40.455 92.115 41.655 ;
        RECT 96.195 40.455 96.595 41.655 ;
        RECT 103.305 41.255 103.805 70.435 ;
        RECT 102.955 40.855 104.155 41.255 ;
        RECT -471.645 37.095 -471.245 38.295 ;
        RECT -462.685 37.095 -462.285 38.295 ;
        RECT -453.725 37.095 -453.325 38.295 ;
        RECT -444.765 37.095 -444.365 38.295 ;
        RECT -435.805 37.095 -435.405 38.295 ;
        RECT -426.845 37.095 -426.445 38.295 ;
        RECT -417.885 37.095 -417.485 38.295 ;
        RECT -408.925 37.095 -408.525 38.295 ;
        RECT -399.965 37.095 -399.565 38.295 ;
        RECT -391.005 37.095 -390.605 38.295 ;
        RECT -382.045 37.095 -381.645 38.295 ;
        RECT -373.085 37.095 -372.685 38.295 ;
        RECT -364.125 37.095 -363.725 38.295 ;
        RECT -355.165 37.095 -354.765 38.295 ;
        RECT -346.205 37.095 -345.805 38.295 ;
        RECT -337.245 37.095 -336.845 38.295 ;
        RECT -328.285 37.095 -327.885 38.295 ;
        RECT -319.325 37.095 -318.925 38.295 ;
        RECT -310.365 37.095 -309.965 38.295 ;
        RECT -301.405 37.095 -301.005 38.295 ;
        RECT -292.445 37.095 -292.045 38.295 ;
        RECT -283.485 37.095 -283.085 38.295 ;
        RECT -274.525 37.095 -274.125 38.295 ;
        RECT -265.565 37.095 -265.165 38.295 ;
        RECT -256.605 37.095 -256.205 38.295 ;
        RECT -247.645 37.095 -247.245 38.295 ;
        RECT -238.685 37.095 -238.285 38.295 ;
        RECT -229.725 37.095 -229.325 38.295 ;
        RECT -220.765 37.095 -220.365 38.295 ;
        RECT -211.805 37.095 -211.405 38.295 ;
        RECT -202.845 37.095 -202.445 38.295 ;
        RECT -193.885 37.095 -193.485 38.295 ;
        RECT -183.805 37.095 -183.405 38.295 ;
        RECT -174.845 37.095 -174.445 38.295 ;
        RECT -165.885 37.095 -165.485 38.295 ;
        RECT -156.925 37.095 -156.525 38.295 ;
        RECT -147.965 37.095 -147.565 38.295 ;
        RECT -139.005 37.095 -138.605 38.295 ;
        RECT -130.045 37.095 -129.645 38.295 ;
        RECT -121.085 37.095 -120.685 38.295 ;
        RECT -112.125 37.095 -111.725 38.295 ;
        RECT -103.165 37.095 -102.765 38.295 ;
        RECT -94.205 37.095 -93.805 38.295 ;
        RECT -85.245 37.095 -84.845 38.295 ;
        RECT -76.285 37.095 -75.885 38.295 ;
        RECT -67.325 37.095 -66.925 38.295 ;
        RECT -58.365 37.095 -57.965 38.295 ;
        RECT -49.405 37.095 -49.005 38.295 ;
        RECT -40.445 37.095 -40.045 38.295 ;
        RECT -31.485 37.095 -31.085 38.295 ;
        RECT -22.525 37.095 -22.125 38.295 ;
        RECT -13.565 37.095 -13.165 38.295 ;
        RECT -4.605 37.095 -4.205 38.295 ;
        RECT 4.355 37.095 4.755 38.295 ;
        RECT 13.315 37.095 13.715 38.295 ;
        RECT 22.275 37.095 22.675 38.295 ;
        RECT 31.235 37.095 31.635 38.295 ;
        RECT 40.195 37.095 40.595 38.295 ;
        RECT 49.155 37.095 49.555 38.295 ;
        RECT 58.115 37.095 58.515 38.295 ;
        RECT 67.075 37.095 67.475 38.295 ;
        RECT 76.035 37.095 76.435 38.295 ;
        RECT 84.995 37.095 85.395 38.295 ;
        RECT 93.955 37.095 94.355 38.295 ;
        RECT 105.105 37.895 105.605 73.795 ;
        RECT 104.755 37.495 105.955 37.895 ;
        RECT -467.165 33.735 -466.765 34.935 ;
        RECT -449.245 33.735 -448.845 34.935 ;
        RECT -431.325 33.735 -430.925 34.935 ;
        RECT -413.405 33.735 -413.005 34.935 ;
        RECT -395.485 33.735 -395.085 34.935 ;
        RECT -377.565 33.735 -377.165 34.935 ;
        RECT -359.645 33.735 -359.245 34.935 ;
        RECT -341.725 33.735 -341.325 34.935 ;
        RECT -323.805 33.735 -323.405 34.935 ;
        RECT -305.885 33.735 -305.485 34.935 ;
        RECT -287.965 33.735 -287.565 34.935 ;
        RECT -270.045 33.735 -269.645 34.935 ;
        RECT -252.125 33.735 -251.725 34.935 ;
        RECT -234.205 33.735 -233.805 34.935 ;
        RECT -216.285 33.735 -215.885 34.935 ;
        RECT -198.365 33.735 -197.965 34.935 ;
        RECT -179.325 33.735 -178.925 34.935 ;
        RECT -161.405 33.735 -161.005 34.935 ;
        RECT -143.485 33.735 -143.085 34.935 ;
        RECT -125.565 33.735 -125.165 34.935 ;
        RECT -107.645 33.735 -107.245 34.935 ;
        RECT -89.725 33.735 -89.325 34.935 ;
        RECT -71.805 33.735 -71.405 34.935 ;
        RECT -53.885 33.735 -53.485 34.935 ;
        RECT -35.965 33.735 -35.565 34.935 ;
        RECT -18.045 33.735 -17.645 34.935 ;
        RECT -0.125 33.735 0.275 34.935 ;
        RECT 17.795 33.735 18.195 34.935 ;
        RECT 35.715 33.735 36.115 34.935 ;
        RECT 53.635 33.735 54.035 34.935 ;
        RECT 71.555 33.735 71.955 34.935 ;
        RECT 89.475 33.735 89.875 34.935 ;
        RECT 106.905 34.535 107.405 77.155 ;
        RECT 106.555 34.135 107.755 34.535 ;
        RECT -458.205 30.375 -457.805 31.575 ;
        RECT -422.365 30.375 -421.965 31.575 ;
        RECT -386.525 30.375 -386.125 31.575 ;
        RECT -350.685 30.375 -350.285 31.575 ;
        RECT -314.845 30.375 -314.445 31.575 ;
        RECT -279.005 30.375 -278.605 31.575 ;
        RECT -243.165 30.375 -242.765 31.575 ;
        RECT -207.325 30.375 -206.925 31.575 ;
        RECT -170.365 30.375 -169.965 31.575 ;
        RECT -134.525 30.375 -134.125 31.575 ;
        RECT -98.685 30.375 -98.285 31.575 ;
        RECT -62.845 30.375 -62.445 31.575 ;
        RECT -27.005 30.375 -26.605 31.575 ;
        RECT 8.835 30.375 9.235 31.575 ;
        RECT 44.675 30.375 45.075 31.575 ;
        RECT 80.515 30.375 80.915 31.575 ;
        RECT 108.705 31.175 109.205 80.515 ;
        RECT 108.355 30.775 109.555 31.175 ;
        RECT -440.285 27.015 -439.885 28.215 ;
        RECT -368.605 27.015 -368.205 28.215 ;
        RECT -296.925 27.015 -296.525 28.215 ;
        RECT -225.245 27.015 -224.845 28.215 ;
        RECT -152.445 27.015 -152.045 28.215 ;
        RECT -80.765 27.015 -80.365 28.215 ;
        RECT -9.085 27.015 -8.685 28.215 ;
        RECT 62.595 27.015 62.995 28.215 ;
        RECT 110.505 27.815 111.005 83.875 ;
        RECT 110.155 27.415 111.355 27.815 ;
        RECT -404.445 23.655 -404.045 24.855 ;
        RECT -261.085 23.655 -260.685 24.855 ;
        RECT -116.605 23.655 -116.205 24.855 ;
        RECT 26.755 23.655 27.155 24.855 ;
        RECT 112.305 24.455 112.805 87.235 ;
        RECT 111.955 24.055 113.155 24.455 ;
        RECT -332.765 20.295 -332.365 21.495 ;
        RECT -44.925 20.295 -44.525 21.495 ;
        RECT 114.105 21.095 114.605 90.595 ;
        RECT 113.755 20.695 114.955 21.095 ;
        RECT -188.285 16.935 -187.885 18.135 ;
        RECT 115.905 17.735 116.405 93.955 ;
        RECT 120.925 93.905 121.925 94.405 ;
        RECT 120.925 90.545 121.925 91.045 ;
        RECT 120.925 87.185 121.925 87.685 ;
        RECT 120.925 83.825 121.925 84.325 ;
        RECT 120.925 80.465 121.925 80.965 ;
        RECT 120.925 77.105 121.925 77.605 ;
        RECT 120.925 73.745 121.925 74.245 ;
        RECT 120.925 70.385 121.925 70.885 ;
        RECT 120.925 67.025 121.925 67.525 ;
        RECT 120.925 63.665 121.925 64.165 ;
        RECT 286.700 55.400 289.200 55.620 ;
        RECT 286.700 55.260 293.200 55.400 ;
        RECT 286.700 54.980 299.750 55.260 ;
        RECT 286.700 54.840 293.200 54.980 ;
        RECT 286.700 54.620 289.200 54.840 ;
        RECT 316.170 52.180 322.710 52.460 ;
        RECT 352.010 47.700 360.230 47.980 ;
        RECT 369.930 47.700 375.350 47.980 ;
        RECT 387.850 47.700 394.390 47.980 ;
        RECT 405.770 47.700 417.350 47.980 ;
        RECT 423.690 47.700 432.470 47.980 ;
        RECT 422.010 46.020 426.870 46.300 ;
        RECT 286.700 45.320 289.200 45.540 ;
        RECT 405.770 45.460 413.430 45.740 ;
        RECT 286.700 45.180 293.200 45.320 ;
        RECT 286.700 44.900 299.190 45.180 ;
        RECT 286.700 44.760 293.200 44.900 ;
        RECT 286.700 44.540 289.200 44.760 ;
        RECT 334.090 43.780 344.550 44.060 ;
        RECT 353.690 43.780 376.470 44.060 ;
        RECT 385.660 43.220 436.390 43.500 ;
        RECT 309.450 42.100 319.910 42.380 ;
        RECT 385.660 41.820 385.940 43.220 ;
        RECT 418.650 42.660 423.510 42.940 ;
        RECT 387.290 42.100 392.150 42.380 ;
        RECT 417.530 42.100 444.790 42.380 ;
        RECT 310.570 41.540 314.870 41.820 ;
        RECT 373.850 41.540 385.990 41.820 ;
        RECT 412.490 41.540 416.790 41.820 ;
        RECT 427.050 41.540 457.670 41.820 ;
        RECT 339.130 39.860 339.510 40.140 ;
        RECT 377.770 39.860 435.270 40.140 ;
        RECT 339.180 39.580 339.460 39.860 ;
        RECT 338.010 39.300 404.980 39.580 ;
        RECT 427.050 39.300 443.110 39.580 ;
        RECT 404.700 39.020 404.980 39.300 ;
        RECT 302.730 38.740 308.710 39.020 ;
        RECT 339.130 38.740 363.590 39.020 ;
        RECT 365.450 38.740 374.230 39.020 ;
        RECT 387.850 38.740 403.860 39.020 ;
        RECT 404.650 38.740 405.030 39.020 ;
        RECT 416.970 38.740 420.150 39.020 ;
        RECT 428.170 38.740 445.910 39.020 ;
        RECT 403.580 38.460 403.860 38.740 ;
        RECT 361.530 38.180 365.270 38.460 ;
        RECT 386.170 38.180 391.030 38.460 ;
        RECT 403.580 38.180 415.670 38.460 ;
        RECT 415.340 36.220 415.620 38.180 ;
        RECT 419.820 37.900 420.100 38.740 ;
        RECT 423.130 38.180 438.070 38.460 ;
        RECT 419.820 37.620 442.550 37.900 ;
        RECT 388.410 35.940 412.870 36.220 ;
        RECT 415.340 35.940 422.340 36.220 ;
        RECT 431.530 35.940 448.710 36.220 ;
        RECT 422.060 35.660 422.340 35.940 ;
        RECT 286.700 35.240 289.200 35.460 ;
        RECT 321.770 35.380 338.390 35.660 ;
        RECT 341.930 35.380 355.750 35.660 ;
        RECT 356.490 35.380 378.150 35.660 ;
        RECT 421.870 35.380 434.150 35.660 ;
        RECT 286.700 35.100 293.200 35.240 ;
        RECT 355.420 35.100 355.700 35.380 ;
        RECT 286.700 34.820 299.190 35.100 ;
        RECT 341.370 34.820 343.990 35.100 ;
        RECT 345.290 34.820 349.590 35.100 ;
        RECT 355.420 34.820 360.790 35.100 ;
        RECT 364.330 34.820 389.910 35.100 ;
        RECT 286.700 34.680 293.200 34.820 ;
        RECT 286.700 34.460 289.200 34.680 ;
        RECT 349.770 34.260 363.590 34.540 ;
        RECT 408.570 33.700 418.470 33.980 ;
        RECT 343.610 32.020 416.230 32.300 ;
        RECT 427.050 32.020 459.350 32.300 ;
        RECT 428.730 31.460 458.790 31.740 ;
        RECT 360.410 30.900 363.590 31.180 ;
        RECT 364.890 30.900 387.110 31.180 ;
        RECT 443.290 30.900 458.230 31.180 ;
        RECT 335.210 30.340 336.710 30.620 ;
        RECT 381.690 30.340 384.310 30.620 ;
        RECT 386.170 30.340 408.950 30.620 ;
        RECT 431.530 30.340 455.990 30.620 ;
        RECT 369.930 29.780 384.870 30.060 ;
        RECT 438.250 29.780 446.470 30.060 ;
        RECT 453.930 29.780 459.910 30.060 ;
        RECT 458.410 29.220 460.470 29.500 ;
        RECT 335.210 28.660 335.590 28.940 ;
        RECT 335.260 28.380 335.540 28.660 ;
        RECT 332.970 28.100 343.990 28.380 ;
        RECT 317.850 26.980 331.340 27.260 ;
        RECT 334.650 26.980 361.910 27.260 ;
        RECT 391.770 26.980 393.830 27.260 ;
        RECT 411.370 26.980 415.670 27.260 ;
        RECT 416.970 26.980 434.710 27.260 ;
        RECT 331.060 26.700 331.340 26.980 ;
        RECT 331.060 26.420 331.670 26.700 ;
        RECT 418.090 26.420 421.830 26.700 ;
        RECT 302.730 25.860 303.110 26.140 ;
        RECT 435.450 25.860 454.870 26.140 ;
        RECT 286.700 25.160 289.200 25.380 ;
        RECT 286.700 25.020 293.200 25.160 ;
        RECT 302.780 25.020 303.060 25.860 ;
        RECT 286.700 24.740 303.060 25.020 ;
        RECT 286.700 24.600 293.200 24.740 ;
        RECT 286.700 24.380 289.200 24.600 ;
        RECT 321.770 24.180 334.470 24.460 ;
        RECT 428.780 23.620 443.670 23.900 ;
        RECT 428.780 23.340 429.060 23.620 ;
        RECT 344.170 23.060 348.470 23.340 ;
        RECT 386.730 23.060 389.910 23.340 ;
        RECT 427.050 23.060 429.110 23.340 ;
        RECT 436.570 23.060 455.990 23.340 ;
        RECT 334.090 22.500 346.790 22.780 ;
        RECT 385.610 22.500 418.470 22.780 ;
        RECT 362.090 21.940 370.310 22.220 ;
        RECT 418.700 21.940 435.270 22.220 ;
        RECT 446.090 21.940 457.670 22.220 ;
        RECT 418.700 21.660 418.980 21.940 ;
        RECT 387.290 21.380 407.830 21.660 ;
        RECT 418.650 21.380 419.030 21.660 ;
        RECT 434.330 21.380 439.190 21.660 ;
        RECT 418.700 20.540 418.980 21.380 ;
        RECT 346.410 20.260 418.980 20.540 ;
        RECT 427.610 20.260 449.830 20.540 ;
        RECT 302.780 19.700 342.870 19.980 ;
        RECT 383.370 19.700 383.750 19.980 ;
        RECT 407.450 19.700 435.830 19.980 ;
        RECT 437.130 19.700 448.150 19.980 ;
        RECT 302.780 19.420 303.060 19.700 ;
        RECT 383.420 19.420 383.700 19.700 ;
        RECT 437.180 19.420 437.460 19.700 ;
        RECT 302.730 19.140 303.110 19.420 ;
        RECT 313.930 19.140 324.390 19.420 ;
        RECT 367.130 19.140 367.510 19.420 ;
        RECT 382.250 19.140 388.230 19.420 ;
        RECT 389.530 19.140 404.470 19.420 ;
        RECT 431.530 19.140 437.460 19.420 ;
        RECT 367.180 18.300 367.460 19.140 ;
        RECT 369.370 18.580 383.750 18.860 ;
        RECT 422.570 18.580 426.310 18.860 ;
        RECT 316.730 18.020 329.430 18.300 ;
        RECT 367.180 18.020 390.140 18.300 ;
        RECT 115.555 17.335 116.755 17.735 ;
        RECT 389.860 16.620 390.140 18.020 ;
        RECT 389.860 16.340 400.550 16.620 ;
        RECT 404.650 16.340 420.100 16.620 ;
        RECT 439.370 16.340 457.670 16.620 ;
        RECT 298.810 15.780 299.190 16.060 ;
        RECT 286.700 15.080 289.200 15.300 ;
        RECT 286.700 14.940 293.200 15.080 ;
        RECT 298.860 14.940 299.140 15.780 ;
        RECT 419.820 15.500 420.100 16.340 ;
        RECT 325.130 15.220 364.150 15.500 ;
        RECT 393.450 15.220 417.350 15.500 ;
        RECT 419.770 15.220 424.070 15.500 ;
        RECT 431.580 15.220 436.390 15.500 ;
        RECT 431.580 14.940 431.860 15.220 ;
        RECT -189.405 13.575 -189.005 14.775 ;
        RECT 286.700 14.660 299.140 14.940 ;
        RECT 326.810 14.660 345.670 14.940 ;
        RECT 349.210 14.660 380.900 14.940 ;
        RECT 286.700 14.520 293.200 14.660 ;
        RECT 286.700 14.300 289.200 14.520 ;
        RECT 320.650 14.100 325.510 14.380 ;
        RECT 343.050 14.100 357.430 14.380 ;
        RECT 380.620 13.820 380.900 14.660 ;
        RECT 384.540 14.660 431.860 14.940 ;
        RECT 435.450 14.660 442.550 14.940 ;
        RECT 384.540 14.380 384.820 14.660 ;
        RECT 381.690 14.100 384.820 14.380 ;
        RECT 389.860 14.100 402.230 14.380 ;
        RECT 429.850 14.100 435.270 14.380 ;
        RECT 389.860 13.820 390.140 14.100 ;
        RECT 380.620 13.540 390.140 13.820 ;
        RECT 404.090 12.980 407.270 13.260 ;
        RECT 423.460 12.980 439.190 13.260 ;
        RECT 423.460 12.700 423.740 12.980 ;
        RECT 312.300 12.420 326.070 12.700 ;
        RECT 381.130 12.420 388.790 12.700 ;
        RECT 389.860 12.420 423.740 12.700 ;
        RECT 426.490 12.420 428.550 12.700 ;
        RECT 312.300 11.580 312.580 12.420 ;
        RECT 389.860 12.140 390.140 12.420 ;
        RECT 426.540 12.140 426.820 12.420 ;
        RECT 324.570 11.860 327.750 12.140 ;
        RECT 344.730 11.860 390.140 12.140 ;
        RECT 392.330 11.860 426.820 12.140 ;
        RECT 297.690 11.300 312.630 11.580 ;
        RECT 318.410 11.300 326.070 11.580 ;
        RECT 346.410 11.300 383.190 11.580 ;
        RECT 359.290 10.740 367.510 11.020 ;
        RECT 359.340 10.460 359.620 10.740 ;
        RECT 355.930 10.180 359.620 10.460 ;
        RECT 369.420 10.460 369.700 11.300 ;
        RECT 401.290 10.740 434.150 11.020 ;
        RECT 447.210 10.740 460.470 11.020 ;
        RECT 369.420 10.180 370.310 10.460 ;
        RECT 407.450 10.180 433.030 10.460 ;
        RECT 308.890 9.620 310.950 9.900 ;
        RECT 322.330 7.940 345.110 8.220 ;
        RECT 433.770 7.940 436.950 8.220 ;
        RECT 235.860 1.720 237.460 7.720 ;
        RECT 299.370 7.380 305.910 7.660 ;
        RECT 310.570 7.380 319.910 7.660 ;
        RECT 403.530 7.380 407.270 7.660 ;
        RECT 303.850 6.820 322.150 7.100 ;
        RECT 407.450 6.820 410.630 7.100 ;
        RECT 423.130 6.820 446.470 7.100 ;
        RECT 312.810 6.260 317.110 6.540 ;
        RECT 327.370 6.260 396.630 6.540 ;
        RECT 402.970 6.260 427.430 6.540 ;
        RECT 286.700 5.000 289.200 5.220 ;
        RECT 308.330 5.140 327.190 5.420 ;
        RECT 286.700 4.860 293.200 5.000 ;
        RECT 286.700 4.580 298.630 4.860 ;
        RECT 303.850 4.580 306.140 4.860 ;
        RECT 321.770 4.580 332.230 4.860 ;
        RECT 364.660 4.580 426.870 4.860 ;
        RECT 286.700 4.440 293.200 4.580 ;
        RECT 286.700 4.220 289.200 4.440 ;
        RECT 305.860 4.300 306.140 4.580 ;
        RECT 364.660 4.300 364.940 4.580 ;
        RECT 305.860 4.020 364.940 4.300 ;
        RECT 392.330 4.020 400.550 4.300 ;
        RECT 428.170 4.020 432.470 4.300 ;
        RECT 301.610 3.460 310.390 3.740 ;
        RECT 330.730 3.460 331.110 3.740 ;
        RECT 394.570 3.460 398.310 3.740 ;
        RECT 454.490 3.460 454.870 3.740 ;
        RECT 312.250 2.900 324.950 3.180 ;
        RECT 330.780 2.620 331.060 3.460 ;
        RECT 346.410 2.900 389.350 3.180 ;
        RECT 454.540 2.620 454.820 3.460 ;
        RECT 330.780 2.340 371.990 2.620 ;
        RECT 373.850 2.340 387.110 2.620 ;
        RECT 442.730 2.340 454.820 2.620 ;
        RECT 409.130 1.220 435.830 1.500 ;
        RECT 304.970 0.660 347.910 0.940 ;
        RECT 356.490 0.660 392.150 0.940 ;
        RECT 437.130 0.660 457.620 0.940 ;
        RECT 351.450 0.100 398.870 0.380 ;
        RECT 457.340 -0.180 457.620 0.660 ;
        RECT 318.460 -0.460 319.910 -0.180 ;
        RECT 364.330 -0.460 368.630 -0.180 ;
        RECT 386.170 -0.460 408.950 -0.180 ;
        RECT 435.450 -0.460 448.940 -0.180 ;
        RECT 457.290 -0.460 457.670 -0.180 ;
        RECT 318.460 -0.740 318.740 -0.460 ;
        RECT 448.660 -0.740 448.940 -0.460 ;
        RECT 316.170 -1.020 318.790 -0.740 ;
        RECT 363.210 -1.020 372.550 -0.740 ;
        RECT 412.490 -1.020 425.190 -0.740 ;
        RECT 448.660 -1.020 459.910 -0.740 ;
        RECT 331.290 -1.580 350.710 -1.300 ;
        RECT 358.730 -1.580 363.030 -1.300 ;
        RECT 384.490 -1.580 388.230 -1.300 ;
        RECT 396.810 -1.580 412.310 -1.300 ;
        RECT 320.650 -2.140 323.830 -1.860 ;
        RECT 388.410 -2.140 390.470 -1.860 ;
        RECT 407.450 -2.140 409.510 -1.860 ;
        RECT 300.490 -3.260 320.470 -2.980 ;
        RECT 325.690 -3.260 405.030 -2.980 ;
        RECT 318.970 -3.820 376.470 -3.540 ;
        RECT 229.700 -5.865 235.700 -4.265 ;
        RECT 299.370 -4.380 304.790 -4.100 ;
        RECT 311.690 -4.380 337.270 -4.100 ;
        RECT 346.970 -4.380 351.270 -4.100 ;
        RECT 383.930 -4.380 394.950 -4.100 ;
        RECT 411.930 -4.380 424.070 -4.100 ;
        RECT 387.900 -4.660 388.180 -4.380 ;
        RECT 286.700 -5.080 289.200 -4.860 ;
        RECT 323.450 -4.940 331.110 -4.660 ;
        RECT 349.210 -4.940 356.870 -4.660 ;
        RECT 387.850 -4.940 388.230 -4.660 ;
        RECT 390.090 -4.940 402.180 -4.660 ;
        RECT 286.700 -5.220 293.200 -5.080 ;
        RECT 286.700 -5.500 299.190 -5.220 ;
        RECT 360.410 -5.500 364.710 -5.220 ;
        RECT 389.860 -5.500 397.750 -5.220 ;
        RECT 286.700 -5.640 293.200 -5.500 ;
        RECT 286.700 -5.860 289.200 -5.640 ;
        RECT 389.860 -5.780 390.140 -5.500 ;
        RECT 361.530 -6.060 390.140 -5.780 ;
        RECT 391.210 -6.060 397.190 -5.780 ;
        RECT 401.900 -6.340 402.180 -4.940 ;
        RECT 349.770 -6.620 354.070 -6.340 ;
        RECT 401.850 -6.620 402.230 -6.340 ;
        RECT 403.530 -6.620 420.150 -6.340 ;
        RECT 432.650 -6.620 437.510 -6.340 ;
        RECT 403.580 -6.900 403.860 -6.620 ;
        RECT 382.250 -7.180 398.820 -6.900 ;
        RECT 399.610 -7.180 403.860 -6.900 ;
        RECT 436.570 -7.180 445.350 -6.900 ;
        RECT 398.540 -7.460 398.820 -7.180 ;
        RECT 345.290 -7.740 389.910 -7.460 ;
        RECT 398.540 -7.740 414.550 -7.460 ;
        RECT 438.250 -7.740 443.670 -7.460 ;
        RECT 305.530 -8.300 308.710 -8.020 ;
        RECT 387.290 -8.300 392.150 -8.020 ;
        RECT 396.250 -8.300 405.030 -8.020 ;
        RECT 422.570 -8.300 427.430 -8.020 ;
        RECT 345.850 -8.860 362.470 -8.580 ;
        RECT 363.210 -8.860 369.750 -8.580 ;
        RECT 385.050 -8.860 396.070 -8.580 ;
        RECT 404.090 -8.860 412.310 -8.580 ;
        RECT 362.650 -9.420 368.630 -9.140 ;
        RECT 372.170 -9.420 377.590 -9.140 ;
        RECT 396.250 -9.420 419.030 -9.140 ;
        RECT 448.660 -9.420 461.030 -9.140 ;
        RECT 448.660 -10.260 448.940 -9.420 ;
        RECT 431.530 -10.540 448.940 -10.260 ;
        RECT 366.570 -11.100 429.110 -10.820 ;
        RECT 443.290 -11.100 446.470 -10.820 ;
        RECT 353.690 -11.660 366.390 -11.380 ;
        RECT 371.050 -11.660 380.390 -11.380 ;
        RECT 404.650 -11.660 424.630 -11.380 ;
        RECT 429.290 -11.660 455.430 -11.380 ;
        RECT 360.970 -12.220 379.830 -11.940 ;
        RECT 390.650 -12.220 412.870 -11.940 ;
        RECT 430.410 -12.220 441.430 -11.940 ;
        RECT 369.370 -12.780 392.710 -12.500 ;
        RECT 393.500 -12.780 419.590 -12.500 ;
        RECT 393.500 -13.060 393.780 -12.780 ;
        RECT 380.010 -13.340 393.780 -13.060 ;
        RECT 394.620 -13.340 401.110 -13.060 ;
        RECT -189.405 -14.775 -189.005 -13.575 ;
        RECT 394.620 -13.620 394.900 -13.340 ;
        RECT 376.090 -13.900 383.750 -13.620 ;
        RECT 389.530 -13.900 394.900 -13.620 ;
        RECT 366.010 -14.460 385.430 -14.180 ;
        RECT 388.970 -14.460 396.070 -14.180 ;
        RECT 401.850 -14.460 411.190 -14.180 ;
        RECT 286.700 -15.160 289.200 -14.940 ;
        RECT 363.210 -15.020 384.870 -14.740 ;
        RECT 385.610 -15.020 398.310 -14.740 ;
        RECT 286.700 -15.300 293.200 -15.160 ;
        RECT 286.700 -15.580 299.190 -15.300 ;
        RECT 305.530 -15.580 313.190 -15.300 ;
        RECT 330.730 -15.580 421.830 -15.300 ;
        RECT 286.700 -15.720 293.200 -15.580 ;
        RECT 286.700 -15.940 289.200 -15.720 ;
        RECT 321.770 -16.140 329.430 -15.860 ;
        RECT 353.130 -16.140 383.700 -15.860 ;
        RECT 384.490 -16.140 390.470 -15.860 ;
        RECT 392.890 -16.140 407.830 -15.860 ;
        RECT 420.890 -16.140 424.070 -15.860 ;
        RECT 383.420 -16.420 383.700 -16.140 ;
        RECT 303.850 -16.700 309.830 -16.420 ;
        RECT 360.410 -16.700 370.870 -16.420 ;
        RECT 372.730 -16.700 382.630 -16.420 ;
        RECT 383.420 -16.700 403.350 -16.420 ;
        RECT 408.570 -16.700 415.110 -16.420 ;
        RECT -188.285 -18.135 -187.885 -16.935 ;
        RECT 420.940 -16.980 421.220 -16.140 ;
        RECT 302.730 -17.260 322.150 -16.980 ;
        RECT 359.290 -17.260 367.510 -16.980 ;
        RECT 375.530 -17.260 385.990 -16.980 ;
        RECT 397.930 -17.260 421.220 -16.980 ;
        RECT 449.450 -17.260 456.550 -16.980 ;
        RECT 115.555 -17.735 116.755 -17.335 ;
        RECT -332.765 -21.495 -332.365 -20.295 ;
        RECT -44.925 -21.495 -44.525 -20.295 ;
        RECT 113.755 -21.095 114.955 -20.695 ;
        RECT -404.445 -24.855 -404.045 -23.655 ;
        RECT -261.085 -24.855 -260.685 -23.655 ;
        RECT -116.605 -24.855 -116.205 -23.655 ;
        RECT 26.755 -24.855 27.155 -23.655 ;
        RECT 111.955 -24.455 113.155 -24.055 ;
        RECT -440.285 -28.215 -439.885 -27.015 ;
        RECT -368.605 -28.215 -368.205 -27.015 ;
        RECT -296.925 -28.215 -296.525 -27.015 ;
        RECT -225.245 -28.215 -224.845 -27.015 ;
        RECT -152.445 -28.215 -152.045 -27.015 ;
        RECT -80.765 -28.215 -80.365 -27.015 ;
        RECT -9.085 -28.215 -8.685 -27.015 ;
        RECT 62.595 -28.215 62.995 -27.015 ;
        RECT 110.155 -27.815 111.355 -27.415 ;
        RECT -458.205 -31.575 -457.805 -30.375 ;
        RECT -422.365 -31.575 -421.965 -30.375 ;
        RECT -386.525 -31.575 -386.125 -30.375 ;
        RECT -350.685 -31.575 -350.285 -30.375 ;
        RECT -314.845 -31.575 -314.445 -30.375 ;
        RECT -279.005 -31.575 -278.605 -30.375 ;
        RECT -243.165 -31.575 -242.765 -30.375 ;
        RECT -207.325 -31.575 -206.925 -30.375 ;
        RECT -170.365 -31.575 -169.965 -30.375 ;
        RECT -134.525 -31.575 -134.125 -30.375 ;
        RECT -98.685 -31.575 -98.285 -30.375 ;
        RECT -62.845 -31.575 -62.445 -30.375 ;
        RECT -27.005 -31.575 -26.605 -30.375 ;
        RECT 8.835 -31.575 9.235 -30.375 ;
        RECT 44.675 -31.575 45.075 -30.375 ;
        RECT 80.515 -31.575 80.915 -30.375 ;
        RECT 108.355 -31.175 109.555 -30.775 ;
        RECT -467.165 -34.935 -466.765 -33.735 ;
        RECT -449.245 -34.935 -448.845 -33.735 ;
        RECT -431.325 -34.935 -430.925 -33.735 ;
        RECT -413.405 -34.935 -413.005 -33.735 ;
        RECT -395.485 -34.935 -395.085 -33.735 ;
        RECT -377.565 -34.935 -377.165 -33.735 ;
        RECT -359.645 -34.935 -359.245 -33.735 ;
        RECT -341.725 -34.935 -341.325 -33.735 ;
        RECT -323.805 -34.935 -323.405 -33.735 ;
        RECT -305.885 -34.935 -305.485 -33.735 ;
        RECT -287.965 -34.935 -287.565 -33.735 ;
        RECT -270.045 -34.935 -269.645 -33.735 ;
        RECT -252.125 -34.935 -251.725 -33.735 ;
        RECT -234.205 -34.935 -233.805 -33.735 ;
        RECT -216.285 -34.935 -215.885 -33.735 ;
        RECT -198.365 -34.935 -197.965 -33.735 ;
        RECT -179.325 -34.935 -178.925 -33.735 ;
        RECT -161.405 -34.935 -161.005 -33.735 ;
        RECT -143.485 -34.935 -143.085 -33.735 ;
        RECT -125.565 -34.935 -125.165 -33.735 ;
        RECT -107.645 -34.935 -107.245 -33.735 ;
        RECT -89.725 -34.935 -89.325 -33.735 ;
        RECT -71.805 -34.935 -71.405 -33.735 ;
        RECT -53.885 -34.935 -53.485 -33.735 ;
        RECT -35.965 -34.935 -35.565 -33.735 ;
        RECT -18.045 -34.935 -17.645 -33.735 ;
        RECT -0.125 -34.935 0.275 -33.735 ;
        RECT 17.795 -34.935 18.195 -33.735 ;
        RECT 35.715 -34.935 36.115 -33.735 ;
        RECT 53.635 -34.935 54.035 -33.735 ;
        RECT 71.555 -34.935 71.955 -33.735 ;
        RECT 89.475 -34.935 89.875 -33.735 ;
        RECT 106.555 -34.535 107.755 -34.135 ;
        RECT -471.645 -38.295 -471.245 -37.095 ;
        RECT -462.685 -38.295 -462.285 -37.095 ;
        RECT -453.725 -38.295 -453.325 -37.095 ;
        RECT -444.765 -38.295 -444.365 -37.095 ;
        RECT -435.805 -38.295 -435.405 -37.095 ;
        RECT -426.845 -38.295 -426.445 -37.095 ;
        RECT -417.885 -38.295 -417.485 -37.095 ;
        RECT -408.925 -38.295 -408.525 -37.095 ;
        RECT -399.965 -38.295 -399.565 -37.095 ;
        RECT -391.005 -38.295 -390.605 -37.095 ;
        RECT -382.045 -38.295 -381.645 -37.095 ;
        RECT -373.085 -38.295 -372.685 -37.095 ;
        RECT -364.125 -38.295 -363.725 -37.095 ;
        RECT -355.165 -38.295 -354.765 -37.095 ;
        RECT -346.205 -38.295 -345.805 -37.095 ;
        RECT -337.245 -38.295 -336.845 -37.095 ;
        RECT -328.285 -38.295 -327.885 -37.095 ;
        RECT -319.325 -38.295 -318.925 -37.095 ;
        RECT -310.365 -38.295 -309.965 -37.095 ;
        RECT -301.405 -38.295 -301.005 -37.095 ;
        RECT -292.445 -38.295 -292.045 -37.095 ;
        RECT -283.485 -38.295 -283.085 -37.095 ;
        RECT -274.525 -38.295 -274.125 -37.095 ;
        RECT -265.565 -38.295 -265.165 -37.095 ;
        RECT -256.605 -38.295 -256.205 -37.095 ;
        RECT -247.645 -38.295 -247.245 -37.095 ;
        RECT -238.685 -38.295 -238.285 -37.095 ;
        RECT -229.725 -38.295 -229.325 -37.095 ;
        RECT -220.765 -38.295 -220.365 -37.095 ;
        RECT -211.805 -38.295 -211.405 -37.095 ;
        RECT -202.845 -38.295 -202.445 -37.095 ;
        RECT -193.885 -38.295 -193.485 -37.095 ;
        RECT -183.805 -38.295 -183.405 -37.095 ;
        RECT -174.845 -38.295 -174.445 -37.095 ;
        RECT -165.885 -38.295 -165.485 -37.095 ;
        RECT -156.925 -38.295 -156.525 -37.095 ;
        RECT -147.965 -38.295 -147.565 -37.095 ;
        RECT -139.005 -38.295 -138.605 -37.095 ;
        RECT -130.045 -38.295 -129.645 -37.095 ;
        RECT -121.085 -38.295 -120.685 -37.095 ;
        RECT -112.125 -38.295 -111.725 -37.095 ;
        RECT -103.165 -38.295 -102.765 -37.095 ;
        RECT -94.205 -38.295 -93.805 -37.095 ;
        RECT -85.245 -38.295 -84.845 -37.095 ;
        RECT -76.285 -38.295 -75.885 -37.095 ;
        RECT -67.325 -38.295 -66.925 -37.095 ;
        RECT -58.365 -38.295 -57.965 -37.095 ;
        RECT -49.405 -38.295 -49.005 -37.095 ;
        RECT -40.445 -38.295 -40.045 -37.095 ;
        RECT -31.485 -38.295 -31.085 -37.095 ;
        RECT -22.525 -38.295 -22.125 -37.095 ;
        RECT -13.565 -38.295 -13.165 -37.095 ;
        RECT -4.605 -38.295 -4.205 -37.095 ;
        RECT 4.355 -38.295 4.755 -37.095 ;
        RECT 13.315 -38.295 13.715 -37.095 ;
        RECT 22.275 -38.295 22.675 -37.095 ;
        RECT 31.235 -38.295 31.635 -37.095 ;
        RECT 40.195 -38.295 40.595 -37.095 ;
        RECT 49.155 -38.295 49.555 -37.095 ;
        RECT 58.115 -38.295 58.515 -37.095 ;
        RECT 67.075 -38.295 67.475 -37.095 ;
        RECT 76.035 -38.295 76.435 -37.095 ;
        RECT 84.995 -38.295 85.395 -37.095 ;
        RECT 93.955 -38.295 94.355 -37.095 ;
        RECT 104.755 -37.895 105.955 -37.495 ;
        RECT -473.885 -41.655 -473.485 -40.455 ;
        RECT -469.405 -41.655 -469.005 -40.455 ;
        RECT -464.925 -41.655 -464.525 -40.455 ;
        RECT -460.445 -41.655 -460.045 -40.455 ;
        RECT -455.965 -41.655 -455.565 -40.455 ;
        RECT -451.485 -41.655 -451.085 -40.455 ;
        RECT -447.005 -41.655 -446.605 -40.455 ;
        RECT -442.525 -41.655 -442.125 -40.455 ;
        RECT -438.045 -41.655 -437.645 -40.455 ;
        RECT -433.565 -41.655 -433.165 -40.455 ;
        RECT -429.085 -41.655 -428.685 -40.455 ;
        RECT -424.605 -41.655 -424.205 -40.455 ;
        RECT -420.125 -41.655 -419.725 -40.455 ;
        RECT -415.645 -41.655 -415.245 -40.455 ;
        RECT -411.165 -41.655 -410.765 -40.455 ;
        RECT -406.685 -41.655 -406.285 -40.455 ;
        RECT -402.205 -41.655 -401.805 -40.455 ;
        RECT -397.725 -41.655 -397.325 -40.455 ;
        RECT -393.245 -41.655 -392.845 -40.455 ;
        RECT -388.765 -41.655 -388.365 -40.455 ;
        RECT -384.285 -41.655 -383.885 -40.455 ;
        RECT -379.805 -41.655 -379.405 -40.455 ;
        RECT -375.325 -41.655 -374.925 -40.455 ;
        RECT -370.845 -41.655 -370.445 -40.455 ;
        RECT -366.365 -41.655 -365.965 -40.455 ;
        RECT -361.885 -41.655 -361.485 -40.455 ;
        RECT -357.405 -41.655 -357.005 -40.455 ;
        RECT -352.925 -41.655 -352.525 -40.455 ;
        RECT -348.445 -41.655 -348.045 -40.455 ;
        RECT -343.965 -41.655 -343.565 -40.455 ;
        RECT -339.485 -41.655 -339.085 -40.455 ;
        RECT -335.005 -41.655 -334.605 -40.455 ;
        RECT -330.525 -41.655 -330.125 -40.455 ;
        RECT -326.045 -41.655 -325.645 -40.455 ;
        RECT -321.565 -41.655 -321.165 -40.455 ;
        RECT -317.085 -41.655 -316.685 -40.455 ;
        RECT -312.605 -41.655 -312.205 -40.455 ;
        RECT -308.125 -41.655 -307.725 -40.455 ;
        RECT -303.645 -41.655 -303.245 -40.455 ;
        RECT -299.165 -41.655 -298.765 -40.455 ;
        RECT -294.685 -41.655 -294.285 -40.455 ;
        RECT -290.205 -41.655 -289.805 -40.455 ;
        RECT -285.725 -41.655 -285.325 -40.455 ;
        RECT -281.245 -41.655 -280.845 -40.455 ;
        RECT -276.765 -41.655 -276.365 -40.455 ;
        RECT -272.285 -41.655 -271.885 -40.455 ;
        RECT -267.805 -41.655 -267.405 -40.455 ;
        RECT -263.325 -41.655 -262.925 -40.455 ;
        RECT -258.845 -41.655 -258.445 -40.455 ;
        RECT -254.365 -41.655 -253.965 -40.455 ;
        RECT -249.885 -41.655 -249.485 -40.455 ;
        RECT -245.405 -41.655 -245.005 -40.455 ;
        RECT -240.925 -41.655 -240.525 -40.455 ;
        RECT -236.445 -41.655 -236.045 -40.455 ;
        RECT -231.965 -41.655 -231.565 -40.455 ;
        RECT -227.485 -41.655 -227.085 -40.455 ;
        RECT -223.005 -41.655 -222.605 -40.455 ;
        RECT -218.525 -41.655 -218.125 -40.455 ;
        RECT -214.045 -41.655 -213.645 -40.455 ;
        RECT -209.565 -41.655 -209.165 -40.455 ;
        RECT -205.085 -41.655 -204.685 -40.455 ;
        RECT -200.605 -41.655 -200.205 -40.455 ;
        RECT -196.125 -41.655 -195.725 -40.455 ;
        RECT -191.645 -41.655 -191.245 -40.455 ;
        RECT -186.045 -41.655 -185.645 -40.455 ;
        RECT -181.565 -41.655 -181.165 -40.455 ;
        RECT -177.085 -41.655 -176.685 -40.455 ;
        RECT -172.605 -41.655 -172.205 -40.455 ;
        RECT -168.125 -41.655 -167.725 -40.455 ;
        RECT -163.645 -41.655 -163.245 -40.455 ;
        RECT -159.165 -41.655 -158.765 -40.455 ;
        RECT -154.685 -41.655 -154.285 -40.455 ;
        RECT -150.205 -41.655 -149.805 -40.455 ;
        RECT -145.725 -41.655 -145.325 -40.455 ;
        RECT -141.245 -41.655 -140.845 -40.455 ;
        RECT -136.765 -41.655 -136.365 -40.455 ;
        RECT -132.285 -41.655 -131.885 -40.455 ;
        RECT -127.805 -41.655 -127.405 -40.455 ;
        RECT -123.325 -41.655 -122.925 -40.455 ;
        RECT -118.845 -41.655 -118.445 -40.455 ;
        RECT -114.365 -41.655 -113.965 -40.455 ;
        RECT -109.885 -41.655 -109.485 -40.455 ;
        RECT -105.405 -41.655 -105.005 -40.455 ;
        RECT -100.925 -41.655 -100.525 -40.455 ;
        RECT -96.445 -41.655 -96.045 -40.455 ;
        RECT -91.965 -41.655 -91.565 -40.455 ;
        RECT -87.485 -41.655 -87.085 -40.455 ;
        RECT -83.005 -41.655 -82.605 -40.455 ;
        RECT -78.525 -41.655 -78.125 -40.455 ;
        RECT -74.045 -41.655 -73.645 -40.455 ;
        RECT -69.565 -41.655 -69.165 -40.455 ;
        RECT -65.085 -41.655 -64.685 -40.455 ;
        RECT -60.605 -41.655 -60.205 -40.455 ;
        RECT -56.125 -41.655 -55.725 -40.455 ;
        RECT -51.645 -41.655 -51.245 -40.455 ;
        RECT -47.165 -41.655 -46.765 -40.455 ;
        RECT -42.685 -41.655 -42.285 -40.455 ;
        RECT -38.205 -41.655 -37.805 -40.455 ;
        RECT -33.725 -41.655 -33.325 -40.455 ;
        RECT -29.245 -41.655 -28.845 -40.455 ;
        RECT -24.765 -41.655 -24.365 -40.455 ;
        RECT -20.285 -41.655 -19.885 -40.455 ;
        RECT -15.805 -41.655 -15.405 -40.455 ;
        RECT -11.325 -41.655 -10.925 -40.455 ;
        RECT -6.845 -41.655 -6.445 -40.455 ;
        RECT -2.365 -41.655 -1.965 -40.455 ;
        RECT 2.115 -41.655 2.515 -40.455 ;
        RECT 6.595 -41.655 6.995 -40.455 ;
        RECT 11.075 -41.655 11.475 -40.455 ;
        RECT 15.555 -41.655 15.955 -40.455 ;
        RECT 20.035 -41.655 20.435 -40.455 ;
        RECT 24.515 -41.655 24.915 -40.455 ;
        RECT 28.995 -41.655 29.395 -40.455 ;
        RECT 33.475 -41.655 33.875 -40.455 ;
        RECT 37.955 -41.655 38.355 -40.455 ;
        RECT 42.435 -41.655 42.835 -40.455 ;
        RECT 46.915 -41.655 47.315 -40.455 ;
        RECT 51.395 -41.655 51.795 -40.455 ;
        RECT 55.875 -41.655 56.275 -40.455 ;
        RECT 60.355 -41.655 60.755 -40.455 ;
        RECT 64.835 -41.655 65.235 -40.455 ;
        RECT 69.315 -41.655 69.715 -40.455 ;
        RECT 73.795 -41.655 74.195 -40.455 ;
        RECT 78.275 -41.655 78.675 -40.455 ;
        RECT 82.755 -41.655 83.155 -40.455 ;
        RECT 87.235 -41.655 87.635 -40.455 ;
        RECT 91.715 -41.655 92.115 -40.455 ;
        RECT 96.195 -41.655 96.595 -40.455 ;
        RECT 102.955 -41.255 104.155 -40.855 ;
        RECT -475.005 -45.015 -474.605 -43.815 ;
        RECT -472.765 -45.015 -472.365 -43.815 ;
        RECT -470.525 -45.015 -470.125 -43.815 ;
        RECT -468.285 -45.015 -467.885 -43.815 ;
        RECT -466.045 -45.015 -465.645 -43.815 ;
        RECT -463.805 -45.015 -463.405 -43.815 ;
        RECT -461.565 -45.015 -461.165 -43.815 ;
        RECT -459.325 -45.015 -458.925 -43.815 ;
        RECT -457.085 -45.015 -456.685 -43.815 ;
        RECT -454.845 -45.015 -454.445 -43.815 ;
        RECT -452.605 -45.015 -452.205 -43.815 ;
        RECT -450.365 -45.015 -449.965 -43.815 ;
        RECT -448.125 -45.015 -447.725 -43.815 ;
        RECT -445.885 -45.015 -445.485 -43.815 ;
        RECT -443.645 -45.015 -443.245 -43.815 ;
        RECT -441.405 -45.015 -441.005 -43.815 ;
        RECT -439.165 -45.015 -438.765 -43.815 ;
        RECT -436.925 -45.015 -436.525 -43.815 ;
        RECT -434.685 -45.015 -434.285 -43.815 ;
        RECT -432.445 -45.015 -432.045 -43.815 ;
        RECT -430.205 -45.015 -429.805 -43.815 ;
        RECT -427.965 -45.015 -427.565 -43.815 ;
        RECT -425.725 -45.015 -425.325 -43.815 ;
        RECT -423.485 -45.015 -423.085 -43.815 ;
        RECT -421.245 -45.015 -420.845 -43.815 ;
        RECT -419.005 -45.015 -418.605 -43.815 ;
        RECT -416.765 -45.015 -416.365 -43.815 ;
        RECT -414.525 -45.015 -414.125 -43.815 ;
        RECT -412.285 -45.015 -411.885 -43.815 ;
        RECT -410.045 -45.015 -409.645 -43.815 ;
        RECT -407.805 -45.015 -407.405 -43.815 ;
        RECT -405.565 -45.015 -405.165 -43.815 ;
        RECT -403.325 -45.015 -402.925 -43.815 ;
        RECT -401.085 -45.015 -400.685 -43.815 ;
        RECT -398.845 -45.015 -398.445 -43.815 ;
        RECT -396.605 -45.015 -396.205 -43.815 ;
        RECT -394.365 -45.015 -393.965 -43.815 ;
        RECT -392.125 -45.015 -391.725 -43.815 ;
        RECT -389.885 -45.015 -389.485 -43.815 ;
        RECT -387.645 -45.015 -387.245 -43.815 ;
        RECT -385.405 -45.015 -385.005 -43.815 ;
        RECT -383.165 -45.015 -382.765 -43.815 ;
        RECT -380.925 -45.015 -380.525 -43.815 ;
        RECT -378.685 -45.015 -378.285 -43.815 ;
        RECT -376.445 -45.015 -376.045 -43.815 ;
        RECT -374.205 -45.015 -373.805 -43.815 ;
        RECT -371.965 -45.015 -371.565 -43.815 ;
        RECT -369.725 -45.015 -369.325 -43.815 ;
        RECT -367.485 -45.015 -367.085 -43.815 ;
        RECT -365.245 -45.015 -364.845 -43.815 ;
        RECT -363.005 -45.015 -362.605 -43.815 ;
        RECT -360.765 -45.015 -360.365 -43.815 ;
        RECT -358.525 -45.015 -358.125 -43.815 ;
        RECT -356.285 -45.015 -355.885 -43.815 ;
        RECT -354.045 -45.015 -353.645 -43.815 ;
        RECT -351.805 -45.015 -351.405 -43.815 ;
        RECT -349.565 -45.015 -349.165 -43.815 ;
        RECT -347.325 -45.015 -346.925 -43.815 ;
        RECT -345.085 -45.015 -344.685 -43.815 ;
        RECT -342.845 -45.015 -342.445 -43.815 ;
        RECT -340.605 -45.015 -340.205 -43.815 ;
        RECT -338.365 -45.015 -337.965 -43.815 ;
        RECT -336.125 -45.015 -335.725 -43.815 ;
        RECT -333.885 -45.015 -333.485 -43.815 ;
        RECT -331.645 -45.015 -331.245 -43.815 ;
        RECT -329.405 -45.015 -329.005 -43.815 ;
        RECT -327.165 -45.015 -326.765 -43.815 ;
        RECT -324.925 -45.015 -324.525 -43.815 ;
        RECT -322.685 -45.015 -322.285 -43.815 ;
        RECT -320.445 -45.015 -320.045 -43.815 ;
        RECT -318.205 -45.015 -317.805 -43.815 ;
        RECT -315.965 -45.015 -315.565 -43.815 ;
        RECT -313.725 -45.015 -313.325 -43.815 ;
        RECT -311.485 -45.015 -311.085 -43.815 ;
        RECT -309.245 -45.015 -308.845 -43.815 ;
        RECT -307.005 -45.015 -306.605 -43.815 ;
        RECT -304.765 -45.015 -304.365 -43.815 ;
        RECT -302.525 -45.015 -302.125 -43.815 ;
        RECT -300.285 -45.015 -299.885 -43.815 ;
        RECT -298.045 -45.015 -297.645 -43.815 ;
        RECT -295.805 -45.015 -295.405 -43.815 ;
        RECT -293.565 -45.015 -293.165 -43.815 ;
        RECT -291.325 -45.015 -290.925 -43.815 ;
        RECT -289.085 -45.015 -288.685 -43.815 ;
        RECT -286.845 -45.015 -286.445 -43.815 ;
        RECT -284.605 -45.015 -284.205 -43.815 ;
        RECT -282.365 -45.015 -281.965 -43.815 ;
        RECT -280.125 -45.015 -279.725 -43.815 ;
        RECT -277.885 -45.015 -277.485 -43.815 ;
        RECT -275.645 -45.015 -275.245 -43.815 ;
        RECT -273.405 -45.015 -273.005 -43.815 ;
        RECT -271.165 -45.015 -270.765 -43.815 ;
        RECT -268.925 -45.015 -268.525 -43.815 ;
        RECT -266.685 -45.015 -266.285 -43.815 ;
        RECT -264.445 -45.015 -264.045 -43.815 ;
        RECT -262.205 -45.015 -261.805 -43.815 ;
        RECT -259.965 -45.015 -259.565 -43.815 ;
        RECT -257.725 -45.015 -257.325 -43.815 ;
        RECT -255.485 -45.015 -255.085 -43.815 ;
        RECT -253.245 -45.015 -252.845 -43.815 ;
        RECT -251.005 -45.015 -250.605 -43.815 ;
        RECT -248.765 -45.015 -248.365 -43.815 ;
        RECT -246.525 -45.015 -246.125 -43.815 ;
        RECT -244.285 -45.015 -243.885 -43.815 ;
        RECT -242.045 -45.015 -241.645 -43.815 ;
        RECT -239.805 -45.015 -239.405 -43.815 ;
        RECT -237.565 -45.015 -237.165 -43.815 ;
        RECT -235.325 -45.015 -234.925 -43.815 ;
        RECT -233.085 -45.015 -232.685 -43.815 ;
        RECT -230.845 -45.015 -230.445 -43.815 ;
        RECT -228.605 -45.015 -228.205 -43.815 ;
        RECT -226.365 -45.015 -225.965 -43.815 ;
        RECT -224.125 -45.015 -223.725 -43.815 ;
        RECT -221.885 -45.015 -221.485 -43.815 ;
        RECT -219.645 -45.015 -219.245 -43.815 ;
        RECT -217.405 -45.015 -217.005 -43.815 ;
        RECT -215.165 -45.015 -214.765 -43.815 ;
        RECT -212.925 -45.015 -212.525 -43.815 ;
        RECT -210.685 -45.015 -210.285 -43.815 ;
        RECT -208.445 -45.015 -208.045 -43.815 ;
        RECT -206.205 -45.015 -205.805 -43.815 ;
        RECT -203.965 -45.015 -203.565 -43.815 ;
        RECT -201.725 -45.015 -201.325 -43.815 ;
        RECT -199.485 -45.015 -199.085 -43.815 ;
        RECT -197.245 -45.015 -196.845 -43.815 ;
        RECT -195.005 -45.015 -194.605 -43.815 ;
        RECT -192.765 -45.015 -192.365 -43.815 ;
        RECT -190.525 -45.015 -190.125 -43.815 ;
        RECT -187.165 -45.015 -186.765 -43.815 ;
        RECT -184.925 -45.015 -184.525 -43.815 ;
        RECT -182.685 -45.015 -182.285 -43.815 ;
        RECT -180.445 -45.015 -180.045 -43.815 ;
        RECT -178.205 -45.015 -177.805 -43.815 ;
        RECT -175.965 -45.015 -175.565 -43.815 ;
        RECT -173.725 -45.015 -173.325 -43.815 ;
        RECT -171.485 -45.015 -171.085 -43.815 ;
        RECT -169.245 -45.015 -168.845 -43.815 ;
        RECT -167.005 -45.015 -166.605 -43.815 ;
        RECT -164.765 -45.015 -164.365 -43.815 ;
        RECT -162.525 -45.015 -162.125 -43.815 ;
        RECT -160.285 -45.015 -159.885 -43.815 ;
        RECT -158.045 -45.015 -157.645 -43.815 ;
        RECT -155.805 -45.015 -155.405 -43.815 ;
        RECT -153.565 -45.015 -153.165 -43.815 ;
        RECT -151.325 -45.015 -150.925 -43.815 ;
        RECT -149.085 -45.015 -148.685 -43.815 ;
        RECT -146.845 -45.015 -146.445 -43.815 ;
        RECT -144.605 -45.015 -144.205 -43.815 ;
        RECT -142.365 -45.015 -141.965 -43.815 ;
        RECT -140.125 -45.015 -139.725 -43.815 ;
        RECT -137.885 -45.015 -137.485 -43.815 ;
        RECT -135.645 -45.015 -135.245 -43.815 ;
        RECT -133.405 -45.015 -133.005 -43.815 ;
        RECT -131.165 -45.015 -130.765 -43.815 ;
        RECT -128.925 -45.015 -128.525 -43.815 ;
        RECT -126.685 -45.015 -126.285 -43.815 ;
        RECT -124.445 -45.015 -124.045 -43.815 ;
        RECT -122.205 -45.015 -121.805 -43.815 ;
        RECT -119.965 -45.015 -119.565 -43.815 ;
        RECT -117.725 -45.015 -117.325 -43.815 ;
        RECT -115.485 -45.015 -115.085 -43.815 ;
        RECT -113.245 -45.015 -112.845 -43.815 ;
        RECT -111.005 -45.015 -110.605 -43.815 ;
        RECT -108.765 -45.015 -108.365 -43.815 ;
        RECT -106.525 -45.015 -106.125 -43.815 ;
        RECT -104.285 -45.015 -103.885 -43.815 ;
        RECT -102.045 -45.015 -101.645 -43.815 ;
        RECT -99.805 -45.015 -99.405 -43.815 ;
        RECT -97.565 -45.015 -97.165 -43.815 ;
        RECT -95.325 -45.015 -94.925 -43.815 ;
        RECT -93.085 -45.015 -92.685 -43.815 ;
        RECT -90.845 -45.015 -90.445 -43.815 ;
        RECT -88.605 -45.015 -88.205 -43.815 ;
        RECT -86.365 -45.015 -85.965 -43.815 ;
        RECT -84.125 -45.015 -83.725 -43.815 ;
        RECT -81.885 -45.015 -81.485 -43.815 ;
        RECT -79.645 -45.015 -79.245 -43.815 ;
        RECT -77.405 -45.015 -77.005 -43.815 ;
        RECT -75.165 -45.015 -74.765 -43.815 ;
        RECT -72.925 -45.015 -72.525 -43.815 ;
        RECT -70.685 -45.015 -70.285 -43.815 ;
        RECT -68.445 -45.015 -68.045 -43.815 ;
        RECT -66.205 -45.015 -65.805 -43.815 ;
        RECT -63.965 -45.015 -63.565 -43.815 ;
        RECT -61.725 -45.015 -61.325 -43.815 ;
        RECT -59.485 -45.015 -59.085 -43.815 ;
        RECT -57.245 -45.015 -56.845 -43.815 ;
        RECT -55.005 -45.015 -54.605 -43.815 ;
        RECT -52.765 -45.015 -52.365 -43.815 ;
        RECT -50.525 -45.015 -50.125 -43.815 ;
        RECT -48.285 -45.015 -47.885 -43.815 ;
        RECT -46.045 -45.015 -45.645 -43.815 ;
        RECT -43.805 -45.015 -43.405 -43.815 ;
        RECT -41.565 -45.015 -41.165 -43.815 ;
        RECT -39.325 -45.015 -38.925 -43.815 ;
        RECT -37.085 -45.015 -36.685 -43.815 ;
        RECT -34.845 -45.015 -34.445 -43.815 ;
        RECT -32.605 -45.015 -32.205 -43.815 ;
        RECT -30.365 -45.015 -29.965 -43.815 ;
        RECT -28.125 -45.015 -27.725 -43.815 ;
        RECT -25.885 -45.015 -25.485 -43.815 ;
        RECT -23.645 -45.015 -23.245 -43.815 ;
        RECT -21.405 -45.015 -21.005 -43.815 ;
        RECT -19.165 -45.015 -18.765 -43.815 ;
        RECT -16.925 -45.015 -16.525 -43.815 ;
        RECT -14.685 -45.015 -14.285 -43.815 ;
        RECT -12.445 -45.015 -12.045 -43.815 ;
        RECT -10.205 -45.015 -9.805 -43.815 ;
        RECT -7.965 -45.015 -7.565 -43.815 ;
        RECT -5.725 -45.015 -5.325 -43.815 ;
        RECT -3.485 -45.015 -3.085 -43.815 ;
        RECT -1.245 -45.015 -0.845 -43.815 ;
        RECT 0.995 -45.015 1.395 -43.815 ;
        RECT 3.235 -45.015 3.635 -43.815 ;
        RECT 5.475 -45.015 5.875 -43.815 ;
        RECT 7.715 -45.015 8.115 -43.815 ;
        RECT 9.955 -45.015 10.355 -43.815 ;
        RECT 12.195 -45.015 12.595 -43.815 ;
        RECT 14.435 -45.015 14.835 -43.815 ;
        RECT 16.675 -45.015 17.075 -43.815 ;
        RECT 18.915 -45.015 19.315 -43.815 ;
        RECT 21.155 -45.015 21.555 -43.815 ;
        RECT 23.395 -45.015 23.795 -43.815 ;
        RECT 25.635 -45.015 26.035 -43.815 ;
        RECT 27.875 -45.015 28.275 -43.815 ;
        RECT 30.115 -45.015 30.515 -43.815 ;
        RECT 32.355 -45.015 32.755 -43.815 ;
        RECT 34.595 -45.015 34.995 -43.815 ;
        RECT 36.835 -45.015 37.235 -43.815 ;
        RECT 39.075 -45.015 39.475 -43.815 ;
        RECT 41.315 -45.015 41.715 -43.815 ;
        RECT 43.555 -45.015 43.955 -43.815 ;
        RECT 45.795 -45.015 46.195 -43.815 ;
        RECT 48.035 -45.015 48.435 -43.815 ;
        RECT 50.275 -45.015 50.675 -43.815 ;
        RECT 52.515 -45.015 52.915 -43.815 ;
        RECT 54.755 -45.015 55.155 -43.815 ;
        RECT 56.995 -45.015 57.395 -43.815 ;
        RECT 59.235 -45.015 59.635 -43.815 ;
        RECT 61.475 -45.015 61.875 -43.815 ;
        RECT 63.715 -45.015 64.115 -43.815 ;
        RECT 65.955 -45.015 66.355 -43.815 ;
        RECT 68.195 -45.015 68.595 -43.815 ;
        RECT 70.435 -45.015 70.835 -43.815 ;
        RECT 72.675 -45.015 73.075 -43.815 ;
        RECT 74.915 -45.015 75.315 -43.815 ;
        RECT 77.155 -45.015 77.555 -43.815 ;
        RECT 79.395 -45.015 79.795 -43.815 ;
        RECT 81.635 -45.015 82.035 -43.815 ;
        RECT 83.875 -45.015 84.275 -43.815 ;
        RECT 86.115 -45.015 86.515 -43.815 ;
        RECT 88.355 -45.015 88.755 -43.815 ;
        RECT 90.595 -45.015 90.995 -43.815 ;
        RECT 92.835 -45.015 93.235 -43.815 ;
        RECT 95.075 -45.015 95.475 -43.815 ;
        RECT 97.315 -45.015 97.715 -43.815 ;
        RECT 101.155 -44.615 102.355 -44.215 ;
        RECT -475.005 -67.875 -474.605 -66.675 ;
        RECT -472.765 -67.875 -472.365 -66.675 ;
        RECT -470.525 -67.875 -470.125 -66.675 ;
        RECT -468.285 -67.875 -467.885 -66.675 ;
        RECT -466.045 -67.875 -465.645 -66.675 ;
        RECT -463.805 -67.875 -463.405 -66.675 ;
        RECT -461.565 -67.875 -461.165 -66.675 ;
        RECT -459.325 -67.875 -458.925 -66.675 ;
        RECT -457.085 -67.875 -456.685 -66.675 ;
        RECT -454.845 -67.875 -454.445 -66.675 ;
        RECT -452.605 -67.875 -452.205 -66.675 ;
        RECT -450.365 -67.875 -449.965 -66.675 ;
        RECT -448.125 -67.875 -447.725 -66.675 ;
        RECT -445.885 -67.875 -445.485 -66.675 ;
        RECT -443.645 -67.875 -443.245 -66.675 ;
        RECT -441.405 -67.875 -441.005 -66.675 ;
        RECT -439.165 -67.875 -438.765 -66.675 ;
        RECT -436.925 -67.875 -436.525 -66.675 ;
        RECT -434.685 -67.875 -434.285 -66.675 ;
        RECT -432.445 -67.875 -432.045 -66.675 ;
        RECT -430.205 -67.875 -429.805 -66.675 ;
        RECT -427.965 -67.875 -427.565 -66.675 ;
        RECT -425.725 -67.875 -425.325 -66.675 ;
        RECT -423.485 -67.875 -423.085 -66.675 ;
        RECT -421.245 -67.875 -420.845 -66.675 ;
        RECT -419.005 -67.875 -418.605 -66.675 ;
        RECT -416.765 -67.875 -416.365 -66.675 ;
        RECT -414.525 -67.875 -414.125 -66.675 ;
        RECT -412.285 -67.875 -411.885 -66.675 ;
        RECT -410.045 -67.875 -409.645 -66.675 ;
        RECT -407.805 -67.875 -407.405 -66.675 ;
        RECT -405.565 -67.875 -405.165 -66.675 ;
        RECT -403.325 -67.875 -402.925 -66.675 ;
        RECT -401.085 -67.875 -400.685 -66.675 ;
        RECT -398.845 -67.875 -398.445 -66.675 ;
        RECT -396.605 -67.875 -396.205 -66.675 ;
        RECT -394.365 -67.875 -393.965 -66.675 ;
        RECT -392.125 -67.875 -391.725 -66.675 ;
        RECT -389.885 -67.875 -389.485 -66.675 ;
        RECT -387.645 -67.875 -387.245 -66.675 ;
        RECT -385.405 -67.875 -385.005 -66.675 ;
        RECT -383.165 -67.875 -382.765 -66.675 ;
        RECT -380.925 -67.875 -380.525 -66.675 ;
        RECT -378.685 -67.875 -378.285 -66.675 ;
        RECT -376.445 -67.875 -376.045 -66.675 ;
        RECT -374.205 -67.875 -373.805 -66.675 ;
        RECT -371.965 -67.875 -371.565 -66.675 ;
        RECT -369.725 -67.875 -369.325 -66.675 ;
        RECT -367.485 -67.875 -367.085 -66.675 ;
        RECT -365.245 -67.875 -364.845 -66.675 ;
        RECT -363.005 -67.875 -362.605 -66.675 ;
        RECT -360.765 -67.875 -360.365 -66.675 ;
        RECT -358.525 -67.875 -358.125 -66.675 ;
        RECT -356.285 -67.875 -355.885 -66.675 ;
        RECT -354.045 -67.875 -353.645 -66.675 ;
        RECT -351.805 -67.875 -351.405 -66.675 ;
        RECT -349.565 -67.875 -349.165 -66.675 ;
        RECT -347.325 -67.875 -346.925 -66.675 ;
        RECT -345.085 -67.875 -344.685 -66.675 ;
        RECT -342.845 -67.875 -342.445 -66.675 ;
        RECT -340.605 -67.875 -340.205 -66.675 ;
        RECT -338.365 -67.875 -337.965 -66.675 ;
        RECT -336.125 -67.875 -335.725 -66.675 ;
        RECT -333.885 -67.875 -333.485 -66.675 ;
        RECT -331.645 -67.875 -331.245 -66.675 ;
        RECT -329.405 -67.875 -329.005 -66.675 ;
        RECT -327.165 -67.875 -326.765 -66.675 ;
        RECT -324.925 -67.875 -324.525 -66.675 ;
        RECT -322.685 -67.875 -322.285 -66.675 ;
        RECT -320.445 -67.875 -320.045 -66.675 ;
        RECT -318.205 -67.875 -317.805 -66.675 ;
        RECT -315.965 -67.875 -315.565 -66.675 ;
        RECT -313.725 -67.875 -313.325 -66.675 ;
        RECT -311.485 -67.875 -311.085 -66.675 ;
        RECT -309.245 -67.875 -308.845 -66.675 ;
        RECT -307.005 -67.875 -306.605 -66.675 ;
        RECT -304.765 -67.875 -304.365 -66.675 ;
        RECT -302.525 -67.875 -302.125 -66.675 ;
        RECT -300.285 -67.875 -299.885 -66.675 ;
        RECT -298.045 -67.875 -297.645 -66.675 ;
        RECT -295.805 -67.875 -295.405 -66.675 ;
        RECT -293.565 -67.875 -293.165 -66.675 ;
        RECT -291.325 -67.875 -290.925 -66.675 ;
        RECT -289.085 -67.875 -288.685 -66.675 ;
        RECT -286.845 -67.875 -286.445 -66.675 ;
        RECT -284.605 -67.875 -284.205 -66.675 ;
        RECT -282.365 -67.875 -281.965 -66.675 ;
        RECT -280.125 -67.875 -279.725 -66.675 ;
        RECT -277.885 -67.875 -277.485 -66.675 ;
        RECT -275.645 -67.875 -275.245 -66.675 ;
        RECT -273.405 -67.875 -273.005 -66.675 ;
        RECT -271.165 -67.875 -270.765 -66.675 ;
        RECT -268.925 -67.875 -268.525 -66.675 ;
        RECT -266.685 -67.875 -266.285 -66.675 ;
        RECT -264.445 -67.875 -264.045 -66.675 ;
        RECT -262.205 -67.875 -261.805 -66.675 ;
        RECT -259.965 -67.875 -259.565 -66.675 ;
        RECT -257.725 -67.875 -257.325 -66.675 ;
        RECT -255.485 -67.875 -255.085 -66.675 ;
        RECT -253.245 -67.875 -252.845 -66.675 ;
        RECT -251.005 -67.875 -250.605 -66.675 ;
        RECT -248.765 -67.875 -248.365 -66.675 ;
        RECT -246.525 -67.875 -246.125 -66.675 ;
        RECT -244.285 -67.875 -243.885 -66.675 ;
        RECT -242.045 -67.875 -241.645 -66.675 ;
        RECT -239.805 -67.875 -239.405 -66.675 ;
        RECT -237.565 -67.875 -237.165 -66.675 ;
        RECT -235.325 -67.875 -234.925 -66.675 ;
        RECT -233.085 -67.875 -232.685 -66.675 ;
        RECT -230.845 -67.875 -230.445 -66.675 ;
        RECT -228.605 -67.875 -228.205 -66.675 ;
        RECT -226.365 -67.875 -225.965 -66.675 ;
        RECT -224.125 -67.875 -223.725 -66.675 ;
        RECT -221.885 -67.875 -221.485 -66.675 ;
        RECT -219.645 -67.875 -219.245 -66.675 ;
        RECT -217.405 -67.875 -217.005 -66.675 ;
        RECT -215.165 -67.875 -214.765 -66.675 ;
        RECT -212.925 -67.875 -212.525 -66.675 ;
        RECT -210.685 -67.875 -210.285 -66.675 ;
        RECT -208.445 -67.875 -208.045 -66.675 ;
        RECT -206.205 -67.875 -205.805 -66.675 ;
        RECT -203.965 -67.875 -203.565 -66.675 ;
        RECT -201.725 -67.875 -201.325 -66.675 ;
        RECT -199.485 -67.875 -199.085 -66.675 ;
        RECT -197.245 -67.875 -196.845 -66.675 ;
        RECT -195.005 -67.875 -194.605 -66.675 ;
        RECT -192.765 -67.875 -192.365 -66.675 ;
        RECT -190.525 -67.875 -190.125 -66.675 ;
        RECT -187.165 -67.875 -186.765 -66.675 ;
        RECT -184.925 -67.875 -184.525 -66.675 ;
        RECT -182.685 -67.875 -182.285 -66.675 ;
        RECT -180.445 -67.875 -180.045 -66.675 ;
        RECT -178.205 -67.875 -177.805 -66.675 ;
        RECT -175.965 -67.875 -175.565 -66.675 ;
        RECT -173.725 -67.875 -173.325 -66.675 ;
        RECT -171.485 -67.875 -171.085 -66.675 ;
        RECT -169.245 -67.875 -168.845 -66.675 ;
        RECT -167.005 -67.875 -166.605 -66.675 ;
        RECT -164.765 -67.875 -164.365 -66.675 ;
        RECT -162.525 -67.875 -162.125 -66.675 ;
        RECT -160.285 -67.875 -159.885 -66.675 ;
        RECT -158.045 -67.875 -157.645 -66.675 ;
        RECT -155.805 -67.875 -155.405 -66.675 ;
        RECT -153.565 -67.875 -153.165 -66.675 ;
        RECT -151.325 -67.875 -150.925 -66.675 ;
        RECT -149.085 -67.875 -148.685 -66.675 ;
        RECT -146.845 -67.875 -146.445 -66.675 ;
        RECT -144.605 -67.875 -144.205 -66.675 ;
        RECT -142.365 -67.875 -141.965 -66.675 ;
        RECT -140.125 -67.875 -139.725 -66.675 ;
        RECT -137.885 -67.875 -137.485 -66.675 ;
        RECT -135.645 -67.875 -135.245 -66.675 ;
        RECT -133.405 -67.875 -133.005 -66.675 ;
        RECT -131.165 -67.875 -130.765 -66.675 ;
        RECT -128.925 -67.875 -128.525 -66.675 ;
        RECT -126.685 -67.875 -126.285 -66.675 ;
        RECT -124.445 -67.875 -124.045 -66.675 ;
        RECT -122.205 -67.875 -121.805 -66.675 ;
        RECT -119.965 -67.875 -119.565 -66.675 ;
        RECT -117.725 -67.875 -117.325 -66.675 ;
        RECT -115.485 -67.875 -115.085 -66.675 ;
        RECT -113.245 -67.875 -112.845 -66.675 ;
        RECT -111.005 -67.875 -110.605 -66.675 ;
        RECT -108.765 -67.875 -108.365 -66.675 ;
        RECT -106.525 -67.875 -106.125 -66.675 ;
        RECT -104.285 -67.875 -103.885 -66.675 ;
        RECT -102.045 -67.875 -101.645 -66.675 ;
        RECT -99.805 -67.875 -99.405 -66.675 ;
        RECT -97.565 -67.875 -97.165 -66.675 ;
        RECT -95.325 -67.875 -94.925 -66.675 ;
        RECT -93.085 -67.875 -92.685 -66.675 ;
        RECT -90.845 -67.875 -90.445 -66.675 ;
        RECT -88.605 -67.875 -88.205 -66.675 ;
        RECT -86.365 -67.875 -85.965 -66.675 ;
        RECT -84.125 -67.875 -83.725 -66.675 ;
        RECT -81.885 -67.875 -81.485 -66.675 ;
        RECT -79.645 -67.875 -79.245 -66.675 ;
        RECT -77.405 -67.875 -77.005 -66.675 ;
        RECT -75.165 -67.875 -74.765 -66.675 ;
        RECT -72.925 -67.875 -72.525 -66.675 ;
        RECT -70.685 -67.875 -70.285 -66.675 ;
        RECT -68.445 -67.875 -68.045 -66.675 ;
        RECT -66.205 -67.875 -65.805 -66.675 ;
        RECT -63.965 -67.875 -63.565 -66.675 ;
        RECT -61.725 -67.875 -61.325 -66.675 ;
        RECT -59.485 -67.875 -59.085 -66.675 ;
        RECT -57.245 -67.875 -56.845 -66.675 ;
        RECT -55.005 -67.875 -54.605 -66.675 ;
        RECT -52.765 -67.875 -52.365 -66.675 ;
        RECT -50.525 -67.875 -50.125 -66.675 ;
        RECT -48.285 -67.875 -47.885 -66.675 ;
        RECT -46.045 -67.875 -45.645 -66.675 ;
        RECT -43.805 -67.875 -43.405 -66.675 ;
        RECT -41.565 -67.875 -41.165 -66.675 ;
        RECT -39.325 -67.875 -38.925 -66.675 ;
        RECT -37.085 -67.875 -36.685 -66.675 ;
        RECT -34.845 -67.875 -34.445 -66.675 ;
        RECT -32.605 -67.875 -32.205 -66.675 ;
        RECT -30.365 -67.875 -29.965 -66.675 ;
        RECT -28.125 -67.875 -27.725 -66.675 ;
        RECT -25.885 -67.875 -25.485 -66.675 ;
        RECT -23.645 -67.875 -23.245 -66.675 ;
        RECT -21.405 -67.875 -21.005 -66.675 ;
        RECT -19.165 -67.875 -18.765 -66.675 ;
        RECT -16.925 -67.875 -16.525 -66.675 ;
        RECT -14.685 -67.875 -14.285 -66.675 ;
        RECT -12.445 -67.875 -12.045 -66.675 ;
        RECT -10.205 -67.875 -9.805 -66.675 ;
        RECT -7.965 -67.875 -7.565 -66.675 ;
        RECT -5.725 -67.875 -5.325 -66.675 ;
        RECT -3.485 -67.875 -3.085 -66.675 ;
        RECT -1.245 -67.875 -0.845 -66.675 ;
        RECT 0.995 -67.875 1.395 -66.675 ;
        RECT 3.235 -67.875 3.635 -66.675 ;
        RECT 5.475 -67.875 5.875 -66.675 ;
        RECT 7.715 -67.875 8.115 -66.675 ;
        RECT 9.955 -67.875 10.355 -66.675 ;
        RECT 12.195 -67.875 12.595 -66.675 ;
        RECT 14.435 -67.875 14.835 -66.675 ;
        RECT 16.675 -67.875 17.075 -66.675 ;
        RECT 18.915 -67.875 19.315 -66.675 ;
        RECT 21.155 -67.875 21.555 -66.675 ;
        RECT 23.395 -67.875 23.795 -66.675 ;
        RECT 25.635 -67.875 26.035 -66.675 ;
        RECT 27.875 -67.875 28.275 -66.675 ;
        RECT 30.115 -67.875 30.515 -66.675 ;
        RECT 32.355 -67.875 32.755 -66.675 ;
        RECT 34.595 -67.875 34.995 -66.675 ;
        RECT 36.835 -67.875 37.235 -66.675 ;
        RECT 39.075 -67.875 39.475 -66.675 ;
        RECT 41.315 -67.875 41.715 -66.675 ;
        RECT 43.555 -67.875 43.955 -66.675 ;
        RECT 45.795 -67.875 46.195 -66.675 ;
        RECT 48.035 -67.875 48.435 -66.675 ;
        RECT 50.275 -67.875 50.675 -66.675 ;
        RECT 52.515 -67.875 52.915 -66.675 ;
        RECT 54.755 -67.875 55.155 -66.675 ;
        RECT 56.995 -67.875 57.395 -66.675 ;
        RECT 59.235 -67.875 59.635 -66.675 ;
        RECT 61.475 -67.875 61.875 -66.675 ;
        RECT 63.715 -67.875 64.115 -66.675 ;
        RECT 65.955 -67.875 66.355 -66.675 ;
        RECT 68.195 -67.875 68.595 -66.675 ;
        RECT 70.435 -67.875 70.835 -66.675 ;
        RECT 72.675 -67.875 73.075 -66.675 ;
        RECT 74.915 -67.875 75.315 -66.675 ;
        RECT 77.155 -67.875 77.555 -66.675 ;
        RECT 79.395 -67.875 79.795 -66.675 ;
        RECT 81.635 -67.875 82.035 -66.675 ;
        RECT 83.875 -67.875 84.275 -66.675 ;
        RECT 86.115 -67.875 86.515 -66.675 ;
        RECT 88.355 -67.875 88.755 -66.675 ;
        RECT 90.595 -67.875 90.995 -66.675 ;
        RECT 92.835 -67.875 93.235 -66.675 ;
        RECT 95.075 -67.875 95.475 -66.675 ;
        RECT 97.315 -67.875 97.715 -66.675 ;
        RECT 101.505 -67.075 102.005 -44.615 ;
        RECT 101.155 -67.475 102.355 -67.075 ;
        RECT -473.885 -71.235 -473.485 -70.035 ;
        RECT -469.405 -71.235 -469.005 -70.035 ;
        RECT -464.925 -71.235 -464.525 -70.035 ;
        RECT -460.445 -71.235 -460.045 -70.035 ;
        RECT -455.965 -71.235 -455.565 -70.035 ;
        RECT -451.485 -71.235 -451.085 -70.035 ;
        RECT -447.005 -71.235 -446.605 -70.035 ;
        RECT -442.525 -71.235 -442.125 -70.035 ;
        RECT -438.045 -71.235 -437.645 -70.035 ;
        RECT -433.565 -71.235 -433.165 -70.035 ;
        RECT -429.085 -71.235 -428.685 -70.035 ;
        RECT -424.605 -71.235 -424.205 -70.035 ;
        RECT -420.125 -71.235 -419.725 -70.035 ;
        RECT -415.645 -71.235 -415.245 -70.035 ;
        RECT -411.165 -71.235 -410.765 -70.035 ;
        RECT -406.685 -71.235 -406.285 -70.035 ;
        RECT -402.205 -71.235 -401.805 -70.035 ;
        RECT -397.725 -71.235 -397.325 -70.035 ;
        RECT -393.245 -71.235 -392.845 -70.035 ;
        RECT -388.765 -71.235 -388.365 -70.035 ;
        RECT -384.285 -71.235 -383.885 -70.035 ;
        RECT -379.805 -71.235 -379.405 -70.035 ;
        RECT -375.325 -71.235 -374.925 -70.035 ;
        RECT -370.845 -71.235 -370.445 -70.035 ;
        RECT -366.365 -71.235 -365.965 -70.035 ;
        RECT -361.885 -71.235 -361.485 -70.035 ;
        RECT -357.405 -71.235 -357.005 -70.035 ;
        RECT -352.925 -71.235 -352.525 -70.035 ;
        RECT -348.445 -71.235 -348.045 -70.035 ;
        RECT -343.965 -71.235 -343.565 -70.035 ;
        RECT -339.485 -71.235 -339.085 -70.035 ;
        RECT -335.005 -71.235 -334.605 -70.035 ;
        RECT -330.525 -71.235 -330.125 -70.035 ;
        RECT -326.045 -71.235 -325.645 -70.035 ;
        RECT -321.565 -71.235 -321.165 -70.035 ;
        RECT -317.085 -71.235 -316.685 -70.035 ;
        RECT -312.605 -71.235 -312.205 -70.035 ;
        RECT -308.125 -71.235 -307.725 -70.035 ;
        RECT -303.645 -71.235 -303.245 -70.035 ;
        RECT -299.165 -71.235 -298.765 -70.035 ;
        RECT -294.685 -71.235 -294.285 -70.035 ;
        RECT -290.205 -71.235 -289.805 -70.035 ;
        RECT -285.725 -71.235 -285.325 -70.035 ;
        RECT -281.245 -71.235 -280.845 -70.035 ;
        RECT -276.765 -71.235 -276.365 -70.035 ;
        RECT -272.285 -71.235 -271.885 -70.035 ;
        RECT -267.805 -71.235 -267.405 -70.035 ;
        RECT -263.325 -71.235 -262.925 -70.035 ;
        RECT -258.845 -71.235 -258.445 -70.035 ;
        RECT -254.365 -71.235 -253.965 -70.035 ;
        RECT -249.885 -71.235 -249.485 -70.035 ;
        RECT -245.405 -71.235 -245.005 -70.035 ;
        RECT -240.925 -71.235 -240.525 -70.035 ;
        RECT -236.445 -71.235 -236.045 -70.035 ;
        RECT -231.965 -71.235 -231.565 -70.035 ;
        RECT -227.485 -71.235 -227.085 -70.035 ;
        RECT -223.005 -71.235 -222.605 -70.035 ;
        RECT -218.525 -71.235 -218.125 -70.035 ;
        RECT -214.045 -71.235 -213.645 -70.035 ;
        RECT -209.565 -71.235 -209.165 -70.035 ;
        RECT -205.085 -71.235 -204.685 -70.035 ;
        RECT -200.605 -71.235 -200.205 -70.035 ;
        RECT -196.125 -71.235 -195.725 -70.035 ;
        RECT -191.645 -71.235 -191.245 -70.035 ;
        RECT -186.045 -71.235 -185.645 -70.035 ;
        RECT -181.565 -71.235 -181.165 -70.035 ;
        RECT -177.085 -71.235 -176.685 -70.035 ;
        RECT -172.605 -71.235 -172.205 -70.035 ;
        RECT -168.125 -71.235 -167.725 -70.035 ;
        RECT -163.645 -71.235 -163.245 -70.035 ;
        RECT -159.165 -71.235 -158.765 -70.035 ;
        RECT -154.685 -71.235 -154.285 -70.035 ;
        RECT -150.205 -71.235 -149.805 -70.035 ;
        RECT -145.725 -71.235 -145.325 -70.035 ;
        RECT -141.245 -71.235 -140.845 -70.035 ;
        RECT -136.765 -71.235 -136.365 -70.035 ;
        RECT -132.285 -71.235 -131.885 -70.035 ;
        RECT -127.805 -71.235 -127.405 -70.035 ;
        RECT -123.325 -71.235 -122.925 -70.035 ;
        RECT -118.845 -71.235 -118.445 -70.035 ;
        RECT -114.365 -71.235 -113.965 -70.035 ;
        RECT -109.885 -71.235 -109.485 -70.035 ;
        RECT -105.405 -71.235 -105.005 -70.035 ;
        RECT -100.925 -71.235 -100.525 -70.035 ;
        RECT -96.445 -71.235 -96.045 -70.035 ;
        RECT -91.965 -71.235 -91.565 -70.035 ;
        RECT -87.485 -71.235 -87.085 -70.035 ;
        RECT -83.005 -71.235 -82.605 -70.035 ;
        RECT -78.525 -71.235 -78.125 -70.035 ;
        RECT -74.045 -71.235 -73.645 -70.035 ;
        RECT -69.565 -71.235 -69.165 -70.035 ;
        RECT -65.085 -71.235 -64.685 -70.035 ;
        RECT -60.605 -71.235 -60.205 -70.035 ;
        RECT -56.125 -71.235 -55.725 -70.035 ;
        RECT -51.645 -71.235 -51.245 -70.035 ;
        RECT -47.165 -71.235 -46.765 -70.035 ;
        RECT -42.685 -71.235 -42.285 -70.035 ;
        RECT -38.205 -71.235 -37.805 -70.035 ;
        RECT -33.725 -71.235 -33.325 -70.035 ;
        RECT -29.245 -71.235 -28.845 -70.035 ;
        RECT -24.765 -71.235 -24.365 -70.035 ;
        RECT -20.285 -71.235 -19.885 -70.035 ;
        RECT -15.805 -71.235 -15.405 -70.035 ;
        RECT -11.325 -71.235 -10.925 -70.035 ;
        RECT -6.845 -71.235 -6.445 -70.035 ;
        RECT -2.365 -71.235 -1.965 -70.035 ;
        RECT 2.115 -71.235 2.515 -70.035 ;
        RECT 6.595 -71.235 6.995 -70.035 ;
        RECT 11.075 -71.235 11.475 -70.035 ;
        RECT 15.555 -71.235 15.955 -70.035 ;
        RECT 20.035 -71.235 20.435 -70.035 ;
        RECT 24.515 -71.235 24.915 -70.035 ;
        RECT 28.995 -71.235 29.395 -70.035 ;
        RECT 33.475 -71.235 33.875 -70.035 ;
        RECT 37.955 -71.235 38.355 -70.035 ;
        RECT 42.435 -71.235 42.835 -70.035 ;
        RECT 46.915 -71.235 47.315 -70.035 ;
        RECT 51.395 -71.235 51.795 -70.035 ;
        RECT 55.875 -71.235 56.275 -70.035 ;
        RECT 60.355 -71.235 60.755 -70.035 ;
        RECT 64.835 -71.235 65.235 -70.035 ;
        RECT 69.315 -71.235 69.715 -70.035 ;
        RECT 73.795 -71.235 74.195 -70.035 ;
        RECT 78.275 -71.235 78.675 -70.035 ;
        RECT 82.755 -71.235 83.155 -70.035 ;
        RECT 87.235 -71.235 87.635 -70.035 ;
        RECT 91.715 -71.235 92.115 -70.035 ;
        RECT 96.195 -71.235 96.595 -70.035 ;
        RECT 103.305 -70.435 103.805 -41.255 ;
        RECT 102.955 -70.835 104.155 -70.435 ;
        RECT -471.645 -74.595 -471.245 -73.395 ;
        RECT -462.685 -74.595 -462.285 -73.395 ;
        RECT -453.725 -74.595 -453.325 -73.395 ;
        RECT -444.765 -74.595 -444.365 -73.395 ;
        RECT -435.805 -74.595 -435.405 -73.395 ;
        RECT -426.845 -74.595 -426.445 -73.395 ;
        RECT -417.885 -74.595 -417.485 -73.395 ;
        RECT -408.925 -74.595 -408.525 -73.395 ;
        RECT -399.965 -74.595 -399.565 -73.395 ;
        RECT -391.005 -74.595 -390.605 -73.395 ;
        RECT -382.045 -74.595 -381.645 -73.395 ;
        RECT -373.085 -74.595 -372.685 -73.395 ;
        RECT -364.125 -74.595 -363.725 -73.395 ;
        RECT -355.165 -74.595 -354.765 -73.395 ;
        RECT -346.205 -74.595 -345.805 -73.395 ;
        RECT -337.245 -74.595 -336.845 -73.395 ;
        RECT -328.285 -74.595 -327.885 -73.395 ;
        RECT -319.325 -74.595 -318.925 -73.395 ;
        RECT -310.365 -74.595 -309.965 -73.395 ;
        RECT -301.405 -74.595 -301.005 -73.395 ;
        RECT -292.445 -74.595 -292.045 -73.395 ;
        RECT -283.485 -74.595 -283.085 -73.395 ;
        RECT -274.525 -74.595 -274.125 -73.395 ;
        RECT -265.565 -74.595 -265.165 -73.395 ;
        RECT -256.605 -74.595 -256.205 -73.395 ;
        RECT -247.645 -74.595 -247.245 -73.395 ;
        RECT -238.685 -74.595 -238.285 -73.395 ;
        RECT -229.725 -74.595 -229.325 -73.395 ;
        RECT -220.765 -74.595 -220.365 -73.395 ;
        RECT -211.805 -74.595 -211.405 -73.395 ;
        RECT -202.845 -74.595 -202.445 -73.395 ;
        RECT -193.885 -74.595 -193.485 -73.395 ;
        RECT -183.805 -74.595 -183.405 -73.395 ;
        RECT -174.845 -74.595 -174.445 -73.395 ;
        RECT -165.885 -74.595 -165.485 -73.395 ;
        RECT -156.925 -74.595 -156.525 -73.395 ;
        RECT -147.965 -74.595 -147.565 -73.395 ;
        RECT -139.005 -74.595 -138.605 -73.395 ;
        RECT -130.045 -74.595 -129.645 -73.395 ;
        RECT -121.085 -74.595 -120.685 -73.395 ;
        RECT -112.125 -74.595 -111.725 -73.395 ;
        RECT -103.165 -74.595 -102.765 -73.395 ;
        RECT -94.205 -74.595 -93.805 -73.395 ;
        RECT -85.245 -74.595 -84.845 -73.395 ;
        RECT -76.285 -74.595 -75.885 -73.395 ;
        RECT -67.325 -74.595 -66.925 -73.395 ;
        RECT -58.365 -74.595 -57.965 -73.395 ;
        RECT -49.405 -74.595 -49.005 -73.395 ;
        RECT -40.445 -74.595 -40.045 -73.395 ;
        RECT -31.485 -74.595 -31.085 -73.395 ;
        RECT -22.525 -74.595 -22.125 -73.395 ;
        RECT -13.565 -74.595 -13.165 -73.395 ;
        RECT -4.605 -74.595 -4.205 -73.395 ;
        RECT 4.355 -74.595 4.755 -73.395 ;
        RECT 13.315 -74.595 13.715 -73.395 ;
        RECT 22.275 -74.595 22.675 -73.395 ;
        RECT 31.235 -74.595 31.635 -73.395 ;
        RECT 40.195 -74.595 40.595 -73.395 ;
        RECT 49.155 -74.595 49.555 -73.395 ;
        RECT 58.115 -74.595 58.515 -73.395 ;
        RECT 67.075 -74.595 67.475 -73.395 ;
        RECT 76.035 -74.595 76.435 -73.395 ;
        RECT 84.995 -74.595 85.395 -73.395 ;
        RECT 93.955 -74.595 94.355 -73.395 ;
        RECT 105.105 -73.795 105.605 -37.895 ;
        RECT 104.755 -74.195 105.955 -73.795 ;
        RECT -467.165 -77.955 -466.765 -76.755 ;
        RECT -449.245 -77.955 -448.845 -76.755 ;
        RECT -431.325 -77.955 -430.925 -76.755 ;
        RECT -413.405 -77.955 -413.005 -76.755 ;
        RECT -395.485 -77.955 -395.085 -76.755 ;
        RECT -377.565 -77.955 -377.165 -76.755 ;
        RECT -359.645 -77.955 -359.245 -76.755 ;
        RECT -341.725 -77.955 -341.325 -76.755 ;
        RECT -323.805 -77.955 -323.405 -76.755 ;
        RECT -305.885 -77.955 -305.485 -76.755 ;
        RECT -287.965 -77.955 -287.565 -76.755 ;
        RECT -270.045 -77.955 -269.645 -76.755 ;
        RECT -252.125 -77.955 -251.725 -76.755 ;
        RECT -234.205 -77.955 -233.805 -76.755 ;
        RECT -216.285 -77.955 -215.885 -76.755 ;
        RECT -198.365 -77.955 -197.965 -76.755 ;
        RECT -179.325 -77.955 -178.925 -76.755 ;
        RECT -161.405 -77.955 -161.005 -76.755 ;
        RECT -143.485 -77.955 -143.085 -76.755 ;
        RECT -125.565 -77.955 -125.165 -76.755 ;
        RECT -107.645 -77.955 -107.245 -76.755 ;
        RECT -89.725 -77.955 -89.325 -76.755 ;
        RECT -71.805 -77.955 -71.405 -76.755 ;
        RECT -53.885 -77.955 -53.485 -76.755 ;
        RECT -35.965 -77.955 -35.565 -76.755 ;
        RECT -18.045 -77.955 -17.645 -76.755 ;
        RECT -0.125 -77.955 0.275 -76.755 ;
        RECT 17.795 -77.955 18.195 -76.755 ;
        RECT 35.715 -77.955 36.115 -76.755 ;
        RECT 53.635 -77.955 54.035 -76.755 ;
        RECT 71.555 -77.955 71.955 -76.755 ;
        RECT 89.475 -77.955 89.875 -76.755 ;
        RECT 106.905 -77.155 107.405 -34.535 ;
        RECT 106.555 -77.555 107.755 -77.155 ;
        RECT -486.955 -83.235 -486.555 -81.155 ;
        RECT -458.205 -81.315 -457.805 -80.115 ;
        RECT -422.365 -81.315 -421.965 -80.115 ;
        RECT -386.525 -81.315 -386.125 -80.115 ;
        RECT -350.685 -81.315 -350.285 -80.115 ;
        RECT -314.845 -81.315 -314.445 -80.115 ;
        RECT -279.005 -81.315 -278.605 -80.115 ;
        RECT -243.165 -81.315 -242.765 -80.115 ;
        RECT -207.325 -81.315 -206.925 -80.115 ;
        RECT -170.365 -81.315 -169.965 -80.115 ;
        RECT -134.525 -81.315 -134.125 -80.115 ;
        RECT -98.685 -81.315 -98.285 -80.115 ;
        RECT -62.845 -81.315 -62.445 -80.115 ;
        RECT -27.005 -81.315 -26.605 -80.115 ;
        RECT 8.835 -81.315 9.235 -80.115 ;
        RECT 44.675 -81.315 45.075 -80.115 ;
        RECT 80.515 -81.315 80.915 -80.115 ;
        RECT 108.705 -80.515 109.205 -31.175 ;
        RECT 108.355 -80.915 109.555 -80.515 ;
        RECT -497.595 -83.765 -495.515 -83.365 ;
        RECT -440.285 -84.675 -439.885 -83.475 ;
        RECT -368.605 -84.675 -368.205 -83.475 ;
        RECT -296.925 -84.675 -296.525 -83.475 ;
        RECT -225.245 -84.675 -224.845 -83.475 ;
        RECT -152.445 -84.675 -152.045 -83.475 ;
        RECT -80.765 -84.675 -80.365 -83.475 ;
        RECT -9.085 -84.675 -8.685 -83.475 ;
        RECT 62.595 -84.675 62.995 -83.475 ;
        RECT 110.505 -83.875 111.005 -27.815 ;
        RECT 110.155 -84.275 111.355 -83.875 ;
        RECT -404.445 -88.035 -404.045 -86.835 ;
        RECT -261.085 -88.035 -260.685 -86.835 ;
        RECT -116.605 -88.035 -116.205 -86.835 ;
        RECT 26.755 -88.035 27.155 -86.835 ;
        RECT 112.305 -87.235 112.805 -24.455 ;
        RECT 111.955 -87.635 113.155 -87.235 ;
        RECT -332.765 -91.395 -332.365 -90.195 ;
        RECT -44.925 -91.395 -44.525 -90.195 ;
        RECT 114.105 -90.595 114.605 -21.095 ;
        RECT 113.755 -90.995 114.955 -90.595 ;
        RECT -188.285 -94.755 -187.885 -93.555 ;
        RECT 115.905 -93.955 116.405 -17.735 ;
        RECT 385.050 -17.820 406.710 -17.540 ;
        RECT 318.970 -18.940 346.790 -18.660 ;
        RECT 372.170 -18.940 452.630 -18.660 ;
        RECT 321.770 -19.500 325.510 -19.220 ;
        RECT 418.650 -19.500 425.750 -19.220 ;
        RECT 468.200 -19.640 469.200 -18.670 ;
        RECT 465.200 -19.780 469.200 -19.640 ;
        RECT 304.410 -20.060 331.110 -19.780 ;
        RECT 360.970 -20.060 365.830 -19.780 ;
        RECT 371.610 -20.060 385.430 -19.780 ;
        RECT 391.770 -20.060 412.310 -19.780 ;
        RECT 432.090 -20.060 436.950 -19.780 ;
        RECT 453.370 -20.060 456.550 -19.780 ;
        RECT 458.970 -20.060 469.200 -19.780 ;
        RECT 465.200 -20.200 469.200 -20.060 ;
        RECT 298.250 -20.620 313.750 -20.340 ;
        RECT 324.570 -20.620 353.510 -20.340 ;
        RECT 367.130 -20.620 376.470 -20.340 ;
        RECT 391.210 -20.620 418.470 -20.340 ;
        RECT 390.650 -21.180 402.180 -20.900 ;
        RECT 421.450 -21.180 436.950 -20.900 ;
        RECT 468.200 -21.170 469.200 -20.200 ;
        RECT 401.900 -21.460 402.180 -21.180 ;
        RECT 401.850 -21.740 433.590 -21.460 ;
        RECT 422.010 -22.860 424.070 -22.580 ;
        RECT 306.650 -23.420 319.910 -23.140 ;
        RECT 335.210 -23.420 359.670 -23.140 ;
        RECT 364.660 -23.420 406.100 -23.140 ;
        RECT 406.890 -23.420 418.470 -23.140 ;
        RECT 431.530 -23.420 435.830 -23.140 ;
        RECT 301.050 -23.980 312.630 -23.700 ;
        RECT 358.170 -23.980 361.910 -23.700 ;
        RECT 364.660 -24.260 364.940 -23.420 ;
        RECT 366.010 -23.980 391.030 -23.700 ;
        RECT 405.820 -24.260 406.100 -23.420 ;
        RECT 412.490 -23.980 419.030 -23.700 ;
        RECT 351.450 -24.540 364.940 -24.260 ;
        RECT 373.900 -24.540 396.070 -24.260 ;
        RECT 405.820 -24.540 418.470 -24.260 ;
        RECT 419.260 -24.540 438.630 -24.260 ;
        RECT 286.700 -25.240 289.200 -25.020 ;
        RECT 313.930 -25.100 322.710 -24.820 ;
        RECT 345.290 -25.100 345.670 -24.820 ;
        RECT 353.690 -25.100 359.110 -24.820 ;
        RECT 286.700 -25.380 293.200 -25.240 ;
        RECT 345.340 -25.380 345.620 -25.100 ;
        RECT 373.900 -25.380 374.180 -24.540 ;
        RECT 387.850 -25.100 392.710 -24.820 ;
        RECT 286.700 -25.660 299.190 -25.380 ;
        RECT 345.340 -25.660 374.180 -25.380 ;
        RECT 386.730 -25.660 413.430 -25.380 ;
        RECT 286.700 -25.800 293.200 -25.660 ;
        RECT 286.700 -26.020 289.200 -25.800 ;
        RECT 419.260 -25.940 419.540 -24.540 ;
        RECT 420.330 -25.100 421.830 -24.820 ;
        RECT 383.930 -26.220 419.540 -25.940 ;
        RECT 349.770 -26.780 354.630 -26.500 ;
        RECT 385.610 -26.780 447.590 -26.500 ;
        RECT 318.970 -27.340 349.590 -27.060 ;
        RECT 353.690 -27.340 358.550 -27.060 ;
        RECT 376.090 -27.340 387.110 -27.060 ;
        RECT 422.010 -27.340 426.310 -27.060 ;
        RECT 318.410 -27.900 324.390 -27.620 ;
        RECT 355.370 -27.900 365.270 -27.620 ;
        RECT 396.810 -27.900 400.550 -27.620 ;
        RECT 413.050 -27.900 435.830 -27.620 ;
        RECT 331.290 -28.460 355.190 -28.180 ;
        RECT 402.970 -28.460 427.990 -28.180 ;
        RECT 431.530 -28.460 450.390 -28.180 ;
        RECT 431.580 -28.740 431.860 -28.460 ;
        RECT 312.810 -29.020 364.940 -28.740 ;
        RECT 399.610 -29.020 431.860 -28.740 ;
        RECT 432.140 -29.020 460.470 -28.740 ;
        RECT 300.490 -30.140 314.870 -29.860 ;
        RECT 364.660 -30.420 364.940 -29.020 ;
        RECT 432.140 -29.300 432.420 -29.020 ;
        RECT 415.290 -29.580 432.420 -29.300 ;
        RECT 369.980 -30.140 388.230 -29.860 ;
        RECT 369.980 -30.420 370.260 -30.140 ;
        RECT 301.610 -30.700 317.670 -30.420 ;
        RECT 352.010 -30.700 356.870 -30.420 ;
        RECT 364.660 -30.700 370.260 -30.420 ;
        RECT 371.050 -30.700 376.470 -30.420 ;
        RECT 434.330 -30.700 448.940 -30.420 ;
        RECT 456.730 -30.700 459.910 -30.420 ;
        RECT 448.660 -30.980 448.940 -30.700 ;
        RECT 303.850 -31.260 321.030 -30.980 ;
        RECT 423.130 -31.260 437.510 -30.980 ;
        RECT 448.660 -31.260 458.790 -30.980 ;
        RECT 299.930 -31.820 331.110 -31.540 ;
        RECT 424.810 -31.820 426.870 -31.540 ;
        RECT 428.730 -31.820 439.190 -31.540 ;
        RECT 439.930 -31.820 445.350 -31.540 ;
        RECT 326.250 -32.380 332.230 -32.100 ;
        RECT 366.570 -32.380 372.550 -32.100 ;
        RECT 405.210 -32.380 422.390 -32.100 ;
        RECT 432.090 -32.380 444.790 -32.100 ;
        RECT 449.450 -32.380 457.110 -32.100 ;
        RECT 315.050 -32.940 345.110 -32.660 ;
        RECT 373.850 -32.940 387.110 -32.660 ;
        RECT 427.610 -32.940 431.350 -32.660 ;
        RECT 437.130 -32.940 461.030 -32.660 ;
        RECT 432.650 -33.500 442.550 -33.220 ;
        RECT 338.570 -34.060 365.830 -33.780 ;
        RECT 317.850 -34.620 337.830 -34.340 ;
        RECT 350.330 -34.620 352.950 -34.340 ;
        RECT 363.210 -34.620 374.230 -34.340 ;
        RECT 377.770 -34.620 382.070 -34.340 ;
        RECT 446.090 -34.620 455.430 -34.340 ;
        RECT 286.700 -35.320 289.200 -35.100 ;
        RECT 323.450 -35.180 342.870 -34.900 ;
        RECT 354.250 -35.180 359.670 -34.900 ;
        RECT 367.130 -35.180 371.990 -34.900 ;
        RECT 380.010 -35.180 389.350 -34.900 ;
        RECT 423.690 -35.180 433.030 -34.900 ;
        RECT 286.700 -35.460 293.200 -35.320 ;
        RECT 286.700 -35.740 301.990 -35.460 ;
        RECT 321.770 -35.740 348.470 -35.460 ;
        RECT 355.370 -35.740 359.110 -35.460 ;
        RECT 372.730 -35.740 390.140 -35.460 ;
        RECT 390.650 -35.740 411.750 -35.460 ;
        RECT 435.450 -35.740 437.510 -35.460 ;
        RECT 286.700 -35.880 293.200 -35.740 ;
        RECT 286.700 -36.100 289.200 -35.880 ;
        RECT 389.860 -36.020 390.140 -35.740 ;
        RECT 308.890 -36.300 325.510 -36.020 ;
        RECT 332.970 -36.300 352.950 -36.020 ;
        RECT 389.860 -36.300 447.030 -36.020 ;
        RECT 455.050 -36.300 460.470 -36.020 ;
        RECT 318.970 -36.860 337.270 -36.580 ;
        RECT 382.250 -36.860 390.470 -36.580 ;
        RECT 422.570 -36.860 443.060 -36.580 ;
        RECT 445.530 -36.860 458.230 -36.580 ;
        RECT 442.780 -37.700 443.060 -36.860 ;
        RECT 442.780 -37.980 457.670 -37.700 ;
        RECT 327.930 -38.540 372.550 -38.260 ;
        RECT 380.010 -38.540 385.430 -38.260 ;
        RECT 418.090 -38.540 423.510 -38.260 ;
        RECT 436.570 -38.540 449.830 -38.260 ;
        RECT 310.010 -39.100 323.270 -38.820 ;
        RECT 391.210 -39.100 453.750 -38.820 ;
        RECT 317.290 -39.660 326.630 -39.380 ;
        RECT 430.970 -39.660 439.140 -39.380 ;
        RECT 438.860 -39.940 439.140 -39.660 ;
        RECT 331.850 -40.220 347.350 -39.940 ;
        RECT 418.650 -40.220 424.070 -39.940 ;
        RECT 438.810 -40.220 439.190 -39.940 ;
        RECT 339.180 -40.500 339.460 -40.220 ;
        RECT 339.130 -40.780 339.510 -40.500 ;
        RECT 359.290 -40.780 370.310 -40.500 ;
        RECT 377.260 -40.780 384.310 -40.500 ;
        RECT 402.410 -40.780 415.110 -40.500 ;
        RECT 377.260 -41.620 377.540 -40.780 ;
        RECT 339.690 -41.900 377.540 -41.620 ;
        RECT 338.570 -42.460 343.430 -42.180 ;
        RECT 386.170 -42.460 402.790 -42.180 ;
        RECT 344.170 -43.020 355.190 -42.740 ;
        RECT 381.130 -43.020 390.140 -42.740 ;
        RECT 389.860 -43.300 390.140 -43.020 ;
        RECT 334.650 -43.580 349.030 -43.300 ;
        RECT 389.860 -43.580 397.750 -43.300 ;
        RECT 421.450 -43.580 432.470 -43.300 ;
        RECT 315.050 -44.140 347.350 -43.860 ;
        RECT 431.530 -44.140 454.870 -43.860 ;
        RECT 298.810 -44.700 299.190 -44.420 ;
        RECT 286.700 -45.400 289.200 -45.180 ;
        RECT 286.700 -45.540 293.200 -45.400 ;
        RECT 298.860 -45.540 299.140 -44.700 ;
        RECT 286.700 -45.820 299.140 -45.540 ;
        RECT 286.700 -45.960 293.200 -45.820 ;
        RECT 286.700 -46.180 289.200 -45.960 ;
        RECT 427.050 -46.380 459.910 -46.100 ;
        RECT 334.090 -46.940 341.190 -46.660 ;
        RECT 352.010 -46.940 360.230 -46.660 ;
        RECT 387.850 -46.940 398.870 -46.660 ;
        RECT 405.770 -46.940 417.350 -46.660 ;
        RECT 423.690 -46.940 436.390 -46.660 ;
        RECT 389.530 -47.500 393.270 -47.220 ;
        RECT 419.210 -47.500 432.470 -47.220 ;
        RECT 316.170 -48.060 322.710 -47.780 ;
        RECT 369.930 -48.060 382.070 -47.780 ;
        RECT 286.700 -55.480 289.200 -55.260 ;
        RECT 286.700 -55.620 293.200 -55.480 ;
        RECT 286.700 -55.900 306.470 -55.620 ;
        RECT 286.700 -56.040 293.200 -55.900 ;
        RECT 286.700 -56.260 289.200 -56.040 ;
        RECT 120.925 -64.165 121.925 -63.665 ;
        RECT 120.925 -67.525 121.925 -67.025 ;
        RECT 120.925 -70.885 121.925 -70.385 ;
        RECT 120.925 -74.245 121.925 -73.745 ;
        RECT 120.925 -77.605 121.925 -77.105 ;
        RECT 120.925 -80.965 121.925 -80.465 ;
        RECT 120.925 -84.325 121.925 -83.825 ;
        RECT 120.925 -87.685 121.925 -87.185 ;
        RECT 120.925 -91.045 121.925 -90.545 ;
        RECT 115.555 -94.355 116.755 -93.955 ;
        RECT 120.925 -94.405 121.925 -93.905 ;
        RECT -189.405 -98.115 -189.005 -96.915 ;
        RECT 120.925 -97.765 121.925 -97.265 ;
        RECT 135.505 -105.625 469.200 -105.525 ;
        RECT -492.150 -106.425 469.200 -105.625 ;
        RECT 135.505 -106.525 469.200 -106.425 ;
      LAYER Via3 ;
        RECT -189.345 97.675 -189.065 97.955 ;
        RECT -189.345 97.075 -189.065 97.355 ;
        RECT 121.025 97.375 121.825 97.655 ;
        RECT -188.225 94.315 -187.945 94.595 ;
        RECT -188.225 93.715 -187.945 93.995 ;
        RECT 115.715 94.015 115.995 94.295 ;
        RECT 116.315 94.015 116.595 94.295 ;
        RECT 121.025 94.015 121.825 94.295 ;
        RECT -332.705 90.955 -332.425 91.235 ;
        RECT -332.705 90.355 -332.425 90.635 ;
        RECT -44.865 90.955 -44.585 91.235 ;
        RECT -44.865 90.355 -44.585 90.635 ;
        RECT 113.915 90.655 114.195 90.935 ;
        RECT 114.515 90.655 114.795 90.935 ;
        RECT -404.385 87.595 -404.105 87.875 ;
        RECT -404.385 86.995 -404.105 87.275 ;
        RECT -261.025 87.595 -260.745 87.875 ;
        RECT -261.025 86.995 -260.745 87.275 ;
        RECT -116.545 87.595 -116.265 87.875 ;
        RECT -116.545 86.995 -116.265 87.275 ;
        RECT 26.815 87.595 27.095 87.875 ;
        RECT 26.815 86.995 27.095 87.275 ;
        RECT 112.115 87.295 112.395 87.575 ;
        RECT 112.715 87.295 112.995 87.575 ;
        RECT -440.225 84.235 -439.945 84.515 ;
        RECT -497.475 83.425 -495.635 83.705 ;
        RECT -440.225 83.635 -439.945 83.915 ;
        RECT -368.545 84.235 -368.265 84.515 ;
        RECT -368.545 83.635 -368.265 83.915 ;
        RECT -296.865 84.235 -296.585 84.515 ;
        RECT -296.865 83.635 -296.585 83.915 ;
        RECT -225.185 84.235 -224.905 84.515 ;
        RECT -225.185 83.635 -224.905 83.915 ;
        RECT -152.385 84.235 -152.105 84.515 ;
        RECT -152.385 83.635 -152.105 83.915 ;
        RECT -80.705 84.235 -80.425 84.515 ;
        RECT -80.705 83.635 -80.425 83.915 ;
        RECT -9.025 84.235 -8.745 84.515 ;
        RECT -9.025 83.635 -8.745 83.915 ;
        RECT 62.655 84.235 62.935 84.515 ;
        RECT 62.655 83.635 62.935 83.915 ;
        RECT 110.315 83.935 110.595 84.215 ;
        RECT 110.915 83.935 111.195 84.215 ;
        RECT -486.895 81.275 -486.615 83.115 ;
        RECT -458.145 80.875 -457.865 81.155 ;
        RECT -458.145 80.275 -457.865 80.555 ;
        RECT -422.305 80.875 -422.025 81.155 ;
        RECT -422.305 80.275 -422.025 80.555 ;
        RECT -386.465 80.875 -386.185 81.155 ;
        RECT -386.465 80.275 -386.185 80.555 ;
        RECT -350.625 80.875 -350.345 81.155 ;
        RECT -350.625 80.275 -350.345 80.555 ;
        RECT -314.785 80.875 -314.505 81.155 ;
        RECT -314.785 80.275 -314.505 80.555 ;
        RECT -278.945 80.875 -278.665 81.155 ;
        RECT -278.945 80.275 -278.665 80.555 ;
        RECT -243.105 80.875 -242.825 81.155 ;
        RECT -243.105 80.275 -242.825 80.555 ;
        RECT -207.265 80.875 -206.985 81.155 ;
        RECT -207.265 80.275 -206.985 80.555 ;
        RECT -170.305 80.875 -170.025 81.155 ;
        RECT -170.305 80.275 -170.025 80.555 ;
        RECT -134.465 80.875 -134.185 81.155 ;
        RECT -134.465 80.275 -134.185 80.555 ;
        RECT -98.625 80.875 -98.345 81.155 ;
        RECT -98.625 80.275 -98.345 80.555 ;
        RECT -62.785 80.875 -62.505 81.155 ;
        RECT -62.785 80.275 -62.505 80.555 ;
        RECT -26.945 80.875 -26.665 81.155 ;
        RECT -26.945 80.275 -26.665 80.555 ;
        RECT 8.895 80.875 9.175 81.155 ;
        RECT 8.895 80.275 9.175 80.555 ;
        RECT 44.735 80.875 45.015 81.155 ;
        RECT 44.735 80.275 45.015 80.555 ;
        RECT 80.575 80.875 80.855 81.155 ;
        RECT 80.575 80.275 80.855 80.555 ;
        RECT 108.515 80.575 108.795 80.855 ;
        RECT 109.115 80.575 109.395 80.855 ;
        RECT -467.105 77.515 -466.825 77.795 ;
        RECT -467.105 76.915 -466.825 77.195 ;
        RECT -449.185 77.515 -448.905 77.795 ;
        RECT -449.185 76.915 -448.905 77.195 ;
        RECT -431.265 77.515 -430.985 77.795 ;
        RECT -431.265 76.915 -430.985 77.195 ;
        RECT -413.345 77.515 -413.065 77.795 ;
        RECT -413.345 76.915 -413.065 77.195 ;
        RECT -395.425 77.515 -395.145 77.795 ;
        RECT -395.425 76.915 -395.145 77.195 ;
        RECT -377.505 77.515 -377.225 77.795 ;
        RECT -377.505 76.915 -377.225 77.195 ;
        RECT -359.585 77.515 -359.305 77.795 ;
        RECT -359.585 76.915 -359.305 77.195 ;
        RECT -341.665 77.515 -341.385 77.795 ;
        RECT -341.665 76.915 -341.385 77.195 ;
        RECT -323.745 77.515 -323.465 77.795 ;
        RECT -323.745 76.915 -323.465 77.195 ;
        RECT -305.825 77.515 -305.545 77.795 ;
        RECT -305.825 76.915 -305.545 77.195 ;
        RECT -287.905 77.515 -287.625 77.795 ;
        RECT -287.905 76.915 -287.625 77.195 ;
        RECT -269.985 77.515 -269.705 77.795 ;
        RECT -269.985 76.915 -269.705 77.195 ;
        RECT -252.065 77.515 -251.785 77.795 ;
        RECT -252.065 76.915 -251.785 77.195 ;
        RECT -234.145 77.515 -233.865 77.795 ;
        RECT -234.145 76.915 -233.865 77.195 ;
        RECT -216.225 77.515 -215.945 77.795 ;
        RECT -216.225 76.915 -215.945 77.195 ;
        RECT -198.305 77.515 -198.025 77.795 ;
        RECT -198.305 76.915 -198.025 77.195 ;
        RECT -179.265 77.515 -178.985 77.795 ;
        RECT -179.265 76.915 -178.985 77.195 ;
        RECT -161.345 77.515 -161.065 77.795 ;
        RECT -161.345 76.915 -161.065 77.195 ;
        RECT -143.425 77.515 -143.145 77.795 ;
        RECT -143.425 76.915 -143.145 77.195 ;
        RECT -125.505 77.515 -125.225 77.795 ;
        RECT -125.505 76.915 -125.225 77.195 ;
        RECT -107.585 77.515 -107.305 77.795 ;
        RECT -107.585 76.915 -107.305 77.195 ;
        RECT -89.665 77.515 -89.385 77.795 ;
        RECT -89.665 76.915 -89.385 77.195 ;
        RECT -71.745 77.515 -71.465 77.795 ;
        RECT -71.745 76.915 -71.465 77.195 ;
        RECT -53.825 77.515 -53.545 77.795 ;
        RECT -53.825 76.915 -53.545 77.195 ;
        RECT -35.905 77.515 -35.625 77.795 ;
        RECT -35.905 76.915 -35.625 77.195 ;
        RECT -17.985 77.515 -17.705 77.795 ;
        RECT -17.985 76.915 -17.705 77.195 ;
        RECT -0.065 77.515 0.215 77.795 ;
        RECT -0.065 76.915 0.215 77.195 ;
        RECT 17.855 77.515 18.135 77.795 ;
        RECT 17.855 76.915 18.135 77.195 ;
        RECT 35.775 77.515 36.055 77.795 ;
        RECT 35.775 76.915 36.055 77.195 ;
        RECT 53.695 77.515 53.975 77.795 ;
        RECT 53.695 76.915 53.975 77.195 ;
        RECT 71.615 77.515 71.895 77.795 ;
        RECT 71.615 76.915 71.895 77.195 ;
        RECT 89.535 77.515 89.815 77.795 ;
        RECT 89.535 76.915 89.815 77.195 ;
        RECT 106.715 77.215 106.995 77.495 ;
        RECT 107.315 77.215 107.595 77.495 ;
        RECT -471.585 74.155 -471.305 74.435 ;
        RECT -471.585 73.555 -471.305 73.835 ;
        RECT -462.625 74.155 -462.345 74.435 ;
        RECT -462.625 73.555 -462.345 73.835 ;
        RECT -453.665 74.155 -453.385 74.435 ;
        RECT -453.665 73.555 -453.385 73.835 ;
        RECT -444.705 74.155 -444.425 74.435 ;
        RECT -444.705 73.555 -444.425 73.835 ;
        RECT -435.745 74.155 -435.465 74.435 ;
        RECT -435.745 73.555 -435.465 73.835 ;
        RECT -426.785 74.155 -426.505 74.435 ;
        RECT -426.785 73.555 -426.505 73.835 ;
        RECT -417.825 74.155 -417.545 74.435 ;
        RECT -417.825 73.555 -417.545 73.835 ;
        RECT -408.865 74.155 -408.585 74.435 ;
        RECT -408.865 73.555 -408.585 73.835 ;
        RECT -399.905 74.155 -399.625 74.435 ;
        RECT -399.905 73.555 -399.625 73.835 ;
        RECT -390.945 74.155 -390.665 74.435 ;
        RECT -390.945 73.555 -390.665 73.835 ;
        RECT -381.985 74.155 -381.705 74.435 ;
        RECT -381.985 73.555 -381.705 73.835 ;
        RECT -373.025 74.155 -372.745 74.435 ;
        RECT -373.025 73.555 -372.745 73.835 ;
        RECT -364.065 74.155 -363.785 74.435 ;
        RECT -364.065 73.555 -363.785 73.835 ;
        RECT -355.105 74.155 -354.825 74.435 ;
        RECT -355.105 73.555 -354.825 73.835 ;
        RECT -346.145 74.155 -345.865 74.435 ;
        RECT -346.145 73.555 -345.865 73.835 ;
        RECT -337.185 74.155 -336.905 74.435 ;
        RECT -337.185 73.555 -336.905 73.835 ;
        RECT -328.225 74.155 -327.945 74.435 ;
        RECT -328.225 73.555 -327.945 73.835 ;
        RECT -319.265 74.155 -318.985 74.435 ;
        RECT -319.265 73.555 -318.985 73.835 ;
        RECT -310.305 74.155 -310.025 74.435 ;
        RECT -310.305 73.555 -310.025 73.835 ;
        RECT -301.345 74.155 -301.065 74.435 ;
        RECT -301.345 73.555 -301.065 73.835 ;
        RECT -292.385 74.155 -292.105 74.435 ;
        RECT -292.385 73.555 -292.105 73.835 ;
        RECT -283.425 74.155 -283.145 74.435 ;
        RECT -283.425 73.555 -283.145 73.835 ;
        RECT -274.465 74.155 -274.185 74.435 ;
        RECT -274.465 73.555 -274.185 73.835 ;
        RECT -265.505 74.155 -265.225 74.435 ;
        RECT -265.505 73.555 -265.225 73.835 ;
        RECT -256.545 74.155 -256.265 74.435 ;
        RECT -256.545 73.555 -256.265 73.835 ;
        RECT -247.585 74.155 -247.305 74.435 ;
        RECT -247.585 73.555 -247.305 73.835 ;
        RECT -238.625 74.155 -238.345 74.435 ;
        RECT -238.625 73.555 -238.345 73.835 ;
        RECT -229.665 74.155 -229.385 74.435 ;
        RECT -229.665 73.555 -229.385 73.835 ;
        RECT -220.705 74.155 -220.425 74.435 ;
        RECT -220.705 73.555 -220.425 73.835 ;
        RECT -211.745 74.155 -211.465 74.435 ;
        RECT -211.745 73.555 -211.465 73.835 ;
        RECT -202.785 74.155 -202.505 74.435 ;
        RECT -202.785 73.555 -202.505 73.835 ;
        RECT -193.825 74.155 -193.545 74.435 ;
        RECT -193.825 73.555 -193.545 73.835 ;
        RECT -183.745 74.155 -183.465 74.435 ;
        RECT -183.745 73.555 -183.465 73.835 ;
        RECT -174.785 74.155 -174.505 74.435 ;
        RECT -174.785 73.555 -174.505 73.835 ;
        RECT -165.825 74.155 -165.545 74.435 ;
        RECT -165.825 73.555 -165.545 73.835 ;
        RECT -156.865 74.155 -156.585 74.435 ;
        RECT -156.865 73.555 -156.585 73.835 ;
        RECT -147.905 74.155 -147.625 74.435 ;
        RECT -147.905 73.555 -147.625 73.835 ;
        RECT -138.945 74.155 -138.665 74.435 ;
        RECT -138.945 73.555 -138.665 73.835 ;
        RECT -129.985 74.155 -129.705 74.435 ;
        RECT -129.985 73.555 -129.705 73.835 ;
        RECT -121.025 74.155 -120.745 74.435 ;
        RECT -121.025 73.555 -120.745 73.835 ;
        RECT -112.065 74.155 -111.785 74.435 ;
        RECT -112.065 73.555 -111.785 73.835 ;
        RECT -103.105 74.155 -102.825 74.435 ;
        RECT -103.105 73.555 -102.825 73.835 ;
        RECT -94.145 74.155 -93.865 74.435 ;
        RECT -94.145 73.555 -93.865 73.835 ;
        RECT -85.185 74.155 -84.905 74.435 ;
        RECT -85.185 73.555 -84.905 73.835 ;
        RECT -76.225 74.155 -75.945 74.435 ;
        RECT -76.225 73.555 -75.945 73.835 ;
        RECT -67.265 74.155 -66.985 74.435 ;
        RECT -67.265 73.555 -66.985 73.835 ;
        RECT -58.305 74.155 -58.025 74.435 ;
        RECT -58.305 73.555 -58.025 73.835 ;
        RECT -49.345 74.155 -49.065 74.435 ;
        RECT -49.345 73.555 -49.065 73.835 ;
        RECT -40.385 74.155 -40.105 74.435 ;
        RECT -40.385 73.555 -40.105 73.835 ;
        RECT -31.425 74.155 -31.145 74.435 ;
        RECT -31.425 73.555 -31.145 73.835 ;
        RECT -22.465 74.155 -22.185 74.435 ;
        RECT -22.465 73.555 -22.185 73.835 ;
        RECT -13.505 74.155 -13.225 74.435 ;
        RECT -13.505 73.555 -13.225 73.835 ;
        RECT -4.545 74.155 -4.265 74.435 ;
        RECT -4.545 73.555 -4.265 73.835 ;
        RECT 4.415 74.155 4.695 74.435 ;
        RECT 4.415 73.555 4.695 73.835 ;
        RECT 13.375 74.155 13.655 74.435 ;
        RECT 13.375 73.555 13.655 73.835 ;
        RECT 22.335 74.155 22.615 74.435 ;
        RECT 22.335 73.555 22.615 73.835 ;
        RECT 31.295 74.155 31.575 74.435 ;
        RECT 31.295 73.555 31.575 73.835 ;
        RECT 40.255 74.155 40.535 74.435 ;
        RECT 40.255 73.555 40.535 73.835 ;
        RECT 49.215 74.155 49.495 74.435 ;
        RECT 49.215 73.555 49.495 73.835 ;
        RECT 58.175 74.155 58.455 74.435 ;
        RECT 58.175 73.555 58.455 73.835 ;
        RECT 67.135 74.155 67.415 74.435 ;
        RECT 67.135 73.555 67.415 73.835 ;
        RECT 76.095 74.155 76.375 74.435 ;
        RECT 76.095 73.555 76.375 73.835 ;
        RECT 85.055 74.155 85.335 74.435 ;
        RECT 85.055 73.555 85.335 73.835 ;
        RECT 94.015 74.155 94.295 74.435 ;
        RECT 94.015 73.555 94.295 73.835 ;
        RECT 104.915 73.855 105.195 74.135 ;
        RECT 105.515 73.855 105.795 74.135 ;
        RECT -473.825 70.795 -473.545 71.075 ;
        RECT -473.825 70.195 -473.545 70.475 ;
        RECT -469.345 70.795 -469.065 71.075 ;
        RECT -469.345 70.195 -469.065 70.475 ;
        RECT -464.865 70.795 -464.585 71.075 ;
        RECT -464.865 70.195 -464.585 70.475 ;
        RECT -460.385 70.795 -460.105 71.075 ;
        RECT -460.385 70.195 -460.105 70.475 ;
        RECT -455.905 70.795 -455.625 71.075 ;
        RECT -455.905 70.195 -455.625 70.475 ;
        RECT -451.425 70.795 -451.145 71.075 ;
        RECT -451.425 70.195 -451.145 70.475 ;
        RECT -446.945 70.795 -446.665 71.075 ;
        RECT -446.945 70.195 -446.665 70.475 ;
        RECT -442.465 70.795 -442.185 71.075 ;
        RECT -442.465 70.195 -442.185 70.475 ;
        RECT -437.985 70.795 -437.705 71.075 ;
        RECT -437.985 70.195 -437.705 70.475 ;
        RECT -433.505 70.795 -433.225 71.075 ;
        RECT -433.505 70.195 -433.225 70.475 ;
        RECT -429.025 70.795 -428.745 71.075 ;
        RECT -429.025 70.195 -428.745 70.475 ;
        RECT -424.545 70.795 -424.265 71.075 ;
        RECT -424.545 70.195 -424.265 70.475 ;
        RECT -420.065 70.795 -419.785 71.075 ;
        RECT -420.065 70.195 -419.785 70.475 ;
        RECT -415.585 70.795 -415.305 71.075 ;
        RECT -415.585 70.195 -415.305 70.475 ;
        RECT -411.105 70.795 -410.825 71.075 ;
        RECT -411.105 70.195 -410.825 70.475 ;
        RECT -406.625 70.795 -406.345 71.075 ;
        RECT -406.625 70.195 -406.345 70.475 ;
        RECT -402.145 70.795 -401.865 71.075 ;
        RECT -402.145 70.195 -401.865 70.475 ;
        RECT -397.665 70.795 -397.385 71.075 ;
        RECT -397.665 70.195 -397.385 70.475 ;
        RECT -393.185 70.795 -392.905 71.075 ;
        RECT -393.185 70.195 -392.905 70.475 ;
        RECT -388.705 70.795 -388.425 71.075 ;
        RECT -388.705 70.195 -388.425 70.475 ;
        RECT -384.225 70.795 -383.945 71.075 ;
        RECT -384.225 70.195 -383.945 70.475 ;
        RECT -379.745 70.795 -379.465 71.075 ;
        RECT -379.745 70.195 -379.465 70.475 ;
        RECT -375.265 70.795 -374.985 71.075 ;
        RECT -375.265 70.195 -374.985 70.475 ;
        RECT -370.785 70.795 -370.505 71.075 ;
        RECT -370.785 70.195 -370.505 70.475 ;
        RECT -366.305 70.795 -366.025 71.075 ;
        RECT -366.305 70.195 -366.025 70.475 ;
        RECT -361.825 70.795 -361.545 71.075 ;
        RECT -361.825 70.195 -361.545 70.475 ;
        RECT -357.345 70.795 -357.065 71.075 ;
        RECT -357.345 70.195 -357.065 70.475 ;
        RECT -352.865 70.795 -352.585 71.075 ;
        RECT -352.865 70.195 -352.585 70.475 ;
        RECT -348.385 70.795 -348.105 71.075 ;
        RECT -348.385 70.195 -348.105 70.475 ;
        RECT -343.905 70.795 -343.625 71.075 ;
        RECT -343.905 70.195 -343.625 70.475 ;
        RECT -339.425 70.795 -339.145 71.075 ;
        RECT -339.425 70.195 -339.145 70.475 ;
        RECT -334.945 70.795 -334.665 71.075 ;
        RECT -334.945 70.195 -334.665 70.475 ;
        RECT -330.465 70.795 -330.185 71.075 ;
        RECT -330.465 70.195 -330.185 70.475 ;
        RECT -325.985 70.795 -325.705 71.075 ;
        RECT -325.985 70.195 -325.705 70.475 ;
        RECT -321.505 70.795 -321.225 71.075 ;
        RECT -321.505 70.195 -321.225 70.475 ;
        RECT -317.025 70.795 -316.745 71.075 ;
        RECT -317.025 70.195 -316.745 70.475 ;
        RECT -312.545 70.795 -312.265 71.075 ;
        RECT -312.545 70.195 -312.265 70.475 ;
        RECT -308.065 70.795 -307.785 71.075 ;
        RECT -308.065 70.195 -307.785 70.475 ;
        RECT -303.585 70.795 -303.305 71.075 ;
        RECT -303.585 70.195 -303.305 70.475 ;
        RECT -299.105 70.795 -298.825 71.075 ;
        RECT -299.105 70.195 -298.825 70.475 ;
        RECT -294.625 70.795 -294.345 71.075 ;
        RECT -294.625 70.195 -294.345 70.475 ;
        RECT -290.145 70.795 -289.865 71.075 ;
        RECT -290.145 70.195 -289.865 70.475 ;
        RECT -285.665 70.795 -285.385 71.075 ;
        RECT -285.665 70.195 -285.385 70.475 ;
        RECT -281.185 70.795 -280.905 71.075 ;
        RECT -281.185 70.195 -280.905 70.475 ;
        RECT -276.705 70.795 -276.425 71.075 ;
        RECT -276.705 70.195 -276.425 70.475 ;
        RECT -272.225 70.795 -271.945 71.075 ;
        RECT -272.225 70.195 -271.945 70.475 ;
        RECT -267.745 70.795 -267.465 71.075 ;
        RECT -267.745 70.195 -267.465 70.475 ;
        RECT -263.265 70.795 -262.985 71.075 ;
        RECT -263.265 70.195 -262.985 70.475 ;
        RECT -258.785 70.795 -258.505 71.075 ;
        RECT -258.785 70.195 -258.505 70.475 ;
        RECT -254.305 70.795 -254.025 71.075 ;
        RECT -254.305 70.195 -254.025 70.475 ;
        RECT -249.825 70.795 -249.545 71.075 ;
        RECT -249.825 70.195 -249.545 70.475 ;
        RECT -245.345 70.795 -245.065 71.075 ;
        RECT -245.345 70.195 -245.065 70.475 ;
        RECT -240.865 70.795 -240.585 71.075 ;
        RECT -240.865 70.195 -240.585 70.475 ;
        RECT -236.385 70.795 -236.105 71.075 ;
        RECT -236.385 70.195 -236.105 70.475 ;
        RECT -231.905 70.795 -231.625 71.075 ;
        RECT -231.905 70.195 -231.625 70.475 ;
        RECT -227.425 70.795 -227.145 71.075 ;
        RECT -227.425 70.195 -227.145 70.475 ;
        RECT -222.945 70.795 -222.665 71.075 ;
        RECT -222.945 70.195 -222.665 70.475 ;
        RECT -218.465 70.795 -218.185 71.075 ;
        RECT -218.465 70.195 -218.185 70.475 ;
        RECT -213.985 70.795 -213.705 71.075 ;
        RECT -213.985 70.195 -213.705 70.475 ;
        RECT -209.505 70.795 -209.225 71.075 ;
        RECT -209.505 70.195 -209.225 70.475 ;
        RECT -205.025 70.795 -204.745 71.075 ;
        RECT -205.025 70.195 -204.745 70.475 ;
        RECT -200.545 70.795 -200.265 71.075 ;
        RECT -200.545 70.195 -200.265 70.475 ;
        RECT -196.065 70.795 -195.785 71.075 ;
        RECT -196.065 70.195 -195.785 70.475 ;
        RECT -191.585 70.795 -191.305 71.075 ;
        RECT -191.585 70.195 -191.305 70.475 ;
        RECT -185.985 70.795 -185.705 71.075 ;
        RECT -185.985 70.195 -185.705 70.475 ;
        RECT -181.505 70.795 -181.225 71.075 ;
        RECT -181.505 70.195 -181.225 70.475 ;
        RECT -177.025 70.795 -176.745 71.075 ;
        RECT -177.025 70.195 -176.745 70.475 ;
        RECT -172.545 70.795 -172.265 71.075 ;
        RECT -172.545 70.195 -172.265 70.475 ;
        RECT -168.065 70.795 -167.785 71.075 ;
        RECT -168.065 70.195 -167.785 70.475 ;
        RECT -163.585 70.795 -163.305 71.075 ;
        RECT -163.585 70.195 -163.305 70.475 ;
        RECT -159.105 70.795 -158.825 71.075 ;
        RECT -159.105 70.195 -158.825 70.475 ;
        RECT -154.625 70.795 -154.345 71.075 ;
        RECT -154.625 70.195 -154.345 70.475 ;
        RECT -150.145 70.795 -149.865 71.075 ;
        RECT -150.145 70.195 -149.865 70.475 ;
        RECT -145.665 70.795 -145.385 71.075 ;
        RECT -145.665 70.195 -145.385 70.475 ;
        RECT -141.185 70.795 -140.905 71.075 ;
        RECT -141.185 70.195 -140.905 70.475 ;
        RECT -136.705 70.795 -136.425 71.075 ;
        RECT -136.705 70.195 -136.425 70.475 ;
        RECT -132.225 70.795 -131.945 71.075 ;
        RECT -132.225 70.195 -131.945 70.475 ;
        RECT -127.745 70.795 -127.465 71.075 ;
        RECT -127.745 70.195 -127.465 70.475 ;
        RECT -123.265 70.795 -122.985 71.075 ;
        RECT -123.265 70.195 -122.985 70.475 ;
        RECT -118.785 70.795 -118.505 71.075 ;
        RECT -118.785 70.195 -118.505 70.475 ;
        RECT -114.305 70.795 -114.025 71.075 ;
        RECT -114.305 70.195 -114.025 70.475 ;
        RECT -109.825 70.795 -109.545 71.075 ;
        RECT -109.825 70.195 -109.545 70.475 ;
        RECT -105.345 70.795 -105.065 71.075 ;
        RECT -105.345 70.195 -105.065 70.475 ;
        RECT -100.865 70.795 -100.585 71.075 ;
        RECT -100.865 70.195 -100.585 70.475 ;
        RECT -96.385 70.795 -96.105 71.075 ;
        RECT -96.385 70.195 -96.105 70.475 ;
        RECT -91.905 70.795 -91.625 71.075 ;
        RECT -91.905 70.195 -91.625 70.475 ;
        RECT -87.425 70.795 -87.145 71.075 ;
        RECT -87.425 70.195 -87.145 70.475 ;
        RECT -82.945 70.795 -82.665 71.075 ;
        RECT -82.945 70.195 -82.665 70.475 ;
        RECT -78.465 70.795 -78.185 71.075 ;
        RECT -78.465 70.195 -78.185 70.475 ;
        RECT -73.985 70.795 -73.705 71.075 ;
        RECT -73.985 70.195 -73.705 70.475 ;
        RECT -69.505 70.795 -69.225 71.075 ;
        RECT -69.505 70.195 -69.225 70.475 ;
        RECT -65.025 70.795 -64.745 71.075 ;
        RECT -65.025 70.195 -64.745 70.475 ;
        RECT -60.545 70.795 -60.265 71.075 ;
        RECT -60.545 70.195 -60.265 70.475 ;
        RECT -56.065 70.795 -55.785 71.075 ;
        RECT -56.065 70.195 -55.785 70.475 ;
        RECT -51.585 70.795 -51.305 71.075 ;
        RECT -51.585 70.195 -51.305 70.475 ;
        RECT -47.105 70.795 -46.825 71.075 ;
        RECT -47.105 70.195 -46.825 70.475 ;
        RECT -42.625 70.795 -42.345 71.075 ;
        RECT -42.625 70.195 -42.345 70.475 ;
        RECT -38.145 70.795 -37.865 71.075 ;
        RECT -38.145 70.195 -37.865 70.475 ;
        RECT -33.665 70.795 -33.385 71.075 ;
        RECT -33.665 70.195 -33.385 70.475 ;
        RECT -29.185 70.795 -28.905 71.075 ;
        RECT -29.185 70.195 -28.905 70.475 ;
        RECT -24.705 70.795 -24.425 71.075 ;
        RECT -24.705 70.195 -24.425 70.475 ;
        RECT -20.225 70.795 -19.945 71.075 ;
        RECT -20.225 70.195 -19.945 70.475 ;
        RECT -15.745 70.795 -15.465 71.075 ;
        RECT -15.745 70.195 -15.465 70.475 ;
        RECT -11.265 70.795 -10.985 71.075 ;
        RECT -11.265 70.195 -10.985 70.475 ;
        RECT -6.785 70.795 -6.505 71.075 ;
        RECT -6.785 70.195 -6.505 70.475 ;
        RECT -2.305 70.795 -2.025 71.075 ;
        RECT -2.305 70.195 -2.025 70.475 ;
        RECT 2.175 70.795 2.455 71.075 ;
        RECT 2.175 70.195 2.455 70.475 ;
        RECT 6.655 70.795 6.935 71.075 ;
        RECT 6.655 70.195 6.935 70.475 ;
        RECT 11.135 70.795 11.415 71.075 ;
        RECT 11.135 70.195 11.415 70.475 ;
        RECT 15.615 70.795 15.895 71.075 ;
        RECT 15.615 70.195 15.895 70.475 ;
        RECT 20.095 70.795 20.375 71.075 ;
        RECT 20.095 70.195 20.375 70.475 ;
        RECT 24.575 70.795 24.855 71.075 ;
        RECT 24.575 70.195 24.855 70.475 ;
        RECT 29.055 70.795 29.335 71.075 ;
        RECT 29.055 70.195 29.335 70.475 ;
        RECT 33.535 70.795 33.815 71.075 ;
        RECT 33.535 70.195 33.815 70.475 ;
        RECT 38.015 70.795 38.295 71.075 ;
        RECT 38.015 70.195 38.295 70.475 ;
        RECT 42.495 70.795 42.775 71.075 ;
        RECT 42.495 70.195 42.775 70.475 ;
        RECT 46.975 70.795 47.255 71.075 ;
        RECT 46.975 70.195 47.255 70.475 ;
        RECT 51.455 70.795 51.735 71.075 ;
        RECT 51.455 70.195 51.735 70.475 ;
        RECT 55.935 70.795 56.215 71.075 ;
        RECT 55.935 70.195 56.215 70.475 ;
        RECT 60.415 70.795 60.695 71.075 ;
        RECT 60.415 70.195 60.695 70.475 ;
        RECT 64.895 70.795 65.175 71.075 ;
        RECT 64.895 70.195 65.175 70.475 ;
        RECT 69.375 70.795 69.655 71.075 ;
        RECT 69.375 70.195 69.655 70.475 ;
        RECT 73.855 70.795 74.135 71.075 ;
        RECT 73.855 70.195 74.135 70.475 ;
        RECT 78.335 70.795 78.615 71.075 ;
        RECT 78.335 70.195 78.615 70.475 ;
        RECT 82.815 70.795 83.095 71.075 ;
        RECT 82.815 70.195 83.095 70.475 ;
        RECT 87.295 70.795 87.575 71.075 ;
        RECT 87.295 70.195 87.575 70.475 ;
        RECT 91.775 70.795 92.055 71.075 ;
        RECT 91.775 70.195 92.055 70.475 ;
        RECT 96.255 70.795 96.535 71.075 ;
        RECT 96.255 70.195 96.535 70.475 ;
        RECT 103.115 70.495 103.395 70.775 ;
        RECT 103.715 70.495 103.995 70.775 ;
        RECT -474.945 67.435 -474.665 67.715 ;
        RECT -474.945 66.835 -474.665 67.115 ;
        RECT -472.705 67.435 -472.425 67.715 ;
        RECT -472.705 66.835 -472.425 67.115 ;
        RECT -470.465 67.435 -470.185 67.715 ;
        RECT -470.465 66.835 -470.185 67.115 ;
        RECT -468.225 67.435 -467.945 67.715 ;
        RECT -468.225 66.835 -467.945 67.115 ;
        RECT -465.985 67.435 -465.705 67.715 ;
        RECT -465.985 66.835 -465.705 67.115 ;
        RECT -463.745 67.435 -463.465 67.715 ;
        RECT -463.745 66.835 -463.465 67.115 ;
        RECT -461.505 67.435 -461.225 67.715 ;
        RECT -461.505 66.835 -461.225 67.115 ;
        RECT -459.265 67.435 -458.985 67.715 ;
        RECT -459.265 66.835 -458.985 67.115 ;
        RECT -457.025 67.435 -456.745 67.715 ;
        RECT -457.025 66.835 -456.745 67.115 ;
        RECT -454.785 67.435 -454.505 67.715 ;
        RECT -454.785 66.835 -454.505 67.115 ;
        RECT -452.545 67.435 -452.265 67.715 ;
        RECT -452.545 66.835 -452.265 67.115 ;
        RECT -450.305 67.435 -450.025 67.715 ;
        RECT -450.305 66.835 -450.025 67.115 ;
        RECT -448.065 67.435 -447.785 67.715 ;
        RECT -448.065 66.835 -447.785 67.115 ;
        RECT -445.825 67.435 -445.545 67.715 ;
        RECT -445.825 66.835 -445.545 67.115 ;
        RECT -443.585 67.435 -443.305 67.715 ;
        RECT -443.585 66.835 -443.305 67.115 ;
        RECT -441.345 67.435 -441.065 67.715 ;
        RECT -441.345 66.835 -441.065 67.115 ;
        RECT -439.105 67.435 -438.825 67.715 ;
        RECT -439.105 66.835 -438.825 67.115 ;
        RECT -436.865 67.435 -436.585 67.715 ;
        RECT -436.865 66.835 -436.585 67.115 ;
        RECT -434.625 67.435 -434.345 67.715 ;
        RECT -434.625 66.835 -434.345 67.115 ;
        RECT -432.385 67.435 -432.105 67.715 ;
        RECT -432.385 66.835 -432.105 67.115 ;
        RECT -430.145 67.435 -429.865 67.715 ;
        RECT -430.145 66.835 -429.865 67.115 ;
        RECT -427.905 67.435 -427.625 67.715 ;
        RECT -427.905 66.835 -427.625 67.115 ;
        RECT -425.665 67.435 -425.385 67.715 ;
        RECT -425.665 66.835 -425.385 67.115 ;
        RECT -423.425 67.435 -423.145 67.715 ;
        RECT -423.425 66.835 -423.145 67.115 ;
        RECT -421.185 67.435 -420.905 67.715 ;
        RECT -421.185 66.835 -420.905 67.115 ;
        RECT -418.945 67.435 -418.665 67.715 ;
        RECT -418.945 66.835 -418.665 67.115 ;
        RECT -416.705 67.435 -416.425 67.715 ;
        RECT -416.705 66.835 -416.425 67.115 ;
        RECT -414.465 67.435 -414.185 67.715 ;
        RECT -414.465 66.835 -414.185 67.115 ;
        RECT -412.225 67.435 -411.945 67.715 ;
        RECT -412.225 66.835 -411.945 67.115 ;
        RECT -409.985 67.435 -409.705 67.715 ;
        RECT -409.985 66.835 -409.705 67.115 ;
        RECT -407.745 67.435 -407.465 67.715 ;
        RECT -407.745 66.835 -407.465 67.115 ;
        RECT -405.505 67.435 -405.225 67.715 ;
        RECT -405.505 66.835 -405.225 67.115 ;
        RECT -403.265 67.435 -402.985 67.715 ;
        RECT -403.265 66.835 -402.985 67.115 ;
        RECT -401.025 67.435 -400.745 67.715 ;
        RECT -401.025 66.835 -400.745 67.115 ;
        RECT -398.785 67.435 -398.505 67.715 ;
        RECT -398.785 66.835 -398.505 67.115 ;
        RECT -396.545 67.435 -396.265 67.715 ;
        RECT -396.545 66.835 -396.265 67.115 ;
        RECT -394.305 67.435 -394.025 67.715 ;
        RECT -394.305 66.835 -394.025 67.115 ;
        RECT -392.065 67.435 -391.785 67.715 ;
        RECT -392.065 66.835 -391.785 67.115 ;
        RECT -389.825 67.435 -389.545 67.715 ;
        RECT -389.825 66.835 -389.545 67.115 ;
        RECT -387.585 67.435 -387.305 67.715 ;
        RECT -387.585 66.835 -387.305 67.115 ;
        RECT -385.345 67.435 -385.065 67.715 ;
        RECT -385.345 66.835 -385.065 67.115 ;
        RECT -383.105 67.435 -382.825 67.715 ;
        RECT -383.105 66.835 -382.825 67.115 ;
        RECT -380.865 67.435 -380.585 67.715 ;
        RECT -380.865 66.835 -380.585 67.115 ;
        RECT -378.625 67.435 -378.345 67.715 ;
        RECT -378.625 66.835 -378.345 67.115 ;
        RECT -376.385 67.435 -376.105 67.715 ;
        RECT -376.385 66.835 -376.105 67.115 ;
        RECT -374.145 67.435 -373.865 67.715 ;
        RECT -374.145 66.835 -373.865 67.115 ;
        RECT -371.905 67.435 -371.625 67.715 ;
        RECT -371.905 66.835 -371.625 67.115 ;
        RECT -369.665 67.435 -369.385 67.715 ;
        RECT -369.665 66.835 -369.385 67.115 ;
        RECT -367.425 67.435 -367.145 67.715 ;
        RECT -367.425 66.835 -367.145 67.115 ;
        RECT -365.185 67.435 -364.905 67.715 ;
        RECT -365.185 66.835 -364.905 67.115 ;
        RECT -362.945 67.435 -362.665 67.715 ;
        RECT -362.945 66.835 -362.665 67.115 ;
        RECT -360.705 67.435 -360.425 67.715 ;
        RECT -360.705 66.835 -360.425 67.115 ;
        RECT -358.465 67.435 -358.185 67.715 ;
        RECT -358.465 66.835 -358.185 67.115 ;
        RECT -356.225 67.435 -355.945 67.715 ;
        RECT -356.225 66.835 -355.945 67.115 ;
        RECT -353.985 67.435 -353.705 67.715 ;
        RECT -353.985 66.835 -353.705 67.115 ;
        RECT -351.745 67.435 -351.465 67.715 ;
        RECT -351.745 66.835 -351.465 67.115 ;
        RECT -349.505 67.435 -349.225 67.715 ;
        RECT -349.505 66.835 -349.225 67.115 ;
        RECT -347.265 67.435 -346.985 67.715 ;
        RECT -347.265 66.835 -346.985 67.115 ;
        RECT -345.025 67.435 -344.745 67.715 ;
        RECT -345.025 66.835 -344.745 67.115 ;
        RECT -342.785 67.435 -342.505 67.715 ;
        RECT -342.785 66.835 -342.505 67.115 ;
        RECT -340.545 67.435 -340.265 67.715 ;
        RECT -340.545 66.835 -340.265 67.115 ;
        RECT -338.305 67.435 -338.025 67.715 ;
        RECT -338.305 66.835 -338.025 67.115 ;
        RECT -336.065 67.435 -335.785 67.715 ;
        RECT -336.065 66.835 -335.785 67.115 ;
        RECT -333.825 67.435 -333.545 67.715 ;
        RECT -333.825 66.835 -333.545 67.115 ;
        RECT -331.585 67.435 -331.305 67.715 ;
        RECT -331.585 66.835 -331.305 67.115 ;
        RECT -329.345 67.435 -329.065 67.715 ;
        RECT -329.345 66.835 -329.065 67.115 ;
        RECT -327.105 67.435 -326.825 67.715 ;
        RECT -327.105 66.835 -326.825 67.115 ;
        RECT -324.865 67.435 -324.585 67.715 ;
        RECT -324.865 66.835 -324.585 67.115 ;
        RECT -322.625 67.435 -322.345 67.715 ;
        RECT -322.625 66.835 -322.345 67.115 ;
        RECT -320.385 67.435 -320.105 67.715 ;
        RECT -320.385 66.835 -320.105 67.115 ;
        RECT -318.145 67.435 -317.865 67.715 ;
        RECT -318.145 66.835 -317.865 67.115 ;
        RECT -315.905 67.435 -315.625 67.715 ;
        RECT -315.905 66.835 -315.625 67.115 ;
        RECT -313.665 67.435 -313.385 67.715 ;
        RECT -313.665 66.835 -313.385 67.115 ;
        RECT -311.425 67.435 -311.145 67.715 ;
        RECT -311.425 66.835 -311.145 67.115 ;
        RECT -309.185 67.435 -308.905 67.715 ;
        RECT -309.185 66.835 -308.905 67.115 ;
        RECT -306.945 67.435 -306.665 67.715 ;
        RECT -306.945 66.835 -306.665 67.115 ;
        RECT -304.705 67.435 -304.425 67.715 ;
        RECT -304.705 66.835 -304.425 67.115 ;
        RECT -302.465 67.435 -302.185 67.715 ;
        RECT -302.465 66.835 -302.185 67.115 ;
        RECT -300.225 67.435 -299.945 67.715 ;
        RECT -300.225 66.835 -299.945 67.115 ;
        RECT -297.985 67.435 -297.705 67.715 ;
        RECT -297.985 66.835 -297.705 67.115 ;
        RECT -295.745 67.435 -295.465 67.715 ;
        RECT -295.745 66.835 -295.465 67.115 ;
        RECT -293.505 67.435 -293.225 67.715 ;
        RECT -293.505 66.835 -293.225 67.115 ;
        RECT -291.265 67.435 -290.985 67.715 ;
        RECT -291.265 66.835 -290.985 67.115 ;
        RECT -289.025 67.435 -288.745 67.715 ;
        RECT -289.025 66.835 -288.745 67.115 ;
        RECT -286.785 67.435 -286.505 67.715 ;
        RECT -286.785 66.835 -286.505 67.115 ;
        RECT -284.545 67.435 -284.265 67.715 ;
        RECT -284.545 66.835 -284.265 67.115 ;
        RECT -282.305 67.435 -282.025 67.715 ;
        RECT -282.305 66.835 -282.025 67.115 ;
        RECT -280.065 67.435 -279.785 67.715 ;
        RECT -280.065 66.835 -279.785 67.115 ;
        RECT -277.825 67.435 -277.545 67.715 ;
        RECT -277.825 66.835 -277.545 67.115 ;
        RECT -275.585 67.435 -275.305 67.715 ;
        RECT -275.585 66.835 -275.305 67.115 ;
        RECT -273.345 67.435 -273.065 67.715 ;
        RECT -273.345 66.835 -273.065 67.115 ;
        RECT -271.105 67.435 -270.825 67.715 ;
        RECT -271.105 66.835 -270.825 67.115 ;
        RECT -268.865 67.435 -268.585 67.715 ;
        RECT -268.865 66.835 -268.585 67.115 ;
        RECT -266.625 67.435 -266.345 67.715 ;
        RECT -266.625 66.835 -266.345 67.115 ;
        RECT -264.385 67.435 -264.105 67.715 ;
        RECT -264.385 66.835 -264.105 67.115 ;
        RECT -262.145 67.435 -261.865 67.715 ;
        RECT -262.145 66.835 -261.865 67.115 ;
        RECT -259.905 67.435 -259.625 67.715 ;
        RECT -259.905 66.835 -259.625 67.115 ;
        RECT -257.665 67.435 -257.385 67.715 ;
        RECT -257.665 66.835 -257.385 67.115 ;
        RECT -255.425 67.435 -255.145 67.715 ;
        RECT -255.425 66.835 -255.145 67.115 ;
        RECT -253.185 67.435 -252.905 67.715 ;
        RECT -253.185 66.835 -252.905 67.115 ;
        RECT -250.945 67.435 -250.665 67.715 ;
        RECT -250.945 66.835 -250.665 67.115 ;
        RECT -248.705 67.435 -248.425 67.715 ;
        RECT -248.705 66.835 -248.425 67.115 ;
        RECT -246.465 67.435 -246.185 67.715 ;
        RECT -246.465 66.835 -246.185 67.115 ;
        RECT -244.225 67.435 -243.945 67.715 ;
        RECT -244.225 66.835 -243.945 67.115 ;
        RECT -241.985 67.435 -241.705 67.715 ;
        RECT -241.985 66.835 -241.705 67.115 ;
        RECT -239.745 67.435 -239.465 67.715 ;
        RECT -239.745 66.835 -239.465 67.115 ;
        RECT -237.505 67.435 -237.225 67.715 ;
        RECT -237.505 66.835 -237.225 67.115 ;
        RECT -235.265 67.435 -234.985 67.715 ;
        RECT -235.265 66.835 -234.985 67.115 ;
        RECT -233.025 67.435 -232.745 67.715 ;
        RECT -233.025 66.835 -232.745 67.115 ;
        RECT -230.785 67.435 -230.505 67.715 ;
        RECT -230.785 66.835 -230.505 67.115 ;
        RECT -228.545 67.435 -228.265 67.715 ;
        RECT -228.545 66.835 -228.265 67.115 ;
        RECT -226.305 67.435 -226.025 67.715 ;
        RECT -226.305 66.835 -226.025 67.115 ;
        RECT -224.065 67.435 -223.785 67.715 ;
        RECT -224.065 66.835 -223.785 67.115 ;
        RECT -221.825 67.435 -221.545 67.715 ;
        RECT -221.825 66.835 -221.545 67.115 ;
        RECT -219.585 67.435 -219.305 67.715 ;
        RECT -219.585 66.835 -219.305 67.115 ;
        RECT -217.345 67.435 -217.065 67.715 ;
        RECT -217.345 66.835 -217.065 67.115 ;
        RECT -215.105 67.435 -214.825 67.715 ;
        RECT -215.105 66.835 -214.825 67.115 ;
        RECT -212.865 67.435 -212.585 67.715 ;
        RECT -212.865 66.835 -212.585 67.115 ;
        RECT -210.625 67.435 -210.345 67.715 ;
        RECT -210.625 66.835 -210.345 67.115 ;
        RECT -208.385 67.435 -208.105 67.715 ;
        RECT -208.385 66.835 -208.105 67.115 ;
        RECT -206.145 67.435 -205.865 67.715 ;
        RECT -206.145 66.835 -205.865 67.115 ;
        RECT -203.905 67.435 -203.625 67.715 ;
        RECT -203.905 66.835 -203.625 67.115 ;
        RECT -201.665 67.435 -201.385 67.715 ;
        RECT -201.665 66.835 -201.385 67.115 ;
        RECT -199.425 67.435 -199.145 67.715 ;
        RECT -199.425 66.835 -199.145 67.115 ;
        RECT -197.185 67.435 -196.905 67.715 ;
        RECT -197.185 66.835 -196.905 67.115 ;
        RECT -194.945 67.435 -194.665 67.715 ;
        RECT -194.945 66.835 -194.665 67.115 ;
        RECT -192.705 67.435 -192.425 67.715 ;
        RECT -192.705 66.835 -192.425 67.115 ;
        RECT -190.465 67.435 -190.185 67.715 ;
        RECT -190.465 66.835 -190.185 67.115 ;
        RECT -187.105 67.435 -186.825 67.715 ;
        RECT -187.105 66.835 -186.825 67.115 ;
        RECT -184.865 67.435 -184.585 67.715 ;
        RECT -184.865 66.835 -184.585 67.115 ;
        RECT -182.625 67.435 -182.345 67.715 ;
        RECT -182.625 66.835 -182.345 67.115 ;
        RECT -180.385 67.435 -180.105 67.715 ;
        RECT -180.385 66.835 -180.105 67.115 ;
        RECT -178.145 67.435 -177.865 67.715 ;
        RECT -178.145 66.835 -177.865 67.115 ;
        RECT -175.905 67.435 -175.625 67.715 ;
        RECT -175.905 66.835 -175.625 67.115 ;
        RECT -173.665 67.435 -173.385 67.715 ;
        RECT -173.665 66.835 -173.385 67.115 ;
        RECT -171.425 67.435 -171.145 67.715 ;
        RECT -171.425 66.835 -171.145 67.115 ;
        RECT -169.185 67.435 -168.905 67.715 ;
        RECT -169.185 66.835 -168.905 67.115 ;
        RECT -166.945 67.435 -166.665 67.715 ;
        RECT -166.945 66.835 -166.665 67.115 ;
        RECT -164.705 67.435 -164.425 67.715 ;
        RECT -164.705 66.835 -164.425 67.115 ;
        RECT -162.465 67.435 -162.185 67.715 ;
        RECT -162.465 66.835 -162.185 67.115 ;
        RECT -160.225 67.435 -159.945 67.715 ;
        RECT -160.225 66.835 -159.945 67.115 ;
        RECT -157.985 67.435 -157.705 67.715 ;
        RECT -157.985 66.835 -157.705 67.115 ;
        RECT -155.745 67.435 -155.465 67.715 ;
        RECT -155.745 66.835 -155.465 67.115 ;
        RECT -153.505 67.435 -153.225 67.715 ;
        RECT -153.505 66.835 -153.225 67.115 ;
        RECT -151.265 67.435 -150.985 67.715 ;
        RECT -151.265 66.835 -150.985 67.115 ;
        RECT -149.025 67.435 -148.745 67.715 ;
        RECT -149.025 66.835 -148.745 67.115 ;
        RECT -146.785 67.435 -146.505 67.715 ;
        RECT -146.785 66.835 -146.505 67.115 ;
        RECT -144.545 67.435 -144.265 67.715 ;
        RECT -144.545 66.835 -144.265 67.115 ;
        RECT -142.305 67.435 -142.025 67.715 ;
        RECT -142.305 66.835 -142.025 67.115 ;
        RECT -140.065 67.435 -139.785 67.715 ;
        RECT -140.065 66.835 -139.785 67.115 ;
        RECT -137.825 67.435 -137.545 67.715 ;
        RECT -137.825 66.835 -137.545 67.115 ;
        RECT -135.585 67.435 -135.305 67.715 ;
        RECT -135.585 66.835 -135.305 67.115 ;
        RECT -133.345 67.435 -133.065 67.715 ;
        RECT -133.345 66.835 -133.065 67.115 ;
        RECT -131.105 67.435 -130.825 67.715 ;
        RECT -131.105 66.835 -130.825 67.115 ;
        RECT -128.865 67.435 -128.585 67.715 ;
        RECT -128.865 66.835 -128.585 67.115 ;
        RECT -126.625 67.435 -126.345 67.715 ;
        RECT -126.625 66.835 -126.345 67.115 ;
        RECT -124.385 67.435 -124.105 67.715 ;
        RECT -124.385 66.835 -124.105 67.115 ;
        RECT -122.145 67.435 -121.865 67.715 ;
        RECT -122.145 66.835 -121.865 67.115 ;
        RECT -119.905 67.435 -119.625 67.715 ;
        RECT -119.905 66.835 -119.625 67.115 ;
        RECT -117.665 67.435 -117.385 67.715 ;
        RECT -117.665 66.835 -117.385 67.115 ;
        RECT -115.425 67.435 -115.145 67.715 ;
        RECT -115.425 66.835 -115.145 67.115 ;
        RECT -113.185 67.435 -112.905 67.715 ;
        RECT -113.185 66.835 -112.905 67.115 ;
        RECT -110.945 67.435 -110.665 67.715 ;
        RECT -110.945 66.835 -110.665 67.115 ;
        RECT -108.705 67.435 -108.425 67.715 ;
        RECT -108.705 66.835 -108.425 67.115 ;
        RECT -106.465 67.435 -106.185 67.715 ;
        RECT -106.465 66.835 -106.185 67.115 ;
        RECT -104.225 67.435 -103.945 67.715 ;
        RECT -104.225 66.835 -103.945 67.115 ;
        RECT -101.985 67.435 -101.705 67.715 ;
        RECT -101.985 66.835 -101.705 67.115 ;
        RECT -99.745 67.435 -99.465 67.715 ;
        RECT -99.745 66.835 -99.465 67.115 ;
        RECT -97.505 67.435 -97.225 67.715 ;
        RECT -97.505 66.835 -97.225 67.115 ;
        RECT -95.265 67.435 -94.985 67.715 ;
        RECT -95.265 66.835 -94.985 67.115 ;
        RECT -93.025 67.435 -92.745 67.715 ;
        RECT -93.025 66.835 -92.745 67.115 ;
        RECT -90.785 67.435 -90.505 67.715 ;
        RECT -90.785 66.835 -90.505 67.115 ;
        RECT -88.545 67.435 -88.265 67.715 ;
        RECT -88.545 66.835 -88.265 67.115 ;
        RECT -86.305 67.435 -86.025 67.715 ;
        RECT -86.305 66.835 -86.025 67.115 ;
        RECT -84.065 67.435 -83.785 67.715 ;
        RECT -84.065 66.835 -83.785 67.115 ;
        RECT -81.825 67.435 -81.545 67.715 ;
        RECT -81.825 66.835 -81.545 67.115 ;
        RECT -79.585 67.435 -79.305 67.715 ;
        RECT -79.585 66.835 -79.305 67.115 ;
        RECT -77.345 67.435 -77.065 67.715 ;
        RECT -77.345 66.835 -77.065 67.115 ;
        RECT -75.105 67.435 -74.825 67.715 ;
        RECT -75.105 66.835 -74.825 67.115 ;
        RECT -72.865 67.435 -72.585 67.715 ;
        RECT -72.865 66.835 -72.585 67.115 ;
        RECT -70.625 67.435 -70.345 67.715 ;
        RECT -70.625 66.835 -70.345 67.115 ;
        RECT -68.385 67.435 -68.105 67.715 ;
        RECT -68.385 66.835 -68.105 67.115 ;
        RECT -66.145 67.435 -65.865 67.715 ;
        RECT -66.145 66.835 -65.865 67.115 ;
        RECT -63.905 67.435 -63.625 67.715 ;
        RECT -63.905 66.835 -63.625 67.115 ;
        RECT -61.665 67.435 -61.385 67.715 ;
        RECT -61.665 66.835 -61.385 67.115 ;
        RECT -59.425 67.435 -59.145 67.715 ;
        RECT -59.425 66.835 -59.145 67.115 ;
        RECT -57.185 67.435 -56.905 67.715 ;
        RECT -57.185 66.835 -56.905 67.115 ;
        RECT -54.945 67.435 -54.665 67.715 ;
        RECT -54.945 66.835 -54.665 67.115 ;
        RECT -52.705 67.435 -52.425 67.715 ;
        RECT -52.705 66.835 -52.425 67.115 ;
        RECT -50.465 67.435 -50.185 67.715 ;
        RECT -50.465 66.835 -50.185 67.115 ;
        RECT -48.225 67.435 -47.945 67.715 ;
        RECT -48.225 66.835 -47.945 67.115 ;
        RECT -45.985 67.435 -45.705 67.715 ;
        RECT -45.985 66.835 -45.705 67.115 ;
        RECT -43.745 67.435 -43.465 67.715 ;
        RECT -43.745 66.835 -43.465 67.115 ;
        RECT -41.505 67.435 -41.225 67.715 ;
        RECT -41.505 66.835 -41.225 67.115 ;
        RECT -39.265 67.435 -38.985 67.715 ;
        RECT -39.265 66.835 -38.985 67.115 ;
        RECT -37.025 67.435 -36.745 67.715 ;
        RECT -37.025 66.835 -36.745 67.115 ;
        RECT -34.785 67.435 -34.505 67.715 ;
        RECT -34.785 66.835 -34.505 67.115 ;
        RECT -32.545 67.435 -32.265 67.715 ;
        RECT -32.545 66.835 -32.265 67.115 ;
        RECT -30.305 67.435 -30.025 67.715 ;
        RECT -30.305 66.835 -30.025 67.115 ;
        RECT -28.065 67.435 -27.785 67.715 ;
        RECT -28.065 66.835 -27.785 67.115 ;
        RECT -25.825 67.435 -25.545 67.715 ;
        RECT -25.825 66.835 -25.545 67.115 ;
        RECT -23.585 67.435 -23.305 67.715 ;
        RECT -23.585 66.835 -23.305 67.115 ;
        RECT -21.345 67.435 -21.065 67.715 ;
        RECT -21.345 66.835 -21.065 67.115 ;
        RECT -19.105 67.435 -18.825 67.715 ;
        RECT -19.105 66.835 -18.825 67.115 ;
        RECT -16.865 67.435 -16.585 67.715 ;
        RECT -16.865 66.835 -16.585 67.115 ;
        RECT -14.625 67.435 -14.345 67.715 ;
        RECT -14.625 66.835 -14.345 67.115 ;
        RECT -12.385 67.435 -12.105 67.715 ;
        RECT -12.385 66.835 -12.105 67.115 ;
        RECT -10.145 67.435 -9.865 67.715 ;
        RECT -10.145 66.835 -9.865 67.115 ;
        RECT -7.905 67.435 -7.625 67.715 ;
        RECT -7.905 66.835 -7.625 67.115 ;
        RECT -5.665 67.435 -5.385 67.715 ;
        RECT -5.665 66.835 -5.385 67.115 ;
        RECT -3.425 67.435 -3.145 67.715 ;
        RECT -3.425 66.835 -3.145 67.115 ;
        RECT -1.185 67.435 -0.905 67.715 ;
        RECT -1.185 66.835 -0.905 67.115 ;
        RECT 1.055 67.435 1.335 67.715 ;
        RECT 1.055 66.835 1.335 67.115 ;
        RECT 3.295 67.435 3.575 67.715 ;
        RECT 3.295 66.835 3.575 67.115 ;
        RECT 5.535 67.435 5.815 67.715 ;
        RECT 5.535 66.835 5.815 67.115 ;
        RECT 7.775 67.435 8.055 67.715 ;
        RECT 7.775 66.835 8.055 67.115 ;
        RECT 10.015 67.435 10.295 67.715 ;
        RECT 10.015 66.835 10.295 67.115 ;
        RECT 12.255 67.435 12.535 67.715 ;
        RECT 12.255 66.835 12.535 67.115 ;
        RECT 14.495 67.435 14.775 67.715 ;
        RECT 14.495 66.835 14.775 67.115 ;
        RECT 16.735 67.435 17.015 67.715 ;
        RECT 16.735 66.835 17.015 67.115 ;
        RECT 18.975 67.435 19.255 67.715 ;
        RECT 18.975 66.835 19.255 67.115 ;
        RECT 21.215 67.435 21.495 67.715 ;
        RECT 21.215 66.835 21.495 67.115 ;
        RECT 23.455 67.435 23.735 67.715 ;
        RECT 23.455 66.835 23.735 67.115 ;
        RECT 25.695 67.435 25.975 67.715 ;
        RECT 25.695 66.835 25.975 67.115 ;
        RECT 27.935 67.435 28.215 67.715 ;
        RECT 27.935 66.835 28.215 67.115 ;
        RECT 30.175 67.435 30.455 67.715 ;
        RECT 30.175 66.835 30.455 67.115 ;
        RECT 32.415 67.435 32.695 67.715 ;
        RECT 32.415 66.835 32.695 67.115 ;
        RECT 34.655 67.435 34.935 67.715 ;
        RECT 34.655 66.835 34.935 67.115 ;
        RECT 36.895 67.435 37.175 67.715 ;
        RECT 36.895 66.835 37.175 67.115 ;
        RECT 39.135 67.435 39.415 67.715 ;
        RECT 39.135 66.835 39.415 67.115 ;
        RECT 41.375 67.435 41.655 67.715 ;
        RECT 41.375 66.835 41.655 67.115 ;
        RECT 43.615 67.435 43.895 67.715 ;
        RECT 43.615 66.835 43.895 67.115 ;
        RECT 45.855 67.435 46.135 67.715 ;
        RECT 45.855 66.835 46.135 67.115 ;
        RECT 48.095 67.435 48.375 67.715 ;
        RECT 48.095 66.835 48.375 67.115 ;
        RECT 50.335 67.435 50.615 67.715 ;
        RECT 50.335 66.835 50.615 67.115 ;
        RECT 52.575 67.435 52.855 67.715 ;
        RECT 52.575 66.835 52.855 67.115 ;
        RECT 54.815 67.435 55.095 67.715 ;
        RECT 54.815 66.835 55.095 67.115 ;
        RECT 57.055 67.435 57.335 67.715 ;
        RECT 57.055 66.835 57.335 67.115 ;
        RECT 59.295 67.435 59.575 67.715 ;
        RECT 59.295 66.835 59.575 67.115 ;
        RECT 61.535 67.435 61.815 67.715 ;
        RECT 61.535 66.835 61.815 67.115 ;
        RECT 63.775 67.435 64.055 67.715 ;
        RECT 63.775 66.835 64.055 67.115 ;
        RECT 66.015 67.435 66.295 67.715 ;
        RECT 66.015 66.835 66.295 67.115 ;
        RECT 68.255 67.435 68.535 67.715 ;
        RECT 68.255 66.835 68.535 67.115 ;
        RECT 70.495 67.435 70.775 67.715 ;
        RECT 70.495 66.835 70.775 67.115 ;
        RECT 72.735 67.435 73.015 67.715 ;
        RECT 72.735 66.835 73.015 67.115 ;
        RECT 74.975 67.435 75.255 67.715 ;
        RECT 74.975 66.835 75.255 67.115 ;
        RECT 77.215 67.435 77.495 67.715 ;
        RECT 77.215 66.835 77.495 67.115 ;
        RECT 79.455 67.435 79.735 67.715 ;
        RECT 79.455 66.835 79.735 67.115 ;
        RECT 81.695 67.435 81.975 67.715 ;
        RECT 81.695 66.835 81.975 67.115 ;
        RECT 83.935 67.435 84.215 67.715 ;
        RECT 83.935 66.835 84.215 67.115 ;
        RECT 86.175 67.435 86.455 67.715 ;
        RECT 86.175 66.835 86.455 67.115 ;
        RECT 88.415 67.435 88.695 67.715 ;
        RECT 88.415 66.835 88.695 67.115 ;
        RECT 90.655 67.435 90.935 67.715 ;
        RECT 90.655 66.835 90.935 67.115 ;
        RECT 92.895 67.435 93.175 67.715 ;
        RECT 92.895 66.835 93.175 67.115 ;
        RECT 95.135 67.435 95.415 67.715 ;
        RECT 95.135 66.835 95.415 67.115 ;
        RECT 97.375 67.435 97.655 67.715 ;
        RECT 97.375 66.835 97.655 67.115 ;
        RECT 101.315 67.135 101.595 67.415 ;
        RECT 101.915 67.135 102.195 67.415 ;
        RECT -474.945 44.575 -474.665 44.855 ;
        RECT -474.945 43.975 -474.665 44.255 ;
        RECT -472.705 44.575 -472.425 44.855 ;
        RECT -472.705 43.975 -472.425 44.255 ;
        RECT -470.465 44.575 -470.185 44.855 ;
        RECT -470.465 43.975 -470.185 44.255 ;
        RECT -468.225 44.575 -467.945 44.855 ;
        RECT -468.225 43.975 -467.945 44.255 ;
        RECT -465.985 44.575 -465.705 44.855 ;
        RECT -465.985 43.975 -465.705 44.255 ;
        RECT -463.745 44.575 -463.465 44.855 ;
        RECT -463.745 43.975 -463.465 44.255 ;
        RECT -461.505 44.575 -461.225 44.855 ;
        RECT -461.505 43.975 -461.225 44.255 ;
        RECT -459.265 44.575 -458.985 44.855 ;
        RECT -459.265 43.975 -458.985 44.255 ;
        RECT -457.025 44.575 -456.745 44.855 ;
        RECT -457.025 43.975 -456.745 44.255 ;
        RECT -454.785 44.575 -454.505 44.855 ;
        RECT -454.785 43.975 -454.505 44.255 ;
        RECT -452.545 44.575 -452.265 44.855 ;
        RECT -452.545 43.975 -452.265 44.255 ;
        RECT -450.305 44.575 -450.025 44.855 ;
        RECT -450.305 43.975 -450.025 44.255 ;
        RECT -448.065 44.575 -447.785 44.855 ;
        RECT -448.065 43.975 -447.785 44.255 ;
        RECT -445.825 44.575 -445.545 44.855 ;
        RECT -445.825 43.975 -445.545 44.255 ;
        RECT -443.585 44.575 -443.305 44.855 ;
        RECT -443.585 43.975 -443.305 44.255 ;
        RECT -441.345 44.575 -441.065 44.855 ;
        RECT -441.345 43.975 -441.065 44.255 ;
        RECT -439.105 44.575 -438.825 44.855 ;
        RECT -439.105 43.975 -438.825 44.255 ;
        RECT -436.865 44.575 -436.585 44.855 ;
        RECT -436.865 43.975 -436.585 44.255 ;
        RECT -434.625 44.575 -434.345 44.855 ;
        RECT -434.625 43.975 -434.345 44.255 ;
        RECT -432.385 44.575 -432.105 44.855 ;
        RECT -432.385 43.975 -432.105 44.255 ;
        RECT -430.145 44.575 -429.865 44.855 ;
        RECT -430.145 43.975 -429.865 44.255 ;
        RECT -427.905 44.575 -427.625 44.855 ;
        RECT -427.905 43.975 -427.625 44.255 ;
        RECT -425.665 44.575 -425.385 44.855 ;
        RECT -425.665 43.975 -425.385 44.255 ;
        RECT -423.425 44.575 -423.145 44.855 ;
        RECT -423.425 43.975 -423.145 44.255 ;
        RECT -421.185 44.575 -420.905 44.855 ;
        RECT -421.185 43.975 -420.905 44.255 ;
        RECT -418.945 44.575 -418.665 44.855 ;
        RECT -418.945 43.975 -418.665 44.255 ;
        RECT -416.705 44.575 -416.425 44.855 ;
        RECT -416.705 43.975 -416.425 44.255 ;
        RECT -414.465 44.575 -414.185 44.855 ;
        RECT -414.465 43.975 -414.185 44.255 ;
        RECT -412.225 44.575 -411.945 44.855 ;
        RECT -412.225 43.975 -411.945 44.255 ;
        RECT -409.985 44.575 -409.705 44.855 ;
        RECT -409.985 43.975 -409.705 44.255 ;
        RECT -407.745 44.575 -407.465 44.855 ;
        RECT -407.745 43.975 -407.465 44.255 ;
        RECT -405.505 44.575 -405.225 44.855 ;
        RECT -405.505 43.975 -405.225 44.255 ;
        RECT -403.265 44.575 -402.985 44.855 ;
        RECT -403.265 43.975 -402.985 44.255 ;
        RECT -401.025 44.575 -400.745 44.855 ;
        RECT -401.025 43.975 -400.745 44.255 ;
        RECT -398.785 44.575 -398.505 44.855 ;
        RECT -398.785 43.975 -398.505 44.255 ;
        RECT -396.545 44.575 -396.265 44.855 ;
        RECT -396.545 43.975 -396.265 44.255 ;
        RECT -394.305 44.575 -394.025 44.855 ;
        RECT -394.305 43.975 -394.025 44.255 ;
        RECT -392.065 44.575 -391.785 44.855 ;
        RECT -392.065 43.975 -391.785 44.255 ;
        RECT -389.825 44.575 -389.545 44.855 ;
        RECT -389.825 43.975 -389.545 44.255 ;
        RECT -387.585 44.575 -387.305 44.855 ;
        RECT -387.585 43.975 -387.305 44.255 ;
        RECT -385.345 44.575 -385.065 44.855 ;
        RECT -385.345 43.975 -385.065 44.255 ;
        RECT -383.105 44.575 -382.825 44.855 ;
        RECT -383.105 43.975 -382.825 44.255 ;
        RECT -380.865 44.575 -380.585 44.855 ;
        RECT -380.865 43.975 -380.585 44.255 ;
        RECT -378.625 44.575 -378.345 44.855 ;
        RECT -378.625 43.975 -378.345 44.255 ;
        RECT -376.385 44.575 -376.105 44.855 ;
        RECT -376.385 43.975 -376.105 44.255 ;
        RECT -374.145 44.575 -373.865 44.855 ;
        RECT -374.145 43.975 -373.865 44.255 ;
        RECT -371.905 44.575 -371.625 44.855 ;
        RECT -371.905 43.975 -371.625 44.255 ;
        RECT -369.665 44.575 -369.385 44.855 ;
        RECT -369.665 43.975 -369.385 44.255 ;
        RECT -367.425 44.575 -367.145 44.855 ;
        RECT -367.425 43.975 -367.145 44.255 ;
        RECT -365.185 44.575 -364.905 44.855 ;
        RECT -365.185 43.975 -364.905 44.255 ;
        RECT -362.945 44.575 -362.665 44.855 ;
        RECT -362.945 43.975 -362.665 44.255 ;
        RECT -360.705 44.575 -360.425 44.855 ;
        RECT -360.705 43.975 -360.425 44.255 ;
        RECT -358.465 44.575 -358.185 44.855 ;
        RECT -358.465 43.975 -358.185 44.255 ;
        RECT -356.225 44.575 -355.945 44.855 ;
        RECT -356.225 43.975 -355.945 44.255 ;
        RECT -353.985 44.575 -353.705 44.855 ;
        RECT -353.985 43.975 -353.705 44.255 ;
        RECT -351.745 44.575 -351.465 44.855 ;
        RECT -351.745 43.975 -351.465 44.255 ;
        RECT -349.505 44.575 -349.225 44.855 ;
        RECT -349.505 43.975 -349.225 44.255 ;
        RECT -347.265 44.575 -346.985 44.855 ;
        RECT -347.265 43.975 -346.985 44.255 ;
        RECT -345.025 44.575 -344.745 44.855 ;
        RECT -345.025 43.975 -344.745 44.255 ;
        RECT -342.785 44.575 -342.505 44.855 ;
        RECT -342.785 43.975 -342.505 44.255 ;
        RECT -340.545 44.575 -340.265 44.855 ;
        RECT -340.545 43.975 -340.265 44.255 ;
        RECT -338.305 44.575 -338.025 44.855 ;
        RECT -338.305 43.975 -338.025 44.255 ;
        RECT -336.065 44.575 -335.785 44.855 ;
        RECT -336.065 43.975 -335.785 44.255 ;
        RECT -333.825 44.575 -333.545 44.855 ;
        RECT -333.825 43.975 -333.545 44.255 ;
        RECT -331.585 44.575 -331.305 44.855 ;
        RECT -331.585 43.975 -331.305 44.255 ;
        RECT -329.345 44.575 -329.065 44.855 ;
        RECT -329.345 43.975 -329.065 44.255 ;
        RECT -327.105 44.575 -326.825 44.855 ;
        RECT -327.105 43.975 -326.825 44.255 ;
        RECT -324.865 44.575 -324.585 44.855 ;
        RECT -324.865 43.975 -324.585 44.255 ;
        RECT -322.625 44.575 -322.345 44.855 ;
        RECT -322.625 43.975 -322.345 44.255 ;
        RECT -320.385 44.575 -320.105 44.855 ;
        RECT -320.385 43.975 -320.105 44.255 ;
        RECT -318.145 44.575 -317.865 44.855 ;
        RECT -318.145 43.975 -317.865 44.255 ;
        RECT -315.905 44.575 -315.625 44.855 ;
        RECT -315.905 43.975 -315.625 44.255 ;
        RECT -313.665 44.575 -313.385 44.855 ;
        RECT -313.665 43.975 -313.385 44.255 ;
        RECT -311.425 44.575 -311.145 44.855 ;
        RECT -311.425 43.975 -311.145 44.255 ;
        RECT -309.185 44.575 -308.905 44.855 ;
        RECT -309.185 43.975 -308.905 44.255 ;
        RECT -306.945 44.575 -306.665 44.855 ;
        RECT -306.945 43.975 -306.665 44.255 ;
        RECT -304.705 44.575 -304.425 44.855 ;
        RECT -304.705 43.975 -304.425 44.255 ;
        RECT -302.465 44.575 -302.185 44.855 ;
        RECT -302.465 43.975 -302.185 44.255 ;
        RECT -300.225 44.575 -299.945 44.855 ;
        RECT -300.225 43.975 -299.945 44.255 ;
        RECT -297.985 44.575 -297.705 44.855 ;
        RECT -297.985 43.975 -297.705 44.255 ;
        RECT -295.745 44.575 -295.465 44.855 ;
        RECT -295.745 43.975 -295.465 44.255 ;
        RECT -293.505 44.575 -293.225 44.855 ;
        RECT -293.505 43.975 -293.225 44.255 ;
        RECT -291.265 44.575 -290.985 44.855 ;
        RECT -291.265 43.975 -290.985 44.255 ;
        RECT -289.025 44.575 -288.745 44.855 ;
        RECT -289.025 43.975 -288.745 44.255 ;
        RECT -286.785 44.575 -286.505 44.855 ;
        RECT -286.785 43.975 -286.505 44.255 ;
        RECT -284.545 44.575 -284.265 44.855 ;
        RECT -284.545 43.975 -284.265 44.255 ;
        RECT -282.305 44.575 -282.025 44.855 ;
        RECT -282.305 43.975 -282.025 44.255 ;
        RECT -280.065 44.575 -279.785 44.855 ;
        RECT -280.065 43.975 -279.785 44.255 ;
        RECT -277.825 44.575 -277.545 44.855 ;
        RECT -277.825 43.975 -277.545 44.255 ;
        RECT -275.585 44.575 -275.305 44.855 ;
        RECT -275.585 43.975 -275.305 44.255 ;
        RECT -273.345 44.575 -273.065 44.855 ;
        RECT -273.345 43.975 -273.065 44.255 ;
        RECT -271.105 44.575 -270.825 44.855 ;
        RECT -271.105 43.975 -270.825 44.255 ;
        RECT -268.865 44.575 -268.585 44.855 ;
        RECT -268.865 43.975 -268.585 44.255 ;
        RECT -266.625 44.575 -266.345 44.855 ;
        RECT -266.625 43.975 -266.345 44.255 ;
        RECT -264.385 44.575 -264.105 44.855 ;
        RECT -264.385 43.975 -264.105 44.255 ;
        RECT -262.145 44.575 -261.865 44.855 ;
        RECT -262.145 43.975 -261.865 44.255 ;
        RECT -259.905 44.575 -259.625 44.855 ;
        RECT -259.905 43.975 -259.625 44.255 ;
        RECT -257.665 44.575 -257.385 44.855 ;
        RECT -257.665 43.975 -257.385 44.255 ;
        RECT -255.425 44.575 -255.145 44.855 ;
        RECT -255.425 43.975 -255.145 44.255 ;
        RECT -253.185 44.575 -252.905 44.855 ;
        RECT -253.185 43.975 -252.905 44.255 ;
        RECT -250.945 44.575 -250.665 44.855 ;
        RECT -250.945 43.975 -250.665 44.255 ;
        RECT -248.705 44.575 -248.425 44.855 ;
        RECT -248.705 43.975 -248.425 44.255 ;
        RECT -246.465 44.575 -246.185 44.855 ;
        RECT -246.465 43.975 -246.185 44.255 ;
        RECT -244.225 44.575 -243.945 44.855 ;
        RECT -244.225 43.975 -243.945 44.255 ;
        RECT -241.985 44.575 -241.705 44.855 ;
        RECT -241.985 43.975 -241.705 44.255 ;
        RECT -239.745 44.575 -239.465 44.855 ;
        RECT -239.745 43.975 -239.465 44.255 ;
        RECT -237.505 44.575 -237.225 44.855 ;
        RECT -237.505 43.975 -237.225 44.255 ;
        RECT -235.265 44.575 -234.985 44.855 ;
        RECT -235.265 43.975 -234.985 44.255 ;
        RECT -233.025 44.575 -232.745 44.855 ;
        RECT -233.025 43.975 -232.745 44.255 ;
        RECT -230.785 44.575 -230.505 44.855 ;
        RECT -230.785 43.975 -230.505 44.255 ;
        RECT -228.545 44.575 -228.265 44.855 ;
        RECT -228.545 43.975 -228.265 44.255 ;
        RECT -226.305 44.575 -226.025 44.855 ;
        RECT -226.305 43.975 -226.025 44.255 ;
        RECT -224.065 44.575 -223.785 44.855 ;
        RECT -224.065 43.975 -223.785 44.255 ;
        RECT -221.825 44.575 -221.545 44.855 ;
        RECT -221.825 43.975 -221.545 44.255 ;
        RECT -219.585 44.575 -219.305 44.855 ;
        RECT -219.585 43.975 -219.305 44.255 ;
        RECT -217.345 44.575 -217.065 44.855 ;
        RECT -217.345 43.975 -217.065 44.255 ;
        RECT -215.105 44.575 -214.825 44.855 ;
        RECT -215.105 43.975 -214.825 44.255 ;
        RECT -212.865 44.575 -212.585 44.855 ;
        RECT -212.865 43.975 -212.585 44.255 ;
        RECT -210.625 44.575 -210.345 44.855 ;
        RECT -210.625 43.975 -210.345 44.255 ;
        RECT -208.385 44.575 -208.105 44.855 ;
        RECT -208.385 43.975 -208.105 44.255 ;
        RECT -206.145 44.575 -205.865 44.855 ;
        RECT -206.145 43.975 -205.865 44.255 ;
        RECT -203.905 44.575 -203.625 44.855 ;
        RECT -203.905 43.975 -203.625 44.255 ;
        RECT -201.665 44.575 -201.385 44.855 ;
        RECT -201.665 43.975 -201.385 44.255 ;
        RECT -199.425 44.575 -199.145 44.855 ;
        RECT -199.425 43.975 -199.145 44.255 ;
        RECT -197.185 44.575 -196.905 44.855 ;
        RECT -197.185 43.975 -196.905 44.255 ;
        RECT -194.945 44.575 -194.665 44.855 ;
        RECT -194.945 43.975 -194.665 44.255 ;
        RECT -192.705 44.575 -192.425 44.855 ;
        RECT -192.705 43.975 -192.425 44.255 ;
        RECT -190.465 44.575 -190.185 44.855 ;
        RECT -190.465 43.975 -190.185 44.255 ;
        RECT -187.105 44.575 -186.825 44.855 ;
        RECT -187.105 43.975 -186.825 44.255 ;
        RECT -184.865 44.575 -184.585 44.855 ;
        RECT -184.865 43.975 -184.585 44.255 ;
        RECT -182.625 44.575 -182.345 44.855 ;
        RECT -182.625 43.975 -182.345 44.255 ;
        RECT -180.385 44.575 -180.105 44.855 ;
        RECT -180.385 43.975 -180.105 44.255 ;
        RECT -178.145 44.575 -177.865 44.855 ;
        RECT -178.145 43.975 -177.865 44.255 ;
        RECT -175.905 44.575 -175.625 44.855 ;
        RECT -175.905 43.975 -175.625 44.255 ;
        RECT -173.665 44.575 -173.385 44.855 ;
        RECT -173.665 43.975 -173.385 44.255 ;
        RECT -171.425 44.575 -171.145 44.855 ;
        RECT -171.425 43.975 -171.145 44.255 ;
        RECT -169.185 44.575 -168.905 44.855 ;
        RECT -169.185 43.975 -168.905 44.255 ;
        RECT -166.945 44.575 -166.665 44.855 ;
        RECT -166.945 43.975 -166.665 44.255 ;
        RECT -164.705 44.575 -164.425 44.855 ;
        RECT -164.705 43.975 -164.425 44.255 ;
        RECT -162.465 44.575 -162.185 44.855 ;
        RECT -162.465 43.975 -162.185 44.255 ;
        RECT -160.225 44.575 -159.945 44.855 ;
        RECT -160.225 43.975 -159.945 44.255 ;
        RECT -157.985 44.575 -157.705 44.855 ;
        RECT -157.985 43.975 -157.705 44.255 ;
        RECT -155.745 44.575 -155.465 44.855 ;
        RECT -155.745 43.975 -155.465 44.255 ;
        RECT -153.505 44.575 -153.225 44.855 ;
        RECT -153.505 43.975 -153.225 44.255 ;
        RECT -151.265 44.575 -150.985 44.855 ;
        RECT -151.265 43.975 -150.985 44.255 ;
        RECT -149.025 44.575 -148.745 44.855 ;
        RECT -149.025 43.975 -148.745 44.255 ;
        RECT -146.785 44.575 -146.505 44.855 ;
        RECT -146.785 43.975 -146.505 44.255 ;
        RECT -144.545 44.575 -144.265 44.855 ;
        RECT -144.545 43.975 -144.265 44.255 ;
        RECT -142.305 44.575 -142.025 44.855 ;
        RECT -142.305 43.975 -142.025 44.255 ;
        RECT -140.065 44.575 -139.785 44.855 ;
        RECT -140.065 43.975 -139.785 44.255 ;
        RECT -137.825 44.575 -137.545 44.855 ;
        RECT -137.825 43.975 -137.545 44.255 ;
        RECT -135.585 44.575 -135.305 44.855 ;
        RECT -135.585 43.975 -135.305 44.255 ;
        RECT -133.345 44.575 -133.065 44.855 ;
        RECT -133.345 43.975 -133.065 44.255 ;
        RECT -131.105 44.575 -130.825 44.855 ;
        RECT -131.105 43.975 -130.825 44.255 ;
        RECT -128.865 44.575 -128.585 44.855 ;
        RECT -128.865 43.975 -128.585 44.255 ;
        RECT -126.625 44.575 -126.345 44.855 ;
        RECT -126.625 43.975 -126.345 44.255 ;
        RECT -124.385 44.575 -124.105 44.855 ;
        RECT -124.385 43.975 -124.105 44.255 ;
        RECT -122.145 44.575 -121.865 44.855 ;
        RECT -122.145 43.975 -121.865 44.255 ;
        RECT -119.905 44.575 -119.625 44.855 ;
        RECT -119.905 43.975 -119.625 44.255 ;
        RECT -117.665 44.575 -117.385 44.855 ;
        RECT -117.665 43.975 -117.385 44.255 ;
        RECT -115.425 44.575 -115.145 44.855 ;
        RECT -115.425 43.975 -115.145 44.255 ;
        RECT -113.185 44.575 -112.905 44.855 ;
        RECT -113.185 43.975 -112.905 44.255 ;
        RECT -110.945 44.575 -110.665 44.855 ;
        RECT -110.945 43.975 -110.665 44.255 ;
        RECT -108.705 44.575 -108.425 44.855 ;
        RECT -108.705 43.975 -108.425 44.255 ;
        RECT -106.465 44.575 -106.185 44.855 ;
        RECT -106.465 43.975 -106.185 44.255 ;
        RECT -104.225 44.575 -103.945 44.855 ;
        RECT -104.225 43.975 -103.945 44.255 ;
        RECT -101.985 44.575 -101.705 44.855 ;
        RECT -101.985 43.975 -101.705 44.255 ;
        RECT -99.745 44.575 -99.465 44.855 ;
        RECT -99.745 43.975 -99.465 44.255 ;
        RECT -97.505 44.575 -97.225 44.855 ;
        RECT -97.505 43.975 -97.225 44.255 ;
        RECT -95.265 44.575 -94.985 44.855 ;
        RECT -95.265 43.975 -94.985 44.255 ;
        RECT -93.025 44.575 -92.745 44.855 ;
        RECT -93.025 43.975 -92.745 44.255 ;
        RECT -90.785 44.575 -90.505 44.855 ;
        RECT -90.785 43.975 -90.505 44.255 ;
        RECT -88.545 44.575 -88.265 44.855 ;
        RECT -88.545 43.975 -88.265 44.255 ;
        RECT -86.305 44.575 -86.025 44.855 ;
        RECT -86.305 43.975 -86.025 44.255 ;
        RECT -84.065 44.575 -83.785 44.855 ;
        RECT -84.065 43.975 -83.785 44.255 ;
        RECT -81.825 44.575 -81.545 44.855 ;
        RECT -81.825 43.975 -81.545 44.255 ;
        RECT -79.585 44.575 -79.305 44.855 ;
        RECT -79.585 43.975 -79.305 44.255 ;
        RECT -77.345 44.575 -77.065 44.855 ;
        RECT -77.345 43.975 -77.065 44.255 ;
        RECT -75.105 44.575 -74.825 44.855 ;
        RECT -75.105 43.975 -74.825 44.255 ;
        RECT -72.865 44.575 -72.585 44.855 ;
        RECT -72.865 43.975 -72.585 44.255 ;
        RECT -70.625 44.575 -70.345 44.855 ;
        RECT -70.625 43.975 -70.345 44.255 ;
        RECT -68.385 44.575 -68.105 44.855 ;
        RECT -68.385 43.975 -68.105 44.255 ;
        RECT -66.145 44.575 -65.865 44.855 ;
        RECT -66.145 43.975 -65.865 44.255 ;
        RECT -63.905 44.575 -63.625 44.855 ;
        RECT -63.905 43.975 -63.625 44.255 ;
        RECT -61.665 44.575 -61.385 44.855 ;
        RECT -61.665 43.975 -61.385 44.255 ;
        RECT -59.425 44.575 -59.145 44.855 ;
        RECT -59.425 43.975 -59.145 44.255 ;
        RECT -57.185 44.575 -56.905 44.855 ;
        RECT -57.185 43.975 -56.905 44.255 ;
        RECT -54.945 44.575 -54.665 44.855 ;
        RECT -54.945 43.975 -54.665 44.255 ;
        RECT -52.705 44.575 -52.425 44.855 ;
        RECT -52.705 43.975 -52.425 44.255 ;
        RECT -50.465 44.575 -50.185 44.855 ;
        RECT -50.465 43.975 -50.185 44.255 ;
        RECT -48.225 44.575 -47.945 44.855 ;
        RECT -48.225 43.975 -47.945 44.255 ;
        RECT -45.985 44.575 -45.705 44.855 ;
        RECT -45.985 43.975 -45.705 44.255 ;
        RECT -43.745 44.575 -43.465 44.855 ;
        RECT -43.745 43.975 -43.465 44.255 ;
        RECT -41.505 44.575 -41.225 44.855 ;
        RECT -41.505 43.975 -41.225 44.255 ;
        RECT -39.265 44.575 -38.985 44.855 ;
        RECT -39.265 43.975 -38.985 44.255 ;
        RECT -37.025 44.575 -36.745 44.855 ;
        RECT -37.025 43.975 -36.745 44.255 ;
        RECT -34.785 44.575 -34.505 44.855 ;
        RECT -34.785 43.975 -34.505 44.255 ;
        RECT -32.545 44.575 -32.265 44.855 ;
        RECT -32.545 43.975 -32.265 44.255 ;
        RECT -30.305 44.575 -30.025 44.855 ;
        RECT -30.305 43.975 -30.025 44.255 ;
        RECT -28.065 44.575 -27.785 44.855 ;
        RECT -28.065 43.975 -27.785 44.255 ;
        RECT -25.825 44.575 -25.545 44.855 ;
        RECT -25.825 43.975 -25.545 44.255 ;
        RECT -23.585 44.575 -23.305 44.855 ;
        RECT -23.585 43.975 -23.305 44.255 ;
        RECT -21.345 44.575 -21.065 44.855 ;
        RECT -21.345 43.975 -21.065 44.255 ;
        RECT -19.105 44.575 -18.825 44.855 ;
        RECT -19.105 43.975 -18.825 44.255 ;
        RECT -16.865 44.575 -16.585 44.855 ;
        RECT -16.865 43.975 -16.585 44.255 ;
        RECT -14.625 44.575 -14.345 44.855 ;
        RECT -14.625 43.975 -14.345 44.255 ;
        RECT -12.385 44.575 -12.105 44.855 ;
        RECT -12.385 43.975 -12.105 44.255 ;
        RECT -10.145 44.575 -9.865 44.855 ;
        RECT -10.145 43.975 -9.865 44.255 ;
        RECT -7.905 44.575 -7.625 44.855 ;
        RECT -7.905 43.975 -7.625 44.255 ;
        RECT -5.665 44.575 -5.385 44.855 ;
        RECT -5.665 43.975 -5.385 44.255 ;
        RECT -3.425 44.575 -3.145 44.855 ;
        RECT -3.425 43.975 -3.145 44.255 ;
        RECT -1.185 44.575 -0.905 44.855 ;
        RECT -1.185 43.975 -0.905 44.255 ;
        RECT 1.055 44.575 1.335 44.855 ;
        RECT 1.055 43.975 1.335 44.255 ;
        RECT 3.295 44.575 3.575 44.855 ;
        RECT 3.295 43.975 3.575 44.255 ;
        RECT 5.535 44.575 5.815 44.855 ;
        RECT 5.535 43.975 5.815 44.255 ;
        RECT 7.775 44.575 8.055 44.855 ;
        RECT 7.775 43.975 8.055 44.255 ;
        RECT 10.015 44.575 10.295 44.855 ;
        RECT 10.015 43.975 10.295 44.255 ;
        RECT 12.255 44.575 12.535 44.855 ;
        RECT 12.255 43.975 12.535 44.255 ;
        RECT 14.495 44.575 14.775 44.855 ;
        RECT 14.495 43.975 14.775 44.255 ;
        RECT 16.735 44.575 17.015 44.855 ;
        RECT 16.735 43.975 17.015 44.255 ;
        RECT 18.975 44.575 19.255 44.855 ;
        RECT 18.975 43.975 19.255 44.255 ;
        RECT 21.215 44.575 21.495 44.855 ;
        RECT 21.215 43.975 21.495 44.255 ;
        RECT 23.455 44.575 23.735 44.855 ;
        RECT 23.455 43.975 23.735 44.255 ;
        RECT 25.695 44.575 25.975 44.855 ;
        RECT 25.695 43.975 25.975 44.255 ;
        RECT 27.935 44.575 28.215 44.855 ;
        RECT 27.935 43.975 28.215 44.255 ;
        RECT 30.175 44.575 30.455 44.855 ;
        RECT 30.175 43.975 30.455 44.255 ;
        RECT 32.415 44.575 32.695 44.855 ;
        RECT 32.415 43.975 32.695 44.255 ;
        RECT 34.655 44.575 34.935 44.855 ;
        RECT 34.655 43.975 34.935 44.255 ;
        RECT 36.895 44.575 37.175 44.855 ;
        RECT 36.895 43.975 37.175 44.255 ;
        RECT 39.135 44.575 39.415 44.855 ;
        RECT 39.135 43.975 39.415 44.255 ;
        RECT 41.375 44.575 41.655 44.855 ;
        RECT 41.375 43.975 41.655 44.255 ;
        RECT 43.615 44.575 43.895 44.855 ;
        RECT 43.615 43.975 43.895 44.255 ;
        RECT 45.855 44.575 46.135 44.855 ;
        RECT 45.855 43.975 46.135 44.255 ;
        RECT 48.095 44.575 48.375 44.855 ;
        RECT 48.095 43.975 48.375 44.255 ;
        RECT 50.335 44.575 50.615 44.855 ;
        RECT 50.335 43.975 50.615 44.255 ;
        RECT 52.575 44.575 52.855 44.855 ;
        RECT 52.575 43.975 52.855 44.255 ;
        RECT 54.815 44.575 55.095 44.855 ;
        RECT 54.815 43.975 55.095 44.255 ;
        RECT 57.055 44.575 57.335 44.855 ;
        RECT 57.055 43.975 57.335 44.255 ;
        RECT 59.295 44.575 59.575 44.855 ;
        RECT 59.295 43.975 59.575 44.255 ;
        RECT 61.535 44.575 61.815 44.855 ;
        RECT 61.535 43.975 61.815 44.255 ;
        RECT 63.775 44.575 64.055 44.855 ;
        RECT 63.775 43.975 64.055 44.255 ;
        RECT 66.015 44.575 66.295 44.855 ;
        RECT 66.015 43.975 66.295 44.255 ;
        RECT 68.255 44.575 68.535 44.855 ;
        RECT 68.255 43.975 68.535 44.255 ;
        RECT 70.495 44.575 70.775 44.855 ;
        RECT 70.495 43.975 70.775 44.255 ;
        RECT 72.735 44.575 73.015 44.855 ;
        RECT 72.735 43.975 73.015 44.255 ;
        RECT 74.975 44.575 75.255 44.855 ;
        RECT 74.975 43.975 75.255 44.255 ;
        RECT 77.215 44.575 77.495 44.855 ;
        RECT 77.215 43.975 77.495 44.255 ;
        RECT 79.455 44.575 79.735 44.855 ;
        RECT 79.455 43.975 79.735 44.255 ;
        RECT 81.695 44.575 81.975 44.855 ;
        RECT 81.695 43.975 81.975 44.255 ;
        RECT 83.935 44.575 84.215 44.855 ;
        RECT 83.935 43.975 84.215 44.255 ;
        RECT 86.175 44.575 86.455 44.855 ;
        RECT 86.175 43.975 86.455 44.255 ;
        RECT 88.415 44.575 88.695 44.855 ;
        RECT 88.415 43.975 88.695 44.255 ;
        RECT 90.655 44.575 90.935 44.855 ;
        RECT 90.655 43.975 90.935 44.255 ;
        RECT 92.895 44.575 93.175 44.855 ;
        RECT 92.895 43.975 93.175 44.255 ;
        RECT 95.135 44.575 95.415 44.855 ;
        RECT 95.135 43.975 95.415 44.255 ;
        RECT 97.375 44.575 97.655 44.855 ;
        RECT 97.375 43.975 97.655 44.255 ;
        RECT 101.315 44.275 101.595 44.555 ;
        RECT 101.915 44.275 102.195 44.555 ;
        RECT -473.825 41.215 -473.545 41.495 ;
        RECT -473.825 40.615 -473.545 40.895 ;
        RECT -469.345 41.215 -469.065 41.495 ;
        RECT -469.345 40.615 -469.065 40.895 ;
        RECT -464.865 41.215 -464.585 41.495 ;
        RECT -464.865 40.615 -464.585 40.895 ;
        RECT -460.385 41.215 -460.105 41.495 ;
        RECT -460.385 40.615 -460.105 40.895 ;
        RECT -455.905 41.215 -455.625 41.495 ;
        RECT -455.905 40.615 -455.625 40.895 ;
        RECT -451.425 41.215 -451.145 41.495 ;
        RECT -451.425 40.615 -451.145 40.895 ;
        RECT -446.945 41.215 -446.665 41.495 ;
        RECT -446.945 40.615 -446.665 40.895 ;
        RECT -442.465 41.215 -442.185 41.495 ;
        RECT -442.465 40.615 -442.185 40.895 ;
        RECT -437.985 41.215 -437.705 41.495 ;
        RECT -437.985 40.615 -437.705 40.895 ;
        RECT -433.505 41.215 -433.225 41.495 ;
        RECT -433.505 40.615 -433.225 40.895 ;
        RECT -429.025 41.215 -428.745 41.495 ;
        RECT -429.025 40.615 -428.745 40.895 ;
        RECT -424.545 41.215 -424.265 41.495 ;
        RECT -424.545 40.615 -424.265 40.895 ;
        RECT -420.065 41.215 -419.785 41.495 ;
        RECT -420.065 40.615 -419.785 40.895 ;
        RECT -415.585 41.215 -415.305 41.495 ;
        RECT -415.585 40.615 -415.305 40.895 ;
        RECT -411.105 41.215 -410.825 41.495 ;
        RECT -411.105 40.615 -410.825 40.895 ;
        RECT -406.625 41.215 -406.345 41.495 ;
        RECT -406.625 40.615 -406.345 40.895 ;
        RECT -402.145 41.215 -401.865 41.495 ;
        RECT -402.145 40.615 -401.865 40.895 ;
        RECT -397.665 41.215 -397.385 41.495 ;
        RECT -397.665 40.615 -397.385 40.895 ;
        RECT -393.185 41.215 -392.905 41.495 ;
        RECT -393.185 40.615 -392.905 40.895 ;
        RECT -388.705 41.215 -388.425 41.495 ;
        RECT -388.705 40.615 -388.425 40.895 ;
        RECT -384.225 41.215 -383.945 41.495 ;
        RECT -384.225 40.615 -383.945 40.895 ;
        RECT -379.745 41.215 -379.465 41.495 ;
        RECT -379.745 40.615 -379.465 40.895 ;
        RECT -375.265 41.215 -374.985 41.495 ;
        RECT -375.265 40.615 -374.985 40.895 ;
        RECT -370.785 41.215 -370.505 41.495 ;
        RECT -370.785 40.615 -370.505 40.895 ;
        RECT -366.305 41.215 -366.025 41.495 ;
        RECT -366.305 40.615 -366.025 40.895 ;
        RECT -361.825 41.215 -361.545 41.495 ;
        RECT -361.825 40.615 -361.545 40.895 ;
        RECT -357.345 41.215 -357.065 41.495 ;
        RECT -357.345 40.615 -357.065 40.895 ;
        RECT -352.865 41.215 -352.585 41.495 ;
        RECT -352.865 40.615 -352.585 40.895 ;
        RECT -348.385 41.215 -348.105 41.495 ;
        RECT -348.385 40.615 -348.105 40.895 ;
        RECT -343.905 41.215 -343.625 41.495 ;
        RECT -343.905 40.615 -343.625 40.895 ;
        RECT -339.425 41.215 -339.145 41.495 ;
        RECT -339.425 40.615 -339.145 40.895 ;
        RECT -334.945 41.215 -334.665 41.495 ;
        RECT -334.945 40.615 -334.665 40.895 ;
        RECT -330.465 41.215 -330.185 41.495 ;
        RECT -330.465 40.615 -330.185 40.895 ;
        RECT -325.985 41.215 -325.705 41.495 ;
        RECT -325.985 40.615 -325.705 40.895 ;
        RECT -321.505 41.215 -321.225 41.495 ;
        RECT -321.505 40.615 -321.225 40.895 ;
        RECT -317.025 41.215 -316.745 41.495 ;
        RECT -317.025 40.615 -316.745 40.895 ;
        RECT -312.545 41.215 -312.265 41.495 ;
        RECT -312.545 40.615 -312.265 40.895 ;
        RECT -308.065 41.215 -307.785 41.495 ;
        RECT -308.065 40.615 -307.785 40.895 ;
        RECT -303.585 41.215 -303.305 41.495 ;
        RECT -303.585 40.615 -303.305 40.895 ;
        RECT -299.105 41.215 -298.825 41.495 ;
        RECT -299.105 40.615 -298.825 40.895 ;
        RECT -294.625 41.215 -294.345 41.495 ;
        RECT -294.625 40.615 -294.345 40.895 ;
        RECT -290.145 41.215 -289.865 41.495 ;
        RECT -290.145 40.615 -289.865 40.895 ;
        RECT -285.665 41.215 -285.385 41.495 ;
        RECT -285.665 40.615 -285.385 40.895 ;
        RECT -281.185 41.215 -280.905 41.495 ;
        RECT -281.185 40.615 -280.905 40.895 ;
        RECT -276.705 41.215 -276.425 41.495 ;
        RECT -276.705 40.615 -276.425 40.895 ;
        RECT -272.225 41.215 -271.945 41.495 ;
        RECT -272.225 40.615 -271.945 40.895 ;
        RECT -267.745 41.215 -267.465 41.495 ;
        RECT -267.745 40.615 -267.465 40.895 ;
        RECT -263.265 41.215 -262.985 41.495 ;
        RECT -263.265 40.615 -262.985 40.895 ;
        RECT -258.785 41.215 -258.505 41.495 ;
        RECT -258.785 40.615 -258.505 40.895 ;
        RECT -254.305 41.215 -254.025 41.495 ;
        RECT -254.305 40.615 -254.025 40.895 ;
        RECT -249.825 41.215 -249.545 41.495 ;
        RECT -249.825 40.615 -249.545 40.895 ;
        RECT -245.345 41.215 -245.065 41.495 ;
        RECT -245.345 40.615 -245.065 40.895 ;
        RECT -240.865 41.215 -240.585 41.495 ;
        RECT -240.865 40.615 -240.585 40.895 ;
        RECT -236.385 41.215 -236.105 41.495 ;
        RECT -236.385 40.615 -236.105 40.895 ;
        RECT -231.905 41.215 -231.625 41.495 ;
        RECT -231.905 40.615 -231.625 40.895 ;
        RECT -227.425 41.215 -227.145 41.495 ;
        RECT -227.425 40.615 -227.145 40.895 ;
        RECT -222.945 41.215 -222.665 41.495 ;
        RECT -222.945 40.615 -222.665 40.895 ;
        RECT -218.465 41.215 -218.185 41.495 ;
        RECT -218.465 40.615 -218.185 40.895 ;
        RECT -213.985 41.215 -213.705 41.495 ;
        RECT -213.985 40.615 -213.705 40.895 ;
        RECT -209.505 41.215 -209.225 41.495 ;
        RECT -209.505 40.615 -209.225 40.895 ;
        RECT -205.025 41.215 -204.745 41.495 ;
        RECT -205.025 40.615 -204.745 40.895 ;
        RECT -200.545 41.215 -200.265 41.495 ;
        RECT -200.545 40.615 -200.265 40.895 ;
        RECT -196.065 41.215 -195.785 41.495 ;
        RECT -196.065 40.615 -195.785 40.895 ;
        RECT -191.585 41.215 -191.305 41.495 ;
        RECT -191.585 40.615 -191.305 40.895 ;
        RECT -185.985 41.215 -185.705 41.495 ;
        RECT -185.985 40.615 -185.705 40.895 ;
        RECT -181.505 41.215 -181.225 41.495 ;
        RECT -181.505 40.615 -181.225 40.895 ;
        RECT -177.025 41.215 -176.745 41.495 ;
        RECT -177.025 40.615 -176.745 40.895 ;
        RECT -172.545 41.215 -172.265 41.495 ;
        RECT -172.545 40.615 -172.265 40.895 ;
        RECT -168.065 41.215 -167.785 41.495 ;
        RECT -168.065 40.615 -167.785 40.895 ;
        RECT -163.585 41.215 -163.305 41.495 ;
        RECT -163.585 40.615 -163.305 40.895 ;
        RECT -159.105 41.215 -158.825 41.495 ;
        RECT -159.105 40.615 -158.825 40.895 ;
        RECT -154.625 41.215 -154.345 41.495 ;
        RECT -154.625 40.615 -154.345 40.895 ;
        RECT -150.145 41.215 -149.865 41.495 ;
        RECT -150.145 40.615 -149.865 40.895 ;
        RECT -145.665 41.215 -145.385 41.495 ;
        RECT -145.665 40.615 -145.385 40.895 ;
        RECT -141.185 41.215 -140.905 41.495 ;
        RECT -141.185 40.615 -140.905 40.895 ;
        RECT -136.705 41.215 -136.425 41.495 ;
        RECT -136.705 40.615 -136.425 40.895 ;
        RECT -132.225 41.215 -131.945 41.495 ;
        RECT -132.225 40.615 -131.945 40.895 ;
        RECT -127.745 41.215 -127.465 41.495 ;
        RECT -127.745 40.615 -127.465 40.895 ;
        RECT -123.265 41.215 -122.985 41.495 ;
        RECT -123.265 40.615 -122.985 40.895 ;
        RECT -118.785 41.215 -118.505 41.495 ;
        RECT -118.785 40.615 -118.505 40.895 ;
        RECT -114.305 41.215 -114.025 41.495 ;
        RECT -114.305 40.615 -114.025 40.895 ;
        RECT -109.825 41.215 -109.545 41.495 ;
        RECT -109.825 40.615 -109.545 40.895 ;
        RECT -105.345 41.215 -105.065 41.495 ;
        RECT -105.345 40.615 -105.065 40.895 ;
        RECT -100.865 41.215 -100.585 41.495 ;
        RECT -100.865 40.615 -100.585 40.895 ;
        RECT -96.385 41.215 -96.105 41.495 ;
        RECT -96.385 40.615 -96.105 40.895 ;
        RECT -91.905 41.215 -91.625 41.495 ;
        RECT -91.905 40.615 -91.625 40.895 ;
        RECT -87.425 41.215 -87.145 41.495 ;
        RECT -87.425 40.615 -87.145 40.895 ;
        RECT -82.945 41.215 -82.665 41.495 ;
        RECT -82.945 40.615 -82.665 40.895 ;
        RECT -78.465 41.215 -78.185 41.495 ;
        RECT -78.465 40.615 -78.185 40.895 ;
        RECT -73.985 41.215 -73.705 41.495 ;
        RECT -73.985 40.615 -73.705 40.895 ;
        RECT -69.505 41.215 -69.225 41.495 ;
        RECT -69.505 40.615 -69.225 40.895 ;
        RECT -65.025 41.215 -64.745 41.495 ;
        RECT -65.025 40.615 -64.745 40.895 ;
        RECT -60.545 41.215 -60.265 41.495 ;
        RECT -60.545 40.615 -60.265 40.895 ;
        RECT -56.065 41.215 -55.785 41.495 ;
        RECT -56.065 40.615 -55.785 40.895 ;
        RECT -51.585 41.215 -51.305 41.495 ;
        RECT -51.585 40.615 -51.305 40.895 ;
        RECT -47.105 41.215 -46.825 41.495 ;
        RECT -47.105 40.615 -46.825 40.895 ;
        RECT -42.625 41.215 -42.345 41.495 ;
        RECT -42.625 40.615 -42.345 40.895 ;
        RECT -38.145 41.215 -37.865 41.495 ;
        RECT -38.145 40.615 -37.865 40.895 ;
        RECT -33.665 41.215 -33.385 41.495 ;
        RECT -33.665 40.615 -33.385 40.895 ;
        RECT -29.185 41.215 -28.905 41.495 ;
        RECT -29.185 40.615 -28.905 40.895 ;
        RECT -24.705 41.215 -24.425 41.495 ;
        RECT -24.705 40.615 -24.425 40.895 ;
        RECT -20.225 41.215 -19.945 41.495 ;
        RECT -20.225 40.615 -19.945 40.895 ;
        RECT -15.745 41.215 -15.465 41.495 ;
        RECT -15.745 40.615 -15.465 40.895 ;
        RECT -11.265 41.215 -10.985 41.495 ;
        RECT -11.265 40.615 -10.985 40.895 ;
        RECT -6.785 41.215 -6.505 41.495 ;
        RECT -6.785 40.615 -6.505 40.895 ;
        RECT -2.305 41.215 -2.025 41.495 ;
        RECT -2.305 40.615 -2.025 40.895 ;
        RECT 2.175 41.215 2.455 41.495 ;
        RECT 2.175 40.615 2.455 40.895 ;
        RECT 6.655 41.215 6.935 41.495 ;
        RECT 6.655 40.615 6.935 40.895 ;
        RECT 11.135 41.215 11.415 41.495 ;
        RECT 11.135 40.615 11.415 40.895 ;
        RECT 15.615 41.215 15.895 41.495 ;
        RECT 15.615 40.615 15.895 40.895 ;
        RECT 20.095 41.215 20.375 41.495 ;
        RECT 20.095 40.615 20.375 40.895 ;
        RECT 24.575 41.215 24.855 41.495 ;
        RECT 24.575 40.615 24.855 40.895 ;
        RECT 29.055 41.215 29.335 41.495 ;
        RECT 29.055 40.615 29.335 40.895 ;
        RECT 33.535 41.215 33.815 41.495 ;
        RECT 33.535 40.615 33.815 40.895 ;
        RECT 38.015 41.215 38.295 41.495 ;
        RECT 38.015 40.615 38.295 40.895 ;
        RECT 42.495 41.215 42.775 41.495 ;
        RECT 42.495 40.615 42.775 40.895 ;
        RECT 46.975 41.215 47.255 41.495 ;
        RECT 46.975 40.615 47.255 40.895 ;
        RECT 51.455 41.215 51.735 41.495 ;
        RECT 51.455 40.615 51.735 40.895 ;
        RECT 55.935 41.215 56.215 41.495 ;
        RECT 55.935 40.615 56.215 40.895 ;
        RECT 60.415 41.215 60.695 41.495 ;
        RECT 60.415 40.615 60.695 40.895 ;
        RECT 64.895 41.215 65.175 41.495 ;
        RECT 64.895 40.615 65.175 40.895 ;
        RECT 69.375 41.215 69.655 41.495 ;
        RECT 69.375 40.615 69.655 40.895 ;
        RECT 73.855 41.215 74.135 41.495 ;
        RECT 73.855 40.615 74.135 40.895 ;
        RECT 78.335 41.215 78.615 41.495 ;
        RECT 78.335 40.615 78.615 40.895 ;
        RECT 82.815 41.215 83.095 41.495 ;
        RECT 82.815 40.615 83.095 40.895 ;
        RECT 87.295 41.215 87.575 41.495 ;
        RECT 87.295 40.615 87.575 40.895 ;
        RECT 91.775 41.215 92.055 41.495 ;
        RECT 91.775 40.615 92.055 40.895 ;
        RECT 96.255 41.215 96.535 41.495 ;
        RECT 96.255 40.615 96.535 40.895 ;
        RECT 103.115 40.915 103.395 41.195 ;
        RECT 103.715 40.915 103.995 41.195 ;
        RECT -471.585 37.855 -471.305 38.135 ;
        RECT -471.585 37.255 -471.305 37.535 ;
        RECT -462.625 37.855 -462.345 38.135 ;
        RECT -462.625 37.255 -462.345 37.535 ;
        RECT -453.665 37.855 -453.385 38.135 ;
        RECT -453.665 37.255 -453.385 37.535 ;
        RECT -444.705 37.855 -444.425 38.135 ;
        RECT -444.705 37.255 -444.425 37.535 ;
        RECT -435.745 37.855 -435.465 38.135 ;
        RECT -435.745 37.255 -435.465 37.535 ;
        RECT -426.785 37.855 -426.505 38.135 ;
        RECT -426.785 37.255 -426.505 37.535 ;
        RECT -417.825 37.855 -417.545 38.135 ;
        RECT -417.825 37.255 -417.545 37.535 ;
        RECT -408.865 37.855 -408.585 38.135 ;
        RECT -408.865 37.255 -408.585 37.535 ;
        RECT -399.905 37.855 -399.625 38.135 ;
        RECT -399.905 37.255 -399.625 37.535 ;
        RECT -390.945 37.855 -390.665 38.135 ;
        RECT -390.945 37.255 -390.665 37.535 ;
        RECT -381.985 37.855 -381.705 38.135 ;
        RECT -381.985 37.255 -381.705 37.535 ;
        RECT -373.025 37.855 -372.745 38.135 ;
        RECT -373.025 37.255 -372.745 37.535 ;
        RECT -364.065 37.855 -363.785 38.135 ;
        RECT -364.065 37.255 -363.785 37.535 ;
        RECT -355.105 37.855 -354.825 38.135 ;
        RECT -355.105 37.255 -354.825 37.535 ;
        RECT -346.145 37.855 -345.865 38.135 ;
        RECT -346.145 37.255 -345.865 37.535 ;
        RECT -337.185 37.855 -336.905 38.135 ;
        RECT -337.185 37.255 -336.905 37.535 ;
        RECT -328.225 37.855 -327.945 38.135 ;
        RECT -328.225 37.255 -327.945 37.535 ;
        RECT -319.265 37.855 -318.985 38.135 ;
        RECT -319.265 37.255 -318.985 37.535 ;
        RECT -310.305 37.855 -310.025 38.135 ;
        RECT -310.305 37.255 -310.025 37.535 ;
        RECT -301.345 37.855 -301.065 38.135 ;
        RECT -301.345 37.255 -301.065 37.535 ;
        RECT -292.385 37.855 -292.105 38.135 ;
        RECT -292.385 37.255 -292.105 37.535 ;
        RECT -283.425 37.855 -283.145 38.135 ;
        RECT -283.425 37.255 -283.145 37.535 ;
        RECT -274.465 37.855 -274.185 38.135 ;
        RECT -274.465 37.255 -274.185 37.535 ;
        RECT -265.505 37.855 -265.225 38.135 ;
        RECT -265.505 37.255 -265.225 37.535 ;
        RECT -256.545 37.855 -256.265 38.135 ;
        RECT -256.545 37.255 -256.265 37.535 ;
        RECT -247.585 37.855 -247.305 38.135 ;
        RECT -247.585 37.255 -247.305 37.535 ;
        RECT -238.625 37.855 -238.345 38.135 ;
        RECT -238.625 37.255 -238.345 37.535 ;
        RECT -229.665 37.855 -229.385 38.135 ;
        RECT -229.665 37.255 -229.385 37.535 ;
        RECT -220.705 37.855 -220.425 38.135 ;
        RECT -220.705 37.255 -220.425 37.535 ;
        RECT -211.745 37.855 -211.465 38.135 ;
        RECT -211.745 37.255 -211.465 37.535 ;
        RECT -202.785 37.855 -202.505 38.135 ;
        RECT -202.785 37.255 -202.505 37.535 ;
        RECT -193.825 37.855 -193.545 38.135 ;
        RECT -193.825 37.255 -193.545 37.535 ;
        RECT -183.745 37.855 -183.465 38.135 ;
        RECT -183.745 37.255 -183.465 37.535 ;
        RECT -174.785 37.855 -174.505 38.135 ;
        RECT -174.785 37.255 -174.505 37.535 ;
        RECT -165.825 37.855 -165.545 38.135 ;
        RECT -165.825 37.255 -165.545 37.535 ;
        RECT -156.865 37.855 -156.585 38.135 ;
        RECT -156.865 37.255 -156.585 37.535 ;
        RECT -147.905 37.855 -147.625 38.135 ;
        RECT -147.905 37.255 -147.625 37.535 ;
        RECT -138.945 37.855 -138.665 38.135 ;
        RECT -138.945 37.255 -138.665 37.535 ;
        RECT -129.985 37.855 -129.705 38.135 ;
        RECT -129.985 37.255 -129.705 37.535 ;
        RECT -121.025 37.855 -120.745 38.135 ;
        RECT -121.025 37.255 -120.745 37.535 ;
        RECT -112.065 37.855 -111.785 38.135 ;
        RECT -112.065 37.255 -111.785 37.535 ;
        RECT -103.105 37.855 -102.825 38.135 ;
        RECT -103.105 37.255 -102.825 37.535 ;
        RECT -94.145 37.855 -93.865 38.135 ;
        RECT -94.145 37.255 -93.865 37.535 ;
        RECT -85.185 37.855 -84.905 38.135 ;
        RECT -85.185 37.255 -84.905 37.535 ;
        RECT -76.225 37.855 -75.945 38.135 ;
        RECT -76.225 37.255 -75.945 37.535 ;
        RECT -67.265 37.855 -66.985 38.135 ;
        RECT -67.265 37.255 -66.985 37.535 ;
        RECT -58.305 37.855 -58.025 38.135 ;
        RECT -58.305 37.255 -58.025 37.535 ;
        RECT -49.345 37.855 -49.065 38.135 ;
        RECT -49.345 37.255 -49.065 37.535 ;
        RECT -40.385 37.855 -40.105 38.135 ;
        RECT -40.385 37.255 -40.105 37.535 ;
        RECT -31.425 37.855 -31.145 38.135 ;
        RECT -31.425 37.255 -31.145 37.535 ;
        RECT -22.465 37.855 -22.185 38.135 ;
        RECT -22.465 37.255 -22.185 37.535 ;
        RECT -13.505 37.855 -13.225 38.135 ;
        RECT -13.505 37.255 -13.225 37.535 ;
        RECT -4.545 37.855 -4.265 38.135 ;
        RECT -4.545 37.255 -4.265 37.535 ;
        RECT 4.415 37.855 4.695 38.135 ;
        RECT 4.415 37.255 4.695 37.535 ;
        RECT 13.375 37.855 13.655 38.135 ;
        RECT 13.375 37.255 13.655 37.535 ;
        RECT 22.335 37.855 22.615 38.135 ;
        RECT 22.335 37.255 22.615 37.535 ;
        RECT 31.295 37.855 31.575 38.135 ;
        RECT 31.295 37.255 31.575 37.535 ;
        RECT 40.255 37.855 40.535 38.135 ;
        RECT 40.255 37.255 40.535 37.535 ;
        RECT 49.215 37.855 49.495 38.135 ;
        RECT 49.215 37.255 49.495 37.535 ;
        RECT 58.175 37.855 58.455 38.135 ;
        RECT 58.175 37.255 58.455 37.535 ;
        RECT 67.135 37.855 67.415 38.135 ;
        RECT 67.135 37.255 67.415 37.535 ;
        RECT 76.095 37.855 76.375 38.135 ;
        RECT 76.095 37.255 76.375 37.535 ;
        RECT 85.055 37.855 85.335 38.135 ;
        RECT 85.055 37.255 85.335 37.535 ;
        RECT 94.015 37.855 94.295 38.135 ;
        RECT 94.015 37.255 94.295 37.535 ;
        RECT 104.915 37.555 105.195 37.835 ;
        RECT 105.515 37.555 105.795 37.835 ;
        RECT -467.105 34.495 -466.825 34.775 ;
        RECT -467.105 33.895 -466.825 34.175 ;
        RECT -449.185 34.495 -448.905 34.775 ;
        RECT -449.185 33.895 -448.905 34.175 ;
        RECT -431.265 34.495 -430.985 34.775 ;
        RECT -431.265 33.895 -430.985 34.175 ;
        RECT -413.345 34.495 -413.065 34.775 ;
        RECT -413.345 33.895 -413.065 34.175 ;
        RECT -395.425 34.495 -395.145 34.775 ;
        RECT -395.425 33.895 -395.145 34.175 ;
        RECT -377.505 34.495 -377.225 34.775 ;
        RECT -377.505 33.895 -377.225 34.175 ;
        RECT -359.585 34.495 -359.305 34.775 ;
        RECT -359.585 33.895 -359.305 34.175 ;
        RECT -341.665 34.495 -341.385 34.775 ;
        RECT -341.665 33.895 -341.385 34.175 ;
        RECT -323.745 34.495 -323.465 34.775 ;
        RECT -323.745 33.895 -323.465 34.175 ;
        RECT -305.825 34.495 -305.545 34.775 ;
        RECT -305.825 33.895 -305.545 34.175 ;
        RECT -287.905 34.495 -287.625 34.775 ;
        RECT -287.905 33.895 -287.625 34.175 ;
        RECT -269.985 34.495 -269.705 34.775 ;
        RECT -269.985 33.895 -269.705 34.175 ;
        RECT -252.065 34.495 -251.785 34.775 ;
        RECT -252.065 33.895 -251.785 34.175 ;
        RECT -234.145 34.495 -233.865 34.775 ;
        RECT -234.145 33.895 -233.865 34.175 ;
        RECT -216.225 34.495 -215.945 34.775 ;
        RECT -216.225 33.895 -215.945 34.175 ;
        RECT -198.305 34.495 -198.025 34.775 ;
        RECT -198.305 33.895 -198.025 34.175 ;
        RECT -179.265 34.495 -178.985 34.775 ;
        RECT -179.265 33.895 -178.985 34.175 ;
        RECT -161.345 34.495 -161.065 34.775 ;
        RECT -161.345 33.895 -161.065 34.175 ;
        RECT -143.425 34.495 -143.145 34.775 ;
        RECT -143.425 33.895 -143.145 34.175 ;
        RECT -125.505 34.495 -125.225 34.775 ;
        RECT -125.505 33.895 -125.225 34.175 ;
        RECT -107.585 34.495 -107.305 34.775 ;
        RECT -107.585 33.895 -107.305 34.175 ;
        RECT -89.665 34.495 -89.385 34.775 ;
        RECT -89.665 33.895 -89.385 34.175 ;
        RECT -71.745 34.495 -71.465 34.775 ;
        RECT -71.745 33.895 -71.465 34.175 ;
        RECT -53.825 34.495 -53.545 34.775 ;
        RECT -53.825 33.895 -53.545 34.175 ;
        RECT -35.905 34.495 -35.625 34.775 ;
        RECT -35.905 33.895 -35.625 34.175 ;
        RECT -17.985 34.495 -17.705 34.775 ;
        RECT -17.985 33.895 -17.705 34.175 ;
        RECT -0.065 34.495 0.215 34.775 ;
        RECT -0.065 33.895 0.215 34.175 ;
        RECT 17.855 34.495 18.135 34.775 ;
        RECT 17.855 33.895 18.135 34.175 ;
        RECT 35.775 34.495 36.055 34.775 ;
        RECT 35.775 33.895 36.055 34.175 ;
        RECT 53.695 34.495 53.975 34.775 ;
        RECT 53.695 33.895 53.975 34.175 ;
        RECT 71.615 34.495 71.895 34.775 ;
        RECT 71.615 33.895 71.895 34.175 ;
        RECT 89.535 34.495 89.815 34.775 ;
        RECT 89.535 33.895 89.815 34.175 ;
        RECT 106.715 34.195 106.995 34.475 ;
        RECT 107.315 34.195 107.595 34.475 ;
        RECT -458.145 31.135 -457.865 31.415 ;
        RECT -458.145 30.535 -457.865 30.815 ;
        RECT -422.305 31.135 -422.025 31.415 ;
        RECT -422.305 30.535 -422.025 30.815 ;
        RECT -386.465 31.135 -386.185 31.415 ;
        RECT -386.465 30.535 -386.185 30.815 ;
        RECT -350.625 31.135 -350.345 31.415 ;
        RECT -350.625 30.535 -350.345 30.815 ;
        RECT -314.785 31.135 -314.505 31.415 ;
        RECT -314.785 30.535 -314.505 30.815 ;
        RECT -278.945 31.135 -278.665 31.415 ;
        RECT -278.945 30.535 -278.665 30.815 ;
        RECT -243.105 31.135 -242.825 31.415 ;
        RECT -243.105 30.535 -242.825 30.815 ;
        RECT -207.265 31.135 -206.985 31.415 ;
        RECT -207.265 30.535 -206.985 30.815 ;
        RECT -170.305 31.135 -170.025 31.415 ;
        RECT -170.305 30.535 -170.025 30.815 ;
        RECT -134.465 31.135 -134.185 31.415 ;
        RECT -134.465 30.535 -134.185 30.815 ;
        RECT -98.625 31.135 -98.345 31.415 ;
        RECT -98.625 30.535 -98.345 30.815 ;
        RECT -62.785 31.135 -62.505 31.415 ;
        RECT -62.785 30.535 -62.505 30.815 ;
        RECT -26.945 31.135 -26.665 31.415 ;
        RECT -26.945 30.535 -26.665 30.815 ;
        RECT 8.895 31.135 9.175 31.415 ;
        RECT 8.895 30.535 9.175 30.815 ;
        RECT 44.735 31.135 45.015 31.415 ;
        RECT 44.735 30.535 45.015 30.815 ;
        RECT 80.575 31.135 80.855 31.415 ;
        RECT 80.575 30.535 80.855 30.815 ;
        RECT 108.515 30.835 108.795 31.115 ;
        RECT 109.115 30.835 109.395 31.115 ;
        RECT -440.225 27.775 -439.945 28.055 ;
        RECT -440.225 27.175 -439.945 27.455 ;
        RECT -368.545 27.775 -368.265 28.055 ;
        RECT -368.545 27.175 -368.265 27.455 ;
        RECT -296.865 27.775 -296.585 28.055 ;
        RECT -296.865 27.175 -296.585 27.455 ;
        RECT -225.185 27.775 -224.905 28.055 ;
        RECT -225.185 27.175 -224.905 27.455 ;
        RECT -152.385 27.775 -152.105 28.055 ;
        RECT -152.385 27.175 -152.105 27.455 ;
        RECT -80.705 27.775 -80.425 28.055 ;
        RECT -80.705 27.175 -80.425 27.455 ;
        RECT -9.025 27.775 -8.745 28.055 ;
        RECT -9.025 27.175 -8.745 27.455 ;
        RECT 62.655 27.775 62.935 28.055 ;
        RECT 62.655 27.175 62.935 27.455 ;
        RECT 110.315 27.475 110.595 27.755 ;
        RECT 110.915 27.475 111.195 27.755 ;
        RECT -404.385 24.415 -404.105 24.695 ;
        RECT -404.385 23.815 -404.105 24.095 ;
        RECT -261.025 24.415 -260.745 24.695 ;
        RECT -261.025 23.815 -260.745 24.095 ;
        RECT -116.545 24.415 -116.265 24.695 ;
        RECT -116.545 23.815 -116.265 24.095 ;
        RECT 26.815 24.415 27.095 24.695 ;
        RECT 26.815 23.815 27.095 24.095 ;
        RECT 112.115 24.115 112.395 24.395 ;
        RECT 112.715 24.115 112.995 24.395 ;
        RECT -332.705 21.055 -332.425 21.335 ;
        RECT -332.705 20.455 -332.425 20.735 ;
        RECT -44.865 21.055 -44.585 21.335 ;
        RECT -44.865 20.455 -44.585 20.735 ;
        RECT 113.915 20.755 114.195 21.035 ;
        RECT 114.515 20.755 114.795 21.035 ;
        RECT -188.225 17.695 -187.945 17.975 ;
        RECT 121.025 90.655 121.825 90.935 ;
        RECT 121.025 87.295 121.825 87.575 ;
        RECT 121.025 83.935 121.825 84.215 ;
        RECT 121.025 80.575 121.825 80.855 ;
        RECT 121.025 77.215 121.825 77.495 ;
        RECT 121.025 73.855 121.825 74.135 ;
        RECT 121.025 70.495 121.825 70.775 ;
        RECT 121.025 67.135 121.825 67.415 ;
        RECT 121.025 63.775 121.825 64.055 ;
        RECT -188.225 17.095 -187.945 17.375 ;
        RECT 115.715 17.395 115.995 17.675 ;
        RECT 116.315 17.395 116.595 17.675 ;
        RECT -189.345 14.335 -189.065 14.615 ;
        RECT -189.345 13.735 -189.065 14.015 ;
        RECT 236.000 5.040 237.320 7.400 ;
        RECT 236.000 2.040 237.320 4.400 ;
        RECT 389.580 0.660 389.860 0.940 ;
        RECT 230.020 -5.725 232.380 -4.405 ;
        RECT 233.020 -5.725 235.380 -4.405 ;
        RECT 389.020 -6.060 389.300 -5.780 ;
        RECT -189.345 -14.015 -189.065 -13.735 ;
        RECT 389.580 -13.900 389.860 -13.620 ;
        RECT -189.345 -14.615 -189.065 -14.335 ;
        RECT 389.020 -14.460 389.300 -14.180 ;
        RECT 385.660 -15.020 385.940 -14.740 ;
        RECT -188.225 -17.375 -187.945 -17.095 ;
        RECT 385.660 -17.260 385.940 -16.980 ;
        RECT -188.225 -17.975 -187.945 -17.695 ;
        RECT 115.715 -17.675 115.995 -17.395 ;
        RECT 116.315 -17.675 116.595 -17.395 ;
        RECT -332.705 -20.735 -332.425 -20.455 ;
        RECT -332.705 -21.335 -332.425 -21.055 ;
        RECT -44.865 -20.735 -44.585 -20.455 ;
        RECT -44.865 -21.335 -44.585 -21.055 ;
        RECT 113.915 -21.035 114.195 -20.755 ;
        RECT 114.515 -21.035 114.795 -20.755 ;
        RECT -404.385 -24.095 -404.105 -23.815 ;
        RECT -404.385 -24.695 -404.105 -24.415 ;
        RECT -261.025 -24.095 -260.745 -23.815 ;
        RECT -261.025 -24.695 -260.745 -24.415 ;
        RECT -116.545 -24.095 -116.265 -23.815 ;
        RECT -116.545 -24.695 -116.265 -24.415 ;
        RECT 26.815 -24.095 27.095 -23.815 ;
        RECT 26.815 -24.695 27.095 -24.415 ;
        RECT 112.115 -24.395 112.395 -24.115 ;
        RECT 112.715 -24.395 112.995 -24.115 ;
        RECT -440.225 -27.455 -439.945 -27.175 ;
        RECT -440.225 -28.055 -439.945 -27.775 ;
        RECT -368.545 -27.455 -368.265 -27.175 ;
        RECT -368.545 -28.055 -368.265 -27.775 ;
        RECT -296.865 -27.455 -296.585 -27.175 ;
        RECT -296.865 -28.055 -296.585 -27.775 ;
        RECT -225.185 -27.455 -224.905 -27.175 ;
        RECT -225.185 -28.055 -224.905 -27.775 ;
        RECT -152.385 -27.455 -152.105 -27.175 ;
        RECT -152.385 -28.055 -152.105 -27.775 ;
        RECT -80.705 -27.455 -80.425 -27.175 ;
        RECT -80.705 -28.055 -80.425 -27.775 ;
        RECT -9.025 -27.455 -8.745 -27.175 ;
        RECT -9.025 -28.055 -8.745 -27.775 ;
        RECT 62.655 -27.455 62.935 -27.175 ;
        RECT 62.655 -28.055 62.935 -27.775 ;
        RECT 110.315 -27.755 110.595 -27.475 ;
        RECT 110.915 -27.755 111.195 -27.475 ;
        RECT -458.145 -30.815 -457.865 -30.535 ;
        RECT -458.145 -31.415 -457.865 -31.135 ;
        RECT -422.305 -30.815 -422.025 -30.535 ;
        RECT -422.305 -31.415 -422.025 -31.135 ;
        RECT -386.465 -30.815 -386.185 -30.535 ;
        RECT -386.465 -31.415 -386.185 -31.135 ;
        RECT -350.625 -30.815 -350.345 -30.535 ;
        RECT -350.625 -31.415 -350.345 -31.135 ;
        RECT -314.785 -30.815 -314.505 -30.535 ;
        RECT -314.785 -31.415 -314.505 -31.135 ;
        RECT -278.945 -30.815 -278.665 -30.535 ;
        RECT -278.945 -31.415 -278.665 -31.135 ;
        RECT -243.105 -30.815 -242.825 -30.535 ;
        RECT -243.105 -31.415 -242.825 -31.135 ;
        RECT -207.265 -30.815 -206.985 -30.535 ;
        RECT -207.265 -31.415 -206.985 -31.135 ;
        RECT -170.305 -30.815 -170.025 -30.535 ;
        RECT -170.305 -31.415 -170.025 -31.135 ;
        RECT -134.465 -30.815 -134.185 -30.535 ;
        RECT -134.465 -31.415 -134.185 -31.135 ;
        RECT -98.625 -30.815 -98.345 -30.535 ;
        RECT -98.625 -31.415 -98.345 -31.135 ;
        RECT -62.785 -30.815 -62.505 -30.535 ;
        RECT -62.785 -31.415 -62.505 -31.135 ;
        RECT -26.945 -30.815 -26.665 -30.535 ;
        RECT -26.945 -31.415 -26.665 -31.135 ;
        RECT 8.895 -30.815 9.175 -30.535 ;
        RECT 8.895 -31.415 9.175 -31.135 ;
        RECT 44.735 -30.815 45.015 -30.535 ;
        RECT 44.735 -31.415 45.015 -31.135 ;
        RECT 80.575 -30.815 80.855 -30.535 ;
        RECT 80.575 -31.415 80.855 -31.135 ;
        RECT 108.515 -31.115 108.795 -30.835 ;
        RECT 109.115 -31.115 109.395 -30.835 ;
        RECT -467.105 -34.175 -466.825 -33.895 ;
        RECT -467.105 -34.775 -466.825 -34.495 ;
        RECT -449.185 -34.175 -448.905 -33.895 ;
        RECT -449.185 -34.775 -448.905 -34.495 ;
        RECT -431.265 -34.175 -430.985 -33.895 ;
        RECT -431.265 -34.775 -430.985 -34.495 ;
        RECT -413.345 -34.175 -413.065 -33.895 ;
        RECT -413.345 -34.775 -413.065 -34.495 ;
        RECT -395.425 -34.175 -395.145 -33.895 ;
        RECT -395.425 -34.775 -395.145 -34.495 ;
        RECT -377.505 -34.175 -377.225 -33.895 ;
        RECT -377.505 -34.775 -377.225 -34.495 ;
        RECT -359.585 -34.175 -359.305 -33.895 ;
        RECT -359.585 -34.775 -359.305 -34.495 ;
        RECT -341.665 -34.175 -341.385 -33.895 ;
        RECT -341.665 -34.775 -341.385 -34.495 ;
        RECT -323.745 -34.175 -323.465 -33.895 ;
        RECT -323.745 -34.775 -323.465 -34.495 ;
        RECT -305.825 -34.175 -305.545 -33.895 ;
        RECT -305.825 -34.775 -305.545 -34.495 ;
        RECT -287.905 -34.175 -287.625 -33.895 ;
        RECT -287.905 -34.775 -287.625 -34.495 ;
        RECT -269.985 -34.175 -269.705 -33.895 ;
        RECT -269.985 -34.775 -269.705 -34.495 ;
        RECT -252.065 -34.175 -251.785 -33.895 ;
        RECT -252.065 -34.775 -251.785 -34.495 ;
        RECT -234.145 -34.175 -233.865 -33.895 ;
        RECT -234.145 -34.775 -233.865 -34.495 ;
        RECT -216.225 -34.175 -215.945 -33.895 ;
        RECT -216.225 -34.775 -215.945 -34.495 ;
        RECT -198.305 -34.175 -198.025 -33.895 ;
        RECT -198.305 -34.775 -198.025 -34.495 ;
        RECT -179.265 -34.175 -178.985 -33.895 ;
        RECT -179.265 -34.775 -178.985 -34.495 ;
        RECT -161.345 -34.175 -161.065 -33.895 ;
        RECT -161.345 -34.775 -161.065 -34.495 ;
        RECT -143.425 -34.175 -143.145 -33.895 ;
        RECT -143.425 -34.775 -143.145 -34.495 ;
        RECT -125.505 -34.175 -125.225 -33.895 ;
        RECT -125.505 -34.775 -125.225 -34.495 ;
        RECT -107.585 -34.175 -107.305 -33.895 ;
        RECT -107.585 -34.775 -107.305 -34.495 ;
        RECT -89.665 -34.175 -89.385 -33.895 ;
        RECT -89.665 -34.775 -89.385 -34.495 ;
        RECT -71.745 -34.175 -71.465 -33.895 ;
        RECT -71.745 -34.775 -71.465 -34.495 ;
        RECT -53.825 -34.175 -53.545 -33.895 ;
        RECT -53.825 -34.775 -53.545 -34.495 ;
        RECT -35.905 -34.175 -35.625 -33.895 ;
        RECT -35.905 -34.775 -35.625 -34.495 ;
        RECT -17.985 -34.175 -17.705 -33.895 ;
        RECT -17.985 -34.775 -17.705 -34.495 ;
        RECT -0.065 -34.175 0.215 -33.895 ;
        RECT -0.065 -34.775 0.215 -34.495 ;
        RECT 17.855 -34.175 18.135 -33.895 ;
        RECT 17.855 -34.775 18.135 -34.495 ;
        RECT 35.775 -34.175 36.055 -33.895 ;
        RECT 35.775 -34.775 36.055 -34.495 ;
        RECT 53.695 -34.175 53.975 -33.895 ;
        RECT 53.695 -34.775 53.975 -34.495 ;
        RECT 71.615 -34.175 71.895 -33.895 ;
        RECT 71.615 -34.775 71.895 -34.495 ;
        RECT 89.535 -34.175 89.815 -33.895 ;
        RECT 89.535 -34.775 89.815 -34.495 ;
        RECT 106.715 -34.475 106.995 -34.195 ;
        RECT 107.315 -34.475 107.595 -34.195 ;
        RECT -471.585 -37.535 -471.305 -37.255 ;
        RECT -471.585 -38.135 -471.305 -37.855 ;
        RECT -462.625 -37.535 -462.345 -37.255 ;
        RECT -462.625 -38.135 -462.345 -37.855 ;
        RECT -453.665 -37.535 -453.385 -37.255 ;
        RECT -453.665 -38.135 -453.385 -37.855 ;
        RECT -444.705 -37.535 -444.425 -37.255 ;
        RECT -444.705 -38.135 -444.425 -37.855 ;
        RECT -435.745 -37.535 -435.465 -37.255 ;
        RECT -435.745 -38.135 -435.465 -37.855 ;
        RECT -426.785 -37.535 -426.505 -37.255 ;
        RECT -426.785 -38.135 -426.505 -37.855 ;
        RECT -417.825 -37.535 -417.545 -37.255 ;
        RECT -417.825 -38.135 -417.545 -37.855 ;
        RECT -408.865 -37.535 -408.585 -37.255 ;
        RECT -408.865 -38.135 -408.585 -37.855 ;
        RECT -399.905 -37.535 -399.625 -37.255 ;
        RECT -399.905 -38.135 -399.625 -37.855 ;
        RECT -390.945 -37.535 -390.665 -37.255 ;
        RECT -390.945 -38.135 -390.665 -37.855 ;
        RECT -381.985 -37.535 -381.705 -37.255 ;
        RECT -381.985 -38.135 -381.705 -37.855 ;
        RECT -373.025 -37.535 -372.745 -37.255 ;
        RECT -373.025 -38.135 -372.745 -37.855 ;
        RECT -364.065 -37.535 -363.785 -37.255 ;
        RECT -364.065 -38.135 -363.785 -37.855 ;
        RECT -355.105 -37.535 -354.825 -37.255 ;
        RECT -355.105 -38.135 -354.825 -37.855 ;
        RECT -346.145 -37.535 -345.865 -37.255 ;
        RECT -346.145 -38.135 -345.865 -37.855 ;
        RECT -337.185 -37.535 -336.905 -37.255 ;
        RECT -337.185 -38.135 -336.905 -37.855 ;
        RECT -328.225 -37.535 -327.945 -37.255 ;
        RECT -328.225 -38.135 -327.945 -37.855 ;
        RECT -319.265 -37.535 -318.985 -37.255 ;
        RECT -319.265 -38.135 -318.985 -37.855 ;
        RECT -310.305 -37.535 -310.025 -37.255 ;
        RECT -310.305 -38.135 -310.025 -37.855 ;
        RECT -301.345 -37.535 -301.065 -37.255 ;
        RECT -301.345 -38.135 -301.065 -37.855 ;
        RECT -292.385 -37.535 -292.105 -37.255 ;
        RECT -292.385 -38.135 -292.105 -37.855 ;
        RECT -283.425 -37.535 -283.145 -37.255 ;
        RECT -283.425 -38.135 -283.145 -37.855 ;
        RECT -274.465 -37.535 -274.185 -37.255 ;
        RECT -274.465 -38.135 -274.185 -37.855 ;
        RECT -265.505 -37.535 -265.225 -37.255 ;
        RECT -265.505 -38.135 -265.225 -37.855 ;
        RECT -256.545 -37.535 -256.265 -37.255 ;
        RECT -256.545 -38.135 -256.265 -37.855 ;
        RECT -247.585 -37.535 -247.305 -37.255 ;
        RECT -247.585 -38.135 -247.305 -37.855 ;
        RECT -238.625 -37.535 -238.345 -37.255 ;
        RECT -238.625 -38.135 -238.345 -37.855 ;
        RECT -229.665 -37.535 -229.385 -37.255 ;
        RECT -229.665 -38.135 -229.385 -37.855 ;
        RECT -220.705 -37.535 -220.425 -37.255 ;
        RECT -220.705 -38.135 -220.425 -37.855 ;
        RECT -211.745 -37.535 -211.465 -37.255 ;
        RECT -211.745 -38.135 -211.465 -37.855 ;
        RECT -202.785 -37.535 -202.505 -37.255 ;
        RECT -202.785 -38.135 -202.505 -37.855 ;
        RECT -193.825 -37.535 -193.545 -37.255 ;
        RECT -193.825 -38.135 -193.545 -37.855 ;
        RECT -183.745 -37.535 -183.465 -37.255 ;
        RECT -183.745 -38.135 -183.465 -37.855 ;
        RECT -174.785 -37.535 -174.505 -37.255 ;
        RECT -174.785 -38.135 -174.505 -37.855 ;
        RECT -165.825 -37.535 -165.545 -37.255 ;
        RECT -165.825 -38.135 -165.545 -37.855 ;
        RECT -156.865 -37.535 -156.585 -37.255 ;
        RECT -156.865 -38.135 -156.585 -37.855 ;
        RECT -147.905 -37.535 -147.625 -37.255 ;
        RECT -147.905 -38.135 -147.625 -37.855 ;
        RECT -138.945 -37.535 -138.665 -37.255 ;
        RECT -138.945 -38.135 -138.665 -37.855 ;
        RECT -129.985 -37.535 -129.705 -37.255 ;
        RECT -129.985 -38.135 -129.705 -37.855 ;
        RECT -121.025 -37.535 -120.745 -37.255 ;
        RECT -121.025 -38.135 -120.745 -37.855 ;
        RECT -112.065 -37.535 -111.785 -37.255 ;
        RECT -112.065 -38.135 -111.785 -37.855 ;
        RECT -103.105 -37.535 -102.825 -37.255 ;
        RECT -103.105 -38.135 -102.825 -37.855 ;
        RECT -94.145 -37.535 -93.865 -37.255 ;
        RECT -94.145 -38.135 -93.865 -37.855 ;
        RECT -85.185 -37.535 -84.905 -37.255 ;
        RECT -85.185 -38.135 -84.905 -37.855 ;
        RECT -76.225 -37.535 -75.945 -37.255 ;
        RECT -76.225 -38.135 -75.945 -37.855 ;
        RECT -67.265 -37.535 -66.985 -37.255 ;
        RECT -67.265 -38.135 -66.985 -37.855 ;
        RECT -58.305 -37.535 -58.025 -37.255 ;
        RECT -58.305 -38.135 -58.025 -37.855 ;
        RECT -49.345 -37.535 -49.065 -37.255 ;
        RECT -49.345 -38.135 -49.065 -37.855 ;
        RECT -40.385 -37.535 -40.105 -37.255 ;
        RECT -40.385 -38.135 -40.105 -37.855 ;
        RECT -31.425 -37.535 -31.145 -37.255 ;
        RECT -31.425 -38.135 -31.145 -37.855 ;
        RECT -22.465 -37.535 -22.185 -37.255 ;
        RECT -22.465 -38.135 -22.185 -37.855 ;
        RECT -13.505 -37.535 -13.225 -37.255 ;
        RECT -13.505 -38.135 -13.225 -37.855 ;
        RECT -4.545 -37.535 -4.265 -37.255 ;
        RECT -4.545 -38.135 -4.265 -37.855 ;
        RECT 4.415 -37.535 4.695 -37.255 ;
        RECT 4.415 -38.135 4.695 -37.855 ;
        RECT 13.375 -37.535 13.655 -37.255 ;
        RECT 13.375 -38.135 13.655 -37.855 ;
        RECT 22.335 -37.535 22.615 -37.255 ;
        RECT 22.335 -38.135 22.615 -37.855 ;
        RECT 31.295 -37.535 31.575 -37.255 ;
        RECT 31.295 -38.135 31.575 -37.855 ;
        RECT 40.255 -37.535 40.535 -37.255 ;
        RECT 40.255 -38.135 40.535 -37.855 ;
        RECT 49.215 -37.535 49.495 -37.255 ;
        RECT 49.215 -38.135 49.495 -37.855 ;
        RECT 58.175 -37.535 58.455 -37.255 ;
        RECT 58.175 -38.135 58.455 -37.855 ;
        RECT 67.135 -37.535 67.415 -37.255 ;
        RECT 67.135 -38.135 67.415 -37.855 ;
        RECT 76.095 -37.535 76.375 -37.255 ;
        RECT 76.095 -38.135 76.375 -37.855 ;
        RECT 85.055 -37.535 85.335 -37.255 ;
        RECT 85.055 -38.135 85.335 -37.855 ;
        RECT 94.015 -37.535 94.295 -37.255 ;
        RECT 94.015 -38.135 94.295 -37.855 ;
        RECT 104.915 -37.835 105.195 -37.555 ;
        RECT 105.515 -37.835 105.795 -37.555 ;
        RECT -473.825 -40.895 -473.545 -40.615 ;
        RECT -473.825 -41.495 -473.545 -41.215 ;
        RECT -469.345 -40.895 -469.065 -40.615 ;
        RECT -469.345 -41.495 -469.065 -41.215 ;
        RECT -464.865 -40.895 -464.585 -40.615 ;
        RECT -464.865 -41.495 -464.585 -41.215 ;
        RECT -460.385 -40.895 -460.105 -40.615 ;
        RECT -460.385 -41.495 -460.105 -41.215 ;
        RECT -455.905 -40.895 -455.625 -40.615 ;
        RECT -455.905 -41.495 -455.625 -41.215 ;
        RECT -451.425 -40.895 -451.145 -40.615 ;
        RECT -451.425 -41.495 -451.145 -41.215 ;
        RECT -446.945 -40.895 -446.665 -40.615 ;
        RECT -446.945 -41.495 -446.665 -41.215 ;
        RECT -442.465 -40.895 -442.185 -40.615 ;
        RECT -442.465 -41.495 -442.185 -41.215 ;
        RECT -437.985 -40.895 -437.705 -40.615 ;
        RECT -437.985 -41.495 -437.705 -41.215 ;
        RECT -433.505 -40.895 -433.225 -40.615 ;
        RECT -433.505 -41.495 -433.225 -41.215 ;
        RECT -429.025 -40.895 -428.745 -40.615 ;
        RECT -429.025 -41.495 -428.745 -41.215 ;
        RECT -424.545 -40.895 -424.265 -40.615 ;
        RECT -424.545 -41.495 -424.265 -41.215 ;
        RECT -420.065 -40.895 -419.785 -40.615 ;
        RECT -420.065 -41.495 -419.785 -41.215 ;
        RECT -415.585 -40.895 -415.305 -40.615 ;
        RECT -415.585 -41.495 -415.305 -41.215 ;
        RECT -411.105 -40.895 -410.825 -40.615 ;
        RECT -411.105 -41.495 -410.825 -41.215 ;
        RECT -406.625 -40.895 -406.345 -40.615 ;
        RECT -406.625 -41.495 -406.345 -41.215 ;
        RECT -402.145 -40.895 -401.865 -40.615 ;
        RECT -402.145 -41.495 -401.865 -41.215 ;
        RECT -397.665 -40.895 -397.385 -40.615 ;
        RECT -397.665 -41.495 -397.385 -41.215 ;
        RECT -393.185 -40.895 -392.905 -40.615 ;
        RECT -393.185 -41.495 -392.905 -41.215 ;
        RECT -388.705 -40.895 -388.425 -40.615 ;
        RECT -388.705 -41.495 -388.425 -41.215 ;
        RECT -384.225 -40.895 -383.945 -40.615 ;
        RECT -384.225 -41.495 -383.945 -41.215 ;
        RECT -379.745 -40.895 -379.465 -40.615 ;
        RECT -379.745 -41.495 -379.465 -41.215 ;
        RECT -375.265 -40.895 -374.985 -40.615 ;
        RECT -375.265 -41.495 -374.985 -41.215 ;
        RECT -370.785 -40.895 -370.505 -40.615 ;
        RECT -370.785 -41.495 -370.505 -41.215 ;
        RECT -366.305 -40.895 -366.025 -40.615 ;
        RECT -366.305 -41.495 -366.025 -41.215 ;
        RECT -361.825 -40.895 -361.545 -40.615 ;
        RECT -361.825 -41.495 -361.545 -41.215 ;
        RECT -357.345 -40.895 -357.065 -40.615 ;
        RECT -357.345 -41.495 -357.065 -41.215 ;
        RECT -352.865 -40.895 -352.585 -40.615 ;
        RECT -352.865 -41.495 -352.585 -41.215 ;
        RECT -348.385 -40.895 -348.105 -40.615 ;
        RECT -348.385 -41.495 -348.105 -41.215 ;
        RECT -343.905 -40.895 -343.625 -40.615 ;
        RECT -343.905 -41.495 -343.625 -41.215 ;
        RECT -339.425 -40.895 -339.145 -40.615 ;
        RECT -339.425 -41.495 -339.145 -41.215 ;
        RECT -334.945 -40.895 -334.665 -40.615 ;
        RECT -334.945 -41.495 -334.665 -41.215 ;
        RECT -330.465 -40.895 -330.185 -40.615 ;
        RECT -330.465 -41.495 -330.185 -41.215 ;
        RECT -325.985 -40.895 -325.705 -40.615 ;
        RECT -325.985 -41.495 -325.705 -41.215 ;
        RECT -321.505 -40.895 -321.225 -40.615 ;
        RECT -321.505 -41.495 -321.225 -41.215 ;
        RECT -317.025 -40.895 -316.745 -40.615 ;
        RECT -317.025 -41.495 -316.745 -41.215 ;
        RECT -312.545 -40.895 -312.265 -40.615 ;
        RECT -312.545 -41.495 -312.265 -41.215 ;
        RECT -308.065 -40.895 -307.785 -40.615 ;
        RECT -308.065 -41.495 -307.785 -41.215 ;
        RECT -303.585 -40.895 -303.305 -40.615 ;
        RECT -303.585 -41.495 -303.305 -41.215 ;
        RECT -299.105 -40.895 -298.825 -40.615 ;
        RECT -299.105 -41.495 -298.825 -41.215 ;
        RECT -294.625 -40.895 -294.345 -40.615 ;
        RECT -294.625 -41.495 -294.345 -41.215 ;
        RECT -290.145 -40.895 -289.865 -40.615 ;
        RECT -290.145 -41.495 -289.865 -41.215 ;
        RECT -285.665 -40.895 -285.385 -40.615 ;
        RECT -285.665 -41.495 -285.385 -41.215 ;
        RECT -281.185 -40.895 -280.905 -40.615 ;
        RECT -281.185 -41.495 -280.905 -41.215 ;
        RECT -276.705 -40.895 -276.425 -40.615 ;
        RECT -276.705 -41.495 -276.425 -41.215 ;
        RECT -272.225 -40.895 -271.945 -40.615 ;
        RECT -272.225 -41.495 -271.945 -41.215 ;
        RECT -267.745 -40.895 -267.465 -40.615 ;
        RECT -267.745 -41.495 -267.465 -41.215 ;
        RECT -263.265 -40.895 -262.985 -40.615 ;
        RECT -263.265 -41.495 -262.985 -41.215 ;
        RECT -258.785 -40.895 -258.505 -40.615 ;
        RECT -258.785 -41.495 -258.505 -41.215 ;
        RECT -254.305 -40.895 -254.025 -40.615 ;
        RECT -254.305 -41.495 -254.025 -41.215 ;
        RECT -249.825 -40.895 -249.545 -40.615 ;
        RECT -249.825 -41.495 -249.545 -41.215 ;
        RECT -245.345 -40.895 -245.065 -40.615 ;
        RECT -245.345 -41.495 -245.065 -41.215 ;
        RECT -240.865 -40.895 -240.585 -40.615 ;
        RECT -240.865 -41.495 -240.585 -41.215 ;
        RECT -236.385 -40.895 -236.105 -40.615 ;
        RECT -236.385 -41.495 -236.105 -41.215 ;
        RECT -231.905 -40.895 -231.625 -40.615 ;
        RECT -231.905 -41.495 -231.625 -41.215 ;
        RECT -227.425 -40.895 -227.145 -40.615 ;
        RECT -227.425 -41.495 -227.145 -41.215 ;
        RECT -222.945 -40.895 -222.665 -40.615 ;
        RECT -222.945 -41.495 -222.665 -41.215 ;
        RECT -218.465 -40.895 -218.185 -40.615 ;
        RECT -218.465 -41.495 -218.185 -41.215 ;
        RECT -213.985 -40.895 -213.705 -40.615 ;
        RECT -213.985 -41.495 -213.705 -41.215 ;
        RECT -209.505 -40.895 -209.225 -40.615 ;
        RECT -209.505 -41.495 -209.225 -41.215 ;
        RECT -205.025 -40.895 -204.745 -40.615 ;
        RECT -205.025 -41.495 -204.745 -41.215 ;
        RECT -200.545 -40.895 -200.265 -40.615 ;
        RECT -200.545 -41.495 -200.265 -41.215 ;
        RECT -196.065 -40.895 -195.785 -40.615 ;
        RECT -196.065 -41.495 -195.785 -41.215 ;
        RECT -191.585 -40.895 -191.305 -40.615 ;
        RECT -191.585 -41.495 -191.305 -41.215 ;
        RECT -185.985 -40.895 -185.705 -40.615 ;
        RECT -185.985 -41.495 -185.705 -41.215 ;
        RECT -181.505 -40.895 -181.225 -40.615 ;
        RECT -181.505 -41.495 -181.225 -41.215 ;
        RECT -177.025 -40.895 -176.745 -40.615 ;
        RECT -177.025 -41.495 -176.745 -41.215 ;
        RECT -172.545 -40.895 -172.265 -40.615 ;
        RECT -172.545 -41.495 -172.265 -41.215 ;
        RECT -168.065 -40.895 -167.785 -40.615 ;
        RECT -168.065 -41.495 -167.785 -41.215 ;
        RECT -163.585 -40.895 -163.305 -40.615 ;
        RECT -163.585 -41.495 -163.305 -41.215 ;
        RECT -159.105 -40.895 -158.825 -40.615 ;
        RECT -159.105 -41.495 -158.825 -41.215 ;
        RECT -154.625 -40.895 -154.345 -40.615 ;
        RECT -154.625 -41.495 -154.345 -41.215 ;
        RECT -150.145 -40.895 -149.865 -40.615 ;
        RECT -150.145 -41.495 -149.865 -41.215 ;
        RECT -145.665 -40.895 -145.385 -40.615 ;
        RECT -145.665 -41.495 -145.385 -41.215 ;
        RECT -141.185 -40.895 -140.905 -40.615 ;
        RECT -141.185 -41.495 -140.905 -41.215 ;
        RECT -136.705 -40.895 -136.425 -40.615 ;
        RECT -136.705 -41.495 -136.425 -41.215 ;
        RECT -132.225 -40.895 -131.945 -40.615 ;
        RECT -132.225 -41.495 -131.945 -41.215 ;
        RECT -127.745 -40.895 -127.465 -40.615 ;
        RECT -127.745 -41.495 -127.465 -41.215 ;
        RECT -123.265 -40.895 -122.985 -40.615 ;
        RECT -123.265 -41.495 -122.985 -41.215 ;
        RECT -118.785 -40.895 -118.505 -40.615 ;
        RECT -118.785 -41.495 -118.505 -41.215 ;
        RECT -114.305 -40.895 -114.025 -40.615 ;
        RECT -114.305 -41.495 -114.025 -41.215 ;
        RECT -109.825 -40.895 -109.545 -40.615 ;
        RECT -109.825 -41.495 -109.545 -41.215 ;
        RECT -105.345 -40.895 -105.065 -40.615 ;
        RECT -105.345 -41.495 -105.065 -41.215 ;
        RECT -100.865 -40.895 -100.585 -40.615 ;
        RECT -100.865 -41.495 -100.585 -41.215 ;
        RECT -96.385 -40.895 -96.105 -40.615 ;
        RECT -96.385 -41.495 -96.105 -41.215 ;
        RECT -91.905 -40.895 -91.625 -40.615 ;
        RECT -91.905 -41.495 -91.625 -41.215 ;
        RECT -87.425 -40.895 -87.145 -40.615 ;
        RECT -87.425 -41.495 -87.145 -41.215 ;
        RECT -82.945 -40.895 -82.665 -40.615 ;
        RECT -82.945 -41.495 -82.665 -41.215 ;
        RECT -78.465 -40.895 -78.185 -40.615 ;
        RECT -78.465 -41.495 -78.185 -41.215 ;
        RECT -73.985 -40.895 -73.705 -40.615 ;
        RECT -73.985 -41.495 -73.705 -41.215 ;
        RECT -69.505 -40.895 -69.225 -40.615 ;
        RECT -69.505 -41.495 -69.225 -41.215 ;
        RECT -65.025 -40.895 -64.745 -40.615 ;
        RECT -65.025 -41.495 -64.745 -41.215 ;
        RECT -60.545 -40.895 -60.265 -40.615 ;
        RECT -60.545 -41.495 -60.265 -41.215 ;
        RECT -56.065 -40.895 -55.785 -40.615 ;
        RECT -56.065 -41.495 -55.785 -41.215 ;
        RECT -51.585 -40.895 -51.305 -40.615 ;
        RECT -51.585 -41.495 -51.305 -41.215 ;
        RECT -47.105 -40.895 -46.825 -40.615 ;
        RECT -47.105 -41.495 -46.825 -41.215 ;
        RECT -42.625 -40.895 -42.345 -40.615 ;
        RECT -42.625 -41.495 -42.345 -41.215 ;
        RECT -38.145 -40.895 -37.865 -40.615 ;
        RECT -38.145 -41.495 -37.865 -41.215 ;
        RECT -33.665 -40.895 -33.385 -40.615 ;
        RECT -33.665 -41.495 -33.385 -41.215 ;
        RECT -29.185 -40.895 -28.905 -40.615 ;
        RECT -29.185 -41.495 -28.905 -41.215 ;
        RECT -24.705 -40.895 -24.425 -40.615 ;
        RECT -24.705 -41.495 -24.425 -41.215 ;
        RECT -20.225 -40.895 -19.945 -40.615 ;
        RECT -20.225 -41.495 -19.945 -41.215 ;
        RECT -15.745 -40.895 -15.465 -40.615 ;
        RECT -15.745 -41.495 -15.465 -41.215 ;
        RECT -11.265 -40.895 -10.985 -40.615 ;
        RECT -11.265 -41.495 -10.985 -41.215 ;
        RECT -6.785 -40.895 -6.505 -40.615 ;
        RECT -6.785 -41.495 -6.505 -41.215 ;
        RECT -2.305 -40.895 -2.025 -40.615 ;
        RECT -2.305 -41.495 -2.025 -41.215 ;
        RECT 2.175 -40.895 2.455 -40.615 ;
        RECT 2.175 -41.495 2.455 -41.215 ;
        RECT 6.655 -40.895 6.935 -40.615 ;
        RECT 6.655 -41.495 6.935 -41.215 ;
        RECT 11.135 -40.895 11.415 -40.615 ;
        RECT 11.135 -41.495 11.415 -41.215 ;
        RECT 15.615 -40.895 15.895 -40.615 ;
        RECT 15.615 -41.495 15.895 -41.215 ;
        RECT 20.095 -40.895 20.375 -40.615 ;
        RECT 20.095 -41.495 20.375 -41.215 ;
        RECT 24.575 -40.895 24.855 -40.615 ;
        RECT 24.575 -41.495 24.855 -41.215 ;
        RECT 29.055 -40.895 29.335 -40.615 ;
        RECT 29.055 -41.495 29.335 -41.215 ;
        RECT 33.535 -40.895 33.815 -40.615 ;
        RECT 33.535 -41.495 33.815 -41.215 ;
        RECT 38.015 -40.895 38.295 -40.615 ;
        RECT 38.015 -41.495 38.295 -41.215 ;
        RECT 42.495 -40.895 42.775 -40.615 ;
        RECT 42.495 -41.495 42.775 -41.215 ;
        RECT 46.975 -40.895 47.255 -40.615 ;
        RECT 46.975 -41.495 47.255 -41.215 ;
        RECT 51.455 -40.895 51.735 -40.615 ;
        RECT 51.455 -41.495 51.735 -41.215 ;
        RECT 55.935 -40.895 56.215 -40.615 ;
        RECT 55.935 -41.495 56.215 -41.215 ;
        RECT 60.415 -40.895 60.695 -40.615 ;
        RECT 60.415 -41.495 60.695 -41.215 ;
        RECT 64.895 -40.895 65.175 -40.615 ;
        RECT 64.895 -41.495 65.175 -41.215 ;
        RECT 69.375 -40.895 69.655 -40.615 ;
        RECT 69.375 -41.495 69.655 -41.215 ;
        RECT 73.855 -40.895 74.135 -40.615 ;
        RECT 73.855 -41.495 74.135 -41.215 ;
        RECT 78.335 -40.895 78.615 -40.615 ;
        RECT 78.335 -41.495 78.615 -41.215 ;
        RECT 82.815 -40.895 83.095 -40.615 ;
        RECT 82.815 -41.495 83.095 -41.215 ;
        RECT 87.295 -40.895 87.575 -40.615 ;
        RECT 87.295 -41.495 87.575 -41.215 ;
        RECT 91.775 -40.895 92.055 -40.615 ;
        RECT 91.775 -41.495 92.055 -41.215 ;
        RECT 96.255 -40.895 96.535 -40.615 ;
        RECT 96.255 -41.495 96.535 -41.215 ;
        RECT 103.115 -41.195 103.395 -40.915 ;
        RECT 103.715 -41.195 103.995 -40.915 ;
        RECT -474.945 -44.255 -474.665 -43.975 ;
        RECT -474.945 -44.855 -474.665 -44.575 ;
        RECT -472.705 -44.255 -472.425 -43.975 ;
        RECT -472.705 -44.855 -472.425 -44.575 ;
        RECT -470.465 -44.255 -470.185 -43.975 ;
        RECT -470.465 -44.855 -470.185 -44.575 ;
        RECT -468.225 -44.255 -467.945 -43.975 ;
        RECT -468.225 -44.855 -467.945 -44.575 ;
        RECT -465.985 -44.255 -465.705 -43.975 ;
        RECT -465.985 -44.855 -465.705 -44.575 ;
        RECT -463.745 -44.255 -463.465 -43.975 ;
        RECT -463.745 -44.855 -463.465 -44.575 ;
        RECT -461.505 -44.255 -461.225 -43.975 ;
        RECT -461.505 -44.855 -461.225 -44.575 ;
        RECT -459.265 -44.255 -458.985 -43.975 ;
        RECT -459.265 -44.855 -458.985 -44.575 ;
        RECT -457.025 -44.255 -456.745 -43.975 ;
        RECT -457.025 -44.855 -456.745 -44.575 ;
        RECT -454.785 -44.255 -454.505 -43.975 ;
        RECT -454.785 -44.855 -454.505 -44.575 ;
        RECT -452.545 -44.255 -452.265 -43.975 ;
        RECT -452.545 -44.855 -452.265 -44.575 ;
        RECT -450.305 -44.255 -450.025 -43.975 ;
        RECT -450.305 -44.855 -450.025 -44.575 ;
        RECT -448.065 -44.255 -447.785 -43.975 ;
        RECT -448.065 -44.855 -447.785 -44.575 ;
        RECT -445.825 -44.255 -445.545 -43.975 ;
        RECT -445.825 -44.855 -445.545 -44.575 ;
        RECT -443.585 -44.255 -443.305 -43.975 ;
        RECT -443.585 -44.855 -443.305 -44.575 ;
        RECT -441.345 -44.255 -441.065 -43.975 ;
        RECT -441.345 -44.855 -441.065 -44.575 ;
        RECT -439.105 -44.255 -438.825 -43.975 ;
        RECT -439.105 -44.855 -438.825 -44.575 ;
        RECT -436.865 -44.255 -436.585 -43.975 ;
        RECT -436.865 -44.855 -436.585 -44.575 ;
        RECT -434.625 -44.255 -434.345 -43.975 ;
        RECT -434.625 -44.855 -434.345 -44.575 ;
        RECT -432.385 -44.255 -432.105 -43.975 ;
        RECT -432.385 -44.855 -432.105 -44.575 ;
        RECT -430.145 -44.255 -429.865 -43.975 ;
        RECT -430.145 -44.855 -429.865 -44.575 ;
        RECT -427.905 -44.255 -427.625 -43.975 ;
        RECT -427.905 -44.855 -427.625 -44.575 ;
        RECT -425.665 -44.255 -425.385 -43.975 ;
        RECT -425.665 -44.855 -425.385 -44.575 ;
        RECT -423.425 -44.255 -423.145 -43.975 ;
        RECT -423.425 -44.855 -423.145 -44.575 ;
        RECT -421.185 -44.255 -420.905 -43.975 ;
        RECT -421.185 -44.855 -420.905 -44.575 ;
        RECT -418.945 -44.255 -418.665 -43.975 ;
        RECT -418.945 -44.855 -418.665 -44.575 ;
        RECT -416.705 -44.255 -416.425 -43.975 ;
        RECT -416.705 -44.855 -416.425 -44.575 ;
        RECT -414.465 -44.255 -414.185 -43.975 ;
        RECT -414.465 -44.855 -414.185 -44.575 ;
        RECT -412.225 -44.255 -411.945 -43.975 ;
        RECT -412.225 -44.855 -411.945 -44.575 ;
        RECT -409.985 -44.255 -409.705 -43.975 ;
        RECT -409.985 -44.855 -409.705 -44.575 ;
        RECT -407.745 -44.255 -407.465 -43.975 ;
        RECT -407.745 -44.855 -407.465 -44.575 ;
        RECT -405.505 -44.255 -405.225 -43.975 ;
        RECT -405.505 -44.855 -405.225 -44.575 ;
        RECT -403.265 -44.255 -402.985 -43.975 ;
        RECT -403.265 -44.855 -402.985 -44.575 ;
        RECT -401.025 -44.255 -400.745 -43.975 ;
        RECT -401.025 -44.855 -400.745 -44.575 ;
        RECT -398.785 -44.255 -398.505 -43.975 ;
        RECT -398.785 -44.855 -398.505 -44.575 ;
        RECT -396.545 -44.255 -396.265 -43.975 ;
        RECT -396.545 -44.855 -396.265 -44.575 ;
        RECT -394.305 -44.255 -394.025 -43.975 ;
        RECT -394.305 -44.855 -394.025 -44.575 ;
        RECT -392.065 -44.255 -391.785 -43.975 ;
        RECT -392.065 -44.855 -391.785 -44.575 ;
        RECT -389.825 -44.255 -389.545 -43.975 ;
        RECT -389.825 -44.855 -389.545 -44.575 ;
        RECT -387.585 -44.255 -387.305 -43.975 ;
        RECT -387.585 -44.855 -387.305 -44.575 ;
        RECT -385.345 -44.255 -385.065 -43.975 ;
        RECT -385.345 -44.855 -385.065 -44.575 ;
        RECT -383.105 -44.255 -382.825 -43.975 ;
        RECT -383.105 -44.855 -382.825 -44.575 ;
        RECT -380.865 -44.255 -380.585 -43.975 ;
        RECT -380.865 -44.855 -380.585 -44.575 ;
        RECT -378.625 -44.255 -378.345 -43.975 ;
        RECT -378.625 -44.855 -378.345 -44.575 ;
        RECT -376.385 -44.255 -376.105 -43.975 ;
        RECT -376.385 -44.855 -376.105 -44.575 ;
        RECT -374.145 -44.255 -373.865 -43.975 ;
        RECT -374.145 -44.855 -373.865 -44.575 ;
        RECT -371.905 -44.255 -371.625 -43.975 ;
        RECT -371.905 -44.855 -371.625 -44.575 ;
        RECT -369.665 -44.255 -369.385 -43.975 ;
        RECT -369.665 -44.855 -369.385 -44.575 ;
        RECT -367.425 -44.255 -367.145 -43.975 ;
        RECT -367.425 -44.855 -367.145 -44.575 ;
        RECT -365.185 -44.255 -364.905 -43.975 ;
        RECT -365.185 -44.855 -364.905 -44.575 ;
        RECT -362.945 -44.255 -362.665 -43.975 ;
        RECT -362.945 -44.855 -362.665 -44.575 ;
        RECT -360.705 -44.255 -360.425 -43.975 ;
        RECT -360.705 -44.855 -360.425 -44.575 ;
        RECT -358.465 -44.255 -358.185 -43.975 ;
        RECT -358.465 -44.855 -358.185 -44.575 ;
        RECT -356.225 -44.255 -355.945 -43.975 ;
        RECT -356.225 -44.855 -355.945 -44.575 ;
        RECT -353.985 -44.255 -353.705 -43.975 ;
        RECT -353.985 -44.855 -353.705 -44.575 ;
        RECT -351.745 -44.255 -351.465 -43.975 ;
        RECT -351.745 -44.855 -351.465 -44.575 ;
        RECT -349.505 -44.255 -349.225 -43.975 ;
        RECT -349.505 -44.855 -349.225 -44.575 ;
        RECT -347.265 -44.255 -346.985 -43.975 ;
        RECT -347.265 -44.855 -346.985 -44.575 ;
        RECT -345.025 -44.255 -344.745 -43.975 ;
        RECT -345.025 -44.855 -344.745 -44.575 ;
        RECT -342.785 -44.255 -342.505 -43.975 ;
        RECT -342.785 -44.855 -342.505 -44.575 ;
        RECT -340.545 -44.255 -340.265 -43.975 ;
        RECT -340.545 -44.855 -340.265 -44.575 ;
        RECT -338.305 -44.255 -338.025 -43.975 ;
        RECT -338.305 -44.855 -338.025 -44.575 ;
        RECT -336.065 -44.255 -335.785 -43.975 ;
        RECT -336.065 -44.855 -335.785 -44.575 ;
        RECT -333.825 -44.255 -333.545 -43.975 ;
        RECT -333.825 -44.855 -333.545 -44.575 ;
        RECT -331.585 -44.255 -331.305 -43.975 ;
        RECT -331.585 -44.855 -331.305 -44.575 ;
        RECT -329.345 -44.255 -329.065 -43.975 ;
        RECT -329.345 -44.855 -329.065 -44.575 ;
        RECT -327.105 -44.255 -326.825 -43.975 ;
        RECT -327.105 -44.855 -326.825 -44.575 ;
        RECT -324.865 -44.255 -324.585 -43.975 ;
        RECT -324.865 -44.855 -324.585 -44.575 ;
        RECT -322.625 -44.255 -322.345 -43.975 ;
        RECT -322.625 -44.855 -322.345 -44.575 ;
        RECT -320.385 -44.255 -320.105 -43.975 ;
        RECT -320.385 -44.855 -320.105 -44.575 ;
        RECT -318.145 -44.255 -317.865 -43.975 ;
        RECT -318.145 -44.855 -317.865 -44.575 ;
        RECT -315.905 -44.255 -315.625 -43.975 ;
        RECT -315.905 -44.855 -315.625 -44.575 ;
        RECT -313.665 -44.255 -313.385 -43.975 ;
        RECT -313.665 -44.855 -313.385 -44.575 ;
        RECT -311.425 -44.255 -311.145 -43.975 ;
        RECT -311.425 -44.855 -311.145 -44.575 ;
        RECT -309.185 -44.255 -308.905 -43.975 ;
        RECT -309.185 -44.855 -308.905 -44.575 ;
        RECT -306.945 -44.255 -306.665 -43.975 ;
        RECT -306.945 -44.855 -306.665 -44.575 ;
        RECT -304.705 -44.255 -304.425 -43.975 ;
        RECT -304.705 -44.855 -304.425 -44.575 ;
        RECT -302.465 -44.255 -302.185 -43.975 ;
        RECT -302.465 -44.855 -302.185 -44.575 ;
        RECT -300.225 -44.255 -299.945 -43.975 ;
        RECT -300.225 -44.855 -299.945 -44.575 ;
        RECT -297.985 -44.255 -297.705 -43.975 ;
        RECT -297.985 -44.855 -297.705 -44.575 ;
        RECT -295.745 -44.255 -295.465 -43.975 ;
        RECT -295.745 -44.855 -295.465 -44.575 ;
        RECT -293.505 -44.255 -293.225 -43.975 ;
        RECT -293.505 -44.855 -293.225 -44.575 ;
        RECT -291.265 -44.255 -290.985 -43.975 ;
        RECT -291.265 -44.855 -290.985 -44.575 ;
        RECT -289.025 -44.255 -288.745 -43.975 ;
        RECT -289.025 -44.855 -288.745 -44.575 ;
        RECT -286.785 -44.255 -286.505 -43.975 ;
        RECT -286.785 -44.855 -286.505 -44.575 ;
        RECT -284.545 -44.255 -284.265 -43.975 ;
        RECT -284.545 -44.855 -284.265 -44.575 ;
        RECT -282.305 -44.255 -282.025 -43.975 ;
        RECT -282.305 -44.855 -282.025 -44.575 ;
        RECT -280.065 -44.255 -279.785 -43.975 ;
        RECT -280.065 -44.855 -279.785 -44.575 ;
        RECT -277.825 -44.255 -277.545 -43.975 ;
        RECT -277.825 -44.855 -277.545 -44.575 ;
        RECT -275.585 -44.255 -275.305 -43.975 ;
        RECT -275.585 -44.855 -275.305 -44.575 ;
        RECT -273.345 -44.255 -273.065 -43.975 ;
        RECT -273.345 -44.855 -273.065 -44.575 ;
        RECT -271.105 -44.255 -270.825 -43.975 ;
        RECT -271.105 -44.855 -270.825 -44.575 ;
        RECT -268.865 -44.255 -268.585 -43.975 ;
        RECT -268.865 -44.855 -268.585 -44.575 ;
        RECT -266.625 -44.255 -266.345 -43.975 ;
        RECT -266.625 -44.855 -266.345 -44.575 ;
        RECT -264.385 -44.255 -264.105 -43.975 ;
        RECT -264.385 -44.855 -264.105 -44.575 ;
        RECT -262.145 -44.255 -261.865 -43.975 ;
        RECT -262.145 -44.855 -261.865 -44.575 ;
        RECT -259.905 -44.255 -259.625 -43.975 ;
        RECT -259.905 -44.855 -259.625 -44.575 ;
        RECT -257.665 -44.255 -257.385 -43.975 ;
        RECT -257.665 -44.855 -257.385 -44.575 ;
        RECT -255.425 -44.255 -255.145 -43.975 ;
        RECT -255.425 -44.855 -255.145 -44.575 ;
        RECT -253.185 -44.255 -252.905 -43.975 ;
        RECT -253.185 -44.855 -252.905 -44.575 ;
        RECT -250.945 -44.255 -250.665 -43.975 ;
        RECT -250.945 -44.855 -250.665 -44.575 ;
        RECT -248.705 -44.255 -248.425 -43.975 ;
        RECT -248.705 -44.855 -248.425 -44.575 ;
        RECT -246.465 -44.255 -246.185 -43.975 ;
        RECT -246.465 -44.855 -246.185 -44.575 ;
        RECT -244.225 -44.255 -243.945 -43.975 ;
        RECT -244.225 -44.855 -243.945 -44.575 ;
        RECT -241.985 -44.255 -241.705 -43.975 ;
        RECT -241.985 -44.855 -241.705 -44.575 ;
        RECT -239.745 -44.255 -239.465 -43.975 ;
        RECT -239.745 -44.855 -239.465 -44.575 ;
        RECT -237.505 -44.255 -237.225 -43.975 ;
        RECT -237.505 -44.855 -237.225 -44.575 ;
        RECT -235.265 -44.255 -234.985 -43.975 ;
        RECT -235.265 -44.855 -234.985 -44.575 ;
        RECT -233.025 -44.255 -232.745 -43.975 ;
        RECT -233.025 -44.855 -232.745 -44.575 ;
        RECT -230.785 -44.255 -230.505 -43.975 ;
        RECT -230.785 -44.855 -230.505 -44.575 ;
        RECT -228.545 -44.255 -228.265 -43.975 ;
        RECT -228.545 -44.855 -228.265 -44.575 ;
        RECT -226.305 -44.255 -226.025 -43.975 ;
        RECT -226.305 -44.855 -226.025 -44.575 ;
        RECT -224.065 -44.255 -223.785 -43.975 ;
        RECT -224.065 -44.855 -223.785 -44.575 ;
        RECT -221.825 -44.255 -221.545 -43.975 ;
        RECT -221.825 -44.855 -221.545 -44.575 ;
        RECT -219.585 -44.255 -219.305 -43.975 ;
        RECT -219.585 -44.855 -219.305 -44.575 ;
        RECT -217.345 -44.255 -217.065 -43.975 ;
        RECT -217.345 -44.855 -217.065 -44.575 ;
        RECT -215.105 -44.255 -214.825 -43.975 ;
        RECT -215.105 -44.855 -214.825 -44.575 ;
        RECT -212.865 -44.255 -212.585 -43.975 ;
        RECT -212.865 -44.855 -212.585 -44.575 ;
        RECT -210.625 -44.255 -210.345 -43.975 ;
        RECT -210.625 -44.855 -210.345 -44.575 ;
        RECT -208.385 -44.255 -208.105 -43.975 ;
        RECT -208.385 -44.855 -208.105 -44.575 ;
        RECT -206.145 -44.255 -205.865 -43.975 ;
        RECT -206.145 -44.855 -205.865 -44.575 ;
        RECT -203.905 -44.255 -203.625 -43.975 ;
        RECT -203.905 -44.855 -203.625 -44.575 ;
        RECT -201.665 -44.255 -201.385 -43.975 ;
        RECT -201.665 -44.855 -201.385 -44.575 ;
        RECT -199.425 -44.255 -199.145 -43.975 ;
        RECT -199.425 -44.855 -199.145 -44.575 ;
        RECT -197.185 -44.255 -196.905 -43.975 ;
        RECT -197.185 -44.855 -196.905 -44.575 ;
        RECT -194.945 -44.255 -194.665 -43.975 ;
        RECT -194.945 -44.855 -194.665 -44.575 ;
        RECT -192.705 -44.255 -192.425 -43.975 ;
        RECT -192.705 -44.855 -192.425 -44.575 ;
        RECT -190.465 -44.255 -190.185 -43.975 ;
        RECT -190.465 -44.855 -190.185 -44.575 ;
        RECT -187.105 -44.255 -186.825 -43.975 ;
        RECT -187.105 -44.855 -186.825 -44.575 ;
        RECT -184.865 -44.255 -184.585 -43.975 ;
        RECT -184.865 -44.855 -184.585 -44.575 ;
        RECT -182.625 -44.255 -182.345 -43.975 ;
        RECT -182.625 -44.855 -182.345 -44.575 ;
        RECT -180.385 -44.255 -180.105 -43.975 ;
        RECT -180.385 -44.855 -180.105 -44.575 ;
        RECT -178.145 -44.255 -177.865 -43.975 ;
        RECT -178.145 -44.855 -177.865 -44.575 ;
        RECT -175.905 -44.255 -175.625 -43.975 ;
        RECT -175.905 -44.855 -175.625 -44.575 ;
        RECT -173.665 -44.255 -173.385 -43.975 ;
        RECT -173.665 -44.855 -173.385 -44.575 ;
        RECT -171.425 -44.255 -171.145 -43.975 ;
        RECT -171.425 -44.855 -171.145 -44.575 ;
        RECT -169.185 -44.255 -168.905 -43.975 ;
        RECT -169.185 -44.855 -168.905 -44.575 ;
        RECT -166.945 -44.255 -166.665 -43.975 ;
        RECT -166.945 -44.855 -166.665 -44.575 ;
        RECT -164.705 -44.255 -164.425 -43.975 ;
        RECT -164.705 -44.855 -164.425 -44.575 ;
        RECT -162.465 -44.255 -162.185 -43.975 ;
        RECT -162.465 -44.855 -162.185 -44.575 ;
        RECT -160.225 -44.255 -159.945 -43.975 ;
        RECT -160.225 -44.855 -159.945 -44.575 ;
        RECT -157.985 -44.255 -157.705 -43.975 ;
        RECT -157.985 -44.855 -157.705 -44.575 ;
        RECT -155.745 -44.255 -155.465 -43.975 ;
        RECT -155.745 -44.855 -155.465 -44.575 ;
        RECT -153.505 -44.255 -153.225 -43.975 ;
        RECT -153.505 -44.855 -153.225 -44.575 ;
        RECT -151.265 -44.255 -150.985 -43.975 ;
        RECT -151.265 -44.855 -150.985 -44.575 ;
        RECT -149.025 -44.255 -148.745 -43.975 ;
        RECT -149.025 -44.855 -148.745 -44.575 ;
        RECT -146.785 -44.255 -146.505 -43.975 ;
        RECT -146.785 -44.855 -146.505 -44.575 ;
        RECT -144.545 -44.255 -144.265 -43.975 ;
        RECT -144.545 -44.855 -144.265 -44.575 ;
        RECT -142.305 -44.255 -142.025 -43.975 ;
        RECT -142.305 -44.855 -142.025 -44.575 ;
        RECT -140.065 -44.255 -139.785 -43.975 ;
        RECT -140.065 -44.855 -139.785 -44.575 ;
        RECT -137.825 -44.255 -137.545 -43.975 ;
        RECT -137.825 -44.855 -137.545 -44.575 ;
        RECT -135.585 -44.255 -135.305 -43.975 ;
        RECT -135.585 -44.855 -135.305 -44.575 ;
        RECT -133.345 -44.255 -133.065 -43.975 ;
        RECT -133.345 -44.855 -133.065 -44.575 ;
        RECT -131.105 -44.255 -130.825 -43.975 ;
        RECT -131.105 -44.855 -130.825 -44.575 ;
        RECT -128.865 -44.255 -128.585 -43.975 ;
        RECT -128.865 -44.855 -128.585 -44.575 ;
        RECT -126.625 -44.255 -126.345 -43.975 ;
        RECT -126.625 -44.855 -126.345 -44.575 ;
        RECT -124.385 -44.255 -124.105 -43.975 ;
        RECT -124.385 -44.855 -124.105 -44.575 ;
        RECT -122.145 -44.255 -121.865 -43.975 ;
        RECT -122.145 -44.855 -121.865 -44.575 ;
        RECT -119.905 -44.255 -119.625 -43.975 ;
        RECT -119.905 -44.855 -119.625 -44.575 ;
        RECT -117.665 -44.255 -117.385 -43.975 ;
        RECT -117.665 -44.855 -117.385 -44.575 ;
        RECT -115.425 -44.255 -115.145 -43.975 ;
        RECT -115.425 -44.855 -115.145 -44.575 ;
        RECT -113.185 -44.255 -112.905 -43.975 ;
        RECT -113.185 -44.855 -112.905 -44.575 ;
        RECT -110.945 -44.255 -110.665 -43.975 ;
        RECT -110.945 -44.855 -110.665 -44.575 ;
        RECT -108.705 -44.255 -108.425 -43.975 ;
        RECT -108.705 -44.855 -108.425 -44.575 ;
        RECT -106.465 -44.255 -106.185 -43.975 ;
        RECT -106.465 -44.855 -106.185 -44.575 ;
        RECT -104.225 -44.255 -103.945 -43.975 ;
        RECT -104.225 -44.855 -103.945 -44.575 ;
        RECT -101.985 -44.255 -101.705 -43.975 ;
        RECT -101.985 -44.855 -101.705 -44.575 ;
        RECT -99.745 -44.255 -99.465 -43.975 ;
        RECT -99.745 -44.855 -99.465 -44.575 ;
        RECT -97.505 -44.255 -97.225 -43.975 ;
        RECT -97.505 -44.855 -97.225 -44.575 ;
        RECT -95.265 -44.255 -94.985 -43.975 ;
        RECT -95.265 -44.855 -94.985 -44.575 ;
        RECT -93.025 -44.255 -92.745 -43.975 ;
        RECT -93.025 -44.855 -92.745 -44.575 ;
        RECT -90.785 -44.255 -90.505 -43.975 ;
        RECT -90.785 -44.855 -90.505 -44.575 ;
        RECT -88.545 -44.255 -88.265 -43.975 ;
        RECT -88.545 -44.855 -88.265 -44.575 ;
        RECT -86.305 -44.255 -86.025 -43.975 ;
        RECT -86.305 -44.855 -86.025 -44.575 ;
        RECT -84.065 -44.255 -83.785 -43.975 ;
        RECT -84.065 -44.855 -83.785 -44.575 ;
        RECT -81.825 -44.255 -81.545 -43.975 ;
        RECT -81.825 -44.855 -81.545 -44.575 ;
        RECT -79.585 -44.255 -79.305 -43.975 ;
        RECT -79.585 -44.855 -79.305 -44.575 ;
        RECT -77.345 -44.255 -77.065 -43.975 ;
        RECT -77.345 -44.855 -77.065 -44.575 ;
        RECT -75.105 -44.255 -74.825 -43.975 ;
        RECT -75.105 -44.855 -74.825 -44.575 ;
        RECT -72.865 -44.255 -72.585 -43.975 ;
        RECT -72.865 -44.855 -72.585 -44.575 ;
        RECT -70.625 -44.255 -70.345 -43.975 ;
        RECT -70.625 -44.855 -70.345 -44.575 ;
        RECT -68.385 -44.255 -68.105 -43.975 ;
        RECT -68.385 -44.855 -68.105 -44.575 ;
        RECT -66.145 -44.255 -65.865 -43.975 ;
        RECT -66.145 -44.855 -65.865 -44.575 ;
        RECT -63.905 -44.255 -63.625 -43.975 ;
        RECT -63.905 -44.855 -63.625 -44.575 ;
        RECT -61.665 -44.255 -61.385 -43.975 ;
        RECT -61.665 -44.855 -61.385 -44.575 ;
        RECT -59.425 -44.255 -59.145 -43.975 ;
        RECT -59.425 -44.855 -59.145 -44.575 ;
        RECT -57.185 -44.255 -56.905 -43.975 ;
        RECT -57.185 -44.855 -56.905 -44.575 ;
        RECT -54.945 -44.255 -54.665 -43.975 ;
        RECT -54.945 -44.855 -54.665 -44.575 ;
        RECT -52.705 -44.255 -52.425 -43.975 ;
        RECT -52.705 -44.855 -52.425 -44.575 ;
        RECT -50.465 -44.255 -50.185 -43.975 ;
        RECT -50.465 -44.855 -50.185 -44.575 ;
        RECT -48.225 -44.255 -47.945 -43.975 ;
        RECT -48.225 -44.855 -47.945 -44.575 ;
        RECT -45.985 -44.255 -45.705 -43.975 ;
        RECT -45.985 -44.855 -45.705 -44.575 ;
        RECT -43.745 -44.255 -43.465 -43.975 ;
        RECT -43.745 -44.855 -43.465 -44.575 ;
        RECT -41.505 -44.255 -41.225 -43.975 ;
        RECT -41.505 -44.855 -41.225 -44.575 ;
        RECT -39.265 -44.255 -38.985 -43.975 ;
        RECT -39.265 -44.855 -38.985 -44.575 ;
        RECT -37.025 -44.255 -36.745 -43.975 ;
        RECT -37.025 -44.855 -36.745 -44.575 ;
        RECT -34.785 -44.255 -34.505 -43.975 ;
        RECT -34.785 -44.855 -34.505 -44.575 ;
        RECT -32.545 -44.255 -32.265 -43.975 ;
        RECT -32.545 -44.855 -32.265 -44.575 ;
        RECT -30.305 -44.255 -30.025 -43.975 ;
        RECT -30.305 -44.855 -30.025 -44.575 ;
        RECT -28.065 -44.255 -27.785 -43.975 ;
        RECT -28.065 -44.855 -27.785 -44.575 ;
        RECT -25.825 -44.255 -25.545 -43.975 ;
        RECT -25.825 -44.855 -25.545 -44.575 ;
        RECT -23.585 -44.255 -23.305 -43.975 ;
        RECT -23.585 -44.855 -23.305 -44.575 ;
        RECT -21.345 -44.255 -21.065 -43.975 ;
        RECT -21.345 -44.855 -21.065 -44.575 ;
        RECT -19.105 -44.255 -18.825 -43.975 ;
        RECT -19.105 -44.855 -18.825 -44.575 ;
        RECT -16.865 -44.255 -16.585 -43.975 ;
        RECT -16.865 -44.855 -16.585 -44.575 ;
        RECT -14.625 -44.255 -14.345 -43.975 ;
        RECT -14.625 -44.855 -14.345 -44.575 ;
        RECT -12.385 -44.255 -12.105 -43.975 ;
        RECT -12.385 -44.855 -12.105 -44.575 ;
        RECT -10.145 -44.255 -9.865 -43.975 ;
        RECT -10.145 -44.855 -9.865 -44.575 ;
        RECT -7.905 -44.255 -7.625 -43.975 ;
        RECT -7.905 -44.855 -7.625 -44.575 ;
        RECT -5.665 -44.255 -5.385 -43.975 ;
        RECT -5.665 -44.855 -5.385 -44.575 ;
        RECT -3.425 -44.255 -3.145 -43.975 ;
        RECT -3.425 -44.855 -3.145 -44.575 ;
        RECT -1.185 -44.255 -0.905 -43.975 ;
        RECT -1.185 -44.855 -0.905 -44.575 ;
        RECT 1.055 -44.255 1.335 -43.975 ;
        RECT 1.055 -44.855 1.335 -44.575 ;
        RECT 3.295 -44.255 3.575 -43.975 ;
        RECT 3.295 -44.855 3.575 -44.575 ;
        RECT 5.535 -44.255 5.815 -43.975 ;
        RECT 5.535 -44.855 5.815 -44.575 ;
        RECT 7.775 -44.255 8.055 -43.975 ;
        RECT 7.775 -44.855 8.055 -44.575 ;
        RECT 10.015 -44.255 10.295 -43.975 ;
        RECT 10.015 -44.855 10.295 -44.575 ;
        RECT 12.255 -44.255 12.535 -43.975 ;
        RECT 12.255 -44.855 12.535 -44.575 ;
        RECT 14.495 -44.255 14.775 -43.975 ;
        RECT 14.495 -44.855 14.775 -44.575 ;
        RECT 16.735 -44.255 17.015 -43.975 ;
        RECT 16.735 -44.855 17.015 -44.575 ;
        RECT 18.975 -44.255 19.255 -43.975 ;
        RECT 18.975 -44.855 19.255 -44.575 ;
        RECT 21.215 -44.255 21.495 -43.975 ;
        RECT 21.215 -44.855 21.495 -44.575 ;
        RECT 23.455 -44.255 23.735 -43.975 ;
        RECT 23.455 -44.855 23.735 -44.575 ;
        RECT 25.695 -44.255 25.975 -43.975 ;
        RECT 25.695 -44.855 25.975 -44.575 ;
        RECT 27.935 -44.255 28.215 -43.975 ;
        RECT 27.935 -44.855 28.215 -44.575 ;
        RECT 30.175 -44.255 30.455 -43.975 ;
        RECT 30.175 -44.855 30.455 -44.575 ;
        RECT 32.415 -44.255 32.695 -43.975 ;
        RECT 32.415 -44.855 32.695 -44.575 ;
        RECT 34.655 -44.255 34.935 -43.975 ;
        RECT 34.655 -44.855 34.935 -44.575 ;
        RECT 36.895 -44.255 37.175 -43.975 ;
        RECT 36.895 -44.855 37.175 -44.575 ;
        RECT 39.135 -44.255 39.415 -43.975 ;
        RECT 39.135 -44.855 39.415 -44.575 ;
        RECT 41.375 -44.255 41.655 -43.975 ;
        RECT 41.375 -44.855 41.655 -44.575 ;
        RECT 43.615 -44.255 43.895 -43.975 ;
        RECT 43.615 -44.855 43.895 -44.575 ;
        RECT 45.855 -44.255 46.135 -43.975 ;
        RECT 45.855 -44.855 46.135 -44.575 ;
        RECT 48.095 -44.255 48.375 -43.975 ;
        RECT 48.095 -44.855 48.375 -44.575 ;
        RECT 50.335 -44.255 50.615 -43.975 ;
        RECT 50.335 -44.855 50.615 -44.575 ;
        RECT 52.575 -44.255 52.855 -43.975 ;
        RECT 52.575 -44.855 52.855 -44.575 ;
        RECT 54.815 -44.255 55.095 -43.975 ;
        RECT 54.815 -44.855 55.095 -44.575 ;
        RECT 57.055 -44.255 57.335 -43.975 ;
        RECT 57.055 -44.855 57.335 -44.575 ;
        RECT 59.295 -44.255 59.575 -43.975 ;
        RECT 59.295 -44.855 59.575 -44.575 ;
        RECT 61.535 -44.255 61.815 -43.975 ;
        RECT 61.535 -44.855 61.815 -44.575 ;
        RECT 63.775 -44.255 64.055 -43.975 ;
        RECT 63.775 -44.855 64.055 -44.575 ;
        RECT 66.015 -44.255 66.295 -43.975 ;
        RECT 66.015 -44.855 66.295 -44.575 ;
        RECT 68.255 -44.255 68.535 -43.975 ;
        RECT 68.255 -44.855 68.535 -44.575 ;
        RECT 70.495 -44.255 70.775 -43.975 ;
        RECT 70.495 -44.855 70.775 -44.575 ;
        RECT 72.735 -44.255 73.015 -43.975 ;
        RECT 72.735 -44.855 73.015 -44.575 ;
        RECT 74.975 -44.255 75.255 -43.975 ;
        RECT 74.975 -44.855 75.255 -44.575 ;
        RECT 77.215 -44.255 77.495 -43.975 ;
        RECT 77.215 -44.855 77.495 -44.575 ;
        RECT 79.455 -44.255 79.735 -43.975 ;
        RECT 79.455 -44.855 79.735 -44.575 ;
        RECT 81.695 -44.255 81.975 -43.975 ;
        RECT 81.695 -44.855 81.975 -44.575 ;
        RECT 83.935 -44.255 84.215 -43.975 ;
        RECT 83.935 -44.855 84.215 -44.575 ;
        RECT 86.175 -44.255 86.455 -43.975 ;
        RECT 86.175 -44.855 86.455 -44.575 ;
        RECT 88.415 -44.255 88.695 -43.975 ;
        RECT 88.415 -44.855 88.695 -44.575 ;
        RECT 90.655 -44.255 90.935 -43.975 ;
        RECT 90.655 -44.855 90.935 -44.575 ;
        RECT 92.895 -44.255 93.175 -43.975 ;
        RECT 92.895 -44.855 93.175 -44.575 ;
        RECT 95.135 -44.255 95.415 -43.975 ;
        RECT 95.135 -44.855 95.415 -44.575 ;
        RECT 97.375 -44.255 97.655 -43.975 ;
        RECT 97.375 -44.855 97.655 -44.575 ;
        RECT 101.315 -44.555 101.595 -44.275 ;
        RECT 101.915 -44.555 102.195 -44.275 ;
        RECT -474.945 -67.115 -474.665 -66.835 ;
        RECT -474.945 -67.715 -474.665 -67.435 ;
        RECT -472.705 -67.115 -472.425 -66.835 ;
        RECT -472.705 -67.715 -472.425 -67.435 ;
        RECT -470.465 -67.115 -470.185 -66.835 ;
        RECT -470.465 -67.715 -470.185 -67.435 ;
        RECT -468.225 -67.115 -467.945 -66.835 ;
        RECT -468.225 -67.715 -467.945 -67.435 ;
        RECT -465.985 -67.115 -465.705 -66.835 ;
        RECT -465.985 -67.715 -465.705 -67.435 ;
        RECT -463.745 -67.115 -463.465 -66.835 ;
        RECT -463.745 -67.715 -463.465 -67.435 ;
        RECT -461.505 -67.115 -461.225 -66.835 ;
        RECT -461.505 -67.715 -461.225 -67.435 ;
        RECT -459.265 -67.115 -458.985 -66.835 ;
        RECT -459.265 -67.715 -458.985 -67.435 ;
        RECT -457.025 -67.115 -456.745 -66.835 ;
        RECT -457.025 -67.715 -456.745 -67.435 ;
        RECT -454.785 -67.115 -454.505 -66.835 ;
        RECT -454.785 -67.715 -454.505 -67.435 ;
        RECT -452.545 -67.115 -452.265 -66.835 ;
        RECT -452.545 -67.715 -452.265 -67.435 ;
        RECT -450.305 -67.115 -450.025 -66.835 ;
        RECT -450.305 -67.715 -450.025 -67.435 ;
        RECT -448.065 -67.115 -447.785 -66.835 ;
        RECT -448.065 -67.715 -447.785 -67.435 ;
        RECT -445.825 -67.115 -445.545 -66.835 ;
        RECT -445.825 -67.715 -445.545 -67.435 ;
        RECT -443.585 -67.115 -443.305 -66.835 ;
        RECT -443.585 -67.715 -443.305 -67.435 ;
        RECT -441.345 -67.115 -441.065 -66.835 ;
        RECT -441.345 -67.715 -441.065 -67.435 ;
        RECT -439.105 -67.115 -438.825 -66.835 ;
        RECT -439.105 -67.715 -438.825 -67.435 ;
        RECT -436.865 -67.115 -436.585 -66.835 ;
        RECT -436.865 -67.715 -436.585 -67.435 ;
        RECT -434.625 -67.115 -434.345 -66.835 ;
        RECT -434.625 -67.715 -434.345 -67.435 ;
        RECT -432.385 -67.115 -432.105 -66.835 ;
        RECT -432.385 -67.715 -432.105 -67.435 ;
        RECT -430.145 -67.115 -429.865 -66.835 ;
        RECT -430.145 -67.715 -429.865 -67.435 ;
        RECT -427.905 -67.115 -427.625 -66.835 ;
        RECT -427.905 -67.715 -427.625 -67.435 ;
        RECT -425.665 -67.115 -425.385 -66.835 ;
        RECT -425.665 -67.715 -425.385 -67.435 ;
        RECT -423.425 -67.115 -423.145 -66.835 ;
        RECT -423.425 -67.715 -423.145 -67.435 ;
        RECT -421.185 -67.115 -420.905 -66.835 ;
        RECT -421.185 -67.715 -420.905 -67.435 ;
        RECT -418.945 -67.115 -418.665 -66.835 ;
        RECT -418.945 -67.715 -418.665 -67.435 ;
        RECT -416.705 -67.115 -416.425 -66.835 ;
        RECT -416.705 -67.715 -416.425 -67.435 ;
        RECT -414.465 -67.115 -414.185 -66.835 ;
        RECT -414.465 -67.715 -414.185 -67.435 ;
        RECT -412.225 -67.115 -411.945 -66.835 ;
        RECT -412.225 -67.715 -411.945 -67.435 ;
        RECT -409.985 -67.115 -409.705 -66.835 ;
        RECT -409.985 -67.715 -409.705 -67.435 ;
        RECT -407.745 -67.115 -407.465 -66.835 ;
        RECT -407.745 -67.715 -407.465 -67.435 ;
        RECT -405.505 -67.115 -405.225 -66.835 ;
        RECT -405.505 -67.715 -405.225 -67.435 ;
        RECT -403.265 -67.115 -402.985 -66.835 ;
        RECT -403.265 -67.715 -402.985 -67.435 ;
        RECT -401.025 -67.115 -400.745 -66.835 ;
        RECT -401.025 -67.715 -400.745 -67.435 ;
        RECT -398.785 -67.115 -398.505 -66.835 ;
        RECT -398.785 -67.715 -398.505 -67.435 ;
        RECT -396.545 -67.115 -396.265 -66.835 ;
        RECT -396.545 -67.715 -396.265 -67.435 ;
        RECT -394.305 -67.115 -394.025 -66.835 ;
        RECT -394.305 -67.715 -394.025 -67.435 ;
        RECT -392.065 -67.115 -391.785 -66.835 ;
        RECT -392.065 -67.715 -391.785 -67.435 ;
        RECT -389.825 -67.115 -389.545 -66.835 ;
        RECT -389.825 -67.715 -389.545 -67.435 ;
        RECT -387.585 -67.115 -387.305 -66.835 ;
        RECT -387.585 -67.715 -387.305 -67.435 ;
        RECT -385.345 -67.115 -385.065 -66.835 ;
        RECT -385.345 -67.715 -385.065 -67.435 ;
        RECT -383.105 -67.115 -382.825 -66.835 ;
        RECT -383.105 -67.715 -382.825 -67.435 ;
        RECT -380.865 -67.115 -380.585 -66.835 ;
        RECT -380.865 -67.715 -380.585 -67.435 ;
        RECT -378.625 -67.115 -378.345 -66.835 ;
        RECT -378.625 -67.715 -378.345 -67.435 ;
        RECT -376.385 -67.115 -376.105 -66.835 ;
        RECT -376.385 -67.715 -376.105 -67.435 ;
        RECT -374.145 -67.115 -373.865 -66.835 ;
        RECT -374.145 -67.715 -373.865 -67.435 ;
        RECT -371.905 -67.115 -371.625 -66.835 ;
        RECT -371.905 -67.715 -371.625 -67.435 ;
        RECT -369.665 -67.115 -369.385 -66.835 ;
        RECT -369.665 -67.715 -369.385 -67.435 ;
        RECT -367.425 -67.115 -367.145 -66.835 ;
        RECT -367.425 -67.715 -367.145 -67.435 ;
        RECT -365.185 -67.115 -364.905 -66.835 ;
        RECT -365.185 -67.715 -364.905 -67.435 ;
        RECT -362.945 -67.115 -362.665 -66.835 ;
        RECT -362.945 -67.715 -362.665 -67.435 ;
        RECT -360.705 -67.115 -360.425 -66.835 ;
        RECT -360.705 -67.715 -360.425 -67.435 ;
        RECT -358.465 -67.115 -358.185 -66.835 ;
        RECT -358.465 -67.715 -358.185 -67.435 ;
        RECT -356.225 -67.115 -355.945 -66.835 ;
        RECT -356.225 -67.715 -355.945 -67.435 ;
        RECT -353.985 -67.115 -353.705 -66.835 ;
        RECT -353.985 -67.715 -353.705 -67.435 ;
        RECT -351.745 -67.115 -351.465 -66.835 ;
        RECT -351.745 -67.715 -351.465 -67.435 ;
        RECT -349.505 -67.115 -349.225 -66.835 ;
        RECT -349.505 -67.715 -349.225 -67.435 ;
        RECT -347.265 -67.115 -346.985 -66.835 ;
        RECT -347.265 -67.715 -346.985 -67.435 ;
        RECT -345.025 -67.115 -344.745 -66.835 ;
        RECT -345.025 -67.715 -344.745 -67.435 ;
        RECT -342.785 -67.115 -342.505 -66.835 ;
        RECT -342.785 -67.715 -342.505 -67.435 ;
        RECT -340.545 -67.115 -340.265 -66.835 ;
        RECT -340.545 -67.715 -340.265 -67.435 ;
        RECT -338.305 -67.115 -338.025 -66.835 ;
        RECT -338.305 -67.715 -338.025 -67.435 ;
        RECT -336.065 -67.115 -335.785 -66.835 ;
        RECT -336.065 -67.715 -335.785 -67.435 ;
        RECT -333.825 -67.115 -333.545 -66.835 ;
        RECT -333.825 -67.715 -333.545 -67.435 ;
        RECT -331.585 -67.115 -331.305 -66.835 ;
        RECT -331.585 -67.715 -331.305 -67.435 ;
        RECT -329.345 -67.115 -329.065 -66.835 ;
        RECT -329.345 -67.715 -329.065 -67.435 ;
        RECT -327.105 -67.115 -326.825 -66.835 ;
        RECT -327.105 -67.715 -326.825 -67.435 ;
        RECT -324.865 -67.115 -324.585 -66.835 ;
        RECT -324.865 -67.715 -324.585 -67.435 ;
        RECT -322.625 -67.115 -322.345 -66.835 ;
        RECT -322.625 -67.715 -322.345 -67.435 ;
        RECT -320.385 -67.115 -320.105 -66.835 ;
        RECT -320.385 -67.715 -320.105 -67.435 ;
        RECT -318.145 -67.115 -317.865 -66.835 ;
        RECT -318.145 -67.715 -317.865 -67.435 ;
        RECT -315.905 -67.115 -315.625 -66.835 ;
        RECT -315.905 -67.715 -315.625 -67.435 ;
        RECT -313.665 -67.115 -313.385 -66.835 ;
        RECT -313.665 -67.715 -313.385 -67.435 ;
        RECT -311.425 -67.115 -311.145 -66.835 ;
        RECT -311.425 -67.715 -311.145 -67.435 ;
        RECT -309.185 -67.115 -308.905 -66.835 ;
        RECT -309.185 -67.715 -308.905 -67.435 ;
        RECT -306.945 -67.115 -306.665 -66.835 ;
        RECT -306.945 -67.715 -306.665 -67.435 ;
        RECT -304.705 -67.115 -304.425 -66.835 ;
        RECT -304.705 -67.715 -304.425 -67.435 ;
        RECT -302.465 -67.115 -302.185 -66.835 ;
        RECT -302.465 -67.715 -302.185 -67.435 ;
        RECT -300.225 -67.115 -299.945 -66.835 ;
        RECT -300.225 -67.715 -299.945 -67.435 ;
        RECT -297.985 -67.115 -297.705 -66.835 ;
        RECT -297.985 -67.715 -297.705 -67.435 ;
        RECT -295.745 -67.115 -295.465 -66.835 ;
        RECT -295.745 -67.715 -295.465 -67.435 ;
        RECT -293.505 -67.115 -293.225 -66.835 ;
        RECT -293.505 -67.715 -293.225 -67.435 ;
        RECT -291.265 -67.115 -290.985 -66.835 ;
        RECT -291.265 -67.715 -290.985 -67.435 ;
        RECT -289.025 -67.115 -288.745 -66.835 ;
        RECT -289.025 -67.715 -288.745 -67.435 ;
        RECT -286.785 -67.115 -286.505 -66.835 ;
        RECT -286.785 -67.715 -286.505 -67.435 ;
        RECT -284.545 -67.115 -284.265 -66.835 ;
        RECT -284.545 -67.715 -284.265 -67.435 ;
        RECT -282.305 -67.115 -282.025 -66.835 ;
        RECT -282.305 -67.715 -282.025 -67.435 ;
        RECT -280.065 -67.115 -279.785 -66.835 ;
        RECT -280.065 -67.715 -279.785 -67.435 ;
        RECT -277.825 -67.115 -277.545 -66.835 ;
        RECT -277.825 -67.715 -277.545 -67.435 ;
        RECT -275.585 -67.115 -275.305 -66.835 ;
        RECT -275.585 -67.715 -275.305 -67.435 ;
        RECT -273.345 -67.115 -273.065 -66.835 ;
        RECT -273.345 -67.715 -273.065 -67.435 ;
        RECT -271.105 -67.115 -270.825 -66.835 ;
        RECT -271.105 -67.715 -270.825 -67.435 ;
        RECT -268.865 -67.115 -268.585 -66.835 ;
        RECT -268.865 -67.715 -268.585 -67.435 ;
        RECT -266.625 -67.115 -266.345 -66.835 ;
        RECT -266.625 -67.715 -266.345 -67.435 ;
        RECT -264.385 -67.115 -264.105 -66.835 ;
        RECT -264.385 -67.715 -264.105 -67.435 ;
        RECT -262.145 -67.115 -261.865 -66.835 ;
        RECT -262.145 -67.715 -261.865 -67.435 ;
        RECT -259.905 -67.115 -259.625 -66.835 ;
        RECT -259.905 -67.715 -259.625 -67.435 ;
        RECT -257.665 -67.115 -257.385 -66.835 ;
        RECT -257.665 -67.715 -257.385 -67.435 ;
        RECT -255.425 -67.115 -255.145 -66.835 ;
        RECT -255.425 -67.715 -255.145 -67.435 ;
        RECT -253.185 -67.115 -252.905 -66.835 ;
        RECT -253.185 -67.715 -252.905 -67.435 ;
        RECT -250.945 -67.115 -250.665 -66.835 ;
        RECT -250.945 -67.715 -250.665 -67.435 ;
        RECT -248.705 -67.115 -248.425 -66.835 ;
        RECT -248.705 -67.715 -248.425 -67.435 ;
        RECT -246.465 -67.115 -246.185 -66.835 ;
        RECT -246.465 -67.715 -246.185 -67.435 ;
        RECT -244.225 -67.115 -243.945 -66.835 ;
        RECT -244.225 -67.715 -243.945 -67.435 ;
        RECT -241.985 -67.115 -241.705 -66.835 ;
        RECT -241.985 -67.715 -241.705 -67.435 ;
        RECT -239.745 -67.115 -239.465 -66.835 ;
        RECT -239.745 -67.715 -239.465 -67.435 ;
        RECT -237.505 -67.115 -237.225 -66.835 ;
        RECT -237.505 -67.715 -237.225 -67.435 ;
        RECT -235.265 -67.115 -234.985 -66.835 ;
        RECT -235.265 -67.715 -234.985 -67.435 ;
        RECT -233.025 -67.115 -232.745 -66.835 ;
        RECT -233.025 -67.715 -232.745 -67.435 ;
        RECT -230.785 -67.115 -230.505 -66.835 ;
        RECT -230.785 -67.715 -230.505 -67.435 ;
        RECT -228.545 -67.115 -228.265 -66.835 ;
        RECT -228.545 -67.715 -228.265 -67.435 ;
        RECT -226.305 -67.115 -226.025 -66.835 ;
        RECT -226.305 -67.715 -226.025 -67.435 ;
        RECT -224.065 -67.115 -223.785 -66.835 ;
        RECT -224.065 -67.715 -223.785 -67.435 ;
        RECT -221.825 -67.115 -221.545 -66.835 ;
        RECT -221.825 -67.715 -221.545 -67.435 ;
        RECT -219.585 -67.115 -219.305 -66.835 ;
        RECT -219.585 -67.715 -219.305 -67.435 ;
        RECT -217.345 -67.115 -217.065 -66.835 ;
        RECT -217.345 -67.715 -217.065 -67.435 ;
        RECT -215.105 -67.115 -214.825 -66.835 ;
        RECT -215.105 -67.715 -214.825 -67.435 ;
        RECT -212.865 -67.115 -212.585 -66.835 ;
        RECT -212.865 -67.715 -212.585 -67.435 ;
        RECT -210.625 -67.115 -210.345 -66.835 ;
        RECT -210.625 -67.715 -210.345 -67.435 ;
        RECT -208.385 -67.115 -208.105 -66.835 ;
        RECT -208.385 -67.715 -208.105 -67.435 ;
        RECT -206.145 -67.115 -205.865 -66.835 ;
        RECT -206.145 -67.715 -205.865 -67.435 ;
        RECT -203.905 -67.115 -203.625 -66.835 ;
        RECT -203.905 -67.715 -203.625 -67.435 ;
        RECT -201.665 -67.115 -201.385 -66.835 ;
        RECT -201.665 -67.715 -201.385 -67.435 ;
        RECT -199.425 -67.115 -199.145 -66.835 ;
        RECT -199.425 -67.715 -199.145 -67.435 ;
        RECT -197.185 -67.115 -196.905 -66.835 ;
        RECT -197.185 -67.715 -196.905 -67.435 ;
        RECT -194.945 -67.115 -194.665 -66.835 ;
        RECT -194.945 -67.715 -194.665 -67.435 ;
        RECT -192.705 -67.115 -192.425 -66.835 ;
        RECT -192.705 -67.715 -192.425 -67.435 ;
        RECT -190.465 -67.115 -190.185 -66.835 ;
        RECT -190.465 -67.715 -190.185 -67.435 ;
        RECT -187.105 -67.115 -186.825 -66.835 ;
        RECT -187.105 -67.715 -186.825 -67.435 ;
        RECT -184.865 -67.115 -184.585 -66.835 ;
        RECT -184.865 -67.715 -184.585 -67.435 ;
        RECT -182.625 -67.115 -182.345 -66.835 ;
        RECT -182.625 -67.715 -182.345 -67.435 ;
        RECT -180.385 -67.115 -180.105 -66.835 ;
        RECT -180.385 -67.715 -180.105 -67.435 ;
        RECT -178.145 -67.115 -177.865 -66.835 ;
        RECT -178.145 -67.715 -177.865 -67.435 ;
        RECT -175.905 -67.115 -175.625 -66.835 ;
        RECT -175.905 -67.715 -175.625 -67.435 ;
        RECT -173.665 -67.115 -173.385 -66.835 ;
        RECT -173.665 -67.715 -173.385 -67.435 ;
        RECT -171.425 -67.115 -171.145 -66.835 ;
        RECT -171.425 -67.715 -171.145 -67.435 ;
        RECT -169.185 -67.115 -168.905 -66.835 ;
        RECT -169.185 -67.715 -168.905 -67.435 ;
        RECT -166.945 -67.115 -166.665 -66.835 ;
        RECT -166.945 -67.715 -166.665 -67.435 ;
        RECT -164.705 -67.115 -164.425 -66.835 ;
        RECT -164.705 -67.715 -164.425 -67.435 ;
        RECT -162.465 -67.115 -162.185 -66.835 ;
        RECT -162.465 -67.715 -162.185 -67.435 ;
        RECT -160.225 -67.115 -159.945 -66.835 ;
        RECT -160.225 -67.715 -159.945 -67.435 ;
        RECT -157.985 -67.115 -157.705 -66.835 ;
        RECT -157.985 -67.715 -157.705 -67.435 ;
        RECT -155.745 -67.115 -155.465 -66.835 ;
        RECT -155.745 -67.715 -155.465 -67.435 ;
        RECT -153.505 -67.115 -153.225 -66.835 ;
        RECT -153.505 -67.715 -153.225 -67.435 ;
        RECT -151.265 -67.115 -150.985 -66.835 ;
        RECT -151.265 -67.715 -150.985 -67.435 ;
        RECT -149.025 -67.115 -148.745 -66.835 ;
        RECT -149.025 -67.715 -148.745 -67.435 ;
        RECT -146.785 -67.115 -146.505 -66.835 ;
        RECT -146.785 -67.715 -146.505 -67.435 ;
        RECT -144.545 -67.115 -144.265 -66.835 ;
        RECT -144.545 -67.715 -144.265 -67.435 ;
        RECT -142.305 -67.115 -142.025 -66.835 ;
        RECT -142.305 -67.715 -142.025 -67.435 ;
        RECT -140.065 -67.115 -139.785 -66.835 ;
        RECT -140.065 -67.715 -139.785 -67.435 ;
        RECT -137.825 -67.115 -137.545 -66.835 ;
        RECT -137.825 -67.715 -137.545 -67.435 ;
        RECT -135.585 -67.115 -135.305 -66.835 ;
        RECT -135.585 -67.715 -135.305 -67.435 ;
        RECT -133.345 -67.115 -133.065 -66.835 ;
        RECT -133.345 -67.715 -133.065 -67.435 ;
        RECT -131.105 -67.115 -130.825 -66.835 ;
        RECT -131.105 -67.715 -130.825 -67.435 ;
        RECT -128.865 -67.115 -128.585 -66.835 ;
        RECT -128.865 -67.715 -128.585 -67.435 ;
        RECT -126.625 -67.115 -126.345 -66.835 ;
        RECT -126.625 -67.715 -126.345 -67.435 ;
        RECT -124.385 -67.115 -124.105 -66.835 ;
        RECT -124.385 -67.715 -124.105 -67.435 ;
        RECT -122.145 -67.115 -121.865 -66.835 ;
        RECT -122.145 -67.715 -121.865 -67.435 ;
        RECT -119.905 -67.115 -119.625 -66.835 ;
        RECT -119.905 -67.715 -119.625 -67.435 ;
        RECT -117.665 -67.115 -117.385 -66.835 ;
        RECT -117.665 -67.715 -117.385 -67.435 ;
        RECT -115.425 -67.115 -115.145 -66.835 ;
        RECT -115.425 -67.715 -115.145 -67.435 ;
        RECT -113.185 -67.115 -112.905 -66.835 ;
        RECT -113.185 -67.715 -112.905 -67.435 ;
        RECT -110.945 -67.115 -110.665 -66.835 ;
        RECT -110.945 -67.715 -110.665 -67.435 ;
        RECT -108.705 -67.115 -108.425 -66.835 ;
        RECT -108.705 -67.715 -108.425 -67.435 ;
        RECT -106.465 -67.115 -106.185 -66.835 ;
        RECT -106.465 -67.715 -106.185 -67.435 ;
        RECT -104.225 -67.115 -103.945 -66.835 ;
        RECT -104.225 -67.715 -103.945 -67.435 ;
        RECT -101.985 -67.115 -101.705 -66.835 ;
        RECT -101.985 -67.715 -101.705 -67.435 ;
        RECT -99.745 -67.115 -99.465 -66.835 ;
        RECT -99.745 -67.715 -99.465 -67.435 ;
        RECT -97.505 -67.115 -97.225 -66.835 ;
        RECT -97.505 -67.715 -97.225 -67.435 ;
        RECT -95.265 -67.115 -94.985 -66.835 ;
        RECT -95.265 -67.715 -94.985 -67.435 ;
        RECT -93.025 -67.115 -92.745 -66.835 ;
        RECT -93.025 -67.715 -92.745 -67.435 ;
        RECT -90.785 -67.115 -90.505 -66.835 ;
        RECT -90.785 -67.715 -90.505 -67.435 ;
        RECT -88.545 -67.115 -88.265 -66.835 ;
        RECT -88.545 -67.715 -88.265 -67.435 ;
        RECT -86.305 -67.115 -86.025 -66.835 ;
        RECT -86.305 -67.715 -86.025 -67.435 ;
        RECT -84.065 -67.115 -83.785 -66.835 ;
        RECT -84.065 -67.715 -83.785 -67.435 ;
        RECT -81.825 -67.115 -81.545 -66.835 ;
        RECT -81.825 -67.715 -81.545 -67.435 ;
        RECT -79.585 -67.115 -79.305 -66.835 ;
        RECT -79.585 -67.715 -79.305 -67.435 ;
        RECT -77.345 -67.115 -77.065 -66.835 ;
        RECT -77.345 -67.715 -77.065 -67.435 ;
        RECT -75.105 -67.115 -74.825 -66.835 ;
        RECT -75.105 -67.715 -74.825 -67.435 ;
        RECT -72.865 -67.115 -72.585 -66.835 ;
        RECT -72.865 -67.715 -72.585 -67.435 ;
        RECT -70.625 -67.115 -70.345 -66.835 ;
        RECT -70.625 -67.715 -70.345 -67.435 ;
        RECT -68.385 -67.115 -68.105 -66.835 ;
        RECT -68.385 -67.715 -68.105 -67.435 ;
        RECT -66.145 -67.115 -65.865 -66.835 ;
        RECT -66.145 -67.715 -65.865 -67.435 ;
        RECT -63.905 -67.115 -63.625 -66.835 ;
        RECT -63.905 -67.715 -63.625 -67.435 ;
        RECT -61.665 -67.115 -61.385 -66.835 ;
        RECT -61.665 -67.715 -61.385 -67.435 ;
        RECT -59.425 -67.115 -59.145 -66.835 ;
        RECT -59.425 -67.715 -59.145 -67.435 ;
        RECT -57.185 -67.115 -56.905 -66.835 ;
        RECT -57.185 -67.715 -56.905 -67.435 ;
        RECT -54.945 -67.115 -54.665 -66.835 ;
        RECT -54.945 -67.715 -54.665 -67.435 ;
        RECT -52.705 -67.115 -52.425 -66.835 ;
        RECT -52.705 -67.715 -52.425 -67.435 ;
        RECT -50.465 -67.115 -50.185 -66.835 ;
        RECT -50.465 -67.715 -50.185 -67.435 ;
        RECT -48.225 -67.115 -47.945 -66.835 ;
        RECT -48.225 -67.715 -47.945 -67.435 ;
        RECT -45.985 -67.115 -45.705 -66.835 ;
        RECT -45.985 -67.715 -45.705 -67.435 ;
        RECT -43.745 -67.115 -43.465 -66.835 ;
        RECT -43.745 -67.715 -43.465 -67.435 ;
        RECT -41.505 -67.115 -41.225 -66.835 ;
        RECT -41.505 -67.715 -41.225 -67.435 ;
        RECT -39.265 -67.115 -38.985 -66.835 ;
        RECT -39.265 -67.715 -38.985 -67.435 ;
        RECT -37.025 -67.115 -36.745 -66.835 ;
        RECT -37.025 -67.715 -36.745 -67.435 ;
        RECT -34.785 -67.115 -34.505 -66.835 ;
        RECT -34.785 -67.715 -34.505 -67.435 ;
        RECT -32.545 -67.115 -32.265 -66.835 ;
        RECT -32.545 -67.715 -32.265 -67.435 ;
        RECT -30.305 -67.115 -30.025 -66.835 ;
        RECT -30.305 -67.715 -30.025 -67.435 ;
        RECT -28.065 -67.115 -27.785 -66.835 ;
        RECT -28.065 -67.715 -27.785 -67.435 ;
        RECT -25.825 -67.115 -25.545 -66.835 ;
        RECT -25.825 -67.715 -25.545 -67.435 ;
        RECT -23.585 -67.115 -23.305 -66.835 ;
        RECT -23.585 -67.715 -23.305 -67.435 ;
        RECT -21.345 -67.115 -21.065 -66.835 ;
        RECT -21.345 -67.715 -21.065 -67.435 ;
        RECT -19.105 -67.115 -18.825 -66.835 ;
        RECT -19.105 -67.715 -18.825 -67.435 ;
        RECT -16.865 -67.115 -16.585 -66.835 ;
        RECT -16.865 -67.715 -16.585 -67.435 ;
        RECT -14.625 -67.115 -14.345 -66.835 ;
        RECT -14.625 -67.715 -14.345 -67.435 ;
        RECT -12.385 -67.115 -12.105 -66.835 ;
        RECT -12.385 -67.715 -12.105 -67.435 ;
        RECT -10.145 -67.115 -9.865 -66.835 ;
        RECT -10.145 -67.715 -9.865 -67.435 ;
        RECT -7.905 -67.115 -7.625 -66.835 ;
        RECT -7.905 -67.715 -7.625 -67.435 ;
        RECT -5.665 -67.115 -5.385 -66.835 ;
        RECT -5.665 -67.715 -5.385 -67.435 ;
        RECT -3.425 -67.115 -3.145 -66.835 ;
        RECT -3.425 -67.715 -3.145 -67.435 ;
        RECT -1.185 -67.115 -0.905 -66.835 ;
        RECT -1.185 -67.715 -0.905 -67.435 ;
        RECT 1.055 -67.115 1.335 -66.835 ;
        RECT 1.055 -67.715 1.335 -67.435 ;
        RECT 3.295 -67.115 3.575 -66.835 ;
        RECT 3.295 -67.715 3.575 -67.435 ;
        RECT 5.535 -67.115 5.815 -66.835 ;
        RECT 5.535 -67.715 5.815 -67.435 ;
        RECT 7.775 -67.115 8.055 -66.835 ;
        RECT 7.775 -67.715 8.055 -67.435 ;
        RECT 10.015 -67.115 10.295 -66.835 ;
        RECT 10.015 -67.715 10.295 -67.435 ;
        RECT 12.255 -67.115 12.535 -66.835 ;
        RECT 12.255 -67.715 12.535 -67.435 ;
        RECT 14.495 -67.115 14.775 -66.835 ;
        RECT 14.495 -67.715 14.775 -67.435 ;
        RECT 16.735 -67.115 17.015 -66.835 ;
        RECT 16.735 -67.715 17.015 -67.435 ;
        RECT 18.975 -67.115 19.255 -66.835 ;
        RECT 18.975 -67.715 19.255 -67.435 ;
        RECT 21.215 -67.115 21.495 -66.835 ;
        RECT 21.215 -67.715 21.495 -67.435 ;
        RECT 23.455 -67.115 23.735 -66.835 ;
        RECT 23.455 -67.715 23.735 -67.435 ;
        RECT 25.695 -67.115 25.975 -66.835 ;
        RECT 25.695 -67.715 25.975 -67.435 ;
        RECT 27.935 -67.115 28.215 -66.835 ;
        RECT 27.935 -67.715 28.215 -67.435 ;
        RECT 30.175 -67.115 30.455 -66.835 ;
        RECT 30.175 -67.715 30.455 -67.435 ;
        RECT 32.415 -67.115 32.695 -66.835 ;
        RECT 32.415 -67.715 32.695 -67.435 ;
        RECT 34.655 -67.115 34.935 -66.835 ;
        RECT 34.655 -67.715 34.935 -67.435 ;
        RECT 36.895 -67.115 37.175 -66.835 ;
        RECT 36.895 -67.715 37.175 -67.435 ;
        RECT 39.135 -67.115 39.415 -66.835 ;
        RECT 39.135 -67.715 39.415 -67.435 ;
        RECT 41.375 -67.115 41.655 -66.835 ;
        RECT 41.375 -67.715 41.655 -67.435 ;
        RECT 43.615 -67.115 43.895 -66.835 ;
        RECT 43.615 -67.715 43.895 -67.435 ;
        RECT 45.855 -67.115 46.135 -66.835 ;
        RECT 45.855 -67.715 46.135 -67.435 ;
        RECT 48.095 -67.115 48.375 -66.835 ;
        RECT 48.095 -67.715 48.375 -67.435 ;
        RECT 50.335 -67.115 50.615 -66.835 ;
        RECT 50.335 -67.715 50.615 -67.435 ;
        RECT 52.575 -67.115 52.855 -66.835 ;
        RECT 52.575 -67.715 52.855 -67.435 ;
        RECT 54.815 -67.115 55.095 -66.835 ;
        RECT 54.815 -67.715 55.095 -67.435 ;
        RECT 57.055 -67.115 57.335 -66.835 ;
        RECT 57.055 -67.715 57.335 -67.435 ;
        RECT 59.295 -67.115 59.575 -66.835 ;
        RECT 59.295 -67.715 59.575 -67.435 ;
        RECT 61.535 -67.115 61.815 -66.835 ;
        RECT 61.535 -67.715 61.815 -67.435 ;
        RECT 63.775 -67.115 64.055 -66.835 ;
        RECT 63.775 -67.715 64.055 -67.435 ;
        RECT 66.015 -67.115 66.295 -66.835 ;
        RECT 66.015 -67.715 66.295 -67.435 ;
        RECT 68.255 -67.115 68.535 -66.835 ;
        RECT 68.255 -67.715 68.535 -67.435 ;
        RECT 70.495 -67.115 70.775 -66.835 ;
        RECT 70.495 -67.715 70.775 -67.435 ;
        RECT 72.735 -67.115 73.015 -66.835 ;
        RECT 72.735 -67.715 73.015 -67.435 ;
        RECT 74.975 -67.115 75.255 -66.835 ;
        RECT 74.975 -67.715 75.255 -67.435 ;
        RECT 77.215 -67.115 77.495 -66.835 ;
        RECT 77.215 -67.715 77.495 -67.435 ;
        RECT 79.455 -67.115 79.735 -66.835 ;
        RECT 79.455 -67.715 79.735 -67.435 ;
        RECT 81.695 -67.115 81.975 -66.835 ;
        RECT 81.695 -67.715 81.975 -67.435 ;
        RECT 83.935 -67.115 84.215 -66.835 ;
        RECT 83.935 -67.715 84.215 -67.435 ;
        RECT 86.175 -67.115 86.455 -66.835 ;
        RECT 86.175 -67.715 86.455 -67.435 ;
        RECT 88.415 -67.115 88.695 -66.835 ;
        RECT 88.415 -67.715 88.695 -67.435 ;
        RECT 90.655 -67.115 90.935 -66.835 ;
        RECT 90.655 -67.715 90.935 -67.435 ;
        RECT 92.895 -67.115 93.175 -66.835 ;
        RECT 92.895 -67.715 93.175 -67.435 ;
        RECT 95.135 -67.115 95.415 -66.835 ;
        RECT 95.135 -67.715 95.415 -67.435 ;
        RECT 97.375 -67.115 97.655 -66.835 ;
        RECT 97.375 -67.715 97.655 -67.435 ;
        RECT 101.315 -67.415 101.595 -67.135 ;
        RECT 101.915 -67.415 102.195 -67.135 ;
        RECT -473.825 -70.475 -473.545 -70.195 ;
        RECT -473.825 -71.075 -473.545 -70.795 ;
        RECT -469.345 -70.475 -469.065 -70.195 ;
        RECT -469.345 -71.075 -469.065 -70.795 ;
        RECT -464.865 -70.475 -464.585 -70.195 ;
        RECT -464.865 -71.075 -464.585 -70.795 ;
        RECT -460.385 -70.475 -460.105 -70.195 ;
        RECT -460.385 -71.075 -460.105 -70.795 ;
        RECT -455.905 -70.475 -455.625 -70.195 ;
        RECT -455.905 -71.075 -455.625 -70.795 ;
        RECT -451.425 -70.475 -451.145 -70.195 ;
        RECT -451.425 -71.075 -451.145 -70.795 ;
        RECT -446.945 -70.475 -446.665 -70.195 ;
        RECT -446.945 -71.075 -446.665 -70.795 ;
        RECT -442.465 -70.475 -442.185 -70.195 ;
        RECT -442.465 -71.075 -442.185 -70.795 ;
        RECT -437.985 -70.475 -437.705 -70.195 ;
        RECT -437.985 -71.075 -437.705 -70.795 ;
        RECT -433.505 -70.475 -433.225 -70.195 ;
        RECT -433.505 -71.075 -433.225 -70.795 ;
        RECT -429.025 -70.475 -428.745 -70.195 ;
        RECT -429.025 -71.075 -428.745 -70.795 ;
        RECT -424.545 -70.475 -424.265 -70.195 ;
        RECT -424.545 -71.075 -424.265 -70.795 ;
        RECT -420.065 -70.475 -419.785 -70.195 ;
        RECT -420.065 -71.075 -419.785 -70.795 ;
        RECT -415.585 -70.475 -415.305 -70.195 ;
        RECT -415.585 -71.075 -415.305 -70.795 ;
        RECT -411.105 -70.475 -410.825 -70.195 ;
        RECT -411.105 -71.075 -410.825 -70.795 ;
        RECT -406.625 -70.475 -406.345 -70.195 ;
        RECT -406.625 -71.075 -406.345 -70.795 ;
        RECT -402.145 -70.475 -401.865 -70.195 ;
        RECT -402.145 -71.075 -401.865 -70.795 ;
        RECT -397.665 -70.475 -397.385 -70.195 ;
        RECT -397.665 -71.075 -397.385 -70.795 ;
        RECT -393.185 -70.475 -392.905 -70.195 ;
        RECT -393.185 -71.075 -392.905 -70.795 ;
        RECT -388.705 -70.475 -388.425 -70.195 ;
        RECT -388.705 -71.075 -388.425 -70.795 ;
        RECT -384.225 -70.475 -383.945 -70.195 ;
        RECT -384.225 -71.075 -383.945 -70.795 ;
        RECT -379.745 -70.475 -379.465 -70.195 ;
        RECT -379.745 -71.075 -379.465 -70.795 ;
        RECT -375.265 -70.475 -374.985 -70.195 ;
        RECT -375.265 -71.075 -374.985 -70.795 ;
        RECT -370.785 -70.475 -370.505 -70.195 ;
        RECT -370.785 -71.075 -370.505 -70.795 ;
        RECT -366.305 -70.475 -366.025 -70.195 ;
        RECT -366.305 -71.075 -366.025 -70.795 ;
        RECT -361.825 -70.475 -361.545 -70.195 ;
        RECT -361.825 -71.075 -361.545 -70.795 ;
        RECT -357.345 -70.475 -357.065 -70.195 ;
        RECT -357.345 -71.075 -357.065 -70.795 ;
        RECT -352.865 -70.475 -352.585 -70.195 ;
        RECT -352.865 -71.075 -352.585 -70.795 ;
        RECT -348.385 -70.475 -348.105 -70.195 ;
        RECT -348.385 -71.075 -348.105 -70.795 ;
        RECT -343.905 -70.475 -343.625 -70.195 ;
        RECT -343.905 -71.075 -343.625 -70.795 ;
        RECT -339.425 -70.475 -339.145 -70.195 ;
        RECT -339.425 -71.075 -339.145 -70.795 ;
        RECT -334.945 -70.475 -334.665 -70.195 ;
        RECT -334.945 -71.075 -334.665 -70.795 ;
        RECT -330.465 -70.475 -330.185 -70.195 ;
        RECT -330.465 -71.075 -330.185 -70.795 ;
        RECT -325.985 -70.475 -325.705 -70.195 ;
        RECT -325.985 -71.075 -325.705 -70.795 ;
        RECT -321.505 -70.475 -321.225 -70.195 ;
        RECT -321.505 -71.075 -321.225 -70.795 ;
        RECT -317.025 -70.475 -316.745 -70.195 ;
        RECT -317.025 -71.075 -316.745 -70.795 ;
        RECT -312.545 -70.475 -312.265 -70.195 ;
        RECT -312.545 -71.075 -312.265 -70.795 ;
        RECT -308.065 -70.475 -307.785 -70.195 ;
        RECT -308.065 -71.075 -307.785 -70.795 ;
        RECT -303.585 -70.475 -303.305 -70.195 ;
        RECT -303.585 -71.075 -303.305 -70.795 ;
        RECT -299.105 -70.475 -298.825 -70.195 ;
        RECT -299.105 -71.075 -298.825 -70.795 ;
        RECT -294.625 -70.475 -294.345 -70.195 ;
        RECT -294.625 -71.075 -294.345 -70.795 ;
        RECT -290.145 -70.475 -289.865 -70.195 ;
        RECT -290.145 -71.075 -289.865 -70.795 ;
        RECT -285.665 -70.475 -285.385 -70.195 ;
        RECT -285.665 -71.075 -285.385 -70.795 ;
        RECT -281.185 -70.475 -280.905 -70.195 ;
        RECT -281.185 -71.075 -280.905 -70.795 ;
        RECT -276.705 -70.475 -276.425 -70.195 ;
        RECT -276.705 -71.075 -276.425 -70.795 ;
        RECT -272.225 -70.475 -271.945 -70.195 ;
        RECT -272.225 -71.075 -271.945 -70.795 ;
        RECT -267.745 -70.475 -267.465 -70.195 ;
        RECT -267.745 -71.075 -267.465 -70.795 ;
        RECT -263.265 -70.475 -262.985 -70.195 ;
        RECT -263.265 -71.075 -262.985 -70.795 ;
        RECT -258.785 -70.475 -258.505 -70.195 ;
        RECT -258.785 -71.075 -258.505 -70.795 ;
        RECT -254.305 -70.475 -254.025 -70.195 ;
        RECT -254.305 -71.075 -254.025 -70.795 ;
        RECT -249.825 -70.475 -249.545 -70.195 ;
        RECT -249.825 -71.075 -249.545 -70.795 ;
        RECT -245.345 -70.475 -245.065 -70.195 ;
        RECT -245.345 -71.075 -245.065 -70.795 ;
        RECT -240.865 -70.475 -240.585 -70.195 ;
        RECT -240.865 -71.075 -240.585 -70.795 ;
        RECT -236.385 -70.475 -236.105 -70.195 ;
        RECT -236.385 -71.075 -236.105 -70.795 ;
        RECT -231.905 -70.475 -231.625 -70.195 ;
        RECT -231.905 -71.075 -231.625 -70.795 ;
        RECT -227.425 -70.475 -227.145 -70.195 ;
        RECT -227.425 -71.075 -227.145 -70.795 ;
        RECT -222.945 -70.475 -222.665 -70.195 ;
        RECT -222.945 -71.075 -222.665 -70.795 ;
        RECT -218.465 -70.475 -218.185 -70.195 ;
        RECT -218.465 -71.075 -218.185 -70.795 ;
        RECT -213.985 -70.475 -213.705 -70.195 ;
        RECT -213.985 -71.075 -213.705 -70.795 ;
        RECT -209.505 -70.475 -209.225 -70.195 ;
        RECT -209.505 -71.075 -209.225 -70.795 ;
        RECT -205.025 -70.475 -204.745 -70.195 ;
        RECT -205.025 -71.075 -204.745 -70.795 ;
        RECT -200.545 -70.475 -200.265 -70.195 ;
        RECT -200.545 -71.075 -200.265 -70.795 ;
        RECT -196.065 -70.475 -195.785 -70.195 ;
        RECT -196.065 -71.075 -195.785 -70.795 ;
        RECT -191.585 -70.475 -191.305 -70.195 ;
        RECT -191.585 -71.075 -191.305 -70.795 ;
        RECT -185.985 -70.475 -185.705 -70.195 ;
        RECT -185.985 -71.075 -185.705 -70.795 ;
        RECT -181.505 -70.475 -181.225 -70.195 ;
        RECT -181.505 -71.075 -181.225 -70.795 ;
        RECT -177.025 -70.475 -176.745 -70.195 ;
        RECT -177.025 -71.075 -176.745 -70.795 ;
        RECT -172.545 -70.475 -172.265 -70.195 ;
        RECT -172.545 -71.075 -172.265 -70.795 ;
        RECT -168.065 -70.475 -167.785 -70.195 ;
        RECT -168.065 -71.075 -167.785 -70.795 ;
        RECT -163.585 -70.475 -163.305 -70.195 ;
        RECT -163.585 -71.075 -163.305 -70.795 ;
        RECT -159.105 -70.475 -158.825 -70.195 ;
        RECT -159.105 -71.075 -158.825 -70.795 ;
        RECT -154.625 -70.475 -154.345 -70.195 ;
        RECT -154.625 -71.075 -154.345 -70.795 ;
        RECT -150.145 -70.475 -149.865 -70.195 ;
        RECT -150.145 -71.075 -149.865 -70.795 ;
        RECT -145.665 -70.475 -145.385 -70.195 ;
        RECT -145.665 -71.075 -145.385 -70.795 ;
        RECT -141.185 -70.475 -140.905 -70.195 ;
        RECT -141.185 -71.075 -140.905 -70.795 ;
        RECT -136.705 -70.475 -136.425 -70.195 ;
        RECT -136.705 -71.075 -136.425 -70.795 ;
        RECT -132.225 -70.475 -131.945 -70.195 ;
        RECT -132.225 -71.075 -131.945 -70.795 ;
        RECT -127.745 -70.475 -127.465 -70.195 ;
        RECT -127.745 -71.075 -127.465 -70.795 ;
        RECT -123.265 -70.475 -122.985 -70.195 ;
        RECT -123.265 -71.075 -122.985 -70.795 ;
        RECT -118.785 -70.475 -118.505 -70.195 ;
        RECT -118.785 -71.075 -118.505 -70.795 ;
        RECT -114.305 -70.475 -114.025 -70.195 ;
        RECT -114.305 -71.075 -114.025 -70.795 ;
        RECT -109.825 -70.475 -109.545 -70.195 ;
        RECT -109.825 -71.075 -109.545 -70.795 ;
        RECT -105.345 -70.475 -105.065 -70.195 ;
        RECT -105.345 -71.075 -105.065 -70.795 ;
        RECT -100.865 -70.475 -100.585 -70.195 ;
        RECT -100.865 -71.075 -100.585 -70.795 ;
        RECT -96.385 -70.475 -96.105 -70.195 ;
        RECT -96.385 -71.075 -96.105 -70.795 ;
        RECT -91.905 -70.475 -91.625 -70.195 ;
        RECT -91.905 -71.075 -91.625 -70.795 ;
        RECT -87.425 -70.475 -87.145 -70.195 ;
        RECT -87.425 -71.075 -87.145 -70.795 ;
        RECT -82.945 -70.475 -82.665 -70.195 ;
        RECT -82.945 -71.075 -82.665 -70.795 ;
        RECT -78.465 -70.475 -78.185 -70.195 ;
        RECT -78.465 -71.075 -78.185 -70.795 ;
        RECT -73.985 -70.475 -73.705 -70.195 ;
        RECT -73.985 -71.075 -73.705 -70.795 ;
        RECT -69.505 -70.475 -69.225 -70.195 ;
        RECT -69.505 -71.075 -69.225 -70.795 ;
        RECT -65.025 -70.475 -64.745 -70.195 ;
        RECT -65.025 -71.075 -64.745 -70.795 ;
        RECT -60.545 -70.475 -60.265 -70.195 ;
        RECT -60.545 -71.075 -60.265 -70.795 ;
        RECT -56.065 -70.475 -55.785 -70.195 ;
        RECT -56.065 -71.075 -55.785 -70.795 ;
        RECT -51.585 -70.475 -51.305 -70.195 ;
        RECT -51.585 -71.075 -51.305 -70.795 ;
        RECT -47.105 -70.475 -46.825 -70.195 ;
        RECT -47.105 -71.075 -46.825 -70.795 ;
        RECT -42.625 -70.475 -42.345 -70.195 ;
        RECT -42.625 -71.075 -42.345 -70.795 ;
        RECT -38.145 -70.475 -37.865 -70.195 ;
        RECT -38.145 -71.075 -37.865 -70.795 ;
        RECT -33.665 -70.475 -33.385 -70.195 ;
        RECT -33.665 -71.075 -33.385 -70.795 ;
        RECT -29.185 -70.475 -28.905 -70.195 ;
        RECT -29.185 -71.075 -28.905 -70.795 ;
        RECT -24.705 -70.475 -24.425 -70.195 ;
        RECT -24.705 -71.075 -24.425 -70.795 ;
        RECT -20.225 -70.475 -19.945 -70.195 ;
        RECT -20.225 -71.075 -19.945 -70.795 ;
        RECT -15.745 -70.475 -15.465 -70.195 ;
        RECT -15.745 -71.075 -15.465 -70.795 ;
        RECT -11.265 -70.475 -10.985 -70.195 ;
        RECT -11.265 -71.075 -10.985 -70.795 ;
        RECT -6.785 -70.475 -6.505 -70.195 ;
        RECT -6.785 -71.075 -6.505 -70.795 ;
        RECT -2.305 -70.475 -2.025 -70.195 ;
        RECT -2.305 -71.075 -2.025 -70.795 ;
        RECT 2.175 -70.475 2.455 -70.195 ;
        RECT 2.175 -71.075 2.455 -70.795 ;
        RECT 6.655 -70.475 6.935 -70.195 ;
        RECT 6.655 -71.075 6.935 -70.795 ;
        RECT 11.135 -70.475 11.415 -70.195 ;
        RECT 11.135 -71.075 11.415 -70.795 ;
        RECT 15.615 -70.475 15.895 -70.195 ;
        RECT 15.615 -71.075 15.895 -70.795 ;
        RECT 20.095 -70.475 20.375 -70.195 ;
        RECT 20.095 -71.075 20.375 -70.795 ;
        RECT 24.575 -70.475 24.855 -70.195 ;
        RECT 24.575 -71.075 24.855 -70.795 ;
        RECT 29.055 -70.475 29.335 -70.195 ;
        RECT 29.055 -71.075 29.335 -70.795 ;
        RECT 33.535 -70.475 33.815 -70.195 ;
        RECT 33.535 -71.075 33.815 -70.795 ;
        RECT 38.015 -70.475 38.295 -70.195 ;
        RECT 38.015 -71.075 38.295 -70.795 ;
        RECT 42.495 -70.475 42.775 -70.195 ;
        RECT 42.495 -71.075 42.775 -70.795 ;
        RECT 46.975 -70.475 47.255 -70.195 ;
        RECT 46.975 -71.075 47.255 -70.795 ;
        RECT 51.455 -70.475 51.735 -70.195 ;
        RECT 51.455 -71.075 51.735 -70.795 ;
        RECT 55.935 -70.475 56.215 -70.195 ;
        RECT 55.935 -71.075 56.215 -70.795 ;
        RECT 60.415 -70.475 60.695 -70.195 ;
        RECT 60.415 -71.075 60.695 -70.795 ;
        RECT 64.895 -70.475 65.175 -70.195 ;
        RECT 64.895 -71.075 65.175 -70.795 ;
        RECT 69.375 -70.475 69.655 -70.195 ;
        RECT 69.375 -71.075 69.655 -70.795 ;
        RECT 73.855 -70.475 74.135 -70.195 ;
        RECT 73.855 -71.075 74.135 -70.795 ;
        RECT 78.335 -70.475 78.615 -70.195 ;
        RECT 78.335 -71.075 78.615 -70.795 ;
        RECT 82.815 -70.475 83.095 -70.195 ;
        RECT 82.815 -71.075 83.095 -70.795 ;
        RECT 87.295 -70.475 87.575 -70.195 ;
        RECT 87.295 -71.075 87.575 -70.795 ;
        RECT 91.775 -70.475 92.055 -70.195 ;
        RECT 91.775 -71.075 92.055 -70.795 ;
        RECT 96.255 -70.475 96.535 -70.195 ;
        RECT 96.255 -71.075 96.535 -70.795 ;
        RECT 103.115 -70.775 103.395 -70.495 ;
        RECT 103.715 -70.775 103.995 -70.495 ;
        RECT -471.585 -73.835 -471.305 -73.555 ;
        RECT -471.585 -74.435 -471.305 -74.155 ;
        RECT -462.625 -73.835 -462.345 -73.555 ;
        RECT -462.625 -74.435 -462.345 -74.155 ;
        RECT -453.665 -73.835 -453.385 -73.555 ;
        RECT -453.665 -74.435 -453.385 -74.155 ;
        RECT -444.705 -73.835 -444.425 -73.555 ;
        RECT -444.705 -74.435 -444.425 -74.155 ;
        RECT -435.745 -73.835 -435.465 -73.555 ;
        RECT -435.745 -74.435 -435.465 -74.155 ;
        RECT -426.785 -73.835 -426.505 -73.555 ;
        RECT -426.785 -74.435 -426.505 -74.155 ;
        RECT -417.825 -73.835 -417.545 -73.555 ;
        RECT -417.825 -74.435 -417.545 -74.155 ;
        RECT -408.865 -73.835 -408.585 -73.555 ;
        RECT -408.865 -74.435 -408.585 -74.155 ;
        RECT -399.905 -73.835 -399.625 -73.555 ;
        RECT -399.905 -74.435 -399.625 -74.155 ;
        RECT -390.945 -73.835 -390.665 -73.555 ;
        RECT -390.945 -74.435 -390.665 -74.155 ;
        RECT -381.985 -73.835 -381.705 -73.555 ;
        RECT -381.985 -74.435 -381.705 -74.155 ;
        RECT -373.025 -73.835 -372.745 -73.555 ;
        RECT -373.025 -74.435 -372.745 -74.155 ;
        RECT -364.065 -73.835 -363.785 -73.555 ;
        RECT -364.065 -74.435 -363.785 -74.155 ;
        RECT -355.105 -73.835 -354.825 -73.555 ;
        RECT -355.105 -74.435 -354.825 -74.155 ;
        RECT -346.145 -73.835 -345.865 -73.555 ;
        RECT -346.145 -74.435 -345.865 -74.155 ;
        RECT -337.185 -73.835 -336.905 -73.555 ;
        RECT -337.185 -74.435 -336.905 -74.155 ;
        RECT -328.225 -73.835 -327.945 -73.555 ;
        RECT -328.225 -74.435 -327.945 -74.155 ;
        RECT -319.265 -73.835 -318.985 -73.555 ;
        RECT -319.265 -74.435 -318.985 -74.155 ;
        RECT -310.305 -73.835 -310.025 -73.555 ;
        RECT -310.305 -74.435 -310.025 -74.155 ;
        RECT -301.345 -73.835 -301.065 -73.555 ;
        RECT -301.345 -74.435 -301.065 -74.155 ;
        RECT -292.385 -73.835 -292.105 -73.555 ;
        RECT -292.385 -74.435 -292.105 -74.155 ;
        RECT -283.425 -73.835 -283.145 -73.555 ;
        RECT -283.425 -74.435 -283.145 -74.155 ;
        RECT -274.465 -73.835 -274.185 -73.555 ;
        RECT -274.465 -74.435 -274.185 -74.155 ;
        RECT -265.505 -73.835 -265.225 -73.555 ;
        RECT -265.505 -74.435 -265.225 -74.155 ;
        RECT -256.545 -73.835 -256.265 -73.555 ;
        RECT -256.545 -74.435 -256.265 -74.155 ;
        RECT -247.585 -73.835 -247.305 -73.555 ;
        RECT -247.585 -74.435 -247.305 -74.155 ;
        RECT -238.625 -73.835 -238.345 -73.555 ;
        RECT -238.625 -74.435 -238.345 -74.155 ;
        RECT -229.665 -73.835 -229.385 -73.555 ;
        RECT -229.665 -74.435 -229.385 -74.155 ;
        RECT -220.705 -73.835 -220.425 -73.555 ;
        RECT -220.705 -74.435 -220.425 -74.155 ;
        RECT -211.745 -73.835 -211.465 -73.555 ;
        RECT -211.745 -74.435 -211.465 -74.155 ;
        RECT -202.785 -73.835 -202.505 -73.555 ;
        RECT -202.785 -74.435 -202.505 -74.155 ;
        RECT -193.825 -73.835 -193.545 -73.555 ;
        RECT -193.825 -74.435 -193.545 -74.155 ;
        RECT -183.745 -73.835 -183.465 -73.555 ;
        RECT -183.745 -74.435 -183.465 -74.155 ;
        RECT -174.785 -73.835 -174.505 -73.555 ;
        RECT -174.785 -74.435 -174.505 -74.155 ;
        RECT -165.825 -73.835 -165.545 -73.555 ;
        RECT -165.825 -74.435 -165.545 -74.155 ;
        RECT -156.865 -73.835 -156.585 -73.555 ;
        RECT -156.865 -74.435 -156.585 -74.155 ;
        RECT -147.905 -73.835 -147.625 -73.555 ;
        RECT -147.905 -74.435 -147.625 -74.155 ;
        RECT -138.945 -73.835 -138.665 -73.555 ;
        RECT -138.945 -74.435 -138.665 -74.155 ;
        RECT -129.985 -73.835 -129.705 -73.555 ;
        RECT -129.985 -74.435 -129.705 -74.155 ;
        RECT -121.025 -73.835 -120.745 -73.555 ;
        RECT -121.025 -74.435 -120.745 -74.155 ;
        RECT -112.065 -73.835 -111.785 -73.555 ;
        RECT -112.065 -74.435 -111.785 -74.155 ;
        RECT -103.105 -73.835 -102.825 -73.555 ;
        RECT -103.105 -74.435 -102.825 -74.155 ;
        RECT -94.145 -73.835 -93.865 -73.555 ;
        RECT -94.145 -74.435 -93.865 -74.155 ;
        RECT -85.185 -73.835 -84.905 -73.555 ;
        RECT -85.185 -74.435 -84.905 -74.155 ;
        RECT -76.225 -73.835 -75.945 -73.555 ;
        RECT -76.225 -74.435 -75.945 -74.155 ;
        RECT -67.265 -73.835 -66.985 -73.555 ;
        RECT -67.265 -74.435 -66.985 -74.155 ;
        RECT -58.305 -73.835 -58.025 -73.555 ;
        RECT -58.305 -74.435 -58.025 -74.155 ;
        RECT -49.345 -73.835 -49.065 -73.555 ;
        RECT -49.345 -74.435 -49.065 -74.155 ;
        RECT -40.385 -73.835 -40.105 -73.555 ;
        RECT -40.385 -74.435 -40.105 -74.155 ;
        RECT -31.425 -73.835 -31.145 -73.555 ;
        RECT -31.425 -74.435 -31.145 -74.155 ;
        RECT -22.465 -73.835 -22.185 -73.555 ;
        RECT -22.465 -74.435 -22.185 -74.155 ;
        RECT -13.505 -73.835 -13.225 -73.555 ;
        RECT -13.505 -74.435 -13.225 -74.155 ;
        RECT -4.545 -73.835 -4.265 -73.555 ;
        RECT -4.545 -74.435 -4.265 -74.155 ;
        RECT 4.415 -73.835 4.695 -73.555 ;
        RECT 4.415 -74.435 4.695 -74.155 ;
        RECT 13.375 -73.835 13.655 -73.555 ;
        RECT 13.375 -74.435 13.655 -74.155 ;
        RECT 22.335 -73.835 22.615 -73.555 ;
        RECT 22.335 -74.435 22.615 -74.155 ;
        RECT 31.295 -73.835 31.575 -73.555 ;
        RECT 31.295 -74.435 31.575 -74.155 ;
        RECT 40.255 -73.835 40.535 -73.555 ;
        RECT 40.255 -74.435 40.535 -74.155 ;
        RECT 49.215 -73.835 49.495 -73.555 ;
        RECT 49.215 -74.435 49.495 -74.155 ;
        RECT 58.175 -73.835 58.455 -73.555 ;
        RECT 58.175 -74.435 58.455 -74.155 ;
        RECT 67.135 -73.835 67.415 -73.555 ;
        RECT 67.135 -74.435 67.415 -74.155 ;
        RECT 76.095 -73.835 76.375 -73.555 ;
        RECT 76.095 -74.435 76.375 -74.155 ;
        RECT 85.055 -73.835 85.335 -73.555 ;
        RECT 85.055 -74.435 85.335 -74.155 ;
        RECT 94.015 -73.835 94.295 -73.555 ;
        RECT 94.015 -74.435 94.295 -74.155 ;
        RECT 104.915 -74.135 105.195 -73.855 ;
        RECT 105.515 -74.135 105.795 -73.855 ;
        RECT -467.105 -77.195 -466.825 -76.915 ;
        RECT -467.105 -77.795 -466.825 -77.515 ;
        RECT -449.185 -77.195 -448.905 -76.915 ;
        RECT -449.185 -77.795 -448.905 -77.515 ;
        RECT -431.265 -77.195 -430.985 -76.915 ;
        RECT -431.265 -77.795 -430.985 -77.515 ;
        RECT -413.345 -77.195 -413.065 -76.915 ;
        RECT -413.345 -77.795 -413.065 -77.515 ;
        RECT -395.425 -77.195 -395.145 -76.915 ;
        RECT -395.425 -77.795 -395.145 -77.515 ;
        RECT -377.505 -77.195 -377.225 -76.915 ;
        RECT -377.505 -77.795 -377.225 -77.515 ;
        RECT -359.585 -77.195 -359.305 -76.915 ;
        RECT -359.585 -77.795 -359.305 -77.515 ;
        RECT -341.665 -77.195 -341.385 -76.915 ;
        RECT -341.665 -77.795 -341.385 -77.515 ;
        RECT -323.745 -77.195 -323.465 -76.915 ;
        RECT -323.745 -77.795 -323.465 -77.515 ;
        RECT -305.825 -77.195 -305.545 -76.915 ;
        RECT -305.825 -77.795 -305.545 -77.515 ;
        RECT -287.905 -77.195 -287.625 -76.915 ;
        RECT -287.905 -77.795 -287.625 -77.515 ;
        RECT -269.985 -77.195 -269.705 -76.915 ;
        RECT -269.985 -77.795 -269.705 -77.515 ;
        RECT -252.065 -77.195 -251.785 -76.915 ;
        RECT -252.065 -77.795 -251.785 -77.515 ;
        RECT -234.145 -77.195 -233.865 -76.915 ;
        RECT -234.145 -77.795 -233.865 -77.515 ;
        RECT -216.225 -77.195 -215.945 -76.915 ;
        RECT -216.225 -77.795 -215.945 -77.515 ;
        RECT -198.305 -77.195 -198.025 -76.915 ;
        RECT -198.305 -77.795 -198.025 -77.515 ;
        RECT -179.265 -77.195 -178.985 -76.915 ;
        RECT -179.265 -77.795 -178.985 -77.515 ;
        RECT -161.345 -77.195 -161.065 -76.915 ;
        RECT -161.345 -77.795 -161.065 -77.515 ;
        RECT -143.425 -77.195 -143.145 -76.915 ;
        RECT -143.425 -77.795 -143.145 -77.515 ;
        RECT -125.505 -77.195 -125.225 -76.915 ;
        RECT -125.505 -77.795 -125.225 -77.515 ;
        RECT -107.585 -77.195 -107.305 -76.915 ;
        RECT -107.585 -77.795 -107.305 -77.515 ;
        RECT -89.665 -77.195 -89.385 -76.915 ;
        RECT -89.665 -77.795 -89.385 -77.515 ;
        RECT -71.745 -77.195 -71.465 -76.915 ;
        RECT -71.745 -77.795 -71.465 -77.515 ;
        RECT -53.825 -77.195 -53.545 -76.915 ;
        RECT -53.825 -77.795 -53.545 -77.515 ;
        RECT -35.905 -77.195 -35.625 -76.915 ;
        RECT -35.905 -77.795 -35.625 -77.515 ;
        RECT -17.985 -77.195 -17.705 -76.915 ;
        RECT -17.985 -77.795 -17.705 -77.515 ;
        RECT -0.065 -77.195 0.215 -76.915 ;
        RECT -0.065 -77.795 0.215 -77.515 ;
        RECT 17.855 -77.195 18.135 -76.915 ;
        RECT 17.855 -77.795 18.135 -77.515 ;
        RECT 35.775 -77.195 36.055 -76.915 ;
        RECT 35.775 -77.795 36.055 -77.515 ;
        RECT 53.695 -77.195 53.975 -76.915 ;
        RECT 53.695 -77.795 53.975 -77.515 ;
        RECT 71.615 -77.195 71.895 -76.915 ;
        RECT 71.615 -77.795 71.895 -77.515 ;
        RECT 89.535 -77.195 89.815 -76.915 ;
        RECT 89.535 -77.795 89.815 -77.515 ;
        RECT 106.715 -77.495 106.995 -77.215 ;
        RECT 107.315 -77.495 107.595 -77.215 ;
        RECT -458.145 -80.555 -457.865 -80.275 ;
        RECT -458.145 -81.155 -457.865 -80.875 ;
        RECT -486.895 -83.115 -486.615 -81.275 ;
        RECT -422.305 -80.555 -422.025 -80.275 ;
        RECT -422.305 -81.155 -422.025 -80.875 ;
        RECT -386.465 -80.555 -386.185 -80.275 ;
        RECT -386.465 -81.155 -386.185 -80.875 ;
        RECT -350.625 -80.555 -350.345 -80.275 ;
        RECT -350.625 -81.155 -350.345 -80.875 ;
        RECT -314.785 -80.555 -314.505 -80.275 ;
        RECT -314.785 -81.155 -314.505 -80.875 ;
        RECT -278.945 -80.555 -278.665 -80.275 ;
        RECT -278.945 -81.155 -278.665 -80.875 ;
        RECT -243.105 -80.555 -242.825 -80.275 ;
        RECT -243.105 -81.155 -242.825 -80.875 ;
        RECT -207.265 -80.555 -206.985 -80.275 ;
        RECT -207.265 -81.155 -206.985 -80.875 ;
        RECT -170.305 -80.555 -170.025 -80.275 ;
        RECT -170.305 -81.155 -170.025 -80.875 ;
        RECT -134.465 -80.555 -134.185 -80.275 ;
        RECT -134.465 -81.155 -134.185 -80.875 ;
        RECT -98.625 -80.555 -98.345 -80.275 ;
        RECT -98.625 -81.155 -98.345 -80.875 ;
        RECT -62.785 -80.555 -62.505 -80.275 ;
        RECT -62.785 -81.155 -62.505 -80.875 ;
        RECT -26.945 -80.555 -26.665 -80.275 ;
        RECT -26.945 -81.155 -26.665 -80.875 ;
        RECT 8.895 -80.555 9.175 -80.275 ;
        RECT 8.895 -81.155 9.175 -80.875 ;
        RECT 44.735 -80.555 45.015 -80.275 ;
        RECT 44.735 -81.155 45.015 -80.875 ;
        RECT 80.575 -80.555 80.855 -80.275 ;
        RECT 80.575 -81.155 80.855 -80.875 ;
        RECT 108.515 -80.855 108.795 -80.575 ;
        RECT 109.115 -80.855 109.395 -80.575 ;
        RECT -497.475 -83.705 -495.635 -83.425 ;
        RECT -440.225 -83.915 -439.945 -83.635 ;
        RECT -440.225 -84.515 -439.945 -84.235 ;
        RECT -368.545 -83.915 -368.265 -83.635 ;
        RECT -368.545 -84.515 -368.265 -84.235 ;
        RECT -296.865 -83.915 -296.585 -83.635 ;
        RECT -296.865 -84.515 -296.585 -84.235 ;
        RECT -225.185 -83.915 -224.905 -83.635 ;
        RECT -225.185 -84.515 -224.905 -84.235 ;
        RECT -152.385 -83.915 -152.105 -83.635 ;
        RECT -152.385 -84.515 -152.105 -84.235 ;
        RECT -80.705 -83.915 -80.425 -83.635 ;
        RECT -80.705 -84.515 -80.425 -84.235 ;
        RECT -9.025 -83.915 -8.745 -83.635 ;
        RECT -9.025 -84.515 -8.745 -84.235 ;
        RECT 62.655 -83.915 62.935 -83.635 ;
        RECT 62.655 -84.515 62.935 -84.235 ;
        RECT 110.315 -84.215 110.595 -83.935 ;
        RECT 110.915 -84.215 111.195 -83.935 ;
        RECT -404.385 -87.275 -404.105 -86.995 ;
        RECT -404.385 -87.875 -404.105 -87.595 ;
        RECT -261.025 -87.275 -260.745 -86.995 ;
        RECT -261.025 -87.875 -260.745 -87.595 ;
        RECT -116.545 -87.275 -116.265 -86.995 ;
        RECT -116.545 -87.875 -116.265 -87.595 ;
        RECT 26.815 -87.275 27.095 -86.995 ;
        RECT 26.815 -87.875 27.095 -87.595 ;
        RECT 112.115 -87.575 112.395 -87.295 ;
        RECT 112.715 -87.575 112.995 -87.295 ;
        RECT -332.705 -90.635 -332.425 -90.355 ;
        RECT -332.705 -91.235 -332.425 -90.955 ;
        RECT -44.865 -90.635 -44.585 -90.355 ;
        RECT -44.865 -91.235 -44.585 -90.955 ;
        RECT 113.915 -90.935 114.195 -90.655 ;
        RECT 114.515 -90.935 114.795 -90.655 ;
        RECT -188.225 -93.995 -187.945 -93.715 ;
        RECT 121.025 -64.055 121.825 -63.775 ;
        RECT 121.025 -67.415 121.825 -67.135 ;
        RECT 121.025 -70.775 121.825 -70.495 ;
        RECT 121.025 -74.135 121.825 -73.855 ;
        RECT 121.025 -77.495 121.825 -77.215 ;
        RECT 121.025 -80.855 121.825 -80.575 ;
        RECT 121.025 -84.215 121.825 -83.935 ;
        RECT 121.025 -87.575 121.825 -87.295 ;
        RECT 121.025 -90.935 121.825 -90.655 ;
        RECT -188.225 -94.595 -187.945 -94.315 ;
        RECT 115.715 -94.295 115.995 -94.015 ;
        RECT 116.315 -94.295 116.595 -94.015 ;
        RECT 121.025 -94.295 121.825 -94.015 ;
        RECT -189.345 -97.355 -189.065 -97.075 ;
        RECT -189.345 -97.955 -189.065 -97.675 ;
        RECT 121.025 -97.655 121.825 -97.375 ;
      LAYER Metal4 ;
        RECT -189.405 97.765 -189.005 98.115 ;
        RECT -189.405 97.265 121.925 97.765 ;
        RECT -189.405 96.915 -189.005 97.265 ;
        RECT -188.285 94.405 -187.885 94.755 ;
        RECT -188.285 93.905 121.925 94.405 ;
        RECT -188.285 93.555 -187.885 93.905 ;
        RECT -332.765 91.045 -332.365 91.395 ;
        RECT -44.925 91.045 -44.525 91.395 ;
        RECT -332.765 90.545 121.925 91.045 ;
        RECT -332.765 90.195 -332.365 90.545 ;
        RECT -44.925 90.195 -44.525 90.545 ;
        RECT -404.445 87.685 -404.045 88.035 ;
        RECT -261.085 87.685 -260.685 88.035 ;
        RECT -116.605 87.685 -116.205 88.035 ;
        RECT 26.755 87.685 27.155 88.035 ;
        RECT -404.445 87.185 121.925 87.685 ;
        RECT -404.445 86.835 -404.045 87.185 ;
        RECT -261.085 86.835 -260.685 87.185 ;
        RECT -116.605 86.835 -116.205 87.185 ;
        RECT 26.755 86.835 27.155 87.185 ;
        RECT -440.285 84.325 -439.885 84.675 ;
        RECT -368.605 84.325 -368.205 84.675 ;
        RECT -296.925 84.325 -296.525 84.675 ;
        RECT -225.245 84.325 -224.845 84.675 ;
        RECT -152.445 84.325 -152.045 84.675 ;
        RECT -80.765 84.325 -80.365 84.675 ;
        RECT -9.085 84.325 -8.685 84.675 ;
        RECT 62.595 84.325 62.995 84.675 ;
        RECT -440.285 83.825 121.925 84.325 ;
        RECT -497.595 83.365 -495.515 83.765 ;
        RECT -440.285 83.475 -439.885 83.825 ;
        RECT -368.605 83.475 -368.205 83.825 ;
        RECT -296.925 83.475 -296.525 83.825 ;
        RECT -225.245 83.475 -224.845 83.825 ;
        RECT -152.445 83.475 -152.045 83.825 ;
        RECT -80.765 83.475 -80.365 83.825 ;
        RECT -9.085 83.475 -8.685 83.825 ;
        RECT 62.595 83.475 62.995 83.825 ;
        RECT -486.955 81.155 -486.555 83.235 ;
        RECT -458.205 80.965 -457.805 81.315 ;
        RECT -422.365 80.965 -421.965 81.315 ;
        RECT -386.525 80.965 -386.125 81.315 ;
        RECT -350.685 80.965 -350.285 81.315 ;
        RECT -314.845 80.965 -314.445 81.315 ;
        RECT -279.005 80.965 -278.605 81.315 ;
        RECT -243.165 80.965 -242.765 81.315 ;
        RECT -207.325 80.965 -206.925 81.315 ;
        RECT -170.365 80.965 -169.965 81.315 ;
        RECT -134.525 80.965 -134.125 81.315 ;
        RECT -98.685 80.965 -98.285 81.315 ;
        RECT -62.845 80.965 -62.445 81.315 ;
        RECT -27.005 80.965 -26.605 81.315 ;
        RECT 8.835 80.965 9.235 81.315 ;
        RECT 44.675 80.965 45.075 81.315 ;
        RECT 80.515 80.965 80.915 81.315 ;
        RECT -458.205 80.465 121.925 80.965 ;
        RECT -458.205 80.115 -457.805 80.465 ;
        RECT -422.365 80.115 -421.965 80.465 ;
        RECT -386.525 80.115 -386.125 80.465 ;
        RECT -350.685 80.115 -350.285 80.465 ;
        RECT -314.845 80.115 -314.445 80.465 ;
        RECT -279.005 80.115 -278.605 80.465 ;
        RECT -243.165 80.115 -242.765 80.465 ;
        RECT -207.325 80.115 -206.925 80.465 ;
        RECT -170.365 80.115 -169.965 80.465 ;
        RECT -134.525 80.115 -134.125 80.465 ;
        RECT -98.685 80.115 -98.285 80.465 ;
        RECT -62.845 80.115 -62.445 80.465 ;
        RECT -27.005 80.115 -26.605 80.465 ;
        RECT 8.835 80.115 9.235 80.465 ;
        RECT 44.675 80.115 45.075 80.465 ;
        RECT 80.515 80.115 80.915 80.465 ;
        RECT -497.305 78.300 -486.905 78.900 ;
        RECT -497.305 70.300 -495.505 78.300 ;
        RECT -487.505 70.300 -486.905 78.300 ;
        RECT -467.165 77.605 -466.765 77.955 ;
        RECT -449.245 77.605 -448.845 77.955 ;
        RECT -431.325 77.605 -430.925 77.955 ;
        RECT -413.405 77.605 -413.005 77.955 ;
        RECT -395.485 77.605 -395.085 77.955 ;
        RECT -377.565 77.605 -377.165 77.955 ;
        RECT -359.645 77.605 -359.245 77.955 ;
        RECT -341.725 77.605 -341.325 77.955 ;
        RECT -323.805 77.605 -323.405 77.955 ;
        RECT -305.885 77.605 -305.485 77.955 ;
        RECT -287.965 77.605 -287.565 77.955 ;
        RECT -270.045 77.605 -269.645 77.955 ;
        RECT -252.125 77.605 -251.725 77.955 ;
        RECT -234.205 77.605 -233.805 77.955 ;
        RECT -216.285 77.605 -215.885 77.955 ;
        RECT -198.365 77.605 -197.965 77.955 ;
        RECT -179.325 77.605 -178.925 77.955 ;
        RECT -161.405 77.605 -161.005 77.955 ;
        RECT -143.485 77.605 -143.085 77.955 ;
        RECT -125.565 77.605 -125.165 77.955 ;
        RECT -107.645 77.605 -107.245 77.955 ;
        RECT -89.725 77.605 -89.325 77.955 ;
        RECT -71.805 77.605 -71.405 77.955 ;
        RECT -53.885 77.605 -53.485 77.955 ;
        RECT -35.965 77.605 -35.565 77.955 ;
        RECT -18.045 77.605 -17.645 77.955 ;
        RECT -0.125 77.605 0.275 77.955 ;
        RECT 17.795 77.605 18.195 77.955 ;
        RECT 35.715 77.605 36.115 77.955 ;
        RECT 53.635 77.605 54.035 77.955 ;
        RECT 71.555 77.605 71.955 77.955 ;
        RECT 89.475 77.605 89.875 77.955 ;
        RECT -467.165 77.105 121.925 77.605 ;
        RECT -467.165 76.755 -466.765 77.105 ;
        RECT -449.245 76.755 -448.845 77.105 ;
        RECT -431.325 76.755 -430.925 77.105 ;
        RECT -413.405 76.755 -413.005 77.105 ;
        RECT -395.485 76.755 -395.085 77.105 ;
        RECT -377.565 76.755 -377.165 77.105 ;
        RECT -359.645 76.755 -359.245 77.105 ;
        RECT -341.725 76.755 -341.325 77.105 ;
        RECT -323.805 76.755 -323.405 77.105 ;
        RECT -305.885 76.755 -305.485 77.105 ;
        RECT -287.965 76.755 -287.565 77.105 ;
        RECT -270.045 76.755 -269.645 77.105 ;
        RECT -252.125 76.755 -251.725 77.105 ;
        RECT -234.205 76.755 -233.805 77.105 ;
        RECT -216.285 76.755 -215.885 77.105 ;
        RECT -198.365 76.755 -197.965 77.105 ;
        RECT -179.325 76.755 -178.925 77.105 ;
        RECT -161.405 76.755 -161.005 77.105 ;
        RECT -143.485 76.755 -143.085 77.105 ;
        RECT -125.565 76.755 -125.165 77.105 ;
        RECT -107.645 76.755 -107.245 77.105 ;
        RECT -89.725 76.755 -89.325 77.105 ;
        RECT -71.805 76.755 -71.405 77.105 ;
        RECT -53.885 76.755 -53.485 77.105 ;
        RECT -35.965 76.755 -35.565 77.105 ;
        RECT -18.045 76.755 -17.645 77.105 ;
        RECT -0.125 76.755 0.275 77.105 ;
        RECT 17.795 76.755 18.195 77.105 ;
        RECT 35.715 76.755 36.115 77.105 ;
        RECT 53.635 76.755 54.035 77.105 ;
        RECT 71.555 76.755 71.955 77.105 ;
        RECT 89.475 76.755 89.875 77.105 ;
        RECT -471.645 74.245 -471.245 74.595 ;
        RECT -462.685 74.245 -462.285 74.595 ;
        RECT -453.725 74.245 -453.325 74.595 ;
        RECT -444.765 74.245 -444.365 74.595 ;
        RECT -435.805 74.245 -435.405 74.595 ;
        RECT -426.845 74.245 -426.445 74.595 ;
        RECT -417.885 74.245 -417.485 74.595 ;
        RECT -408.925 74.245 -408.525 74.595 ;
        RECT -399.965 74.245 -399.565 74.595 ;
        RECT -391.005 74.245 -390.605 74.595 ;
        RECT -382.045 74.245 -381.645 74.595 ;
        RECT -373.085 74.245 -372.685 74.595 ;
        RECT -364.125 74.245 -363.725 74.595 ;
        RECT -355.165 74.245 -354.765 74.595 ;
        RECT -346.205 74.245 -345.805 74.595 ;
        RECT -337.245 74.245 -336.845 74.595 ;
        RECT -328.285 74.245 -327.885 74.595 ;
        RECT -319.325 74.245 -318.925 74.595 ;
        RECT -310.365 74.245 -309.965 74.595 ;
        RECT -301.405 74.245 -301.005 74.595 ;
        RECT -292.445 74.245 -292.045 74.595 ;
        RECT -283.485 74.245 -283.085 74.595 ;
        RECT -274.525 74.245 -274.125 74.595 ;
        RECT -265.565 74.245 -265.165 74.595 ;
        RECT -256.605 74.245 -256.205 74.595 ;
        RECT -247.645 74.245 -247.245 74.595 ;
        RECT -238.685 74.245 -238.285 74.595 ;
        RECT -229.725 74.245 -229.325 74.595 ;
        RECT -220.765 74.245 -220.365 74.595 ;
        RECT -211.805 74.245 -211.405 74.595 ;
        RECT -202.845 74.245 -202.445 74.595 ;
        RECT -193.885 74.245 -193.485 74.595 ;
        RECT -183.805 74.245 -183.405 74.595 ;
        RECT -174.845 74.245 -174.445 74.595 ;
        RECT -165.885 74.245 -165.485 74.595 ;
        RECT -156.925 74.245 -156.525 74.595 ;
        RECT -147.965 74.245 -147.565 74.595 ;
        RECT -139.005 74.245 -138.605 74.595 ;
        RECT -130.045 74.245 -129.645 74.595 ;
        RECT -121.085 74.245 -120.685 74.595 ;
        RECT -112.125 74.245 -111.725 74.595 ;
        RECT -103.165 74.245 -102.765 74.595 ;
        RECT -94.205 74.245 -93.805 74.595 ;
        RECT -85.245 74.245 -84.845 74.595 ;
        RECT -76.285 74.245 -75.885 74.595 ;
        RECT -67.325 74.245 -66.925 74.595 ;
        RECT -58.365 74.245 -57.965 74.595 ;
        RECT -49.405 74.245 -49.005 74.595 ;
        RECT -40.445 74.245 -40.045 74.595 ;
        RECT -31.485 74.245 -31.085 74.595 ;
        RECT -22.525 74.245 -22.125 74.595 ;
        RECT -13.565 74.245 -13.165 74.595 ;
        RECT -4.605 74.245 -4.205 74.595 ;
        RECT 4.355 74.245 4.755 74.595 ;
        RECT 13.315 74.245 13.715 74.595 ;
        RECT 22.275 74.245 22.675 74.595 ;
        RECT 31.235 74.245 31.635 74.595 ;
        RECT 40.195 74.245 40.595 74.595 ;
        RECT 49.155 74.245 49.555 74.595 ;
        RECT 58.115 74.245 58.515 74.595 ;
        RECT 67.075 74.245 67.475 74.595 ;
        RECT 76.035 74.245 76.435 74.595 ;
        RECT 84.995 74.245 85.395 74.595 ;
        RECT 93.955 74.245 94.355 74.595 ;
        RECT -471.645 73.745 121.925 74.245 ;
        RECT -471.645 73.395 -471.245 73.745 ;
        RECT -462.685 73.395 -462.285 73.745 ;
        RECT -453.725 73.395 -453.325 73.745 ;
        RECT -444.765 73.395 -444.365 73.745 ;
        RECT -435.805 73.395 -435.405 73.745 ;
        RECT -426.845 73.395 -426.445 73.745 ;
        RECT -417.885 73.395 -417.485 73.745 ;
        RECT -408.925 73.395 -408.525 73.745 ;
        RECT -399.965 73.395 -399.565 73.745 ;
        RECT -391.005 73.395 -390.605 73.745 ;
        RECT -382.045 73.395 -381.645 73.745 ;
        RECT -373.085 73.395 -372.685 73.745 ;
        RECT -364.125 73.395 -363.725 73.745 ;
        RECT -355.165 73.395 -354.765 73.745 ;
        RECT -346.205 73.395 -345.805 73.745 ;
        RECT -337.245 73.395 -336.845 73.745 ;
        RECT -328.285 73.395 -327.885 73.745 ;
        RECT -319.325 73.395 -318.925 73.745 ;
        RECT -310.365 73.395 -309.965 73.745 ;
        RECT -301.405 73.395 -301.005 73.745 ;
        RECT -292.445 73.395 -292.045 73.745 ;
        RECT -283.485 73.395 -283.085 73.745 ;
        RECT -274.525 73.395 -274.125 73.745 ;
        RECT -265.565 73.395 -265.165 73.745 ;
        RECT -256.605 73.395 -256.205 73.745 ;
        RECT -247.645 73.395 -247.245 73.745 ;
        RECT -238.685 73.395 -238.285 73.745 ;
        RECT -229.725 73.395 -229.325 73.745 ;
        RECT -220.765 73.395 -220.365 73.745 ;
        RECT -211.805 73.395 -211.405 73.745 ;
        RECT -202.845 73.395 -202.445 73.745 ;
        RECT -193.885 73.395 -193.485 73.745 ;
        RECT -183.805 73.395 -183.405 73.745 ;
        RECT -174.845 73.395 -174.445 73.745 ;
        RECT -165.885 73.395 -165.485 73.745 ;
        RECT -156.925 73.395 -156.525 73.745 ;
        RECT -147.965 73.395 -147.565 73.745 ;
        RECT -139.005 73.395 -138.605 73.745 ;
        RECT -130.045 73.395 -129.645 73.745 ;
        RECT -121.085 73.395 -120.685 73.745 ;
        RECT -112.125 73.395 -111.725 73.745 ;
        RECT -103.165 73.395 -102.765 73.745 ;
        RECT -94.205 73.395 -93.805 73.745 ;
        RECT -85.245 73.395 -84.845 73.745 ;
        RECT -76.285 73.395 -75.885 73.745 ;
        RECT -67.325 73.395 -66.925 73.745 ;
        RECT -58.365 73.395 -57.965 73.745 ;
        RECT -49.405 73.395 -49.005 73.745 ;
        RECT -40.445 73.395 -40.045 73.745 ;
        RECT -31.485 73.395 -31.085 73.745 ;
        RECT -22.525 73.395 -22.125 73.745 ;
        RECT -13.565 73.395 -13.165 73.745 ;
        RECT -4.605 73.395 -4.205 73.745 ;
        RECT 4.355 73.395 4.755 73.745 ;
        RECT 13.315 73.395 13.715 73.745 ;
        RECT 22.275 73.395 22.675 73.745 ;
        RECT 31.235 73.395 31.635 73.745 ;
        RECT 40.195 73.395 40.595 73.745 ;
        RECT 49.155 73.395 49.555 73.745 ;
        RECT 58.115 73.395 58.515 73.745 ;
        RECT 67.075 73.395 67.475 73.745 ;
        RECT 76.035 73.395 76.435 73.745 ;
        RECT 84.995 73.395 85.395 73.745 ;
        RECT 93.955 73.395 94.355 73.745 ;
        RECT -497.305 69.700 -486.905 70.300 ;
        RECT -473.885 70.885 -473.485 71.235 ;
        RECT -469.405 70.885 -469.005 71.235 ;
        RECT -464.925 70.885 -464.525 71.235 ;
        RECT -460.445 70.885 -460.045 71.235 ;
        RECT -455.965 70.885 -455.565 71.235 ;
        RECT -451.485 70.885 -451.085 71.235 ;
        RECT -447.005 70.885 -446.605 71.235 ;
        RECT -442.525 70.885 -442.125 71.235 ;
        RECT -438.045 70.885 -437.645 71.235 ;
        RECT -433.565 70.885 -433.165 71.235 ;
        RECT -429.085 70.885 -428.685 71.235 ;
        RECT -424.605 70.885 -424.205 71.235 ;
        RECT -420.125 70.885 -419.725 71.235 ;
        RECT -415.645 70.885 -415.245 71.235 ;
        RECT -411.165 70.885 -410.765 71.235 ;
        RECT -406.685 70.885 -406.285 71.235 ;
        RECT -402.205 70.885 -401.805 71.235 ;
        RECT -397.725 70.885 -397.325 71.235 ;
        RECT -393.245 70.885 -392.845 71.235 ;
        RECT -388.765 70.885 -388.365 71.235 ;
        RECT -384.285 70.885 -383.885 71.235 ;
        RECT -379.805 70.885 -379.405 71.235 ;
        RECT -375.325 70.885 -374.925 71.235 ;
        RECT -370.845 70.885 -370.445 71.235 ;
        RECT -366.365 70.885 -365.965 71.235 ;
        RECT -361.885 70.885 -361.485 71.235 ;
        RECT -357.405 70.885 -357.005 71.235 ;
        RECT -352.925 70.885 -352.525 71.235 ;
        RECT -348.445 70.885 -348.045 71.235 ;
        RECT -343.965 70.885 -343.565 71.235 ;
        RECT -339.485 70.885 -339.085 71.235 ;
        RECT -335.005 70.885 -334.605 71.235 ;
        RECT -330.525 70.885 -330.125 71.235 ;
        RECT -326.045 70.885 -325.645 71.235 ;
        RECT -321.565 70.885 -321.165 71.235 ;
        RECT -317.085 70.885 -316.685 71.235 ;
        RECT -312.605 70.885 -312.205 71.235 ;
        RECT -308.125 70.885 -307.725 71.235 ;
        RECT -303.645 70.885 -303.245 71.235 ;
        RECT -299.165 70.885 -298.765 71.235 ;
        RECT -294.685 70.885 -294.285 71.235 ;
        RECT -290.205 70.885 -289.805 71.235 ;
        RECT -285.725 70.885 -285.325 71.235 ;
        RECT -281.245 70.885 -280.845 71.235 ;
        RECT -276.765 70.885 -276.365 71.235 ;
        RECT -272.285 70.885 -271.885 71.235 ;
        RECT -267.805 70.885 -267.405 71.235 ;
        RECT -263.325 70.885 -262.925 71.235 ;
        RECT -258.845 70.885 -258.445 71.235 ;
        RECT -254.365 70.885 -253.965 71.235 ;
        RECT -249.885 70.885 -249.485 71.235 ;
        RECT -245.405 70.885 -245.005 71.235 ;
        RECT -240.925 70.885 -240.525 71.235 ;
        RECT -236.445 70.885 -236.045 71.235 ;
        RECT -231.965 70.885 -231.565 71.235 ;
        RECT -227.485 70.885 -227.085 71.235 ;
        RECT -223.005 70.885 -222.605 71.235 ;
        RECT -218.525 70.885 -218.125 71.235 ;
        RECT -214.045 70.885 -213.645 71.235 ;
        RECT -209.565 70.885 -209.165 71.235 ;
        RECT -205.085 70.885 -204.685 71.235 ;
        RECT -200.605 70.885 -200.205 71.235 ;
        RECT -196.125 70.885 -195.725 71.235 ;
        RECT -191.645 70.885 -191.245 71.235 ;
        RECT -186.045 70.885 -185.645 71.235 ;
        RECT -181.565 70.885 -181.165 71.235 ;
        RECT -177.085 70.885 -176.685 71.235 ;
        RECT -172.605 70.885 -172.205 71.235 ;
        RECT -168.125 70.885 -167.725 71.235 ;
        RECT -163.645 70.885 -163.245 71.235 ;
        RECT -159.165 70.885 -158.765 71.235 ;
        RECT -154.685 70.885 -154.285 71.235 ;
        RECT -150.205 70.885 -149.805 71.235 ;
        RECT -145.725 70.885 -145.325 71.235 ;
        RECT -141.245 70.885 -140.845 71.235 ;
        RECT -136.765 70.885 -136.365 71.235 ;
        RECT -132.285 70.885 -131.885 71.235 ;
        RECT -127.805 70.885 -127.405 71.235 ;
        RECT -123.325 70.885 -122.925 71.235 ;
        RECT -118.845 70.885 -118.445 71.235 ;
        RECT -114.365 70.885 -113.965 71.235 ;
        RECT -109.885 70.885 -109.485 71.235 ;
        RECT -105.405 70.885 -105.005 71.235 ;
        RECT -100.925 70.885 -100.525 71.235 ;
        RECT -96.445 70.885 -96.045 71.235 ;
        RECT -91.965 70.885 -91.565 71.235 ;
        RECT -87.485 70.885 -87.085 71.235 ;
        RECT -83.005 70.885 -82.605 71.235 ;
        RECT -78.525 70.885 -78.125 71.235 ;
        RECT -74.045 70.885 -73.645 71.235 ;
        RECT -69.565 70.885 -69.165 71.235 ;
        RECT -65.085 70.885 -64.685 71.235 ;
        RECT -60.605 70.885 -60.205 71.235 ;
        RECT -56.125 70.885 -55.725 71.235 ;
        RECT -51.645 70.885 -51.245 71.235 ;
        RECT -47.165 70.885 -46.765 71.235 ;
        RECT -42.685 70.885 -42.285 71.235 ;
        RECT -38.205 70.885 -37.805 71.235 ;
        RECT -33.725 70.885 -33.325 71.235 ;
        RECT -29.245 70.885 -28.845 71.235 ;
        RECT -24.765 70.885 -24.365 71.235 ;
        RECT -20.285 70.885 -19.885 71.235 ;
        RECT -15.805 70.885 -15.405 71.235 ;
        RECT -11.325 70.885 -10.925 71.235 ;
        RECT -6.845 70.885 -6.445 71.235 ;
        RECT -2.365 70.885 -1.965 71.235 ;
        RECT 2.115 70.885 2.515 71.235 ;
        RECT 6.595 70.885 6.995 71.235 ;
        RECT 11.075 70.885 11.475 71.235 ;
        RECT 15.555 70.885 15.955 71.235 ;
        RECT 20.035 70.885 20.435 71.235 ;
        RECT 24.515 70.885 24.915 71.235 ;
        RECT 28.995 70.885 29.395 71.235 ;
        RECT 33.475 70.885 33.875 71.235 ;
        RECT 37.955 70.885 38.355 71.235 ;
        RECT 42.435 70.885 42.835 71.235 ;
        RECT 46.915 70.885 47.315 71.235 ;
        RECT 51.395 70.885 51.795 71.235 ;
        RECT 55.875 70.885 56.275 71.235 ;
        RECT 60.355 70.885 60.755 71.235 ;
        RECT 64.835 70.885 65.235 71.235 ;
        RECT 69.315 70.885 69.715 71.235 ;
        RECT 73.795 70.885 74.195 71.235 ;
        RECT 78.275 70.885 78.675 71.235 ;
        RECT 82.755 70.885 83.155 71.235 ;
        RECT 87.235 70.885 87.635 71.235 ;
        RECT 91.715 70.885 92.115 71.235 ;
        RECT 96.195 70.885 96.595 71.235 ;
        RECT -473.885 70.385 121.925 70.885 ;
        RECT -473.885 70.035 -473.485 70.385 ;
        RECT -469.405 70.035 -469.005 70.385 ;
        RECT -464.925 70.035 -464.525 70.385 ;
        RECT -460.445 70.035 -460.045 70.385 ;
        RECT -455.965 70.035 -455.565 70.385 ;
        RECT -451.485 70.035 -451.085 70.385 ;
        RECT -447.005 70.035 -446.605 70.385 ;
        RECT -442.525 70.035 -442.125 70.385 ;
        RECT -438.045 70.035 -437.645 70.385 ;
        RECT -433.565 70.035 -433.165 70.385 ;
        RECT -429.085 70.035 -428.685 70.385 ;
        RECT -424.605 70.035 -424.205 70.385 ;
        RECT -420.125 70.035 -419.725 70.385 ;
        RECT -415.645 70.035 -415.245 70.385 ;
        RECT -411.165 70.035 -410.765 70.385 ;
        RECT -406.685 70.035 -406.285 70.385 ;
        RECT -402.205 70.035 -401.805 70.385 ;
        RECT -397.725 70.035 -397.325 70.385 ;
        RECT -393.245 70.035 -392.845 70.385 ;
        RECT -388.765 70.035 -388.365 70.385 ;
        RECT -384.285 70.035 -383.885 70.385 ;
        RECT -379.805 70.035 -379.405 70.385 ;
        RECT -375.325 70.035 -374.925 70.385 ;
        RECT -370.845 70.035 -370.445 70.385 ;
        RECT -366.365 70.035 -365.965 70.385 ;
        RECT -361.885 70.035 -361.485 70.385 ;
        RECT -357.405 70.035 -357.005 70.385 ;
        RECT -352.925 70.035 -352.525 70.385 ;
        RECT -348.445 70.035 -348.045 70.385 ;
        RECT -343.965 70.035 -343.565 70.385 ;
        RECT -339.485 70.035 -339.085 70.385 ;
        RECT -335.005 70.035 -334.605 70.385 ;
        RECT -330.525 70.035 -330.125 70.385 ;
        RECT -326.045 70.035 -325.645 70.385 ;
        RECT -321.565 70.035 -321.165 70.385 ;
        RECT -317.085 70.035 -316.685 70.385 ;
        RECT -312.605 70.035 -312.205 70.385 ;
        RECT -308.125 70.035 -307.725 70.385 ;
        RECT -303.645 70.035 -303.245 70.385 ;
        RECT -299.165 70.035 -298.765 70.385 ;
        RECT -294.685 70.035 -294.285 70.385 ;
        RECT -290.205 70.035 -289.805 70.385 ;
        RECT -285.725 70.035 -285.325 70.385 ;
        RECT -281.245 70.035 -280.845 70.385 ;
        RECT -276.765 70.035 -276.365 70.385 ;
        RECT -272.285 70.035 -271.885 70.385 ;
        RECT -267.805 70.035 -267.405 70.385 ;
        RECT -263.325 70.035 -262.925 70.385 ;
        RECT -258.845 70.035 -258.445 70.385 ;
        RECT -254.365 70.035 -253.965 70.385 ;
        RECT -249.885 70.035 -249.485 70.385 ;
        RECT -245.405 70.035 -245.005 70.385 ;
        RECT -240.925 70.035 -240.525 70.385 ;
        RECT -236.445 70.035 -236.045 70.385 ;
        RECT -231.965 70.035 -231.565 70.385 ;
        RECT -227.485 70.035 -227.085 70.385 ;
        RECT -223.005 70.035 -222.605 70.385 ;
        RECT -218.525 70.035 -218.125 70.385 ;
        RECT -214.045 70.035 -213.645 70.385 ;
        RECT -209.565 70.035 -209.165 70.385 ;
        RECT -205.085 70.035 -204.685 70.385 ;
        RECT -200.605 70.035 -200.205 70.385 ;
        RECT -196.125 70.035 -195.725 70.385 ;
        RECT -191.645 70.035 -191.245 70.385 ;
        RECT -186.045 70.035 -185.645 70.385 ;
        RECT -181.565 70.035 -181.165 70.385 ;
        RECT -177.085 70.035 -176.685 70.385 ;
        RECT -172.605 70.035 -172.205 70.385 ;
        RECT -168.125 70.035 -167.725 70.385 ;
        RECT -163.645 70.035 -163.245 70.385 ;
        RECT -159.165 70.035 -158.765 70.385 ;
        RECT -154.685 70.035 -154.285 70.385 ;
        RECT -150.205 70.035 -149.805 70.385 ;
        RECT -145.725 70.035 -145.325 70.385 ;
        RECT -141.245 70.035 -140.845 70.385 ;
        RECT -136.765 70.035 -136.365 70.385 ;
        RECT -132.285 70.035 -131.885 70.385 ;
        RECT -127.805 70.035 -127.405 70.385 ;
        RECT -123.325 70.035 -122.925 70.385 ;
        RECT -118.845 70.035 -118.445 70.385 ;
        RECT -114.365 70.035 -113.965 70.385 ;
        RECT -109.885 70.035 -109.485 70.385 ;
        RECT -105.405 70.035 -105.005 70.385 ;
        RECT -100.925 70.035 -100.525 70.385 ;
        RECT -96.445 70.035 -96.045 70.385 ;
        RECT -91.965 70.035 -91.565 70.385 ;
        RECT -87.485 70.035 -87.085 70.385 ;
        RECT -83.005 70.035 -82.605 70.385 ;
        RECT -78.525 70.035 -78.125 70.385 ;
        RECT -74.045 70.035 -73.645 70.385 ;
        RECT -69.565 70.035 -69.165 70.385 ;
        RECT -65.085 70.035 -64.685 70.385 ;
        RECT -60.605 70.035 -60.205 70.385 ;
        RECT -56.125 70.035 -55.725 70.385 ;
        RECT -51.645 70.035 -51.245 70.385 ;
        RECT -47.165 70.035 -46.765 70.385 ;
        RECT -42.685 70.035 -42.285 70.385 ;
        RECT -38.205 70.035 -37.805 70.385 ;
        RECT -33.725 70.035 -33.325 70.385 ;
        RECT -29.245 70.035 -28.845 70.385 ;
        RECT -24.765 70.035 -24.365 70.385 ;
        RECT -20.285 70.035 -19.885 70.385 ;
        RECT -15.805 70.035 -15.405 70.385 ;
        RECT -11.325 70.035 -10.925 70.385 ;
        RECT -6.845 70.035 -6.445 70.385 ;
        RECT -2.365 70.035 -1.965 70.385 ;
        RECT 2.115 70.035 2.515 70.385 ;
        RECT 6.595 70.035 6.995 70.385 ;
        RECT 11.075 70.035 11.475 70.385 ;
        RECT 15.555 70.035 15.955 70.385 ;
        RECT 20.035 70.035 20.435 70.385 ;
        RECT 24.515 70.035 24.915 70.385 ;
        RECT 28.995 70.035 29.395 70.385 ;
        RECT 33.475 70.035 33.875 70.385 ;
        RECT 37.955 70.035 38.355 70.385 ;
        RECT 42.435 70.035 42.835 70.385 ;
        RECT 46.915 70.035 47.315 70.385 ;
        RECT 51.395 70.035 51.795 70.385 ;
        RECT 55.875 70.035 56.275 70.385 ;
        RECT 60.355 70.035 60.755 70.385 ;
        RECT 64.835 70.035 65.235 70.385 ;
        RECT 69.315 70.035 69.715 70.385 ;
        RECT 73.795 70.035 74.195 70.385 ;
        RECT 78.275 70.035 78.675 70.385 ;
        RECT 82.755 70.035 83.155 70.385 ;
        RECT 87.235 70.035 87.635 70.385 ;
        RECT 91.715 70.035 92.115 70.385 ;
        RECT 96.195 70.035 96.595 70.385 ;
        RECT -475.005 67.525 -474.605 67.875 ;
        RECT -472.765 67.525 -472.365 67.875 ;
        RECT -470.525 67.525 -470.125 67.875 ;
        RECT -468.285 67.525 -467.885 67.875 ;
        RECT -466.045 67.525 -465.645 67.875 ;
        RECT -463.805 67.525 -463.405 67.875 ;
        RECT -461.565 67.525 -461.165 67.875 ;
        RECT -459.325 67.525 -458.925 67.875 ;
        RECT -457.085 67.525 -456.685 67.875 ;
        RECT -454.845 67.525 -454.445 67.875 ;
        RECT -452.605 67.525 -452.205 67.875 ;
        RECT -450.365 67.525 -449.965 67.875 ;
        RECT -448.125 67.525 -447.725 67.875 ;
        RECT -445.885 67.525 -445.485 67.875 ;
        RECT -443.645 67.525 -443.245 67.875 ;
        RECT -441.405 67.525 -441.005 67.875 ;
        RECT -439.165 67.525 -438.765 67.875 ;
        RECT -436.925 67.525 -436.525 67.875 ;
        RECT -434.685 67.525 -434.285 67.875 ;
        RECT -432.445 67.525 -432.045 67.875 ;
        RECT -430.205 67.525 -429.805 67.875 ;
        RECT -427.965 67.525 -427.565 67.875 ;
        RECT -425.725 67.525 -425.325 67.875 ;
        RECT -423.485 67.525 -423.085 67.875 ;
        RECT -421.245 67.525 -420.845 67.875 ;
        RECT -419.005 67.525 -418.605 67.875 ;
        RECT -416.765 67.525 -416.365 67.875 ;
        RECT -414.525 67.525 -414.125 67.875 ;
        RECT -412.285 67.525 -411.885 67.875 ;
        RECT -410.045 67.525 -409.645 67.875 ;
        RECT -407.805 67.525 -407.405 67.875 ;
        RECT -405.565 67.525 -405.165 67.875 ;
        RECT -403.325 67.525 -402.925 67.875 ;
        RECT -401.085 67.525 -400.685 67.875 ;
        RECT -398.845 67.525 -398.445 67.875 ;
        RECT -396.605 67.525 -396.205 67.875 ;
        RECT -394.365 67.525 -393.965 67.875 ;
        RECT -392.125 67.525 -391.725 67.875 ;
        RECT -389.885 67.525 -389.485 67.875 ;
        RECT -387.645 67.525 -387.245 67.875 ;
        RECT -385.405 67.525 -385.005 67.875 ;
        RECT -383.165 67.525 -382.765 67.875 ;
        RECT -380.925 67.525 -380.525 67.875 ;
        RECT -378.685 67.525 -378.285 67.875 ;
        RECT -376.445 67.525 -376.045 67.875 ;
        RECT -374.205 67.525 -373.805 67.875 ;
        RECT -371.965 67.525 -371.565 67.875 ;
        RECT -369.725 67.525 -369.325 67.875 ;
        RECT -367.485 67.525 -367.085 67.875 ;
        RECT -365.245 67.525 -364.845 67.875 ;
        RECT -363.005 67.525 -362.605 67.875 ;
        RECT -360.765 67.525 -360.365 67.875 ;
        RECT -358.525 67.525 -358.125 67.875 ;
        RECT -356.285 67.525 -355.885 67.875 ;
        RECT -354.045 67.525 -353.645 67.875 ;
        RECT -351.805 67.525 -351.405 67.875 ;
        RECT -349.565 67.525 -349.165 67.875 ;
        RECT -347.325 67.525 -346.925 67.875 ;
        RECT -345.085 67.525 -344.685 67.875 ;
        RECT -342.845 67.525 -342.445 67.875 ;
        RECT -340.605 67.525 -340.205 67.875 ;
        RECT -338.365 67.525 -337.965 67.875 ;
        RECT -336.125 67.525 -335.725 67.875 ;
        RECT -333.885 67.525 -333.485 67.875 ;
        RECT -331.645 67.525 -331.245 67.875 ;
        RECT -329.405 67.525 -329.005 67.875 ;
        RECT -327.165 67.525 -326.765 67.875 ;
        RECT -324.925 67.525 -324.525 67.875 ;
        RECT -322.685 67.525 -322.285 67.875 ;
        RECT -320.445 67.525 -320.045 67.875 ;
        RECT -318.205 67.525 -317.805 67.875 ;
        RECT -315.965 67.525 -315.565 67.875 ;
        RECT -313.725 67.525 -313.325 67.875 ;
        RECT -311.485 67.525 -311.085 67.875 ;
        RECT -309.245 67.525 -308.845 67.875 ;
        RECT -307.005 67.525 -306.605 67.875 ;
        RECT -304.765 67.525 -304.365 67.875 ;
        RECT -302.525 67.525 -302.125 67.875 ;
        RECT -300.285 67.525 -299.885 67.875 ;
        RECT -298.045 67.525 -297.645 67.875 ;
        RECT -295.805 67.525 -295.405 67.875 ;
        RECT -293.565 67.525 -293.165 67.875 ;
        RECT -291.325 67.525 -290.925 67.875 ;
        RECT -289.085 67.525 -288.685 67.875 ;
        RECT -286.845 67.525 -286.445 67.875 ;
        RECT -284.605 67.525 -284.205 67.875 ;
        RECT -282.365 67.525 -281.965 67.875 ;
        RECT -280.125 67.525 -279.725 67.875 ;
        RECT -277.885 67.525 -277.485 67.875 ;
        RECT -275.645 67.525 -275.245 67.875 ;
        RECT -273.405 67.525 -273.005 67.875 ;
        RECT -271.165 67.525 -270.765 67.875 ;
        RECT -268.925 67.525 -268.525 67.875 ;
        RECT -266.685 67.525 -266.285 67.875 ;
        RECT -264.445 67.525 -264.045 67.875 ;
        RECT -262.205 67.525 -261.805 67.875 ;
        RECT -259.965 67.525 -259.565 67.875 ;
        RECT -257.725 67.525 -257.325 67.875 ;
        RECT -255.485 67.525 -255.085 67.875 ;
        RECT -253.245 67.525 -252.845 67.875 ;
        RECT -251.005 67.525 -250.605 67.875 ;
        RECT -248.765 67.525 -248.365 67.875 ;
        RECT -246.525 67.525 -246.125 67.875 ;
        RECT -244.285 67.525 -243.885 67.875 ;
        RECT -242.045 67.525 -241.645 67.875 ;
        RECT -239.805 67.525 -239.405 67.875 ;
        RECT -237.565 67.525 -237.165 67.875 ;
        RECT -235.325 67.525 -234.925 67.875 ;
        RECT -233.085 67.525 -232.685 67.875 ;
        RECT -230.845 67.525 -230.445 67.875 ;
        RECT -228.605 67.525 -228.205 67.875 ;
        RECT -226.365 67.525 -225.965 67.875 ;
        RECT -224.125 67.525 -223.725 67.875 ;
        RECT -221.885 67.525 -221.485 67.875 ;
        RECT -219.645 67.525 -219.245 67.875 ;
        RECT -217.405 67.525 -217.005 67.875 ;
        RECT -215.165 67.525 -214.765 67.875 ;
        RECT -212.925 67.525 -212.525 67.875 ;
        RECT -210.685 67.525 -210.285 67.875 ;
        RECT -208.445 67.525 -208.045 67.875 ;
        RECT -206.205 67.525 -205.805 67.875 ;
        RECT -203.965 67.525 -203.565 67.875 ;
        RECT -201.725 67.525 -201.325 67.875 ;
        RECT -199.485 67.525 -199.085 67.875 ;
        RECT -197.245 67.525 -196.845 67.875 ;
        RECT -195.005 67.525 -194.605 67.875 ;
        RECT -192.765 67.525 -192.365 67.875 ;
        RECT -190.525 67.525 -190.125 67.875 ;
        RECT -187.165 67.525 -186.765 67.875 ;
        RECT -184.925 67.525 -184.525 67.875 ;
        RECT -182.685 67.525 -182.285 67.875 ;
        RECT -180.445 67.525 -180.045 67.875 ;
        RECT -178.205 67.525 -177.805 67.875 ;
        RECT -175.965 67.525 -175.565 67.875 ;
        RECT -173.725 67.525 -173.325 67.875 ;
        RECT -171.485 67.525 -171.085 67.875 ;
        RECT -169.245 67.525 -168.845 67.875 ;
        RECT -167.005 67.525 -166.605 67.875 ;
        RECT -164.765 67.525 -164.365 67.875 ;
        RECT -162.525 67.525 -162.125 67.875 ;
        RECT -160.285 67.525 -159.885 67.875 ;
        RECT -158.045 67.525 -157.645 67.875 ;
        RECT -155.805 67.525 -155.405 67.875 ;
        RECT -153.565 67.525 -153.165 67.875 ;
        RECT -151.325 67.525 -150.925 67.875 ;
        RECT -149.085 67.525 -148.685 67.875 ;
        RECT -146.845 67.525 -146.445 67.875 ;
        RECT -144.605 67.525 -144.205 67.875 ;
        RECT -142.365 67.525 -141.965 67.875 ;
        RECT -140.125 67.525 -139.725 67.875 ;
        RECT -137.885 67.525 -137.485 67.875 ;
        RECT -135.645 67.525 -135.245 67.875 ;
        RECT -133.405 67.525 -133.005 67.875 ;
        RECT -131.165 67.525 -130.765 67.875 ;
        RECT -128.925 67.525 -128.525 67.875 ;
        RECT -126.685 67.525 -126.285 67.875 ;
        RECT -124.445 67.525 -124.045 67.875 ;
        RECT -122.205 67.525 -121.805 67.875 ;
        RECT -119.965 67.525 -119.565 67.875 ;
        RECT -117.725 67.525 -117.325 67.875 ;
        RECT -115.485 67.525 -115.085 67.875 ;
        RECT -113.245 67.525 -112.845 67.875 ;
        RECT -111.005 67.525 -110.605 67.875 ;
        RECT -108.765 67.525 -108.365 67.875 ;
        RECT -106.525 67.525 -106.125 67.875 ;
        RECT -104.285 67.525 -103.885 67.875 ;
        RECT -102.045 67.525 -101.645 67.875 ;
        RECT -99.805 67.525 -99.405 67.875 ;
        RECT -97.565 67.525 -97.165 67.875 ;
        RECT -95.325 67.525 -94.925 67.875 ;
        RECT -93.085 67.525 -92.685 67.875 ;
        RECT -90.845 67.525 -90.445 67.875 ;
        RECT -88.605 67.525 -88.205 67.875 ;
        RECT -86.365 67.525 -85.965 67.875 ;
        RECT -84.125 67.525 -83.725 67.875 ;
        RECT -81.885 67.525 -81.485 67.875 ;
        RECT -79.645 67.525 -79.245 67.875 ;
        RECT -77.405 67.525 -77.005 67.875 ;
        RECT -75.165 67.525 -74.765 67.875 ;
        RECT -72.925 67.525 -72.525 67.875 ;
        RECT -70.685 67.525 -70.285 67.875 ;
        RECT -68.445 67.525 -68.045 67.875 ;
        RECT -66.205 67.525 -65.805 67.875 ;
        RECT -63.965 67.525 -63.565 67.875 ;
        RECT -61.725 67.525 -61.325 67.875 ;
        RECT -59.485 67.525 -59.085 67.875 ;
        RECT -57.245 67.525 -56.845 67.875 ;
        RECT -55.005 67.525 -54.605 67.875 ;
        RECT -52.765 67.525 -52.365 67.875 ;
        RECT -50.525 67.525 -50.125 67.875 ;
        RECT -48.285 67.525 -47.885 67.875 ;
        RECT -46.045 67.525 -45.645 67.875 ;
        RECT -43.805 67.525 -43.405 67.875 ;
        RECT -41.565 67.525 -41.165 67.875 ;
        RECT -39.325 67.525 -38.925 67.875 ;
        RECT -37.085 67.525 -36.685 67.875 ;
        RECT -34.845 67.525 -34.445 67.875 ;
        RECT -32.605 67.525 -32.205 67.875 ;
        RECT -30.365 67.525 -29.965 67.875 ;
        RECT -28.125 67.525 -27.725 67.875 ;
        RECT -25.885 67.525 -25.485 67.875 ;
        RECT -23.645 67.525 -23.245 67.875 ;
        RECT -21.405 67.525 -21.005 67.875 ;
        RECT -19.165 67.525 -18.765 67.875 ;
        RECT -16.925 67.525 -16.525 67.875 ;
        RECT -14.685 67.525 -14.285 67.875 ;
        RECT -12.445 67.525 -12.045 67.875 ;
        RECT -10.205 67.525 -9.805 67.875 ;
        RECT -7.965 67.525 -7.565 67.875 ;
        RECT -5.725 67.525 -5.325 67.875 ;
        RECT -3.485 67.525 -3.085 67.875 ;
        RECT -1.245 67.525 -0.845 67.875 ;
        RECT 0.995 67.525 1.395 67.875 ;
        RECT 3.235 67.525 3.635 67.875 ;
        RECT 5.475 67.525 5.875 67.875 ;
        RECT 7.715 67.525 8.115 67.875 ;
        RECT 9.955 67.525 10.355 67.875 ;
        RECT 12.195 67.525 12.595 67.875 ;
        RECT 14.435 67.525 14.835 67.875 ;
        RECT 16.675 67.525 17.075 67.875 ;
        RECT 18.915 67.525 19.315 67.875 ;
        RECT 21.155 67.525 21.555 67.875 ;
        RECT 23.395 67.525 23.795 67.875 ;
        RECT 25.635 67.525 26.035 67.875 ;
        RECT 27.875 67.525 28.275 67.875 ;
        RECT 30.115 67.525 30.515 67.875 ;
        RECT 32.355 67.525 32.755 67.875 ;
        RECT 34.595 67.525 34.995 67.875 ;
        RECT 36.835 67.525 37.235 67.875 ;
        RECT 39.075 67.525 39.475 67.875 ;
        RECT 41.315 67.525 41.715 67.875 ;
        RECT 43.555 67.525 43.955 67.875 ;
        RECT 45.795 67.525 46.195 67.875 ;
        RECT 48.035 67.525 48.435 67.875 ;
        RECT 50.275 67.525 50.675 67.875 ;
        RECT 52.515 67.525 52.915 67.875 ;
        RECT 54.755 67.525 55.155 67.875 ;
        RECT 56.995 67.525 57.395 67.875 ;
        RECT 59.235 67.525 59.635 67.875 ;
        RECT 61.475 67.525 61.875 67.875 ;
        RECT 63.715 67.525 64.115 67.875 ;
        RECT 65.955 67.525 66.355 67.875 ;
        RECT 68.195 67.525 68.595 67.875 ;
        RECT 70.435 67.525 70.835 67.875 ;
        RECT 72.675 67.525 73.075 67.875 ;
        RECT 74.915 67.525 75.315 67.875 ;
        RECT 77.155 67.525 77.555 67.875 ;
        RECT 79.395 67.525 79.795 67.875 ;
        RECT 81.635 67.525 82.035 67.875 ;
        RECT 83.875 67.525 84.275 67.875 ;
        RECT 86.115 67.525 86.515 67.875 ;
        RECT 88.355 67.525 88.755 67.875 ;
        RECT 90.595 67.525 90.995 67.875 ;
        RECT 92.835 67.525 93.235 67.875 ;
        RECT 95.075 67.525 95.475 67.875 ;
        RECT 97.315 67.525 97.715 67.875 ;
        RECT -475.005 67.025 121.925 67.525 ;
        RECT -497.305 66.300 -486.905 66.900 ;
        RECT -475.005 66.675 -474.605 67.025 ;
        RECT -472.765 66.675 -472.365 67.025 ;
        RECT -470.525 66.675 -470.125 67.025 ;
        RECT -468.285 66.675 -467.885 67.025 ;
        RECT -466.045 66.675 -465.645 67.025 ;
        RECT -463.805 66.675 -463.405 67.025 ;
        RECT -461.565 66.675 -461.165 67.025 ;
        RECT -459.325 66.675 -458.925 67.025 ;
        RECT -457.085 66.675 -456.685 67.025 ;
        RECT -454.845 66.675 -454.445 67.025 ;
        RECT -452.605 66.675 -452.205 67.025 ;
        RECT -450.365 66.675 -449.965 67.025 ;
        RECT -448.125 66.675 -447.725 67.025 ;
        RECT -445.885 66.675 -445.485 67.025 ;
        RECT -443.645 66.675 -443.245 67.025 ;
        RECT -441.405 66.675 -441.005 67.025 ;
        RECT -439.165 66.675 -438.765 67.025 ;
        RECT -436.925 66.675 -436.525 67.025 ;
        RECT -434.685 66.675 -434.285 67.025 ;
        RECT -432.445 66.675 -432.045 67.025 ;
        RECT -430.205 66.675 -429.805 67.025 ;
        RECT -427.965 66.675 -427.565 67.025 ;
        RECT -425.725 66.675 -425.325 67.025 ;
        RECT -423.485 66.675 -423.085 67.025 ;
        RECT -421.245 66.675 -420.845 67.025 ;
        RECT -419.005 66.675 -418.605 67.025 ;
        RECT -416.765 66.675 -416.365 67.025 ;
        RECT -414.525 66.675 -414.125 67.025 ;
        RECT -412.285 66.675 -411.885 67.025 ;
        RECT -410.045 66.675 -409.645 67.025 ;
        RECT -407.805 66.675 -407.405 67.025 ;
        RECT -405.565 66.675 -405.165 67.025 ;
        RECT -403.325 66.675 -402.925 67.025 ;
        RECT -401.085 66.675 -400.685 67.025 ;
        RECT -398.845 66.675 -398.445 67.025 ;
        RECT -396.605 66.675 -396.205 67.025 ;
        RECT -394.365 66.675 -393.965 67.025 ;
        RECT -392.125 66.675 -391.725 67.025 ;
        RECT -389.885 66.675 -389.485 67.025 ;
        RECT -387.645 66.675 -387.245 67.025 ;
        RECT -385.405 66.675 -385.005 67.025 ;
        RECT -383.165 66.675 -382.765 67.025 ;
        RECT -380.925 66.675 -380.525 67.025 ;
        RECT -378.685 66.675 -378.285 67.025 ;
        RECT -376.445 66.675 -376.045 67.025 ;
        RECT -374.205 66.675 -373.805 67.025 ;
        RECT -371.965 66.675 -371.565 67.025 ;
        RECT -369.725 66.675 -369.325 67.025 ;
        RECT -367.485 66.675 -367.085 67.025 ;
        RECT -365.245 66.675 -364.845 67.025 ;
        RECT -363.005 66.675 -362.605 67.025 ;
        RECT -360.765 66.675 -360.365 67.025 ;
        RECT -358.525 66.675 -358.125 67.025 ;
        RECT -356.285 66.675 -355.885 67.025 ;
        RECT -354.045 66.675 -353.645 67.025 ;
        RECT -351.805 66.675 -351.405 67.025 ;
        RECT -349.565 66.675 -349.165 67.025 ;
        RECT -347.325 66.675 -346.925 67.025 ;
        RECT -345.085 66.675 -344.685 67.025 ;
        RECT -342.845 66.675 -342.445 67.025 ;
        RECT -340.605 66.675 -340.205 67.025 ;
        RECT -338.365 66.675 -337.965 67.025 ;
        RECT -336.125 66.675 -335.725 67.025 ;
        RECT -333.885 66.675 -333.485 67.025 ;
        RECT -331.645 66.675 -331.245 67.025 ;
        RECT -329.405 66.675 -329.005 67.025 ;
        RECT -327.165 66.675 -326.765 67.025 ;
        RECT -324.925 66.675 -324.525 67.025 ;
        RECT -322.685 66.675 -322.285 67.025 ;
        RECT -320.445 66.675 -320.045 67.025 ;
        RECT -318.205 66.675 -317.805 67.025 ;
        RECT -315.965 66.675 -315.565 67.025 ;
        RECT -313.725 66.675 -313.325 67.025 ;
        RECT -311.485 66.675 -311.085 67.025 ;
        RECT -309.245 66.675 -308.845 67.025 ;
        RECT -307.005 66.675 -306.605 67.025 ;
        RECT -304.765 66.675 -304.365 67.025 ;
        RECT -302.525 66.675 -302.125 67.025 ;
        RECT -300.285 66.675 -299.885 67.025 ;
        RECT -298.045 66.675 -297.645 67.025 ;
        RECT -295.805 66.675 -295.405 67.025 ;
        RECT -293.565 66.675 -293.165 67.025 ;
        RECT -291.325 66.675 -290.925 67.025 ;
        RECT -289.085 66.675 -288.685 67.025 ;
        RECT -286.845 66.675 -286.445 67.025 ;
        RECT -284.605 66.675 -284.205 67.025 ;
        RECT -282.365 66.675 -281.965 67.025 ;
        RECT -280.125 66.675 -279.725 67.025 ;
        RECT -277.885 66.675 -277.485 67.025 ;
        RECT -275.645 66.675 -275.245 67.025 ;
        RECT -273.405 66.675 -273.005 67.025 ;
        RECT -271.165 66.675 -270.765 67.025 ;
        RECT -268.925 66.675 -268.525 67.025 ;
        RECT -266.685 66.675 -266.285 67.025 ;
        RECT -264.445 66.675 -264.045 67.025 ;
        RECT -262.205 66.675 -261.805 67.025 ;
        RECT -259.965 66.675 -259.565 67.025 ;
        RECT -257.725 66.675 -257.325 67.025 ;
        RECT -255.485 66.675 -255.085 67.025 ;
        RECT -253.245 66.675 -252.845 67.025 ;
        RECT -251.005 66.675 -250.605 67.025 ;
        RECT -248.765 66.675 -248.365 67.025 ;
        RECT -246.525 66.675 -246.125 67.025 ;
        RECT -244.285 66.675 -243.885 67.025 ;
        RECT -242.045 66.675 -241.645 67.025 ;
        RECT -239.805 66.675 -239.405 67.025 ;
        RECT -237.565 66.675 -237.165 67.025 ;
        RECT -235.325 66.675 -234.925 67.025 ;
        RECT -233.085 66.675 -232.685 67.025 ;
        RECT -230.845 66.675 -230.445 67.025 ;
        RECT -228.605 66.675 -228.205 67.025 ;
        RECT -226.365 66.675 -225.965 67.025 ;
        RECT -224.125 66.675 -223.725 67.025 ;
        RECT -221.885 66.675 -221.485 67.025 ;
        RECT -219.645 66.675 -219.245 67.025 ;
        RECT -217.405 66.675 -217.005 67.025 ;
        RECT -215.165 66.675 -214.765 67.025 ;
        RECT -212.925 66.675 -212.525 67.025 ;
        RECT -210.685 66.675 -210.285 67.025 ;
        RECT -208.445 66.675 -208.045 67.025 ;
        RECT -206.205 66.675 -205.805 67.025 ;
        RECT -203.965 66.675 -203.565 67.025 ;
        RECT -201.725 66.675 -201.325 67.025 ;
        RECT -199.485 66.675 -199.085 67.025 ;
        RECT -197.245 66.675 -196.845 67.025 ;
        RECT -195.005 66.675 -194.605 67.025 ;
        RECT -192.765 66.675 -192.365 67.025 ;
        RECT -190.525 66.675 -190.125 67.025 ;
        RECT -187.165 66.675 -186.765 67.025 ;
        RECT -184.925 66.675 -184.525 67.025 ;
        RECT -182.685 66.675 -182.285 67.025 ;
        RECT -180.445 66.675 -180.045 67.025 ;
        RECT -178.205 66.675 -177.805 67.025 ;
        RECT -175.965 66.675 -175.565 67.025 ;
        RECT -173.725 66.675 -173.325 67.025 ;
        RECT -171.485 66.675 -171.085 67.025 ;
        RECT -169.245 66.675 -168.845 67.025 ;
        RECT -167.005 66.675 -166.605 67.025 ;
        RECT -164.765 66.675 -164.365 67.025 ;
        RECT -162.525 66.675 -162.125 67.025 ;
        RECT -160.285 66.675 -159.885 67.025 ;
        RECT -158.045 66.675 -157.645 67.025 ;
        RECT -155.805 66.675 -155.405 67.025 ;
        RECT -153.565 66.675 -153.165 67.025 ;
        RECT -151.325 66.675 -150.925 67.025 ;
        RECT -149.085 66.675 -148.685 67.025 ;
        RECT -146.845 66.675 -146.445 67.025 ;
        RECT -144.605 66.675 -144.205 67.025 ;
        RECT -142.365 66.675 -141.965 67.025 ;
        RECT -140.125 66.675 -139.725 67.025 ;
        RECT -137.885 66.675 -137.485 67.025 ;
        RECT -135.645 66.675 -135.245 67.025 ;
        RECT -133.405 66.675 -133.005 67.025 ;
        RECT -131.165 66.675 -130.765 67.025 ;
        RECT -128.925 66.675 -128.525 67.025 ;
        RECT -126.685 66.675 -126.285 67.025 ;
        RECT -124.445 66.675 -124.045 67.025 ;
        RECT -122.205 66.675 -121.805 67.025 ;
        RECT -119.965 66.675 -119.565 67.025 ;
        RECT -117.725 66.675 -117.325 67.025 ;
        RECT -115.485 66.675 -115.085 67.025 ;
        RECT -113.245 66.675 -112.845 67.025 ;
        RECT -111.005 66.675 -110.605 67.025 ;
        RECT -108.765 66.675 -108.365 67.025 ;
        RECT -106.525 66.675 -106.125 67.025 ;
        RECT -104.285 66.675 -103.885 67.025 ;
        RECT -102.045 66.675 -101.645 67.025 ;
        RECT -99.805 66.675 -99.405 67.025 ;
        RECT -97.565 66.675 -97.165 67.025 ;
        RECT -95.325 66.675 -94.925 67.025 ;
        RECT -93.085 66.675 -92.685 67.025 ;
        RECT -90.845 66.675 -90.445 67.025 ;
        RECT -88.605 66.675 -88.205 67.025 ;
        RECT -86.365 66.675 -85.965 67.025 ;
        RECT -84.125 66.675 -83.725 67.025 ;
        RECT -81.885 66.675 -81.485 67.025 ;
        RECT -79.645 66.675 -79.245 67.025 ;
        RECT -77.405 66.675 -77.005 67.025 ;
        RECT -75.165 66.675 -74.765 67.025 ;
        RECT -72.925 66.675 -72.525 67.025 ;
        RECT -70.685 66.675 -70.285 67.025 ;
        RECT -68.445 66.675 -68.045 67.025 ;
        RECT -66.205 66.675 -65.805 67.025 ;
        RECT -63.965 66.675 -63.565 67.025 ;
        RECT -61.725 66.675 -61.325 67.025 ;
        RECT -59.485 66.675 -59.085 67.025 ;
        RECT -57.245 66.675 -56.845 67.025 ;
        RECT -55.005 66.675 -54.605 67.025 ;
        RECT -52.765 66.675 -52.365 67.025 ;
        RECT -50.525 66.675 -50.125 67.025 ;
        RECT -48.285 66.675 -47.885 67.025 ;
        RECT -46.045 66.675 -45.645 67.025 ;
        RECT -43.805 66.675 -43.405 67.025 ;
        RECT -41.565 66.675 -41.165 67.025 ;
        RECT -39.325 66.675 -38.925 67.025 ;
        RECT -37.085 66.675 -36.685 67.025 ;
        RECT -34.845 66.675 -34.445 67.025 ;
        RECT -32.605 66.675 -32.205 67.025 ;
        RECT -30.365 66.675 -29.965 67.025 ;
        RECT -28.125 66.675 -27.725 67.025 ;
        RECT -25.885 66.675 -25.485 67.025 ;
        RECT -23.645 66.675 -23.245 67.025 ;
        RECT -21.405 66.675 -21.005 67.025 ;
        RECT -19.165 66.675 -18.765 67.025 ;
        RECT -16.925 66.675 -16.525 67.025 ;
        RECT -14.685 66.675 -14.285 67.025 ;
        RECT -12.445 66.675 -12.045 67.025 ;
        RECT -10.205 66.675 -9.805 67.025 ;
        RECT -7.965 66.675 -7.565 67.025 ;
        RECT -5.725 66.675 -5.325 67.025 ;
        RECT -3.485 66.675 -3.085 67.025 ;
        RECT -1.245 66.675 -0.845 67.025 ;
        RECT 0.995 66.675 1.395 67.025 ;
        RECT 3.235 66.675 3.635 67.025 ;
        RECT 5.475 66.675 5.875 67.025 ;
        RECT 7.715 66.675 8.115 67.025 ;
        RECT 9.955 66.675 10.355 67.025 ;
        RECT 12.195 66.675 12.595 67.025 ;
        RECT 14.435 66.675 14.835 67.025 ;
        RECT 16.675 66.675 17.075 67.025 ;
        RECT 18.915 66.675 19.315 67.025 ;
        RECT 21.155 66.675 21.555 67.025 ;
        RECT 23.395 66.675 23.795 67.025 ;
        RECT 25.635 66.675 26.035 67.025 ;
        RECT 27.875 66.675 28.275 67.025 ;
        RECT 30.115 66.675 30.515 67.025 ;
        RECT 32.355 66.675 32.755 67.025 ;
        RECT 34.595 66.675 34.995 67.025 ;
        RECT 36.835 66.675 37.235 67.025 ;
        RECT 39.075 66.675 39.475 67.025 ;
        RECT 41.315 66.675 41.715 67.025 ;
        RECT 43.555 66.675 43.955 67.025 ;
        RECT 45.795 66.675 46.195 67.025 ;
        RECT 48.035 66.675 48.435 67.025 ;
        RECT 50.275 66.675 50.675 67.025 ;
        RECT 52.515 66.675 52.915 67.025 ;
        RECT 54.755 66.675 55.155 67.025 ;
        RECT 56.995 66.675 57.395 67.025 ;
        RECT 59.235 66.675 59.635 67.025 ;
        RECT 61.475 66.675 61.875 67.025 ;
        RECT 63.715 66.675 64.115 67.025 ;
        RECT 65.955 66.675 66.355 67.025 ;
        RECT 68.195 66.675 68.595 67.025 ;
        RECT 70.435 66.675 70.835 67.025 ;
        RECT 72.675 66.675 73.075 67.025 ;
        RECT 74.915 66.675 75.315 67.025 ;
        RECT 77.155 66.675 77.555 67.025 ;
        RECT 79.395 66.675 79.795 67.025 ;
        RECT 81.635 66.675 82.035 67.025 ;
        RECT 83.875 66.675 84.275 67.025 ;
        RECT 86.115 66.675 86.515 67.025 ;
        RECT 88.355 66.675 88.755 67.025 ;
        RECT 90.595 66.675 90.995 67.025 ;
        RECT 92.835 66.675 93.235 67.025 ;
        RECT 95.075 66.675 95.475 67.025 ;
        RECT 97.315 66.675 97.715 67.025 ;
        RECT -497.305 58.300 -495.505 66.300 ;
        RECT -487.505 58.300 -486.905 66.300 ;
        RECT -497.305 57.700 -486.905 58.300 ;
        RECT 117.705 63.665 121.925 64.165 ;
        RECT -497.305 54.300 -486.905 54.900 ;
        RECT -497.305 46.300 -495.505 54.300 ;
        RECT -487.505 46.300 -486.905 54.300 ;
        RECT -497.305 45.700 -486.905 46.300 ;
        RECT -475.005 44.665 -474.605 45.015 ;
        RECT -472.765 44.665 -472.365 45.015 ;
        RECT -470.525 44.665 -470.125 45.015 ;
        RECT -468.285 44.665 -467.885 45.015 ;
        RECT -466.045 44.665 -465.645 45.015 ;
        RECT -463.805 44.665 -463.405 45.015 ;
        RECT -461.565 44.665 -461.165 45.015 ;
        RECT -459.325 44.665 -458.925 45.015 ;
        RECT -457.085 44.665 -456.685 45.015 ;
        RECT -454.845 44.665 -454.445 45.015 ;
        RECT -452.605 44.665 -452.205 45.015 ;
        RECT -450.365 44.665 -449.965 45.015 ;
        RECT -448.125 44.665 -447.725 45.015 ;
        RECT -445.885 44.665 -445.485 45.015 ;
        RECT -443.645 44.665 -443.245 45.015 ;
        RECT -441.405 44.665 -441.005 45.015 ;
        RECT -439.165 44.665 -438.765 45.015 ;
        RECT -436.925 44.665 -436.525 45.015 ;
        RECT -434.685 44.665 -434.285 45.015 ;
        RECT -432.445 44.665 -432.045 45.015 ;
        RECT -430.205 44.665 -429.805 45.015 ;
        RECT -427.965 44.665 -427.565 45.015 ;
        RECT -425.725 44.665 -425.325 45.015 ;
        RECT -423.485 44.665 -423.085 45.015 ;
        RECT -421.245 44.665 -420.845 45.015 ;
        RECT -419.005 44.665 -418.605 45.015 ;
        RECT -416.765 44.665 -416.365 45.015 ;
        RECT -414.525 44.665 -414.125 45.015 ;
        RECT -412.285 44.665 -411.885 45.015 ;
        RECT -410.045 44.665 -409.645 45.015 ;
        RECT -407.805 44.665 -407.405 45.015 ;
        RECT -405.565 44.665 -405.165 45.015 ;
        RECT -403.325 44.665 -402.925 45.015 ;
        RECT -401.085 44.665 -400.685 45.015 ;
        RECT -398.845 44.665 -398.445 45.015 ;
        RECT -396.605 44.665 -396.205 45.015 ;
        RECT -394.365 44.665 -393.965 45.015 ;
        RECT -392.125 44.665 -391.725 45.015 ;
        RECT -389.885 44.665 -389.485 45.015 ;
        RECT -387.645 44.665 -387.245 45.015 ;
        RECT -385.405 44.665 -385.005 45.015 ;
        RECT -383.165 44.665 -382.765 45.015 ;
        RECT -380.925 44.665 -380.525 45.015 ;
        RECT -378.685 44.665 -378.285 45.015 ;
        RECT -376.445 44.665 -376.045 45.015 ;
        RECT -374.205 44.665 -373.805 45.015 ;
        RECT -371.965 44.665 -371.565 45.015 ;
        RECT -369.725 44.665 -369.325 45.015 ;
        RECT -367.485 44.665 -367.085 45.015 ;
        RECT -365.245 44.665 -364.845 45.015 ;
        RECT -363.005 44.665 -362.605 45.015 ;
        RECT -360.765 44.665 -360.365 45.015 ;
        RECT -358.525 44.665 -358.125 45.015 ;
        RECT -356.285 44.665 -355.885 45.015 ;
        RECT -354.045 44.665 -353.645 45.015 ;
        RECT -351.805 44.665 -351.405 45.015 ;
        RECT -349.565 44.665 -349.165 45.015 ;
        RECT -347.325 44.665 -346.925 45.015 ;
        RECT -345.085 44.665 -344.685 45.015 ;
        RECT -342.845 44.665 -342.445 45.015 ;
        RECT -340.605 44.665 -340.205 45.015 ;
        RECT -338.365 44.665 -337.965 45.015 ;
        RECT -336.125 44.665 -335.725 45.015 ;
        RECT -333.885 44.665 -333.485 45.015 ;
        RECT -331.645 44.665 -331.245 45.015 ;
        RECT -329.405 44.665 -329.005 45.015 ;
        RECT -327.165 44.665 -326.765 45.015 ;
        RECT -324.925 44.665 -324.525 45.015 ;
        RECT -322.685 44.665 -322.285 45.015 ;
        RECT -320.445 44.665 -320.045 45.015 ;
        RECT -318.205 44.665 -317.805 45.015 ;
        RECT -315.965 44.665 -315.565 45.015 ;
        RECT -313.725 44.665 -313.325 45.015 ;
        RECT -311.485 44.665 -311.085 45.015 ;
        RECT -309.245 44.665 -308.845 45.015 ;
        RECT -307.005 44.665 -306.605 45.015 ;
        RECT -304.765 44.665 -304.365 45.015 ;
        RECT -302.525 44.665 -302.125 45.015 ;
        RECT -300.285 44.665 -299.885 45.015 ;
        RECT -298.045 44.665 -297.645 45.015 ;
        RECT -295.805 44.665 -295.405 45.015 ;
        RECT -293.565 44.665 -293.165 45.015 ;
        RECT -291.325 44.665 -290.925 45.015 ;
        RECT -289.085 44.665 -288.685 45.015 ;
        RECT -286.845 44.665 -286.445 45.015 ;
        RECT -284.605 44.665 -284.205 45.015 ;
        RECT -282.365 44.665 -281.965 45.015 ;
        RECT -280.125 44.665 -279.725 45.015 ;
        RECT -277.885 44.665 -277.485 45.015 ;
        RECT -275.645 44.665 -275.245 45.015 ;
        RECT -273.405 44.665 -273.005 45.015 ;
        RECT -271.165 44.665 -270.765 45.015 ;
        RECT -268.925 44.665 -268.525 45.015 ;
        RECT -266.685 44.665 -266.285 45.015 ;
        RECT -264.445 44.665 -264.045 45.015 ;
        RECT -262.205 44.665 -261.805 45.015 ;
        RECT -259.965 44.665 -259.565 45.015 ;
        RECT -257.725 44.665 -257.325 45.015 ;
        RECT -255.485 44.665 -255.085 45.015 ;
        RECT -253.245 44.665 -252.845 45.015 ;
        RECT -251.005 44.665 -250.605 45.015 ;
        RECT -248.765 44.665 -248.365 45.015 ;
        RECT -246.525 44.665 -246.125 45.015 ;
        RECT -244.285 44.665 -243.885 45.015 ;
        RECT -242.045 44.665 -241.645 45.015 ;
        RECT -239.805 44.665 -239.405 45.015 ;
        RECT -237.565 44.665 -237.165 45.015 ;
        RECT -235.325 44.665 -234.925 45.015 ;
        RECT -233.085 44.665 -232.685 45.015 ;
        RECT -230.845 44.665 -230.445 45.015 ;
        RECT -228.605 44.665 -228.205 45.015 ;
        RECT -226.365 44.665 -225.965 45.015 ;
        RECT -224.125 44.665 -223.725 45.015 ;
        RECT -221.885 44.665 -221.485 45.015 ;
        RECT -219.645 44.665 -219.245 45.015 ;
        RECT -217.405 44.665 -217.005 45.015 ;
        RECT -215.165 44.665 -214.765 45.015 ;
        RECT -212.925 44.665 -212.525 45.015 ;
        RECT -210.685 44.665 -210.285 45.015 ;
        RECT -208.445 44.665 -208.045 45.015 ;
        RECT -206.205 44.665 -205.805 45.015 ;
        RECT -203.965 44.665 -203.565 45.015 ;
        RECT -201.725 44.665 -201.325 45.015 ;
        RECT -199.485 44.665 -199.085 45.015 ;
        RECT -197.245 44.665 -196.845 45.015 ;
        RECT -195.005 44.665 -194.605 45.015 ;
        RECT -192.765 44.665 -192.365 45.015 ;
        RECT -190.525 44.665 -190.125 45.015 ;
        RECT -187.165 44.665 -186.765 45.015 ;
        RECT -184.925 44.665 -184.525 45.015 ;
        RECT -182.685 44.665 -182.285 45.015 ;
        RECT -180.445 44.665 -180.045 45.015 ;
        RECT -178.205 44.665 -177.805 45.015 ;
        RECT -175.965 44.665 -175.565 45.015 ;
        RECT -173.725 44.665 -173.325 45.015 ;
        RECT -171.485 44.665 -171.085 45.015 ;
        RECT -169.245 44.665 -168.845 45.015 ;
        RECT -167.005 44.665 -166.605 45.015 ;
        RECT -164.765 44.665 -164.365 45.015 ;
        RECT -162.525 44.665 -162.125 45.015 ;
        RECT -160.285 44.665 -159.885 45.015 ;
        RECT -158.045 44.665 -157.645 45.015 ;
        RECT -155.805 44.665 -155.405 45.015 ;
        RECT -153.565 44.665 -153.165 45.015 ;
        RECT -151.325 44.665 -150.925 45.015 ;
        RECT -149.085 44.665 -148.685 45.015 ;
        RECT -146.845 44.665 -146.445 45.015 ;
        RECT -144.605 44.665 -144.205 45.015 ;
        RECT -142.365 44.665 -141.965 45.015 ;
        RECT -140.125 44.665 -139.725 45.015 ;
        RECT -137.885 44.665 -137.485 45.015 ;
        RECT -135.645 44.665 -135.245 45.015 ;
        RECT -133.405 44.665 -133.005 45.015 ;
        RECT -131.165 44.665 -130.765 45.015 ;
        RECT -128.925 44.665 -128.525 45.015 ;
        RECT -126.685 44.665 -126.285 45.015 ;
        RECT -124.445 44.665 -124.045 45.015 ;
        RECT -122.205 44.665 -121.805 45.015 ;
        RECT -119.965 44.665 -119.565 45.015 ;
        RECT -117.725 44.665 -117.325 45.015 ;
        RECT -115.485 44.665 -115.085 45.015 ;
        RECT -113.245 44.665 -112.845 45.015 ;
        RECT -111.005 44.665 -110.605 45.015 ;
        RECT -108.765 44.665 -108.365 45.015 ;
        RECT -106.525 44.665 -106.125 45.015 ;
        RECT -104.285 44.665 -103.885 45.015 ;
        RECT -102.045 44.665 -101.645 45.015 ;
        RECT -99.805 44.665 -99.405 45.015 ;
        RECT -97.565 44.665 -97.165 45.015 ;
        RECT -95.325 44.665 -94.925 45.015 ;
        RECT -93.085 44.665 -92.685 45.015 ;
        RECT -90.845 44.665 -90.445 45.015 ;
        RECT -88.605 44.665 -88.205 45.015 ;
        RECT -86.365 44.665 -85.965 45.015 ;
        RECT -84.125 44.665 -83.725 45.015 ;
        RECT -81.885 44.665 -81.485 45.015 ;
        RECT -79.645 44.665 -79.245 45.015 ;
        RECT -77.405 44.665 -77.005 45.015 ;
        RECT -75.165 44.665 -74.765 45.015 ;
        RECT -72.925 44.665 -72.525 45.015 ;
        RECT -70.685 44.665 -70.285 45.015 ;
        RECT -68.445 44.665 -68.045 45.015 ;
        RECT -66.205 44.665 -65.805 45.015 ;
        RECT -63.965 44.665 -63.565 45.015 ;
        RECT -61.725 44.665 -61.325 45.015 ;
        RECT -59.485 44.665 -59.085 45.015 ;
        RECT -57.245 44.665 -56.845 45.015 ;
        RECT -55.005 44.665 -54.605 45.015 ;
        RECT -52.765 44.665 -52.365 45.015 ;
        RECT -50.525 44.665 -50.125 45.015 ;
        RECT -48.285 44.665 -47.885 45.015 ;
        RECT -46.045 44.665 -45.645 45.015 ;
        RECT -43.805 44.665 -43.405 45.015 ;
        RECT -41.565 44.665 -41.165 45.015 ;
        RECT -39.325 44.665 -38.925 45.015 ;
        RECT -37.085 44.665 -36.685 45.015 ;
        RECT -34.845 44.665 -34.445 45.015 ;
        RECT -32.605 44.665 -32.205 45.015 ;
        RECT -30.365 44.665 -29.965 45.015 ;
        RECT -28.125 44.665 -27.725 45.015 ;
        RECT -25.885 44.665 -25.485 45.015 ;
        RECT -23.645 44.665 -23.245 45.015 ;
        RECT -21.405 44.665 -21.005 45.015 ;
        RECT -19.165 44.665 -18.765 45.015 ;
        RECT -16.925 44.665 -16.525 45.015 ;
        RECT -14.685 44.665 -14.285 45.015 ;
        RECT -12.445 44.665 -12.045 45.015 ;
        RECT -10.205 44.665 -9.805 45.015 ;
        RECT -7.965 44.665 -7.565 45.015 ;
        RECT -5.725 44.665 -5.325 45.015 ;
        RECT -3.485 44.665 -3.085 45.015 ;
        RECT -1.245 44.665 -0.845 45.015 ;
        RECT 0.995 44.665 1.395 45.015 ;
        RECT 3.235 44.665 3.635 45.015 ;
        RECT 5.475 44.665 5.875 45.015 ;
        RECT 7.715 44.665 8.115 45.015 ;
        RECT 9.955 44.665 10.355 45.015 ;
        RECT 12.195 44.665 12.595 45.015 ;
        RECT 14.435 44.665 14.835 45.015 ;
        RECT 16.675 44.665 17.075 45.015 ;
        RECT 18.915 44.665 19.315 45.015 ;
        RECT 21.155 44.665 21.555 45.015 ;
        RECT 23.395 44.665 23.795 45.015 ;
        RECT 25.635 44.665 26.035 45.015 ;
        RECT 27.875 44.665 28.275 45.015 ;
        RECT 30.115 44.665 30.515 45.015 ;
        RECT 32.355 44.665 32.755 45.015 ;
        RECT 34.595 44.665 34.995 45.015 ;
        RECT 36.835 44.665 37.235 45.015 ;
        RECT 39.075 44.665 39.475 45.015 ;
        RECT 41.315 44.665 41.715 45.015 ;
        RECT 43.555 44.665 43.955 45.015 ;
        RECT 45.795 44.665 46.195 45.015 ;
        RECT 48.035 44.665 48.435 45.015 ;
        RECT 50.275 44.665 50.675 45.015 ;
        RECT 52.515 44.665 52.915 45.015 ;
        RECT 54.755 44.665 55.155 45.015 ;
        RECT 56.995 44.665 57.395 45.015 ;
        RECT 59.235 44.665 59.635 45.015 ;
        RECT 61.475 44.665 61.875 45.015 ;
        RECT 63.715 44.665 64.115 45.015 ;
        RECT 65.955 44.665 66.355 45.015 ;
        RECT 68.195 44.665 68.595 45.015 ;
        RECT 70.435 44.665 70.835 45.015 ;
        RECT 72.675 44.665 73.075 45.015 ;
        RECT 74.915 44.665 75.315 45.015 ;
        RECT 77.155 44.665 77.555 45.015 ;
        RECT 79.395 44.665 79.795 45.015 ;
        RECT 81.635 44.665 82.035 45.015 ;
        RECT 83.875 44.665 84.275 45.015 ;
        RECT 86.115 44.665 86.515 45.015 ;
        RECT 88.355 44.665 88.755 45.015 ;
        RECT 90.595 44.665 90.995 45.015 ;
        RECT 92.835 44.665 93.235 45.015 ;
        RECT 95.075 44.665 95.475 45.015 ;
        RECT 97.315 44.665 97.715 45.015 ;
        RECT -475.005 44.615 101.955 44.665 ;
        RECT -475.005 44.215 102.355 44.615 ;
        RECT -475.005 44.165 101.955 44.215 ;
        RECT -475.005 43.815 -474.605 44.165 ;
        RECT -472.765 43.815 -472.365 44.165 ;
        RECT -470.525 43.815 -470.125 44.165 ;
        RECT -468.285 43.815 -467.885 44.165 ;
        RECT -466.045 43.815 -465.645 44.165 ;
        RECT -463.805 43.815 -463.405 44.165 ;
        RECT -461.565 43.815 -461.165 44.165 ;
        RECT -459.325 43.815 -458.925 44.165 ;
        RECT -457.085 43.815 -456.685 44.165 ;
        RECT -454.845 43.815 -454.445 44.165 ;
        RECT -452.605 43.815 -452.205 44.165 ;
        RECT -450.365 43.815 -449.965 44.165 ;
        RECT -448.125 43.815 -447.725 44.165 ;
        RECT -445.885 43.815 -445.485 44.165 ;
        RECT -443.645 43.815 -443.245 44.165 ;
        RECT -441.405 43.815 -441.005 44.165 ;
        RECT -439.165 43.815 -438.765 44.165 ;
        RECT -436.925 43.815 -436.525 44.165 ;
        RECT -434.685 43.815 -434.285 44.165 ;
        RECT -432.445 43.815 -432.045 44.165 ;
        RECT -430.205 43.815 -429.805 44.165 ;
        RECT -427.965 43.815 -427.565 44.165 ;
        RECT -425.725 43.815 -425.325 44.165 ;
        RECT -423.485 43.815 -423.085 44.165 ;
        RECT -421.245 43.815 -420.845 44.165 ;
        RECT -419.005 43.815 -418.605 44.165 ;
        RECT -416.765 43.815 -416.365 44.165 ;
        RECT -414.525 43.815 -414.125 44.165 ;
        RECT -412.285 43.815 -411.885 44.165 ;
        RECT -410.045 43.815 -409.645 44.165 ;
        RECT -407.805 43.815 -407.405 44.165 ;
        RECT -405.565 43.815 -405.165 44.165 ;
        RECT -403.325 43.815 -402.925 44.165 ;
        RECT -401.085 43.815 -400.685 44.165 ;
        RECT -398.845 43.815 -398.445 44.165 ;
        RECT -396.605 43.815 -396.205 44.165 ;
        RECT -394.365 43.815 -393.965 44.165 ;
        RECT -392.125 43.815 -391.725 44.165 ;
        RECT -389.885 43.815 -389.485 44.165 ;
        RECT -387.645 43.815 -387.245 44.165 ;
        RECT -385.405 43.815 -385.005 44.165 ;
        RECT -383.165 43.815 -382.765 44.165 ;
        RECT -380.925 43.815 -380.525 44.165 ;
        RECT -378.685 43.815 -378.285 44.165 ;
        RECT -376.445 43.815 -376.045 44.165 ;
        RECT -374.205 43.815 -373.805 44.165 ;
        RECT -371.965 43.815 -371.565 44.165 ;
        RECT -369.725 43.815 -369.325 44.165 ;
        RECT -367.485 43.815 -367.085 44.165 ;
        RECT -365.245 43.815 -364.845 44.165 ;
        RECT -363.005 43.815 -362.605 44.165 ;
        RECT -360.765 43.815 -360.365 44.165 ;
        RECT -358.525 43.815 -358.125 44.165 ;
        RECT -356.285 43.815 -355.885 44.165 ;
        RECT -354.045 43.815 -353.645 44.165 ;
        RECT -351.805 43.815 -351.405 44.165 ;
        RECT -349.565 43.815 -349.165 44.165 ;
        RECT -347.325 43.815 -346.925 44.165 ;
        RECT -345.085 43.815 -344.685 44.165 ;
        RECT -342.845 43.815 -342.445 44.165 ;
        RECT -340.605 43.815 -340.205 44.165 ;
        RECT -338.365 43.815 -337.965 44.165 ;
        RECT -336.125 43.815 -335.725 44.165 ;
        RECT -333.885 43.815 -333.485 44.165 ;
        RECT -331.645 43.815 -331.245 44.165 ;
        RECT -329.405 43.815 -329.005 44.165 ;
        RECT -327.165 43.815 -326.765 44.165 ;
        RECT -324.925 43.815 -324.525 44.165 ;
        RECT -322.685 43.815 -322.285 44.165 ;
        RECT -320.445 43.815 -320.045 44.165 ;
        RECT -318.205 43.815 -317.805 44.165 ;
        RECT -315.965 43.815 -315.565 44.165 ;
        RECT -313.725 43.815 -313.325 44.165 ;
        RECT -311.485 43.815 -311.085 44.165 ;
        RECT -309.245 43.815 -308.845 44.165 ;
        RECT -307.005 43.815 -306.605 44.165 ;
        RECT -304.765 43.815 -304.365 44.165 ;
        RECT -302.525 43.815 -302.125 44.165 ;
        RECT -300.285 43.815 -299.885 44.165 ;
        RECT -298.045 43.815 -297.645 44.165 ;
        RECT -295.805 43.815 -295.405 44.165 ;
        RECT -293.565 43.815 -293.165 44.165 ;
        RECT -291.325 43.815 -290.925 44.165 ;
        RECT -289.085 43.815 -288.685 44.165 ;
        RECT -286.845 43.815 -286.445 44.165 ;
        RECT -284.605 43.815 -284.205 44.165 ;
        RECT -282.365 43.815 -281.965 44.165 ;
        RECT -280.125 43.815 -279.725 44.165 ;
        RECT -277.885 43.815 -277.485 44.165 ;
        RECT -275.645 43.815 -275.245 44.165 ;
        RECT -273.405 43.815 -273.005 44.165 ;
        RECT -271.165 43.815 -270.765 44.165 ;
        RECT -268.925 43.815 -268.525 44.165 ;
        RECT -266.685 43.815 -266.285 44.165 ;
        RECT -264.445 43.815 -264.045 44.165 ;
        RECT -262.205 43.815 -261.805 44.165 ;
        RECT -259.965 43.815 -259.565 44.165 ;
        RECT -257.725 43.815 -257.325 44.165 ;
        RECT -255.485 43.815 -255.085 44.165 ;
        RECT -253.245 43.815 -252.845 44.165 ;
        RECT -251.005 43.815 -250.605 44.165 ;
        RECT -248.765 43.815 -248.365 44.165 ;
        RECT -246.525 43.815 -246.125 44.165 ;
        RECT -244.285 43.815 -243.885 44.165 ;
        RECT -242.045 43.815 -241.645 44.165 ;
        RECT -239.805 43.815 -239.405 44.165 ;
        RECT -237.565 43.815 -237.165 44.165 ;
        RECT -235.325 43.815 -234.925 44.165 ;
        RECT -233.085 43.815 -232.685 44.165 ;
        RECT -230.845 43.815 -230.445 44.165 ;
        RECT -228.605 43.815 -228.205 44.165 ;
        RECT -226.365 43.815 -225.965 44.165 ;
        RECT -224.125 43.815 -223.725 44.165 ;
        RECT -221.885 43.815 -221.485 44.165 ;
        RECT -219.645 43.815 -219.245 44.165 ;
        RECT -217.405 43.815 -217.005 44.165 ;
        RECT -215.165 43.815 -214.765 44.165 ;
        RECT -212.925 43.815 -212.525 44.165 ;
        RECT -210.685 43.815 -210.285 44.165 ;
        RECT -208.445 43.815 -208.045 44.165 ;
        RECT -206.205 43.815 -205.805 44.165 ;
        RECT -203.965 43.815 -203.565 44.165 ;
        RECT -201.725 43.815 -201.325 44.165 ;
        RECT -199.485 43.815 -199.085 44.165 ;
        RECT -197.245 43.815 -196.845 44.165 ;
        RECT -195.005 43.815 -194.605 44.165 ;
        RECT -192.765 43.815 -192.365 44.165 ;
        RECT -190.525 43.815 -190.125 44.165 ;
        RECT -187.165 43.815 -186.765 44.165 ;
        RECT -184.925 43.815 -184.525 44.165 ;
        RECT -182.685 43.815 -182.285 44.165 ;
        RECT -180.445 43.815 -180.045 44.165 ;
        RECT -178.205 43.815 -177.805 44.165 ;
        RECT -175.965 43.815 -175.565 44.165 ;
        RECT -173.725 43.815 -173.325 44.165 ;
        RECT -171.485 43.815 -171.085 44.165 ;
        RECT -169.245 43.815 -168.845 44.165 ;
        RECT -167.005 43.815 -166.605 44.165 ;
        RECT -164.765 43.815 -164.365 44.165 ;
        RECT -162.525 43.815 -162.125 44.165 ;
        RECT -160.285 43.815 -159.885 44.165 ;
        RECT -158.045 43.815 -157.645 44.165 ;
        RECT -155.805 43.815 -155.405 44.165 ;
        RECT -153.565 43.815 -153.165 44.165 ;
        RECT -151.325 43.815 -150.925 44.165 ;
        RECT -149.085 43.815 -148.685 44.165 ;
        RECT -146.845 43.815 -146.445 44.165 ;
        RECT -144.605 43.815 -144.205 44.165 ;
        RECT -142.365 43.815 -141.965 44.165 ;
        RECT -140.125 43.815 -139.725 44.165 ;
        RECT -137.885 43.815 -137.485 44.165 ;
        RECT -135.645 43.815 -135.245 44.165 ;
        RECT -133.405 43.815 -133.005 44.165 ;
        RECT -131.165 43.815 -130.765 44.165 ;
        RECT -128.925 43.815 -128.525 44.165 ;
        RECT -126.685 43.815 -126.285 44.165 ;
        RECT -124.445 43.815 -124.045 44.165 ;
        RECT -122.205 43.815 -121.805 44.165 ;
        RECT -119.965 43.815 -119.565 44.165 ;
        RECT -117.725 43.815 -117.325 44.165 ;
        RECT -115.485 43.815 -115.085 44.165 ;
        RECT -113.245 43.815 -112.845 44.165 ;
        RECT -111.005 43.815 -110.605 44.165 ;
        RECT -108.765 43.815 -108.365 44.165 ;
        RECT -106.525 43.815 -106.125 44.165 ;
        RECT -104.285 43.815 -103.885 44.165 ;
        RECT -102.045 43.815 -101.645 44.165 ;
        RECT -99.805 43.815 -99.405 44.165 ;
        RECT -97.565 43.815 -97.165 44.165 ;
        RECT -95.325 43.815 -94.925 44.165 ;
        RECT -93.085 43.815 -92.685 44.165 ;
        RECT -90.845 43.815 -90.445 44.165 ;
        RECT -88.605 43.815 -88.205 44.165 ;
        RECT -86.365 43.815 -85.965 44.165 ;
        RECT -84.125 43.815 -83.725 44.165 ;
        RECT -81.885 43.815 -81.485 44.165 ;
        RECT -79.645 43.815 -79.245 44.165 ;
        RECT -77.405 43.815 -77.005 44.165 ;
        RECT -75.165 43.815 -74.765 44.165 ;
        RECT -72.925 43.815 -72.525 44.165 ;
        RECT -70.685 43.815 -70.285 44.165 ;
        RECT -68.445 43.815 -68.045 44.165 ;
        RECT -66.205 43.815 -65.805 44.165 ;
        RECT -63.965 43.815 -63.565 44.165 ;
        RECT -61.725 43.815 -61.325 44.165 ;
        RECT -59.485 43.815 -59.085 44.165 ;
        RECT -57.245 43.815 -56.845 44.165 ;
        RECT -55.005 43.815 -54.605 44.165 ;
        RECT -52.765 43.815 -52.365 44.165 ;
        RECT -50.525 43.815 -50.125 44.165 ;
        RECT -48.285 43.815 -47.885 44.165 ;
        RECT -46.045 43.815 -45.645 44.165 ;
        RECT -43.805 43.815 -43.405 44.165 ;
        RECT -41.565 43.815 -41.165 44.165 ;
        RECT -39.325 43.815 -38.925 44.165 ;
        RECT -37.085 43.815 -36.685 44.165 ;
        RECT -34.845 43.815 -34.445 44.165 ;
        RECT -32.605 43.815 -32.205 44.165 ;
        RECT -30.365 43.815 -29.965 44.165 ;
        RECT -28.125 43.815 -27.725 44.165 ;
        RECT -25.885 43.815 -25.485 44.165 ;
        RECT -23.645 43.815 -23.245 44.165 ;
        RECT -21.405 43.815 -21.005 44.165 ;
        RECT -19.165 43.815 -18.765 44.165 ;
        RECT -16.925 43.815 -16.525 44.165 ;
        RECT -14.685 43.815 -14.285 44.165 ;
        RECT -12.445 43.815 -12.045 44.165 ;
        RECT -10.205 43.815 -9.805 44.165 ;
        RECT -7.965 43.815 -7.565 44.165 ;
        RECT -5.725 43.815 -5.325 44.165 ;
        RECT -3.485 43.815 -3.085 44.165 ;
        RECT -1.245 43.815 -0.845 44.165 ;
        RECT 0.995 43.815 1.395 44.165 ;
        RECT 3.235 43.815 3.635 44.165 ;
        RECT 5.475 43.815 5.875 44.165 ;
        RECT 7.715 43.815 8.115 44.165 ;
        RECT 9.955 43.815 10.355 44.165 ;
        RECT 12.195 43.815 12.595 44.165 ;
        RECT 14.435 43.815 14.835 44.165 ;
        RECT 16.675 43.815 17.075 44.165 ;
        RECT 18.915 43.815 19.315 44.165 ;
        RECT 21.155 43.815 21.555 44.165 ;
        RECT 23.395 43.815 23.795 44.165 ;
        RECT 25.635 43.815 26.035 44.165 ;
        RECT 27.875 43.815 28.275 44.165 ;
        RECT 30.115 43.815 30.515 44.165 ;
        RECT 32.355 43.815 32.755 44.165 ;
        RECT 34.595 43.815 34.995 44.165 ;
        RECT 36.835 43.815 37.235 44.165 ;
        RECT 39.075 43.815 39.475 44.165 ;
        RECT 41.315 43.815 41.715 44.165 ;
        RECT 43.555 43.815 43.955 44.165 ;
        RECT 45.795 43.815 46.195 44.165 ;
        RECT 48.035 43.815 48.435 44.165 ;
        RECT 50.275 43.815 50.675 44.165 ;
        RECT 52.515 43.815 52.915 44.165 ;
        RECT 54.755 43.815 55.155 44.165 ;
        RECT 56.995 43.815 57.395 44.165 ;
        RECT 59.235 43.815 59.635 44.165 ;
        RECT 61.475 43.815 61.875 44.165 ;
        RECT 63.715 43.815 64.115 44.165 ;
        RECT 65.955 43.815 66.355 44.165 ;
        RECT 68.195 43.815 68.595 44.165 ;
        RECT 70.435 43.815 70.835 44.165 ;
        RECT 72.675 43.815 73.075 44.165 ;
        RECT 74.915 43.815 75.315 44.165 ;
        RECT 77.155 43.815 77.555 44.165 ;
        RECT 79.395 43.815 79.795 44.165 ;
        RECT 81.635 43.815 82.035 44.165 ;
        RECT 83.875 43.815 84.275 44.165 ;
        RECT 86.115 43.815 86.515 44.165 ;
        RECT 88.355 43.815 88.755 44.165 ;
        RECT 90.595 43.815 90.995 44.165 ;
        RECT 92.835 43.815 93.235 44.165 ;
        RECT 95.075 43.815 95.475 44.165 ;
        RECT 97.315 43.815 97.715 44.165 ;
        RECT -497.305 42.300 -486.905 42.900 ;
        RECT -497.305 34.300 -495.505 42.300 ;
        RECT -487.505 34.300 -486.905 42.300 ;
        RECT -473.885 41.305 -473.485 41.655 ;
        RECT -469.405 41.305 -469.005 41.655 ;
        RECT -464.925 41.305 -464.525 41.655 ;
        RECT -460.445 41.305 -460.045 41.655 ;
        RECT -455.965 41.305 -455.565 41.655 ;
        RECT -451.485 41.305 -451.085 41.655 ;
        RECT -447.005 41.305 -446.605 41.655 ;
        RECT -442.525 41.305 -442.125 41.655 ;
        RECT -438.045 41.305 -437.645 41.655 ;
        RECT -433.565 41.305 -433.165 41.655 ;
        RECT -429.085 41.305 -428.685 41.655 ;
        RECT -424.605 41.305 -424.205 41.655 ;
        RECT -420.125 41.305 -419.725 41.655 ;
        RECT -415.645 41.305 -415.245 41.655 ;
        RECT -411.165 41.305 -410.765 41.655 ;
        RECT -406.685 41.305 -406.285 41.655 ;
        RECT -402.205 41.305 -401.805 41.655 ;
        RECT -397.725 41.305 -397.325 41.655 ;
        RECT -393.245 41.305 -392.845 41.655 ;
        RECT -388.765 41.305 -388.365 41.655 ;
        RECT -384.285 41.305 -383.885 41.655 ;
        RECT -379.805 41.305 -379.405 41.655 ;
        RECT -375.325 41.305 -374.925 41.655 ;
        RECT -370.845 41.305 -370.445 41.655 ;
        RECT -366.365 41.305 -365.965 41.655 ;
        RECT -361.885 41.305 -361.485 41.655 ;
        RECT -357.405 41.305 -357.005 41.655 ;
        RECT -352.925 41.305 -352.525 41.655 ;
        RECT -348.445 41.305 -348.045 41.655 ;
        RECT -343.965 41.305 -343.565 41.655 ;
        RECT -339.485 41.305 -339.085 41.655 ;
        RECT -335.005 41.305 -334.605 41.655 ;
        RECT -330.525 41.305 -330.125 41.655 ;
        RECT -326.045 41.305 -325.645 41.655 ;
        RECT -321.565 41.305 -321.165 41.655 ;
        RECT -317.085 41.305 -316.685 41.655 ;
        RECT -312.605 41.305 -312.205 41.655 ;
        RECT -308.125 41.305 -307.725 41.655 ;
        RECT -303.645 41.305 -303.245 41.655 ;
        RECT -299.165 41.305 -298.765 41.655 ;
        RECT -294.685 41.305 -294.285 41.655 ;
        RECT -290.205 41.305 -289.805 41.655 ;
        RECT -285.725 41.305 -285.325 41.655 ;
        RECT -281.245 41.305 -280.845 41.655 ;
        RECT -276.765 41.305 -276.365 41.655 ;
        RECT -272.285 41.305 -271.885 41.655 ;
        RECT -267.805 41.305 -267.405 41.655 ;
        RECT -263.325 41.305 -262.925 41.655 ;
        RECT -258.845 41.305 -258.445 41.655 ;
        RECT -254.365 41.305 -253.965 41.655 ;
        RECT -249.885 41.305 -249.485 41.655 ;
        RECT -245.405 41.305 -245.005 41.655 ;
        RECT -240.925 41.305 -240.525 41.655 ;
        RECT -236.445 41.305 -236.045 41.655 ;
        RECT -231.965 41.305 -231.565 41.655 ;
        RECT -227.485 41.305 -227.085 41.655 ;
        RECT -223.005 41.305 -222.605 41.655 ;
        RECT -218.525 41.305 -218.125 41.655 ;
        RECT -214.045 41.305 -213.645 41.655 ;
        RECT -209.565 41.305 -209.165 41.655 ;
        RECT -205.085 41.305 -204.685 41.655 ;
        RECT -200.605 41.305 -200.205 41.655 ;
        RECT -196.125 41.305 -195.725 41.655 ;
        RECT -191.645 41.305 -191.245 41.655 ;
        RECT -186.045 41.305 -185.645 41.655 ;
        RECT -181.565 41.305 -181.165 41.655 ;
        RECT -177.085 41.305 -176.685 41.655 ;
        RECT -172.605 41.305 -172.205 41.655 ;
        RECT -168.125 41.305 -167.725 41.655 ;
        RECT -163.645 41.305 -163.245 41.655 ;
        RECT -159.165 41.305 -158.765 41.655 ;
        RECT -154.685 41.305 -154.285 41.655 ;
        RECT -150.205 41.305 -149.805 41.655 ;
        RECT -145.725 41.305 -145.325 41.655 ;
        RECT -141.245 41.305 -140.845 41.655 ;
        RECT -136.765 41.305 -136.365 41.655 ;
        RECT -132.285 41.305 -131.885 41.655 ;
        RECT -127.805 41.305 -127.405 41.655 ;
        RECT -123.325 41.305 -122.925 41.655 ;
        RECT -118.845 41.305 -118.445 41.655 ;
        RECT -114.365 41.305 -113.965 41.655 ;
        RECT -109.885 41.305 -109.485 41.655 ;
        RECT -105.405 41.305 -105.005 41.655 ;
        RECT -100.925 41.305 -100.525 41.655 ;
        RECT -96.445 41.305 -96.045 41.655 ;
        RECT -91.965 41.305 -91.565 41.655 ;
        RECT -87.485 41.305 -87.085 41.655 ;
        RECT -83.005 41.305 -82.605 41.655 ;
        RECT -78.525 41.305 -78.125 41.655 ;
        RECT -74.045 41.305 -73.645 41.655 ;
        RECT -69.565 41.305 -69.165 41.655 ;
        RECT -65.085 41.305 -64.685 41.655 ;
        RECT -60.605 41.305 -60.205 41.655 ;
        RECT -56.125 41.305 -55.725 41.655 ;
        RECT -51.645 41.305 -51.245 41.655 ;
        RECT -47.165 41.305 -46.765 41.655 ;
        RECT -42.685 41.305 -42.285 41.655 ;
        RECT -38.205 41.305 -37.805 41.655 ;
        RECT -33.725 41.305 -33.325 41.655 ;
        RECT -29.245 41.305 -28.845 41.655 ;
        RECT -24.765 41.305 -24.365 41.655 ;
        RECT -20.285 41.305 -19.885 41.655 ;
        RECT -15.805 41.305 -15.405 41.655 ;
        RECT -11.325 41.305 -10.925 41.655 ;
        RECT -6.845 41.305 -6.445 41.655 ;
        RECT -2.365 41.305 -1.965 41.655 ;
        RECT 2.115 41.305 2.515 41.655 ;
        RECT 6.595 41.305 6.995 41.655 ;
        RECT 11.075 41.305 11.475 41.655 ;
        RECT 15.555 41.305 15.955 41.655 ;
        RECT 20.035 41.305 20.435 41.655 ;
        RECT 24.515 41.305 24.915 41.655 ;
        RECT 28.995 41.305 29.395 41.655 ;
        RECT 33.475 41.305 33.875 41.655 ;
        RECT 37.955 41.305 38.355 41.655 ;
        RECT 42.435 41.305 42.835 41.655 ;
        RECT 46.915 41.305 47.315 41.655 ;
        RECT 51.395 41.305 51.795 41.655 ;
        RECT 55.875 41.305 56.275 41.655 ;
        RECT 60.355 41.305 60.755 41.655 ;
        RECT 64.835 41.305 65.235 41.655 ;
        RECT 69.315 41.305 69.715 41.655 ;
        RECT 73.795 41.305 74.195 41.655 ;
        RECT 78.275 41.305 78.675 41.655 ;
        RECT 82.755 41.305 83.155 41.655 ;
        RECT 87.235 41.305 87.635 41.655 ;
        RECT 91.715 41.305 92.115 41.655 ;
        RECT 96.195 41.305 96.595 41.655 ;
        RECT -473.885 41.255 103.755 41.305 ;
        RECT -473.885 40.855 104.155 41.255 ;
        RECT -473.885 40.805 103.755 40.855 ;
        RECT -473.885 40.455 -473.485 40.805 ;
        RECT -469.405 40.455 -469.005 40.805 ;
        RECT -464.925 40.455 -464.525 40.805 ;
        RECT -460.445 40.455 -460.045 40.805 ;
        RECT -455.965 40.455 -455.565 40.805 ;
        RECT -451.485 40.455 -451.085 40.805 ;
        RECT -447.005 40.455 -446.605 40.805 ;
        RECT -442.525 40.455 -442.125 40.805 ;
        RECT -438.045 40.455 -437.645 40.805 ;
        RECT -433.565 40.455 -433.165 40.805 ;
        RECT -429.085 40.455 -428.685 40.805 ;
        RECT -424.605 40.455 -424.205 40.805 ;
        RECT -420.125 40.455 -419.725 40.805 ;
        RECT -415.645 40.455 -415.245 40.805 ;
        RECT -411.165 40.455 -410.765 40.805 ;
        RECT -406.685 40.455 -406.285 40.805 ;
        RECT -402.205 40.455 -401.805 40.805 ;
        RECT -397.725 40.455 -397.325 40.805 ;
        RECT -393.245 40.455 -392.845 40.805 ;
        RECT -388.765 40.455 -388.365 40.805 ;
        RECT -384.285 40.455 -383.885 40.805 ;
        RECT -379.805 40.455 -379.405 40.805 ;
        RECT -375.325 40.455 -374.925 40.805 ;
        RECT -370.845 40.455 -370.445 40.805 ;
        RECT -366.365 40.455 -365.965 40.805 ;
        RECT -361.885 40.455 -361.485 40.805 ;
        RECT -357.405 40.455 -357.005 40.805 ;
        RECT -352.925 40.455 -352.525 40.805 ;
        RECT -348.445 40.455 -348.045 40.805 ;
        RECT -343.965 40.455 -343.565 40.805 ;
        RECT -339.485 40.455 -339.085 40.805 ;
        RECT -335.005 40.455 -334.605 40.805 ;
        RECT -330.525 40.455 -330.125 40.805 ;
        RECT -326.045 40.455 -325.645 40.805 ;
        RECT -321.565 40.455 -321.165 40.805 ;
        RECT -317.085 40.455 -316.685 40.805 ;
        RECT -312.605 40.455 -312.205 40.805 ;
        RECT -308.125 40.455 -307.725 40.805 ;
        RECT -303.645 40.455 -303.245 40.805 ;
        RECT -299.165 40.455 -298.765 40.805 ;
        RECT -294.685 40.455 -294.285 40.805 ;
        RECT -290.205 40.455 -289.805 40.805 ;
        RECT -285.725 40.455 -285.325 40.805 ;
        RECT -281.245 40.455 -280.845 40.805 ;
        RECT -276.765 40.455 -276.365 40.805 ;
        RECT -272.285 40.455 -271.885 40.805 ;
        RECT -267.805 40.455 -267.405 40.805 ;
        RECT -263.325 40.455 -262.925 40.805 ;
        RECT -258.845 40.455 -258.445 40.805 ;
        RECT -254.365 40.455 -253.965 40.805 ;
        RECT -249.885 40.455 -249.485 40.805 ;
        RECT -245.405 40.455 -245.005 40.805 ;
        RECT -240.925 40.455 -240.525 40.805 ;
        RECT -236.445 40.455 -236.045 40.805 ;
        RECT -231.965 40.455 -231.565 40.805 ;
        RECT -227.485 40.455 -227.085 40.805 ;
        RECT -223.005 40.455 -222.605 40.805 ;
        RECT -218.525 40.455 -218.125 40.805 ;
        RECT -214.045 40.455 -213.645 40.805 ;
        RECT -209.565 40.455 -209.165 40.805 ;
        RECT -205.085 40.455 -204.685 40.805 ;
        RECT -200.605 40.455 -200.205 40.805 ;
        RECT -196.125 40.455 -195.725 40.805 ;
        RECT -191.645 40.455 -191.245 40.805 ;
        RECT -186.045 40.455 -185.645 40.805 ;
        RECT -181.565 40.455 -181.165 40.805 ;
        RECT -177.085 40.455 -176.685 40.805 ;
        RECT -172.605 40.455 -172.205 40.805 ;
        RECT -168.125 40.455 -167.725 40.805 ;
        RECT -163.645 40.455 -163.245 40.805 ;
        RECT -159.165 40.455 -158.765 40.805 ;
        RECT -154.685 40.455 -154.285 40.805 ;
        RECT -150.205 40.455 -149.805 40.805 ;
        RECT -145.725 40.455 -145.325 40.805 ;
        RECT -141.245 40.455 -140.845 40.805 ;
        RECT -136.765 40.455 -136.365 40.805 ;
        RECT -132.285 40.455 -131.885 40.805 ;
        RECT -127.805 40.455 -127.405 40.805 ;
        RECT -123.325 40.455 -122.925 40.805 ;
        RECT -118.845 40.455 -118.445 40.805 ;
        RECT -114.365 40.455 -113.965 40.805 ;
        RECT -109.885 40.455 -109.485 40.805 ;
        RECT -105.405 40.455 -105.005 40.805 ;
        RECT -100.925 40.455 -100.525 40.805 ;
        RECT -96.445 40.455 -96.045 40.805 ;
        RECT -91.965 40.455 -91.565 40.805 ;
        RECT -87.485 40.455 -87.085 40.805 ;
        RECT -83.005 40.455 -82.605 40.805 ;
        RECT -78.525 40.455 -78.125 40.805 ;
        RECT -74.045 40.455 -73.645 40.805 ;
        RECT -69.565 40.455 -69.165 40.805 ;
        RECT -65.085 40.455 -64.685 40.805 ;
        RECT -60.605 40.455 -60.205 40.805 ;
        RECT -56.125 40.455 -55.725 40.805 ;
        RECT -51.645 40.455 -51.245 40.805 ;
        RECT -47.165 40.455 -46.765 40.805 ;
        RECT -42.685 40.455 -42.285 40.805 ;
        RECT -38.205 40.455 -37.805 40.805 ;
        RECT -33.725 40.455 -33.325 40.805 ;
        RECT -29.245 40.455 -28.845 40.805 ;
        RECT -24.765 40.455 -24.365 40.805 ;
        RECT -20.285 40.455 -19.885 40.805 ;
        RECT -15.805 40.455 -15.405 40.805 ;
        RECT -11.325 40.455 -10.925 40.805 ;
        RECT -6.845 40.455 -6.445 40.805 ;
        RECT -2.365 40.455 -1.965 40.805 ;
        RECT 2.115 40.455 2.515 40.805 ;
        RECT 6.595 40.455 6.995 40.805 ;
        RECT 11.075 40.455 11.475 40.805 ;
        RECT 15.555 40.455 15.955 40.805 ;
        RECT 20.035 40.455 20.435 40.805 ;
        RECT 24.515 40.455 24.915 40.805 ;
        RECT 28.995 40.455 29.395 40.805 ;
        RECT 33.475 40.455 33.875 40.805 ;
        RECT 37.955 40.455 38.355 40.805 ;
        RECT 42.435 40.455 42.835 40.805 ;
        RECT 46.915 40.455 47.315 40.805 ;
        RECT 51.395 40.455 51.795 40.805 ;
        RECT 55.875 40.455 56.275 40.805 ;
        RECT 60.355 40.455 60.755 40.805 ;
        RECT 64.835 40.455 65.235 40.805 ;
        RECT 69.315 40.455 69.715 40.805 ;
        RECT 73.795 40.455 74.195 40.805 ;
        RECT 78.275 40.455 78.675 40.805 ;
        RECT 82.755 40.455 83.155 40.805 ;
        RECT 87.235 40.455 87.635 40.805 ;
        RECT 91.715 40.455 92.115 40.805 ;
        RECT 96.195 40.455 96.595 40.805 ;
        RECT -471.645 37.945 -471.245 38.295 ;
        RECT -462.685 37.945 -462.285 38.295 ;
        RECT -453.725 37.945 -453.325 38.295 ;
        RECT -444.765 37.945 -444.365 38.295 ;
        RECT -435.805 37.945 -435.405 38.295 ;
        RECT -426.845 37.945 -426.445 38.295 ;
        RECT -417.885 37.945 -417.485 38.295 ;
        RECT -408.925 37.945 -408.525 38.295 ;
        RECT -399.965 37.945 -399.565 38.295 ;
        RECT -391.005 37.945 -390.605 38.295 ;
        RECT -382.045 37.945 -381.645 38.295 ;
        RECT -373.085 37.945 -372.685 38.295 ;
        RECT -364.125 37.945 -363.725 38.295 ;
        RECT -355.165 37.945 -354.765 38.295 ;
        RECT -346.205 37.945 -345.805 38.295 ;
        RECT -337.245 37.945 -336.845 38.295 ;
        RECT -328.285 37.945 -327.885 38.295 ;
        RECT -319.325 37.945 -318.925 38.295 ;
        RECT -310.365 37.945 -309.965 38.295 ;
        RECT -301.405 37.945 -301.005 38.295 ;
        RECT -292.445 37.945 -292.045 38.295 ;
        RECT -283.485 37.945 -283.085 38.295 ;
        RECT -274.525 37.945 -274.125 38.295 ;
        RECT -265.565 37.945 -265.165 38.295 ;
        RECT -256.605 37.945 -256.205 38.295 ;
        RECT -247.645 37.945 -247.245 38.295 ;
        RECT -238.685 37.945 -238.285 38.295 ;
        RECT -229.725 37.945 -229.325 38.295 ;
        RECT -220.765 37.945 -220.365 38.295 ;
        RECT -211.805 37.945 -211.405 38.295 ;
        RECT -202.845 37.945 -202.445 38.295 ;
        RECT -193.885 37.945 -193.485 38.295 ;
        RECT -183.805 37.945 -183.405 38.295 ;
        RECT -174.845 37.945 -174.445 38.295 ;
        RECT -165.885 37.945 -165.485 38.295 ;
        RECT -156.925 37.945 -156.525 38.295 ;
        RECT -147.965 37.945 -147.565 38.295 ;
        RECT -139.005 37.945 -138.605 38.295 ;
        RECT -130.045 37.945 -129.645 38.295 ;
        RECT -121.085 37.945 -120.685 38.295 ;
        RECT -112.125 37.945 -111.725 38.295 ;
        RECT -103.165 37.945 -102.765 38.295 ;
        RECT -94.205 37.945 -93.805 38.295 ;
        RECT -85.245 37.945 -84.845 38.295 ;
        RECT -76.285 37.945 -75.885 38.295 ;
        RECT -67.325 37.945 -66.925 38.295 ;
        RECT -58.365 37.945 -57.965 38.295 ;
        RECT -49.405 37.945 -49.005 38.295 ;
        RECT -40.445 37.945 -40.045 38.295 ;
        RECT -31.485 37.945 -31.085 38.295 ;
        RECT -22.525 37.945 -22.125 38.295 ;
        RECT -13.565 37.945 -13.165 38.295 ;
        RECT -4.605 37.945 -4.205 38.295 ;
        RECT 4.355 37.945 4.755 38.295 ;
        RECT 13.315 37.945 13.715 38.295 ;
        RECT 22.275 37.945 22.675 38.295 ;
        RECT 31.235 37.945 31.635 38.295 ;
        RECT 40.195 37.945 40.595 38.295 ;
        RECT 49.155 37.945 49.555 38.295 ;
        RECT 58.115 37.945 58.515 38.295 ;
        RECT 67.075 37.945 67.475 38.295 ;
        RECT 76.035 37.945 76.435 38.295 ;
        RECT 84.995 37.945 85.395 38.295 ;
        RECT 93.955 37.945 94.355 38.295 ;
        RECT -471.645 37.895 105.555 37.945 ;
        RECT -471.645 37.495 105.955 37.895 ;
        RECT -471.645 37.445 105.555 37.495 ;
        RECT -471.645 37.095 -471.245 37.445 ;
        RECT -462.685 37.095 -462.285 37.445 ;
        RECT -453.725 37.095 -453.325 37.445 ;
        RECT -444.765 37.095 -444.365 37.445 ;
        RECT -435.805 37.095 -435.405 37.445 ;
        RECT -426.845 37.095 -426.445 37.445 ;
        RECT -417.885 37.095 -417.485 37.445 ;
        RECT -408.925 37.095 -408.525 37.445 ;
        RECT -399.965 37.095 -399.565 37.445 ;
        RECT -391.005 37.095 -390.605 37.445 ;
        RECT -382.045 37.095 -381.645 37.445 ;
        RECT -373.085 37.095 -372.685 37.445 ;
        RECT -364.125 37.095 -363.725 37.445 ;
        RECT -355.165 37.095 -354.765 37.445 ;
        RECT -346.205 37.095 -345.805 37.445 ;
        RECT -337.245 37.095 -336.845 37.445 ;
        RECT -328.285 37.095 -327.885 37.445 ;
        RECT -319.325 37.095 -318.925 37.445 ;
        RECT -310.365 37.095 -309.965 37.445 ;
        RECT -301.405 37.095 -301.005 37.445 ;
        RECT -292.445 37.095 -292.045 37.445 ;
        RECT -283.485 37.095 -283.085 37.445 ;
        RECT -274.525 37.095 -274.125 37.445 ;
        RECT -265.565 37.095 -265.165 37.445 ;
        RECT -256.605 37.095 -256.205 37.445 ;
        RECT -247.645 37.095 -247.245 37.445 ;
        RECT -238.685 37.095 -238.285 37.445 ;
        RECT -229.725 37.095 -229.325 37.445 ;
        RECT -220.765 37.095 -220.365 37.445 ;
        RECT -211.805 37.095 -211.405 37.445 ;
        RECT -202.845 37.095 -202.445 37.445 ;
        RECT -193.885 37.095 -193.485 37.445 ;
        RECT -183.805 37.095 -183.405 37.445 ;
        RECT -174.845 37.095 -174.445 37.445 ;
        RECT -165.885 37.095 -165.485 37.445 ;
        RECT -156.925 37.095 -156.525 37.445 ;
        RECT -147.965 37.095 -147.565 37.445 ;
        RECT -139.005 37.095 -138.605 37.445 ;
        RECT -130.045 37.095 -129.645 37.445 ;
        RECT -121.085 37.095 -120.685 37.445 ;
        RECT -112.125 37.095 -111.725 37.445 ;
        RECT -103.165 37.095 -102.765 37.445 ;
        RECT -94.205 37.095 -93.805 37.445 ;
        RECT -85.245 37.095 -84.845 37.445 ;
        RECT -76.285 37.095 -75.885 37.445 ;
        RECT -67.325 37.095 -66.925 37.445 ;
        RECT -58.365 37.095 -57.965 37.445 ;
        RECT -49.405 37.095 -49.005 37.445 ;
        RECT -40.445 37.095 -40.045 37.445 ;
        RECT -31.485 37.095 -31.085 37.445 ;
        RECT -22.525 37.095 -22.125 37.445 ;
        RECT -13.565 37.095 -13.165 37.445 ;
        RECT -4.605 37.095 -4.205 37.445 ;
        RECT 4.355 37.095 4.755 37.445 ;
        RECT 13.315 37.095 13.715 37.445 ;
        RECT 22.275 37.095 22.675 37.445 ;
        RECT 31.235 37.095 31.635 37.445 ;
        RECT 40.195 37.095 40.595 37.445 ;
        RECT 49.155 37.095 49.555 37.445 ;
        RECT 58.115 37.095 58.515 37.445 ;
        RECT 67.075 37.095 67.475 37.445 ;
        RECT 76.035 37.095 76.435 37.445 ;
        RECT 84.995 37.095 85.395 37.445 ;
        RECT 93.955 37.095 94.355 37.445 ;
        RECT -497.305 33.700 -486.905 34.300 ;
        RECT -467.165 34.585 -466.765 34.935 ;
        RECT -449.245 34.585 -448.845 34.935 ;
        RECT -431.325 34.585 -430.925 34.935 ;
        RECT -413.405 34.585 -413.005 34.935 ;
        RECT -395.485 34.585 -395.085 34.935 ;
        RECT -377.565 34.585 -377.165 34.935 ;
        RECT -359.645 34.585 -359.245 34.935 ;
        RECT -341.725 34.585 -341.325 34.935 ;
        RECT -323.805 34.585 -323.405 34.935 ;
        RECT -305.885 34.585 -305.485 34.935 ;
        RECT -287.965 34.585 -287.565 34.935 ;
        RECT -270.045 34.585 -269.645 34.935 ;
        RECT -252.125 34.585 -251.725 34.935 ;
        RECT -234.205 34.585 -233.805 34.935 ;
        RECT -216.285 34.585 -215.885 34.935 ;
        RECT -198.365 34.585 -197.965 34.935 ;
        RECT -179.325 34.585 -178.925 34.935 ;
        RECT -161.405 34.585 -161.005 34.935 ;
        RECT -143.485 34.585 -143.085 34.935 ;
        RECT -125.565 34.585 -125.165 34.935 ;
        RECT -107.645 34.585 -107.245 34.935 ;
        RECT -89.725 34.585 -89.325 34.935 ;
        RECT -71.805 34.585 -71.405 34.935 ;
        RECT -53.885 34.585 -53.485 34.935 ;
        RECT -35.965 34.585 -35.565 34.935 ;
        RECT -18.045 34.585 -17.645 34.935 ;
        RECT -0.125 34.585 0.275 34.935 ;
        RECT 17.795 34.585 18.195 34.935 ;
        RECT 35.715 34.585 36.115 34.935 ;
        RECT 53.635 34.585 54.035 34.935 ;
        RECT 71.555 34.585 71.955 34.935 ;
        RECT 89.475 34.585 89.875 34.935 ;
        RECT -467.165 34.535 107.355 34.585 ;
        RECT -467.165 34.135 107.755 34.535 ;
        RECT -467.165 34.085 107.355 34.135 ;
        RECT -467.165 33.735 -466.765 34.085 ;
        RECT -449.245 33.735 -448.845 34.085 ;
        RECT -431.325 33.735 -430.925 34.085 ;
        RECT -413.405 33.735 -413.005 34.085 ;
        RECT -395.485 33.735 -395.085 34.085 ;
        RECT -377.565 33.735 -377.165 34.085 ;
        RECT -359.645 33.735 -359.245 34.085 ;
        RECT -341.725 33.735 -341.325 34.085 ;
        RECT -323.805 33.735 -323.405 34.085 ;
        RECT -305.885 33.735 -305.485 34.085 ;
        RECT -287.965 33.735 -287.565 34.085 ;
        RECT -270.045 33.735 -269.645 34.085 ;
        RECT -252.125 33.735 -251.725 34.085 ;
        RECT -234.205 33.735 -233.805 34.085 ;
        RECT -216.285 33.735 -215.885 34.085 ;
        RECT -198.365 33.735 -197.965 34.085 ;
        RECT -179.325 33.735 -178.925 34.085 ;
        RECT -161.405 33.735 -161.005 34.085 ;
        RECT -143.485 33.735 -143.085 34.085 ;
        RECT -125.565 33.735 -125.165 34.085 ;
        RECT -107.645 33.735 -107.245 34.085 ;
        RECT -89.725 33.735 -89.325 34.085 ;
        RECT -71.805 33.735 -71.405 34.085 ;
        RECT -53.885 33.735 -53.485 34.085 ;
        RECT -35.965 33.735 -35.565 34.085 ;
        RECT -18.045 33.735 -17.645 34.085 ;
        RECT -0.125 33.735 0.275 34.085 ;
        RECT 17.795 33.735 18.195 34.085 ;
        RECT 35.715 33.735 36.115 34.085 ;
        RECT 53.635 33.735 54.035 34.085 ;
        RECT 71.555 33.735 71.955 34.085 ;
        RECT 89.475 33.735 89.875 34.085 ;
        RECT -458.205 31.225 -457.805 31.575 ;
        RECT -422.365 31.225 -421.965 31.575 ;
        RECT -386.525 31.225 -386.125 31.575 ;
        RECT -350.685 31.225 -350.285 31.575 ;
        RECT -314.845 31.225 -314.445 31.575 ;
        RECT -279.005 31.225 -278.605 31.575 ;
        RECT -243.165 31.225 -242.765 31.575 ;
        RECT -207.325 31.225 -206.925 31.575 ;
        RECT -170.365 31.225 -169.965 31.575 ;
        RECT -134.525 31.225 -134.125 31.575 ;
        RECT -98.685 31.225 -98.285 31.575 ;
        RECT -62.845 31.225 -62.445 31.575 ;
        RECT -27.005 31.225 -26.605 31.575 ;
        RECT 8.835 31.225 9.235 31.575 ;
        RECT 44.675 31.225 45.075 31.575 ;
        RECT 80.515 31.225 80.915 31.575 ;
        RECT -458.205 31.175 109.155 31.225 ;
        RECT -497.305 30.300 -486.905 30.900 ;
        RECT -458.205 30.775 109.555 31.175 ;
        RECT -458.205 30.725 109.155 30.775 ;
        RECT -458.205 30.375 -457.805 30.725 ;
        RECT -422.365 30.375 -421.965 30.725 ;
        RECT -386.525 30.375 -386.125 30.725 ;
        RECT -350.685 30.375 -350.285 30.725 ;
        RECT -314.845 30.375 -314.445 30.725 ;
        RECT -279.005 30.375 -278.605 30.725 ;
        RECT -243.165 30.375 -242.765 30.725 ;
        RECT -207.325 30.375 -206.925 30.725 ;
        RECT -170.365 30.375 -169.965 30.725 ;
        RECT -134.525 30.375 -134.125 30.725 ;
        RECT -98.685 30.375 -98.285 30.725 ;
        RECT -62.845 30.375 -62.445 30.725 ;
        RECT -27.005 30.375 -26.605 30.725 ;
        RECT 8.835 30.375 9.235 30.725 ;
        RECT 44.675 30.375 45.075 30.725 ;
        RECT 80.515 30.375 80.915 30.725 ;
        RECT -497.305 22.300 -495.505 30.300 ;
        RECT -487.505 22.300 -486.905 30.300 ;
        RECT -440.285 27.865 -439.885 28.215 ;
        RECT -368.605 27.865 -368.205 28.215 ;
        RECT -296.925 27.865 -296.525 28.215 ;
        RECT -225.245 27.865 -224.845 28.215 ;
        RECT -152.445 27.865 -152.045 28.215 ;
        RECT -80.765 27.865 -80.365 28.215 ;
        RECT -9.085 27.865 -8.685 28.215 ;
        RECT 62.595 27.865 62.995 28.215 ;
        RECT -440.285 27.815 110.955 27.865 ;
        RECT -440.285 27.415 111.355 27.815 ;
        RECT -440.285 27.365 110.955 27.415 ;
        RECT -440.285 27.015 -439.885 27.365 ;
        RECT -368.605 27.015 -368.205 27.365 ;
        RECT -296.925 27.015 -296.525 27.365 ;
        RECT -225.245 27.015 -224.845 27.365 ;
        RECT -152.445 27.015 -152.045 27.365 ;
        RECT -80.765 27.015 -80.365 27.365 ;
        RECT -9.085 27.015 -8.685 27.365 ;
        RECT 62.595 27.015 62.995 27.365 ;
        RECT -404.445 24.505 -404.045 24.855 ;
        RECT -261.085 24.505 -260.685 24.855 ;
        RECT -116.605 24.505 -116.205 24.855 ;
        RECT 26.755 24.505 27.155 24.855 ;
        RECT -404.445 24.455 112.755 24.505 ;
        RECT -404.445 24.055 113.155 24.455 ;
        RECT -404.445 24.005 112.755 24.055 ;
        RECT -404.445 23.655 -404.045 24.005 ;
        RECT -261.085 23.655 -260.685 24.005 ;
        RECT -116.605 23.655 -116.205 24.005 ;
        RECT 26.755 23.655 27.155 24.005 ;
        RECT -497.305 21.700 -486.905 22.300 ;
        RECT -332.765 21.145 -332.365 21.495 ;
        RECT -44.925 21.145 -44.525 21.495 ;
        RECT -332.765 21.095 114.555 21.145 ;
        RECT -332.765 20.695 114.955 21.095 ;
        RECT -332.765 20.645 114.555 20.695 ;
        RECT -332.765 20.295 -332.365 20.645 ;
        RECT -44.925 20.295 -44.525 20.645 ;
        RECT -188.285 17.785 -187.885 18.135 ;
        RECT -188.285 17.735 116.355 17.785 ;
        RECT -188.285 17.335 116.755 17.735 ;
        RECT -188.285 17.285 116.355 17.335 ;
        RECT -188.285 16.935 -187.885 17.285 ;
        RECT -189.405 14.425 -189.005 14.775 ;
        RECT 117.705 14.425 118.205 63.665 ;
        RECT -189.405 14.175 118.205 14.425 ;
        RECT -189.405 13.925 118.155 14.175 ;
        RECT -189.405 13.575 -189.005 13.925 ;
        RECT 239.520 7.720 243.520 117.620 ;
        RECT 235.860 1.720 243.520 7.720 ;
        RECT 239.520 -4.265 243.520 1.720 ;
        RECT 229.700 -5.865 243.520 -4.265 ;
        RECT -189.405 -13.925 -189.005 -13.575 ;
        RECT -189.405 -14.175 118.155 -13.925 ;
        RECT -189.405 -14.425 118.205 -14.175 ;
        RECT -189.405 -14.775 -189.005 -14.425 ;
        RECT -188.285 -17.285 -187.885 -16.935 ;
        RECT -188.285 -17.335 116.355 -17.285 ;
        RECT -188.285 -17.735 116.755 -17.335 ;
        RECT -188.285 -17.785 116.355 -17.735 ;
        RECT -188.285 -18.135 -187.885 -17.785 ;
        RECT -332.765 -20.645 -332.365 -20.295 ;
        RECT -44.925 -20.645 -44.525 -20.295 ;
        RECT -332.765 -20.695 114.555 -20.645 ;
        RECT -332.765 -21.095 114.955 -20.695 ;
        RECT -332.765 -21.145 114.555 -21.095 ;
        RECT -332.765 -21.495 -332.365 -21.145 ;
        RECT -44.925 -21.495 -44.525 -21.145 ;
        RECT -497.305 -22.300 -486.905 -21.700 ;
        RECT -497.305 -30.300 -495.505 -22.300 ;
        RECT -487.505 -30.300 -486.905 -22.300 ;
        RECT -404.445 -24.005 -404.045 -23.655 ;
        RECT -261.085 -24.005 -260.685 -23.655 ;
        RECT -116.605 -24.005 -116.205 -23.655 ;
        RECT 26.755 -24.005 27.155 -23.655 ;
        RECT -404.445 -24.055 112.755 -24.005 ;
        RECT -404.445 -24.455 113.155 -24.055 ;
        RECT -404.445 -24.505 112.755 -24.455 ;
        RECT -404.445 -24.855 -404.045 -24.505 ;
        RECT -261.085 -24.855 -260.685 -24.505 ;
        RECT -116.605 -24.855 -116.205 -24.505 ;
        RECT 26.755 -24.855 27.155 -24.505 ;
        RECT -440.285 -27.365 -439.885 -27.015 ;
        RECT -368.605 -27.365 -368.205 -27.015 ;
        RECT -296.925 -27.365 -296.525 -27.015 ;
        RECT -225.245 -27.365 -224.845 -27.015 ;
        RECT -152.445 -27.365 -152.045 -27.015 ;
        RECT -80.765 -27.365 -80.365 -27.015 ;
        RECT -9.085 -27.365 -8.685 -27.015 ;
        RECT 62.595 -27.365 62.995 -27.015 ;
        RECT -440.285 -27.415 110.955 -27.365 ;
        RECT -440.285 -27.815 111.355 -27.415 ;
        RECT -440.285 -27.865 110.955 -27.815 ;
        RECT -440.285 -28.215 -439.885 -27.865 ;
        RECT -368.605 -28.215 -368.205 -27.865 ;
        RECT -296.925 -28.215 -296.525 -27.865 ;
        RECT -225.245 -28.215 -224.845 -27.865 ;
        RECT -152.445 -28.215 -152.045 -27.865 ;
        RECT -80.765 -28.215 -80.365 -27.865 ;
        RECT -9.085 -28.215 -8.685 -27.865 ;
        RECT 62.595 -28.215 62.995 -27.865 ;
        RECT -497.305 -30.900 -486.905 -30.300 ;
        RECT -458.205 -30.725 -457.805 -30.375 ;
        RECT -422.365 -30.725 -421.965 -30.375 ;
        RECT -386.525 -30.725 -386.125 -30.375 ;
        RECT -350.685 -30.725 -350.285 -30.375 ;
        RECT -314.845 -30.725 -314.445 -30.375 ;
        RECT -279.005 -30.725 -278.605 -30.375 ;
        RECT -243.165 -30.725 -242.765 -30.375 ;
        RECT -207.325 -30.725 -206.925 -30.375 ;
        RECT -170.365 -30.725 -169.965 -30.375 ;
        RECT -134.525 -30.725 -134.125 -30.375 ;
        RECT -98.685 -30.725 -98.285 -30.375 ;
        RECT -62.845 -30.725 -62.445 -30.375 ;
        RECT -27.005 -30.725 -26.605 -30.375 ;
        RECT 8.835 -30.725 9.235 -30.375 ;
        RECT 44.675 -30.725 45.075 -30.375 ;
        RECT 80.515 -30.725 80.915 -30.375 ;
        RECT -458.205 -30.775 109.155 -30.725 ;
        RECT -458.205 -31.175 109.555 -30.775 ;
        RECT -458.205 -31.225 109.155 -31.175 ;
        RECT -458.205 -31.575 -457.805 -31.225 ;
        RECT -422.365 -31.575 -421.965 -31.225 ;
        RECT -386.525 -31.575 -386.125 -31.225 ;
        RECT -350.685 -31.575 -350.285 -31.225 ;
        RECT -314.845 -31.575 -314.445 -31.225 ;
        RECT -279.005 -31.575 -278.605 -31.225 ;
        RECT -243.165 -31.575 -242.765 -31.225 ;
        RECT -207.325 -31.575 -206.925 -31.225 ;
        RECT -170.365 -31.575 -169.965 -31.225 ;
        RECT -134.525 -31.575 -134.125 -31.225 ;
        RECT -98.685 -31.575 -98.285 -31.225 ;
        RECT -62.845 -31.575 -62.445 -31.225 ;
        RECT -27.005 -31.575 -26.605 -31.225 ;
        RECT 8.835 -31.575 9.235 -31.225 ;
        RECT 44.675 -31.575 45.075 -31.225 ;
        RECT 80.515 -31.575 80.915 -31.225 ;
        RECT -497.305 -34.300 -486.905 -33.700 ;
        RECT -497.305 -42.300 -495.505 -34.300 ;
        RECT -487.505 -42.300 -486.905 -34.300 ;
        RECT -467.165 -34.085 -466.765 -33.735 ;
        RECT -449.245 -34.085 -448.845 -33.735 ;
        RECT -431.325 -34.085 -430.925 -33.735 ;
        RECT -413.405 -34.085 -413.005 -33.735 ;
        RECT -395.485 -34.085 -395.085 -33.735 ;
        RECT -377.565 -34.085 -377.165 -33.735 ;
        RECT -359.645 -34.085 -359.245 -33.735 ;
        RECT -341.725 -34.085 -341.325 -33.735 ;
        RECT -323.805 -34.085 -323.405 -33.735 ;
        RECT -305.885 -34.085 -305.485 -33.735 ;
        RECT -287.965 -34.085 -287.565 -33.735 ;
        RECT -270.045 -34.085 -269.645 -33.735 ;
        RECT -252.125 -34.085 -251.725 -33.735 ;
        RECT -234.205 -34.085 -233.805 -33.735 ;
        RECT -216.285 -34.085 -215.885 -33.735 ;
        RECT -198.365 -34.085 -197.965 -33.735 ;
        RECT -179.325 -34.085 -178.925 -33.735 ;
        RECT -161.405 -34.085 -161.005 -33.735 ;
        RECT -143.485 -34.085 -143.085 -33.735 ;
        RECT -125.565 -34.085 -125.165 -33.735 ;
        RECT -107.645 -34.085 -107.245 -33.735 ;
        RECT -89.725 -34.085 -89.325 -33.735 ;
        RECT -71.805 -34.085 -71.405 -33.735 ;
        RECT -53.885 -34.085 -53.485 -33.735 ;
        RECT -35.965 -34.085 -35.565 -33.735 ;
        RECT -18.045 -34.085 -17.645 -33.735 ;
        RECT -0.125 -34.085 0.275 -33.735 ;
        RECT 17.795 -34.085 18.195 -33.735 ;
        RECT 35.715 -34.085 36.115 -33.735 ;
        RECT 53.635 -34.085 54.035 -33.735 ;
        RECT 71.555 -34.085 71.955 -33.735 ;
        RECT 89.475 -34.085 89.875 -33.735 ;
        RECT -467.165 -34.135 107.355 -34.085 ;
        RECT -467.165 -34.535 107.755 -34.135 ;
        RECT -467.165 -34.585 107.355 -34.535 ;
        RECT -467.165 -34.935 -466.765 -34.585 ;
        RECT -449.245 -34.935 -448.845 -34.585 ;
        RECT -431.325 -34.935 -430.925 -34.585 ;
        RECT -413.405 -34.935 -413.005 -34.585 ;
        RECT -395.485 -34.935 -395.085 -34.585 ;
        RECT -377.565 -34.935 -377.165 -34.585 ;
        RECT -359.645 -34.935 -359.245 -34.585 ;
        RECT -341.725 -34.935 -341.325 -34.585 ;
        RECT -323.805 -34.935 -323.405 -34.585 ;
        RECT -305.885 -34.935 -305.485 -34.585 ;
        RECT -287.965 -34.935 -287.565 -34.585 ;
        RECT -270.045 -34.935 -269.645 -34.585 ;
        RECT -252.125 -34.935 -251.725 -34.585 ;
        RECT -234.205 -34.935 -233.805 -34.585 ;
        RECT -216.285 -34.935 -215.885 -34.585 ;
        RECT -198.365 -34.935 -197.965 -34.585 ;
        RECT -179.325 -34.935 -178.925 -34.585 ;
        RECT -161.405 -34.935 -161.005 -34.585 ;
        RECT -143.485 -34.935 -143.085 -34.585 ;
        RECT -125.565 -34.935 -125.165 -34.585 ;
        RECT -107.645 -34.935 -107.245 -34.585 ;
        RECT -89.725 -34.935 -89.325 -34.585 ;
        RECT -71.805 -34.935 -71.405 -34.585 ;
        RECT -53.885 -34.935 -53.485 -34.585 ;
        RECT -35.965 -34.935 -35.565 -34.585 ;
        RECT -18.045 -34.935 -17.645 -34.585 ;
        RECT -0.125 -34.935 0.275 -34.585 ;
        RECT 17.795 -34.935 18.195 -34.585 ;
        RECT 35.715 -34.935 36.115 -34.585 ;
        RECT 53.635 -34.935 54.035 -34.585 ;
        RECT 71.555 -34.935 71.955 -34.585 ;
        RECT 89.475 -34.935 89.875 -34.585 ;
        RECT -471.645 -37.445 -471.245 -37.095 ;
        RECT -462.685 -37.445 -462.285 -37.095 ;
        RECT -453.725 -37.445 -453.325 -37.095 ;
        RECT -444.765 -37.445 -444.365 -37.095 ;
        RECT -435.805 -37.445 -435.405 -37.095 ;
        RECT -426.845 -37.445 -426.445 -37.095 ;
        RECT -417.885 -37.445 -417.485 -37.095 ;
        RECT -408.925 -37.445 -408.525 -37.095 ;
        RECT -399.965 -37.445 -399.565 -37.095 ;
        RECT -391.005 -37.445 -390.605 -37.095 ;
        RECT -382.045 -37.445 -381.645 -37.095 ;
        RECT -373.085 -37.445 -372.685 -37.095 ;
        RECT -364.125 -37.445 -363.725 -37.095 ;
        RECT -355.165 -37.445 -354.765 -37.095 ;
        RECT -346.205 -37.445 -345.805 -37.095 ;
        RECT -337.245 -37.445 -336.845 -37.095 ;
        RECT -328.285 -37.445 -327.885 -37.095 ;
        RECT -319.325 -37.445 -318.925 -37.095 ;
        RECT -310.365 -37.445 -309.965 -37.095 ;
        RECT -301.405 -37.445 -301.005 -37.095 ;
        RECT -292.445 -37.445 -292.045 -37.095 ;
        RECT -283.485 -37.445 -283.085 -37.095 ;
        RECT -274.525 -37.445 -274.125 -37.095 ;
        RECT -265.565 -37.445 -265.165 -37.095 ;
        RECT -256.605 -37.445 -256.205 -37.095 ;
        RECT -247.645 -37.445 -247.245 -37.095 ;
        RECT -238.685 -37.445 -238.285 -37.095 ;
        RECT -229.725 -37.445 -229.325 -37.095 ;
        RECT -220.765 -37.445 -220.365 -37.095 ;
        RECT -211.805 -37.445 -211.405 -37.095 ;
        RECT -202.845 -37.445 -202.445 -37.095 ;
        RECT -193.885 -37.445 -193.485 -37.095 ;
        RECT -183.805 -37.445 -183.405 -37.095 ;
        RECT -174.845 -37.445 -174.445 -37.095 ;
        RECT -165.885 -37.445 -165.485 -37.095 ;
        RECT -156.925 -37.445 -156.525 -37.095 ;
        RECT -147.965 -37.445 -147.565 -37.095 ;
        RECT -139.005 -37.445 -138.605 -37.095 ;
        RECT -130.045 -37.445 -129.645 -37.095 ;
        RECT -121.085 -37.445 -120.685 -37.095 ;
        RECT -112.125 -37.445 -111.725 -37.095 ;
        RECT -103.165 -37.445 -102.765 -37.095 ;
        RECT -94.205 -37.445 -93.805 -37.095 ;
        RECT -85.245 -37.445 -84.845 -37.095 ;
        RECT -76.285 -37.445 -75.885 -37.095 ;
        RECT -67.325 -37.445 -66.925 -37.095 ;
        RECT -58.365 -37.445 -57.965 -37.095 ;
        RECT -49.405 -37.445 -49.005 -37.095 ;
        RECT -40.445 -37.445 -40.045 -37.095 ;
        RECT -31.485 -37.445 -31.085 -37.095 ;
        RECT -22.525 -37.445 -22.125 -37.095 ;
        RECT -13.565 -37.445 -13.165 -37.095 ;
        RECT -4.605 -37.445 -4.205 -37.095 ;
        RECT 4.355 -37.445 4.755 -37.095 ;
        RECT 13.315 -37.445 13.715 -37.095 ;
        RECT 22.275 -37.445 22.675 -37.095 ;
        RECT 31.235 -37.445 31.635 -37.095 ;
        RECT 40.195 -37.445 40.595 -37.095 ;
        RECT 49.155 -37.445 49.555 -37.095 ;
        RECT 58.115 -37.445 58.515 -37.095 ;
        RECT 67.075 -37.445 67.475 -37.095 ;
        RECT 76.035 -37.445 76.435 -37.095 ;
        RECT 84.995 -37.445 85.395 -37.095 ;
        RECT 93.955 -37.445 94.355 -37.095 ;
        RECT -471.645 -37.495 105.555 -37.445 ;
        RECT -471.645 -37.895 105.955 -37.495 ;
        RECT -471.645 -37.945 105.555 -37.895 ;
        RECT -471.645 -38.295 -471.245 -37.945 ;
        RECT -462.685 -38.295 -462.285 -37.945 ;
        RECT -453.725 -38.295 -453.325 -37.945 ;
        RECT -444.765 -38.295 -444.365 -37.945 ;
        RECT -435.805 -38.295 -435.405 -37.945 ;
        RECT -426.845 -38.295 -426.445 -37.945 ;
        RECT -417.885 -38.295 -417.485 -37.945 ;
        RECT -408.925 -38.295 -408.525 -37.945 ;
        RECT -399.965 -38.295 -399.565 -37.945 ;
        RECT -391.005 -38.295 -390.605 -37.945 ;
        RECT -382.045 -38.295 -381.645 -37.945 ;
        RECT -373.085 -38.295 -372.685 -37.945 ;
        RECT -364.125 -38.295 -363.725 -37.945 ;
        RECT -355.165 -38.295 -354.765 -37.945 ;
        RECT -346.205 -38.295 -345.805 -37.945 ;
        RECT -337.245 -38.295 -336.845 -37.945 ;
        RECT -328.285 -38.295 -327.885 -37.945 ;
        RECT -319.325 -38.295 -318.925 -37.945 ;
        RECT -310.365 -38.295 -309.965 -37.945 ;
        RECT -301.405 -38.295 -301.005 -37.945 ;
        RECT -292.445 -38.295 -292.045 -37.945 ;
        RECT -283.485 -38.295 -283.085 -37.945 ;
        RECT -274.525 -38.295 -274.125 -37.945 ;
        RECT -265.565 -38.295 -265.165 -37.945 ;
        RECT -256.605 -38.295 -256.205 -37.945 ;
        RECT -247.645 -38.295 -247.245 -37.945 ;
        RECT -238.685 -38.295 -238.285 -37.945 ;
        RECT -229.725 -38.295 -229.325 -37.945 ;
        RECT -220.765 -38.295 -220.365 -37.945 ;
        RECT -211.805 -38.295 -211.405 -37.945 ;
        RECT -202.845 -38.295 -202.445 -37.945 ;
        RECT -193.885 -38.295 -193.485 -37.945 ;
        RECT -183.805 -38.295 -183.405 -37.945 ;
        RECT -174.845 -38.295 -174.445 -37.945 ;
        RECT -165.885 -38.295 -165.485 -37.945 ;
        RECT -156.925 -38.295 -156.525 -37.945 ;
        RECT -147.965 -38.295 -147.565 -37.945 ;
        RECT -139.005 -38.295 -138.605 -37.945 ;
        RECT -130.045 -38.295 -129.645 -37.945 ;
        RECT -121.085 -38.295 -120.685 -37.945 ;
        RECT -112.125 -38.295 -111.725 -37.945 ;
        RECT -103.165 -38.295 -102.765 -37.945 ;
        RECT -94.205 -38.295 -93.805 -37.945 ;
        RECT -85.245 -38.295 -84.845 -37.945 ;
        RECT -76.285 -38.295 -75.885 -37.945 ;
        RECT -67.325 -38.295 -66.925 -37.945 ;
        RECT -58.365 -38.295 -57.965 -37.945 ;
        RECT -49.405 -38.295 -49.005 -37.945 ;
        RECT -40.445 -38.295 -40.045 -37.945 ;
        RECT -31.485 -38.295 -31.085 -37.945 ;
        RECT -22.525 -38.295 -22.125 -37.945 ;
        RECT -13.565 -38.295 -13.165 -37.945 ;
        RECT -4.605 -38.295 -4.205 -37.945 ;
        RECT 4.355 -38.295 4.755 -37.945 ;
        RECT 13.315 -38.295 13.715 -37.945 ;
        RECT 22.275 -38.295 22.675 -37.945 ;
        RECT 31.235 -38.295 31.635 -37.945 ;
        RECT 40.195 -38.295 40.595 -37.945 ;
        RECT 49.155 -38.295 49.555 -37.945 ;
        RECT 58.115 -38.295 58.515 -37.945 ;
        RECT 67.075 -38.295 67.475 -37.945 ;
        RECT 76.035 -38.295 76.435 -37.945 ;
        RECT 84.995 -38.295 85.395 -37.945 ;
        RECT 93.955 -38.295 94.355 -37.945 ;
        RECT -473.885 -40.805 -473.485 -40.455 ;
        RECT -469.405 -40.805 -469.005 -40.455 ;
        RECT -464.925 -40.805 -464.525 -40.455 ;
        RECT -460.445 -40.805 -460.045 -40.455 ;
        RECT -455.965 -40.805 -455.565 -40.455 ;
        RECT -451.485 -40.805 -451.085 -40.455 ;
        RECT -447.005 -40.805 -446.605 -40.455 ;
        RECT -442.525 -40.805 -442.125 -40.455 ;
        RECT -438.045 -40.805 -437.645 -40.455 ;
        RECT -433.565 -40.805 -433.165 -40.455 ;
        RECT -429.085 -40.805 -428.685 -40.455 ;
        RECT -424.605 -40.805 -424.205 -40.455 ;
        RECT -420.125 -40.805 -419.725 -40.455 ;
        RECT -415.645 -40.805 -415.245 -40.455 ;
        RECT -411.165 -40.805 -410.765 -40.455 ;
        RECT -406.685 -40.805 -406.285 -40.455 ;
        RECT -402.205 -40.805 -401.805 -40.455 ;
        RECT -397.725 -40.805 -397.325 -40.455 ;
        RECT -393.245 -40.805 -392.845 -40.455 ;
        RECT -388.765 -40.805 -388.365 -40.455 ;
        RECT -384.285 -40.805 -383.885 -40.455 ;
        RECT -379.805 -40.805 -379.405 -40.455 ;
        RECT -375.325 -40.805 -374.925 -40.455 ;
        RECT -370.845 -40.805 -370.445 -40.455 ;
        RECT -366.365 -40.805 -365.965 -40.455 ;
        RECT -361.885 -40.805 -361.485 -40.455 ;
        RECT -357.405 -40.805 -357.005 -40.455 ;
        RECT -352.925 -40.805 -352.525 -40.455 ;
        RECT -348.445 -40.805 -348.045 -40.455 ;
        RECT -343.965 -40.805 -343.565 -40.455 ;
        RECT -339.485 -40.805 -339.085 -40.455 ;
        RECT -335.005 -40.805 -334.605 -40.455 ;
        RECT -330.525 -40.805 -330.125 -40.455 ;
        RECT -326.045 -40.805 -325.645 -40.455 ;
        RECT -321.565 -40.805 -321.165 -40.455 ;
        RECT -317.085 -40.805 -316.685 -40.455 ;
        RECT -312.605 -40.805 -312.205 -40.455 ;
        RECT -308.125 -40.805 -307.725 -40.455 ;
        RECT -303.645 -40.805 -303.245 -40.455 ;
        RECT -299.165 -40.805 -298.765 -40.455 ;
        RECT -294.685 -40.805 -294.285 -40.455 ;
        RECT -290.205 -40.805 -289.805 -40.455 ;
        RECT -285.725 -40.805 -285.325 -40.455 ;
        RECT -281.245 -40.805 -280.845 -40.455 ;
        RECT -276.765 -40.805 -276.365 -40.455 ;
        RECT -272.285 -40.805 -271.885 -40.455 ;
        RECT -267.805 -40.805 -267.405 -40.455 ;
        RECT -263.325 -40.805 -262.925 -40.455 ;
        RECT -258.845 -40.805 -258.445 -40.455 ;
        RECT -254.365 -40.805 -253.965 -40.455 ;
        RECT -249.885 -40.805 -249.485 -40.455 ;
        RECT -245.405 -40.805 -245.005 -40.455 ;
        RECT -240.925 -40.805 -240.525 -40.455 ;
        RECT -236.445 -40.805 -236.045 -40.455 ;
        RECT -231.965 -40.805 -231.565 -40.455 ;
        RECT -227.485 -40.805 -227.085 -40.455 ;
        RECT -223.005 -40.805 -222.605 -40.455 ;
        RECT -218.525 -40.805 -218.125 -40.455 ;
        RECT -214.045 -40.805 -213.645 -40.455 ;
        RECT -209.565 -40.805 -209.165 -40.455 ;
        RECT -205.085 -40.805 -204.685 -40.455 ;
        RECT -200.605 -40.805 -200.205 -40.455 ;
        RECT -196.125 -40.805 -195.725 -40.455 ;
        RECT -191.645 -40.805 -191.245 -40.455 ;
        RECT -186.045 -40.805 -185.645 -40.455 ;
        RECT -181.565 -40.805 -181.165 -40.455 ;
        RECT -177.085 -40.805 -176.685 -40.455 ;
        RECT -172.605 -40.805 -172.205 -40.455 ;
        RECT -168.125 -40.805 -167.725 -40.455 ;
        RECT -163.645 -40.805 -163.245 -40.455 ;
        RECT -159.165 -40.805 -158.765 -40.455 ;
        RECT -154.685 -40.805 -154.285 -40.455 ;
        RECT -150.205 -40.805 -149.805 -40.455 ;
        RECT -145.725 -40.805 -145.325 -40.455 ;
        RECT -141.245 -40.805 -140.845 -40.455 ;
        RECT -136.765 -40.805 -136.365 -40.455 ;
        RECT -132.285 -40.805 -131.885 -40.455 ;
        RECT -127.805 -40.805 -127.405 -40.455 ;
        RECT -123.325 -40.805 -122.925 -40.455 ;
        RECT -118.845 -40.805 -118.445 -40.455 ;
        RECT -114.365 -40.805 -113.965 -40.455 ;
        RECT -109.885 -40.805 -109.485 -40.455 ;
        RECT -105.405 -40.805 -105.005 -40.455 ;
        RECT -100.925 -40.805 -100.525 -40.455 ;
        RECT -96.445 -40.805 -96.045 -40.455 ;
        RECT -91.965 -40.805 -91.565 -40.455 ;
        RECT -87.485 -40.805 -87.085 -40.455 ;
        RECT -83.005 -40.805 -82.605 -40.455 ;
        RECT -78.525 -40.805 -78.125 -40.455 ;
        RECT -74.045 -40.805 -73.645 -40.455 ;
        RECT -69.565 -40.805 -69.165 -40.455 ;
        RECT -65.085 -40.805 -64.685 -40.455 ;
        RECT -60.605 -40.805 -60.205 -40.455 ;
        RECT -56.125 -40.805 -55.725 -40.455 ;
        RECT -51.645 -40.805 -51.245 -40.455 ;
        RECT -47.165 -40.805 -46.765 -40.455 ;
        RECT -42.685 -40.805 -42.285 -40.455 ;
        RECT -38.205 -40.805 -37.805 -40.455 ;
        RECT -33.725 -40.805 -33.325 -40.455 ;
        RECT -29.245 -40.805 -28.845 -40.455 ;
        RECT -24.765 -40.805 -24.365 -40.455 ;
        RECT -20.285 -40.805 -19.885 -40.455 ;
        RECT -15.805 -40.805 -15.405 -40.455 ;
        RECT -11.325 -40.805 -10.925 -40.455 ;
        RECT -6.845 -40.805 -6.445 -40.455 ;
        RECT -2.365 -40.805 -1.965 -40.455 ;
        RECT 2.115 -40.805 2.515 -40.455 ;
        RECT 6.595 -40.805 6.995 -40.455 ;
        RECT 11.075 -40.805 11.475 -40.455 ;
        RECT 15.555 -40.805 15.955 -40.455 ;
        RECT 20.035 -40.805 20.435 -40.455 ;
        RECT 24.515 -40.805 24.915 -40.455 ;
        RECT 28.995 -40.805 29.395 -40.455 ;
        RECT 33.475 -40.805 33.875 -40.455 ;
        RECT 37.955 -40.805 38.355 -40.455 ;
        RECT 42.435 -40.805 42.835 -40.455 ;
        RECT 46.915 -40.805 47.315 -40.455 ;
        RECT 51.395 -40.805 51.795 -40.455 ;
        RECT 55.875 -40.805 56.275 -40.455 ;
        RECT 60.355 -40.805 60.755 -40.455 ;
        RECT 64.835 -40.805 65.235 -40.455 ;
        RECT 69.315 -40.805 69.715 -40.455 ;
        RECT 73.795 -40.805 74.195 -40.455 ;
        RECT 78.275 -40.805 78.675 -40.455 ;
        RECT 82.755 -40.805 83.155 -40.455 ;
        RECT 87.235 -40.805 87.635 -40.455 ;
        RECT 91.715 -40.805 92.115 -40.455 ;
        RECT 96.195 -40.805 96.595 -40.455 ;
        RECT -473.885 -40.855 103.755 -40.805 ;
        RECT -473.885 -41.255 104.155 -40.855 ;
        RECT -473.885 -41.305 103.755 -41.255 ;
        RECT -473.885 -41.655 -473.485 -41.305 ;
        RECT -469.405 -41.655 -469.005 -41.305 ;
        RECT -464.925 -41.655 -464.525 -41.305 ;
        RECT -460.445 -41.655 -460.045 -41.305 ;
        RECT -455.965 -41.655 -455.565 -41.305 ;
        RECT -451.485 -41.655 -451.085 -41.305 ;
        RECT -447.005 -41.655 -446.605 -41.305 ;
        RECT -442.525 -41.655 -442.125 -41.305 ;
        RECT -438.045 -41.655 -437.645 -41.305 ;
        RECT -433.565 -41.655 -433.165 -41.305 ;
        RECT -429.085 -41.655 -428.685 -41.305 ;
        RECT -424.605 -41.655 -424.205 -41.305 ;
        RECT -420.125 -41.655 -419.725 -41.305 ;
        RECT -415.645 -41.655 -415.245 -41.305 ;
        RECT -411.165 -41.655 -410.765 -41.305 ;
        RECT -406.685 -41.655 -406.285 -41.305 ;
        RECT -402.205 -41.655 -401.805 -41.305 ;
        RECT -397.725 -41.655 -397.325 -41.305 ;
        RECT -393.245 -41.655 -392.845 -41.305 ;
        RECT -388.765 -41.655 -388.365 -41.305 ;
        RECT -384.285 -41.655 -383.885 -41.305 ;
        RECT -379.805 -41.655 -379.405 -41.305 ;
        RECT -375.325 -41.655 -374.925 -41.305 ;
        RECT -370.845 -41.655 -370.445 -41.305 ;
        RECT -366.365 -41.655 -365.965 -41.305 ;
        RECT -361.885 -41.655 -361.485 -41.305 ;
        RECT -357.405 -41.655 -357.005 -41.305 ;
        RECT -352.925 -41.655 -352.525 -41.305 ;
        RECT -348.445 -41.655 -348.045 -41.305 ;
        RECT -343.965 -41.655 -343.565 -41.305 ;
        RECT -339.485 -41.655 -339.085 -41.305 ;
        RECT -335.005 -41.655 -334.605 -41.305 ;
        RECT -330.525 -41.655 -330.125 -41.305 ;
        RECT -326.045 -41.655 -325.645 -41.305 ;
        RECT -321.565 -41.655 -321.165 -41.305 ;
        RECT -317.085 -41.655 -316.685 -41.305 ;
        RECT -312.605 -41.655 -312.205 -41.305 ;
        RECT -308.125 -41.655 -307.725 -41.305 ;
        RECT -303.645 -41.655 -303.245 -41.305 ;
        RECT -299.165 -41.655 -298.765 -41.305 ;
        RECT -294.685 -41.655 -294.285 -41.305 ;
        RECT -290.205 -41.655 -289.805 -41.305 ;
        RECT -285.725 -41.655 -285.325 -41.305 ;
        RECT -281.245 -41.655 -280.845 -41.305 ;
        RECT -276.765 -41.655 -276.365 -41.305 ;
        RECT -272.285 -41.655 -271.885 -41.305 ;
        RECT -267.805 -41.655 -267.405 -41.305 ;
        RECT -263.325 -41.655 -262.925 -41.305 ;
        RECT -258.845 -41.655 -258.445 -41.305 ;
        RECT -254.365 -41.655 -253.965 -41.305 ;
        RECT -249.885 -41.655 -249.485 -41.305 ;
        RECT -245.405 -41.655 -245.005 -41.305 ;
        RECT -240.925 -41.655 -240.525 -41.305 ;
        RECT -236.445 -41.655 -236.045 -41.305 ;
        RECT -231.965 -41.655 -231.565 -41.305 ;
        RECT -227.485 -41.655 -227.085 -41.305 ;
        RECT -223.005 -41.655 -222.605 -41.305 ;
        RECT -218.525 -41.655 -218.125 -41.305 ;
        RECT -214.045 -41.655 -213.645 -41.305 ;
        RECT -209.565 -41.655 -209.165 -41.305 ;
        RECT -205.085 -41.655 -204.685 -41.305 ;
        RECT -200.605 -41.655 -200.205 -41.305 ;
        RECT -196.125 -41.655 -195.725 -41.305 ;
        RECT -191.645 -41.655 -191.245 -41.305 ;
        RECT -186.045 -41.655 -185.645 -41.305 ;
        RECT -181.565 -41.655 -181.165 -41.305 ;
        RECT -177.085 -41.655 -176.685 -41.305 ;
        RECT -172.605 -41.655 -172.205 -41.305 ;
        RECT -168.125 -41.655 -167.725 -41.305 ;
        RECT -163.645 -41.655 -163.245 -41.305 ;
        RECT -159.165 -41.655 -158.765 -41.305 ;
        RECT -154.685 -41.655 -154.285 -41.305 ;
        RECT -150.205 -41.655 -149.805 -41.305 ;
        RECT -145.725 -41.655 -145.325 -41.305 ;
        RECT -141.245 -41.655 -140.845 -41.305 ;
        RECT -136.765 -41.655 -136.365 -41.305 ;
        RECT -132.285 -41.655 -131.885 -41.305 ;
        RECT -127.805 -41.655 -127.405 -41.305 ;
        RECT -123.325 -41.655 -122.925 -41.305 ;
        RECT -118.845 -41.655 -118.445 -41.305 ;
        RECT -114.365 -41.655 -113.965 -41.305 ;
        RECT -109.885 -41.655 -109.485 -41.305 ;
        RECT -105.405 -41.655 -105.005 -41.305 ;
        RECT -100.925 -41.655 -100.525 -41.305 ;
        RECT -96.445 -41.655 -96.045 -41.305 ;
        RECT -91.965 -41.655 -91.565 -41.305 ;
        RECT -87.485 -41.655 -87.085 -41.305 ;
        RECT -83.005 -41.655 -82.605 -41.305 ;
        RECT -78.525 -41.655 -78.125 -41.305 ;
        RECT -74.045 -41.655 -73.645 -41.305 ;
        RECT -69.565 -41.655 -69.165 -41.305 ;
        RECT -65.085 -41.655 -64.685 -41.305 ;
        RECT -60.605 -41.655 -60.205 -41.305 ;
        RECT -56.125 -41.655 -55.725 -41.305 ;
        RECT -51.645 -41.655 -51.245 -41.305 ;
        RECT -47.165 -41.655 -46.765 -41.305 ;
        RECT -42.685 -41.655 -42.285 -41.305 ;
        RECT -38.205 -41.655 -37.805 -41.305 ;
        RECT -33.725 -41.655 -33.325 -41.305 ;
        RECT -29.245 -41.655 -28.845 -41.305 ;
        RECT -24.765 -41.655 -24.365 -41.305 ;
        RECT -20.285 -41.655 -19.885 -41.305 ;
        RECT -15.805 -41.655 -15.405 -41.305 ;
        RECT -11.325 -41.655 -10.925 -41.305 ;
        RECT -6.845 -41.655 -6.445 -41.305 ;
        RECT -2.365 -41.655 -1.965 -41.305 ;
        RECT 2.115 -41.655 2.515 -41.305 ;
        RECT 6.595 -41.655 6.995 -41.305 ;
        RECT 11.075 -41.655 11.475 -41.305 ;
        RECT 15.555 -41.655 15.955 -41.305 ;
        RECT 20.035 -41.655 20.435 -41.305 ;
        RECT 24.515 -41.655 24.915 -41.305 ;
        RECT 28.995 -41.655 29.395 -41.305 ;
        RECT 33.475 -41.655 33.875 -41.305 ;
        RECT 37.955 -41.655 38.355 -41.305 ;
        RECT 42.435 -41.655 42.835 -41.305 ;
        RECT 46.915 -41.655 47.315 -41.305 ;
        RECT 51.395 -41.655 51.795 -41.305 ;
        RECT 55.875 -41.655 56.275 -41.305 ;
        RECT 60.355 -41.655 60.755 -41.305 ;
        RECT 64.835 -41.655 65.235 -41.305 ;
        RECT 69.315 -41.655 69.715 -41.305 ;
        RECT 73.795 -41.655 74.195 -41.305 ;
        RECT 78.275 -41.655 78.675 -41.305 ;
        RECT 82.755 -41.655 83.155 -41.305 ;
        RECT 87.235 -41.655 87.635 -41.305 ;
        RECT 91.715 -41.655 92.115 -41.305 ;
        RECT 96.195 -41.655 96.595 -41.305 ;
        RECT -497.305 -42.900 -486.905 -42.300 ;
        RECT -475.005 -44.165 -474.605 -43.815 ;
        RECT -472.765 -44.165 -472.365 -43.815 ;
        RECT -470.525 -44.165 -470.125 -43.815 ;
        RECT -468.285 -44.165 -467.885 -43.815 ;
        RECT -466.045 -44.165 -465.645 -43.815 ;
        RECT -463.805 -44.165 -463.405 -43.815 ;
        RECT -461.565 -44.165 -461.165 -43.815 ;
        RECT -459.325 -44.165 -458.925 -43.815 ;
        RECT -457.085 -44.165 -456.685 -43.815 ;
        RECT -454.845 -44.165 -454.445 -43.815 ;
        RECT -452.605 -44.165 -452.205 -43.815 ;
        RECT -450.365 -44.165 -449.965 -43.815 ;
        RECT -448.125 -44.165 -447.725 -43.815 ;
        RECT -445.885 -44.165 -445.485 -43.815 ;
        RECT -443.645 -44.165 -443.245 -43.815 ;
        RECT -441.405 -44.165 -441.005 -43.815 ;
        RECT -439.165 -44.165 -438.765 -43.815 ;
        RECT -436.925 -44.165 -436.525 -43.815 ;
        RECT -434.685 -44.165 -434.285 -43.815 ;
        RECT -432.445 -44.165 -432.045 -43.815 ;
        RECT -430.205 -44.165 -429.805 -43.815 ;
        RECT -427.965 -44.165 -427.565 -43.815 ;
        RECT -425.725 -44.165 -425.325 -43.815 ;
        RECT -423.485 -44.165 -423.085 -43.815 ;
        RECT -421.245 -44.165 -420.845 -43.815 ;
        RECT -419.005 -44.165 -418.605 -43.815 ;
        RECT -416.765 -44.165 -416.365 -43.815 ;
        RECT -414.525 -44.165 -414.125 -43.815 ;
        RECT -412.285 -44.165 -411.885 -43.815 ;
        RECT -410.045 -44.165 -409.645 -43.815 ;
        RECT -407.805 -44.165 -407.405 -43.815 ;
        RECT -405.565 -44.165 -405.165 -43.815 ;
        RECT -403.325 -44.165 -402.925 -43.815 ;
        RECT -401.085 -44.165 -400.685 -43.815 ;
        RECT -398.845 -44.165 -398.445 -43.815 ;
        RECT -396.605 -44.165 -396.205 -43.815 ;
        RECT -394.365 -44.165 -393.965 -43.815 ;
        RECT -392.125 -44.165 -391.725 -43.815 ;
        RECT -389.885 -44.165 -389.485 -43.815 ;
        RECT -387.645 -44.165 -387.245 -43.815 ;
        RECT -385.405 -44.165 -385.005 -43.815 ;
        RECT -383.165 -44.165 -382.765 -43.815 ;
        RECT -380.925 -44.165 -380.525 -43.815 ;
        RECT -378.685 -44.165 -378.285 -43.815 ;
        RECT -376.445 -44.165 -376.045 -43.815 ;
        RECT -374.205 -44.165 -373.805 -43.815 ;
        RECT -371.965 -44.165 -371.565 -43.815 ;
        RECT -369.725 -44.165 -369.325 -43.815 ;
        RECT -367.485 -44.165 -367.085 -43.815 ;
        RECT -365.245 -44.165 -364.845 -43.815 ;
        RECT -363.005 -44.165 -362.605 -43.815 ;
        RECT -360.765 -44.165 -360.365 -43.815 ;
        RECT -358.525 -44.165 -358.125 -43.815 ;
        RECT -356.285 -44.165 -355.885 -43.815 ;
        RECT -354.045 -44.165 -353.645 -43.815 ;
        RECT -351.805 -44.165 -351.405 -43.815 ;
        RECT -349.565 -44.165 -349.165 -43.815 ;
        RECT -347.325 -44.165 -346.925 -43.815 ;
        RECT -345.085 -44.165 -344.685 -43.815 ;
        RECT -342.845 -44.165 -342.445 -43.815 ;
        RECT -340.605 -44.165 -340.205 -43.815 ;
        RECT -338.365 -44.165 -337.965 -43.815 ;
        RECT -336.125 -44.165 -335.725 -43.815 ;
        RECT -333.885 -44.165 -333.485 -43.815 ;
        RECT -331.645 -44.165 -331.245 -43.815 ;
        RECT -329.405 -44.165 -329.005 -43.815 ;
        RECT -327.165 -44.165 -326.765 -43.815 ;
        RECT -324.925 -44.165 -324.525 -43.815 ;
        RECT -322.685 -44.165 -322.285 -43.815 ;
        RECT -320.445 -44.165 -320.045 -43.815 ;
        RECT -318.205 -44.165 -317.805 -43.815 ;
        RECT -315.965 -44.165 -315.565 -43.815 ;
        RECT -313.725 -44.165 -313.325 -43.815 ;
        RECT -311.485 -44.165 -311.085 -43.815 ;
        RECT -309.245 -44.165 -308.845 -43.815 ;
        RECT -307.005 -44.165 -306.605 -43.815 ;
        RECT -304.765 -44.165 -304.365 -43.815 ;
        RECT -302.525 -44.165 -302.125 -43.815 ;
        RECT -300.285 -44.165 -299.885 -43.815 ;
        RECT -298.045 -44.165 -297.645 -43.815 ;
        RECT -295.805 -44.165 -295.405 -43.815 ;
        RECT -293.565 -44.165 -293.165 -43.815 ;
        RECT -291.325 -44.165 -290.925 -43.815 ;
        RECT -289.085 -44.165 -288.685 -43.815 ;
        RECT -286.845 -44.165 -286.445 -43.815 ;
        RECT -284.605 -44.165 -284.205 -43.815 ;
        RECT -282.365 -44.165 -281.965 -43.815 ;
        RECT -280.125 -44.165 -279.725 -43.815 ;
        RECT -277.885 -44.165 -277.485 -43.815 ;
        RECT -275.645 -44.165 -275.245 -43.815 ;
        RECT -273.405 -44.165 -273.005 -43.815 ;
        RECT -271.165 -44.165 -270.765 -43.815 ;
        RECT -268.925 -44.165 -268.525 -43.815 ;
        RECT -266.685 -44.165 -266.285 -43.815 ;
        RECT -264.445 -44.165 -264.045 -43.815 ;
        RECT -262.205 -44.165 -261.805 -43.815 ;
        RECT -259.965 -44.165 -259.565 -43.815 ;
        RECT -257.725 -44.165 -257.325 -43.815 ;
        RECT -255.485 -44.165 -255.085 -43.815 ;
        RECT -253.245 -44.165 -252.845 -43.815 ;
        RECT -251.005 -44.165 -250.605 -43.815 ;
        RECT -248.765 -44.165 -248.365 -43.815 ;
        RECT -246.525 -44.165 -246.125 -43.815 ;
        RECT -244.285 -44.165 -243.885 -43.815 ;
        RECT -242.045 -44.165 -241.645 -43.815 ;
        RECT -239.805 -44.165 -239.405 -43.815 ;
        RECT -237.565 -44.165 -237.165 -43.815 ;
        RECT -235.325 -44.165 -234.925 -43.815 ;
        RECT -233.085 -44.165 -232.685 -43.815 ;
        RECT -230.845 -44.165 -230.445 -43.815 ;
        RECT -228.605 -44.165 -228.205 -43.815 ;
        RECT -226.365 -44.165 -225.965 -43.815 ;
        RECT -224.125 -44.165 -223.725 -43.815 ;
        RECT -221.885 -44.165 -221.485 -43.815 ;
        RECT -219.645 -44.165 -219.245 -43.815 ;
        RECT -217.405 -44.165 -217.005 -43.815 ;
        RECT -215.165 -44.165 -214.765 -43.815 ;
        RECT -212.925 -44.165 -212.525 -43.815 ;
        RECT -210.685 -44.165 -210.285 -43.815 ;
        RECT -208.445 -44.165 -208.045 -43.815 ;
        RECT -206.205 -44.165 -205.805 -43.815 ;
        RECT -203.965 -44.165 -203.565 -43.815 ;
        RECT -201.725 -44.165 -201.325 -43.815 ;
        RECT -199.485 -44.165 -199.085 -43.815 ;
        RECT -197.245 -44.165 -196.845 -43.815 ;
        RECT -195.005 -44.165 -194.605 -43.815 ;
        RECT -192.765 -44.165 -192.365 -43.815 ;
        RECT -190.525 -44.165 -190.125 -43.815 ;
        RECT -187.165 -44.165 -186.765 -43.815 ;
        RECT -184.925 -44.165 -184.525 -43.815 ;
        RECT -182.685 -44.165 -182.285 -43.815 ;
        RECT -180.445 -44.165 -180.045 -43.815 ;
        RECT -178.205 -44.165 -177.805 -43.815 ;
        RECT -175.965 -44.165 -175.565 -43.815 ;
        RECT -173.725 -44.165 -173.325 -43.815 ;
        RECT -171.485 -44.165 -171.085 -43.815 ;
        RECT -169.245 -44.165 -168.845 -43.815 ;
        RECT -167.005 -44.165 -166.605 -43.815 ;
        RECT -164.765 -44.165 -164.365 -43.815 ;
        RECT -162.525 -44.165 -162.125 -43.815 ;
        RECT -160.285 -44.165 -159.885 -43.815 ;
        RECT -158.045 -44.165 -157.645 -43.815 ;
        RECT -155.805 -44.165 -155.405 -43.815 ;
        RECT -153.565 -44.165 -153.165 -43.815 ;
        RECT -151.325 -44.165 -150.925 -43.815 ;
        RECT -149.085 -44.165 -148.685 -43.815 ;
        RECT -146.845 -44.165 -146.445 -43.815 ;
        RECT -144.605 -44.165 -144.205 -43.815 ;
        RECT -142.365 -44.165 -141.965 -43.815 ;
        RECT -140.125 -44.165 -139.725 -43.815 ;
        RECT -137.885 -44.165 -137.485 -43.815 ;
        RECT -135.645 -44.165 -135.245 -43.815 ;
        RECT -133.405 -44.165 -133.005 -43.815 ;
        RECT -131.165 -44.165 -130.765 -43.815 ;
        RECT -128.925 -44.165 -128.525 -43.815 ;
        RECT -126.685 -44.165 -126.285 -43.815 ;
        RECT -124.445 -44.165 -124.045 -43.815 ;
        RECT -122.205 -44.165 -121.805 -43.815 ;
        RECT -119.965 -44.165 -119.565 -43.815 ;
        RECT -117.725 -44.165 -117.325 -43.815 ;
        RECT -115.485 -44.165 -115.085 -43.815 ;
        RECT -113.245 -44.165 -112.845 -43.815 ;
        RECT -111.005 -44.165 -110.605 -43.815 ;
        RECT -108.765 -44.165 -108.365 -43.815 ;
        RECT -106.525 -44.165 -106.125 -43.815 ;
        RECT -104.285 -44.165 -103.885 -43.815 ;
        RECT -102.045 -44.165 -101.645 -43.815 ;
        RECT -99.805 -44.165 -99.405 -43.815 ;
        RECT -97.565 -44.165 -97.165 -43.815 ;
        RECT -95.325 -44.165 -94.925 -43.815 ;
        RECT -93.085 -44.165 -92.685 -43.815 ;
        RECT -90.845 -44.165 -90.445 -43.815 ;
        RECT -88.605 -44.165 -88.205 -43.815 ;
        RECT -86.365 -44.165 -85.965 -43.815 ;
        RECT -84.125 -44.165 -83.725 -43.815 ;
        RECT -81.885 -44.165 -81.485 -43.815 ;
        RECT -79.645 -44.165 -79.245 -43.815 ;
        RECT -77.405 -44.165 -77.005 -43.815 ;
        RECT -75.165 -44.165 -74.765 -43.815 ;
        RECT -72.925 -44.165 -72.525 -43.815 ;
        RECT -70.685 -44.165 -70.285 -43.815 ;
        RECT -68.445 -44.165 -68.045 -43.815 ;
        RECT -66.205 -44.165 -65.805 -43.815 ;
        RECT -63.965 -44.165 -63.565 -43.815 ;
        RECT -61.725 -44.165 -61.325 -43.815 ;
        RECT -59.485 -44.165 -59.085 -43.815 ;
        RECT -57.245 -44.165 -56.845 -43.815 ;
        RECT -55.005 -44.165 -54.605 -43.815 ;
        RECT -52.765 -44.165 -52.365 -43.815 ;
        RECT -50.525 -44.165 -50.125 -43.815 ;
        RECT -48.285 -44.165 -47.885 -43.815 ;
        RECT -46.045 -44.165 -45.645 -43.815 ;
        RECT -43.805 -44.165 -43.405 -43.815 ;
        RECT -41.565 -44.165 -41.165 -43.815 ;
        RECT -39.325 -44.165 -38.925 -43.815 ;
        RECT -37.085 -44.165 -36.685 -43.815 ;
        RECT -34.845 -44.165 -34.445 -43.815 ;
        RECT -32.605 -44.165 -32.205 -43.815 ;
        RECT -30.365 -44.165 -29.965 -43.815 ;
        RECT -28.125 -44.165 -27.725 -43.815 ;
        RECT -25.885 -44.165 -25.485 -43.815 ;
        RECT -23.645 -44.165 -23.245 -43.815 ;
        RECT -21.405 -44.165 -21.005 -43.815 ;
        RECT -19.165 -44.165 -18.765 -43.815 ;
        RECT -16.925 -44.165 -16.525 -43.815 ;
        RECT -14.685 -44.165 -14.285 -43.815 ;
        RECT -12.445 -44.165 -12.045 -43.815 ;
        RECT -10.205 -44.165 -9.805 -43.815 ;
        RECT -7.965 -44.165 -7.565 -43.815 ;
        RECT -5.725 -44.165 -5.325 -43.815 ;
        RECT -3.485 -44.165 -3.085 -43.815 ;
        RECT -1.245 -44.165 -0.845 -43.815 ;
        RECT 0.995 -44.165 1.395 -43.815 ;
        RECT 3.235 -44.165 3.635 -43.815 ;
        RECT 5.475 -44.165 5.875 -43.815 ;
        RECT 7.715 -44.165 8.115 -43.815 ;
        RECT 9.955 -44.165 10.355 -43.815 ;
        RECT 12.195 -44.165 12.595 -43.815 ;
        RECT 14.435 -44.165 14.835 -43.815 ;
        RECT 16.675 -44.165 17.075 -43.815 ;
        RECT 18.915 -44.165 19.315 -43.815 ;
        RECT 21.155 -44.165 21.555 -43.815 ;
        RECT 23.395 -44.165 23.795 -43.815 ;
        RECT 25.635 -44.165 26.035 -43.815 ;
        RECT 27.875 -44.165 28.275 -43.815 ;
        RECT 30.115 -44.165 30.515 -43.815 ;
        RECT 32.355 -44.165 32.755 -43.815 ;
        RECT 34.595 -44.165 34.995 -43.815 ;
        RECT 36.835 -44.165 37.235 -43.815 ;
        RECT 39.075 -44.165 39.475 -43.815 ;
        RECT 41.315 -44.165 41.715 -43.815 ;
        RECT 43.555 -44.165 43.955 -43.815 ;
        RECT 45.795 -44.165 46.195 -43.815 ;
        RECT 48.035 -44.165 48.435 -43.815 ;
        RECT 50.275 -44.165 50.675 -43.815 ;
        RECT 52.515 -44.165 52.915 -43.815 ;
        RECT 54.755 -44.165 55.155 -43.815 ;
        RECT 56.995 -44.165 57.395 -43.815 ;
        RECT 59.235 -44.165 59.635 -43.815 ;
        RECT 61.475 -44.165 61.875 -43.815 ;
        RECT 63.715 -44.165 64.115 -43.815 ;
        RECT 65.955 -44.165 66.355 -43.815 ;
        RECT 68.195 -44.165 68.595 -43.815 ;
        RECT 70.435 -44.165 70.835 -43.815 ;
        RECT 72.675 -44.165 73.075 -43.815 ;
        RECT 74.915 -44.165 75.315 -43.815 ;
        RECT 77.155 -44.165 77.555 -43.815 ;
        RECT 79.395 -44.165 79.795 -43.815 ;
        RECT 81.635 -44.165 82.035 -43.815 ;
        RECT 83.875 -44.165 84.275 -43.815 ;
        RECT 86.115 -44.165 86.515 -43.815 ;
        RECT 88.355 -44.165 88.755 -43.815 ;
        RECT 90.595 -44.165 90.995 -43.815 ;
        RECT 92.835 -44.165 93.235 -43.815 ;
        RECT 95.075 -44.165 95.475 -43.815 ;
        RECT 97.315 -44.165 97.715 -43.815 ;
        RECT -475.005 -44.215 101.955 -44.165 ;
        RECT -475.005 -44.615 102.355 -44.215 ;
        RECT -475.005 -44.665 101.955 -44.615 ;
        RECT -475.005 -45.015 -474.605 -44.665 ;
        RECT -472.765 -45.015 -472.365 -44.665 ;
        RECT -470.525 -45.015 -470.125 -44.665 ;
        RECT -468.285 -45.015 -467.885 -44.665 ;
        RECT -466.045 -45.015 -465.645 -44.665 ;
        RECT -463.805 -45.015 -463.405 -44.665 ;
        RECT -461.565 -45.015 -461.165 -44.665 ;
        RECT -459.325 -45.015 -458.925 -44.665 ;
        RECT -457.085 -45.015 -456.685 -44.665 ;
        RECT -454.845 -45.015 -454.445 -44.665 ;
        RECT -452.605 -45.015 -452.205 -44.665 ;
        RECT -450.365 -45.015 -449.965 -44.665 ;
        RECT -448.125 -45.015 -447.725 -44.665 ;
        RECT -445.885 -45.015 -445.485 -44.665 ;
        RECT -443.645 -45.015 -443.245 -44.665 ;
        RECT -441.405 -45.015 -441.005 -44.665 ;
        RECT -439.165 -45.015 -438.765 -44.665 ;
        RECT -436.925 -45.015 -436.525 -44.665 ;
        RECT -434.685 -45.015 -434.285 -44.665 ;
        RECT -432.445 -45.015 -432.045 -44.665 ;
        RECT -430.205 -45.015 -429.805 -44.665 ;
        RECT -427.965 -45.015 -427.565 -44.665 ;
        RECT -425.725 -45.015 -425.325 -44.665 ;
        RECT -423.485 -45.015 -423.085 -44.665 ;
        RECT -421.245 -45.015 -420.845 -44.665 ;
        RECT -419.005 -45.015 -418.605 -44.665 ;
        RECT -416.765 -45.015 -416.365 -44.665 ;
        RECT -414.525 -45.015 -414.125 -44.665 ;
        RECT -412.285 -45.015 -411.885 -44.665 ;
        RECT -410.045 -45.015 -409.645 -44.665 ;
        RECT -407.805 -45.015 -407.405 -44.665 ;
        RECT -405.565 -45.015 -405.165 -44.665 ;
        RECT -403.325 -45.015 -402.925 -44.665 ;
        RECT -401.085 -45.015 -400.685 -44.665 ;
        RECT -398.845 -45.015 -398.445 -44.665 ;
        RECT -396.605 -45.015 -396.205 -44.665 ;
        RECT -394.365 -45.015 -393.965 -44.665 ;
        RECT -392.125 -45.015 -391.725 -44.665 ;
        RECT -389.885 -45.015 -389.485 -44.665 ;
        RECT -387.645 -45.015 -387.245 -44.665 ;
        RECT -385.405 -45.015 -385.005 -44.665 ;
        RECT -383.165 -45.015 -382.765 -44.665 ;
        RECT -380.925 -45.015 -380.525 -44.665 ;
        RECT -378.685 -45.015 -378.285 -44.665 ;
        RECT -376.445 -45.015 -376.045 -44.665 ;
        RECT -374.205 -45.015 -373.805 -44.665 ;
        RECT -371.965 -45.015 -371.565 -44.665 ;
        RECT -369.725 -45.015 -369.325 -44.665 ;
        RECT -367.485 -45.015 -367.085 -44.665 ;
        RECT -365.245 -45.015 -364.845 -44.665 ;
        RECT -363.005 -45.015 -362.605 -44.665 ;
        RECT -360.765 -45.015 -360.365 -44.665 ;
        RECT -358.525 -45.015 -358.125 -44.665 ;
        RECT -356.285 -45.015 -355.885 -44.665 ;
        RECT -354.045 -45.015 -353.645 -44.665 ;
        RECT -351.805 -45.015 -351.405 -44.665 ;
        RECT -349.565 -45.015 -349.165 -44.665 ;
        RECT -347.325 -45.015 -346.925 -44.665 ;
        RECT -345.085 -45.015 -344.685 -44.665 ;
        RECT -342.845 -45.015 -342.445 -44.665 ;
        RECT -340.605 -45.015 -340.205 -44.665 ;
        RECT -338.365 -45.015 -337.965 -44.665 ;
        RECT -336.125 -45.015 -335.725 -44.665 ;
        RECT -333.885 -45.015 -333.485 -44.665 ;
        RECT -331.645 -45.015 -331.245 -44.665 ;
        RECT -329.405 -45.015 -329.005 -44.665 ;
        RECT -327.165 -45.015 -326.765 -44.665 ;
        RECT -324.925 -45.015 -324.525 -44.665 ;
        RECT -322.685 -45.015 -322.285 -44.665 ;
        RECT -320.445 -45.015 -320.045 -44.665 ;
        RECT -318.205 -45.015 -317.805 -44.665 ;
        RECT -315.965 -45.015 -315.565 -44.665 ;
        RECT -313.725 -45.015 -313.325 -44.665 ;
        RECT -311.485 -45.015 -311.085 -44.665 ;
        RECT -309.245 -45.015 -308.845 -44.665 ;
        RECT -307.005 -45.015 -306.605 -44.665 ;
        RECT -304.765 -45.015 -304.365 -44.665 ;
        RECT -302.525 -45.015 -302.125 -44.665 ;
        RECT -300.285 -45.015 -299.885 -44.665 ;
        RECT -298.045 -45.015 -297.645 -44.665 ;
        RECT -295.805 -45.015 -295.405 -44.665 ;
        RECT -293.565 -45.015 -293.165 -44.665 ;
        RECT -291.325 -45.015 -290.925 -44.665 ;
        RECT -289.085 -45.015 -288.685 -44.665 ;
        RECT -286.845 -45.015 -286.445 -44.665 ;
        RECT -284.605 -45.015 -284.205 -44.665 ;
        RECT -282.365 -45.015 -281.965 -44.665 ;
        RECT -280.125 -45.015 -279.725 -44.665 ;
        RECT -277.885 -45.015 -277.485 -44.665 ;
        RECT -275.645 -45.015 -275.245 -44.665 ;
        RECT -273.405 -45.015 -273.005 -44.665 ;
        RECT -271.165 -45.015 -270.765 -44.665 ;
        RECT -268.925 -45.015 -268.525 -44.665 ;
        RECT -266.685 -45.015 -266.285 -44.665 ;
        RECT -264.445 -45.015 -264.045 -44.665 ;
        RECT -262.205 -45.015 -261.805 -44.665 ;
        RECT -259.965 -45.015 -259.565 -44.665 ;
        RECT -257.725 -45.015 -257.325 -44.665 ;
        RECT -255.485 -45.015 -255.085 -44.665 ;
        RECT -253.245 -45.015 -252.845 -44.665 ;
        RECT -251.005 -45.015 -250.605 -44.665 ;
        RECT -248.765 -45.015 -248.365 -44.665 ;
        RECT -246.525 -45.015 -246.125 -44.665 ;
        RECT -244.285 -45.015 -243.885 -44.665 ;
        RECT -242.045 -45.015 -241.645 -44.665 ;
        RECT -239.805 -45.015 -239.405 -44.665 ;
        RECT -237.565 -45.015 -237.165 -44.665 ;
        RECT -235.325 -45.015 -234.925 -44.665 ;
        RECT -233.085 -45.015 -232.685 -44.665 ;
        RECT -230.845 -45.015 -230.445 -44.665 ;
        RECT -228.605 -45.015 -228.205 -44.665 ;
        RECT -226.365 -45.015 -225.965 -44.665 ;
        RECT -224.125 -45.015 -223.725 -44.665 ;
        RECT -221.885 -45.015 -221.485 -44.665 ;
        RECT -219.645 -45.015 -219.245 -44.665 ;
        RECT -217.405 -45.015 -217.005 -44.665 ;
        RECT -215.165 -45.015 -214.765 -44.665 ;
        RECT -212.925 -45.015 -212.525 -44.665 ;
        RECT -210.685 -45.015 -210.285 -44.665 ;
        RECT -208.445 -45.015 -208.045 -44.665 ;
        RECT -206.205 -45.015 -205.805 -44.665 ;
        RECT -203.965 -45.015 -203.565 -44.665 ;
        RECT -201.725 -45.015 -201.325 -44.665 ;
        RECT -199.485 -45.015 -199.085 -44.665 ;
        RECT -197.245 -45.015 -196.845 -44.665 ;
        RECT -195.005 -45.015 -194.605 -44.665 ;
        RECT -192.765 -45.015 -192.365 -44.665 ;
        RECT -190.525 -45.015 -190.125 -44.665 ;
        RECT -187.165 -45.015 -186.765 -44.665 ;
        RECT -184.925 -45.015 -184.525 -44.665 ;
        RECT -182.685 -45.015 -182.285 -44.665 ;
        RECT -180.445 -45.015 -180.045 -44.665 ;
        RECT -178.205 -45.015 -177.805 -44.665 ;
        RECT -175.965 -45.015 -175.565 -44.665 ;
        RECT -173.725 -45.015 -173.325 -44.665 ;
        RECT -171.485 -45.015 -171.085 -44.665 ;
        RECT -169.245 -45.015 -168.845 -44.665 ;
        RECT -167.005 -45.015 -166.605 -44.665 ;
        RECT -164.765 -45.015 -164.365 -44.665 ;
        RECT -162.525 -45.015 -162.125 -44.665 ;
        RECT -160.285 -45.015 -159.885 -44.665 ;
        RECT -158.045 -45.015 -157.645 -44.665 ;
        RECT -155.805 -45.015 -155.405 -44.665 ;
        RECT -153.565 -45.015 -153.165 -44.665 ;
        RECT -151.325 -45.015 -150.925 -44.665 ;
        RECT -149.085 -45.015 -148.685 -44.665 ;
        RECT -146.845 -45.015 -146.445 -44.665 ;
        RECT -144.605 -45.015 -144.205 -44.665 ;
        RECT -142.365 -45.015 -141.965 -44.665 ;
        RECT -140.125 -45.015 -139.725 -44.665 ;
        RECT -137.885 -45.015 -137.485 -44.665 ;
        RECT -135.645 -45.015 -135.245 -44.665 ;
        RECT -133.405 -45.015 -133.005 -44.665 ;
        RECT -131.165 -45.015 -130.765 -44.665 ;
        RECT -128.925 -45.015 -128.525 -44.665 ;
        RECT -126.685 -45.015 -126.285 -44.665 ;
        RECT -124.445 -45.015 -124.045 -44.665 ;
        RECT -122.205 -45.015 -121.805 -44.665 ;
        RECT -119.965 -45.015 -119.565 -44.665 ;
        RECT -117.725 -45.015 -117.325 -44.665 ;
        RECT -115.485 -45.015 -115.085 -44.665 ;
        RECT -113.245 -45.015 -112.845 -44.665 ;
        RECT -111.005 -45.015 -110.605 -44.665 ;
        RECT -108.765 -45.015 -108.365 -44.665 ;
        RECT -106.525 -45.015 -106.125 -44.665 ;
        RECT -104.285 -45.015 -103.885 -44.665 ;
        RECT -102.045 -45.015 -101.645 -44.665 ;
        RECT -99.805 -45.015 -99.405 -44.665 ;
        RECT -97.565 -45.015 -97.165 -44.665 ;
        RECT -95.325 -45.015 -94.925 -44.665 ;
        RECT -93.085 -45.015 -92.685 -44.665 ;
        RECT -90.845 -45.015 -90.445 -44.665 ;
        RECT -88.605 -45.015 -88.205 -44.665 ;
        RECT -86.365 -45.015 -85.965 -44.665 ;
        RECT -84.125 -45.015 -83.725 -44.665 ;
        RECT -81.885 -45.015 -81.485 -44.665 ;
        RECT -79.645 -45.015 -79.245 -44.665 ;
        RECT -77.405 -45.015 -77.005 -44.665 ;
        RECT -75.165 -45.015 -74.765 -44.665 ;
        RECT -72.925 -45.015 -72.525 -44.665 ;
        RECT -70.685 -45.015 -70.285 -44.665 ;
        RECT -68.445 -45.015 -68.045 -44.665 ;
        RECT -66.205 -45.015 -65.805 -44.665 ;
        RECT -63.965 -45.015 -63.565 -44.665 ;
        RECT -61.725 -45.015 -61.325 -44.665 ;
        RECT -59.485 -45.015 -59.085 -44.665 ;
        RECT -57.245 -45.015 -56.845 -44.665 ;
        RECT -55.005 -45.015 -54.605 -44.665 ;
        RECT -52.765 -45.015 -52.365 -44.665 ;
        RECT -50.525 -45.015 -50.125 -44.665 ;
        RECT -48.285 -45.015 -47.885 -44.665 ;
        RECT -46.045 -45.015 -45.645 -44.665 ;
        RECT -43.805 -45.015 -43.405 -44.665 ;
        RECT -41.565 -45.015 -41.165 -44.665 ;
        RECT -39.325 -45.015 -38.925 -44.665 ;
        RECT -37.085 -45.015 -36.685 -44.665 ;
        RECT -34.845 -45.015 -34.445 -44.665 ;
        RECT -32.605 -45.015 -32.205 -44.665 ;
        RECT -30.365 -45.015 -29.965 -44.665 ;
        RECT -28.125 -45.015 -27.725 -44.665 ;
        RECT -25.885 -45.015 -25.485 -44.665 ;
        RECT -23.645 -45.015 -23.245 -44.665 ;
        RECT -21.405 -45.015 -21.005 -44.665 ;
        RECT -19.165 -45.015 -18.765 -44.665 ;
        RECT -16.925 -45.015 -16.525 -44.665 ;
        RECT -14.685 -45.015 -14.285 -44.665 ;
        RECT -12.445 -45.015 -12.045 -44.665 ;
        RECT -10.205 -45.015 -9.805 -44.665 ;
        RECT -7.965 -45.015 -7.565 -44.665 ;
        RECT -5.725 -45.015 -5.325 -44.665 ;
        RECT -3.485 -45.015 -3.085 -44.665 ;
        RECT -1.245 -45.015 -0.845 -44.665 ;
        RECT 0.995 -45.015 1.395 -44.665 ;
        RECT 3.235 -45.015 3.635 -44.665 ;
        RECT 5.475 -45.015 5.875 -44.665 ;
        RECT 7.715 -45.015 8.115 -44.665 ;
        RECT 9.955 -45.015 10.355 -44.665 ;
        RECT 12.195 -45.015 12.595 -44.665 ;
        RECT 14.435 -45.015 14.835 -44.665 ;
        RECT 16.675 -45.015 17.075 -44.665 ;
        RECT 18.915 -45.015 19.315 -44.665 ;
        RECT 21.155 -45.015 21.555 -44.665 ;
        RECT 23.395 -45.015 23.795 -44.665 ;
        RECT 25.635 -45.015 26.035 -44.665 ;
        RECT 27.875 -45.015 28.275 -44.665 ;
        RECT 30.115 -45.015 30.515 -44.665 ;
        RECT 32.355 -45.015 32.755 -44.665 ;
        RECT 34.595 -45.015 34.995 -44.665 ;
        RECT 36.835 -45.015 37.235 -44.665 ;
        RECT 39.075 -45.015 39.475 -44.665 ;
        RECT 41.315 -45.015 41.715 -44.665 ;
        RECT 43.555 -45.015 43.955 -44.665 ;
        RECT 45.795 -45.015 46.195 -44.665 ;
        RECT 48.035 -45.015 48.435 -44.665 ;
        RECT 50.275 -45.015 50.675 -44.665 ;
        RECT 52.515 -45.015 52.915 -44.665 ;
        RECT 54.755 -45.015 55.155 -44.665 ;
        RECT 56.995 -45.015 57.395 -44.665 ;
        RECT 59.235 -45.015 59.635 -44.665 ;
        RECT 61.475 -45.015 61.875 -44.665 ;
        RECT 63.715 -45.015 64.115 -44.665 ;
        RECT 65.955 -45.015 66.355 -44.665 ;
        RECT 68.195 -45.015 68.595 -44.665 ;
        RECT 70.435 -45.015 70.835 -44.665 ;
        RECT 72.675 -45.015 73.075 -44.665 ;
        RECT 74.915 -45.015 75.315 -44.665 ;
        RECT 77.155 -45.015 77.555 -44.665 ;
        RECT 79.395 -45.015 79.795 -44.665 ;
        RECT 81.635 -45.015 82.035 -44.665 ;
        RECT 83.875 -45.015 84.275 -44.665 ;
        RECT 86.115 -45.015 86.515 -44.665 ;
        RECT 88.355 -45.015 88.755 -44.665 ;
        RECT 90.595 -45.015 90.995 -44.665 ;
        RECT 92.835 -45.015 93.235 -44.665 ;
        RECT 95.075 -45.015 95.475 -44.665 ;
        RECT 97.315 -45.015 97.715 -44.665 ;
        RECT -497.305 -46.300 -486.905 -45.700 ;
        RECT -497.305 -54.300 -495.505 -46.300 ;
        RECT -487.505 -54.300 -486.905 -46.300 ;
        RECT -497.305 -54.900 -486.905 -54.300 ;
        RECT -497.305 -58.300 -486.905 -57.700 ;
        RECT -497.305 -66.300 -495.505 -58.300 ;
        RECT -487.505 -66.300 -486.905 -58.300 ;
        RECT 117.705 -63.665 118.205 -14.425 ;
        RECT 117.705 -64.165 121.925 -63.665 ;
        RECT -497.305 -66.900 -486.905 -66.300 ;
        RECT -475.005 -67.025 -474.605 -66.675 ;
        RECT -472.765 -67.025 -472.365 -66.675 ;
        RECT -470.525 -67.025 -470.125 -66.675 ;
        RECT -468.285 -67.025 -467.885 -66.675 ;
        RECT -466.045 -67.025 -465.645 -66.675 ;
        RECT -463.805 -67.025 -463.405 -66.675 ;
        RECT -461.565 -67.025 -461.165 -66.675 ;
        RECT -459.325 -67.025 -458.925 -66.675 ;
        RECT -457.085 -67.025 -456.685 -66.675 ;
        RECT -454.845 -67.025 -454.445 -66.675 ;
        RECT -452.605 -67.025 -452.205 -66.675 ;
        RECT -450.365 -67.025 -449.965 -66.675 ;
        RECT -448.125 -67.025 -447.725 -66.675 ;
        RECT -445.885 -67.025 -445.485 -66.675 ;
        RECT -443.645 -67.025 -443.245 -66.675 ;
        RECT -441.405 -67.025 -441.005 -66.675 ;
        RECT -439.165 -67.025 -438.765 -66.675 ;
        RECT -436.925 -67.025 -436.525 -66.675 ;
        RECT -434.685 -67.025 -434.285 -66.675 ;
        RECT -432.445 -67.025 -432.045 -66.675 ;
        RECT -430.205 -67.025 -429.805 -66.675 ;
        RECT -427.965 -67.025 -427.565 -66.675 ;
        RECT -425.725 -67.025 -425.325 -66.675 ;
        RECT -423.485 -67.025 -423.085 -66.675 ;
        RECT -421.245 -67.025 -420.845 -66.675 ;
        RECT -419.005 -67.025 -418.605 -66.675 ;
        RECT -416.765 -67.025 -416.365 -66.675 ;
        RECT -414.525 -67.025 -414.125 -66.675 ;
        RECT -412.285 -67.025 -411.885 -66.675 ;
        RECT -410.045 -67.025 -409.645 -66.675 ;
        RECT -407.805 -67.025 -407.405 -66.675 ;
        RECT -405.565 -67.025 -405.165 -66.675 ;
        RECT -403.325 -67.025 -402.925 -66.675 ;
        RECT -401.085 -67.025 -400.685 -66.675 ;
        RECT -398.845 -67.025 -398.445 -66.675 ;
        RECT -396.605 -67.025 -396.205 -66.675 ;
        RECT -394.365 -67.025 -393.965 -66.675 ;
        RECT -392.125 -67.025 -391.725 -66.675 ;
        RECT -389.885 -67.025 -389.485 -66.675 ;
        RECT -387.645 -67.025 -387.245 -66.675 ;
        RECT -385.405 -67.025 -385.005 -66.675 ;
        RECT -383.165 -67.025 -382.765 -66.675 ;
        RECT -380.925 -67.025 -380.525 -66.675 ;
        RECT -378.685 -67.025 -378.285 -66.675 ;
        RECT -376.445 -67.025 -376.045 -66.675 ;
        RECT -374.205 -67.025 -373.805 -66.675 ;
        RECT -371.965 -67.025 -371.565 -66.675 ;
        RECT -369.725 -67.025 -369.325 -66.675 ;
        RECT -367.485 -67.025 -367.085 -66.675 ;
        RECT -365.245 -67.025 -364.845 -66.675 ;
        RECT -363.005 -67.025 -362.605 -66.675 ;
        RECT -360.765 -67.025 -360.365 -66.675 ;
        RECT -358.525 -67.025 -358.125 -66.675 ;
        RECT -356.285 -67.025 -355.885 -66.675 ;
        RECT -354.045 -67.025 -353.645 -66.675 ;
        RECT -351.805 -67.025 -351.405 -66.675 ;
        RECT -349.565 -67.025 -349.165 -66.675 ;
        RECT -347.325 -67.025 -346.925 -66.675 ;
        RECT -345.085 -67.025 -344.685 -66.675 ;
        RECT -342.845 -67.025 -342.445 -66.675 ;
        RECT -340.605 -67.025 -340.205 -66.675 ;
        RECT -338.365 -67.025 -337.965 -66.675 ;
        RECT -336.125 -67.025 -335.725 -66.675 ;
        RECT -333.885 -67.025 -333.485 -66.675 ;
        RECT -331.645 -67.025 -331.245 -66.675 ;
        RECT -329.405 -67.025 -329.005 -66.675 ;
        RECT -327.165 -67.025 -326.765 -66.675 ;
        RECT -324.925 -67.025 -324.525 -66.675 ;
        RECT -322.685 -67.025 -322.285 -66.675 ;
        RECT -320.445 -67.025 -320.045 -66.675 ;
        RECT -318.205 -67.025 -317.805 -66.675 ;
        RECT -315.965 -67.025 -315.565 -66.675 ;
        RECT -313.725 -67.025 -313.325 -66.675 ;
        RECT -311.485 -67.025 -311.085 -66.675 ;
        RECT -309.245 -67.025 -308.845 -66.675 ;
        RECT -307.005 -67.025 -306.605 -66.675 ;
        RECT -304.765 -67.025 -304.365 -66.675 ;
        RECT -302.525 -67.025 -302.125 -66.675 ;
        RECT -300.285 -67.025 -299.885 -66.675 ;
        RECT -298.045 -67.025 -297.645 -66.675 ;
        RECT -295.805 -67.025 -295.405 -66.675 ;
        RECT -293.565 -67.025 -293.165 -66.675 ;
        RECT -291.325 -67.025 -290.925 -66.675 ;
        RECT -289.085 -67.025 -288.685 -66.675 ;
        RECT -286.845 -67.025 -286.445 -66.675 ;
        RECT -284.605 -67.025 -284.205 -66.675 ;
        RECT -282.365 -67.025 -281.965 -66.675 ;
        RECT -280.125 -67.025 -279.725 -66.675 ;
        RECT -277.885 -67.025 -277.485 -66.675 ;
        RECT -275.645 -67.025 -275.245 -66.675 ;
        RECT -273.405 -67.025 -273.005 -66.675 ;
        RECT -271.165 -67.025 -270.765 -66.675 ;
        RECT -268.925 -67.025 -268.525 -66.675 ;
        RECT -266.685 -67.025 -266.285 -66.675 ;
        RECT -264.445 -67.025 -264.045 -66.675 ;
        RECT -262.205 -67.025 -261.805 -66.675 ;
        RECT -259.965 -67.025 -259.565 -66.675 ;
        RECT -257.725 -67.025 -257.325 -66.675 ;
        RECT -255.485 -67.025 -255.085 -66.675 ;
        RECT -253.245 -67.025 -252.845 -66.675 ;
        RECT -251.005 -67.025 -250.605 -66.675 ;
        RECT -248.765 -67.025 -248.365 -66.675 ;
        RECT -246.525 -67.025 -246.125 -66.675 ;
        RECT -244.285 -67.025 -243.885 -66.675 ;
        RECT -242.045 -67.025 -241.645 -66.675 ;
        RECT -239.805 -67.025 -239.405 -66.675 ;
        RECT -237.565 -67.025 -237.165 -66.675 ;
        RECT -235.325 -67.025 -234.925 -66.675 ;
        RECT -233.085 -67.025 -232.685 -66.675 ;
        RECT -230.845 -67.025 -230.445 -66.675 ;
        RECT -228.605 -67.025 -228.205 -66.675 ;
        RECT -226.365 -67.025 -225.965 -66.675 ;
        RECT -224.125 -67.025 -223.725 -66.675 ;
        RECT -221.885 -67.025 -221.485 -66.675 ;
        RECT -219.645 -67.025 -219.245 -66.675 ;
        RECT -217.405 -67.025 -217.005 -66.675 ;
        RECT -215.165 -67.025 -214.765 -66.675 ;
        RECT -212.925 -67.025 -212.525 -66.675 ;
        RECT -210.685 -67.025 -210.285 -66.675 ;
        RECT -208.445 -67.025 -208.045 -66.675 ;
        RECT -206.205 -67.025 -205.805 -66.675 ;
        RECT -203.965 -67.025 -203.565 -66.675 ;
        RECT -201.725 -67.025 -201.325 -66.675 ;
        RECT -199.485 -67.025 -199.085 -66.675 ;
        RECT -197.245 -67.025 -196.845 -66.675 ;
        RECT -195.005 -67.025 -194.605 -66.675 ;
        RECT -192.765 -67.025 -192.365 -66.675 ;
        RECT -190.525 -67.025 -190.125 -66.675 ;
        RECT -187.165 -67.025 -186.765 -66.675 ;
        RECT -184.925 -67.025 -184.525 -66.675 ;
        RECT -182.685 -67.025 -182.285 -66.675 ;
        RECT -180.445 -67.025 -180.045 -66.675 ;
        RECT -178.205 -67.025 -177.805 -66.675 ;
        RECT -175.965 -67.025 -175.565 -66.675 ;
        RECT -173.725 -67.025 -173.325 -66.675 ;
        RECT -171.485 -67.025 -171.085 -66.675 ;
        RECT -169.245 -67.025 -168.845 -66.675 ;
        RECT -167.005 -67.025 -166.605 -66.675 ;
        RECT -164.765 -67.025 -164.365 -66.675 ;
        RECT -162.525 -67.025 -162.125 -66.675 ;
        RECT -160.285 -67.025 -159.885 -66.675 ;
        RECT -158.045 -67.025 -157.645 -66.675 ;
        RECT -155.805 -67.025 -155.405 -66.675 ;
        RECT -153.565 -67.025 -153.165 -66.675 ;
        RECT -151.325 -67.025 -150.925 -66.675 ;
        RECT -149.085 -67.025 -148.685 -66.675 ;
        RECT -146.845 -67.025 -146.445 -66.675 ;
        RECT -144.605 -67.025 -144.205 -66.675 ;
        RECT -142.365 -67.025 -141.965 -66.675 ;
        RECT -140.125 -67.025 -139.725 -66.675 ;
        RECT -137.885 -67.025 -137.485 -66.675 ;
        RECT -135.645 -67.025 -135.245 -66.675 ;
        RECT -133.405 -67.025 -133.005 -66.675 ;
        RECT -131.165 -67.025 -130.765 -66.675 ;
        RECT -128.925 -67.025 -128.525 -66.675 ;
        RECT -126.685 -67.025 -126.285 -66.675 ;
        RECT -124.445 -67.025 -124.045 -66.675 ;
        RECT -122.205 -67.025 -121.805 -66.675 ;
        RECT -119.965 -67.025 -119.565 -66.675 ;
        RECT -117.725 -67.025 -117.325 -66.675 ;
        RECT -115.485 -67.025 -115.085 -66.675 ;
        RECT -113.245 -67.025 -112.845 -66.675 ;
        RECT -111.005 -67.025 -110.605 -66.675 ;
        RECT -108.765 -67.025 -108.365 -66.675 ;
        RECT -106.525 -67.025 -106.125 -66.675 ;
        RECT -104.285 -67.025 -103.885 -66.675 ;
        RECT -102.045 -67.025 -101.645 -66.675 ;
        RECT -99.805 -67.025 -99.405 -66.675 ;
        RECT -97.565 -67.025 -97.165 -66.675 ;
        RECT -95.325 -67.025 -94.925 -66.675 ;
        RECT -93.085 -67.025 -92.685 -66.675 ;
        RECT -90.845 -67.025 -90.445 -66.675 ;
        RECT -88.605 -67.025 -88.205 -66.675 ;
        RECT -86.365 -67.025 -85.965 -66.675 ;
        RECT -84.125 -67.025 -83.725 -66.675 ;
        RECT -81.885 -67.025 -81.485 -66.675 ;
        RECT -79.645 -67.025 -79.245 -66.675 ;
        RECT -77.405 -67.025 -77.005 -66.675 ;
        RECT -75.165 -67.025 -74.765 -66.675 ;
        RECT -72.925 -67.025 -72.525 -66.675 ;
        RECT -70.685 -67.025 -70.285 -66.675 ;
        RECT -68.445 -67.025 -68.045 -66.675 ;
        RECT -66.205 -67.025 -65.805 -66.675 ;
        RECT -63.965 -67.025 -63.565 -66.675 ;
        RECT -61.725 -67.025 -61.325 -66.675 ;
        RECT -59.485 -67.025 -59.085 -66.675 ;
        RECT -57.245 -67.025 -56.845 -66.675 ;
        RECT -55.005 -67.025 -54.605 -66.675 ;
        RECT -52.765 -67.025 -52.365 -66.675 ;
        RECT -50.525 -67.025 -50.125 -66.675 ;
        RECT -48.285 -67.025 -47.885 -66.675 ;
        RECT -46.045 -67.025 -45.645 -66.675 ;
        RECT -43.805 -67.025 -43.405 -66.675 ;
        RECT -41.565 -67.025 -41.165 -66.675 ;
        RECT -39.325 -67.025 -38.925 -66.675 ;
        RECT -37.085 -67.025 -36.685 -66.675 ;
        RECT -34.845 -67.025 -34.445 -66.675 ;
        RECT -32.605 -67.025 -32.205 -66.675 ;
        RECT -30.365 -67.025 -29.965 -66.675 ;
        RECT -28.125 -67.025 -27.725 -66.675 ;
        RECT -25.885 -67.025 -25.485 -66.675 ;
        RECT -23.645 -67.025 -23.245 -66.675 ;
        RECT -21.405 -67.025 -21.005 -66.675 ;
        RECT -19.165 -67.025 -18.765 -66.675 ;
        RECT -16.925 -67.025 -16.525 -66.675 ;
        RECT -14.685 -67.025 -14.285 -66.675 ;
        RECT -12.445 -67.025 -12.045 -66.675 ;
        RECT -10.205 -67.025 -9.805 -66.675 ;
        RECT -7.965 -67.025 -7.565 -66.675 ;
        RECT -5.725 -67.025 -5.325 -66.675 ;
        RECT -3.485 -67.025 -3.085 -66.675 ;
        RECT -1.245 -67.025 -0.845 -66.675 ;
        RECT 0.995 -67.025 1.395 -66.675 ;
        RECT 3.235 -67.025 3.635 -66.675 ;
        RECT 5.475 -67.025 5.875 -66.675 ;
        RECT 7.715 -67.025 8.115 -66.675 ;
        RECT 9.955 -67.025 10.355 -66.675 ;
        RECT 12.195 -67.025 12.595 -66.675 ;
        RECT 14.435 -67.025 14.835 -66.675 ;
        RECT 16.675 -67.025 17.075 -66.675 ;
        RECT 18.915 -67.025 19.315 -66.675 ;
        RECT 21.155 -67.025 21.555 -66.675 ;
        RECT 23.395 -67.025 23.795 -66.675 ;
        RECT 25.635 -67.025 26.035 -66.675 ;
        RECT 27.875 -67.025 28.275 -66.675 ;
        RECT 30.115 -67.025 30.515 -66.675 ;
        RECT 32.355 -67.025 32.755 -66.675 ;
        RECT 34.595 -67.025 34.995 -66.675 ;
        RECT 36.835 -67.025 37.235 -66.675 ;
        RECT 39.075 -67.025 39.475 -66.675 ;
        RECT 41.315 -67.025 41.715 -66.675 ;
        RECT 43.555 -67.025 43.955 -66.675 ;
        RECT 45.795 -67.025 46.195 -66.675 ;
        RECT 48.035 -67.025 48.435 -66.675 ;
        RECT 50.275 -67.025 50.675 -66.675 ;
        RECT 52.515 -67.025 52.915 -66.675 ;
        RECT 54.755 -67.025 55.155 -66.675 ;
        RECT 56.995 -67.025 57.395 -66.675 ;
        RECT 59.235 -67.025 59.635 -66.675 ;
        RECT 61.475 -67.025 61.875 -66.675 ;
        RECT 63.715 -67.025 64.115 -66.675 ;
        RECT 65.955 -67.025 66.355 -66.675 ;
        RECT 68.195 -67.025 68.595 -66.675 ;
        RECT 70.435 -67.025 70.835 -66.675 ;
        RECT 72.675 -67.025 73.075 -66.675 ;
        RECT 74.915 -67.025 75.315 -66.675 ;
        RECT 77.155 -67.025 77.555 -66.675 ;
        RECT 79.395 -67.025 79.795 -66.675 ;
        RECT 81.635 -67.025 82.035 -66.675 ;
        RECT 83.875 -67.025 84.275 -66.675 ;
        RECT 86.115 -67.025 86.515 -66.675 ;
        RECT 88.355 -67.025 88.755 -66.675 ;
        RECT 90.595 -67.025 90.995 -66.675 ;
        RECT 92.835 -67.025 93.235 -66.675 ;
        RECT 95.075 -67.025 95.475 -66.675 ;
        RECT 97.315 -67.025 97.715 -66.675 ;
        RECT -475.005 -67.525 121.925 -67.025 ;
        RECT -475.005 -67.875 -474.605 -67.525 ;
        RECT -472.765 -67.875 -472.365 -67.525 ;
        RECT -470.525 -67.875 -470.125 -67.525 ;
        RECT -468.285 -67.875 -467.885 -67.525 ;
        RECT -466.045 -67.875 -465.645 -67.525 ;
        RECT -463.805 -67.875 -463.405 -67.525 ;
        RECT -461.565 -67.875 -461.165 -67.525 ;
        RECT -459.325 -67.875 -458.925 -67.525 ;
        RECT -457.085 -67.875 -456.685 -67.525 ;
        RECT -454.845 -67.875 -454.445 -67.525 ;
        RECT -452.605 -67.875 -452.205 -67.525 ;
        RECT -450.365 -67.875 -449.965 -67.525 ;
        RECT -448.125 -67.875 -447.725 -67.525 ;
        RECT -445.885 -67.875 -445.485 -67.525 ;
        RECT -443.645 -67.875 -443.245 -67.525 ;
        RECT -441.405 -67.875 -441.005 -67.525 ;
        RECT -439.165 -67.875 -438.765 -67.525 ;
        RECT -436.925 -67.875 -436.525 -67.525 ;
        RECT -434.685 -67.875 -434.285 -67.525 ;
        RECT -432.445 -67.875 -432.045 -67.525 ;
        RECT -430.205 -67.875 -429.805 -67.525 ;
        RECT -427.965 -67.875 -427.565 -67.525 ;
        RECT -425.725 -67.875 -425.325 -67.525 ;
        RECT -423.485 -67.875 -423.085 -67.525 ;
        RECT -421.245 -67.875 -420.845 -67.525 ;
        RECT -419.005 -67.875 -418.605 -67.525 ;
        RECT -416.765 -67.875 -416.365 -67.525 ;
        RECT -414.525 -67.875 -414.125 -67.525 ;
        RECT -412.285 -67.875 -411.885 -67.525 ;
        RECT -410.045 -67.875 -409.645 -67.525 ;
        RECT -407.805 -67.875 -407.405 -67.525 ;
        RECT -405.565 -67.875 -405.165 -67.525 ;
        RECT -403.325 -67.875 -402.925 -67.525 ;
        RECT -401.085 -67.875 -400.685 -67.525 ;
        RECT -398.845 -67.875 -398.445 -67.525 ;
        RECT -396.605 -67.875 -396.205 -67.525 ;
        RECT -394.365 -67.875 -393.965 -67.525 ;
        RECT -392.125 -67.875 -391.725 -67.525 ;
        RECT -389.885 -67.875 -389.485 -67.525 ;
        RECT -387.645 -67.875 -387.245 -67.525 ;
        RECT -385.405 -67.875 -385.005 -67.525 ;
        RECT -383.165 -67.875 -382.765 -67.525 ;
        RECT -380.925 -67.875 -380.525 -67.525 ;
        RECT -378.685 -67.875 -378.285 -67.525 ;
        RECT -376.445 -67.875 -376.045 -67.525 ;
        RECT -374.205 -67.875 -373.805 -67.525 ;
        RECT -371.965 -67.875 -371.565 -67.525 ;
        RECT -369.725 -67.875 -369.325 -67.525 ;
        RECT -367.485 -67.875 -367.085 -67.525 ;
        RECT -365.245 -67.875 -364.845 -67.525 ;
        RECT -363.005 -67.875 -362.605 -67.525 ;
        RECT -360.765 -67.875 -360.365 -67.525 ;
        RECT -358.525 -67.875 -358.125 -67.525 ;
        RECT -356.285 -67.875 -355.885 -67.525 ;
        RECT -354.045 -67.875 -353.645 -67.525 ;
        RECT -351.805 -67.875 -351.405 -67.525 ;
        RECT -349.565 -67.875 -349.165 -67.525 ;
        RECT -347.325 -67.875 -346.925 -67.525 ;
        RECT -345.085 -67.875 -344.685 -67.525 ;
        RECT -342.845 -67.875 -342.445 -67.525 ;
        RECT -340.605 -67.875 -340.205 -67.525 ;
        RECT -338.365 -67.875 -337.965 -67.525 ;
        RECT -336.125 -67.875 -335.725 -67.525 ;
        RECT -333.885 -67.875 -333.485 -67.525 ;
        RECT -331.645 -67.875 -331.245 -67.525 ;
        RECT -329.405 -67.875 -329.005 -67.525 ;
        RECT -327.165 -67.875 -326.765 -67.525 ;
        RECT -324.925 -67.875 -324.525 -67.525 ;
        RECT -322.685 -67.875 -322.285 -67.525 ;
        RECT -320.445 -67.875 -320.045 -67.525 ;
        RECT -318.205 -67.875 -317.805 -67.525 ;
        RECT -315.965 -67.875 -315.565 -67.525 ;
        RECT -313.725 -67.875 -313.325 -67.525 ;
        RECT -311.485 -67.875 -311.085 -67.525 ;
        RECT -309.245 -67.875 -308.845 -67.525 ;
        RECT -307.005 -67.875 -306.605 -67.525 ;
        RECT -304.765 -67.875 -304.365 -67.525 ;
        RECT -302.525 -67.875 -302.125 -67.525 ;
        RECT -300.285 -67.875 -299.885 -67.525 ;
        RECT -298.045 -67.875 -297.645 -67.525 ;
        RECT -295.805 -67.875 -295.405 -67.525 ;
        RECT -293.565 -67.875 -293.165 -67.525 ;
        RECT -291.325 -67.875 -290.925 -67.525 ;
        RECT -289.085 -67.875 -288.685 -67.525 ;
        RECT -286.845 -67.875 -286.445 -67.525 ;
        RECT -284.605 -67.875 -284.205 -67.525 ;
        RECT -282.365 -67.875 -281.965 -67.525 ;
        RECT -280.125 -67.875 -279.725 -67.525 ;
        RECT -277.885 -67.875 -277.485 -67.525 ;
        RECT -275.645 -67.875 -275.245 -67.525 ;
        RECT -273.405 -67.875 -273.005 -67.525 ;
        RECT -271.165 -67.875 -270.765 -67.525 ;
        RECT -268.925 -67.875 -268.525 -67.525 ;
        RECT -266.685 -67.875 -266.285 -67.525 ;
        RECT -264.445 -67.875 -264.045 -67.525 ;
        RECT -262.205 -67.875 -261.805 -67.525 ;
        RECT -259.965 -67.875 -259.565 -67.525 ;
        RECT -257.725 -67.875 -257.325 -67.525 ;
        RECT -255.485 -67.875 -255.085 -67.525 ;
        RECT -253.245 -67.875 -252.845 -67.525 ;
        RECT -251.005 -67.875 -250.605 -67.525 ;
        RECT -248.765 -67.875 -248.365 -67.525 ;
        RECT -246.525 -67.875 -246.125 -67.525 ;
        RECT -244.285 -67.875 -243.885 -67.525 ;
        RECT -242.045 -67.875 -241.645 -67.525 ;
        RECT -239.805 -67.875 -239.405 -67.525 ;
        RECT -237.565 -67.875 -237.165 -67.525 ;
        RECT -235.325 -67.875 -234.925 -67.525 ;
        RECT -233.085 -67.875 -232.685 -67.525 ;
        RECT -230.845 -67.875 -230.445 -67.525 ;
        RECT -228.605 -67.875 -228.205 -67.525 ;
        RECT -226.365 -67.875 -225.965 -67.525 ;
        RECT -224.125 -67.875 -223.725 -67.525 ;
        RECT -221.885 -67.875 -221.485 -67.525 ;
        RECT -219.645 -67.875 -219.245 -67.525 ;
        RECT -217.405 -67.875 -217.005 -67.525 ;
        RECT -215.165 -67.875 -214.765 -67.525 ;
        RECT -212.925 -67.875 -212.525 -67.525 ;
        RECT -210.685 -67.875 -210.285 -67.525 ;
        RECT -208.445 -67.875 -208.045 -67.525 ;
        RECT -206.205 -67.875 -205.805 -67.525 ;
        RECT -203.965 -67.875 -203.565 -67.525 ;
        RECT -201.725 -67.875 -201.325 -67.525 ;
        RECT -199.485 -67.875 -199.085 -67.525 ;
        RECT -197.245 -67.875 -196.845 -67.525 ;
        RECT -195.005 -67.875 -194.605 -67.525 ;
        RECT -192.765 -67.875 -192.365 -67.525 ;
        RECT -190.525 -67.875 -190.125 -67.525 ;
        RECT -187.165 -67.875 -186.765 -67.525 ;
        RECT -184.925 -67.875 -184.525 -67.525 ;
        RECT -182.685 -67.875 -182.285 -67.525 ;
        RECT -180.445 -67.875 -180.045 -67.525 ;
        RECT -178.205 -67.875 -177.805 -67.525 ;
        RECT -175.965 -67.875 -175.565 -67.525 ;
        RECT -173.725 -67.875 -173.325 -67.525 ;
        RECT -171.485 -67.875 -171.085 -67.525 ;
        RECT -169.245 -67.875 -168.845 -67.525 ;
        RECT -167.005 -67.875 -166.605 -67.525 ;
        RECT -164.765 -67.875 -164.365 -67.525 ;
        RECT -162.525 -67.875 -162.125 -67.525 ;
        RECT -160.285 -67.875 -159.885 -67.525 ;
        RECT -158.045 -67.875 -157.645 -67.525 ;
        RECT -155.805 -67.875 -155.405 -67.525 ;
        RECT -153.565 -67.875 -153.165 -67.525 ;
        RECT -151.325 -67.875 -150.925 -67.525 ;
        RECT -149.085 -67.875 -148.685 -67.525 ;
        RECT -146.845 -67.875 -146.445 -67.525 ;
        RECT -144.605 -67.875 -144.205 -67.525 ;
        RECT -142.365 -67.875 -141.965 -67.525 ;
        RECT -140.125 -67.875 -139.725 -67.525 ;
        RECT -137.885 -67.875 -137.485 -67.525 ;
        RECT -135.645 -67.875 -135.245 -67.525 ;
        RECT -133.405 -67.875 -133.005 -67.525 ;
        RECT -131.165 -67.875 -130.765 -67.525 ;
        RECT -128.925 -67.875 -128.525 -67.525 ;
        RECT -126.685 -67.875 -126.285 -67.525 ;
        RECT -124.445 -67.875 -124.045 -67.525 ;
        RECT -122.205 -67.875 -121.805 -67.525 ;
        RECT -119.965 -67.875 -119.565 -67.525 ;
        RECT -117.725 -67.875 -117.325 -67.525 ;
        RECT -115.485 -67.875 -115.085 -67.525 ;
        RECT -113.245 -67.875 -112.845 -67.525 ;
        RECT -111.005 -67.875 -110.605 -67.525 ;
        RECT -108.765 -67.875 -108.365 -67.525 ;
        RECT -106.525 -67.875 -106.125 -67.525 ;
        RECT -104.285 -67.875 -103.885 -67.525 ;
        RECT -102.045 -67.875 -101.645 -67.525 ;
        RECT -99.805 -67.875 -99.405 -67.525 ;
        RECT -97.565 -67.875 -97.165 -67.525 ;
        RECT -95.325 -67.875 -94.925 -67.525 ;
        RECT -93.085 -67.875 -92.685 -67.525 ;
        RECT -90.845 -67.875 -90.445 -67.525 ;
        RECT -88.605 -67.875 -88.205 -67.525 ;
        RECT -86.365 -67.875 -85.965 -67.525 ;
        RECT -84.125 -67.875 -83.725 -67.525 ;
        RECT -81.885 -67.875 -81.485 -67.525 ;
        RECT -79.645 -67.875 -79.245 -67.525 ;
        RECT -77.405 -67.875 -77.005 -67.525 ;
        RECT -75.165 -67.875 -74.765 -67.525 ;
        RECT -72.925 -67.875 -72.525 -67.525 ;
        RECT -70.685 -67.875 -70.285 -67.525 ;
        RECT -68.445 -67.875 -68.045 -67.525 ;
        RECT -66.205 -67.875 -65.805 -67.525 ;
        RECT -63.965 -67.875 -63.565 -67.525 ;
        RECT -61.725 -67.875 -61.325 -67.525 ;
        RECT -59.485 -67.875 -59.085 -67.525 ;
        RECT -57.245 -67.875 -56.845 -67.525 ;
        RECT -55.005 -67.875 -54.605 -67.525 ;
        RECT -52.765 -67.875 -52.365 -67.525 ;
        RECT -50.525 -67.875 -50.125 -67.525 ;
        RECT -48.285 -67.875 -47.885 -67.525 ;
        RECT -46.045 -67.875 -45.645 -67.525 ;
        RECT -43.805 -67.875 -43.405 -67.525 ;
        RECT -41.565 -67.875 -41.165 -67.525 ;
        RECT -39.325 -67.875 -38.925 -67.525 ;
        RECT -37.085 -67.875 -36.685 -67.525 ;
        RECT -34.845 -67.875 -34.445 -67.525 ;
        RECT -32.605 -67.875 -32.205 -67.525 ;
        RECT -30.365 -67.875 -29.965 -67.525 ;
        RECT -28.125 -67.875 -27.725 -67.525 ;
        RECT -25.885 -67.875 -25.485 -67.525 ;
        RECT -23.645 -67.875 -23.245 -67.525 ;
        RECT -21.405 -67.875 -21.005 -67.525 ;
        RECT -19.165 -67.875 -18.765 -67.525 ;
        RECT -16.925 -67.875 -16.525 -67.525 ;
        RECT -14.685 -67.875 -14.285 -67.525 ;
        RECT -12.445 -67.875 -12.045 -67.525 ;
        RECT -10.205 -67.875 -9.805 -67.525 ;
        RECT -7.965 -67.875 -7.565 -67.525 ;
        RECT -5.725 -67.875 -5.325 -67.525 ;
        RECT -3.485 -67.875 -3.085 -67.525 ;
        RECT -1.245 -67.875 -0.845 -67.525 ;
        RECT 0.995 -67.875 1.395 -67.525 ;
        RECT 3.235 -67.875 3.635 -67.525 ;
        RECT 5.475 -67.875 5.875 -67.525 ;
        RECT 7.715 -67.875 8.115 -67.525 ;
        RECT 9.955 -67.875 10.355 -67.525 ;
        RECT 12.195 -67.875 12.595 -67.525 ;
        RECT 14.435 -67.875 14.835 -67.525 ;
        RECT 16.675 -67.875 17.075 -67.525 ;
        RECT 18.915 -67.875 19.315 -67.525 ;
        RECT 21.155 -67.875 21.555 -67.525 ;
        RECT 23.395 -67.875 23.795 -67.525 ;
        RECT 25.635 -67.875 26.035 -67.525 ;
        RECT 27.875 -67.875 28.275 -67.525 ;
        RECT 30.115 -67.875 30.515 -67.525 ;
        RECT 32.355 -67.875 32.755 -67.525 ;
        RECT 34.595 -67.875 34.995 -67.525 ;
        RECT 36.835 -67.875 37.235 -67.525 ;
        RECT 39.075 -67.875 39.475 -67.525 ;
        RECT 41.315 -67.875 41.715 -67.525 ;
        RECT 43.555 -67.875 43.955 -67.525 ;
        RECT 45.795 -67.875 46.195 -67.525 ;
        RECT 48.035 -67.875 48.435 -67.525 ;
        RECT 50.275 -67.875 50.675 -67.525 ;
        RECT 52.515 -67.875 52.915 -67.525 ;
        RECT 54.755 -67.875 55.155 -67.525 ;
        RECT 56.995 -67.875 57.395 -67.525 ;
        RECT 59.235 -67.875 59.635 -67.525 ;
        RECT 61.475 -67.875 61.875 -67.525 ;
        RECT 63.715 -67.875 64.115 -67.525 ;
        RECT 65.955 -67.875 66.355 -67.525 ;
        RECT 68.195 -67.875 68.595 -67.525 ;
        RECT 70.435 -67.875 70.835 -67.525 ;
        RECT 72.675 -67.875 73.075 -67.525 ;
        RECT 74.915 -67.875 75.315 -67.525 ;
        RECT 77.155 -67.875 77.555 -67.525 ;
        RECT 79.395 -67.875 79.795 -67.525 ;
        RECT 81.635 -67.875 82.035 -67.525 ;
        RECT 83.875 -67.875 84.275 -67.525 ;
        RECT 86.115 -67.875 86.515 -67.525 ;
        RECT 88.355 -67.875 88.755 -67.525 ;
        RECT 90.595 -67.875 90.995 -67.525 ;
        RECT 92.835 -67.875 93.235 -67.525 ;
        RECT 95.075 -67.875 95.475 -67.525 ;
        RECT 97.315 -67.875 97.715 -67.525 ;
        RECT -497.305 -70.300 -486.905 -69.700 ;
        RECT -497.305 -78.300 -495.505 -70.300 ;
        RECT -487.505 -78.300 -486.905 -70.300 ;
        RECT -473.885 -70.385 -473.485 -70.035 ;
        RECT -469.405 -70.385 -469.005 -70.035 ;
        RECT -464.925 -70.385 -464.525 -70.035 ;
        RECT -460.445 -70.385 -460.045 -70.035 ;
        RECT -455.965 -70.385 -455.565 -70.035 ;
        RECT -451.485 -70.385 -451.085 -70.035 ;
        RECT -447.005 -70.385 -446.605 -70.035 ;
        RECT -442.525 -70.385 -442.125 -70.035 ;
        RECT -438.045 -70.385 -437.645 -70.035 ;
        RECT -433.565 -70.385 -433.165 -70.035 ;
        RECT -429.085 -70.385 -428.685 -70.035 ;
        RECT -424.605 -70.385 -424.205 -70.035 ;
        RECT -420.125 -70.385 -419.725 -70.035 ;
        RECT -415.645 -70.385 -415.245 -70.035 ;
        RECT -411.165 -70.385 -410.765 -70.035 ;
        RECT -406.685 -70.385 -406.285 -70.035 ;
        RECT -402.205 -70.385 -401.805 -70.035 ;
        RECT -397.725 -70.385 -397.325 -70.035 ;
        RECT -393.245 -70.385 -392.845 -70.035 ;
        RECT -388.765 -70.385 -388.365 -70.035 ;
        RECT -384.285 -70.385 -383.885 -70.035 ;
        RECT -379.805 -70.385 -379.405 -70.035 ;
        RECT -375.325 -70.385 -374.925 -70.035 ;
        RECT -370.845 -70.385 -370.445 -70.035 ;
        RECT -366.365 -70.385 -365.965 -70.035 ;
        RECT -361.885 -70.385 -361.485 -70.035 ;
        RECT -357.405 -70.385 -357.005 -70.035 ;
        RECT -352.925 -70.385 -352.525 -70.035 ;
        RECT -348.445 -70.385 -348.045 -70.035 ;
        RECT -343.965 -70.385 -343.565 -70.035 ;
        RECT -339.485 -70.385 -339.085 -70.035 ;
        RECT -335.005 -70.385 -334.605 -70.035 ;
        RECT -330.525 -70.385 -330.125 -70.035 ;
        RECT -326.045 -70.385 -325.645 -70.035 ;
        RECT -321.565 -70.385 -321.165 -70.035 ;
        RECT -317.085 -70.385 -316.685 -70.035 ;
        RECT -312.605 -70.385 -312.205 -70.035 ;
        RECT -308.125 -70.385 -307.725 -70.035 ;
        RECT -303.645 -70.385 -303.245 -70.035 ;
        RECT -299.165 -70.385 -298.765 -70.035 ;
        RECT -294.685 -70.385 -294.285 -70.035 ;
        RECT -290.205 -70.385 -289.805 -70.035 ;
        RECT -285.725 -70.385 -285.325 -70.035 ;
        RECT -281.245 -70.385 -280.845 -70.035 ;
        RECT -276.765 -70.385 -276.365 -70.035 ;
        RECT -272.285 -70.385 -271.885 -70.035 ;
        RECT -267.805 -70.385 -267.405 -70.035 ;
        RECT -263.325 -70.385 -262.925 -70.035 ;
        RECT -258.845 -70.385 -258.445 -70.035 ;
        RECT -254.365 -70.385 -253.965 -70.035 ;
        RECT -249.885 -70.385 -249.485 -70.035 ;
        RECT -245.405 -70.385 -245.005 -70.035 ;
        RECT -240.925 -70.385 -240.525 -70.035 ;
        RECT -236.445 -70.385 -236.045 -70.035 ;
        RECT -231.965 -70.385 -231.565 -70.035 ;
        RECT -227.485 -70.385 -227.085 -70.035 ;
        RECT -223.005 -70.385 -222.605 -70.035 ;
        RECT -218.525 -70.385 -218.125 -70.035 ;
        RECT -214.045 -70.385 -213.645 -70.035 ;
        RECT -209.565 -70.385 -209.165 -70.035 ;
        RECT -205.085 -70.385 -204.685 -70.035 ;
        RECT -200.605 -70.385 -200.205 -70.035 ;
        RECT -196.125 -70.385 -195.725 -70.035 ;
        RECT -191.645 -70.385 -191.245 -70.035 ;
        RECT -186.045 -70.385 -185.645 -70.035 ;
        RECT -181.565 -70.385 -181.165 -70.035 ;
        RECT -177.085 -70.385 -176.685 -70.035 ;
        RECT -172.605 -70.385 -172.205 -70.035 ;
        RECT -168.125 -70.385 -167.725 -70.035 ;
        RECT -163.645 -70.385 -163.245 -70.035 ;
        RECT -159.165 -70.385 -158.765 -70.035 ;
        RECT -154.685 -70.385 -154.285 -70.035 ;
        RECT -150.205 -70.385 -149.805 -70.035 ;
        RECT -145.725 -70.385 -145.325 -70.035 ;
        RECT -141.245 -70.385 -140.845 -70.035 ;
        RECT -136.765 -70.385 -136.365 -70.035 ;
        RECT -132.285 -70.385 -131.885 -70.035 ;
        RECT -127.805 -70.385 -127.405 -70.035 ;
        RECT -123.325 -70.385 -122.925 -70.035 ;
        RECT -118.845 -70.385 -118.445 -70.035 ;
        RECT -114.365 -70.385 -113.965 -70.035 ;
        RECT -109.885 -70.385 -109.485 -70.035 ;
        RECT -105.405 -70.385 -105.005 -70.035 ;
        RECT -100.925 -70.385 -100.525 -70.035 ;
        RECT -96.445 -70.385 -96.045 -70.035 ;
        RECT -91.965 -70.385 -91.565 -70.035 ;
        RECT -87.485 -70.385 -87.085 -70.035 ;
        RECT -83.005 -70.385 -82.605 -70.035 ;
        RECT -78.525 -70.385 -78.125 -70.035 ;
        RECT -74.045 -70.385 -73.645 -70.035 ;
        RECT -69.565 -70.385 -69.165 -70.035 ;
        RECT -65.085 -70.385 -64.685 -70.035 ;
        RECT -60.605 -70.385 -60.205 -70.035 ;
        RECT -56.125 -70.385 -55.725 -70.035 ;
        RECT -51.645 -70.385 -51.245 -70.035 ;
        RECT -47.165 -70.385 -46.765 -70.035 ;
        RECT -42.685 -70.385 -42.285 -70.035 ;
        RECT -38.205 -70.385 -37.805 -70.035 ;
        RECT -33.725 -70.385 -33.325 -70.035 ;
        RECT -29.245 -70.385 -28.845 -70.035 ;
        RECT -24.765 -70.385 -24.365 -70.035 ;
        RECT -20.285 -70.385 -19.885 -70.035 ;
        RECT -15.805 -70.385 -15.405 -70.035 ;
        RECT -11.325 -70.385 -10.925 -70.035 ;
        RECT -6.845 -70.385 -6.445 -70.035 ;
        RECT -2.365 -70.385 -1.965 -70.035 ;
        RECT 2.115 -70.385 2.515 -70.035 ;
        RECT 6.595 -70.385 6.995 -70.035 ;
        RECT 11.075 -70.385 11.475 -70.035 ;
        RECT 15.555 -70.385 15.955 -70.035 ;
        RECT 20.035 -70.385 20.435 -70.035 ;
        RECT 24.515 -70.385 24.915 -70.035 ;
        RECT 28.995 -70.385 29.395 -70.035 ;
        RECT 33.475 -70.385 33.875 -70.035 ;
        RECT 37.955 -70.385 38.355 -70.035 ;
        RECT 42.435 -70.385 42.835 -70.035 ;
        RECT 46.915 -70.385 47.315 -70.035 ;
        RECT 51.395 -70.385 51.795 -70.035 ;
        RECT 55.875 -70.385 56.275 -70.035 ;
        RECT 60.355 -70.385 60.755 -70.035 ;
        RECT 64.835 -70.385 65.235 -70.035 ;
        RECT 69.315 -70.385 69.715 -70.035 ;
        RECT 73.795 -70.385 74.195 -70.035 ;
        RECT 78.275 -70.385 78.675 -70.035 ;
        RECT 82.755 -70.385 83.155 -70.035 ;
        RECT 87.235 -70.385 87.635 -70.035 ;
        RECT 91.715 -70.385 92.115 -70.035 ;
        RECT 96.195 -70.385 96.595 -70.035 ;
        RECT -473.885 -70.885 121.925 -70.385 ;
        RECT -473.885 -71.235 -473.485 -70.885 ;
        RECT -469.405 -71.235 -469.005 -70.885 ;
        RECT -464.925 -71.235 -464.525 -70.885 ;
        RECT -460.445 -71.235 -460.045 -70.885 ;
        RECT -455.965 -71.235 -455.565 -70.885 ;
        RECT -451.485 -71.235 -451.085 -70.885 ;
        RECT -447.005 -71.235 -446.605 -70.885 ;
        RECT -442.525 -71.235 -442.125 -70.885 ;
        RECT -438.045 -71.235 -437.645 -70.885 ;
        RECT -433.565 -71.235 -433.165 -70.885 ;
        RECT -429.085 -71.235 -428.685 -70.885 ;
        RECT -424.605 -71.235 -424.205 -70.885 ;
        RECT -420.125 -71.235 -419.725 -70.885 ;
        RECT -415.645 -71.235 -415.245 -70.885 ;
        RECT -411.165 -71.235 -410.765 -70.885 ;
        RECT -406.685 -71.235 -406.285 -70.885 ;
        RECT -402.205 -71.235 -401.805 -70.885 ;
        RECT -397.725 -71.235 -397.325 -70.885 ;
        RECT -393.245 -71.235 -392.845 -70.885 ;
        RECT -388.765 -71.235 -388.365 -70.885 ;
        RECT -384.285 -71.235 -383.885 -70.885 ;
        RECT -379.805 -71.235 -379.405 -70.885 ;
        RECT -375.325 -71.235 -374.925 -70.885 ;
        RECT -370.845 -71.235 -370.445 -70.885 ;
        RECT -366.365 -71.235 -365.965 -70.885 ;
        RECT -361.885 -71.235 -361.485 -70.885 ;
        RECT -357.405 -71.235 -357.005 -70.885 ;
        RECT -352.925 -71.235 -352.525 -70.885 ;
        RECT -348.445 -71.235 -348.045 -70.885 ;
        RECT -343.965 -71.235 -343.565 -70.885 ;
        RECT -339.485 -71.235 -339.085 -70.885 ;
        RECT -335.005 -71.235 -334.605 -70.885 ;
        RECT -330.525 -71.235 -330.125 -70.885 ;
        RECT -326.045 -71.235 -325.645 -70.885 ;
        RECT -321.565 -71.235 -321.165 -70.885 ;
        RECT -317.085 -71.235 -316.685 -70.885 ;
        RECT -312.605 -71.235 -312.205 -70.885 ;
        RECT -308.125 -71.235 -307.725 -70.885 ;
        RECT -303.645 -71.235 -303.245 -70.885 ;
        RECT -299.165 -71.235 -298.765 -70.885 ;
        RECT -294.685 -71.235 -294.285 -70.885 ;
        RECT -290.205 -71.235 -289.805 -70.885 ;
        RECT -285.725 -71.235 -285.325 -70.885 ;
        RECT -281.245 -71.235 -280.845 -70.885 ;
        RECT -276.765 -71.235 -276.365 -70.885 ;
        RECT -272.285 -71.235 -271.885 -70.885 ;
        RECT -267.805 -71.235 -267.405 -70.885 ;
        RECT -263.325 -71.235 -262.925 -70.885 ;
        RECT -258.845 -71.235 -258.445 -70.885 ;
        RECT -254.365 -71.235 -253.965 -70.885 ;
        RECT -249.885 -71.235 -249.485 -70.885 ;
        RECT -245.405 -71.235 -245.005 -70.885 ;
        RECT -240.925 -71.235 -240.525 -70.885 ;
        RECT -236.445 -71.235 -236.045 -70.885 ;
        RECT -231.965 -71.235 -231.565 -70.885 ;
        RECT -227.485 -71.235 -227.085 -70.885 ;
        RECT -223.005 -71.235 -222.605 -70.885 ;
        RECT -218.525 -71.235 -218.125 -70.885 ;
        RECT -214.045 -71.235 -213.645 -70.885 ;
        RECT -209.565 -71.235 -209.165 -70.885 ;
        RECT -205.085 -71.235 -204.685 -70.885 ;
        RECT -200.605 -71.235 -200.205 -70.885 ;
        RECT -196.125 -71.235 -195.725 -70.885 ;
        RECT -191.645 -71.235 -191.245 -70.885 ;
        RECT -186.045 -71.235 -185.645 -70.885 ;
        RECT -181.565 -71.235 -181.165 -70.885 ;
        RECT -177.085 -71.235 -176.685 -70.885 ;
        RECT -172.605 -71.235 -172.205 -70.885 ;
        RECT -168.125 -71.235 -167.725 -70.885 ;
        RECT -163.645 -71.235 -163.245 -70.885 ;
        RECT -159.165 -71.235 -158.765 -70.885 ;
        RECT -154.685 -71.235 -154.285 -70.885 ;
        RECT -150.205 -71.235 -149.805 -70.885 ;
        RECT -145.725 -71.235 -145.325 -70.885 ;
        RECT -141.245 -71.235 -140.845 -70.885 ;
        RECT -136.765 -71.235 -136.365 -70.885 ;
        RECT -132.285 -71.235 -131.885 -70.885 ;
        RECT -127.805 -71.235 -127.405 -70.885 ;
        RECT -123.325 -71.235 -122.925 -70.885 ;
        RECT -118.845 -71.235 -118.445 -70.885 ;
        RECT -114.365 -71.235 -113.965 -70.885 ;
        RECT -109.885 -71.235 -109.485 -70.885 ;
        RECT -105.405 -71.235 -105.005 -70.885 ;
        RECT -100.925 -71.235 -100.525 -70.885 ;
        RECT -96.445 -71.235 -96.045 -70.885 ;
        RECT -91.965 -71.235 -91.565 -70.885 ;
        RECT -87.485 -71.235 -87.085 -70.885 ;
        RECT -83.005 -71.235 -82.605 -70.885 ;
        RECT -78.525 -71.235 -78.125 -70.885 ;
        RECT -74.045 -71.235 -73.645 -70.885 ;
        RECT -69.565 -71.235 -69.165 -70.885 ;
        RECT -65.085 -71.235 -64.685 -70.885 ;
        RECT -60.605 -71.235 -60.205 -70.885 ;
        RECT -56.125 -71.235 -55.725 -70.885 ;
        RECT -51.645 -71.235 -51.245 -70.885 ;
        RECT -47.165 -71.235 -46.765 -70.885 ;
        RECT -42.685 -71.235 -42.285 -70.885 ;
        RECT -38.205 -71.235 -37.805 -70.885 ;
        RECT -33.725 -71.235 -33.325 -70.885 ;
        RECT -29.245 -71.235 -28.845 -70.885 ;
        RECT -24.765 -71.235 -24.365 -70.885 ;
        RECT -20.285 -71.235 -19.885 -70.885 ;
        RECT -15.805 -71.235 -15.405 -70.885 ;
        RECT -11.325 -71.235 -10.925 -70.885 ;
        RECT -6.845 -71.235 -6.445 -70.885 ;
        RECT -2.365 -71.235 -1.965 -70.885 ;
        RECT 2.115 -71.235 2.515 -70.885 ;
        RECT 6.595 -71.235 6.995 -70.885 ;
        RECT 11.075 -71.235 11.475 -70.885 ;
        RECT 15.555 -71.235 15.955 -70.885 ;
        RECT 20.035 -71.235 20.435 -70.885 ;
        RECT 24.515 -71.235 24.915 -70.885 ;
        RECT 28.995 -71.235 29.395 -70.885 ;
        RECT 33.475 -71.235 33.875 -70.885 ;
        RECT 37.955 -71.235 38.355 -70.885 ;
        RECT 42.435 -71.235 42.835 -70.885 ;
        RECT 46.915 -71.235 47.315 -70.885 ;
        RECT 51.395 -71.235 51.795 -70.885 ;
        RECT 55.875 -71.235 56.275 -70.885 ;
        RECT 60.355 -71.235 60.755 -70.885 ;
        RECT 64.835 -71.235 65.235 -70.885 ;
        RECT 69.315 -71.235 69.715 -70.885 ;
        RECT 73.795 -71.235 74.195 -70.885 ;
        RECT 78.275 -71.235 78.675 -70.885 ;
        RECT 82.755 -71.235 83.155 -70.885 ;
        RECT 87.235 -71.235 87.635 -70.885 ;
        RECT 91.715 -71.235 92.115 -70.885 ;
        RECT 96.195 -71.235 96.595 -70.885 ;
        RECT -471.645 -73.745 -471.245 -73.395 ;
        RECT -462.685 -73.745 -462.285 -73.395 ;
        RECT -453.725 -73.745 -453.325 -73.395 ;
        RECT -444.765 -73.745 -444.365 -73.395 ;
        RECT -435.805 -73.745 -435.405 -73.395 ;
        RECT -426.845 -73.745 -426.445 -73.395 ;
        RECT -417.885 -73.745 -417.485 -73.395 ;
        RECT -408.925 -73.745 -408.525 -73.395 ;
        RECT -399.965 -73.745 -399.565 -73.395 ;
        RECT -391.005 -73.745 -390.605 -73.395 ;
        RECT -382.045 -73.745 -381.645 -73.395 ;
        RECT -373.085 -73.745 -372.685 -73.395 ;
        RECT -364.125 -73.745 -363.725 -73.395 ;
        RECT -355.165 -73.745 -354.765 -73.395 ;
        RECT -346.205 -73.745 -345.805 -73.395 ;
        RECT -337.245 -73.745 -336.845 -73.395 ;
        RECT -328.285 -73.745 -327.885 -73.395 ;
        RECT -319.325 -73.745 -318.925 -73.395 ;
        RECT -310.365 -73.745 -309.965 -73.395 ;
        RECT -301.405 -73.745 -301.005 -73.395 ;
        RECT -292.445 -73.745 -292.045 -73.395 ;
        RECT -283.485 -73.745 -283.085 -73.395 ;
        RECT -274.525 -73.745 -274.125 -73.395 ;
        RECT -265.565 -73.745 -265.165 -73.395 ;
        RECT -256.605 -73.745 -256.205 -73.395 ;
        RECT -247.645 -73.745 -247.245 -73.395 ;
        RECT -238.685 -73.745 -238.285 -73.395 ;
        RECT -229.725 -73.745 -229.325 -73.395 ;
        RECT -220.765 -73.745 -220.365 -73.395 ;
        RECT -211.805 -73.745 -211.405 -73.395 ;
        RECT -202.845 -73.745 -202.445 -73.395 ;
        RECT -193.885 -73.745 -193.485 -73.395 ;
        RECT -183.805 -73.745 -183.405 -73.395 ;
        RECT -174.845 -73.745 -174.445 -73.395 ;
        RECT -165.885 -73.745 -165.485 -73.395 ;
        RECT -156.925 -73.745 -156.525 -73.395 ;
        RECT -147.965 -73.745 -147.565 -73.395 ;
        RECT -139.005 -73.745 -138.605 -73.395 ;
        RECT -130.045 -73.745 -129.645 -73.395 ;
        RECT -121.085 -73.745 -120.685 -73.395 ;
        RECT -112.125 -73.745 -111.725 -73.395 ;
        RECT -103.165 -73.745 -102.765 -73.395 ;
        RECT -94.205 -73.745 -93.805 -73.395 ;
        RECT -85.245 -73.745 -84.845 -73.395 ;
        RECT -76.285 -73.745 -75.885 -73.395 ;
        RECT -67.325 -73.745 -66.925 -73.395 ;
        RECT -58.365 -73.745 -57.965 -73.395 ;
        RECT -49.405 -73.745 -49.005 -73.395 ;
        RECT -40.445 -73.745 -40.045 -73.395 ;
        RECT -31.485 -73.745 -31.085 -73.395 ;
        RECT -22.525 -73.745 -22.125 -73.395 ;
        RECT -13.565 -73.745 -13.165 -73.395 ;
        RECT -4.605 -73.745 -4.205 -73.395 ;
        RECT 4.355 -73.745 4.755 -73.395 ;
        RECT 13.315 -73.745 13.715 -73.395 ;
        RECT 22.275 -73.745 22.675 -73.395 ;
        RECT 31.235 -73.745 31.635 -73.395 ;
        RECT 40.195 -73.745 40.595 -73.395 ;
        RECT 49.155 -73.745 49.555 -73.395 ;
        RECT 58.115 -73.745 58.515 -73.395 ;
        RECT 67.075 -73.745 67.475 -73.395 ;
        RECT 76.035 -73.745 76.435 -73.395 ;
        RECT 84.995 -73.745 85.395 -73.395 ;
        RECT 93.955 -73.745 94.355 -73.395 ;
        RECT -471.645 -74.245 121.925 -73.745 ;
        RECT -471.645 -74.595 -471.245 -74.245 ;
        RECT -462.685 -74.595 -462.285 -74.245 ;
        RECT -453.725 -74.595 -453.325 -74.245 ;
        RECT -444.765 -74.595 -444.365 -74.245 ;
        RECT -435.805 -74.595 -435.405 -74.245 ;
        RECT -426.845 -74.595 -426.445 -74.245 ;
        RECT -417.885 -74.595 -417.485 -74.245 ;
        RECT -408.925 -74.595 -408.525 -74.245 ;
        RECT -399.965 -74.595 -399.565 -74.245 ;
        RECT -391.005 -74.595 -390.605 -74.245 ;
        RECT -382.045 -74.595 -381.645 -74.245 ;
        RECT -373.085 -74.595 -372.685 -74.245 ;
        RECT -364.125 -74.595 -363.725 -74.245 ;
        RECT -355.165 -74.595 -354.765 -74.245 ;
        RECT -346.205 -74.595 -345.805 -74.245 ;
        RECT -337.245 -74.595 -336.845 -74.245 ;
        RECT -328.285 -74.595 -327.885 -74.245 ;
        RECT -319.325 -74.595 -318.925 -74.245 ;
        RECT -310.365 -74.595 -309.965 -74.245 ;
        RECT -301.405 -74.595 -301.005 -74.245 ;
        RECT -292.445 -74.595 -292.045 -74.245 ;
        RECT -283.485 -74.595 -283.085 -74.245 ;
        RECT -274.525 -74.595 -274.125 -74.245 ;
        RECT -265.565 -74.595 -265.165 -74.245 ;
        RECT -256.605 -74.595 -256.205 -74.245 ;
        RECT -247.645 -74.595 -247.245 -74.245 ;
        RECT -238.685 -74.595 -238.285 -74.245 ;
        RECT -229.725 -74.595 -229.325 -74.245 ;
        RECT -220.765 -74.595 -220.365 -74.245 ;
        RECT -211.805 -74.595 -211.405 -74.245 ;
        RECT -202.845 -74.595 -202.445 -74.245 ;
        RECT -193.885 -74.595 -193.485 -74.245 ;
        RECT -183.805 -74.595 -183.405 -74.245 ;
        RECT -174.845 -74.595 -174.445 -74.245 ;
        RECT -165.885 -74.595 -165.485 -74.245 ;
        RECT -156.925 -74.595 -156.525 -74.245 ;
        RECT -147.965 -74.595 -147.565 -74.245 ;
        RECT -139.005 -74.595 -138.605 -74.245 ;
        RECT -130.045 -74.595 -129.645 -74.245 ;
        RECT -121.085 -74.595 -120.685 -74.245 ;
        RECT -112.125 -74.595 -111.725 -74.245 ;
        RECT -103.165 -74.595 -102.765 -74.245 ;
        RECT -94.205 -74.595 -93.805 -74.245 ;
        RECT -85.245 -74.595 -84.845 -74.245 ;
        RECT -76.285 -74.595 -75.885 -74.245 ;
        RECT -67.325 -74.595 -66.925 -74.245 ;
        RECT -58.365 -74.595 -57.965 -74.245 ;
        RECT -49.405 -74.595 -49.005 -74.245 ;
        RECT -40.445 -74.595 -40.045 -74.245 ;
        RECT -31.485 -74.595 -31.085 -74.245 ;
        RECT -22.525 -74.595 -22.125 -74.245 ;
        RECT -13.565 -74.595 -13.165 -74.245 ;
        RECT -4.605 -74.595 -4.205 -74.245 ;
        RECT 4.355 -74.595 4.755 -74.245 ;
        RECT 13.315 -74.595 13.715 -74.245 ;
        RECT 22.275 -74.595 22.675 -74.245 ;
        RECT 31.235 -74.595 31.635 -74.245 ;
        RECT 40.195 -74.595 40.595 -74.245 ;
        RECT 49.155 -74.595 49.555 -74.245 ;
        RECT 58.115 -74.595 58.515 -74.245 ;
        RECT 67.075 -74.595 67.475 -74.245 ;
        RECT 76.035 -74.595 76.435 -74.245 ;
        RECT 84.995 -74.595 85.395 -74.245 ;
        RECT 93.955 -74.595 94.355 -74.245 ;
        RECT -467.165 -77.105 -466.765 -76.755 ;
        RECT -449.245 -77.105 -448.845 -76.755 ;
        RECT -431.325 -77.105 -430.925 -76.755 ;
        RECT -413.405 -77.105 -413.005 -76.755 ;
        RECT -395.485 -77.105 -395.085 -76.755 ;
        RECT -377.565 -77.105 -377.165 -76.755 ;
        RECT -359.645 -77.105 -359.245 -76.755 ;
        RECT -341.725 -77.105 -341.325 -76.755 ;
        RECT -323.805 -77.105 -323.405 -76.755 ;
        RECT -305.885 -77.105 -305.485 -76.755 ;
        RECT -287.965 -77.105 -287.565 -76.755 ;
        RECT -270.045 -77.105 -269.645 -76.755 ;
        RECT -252.125 -77.105 -251.725 -76.755 ;
        RECT -234.205 -77.105 -233.805 -76.755 ;
        RECT -216.285 -77.105 -215.885 -76.755 ;
        RECT -198.365 -77.105 -197.965 -76.755 ;
        RECT -179.325 -77.105 -178.925 -76.755 ;
        RECT -161.405 -77.105 -161.005 -76.755 ;
        RECT -143.485 -77.105 -143.085 -76.755 ;
        RECT -125.565 -77.105 -125.165 -76.755 ;
        RECT -107.645 -77.105 -107.245 -76.755 ;
        RECT -89.725 -77.105 -89.325 -76.755 ;
        RECT -71.805 -77.105 -71.405 -76.755 ;
        RECT -53.885 -77.105 -53.485 -76.755 ;
        RECT -35.965 -77.105 -35.565 -76.755 ;
        RECT -18.045 -77.105 -17.645 -76.755 ;
        RECT -0.125 -77.105 0.275 -76.755 ;
        RECT 17.795 -77.105 18.195 -76.755 ;
        RECT 35.715 -77.105 36.115 -76.755 ;
        RECT 53.635 -77.105 54.035 -76.755 ;
        RECT 71.555 -77.105 71.955 -76.755 ;
        RECT 89.475 -77.105 89.875 -76.755 ;
        RECT -467.165 -77.605 121.925 -77.105 ;
        RECT -467.165 -77.955 -466.765 -77.605 ;
        RECT -449.245 -77.955 -448.845 -77.605 ;
        RECT -431.325 -77.955 -430.925 -77.605 ;
        RECT -413.405 -77.955 -413.005 -77.605 ;
        RECT -395.485 -77.955 -395.085 -77.605 ;
        RECT -377.565 -77.955 -377.165 -77.605 ;
        RECT -359.645 -77.955 -359.245 -77.605 ;
        RECT -341.725 -77.955 -341.325 -77.605 ;
        RECT -323.805 -77.955 -323.405 -77.605 ;
        RECT -305.885 -77.955 -305.485 -77.605 ;
        RECT -287.965 -77.955 -287.565 -77.605 ;
        RECT -270.045 -77.955 -269.645 -77.605 ;
        RECT -252.125 -77.955 -251.725 -77.605 ;
        RECT -234.205 -77.955 -233.805 -77.605 ;
        RECT -216.285 -77.955 -215.885 -77.605 ;
        RECT -198.365 -77.955 -197.965 -77.605 ;
        RECT -179.325 -77.955 -178.925 -77.605 ;
        RECT -161.405 -77.955 -161.005 -77.605 ;
        RECT -143.485 -77.955 -143.085 -77.605 ;
        RECT -125.565 -77.955 -125.165 -77.605 ;
        RECT -107.645 -77.955 -107.245 -77.605 ;
        RECT -89.725 -77.955 -89.325 -77.605 ;
        RECT -71.805 -77.955 -71.405 -77.605 ;
        RECT -53.885 -77.955 -53.485 -77.605 ;
        RECT -35.965 -77.955 -35.565 -77.605 ;
        RECT -18.045 -77.955 -17.645 -77.605 ;
        RECT -0.125 -77.955 0.275 -77.605 ;
        RECT 17.795 -77.955 18.195 -77.605 ;
        RECT 35.715 -77.955 36.115 -77.605 ;
        RECT 53.635 -77.955 54.035 -77.605 ;
        RECT 71.555 -77.955 71.955 -77.605 ;
        RECT 89.475 -77.955 89.875 -77.605 ;
        RECT -497.305 -78.900 -486.905 -78.300 ;
        RECT -458.205 -80.465 -457.805 -80.115 ;
        RECT -422.365 -80.465 -421.965 -80.115 ;
        RECT -386.525 -80.465 -386.125 -80.115 ;
        RECT -350.685 -80.465 -350.285 -80.115 ;
        RECT -314.845 -80.465 -314.445 -80.115 ;
        RECT -279.005 -80.465 -278.605 -80.115 ;
        RECT -243.165 -80.465 -242.765 -80.115 ;
        RECT -207.325 -80.465 -206.925 -80.115 ;
        RECT -170.365 -80.465 -169.965 -80.115 ;
        RECT -134.525 -80.465 -134.125 -80.115 ;
        RECT -98.685 -80.465 -98.285 -80.115 ;
        RECT -62.845 -80.465 -62.445 -80.115 ;
        RECT -27.005 -80.465 -26.605 -80.115 ;
        RECT 8.835 -80.465 9.235 -80.115 ;
        RECT 44.675 -80.465 45.075 -80.115 ;
        RECT 80.515 -80.465 80.915 -80.115 ;
        RECT -458.205 -80.965 121.925 -80.465 ;
        RECT -486.955 -83.235 -486.555 -81.155 ;
        RECT -458.205 -81.315 -457.805 -80.965 ;
        RECT -422.365 -81.315 -421.965 -80.965 ;
        RECT -386.525 -81.315 -386.125 -80.965 ;
        RECT -350.685 -81.315 -350.285 -80.965 ;
        RECT -314.845 -81.315 -314.445 -80.965 ;
        RECT -279.005 -81.315 -278.605 -80.965 ;
        RECT -243.165 -81.315 -242.765 -80.965 ;
        RECT -207.325 -81.315 -206.925 -80.965 ;
        RECT -170.365 -81.315 -169.965 -80.965 ;
        RECT -134.525 -81.315 -134.125 -80.965 ;
        RECT -98.685 -81.315 -98.285 -80.965 ;
        RECT -62.845 -81.315 -62.445 -80.965 ;
        RECT -27.005 -81.315 -26.605 -80.965 ;
        RECT 8.835 -81.315 9.235 -80.965 ;
        RECT 44.675 -81.315 45.075 -80.965 ;
        RECT 80.515 -81.315 80.915 -80.965 ;
        RECT -497.595 -83.765 -495.515 -83.365 ;
        RECT -440.285 -83.825 -439.885 -83.475 ;
        RECT -368.605 -83.825 -368.205 -83.475 ;
        RECT -296.925 -83.825 -296.525 -83.475 ;
        RECT -225.245 -83.825 -224.845 -83.475 ;
        RECT -152.445 -83.825 -152.045 -83.475 ;
        RECT -80.765 -83.825 -80.365 -83.475 ;
        RECT -9.085 -83.825 -8.685 -83.475 ;
        RECT 62.595 -83.825 62.995 -83.475 ;
        RECT -440.285 -84.325 121.925 -83.825 ;
        RECT -440.285 -84.675 -439.885 -84.325 ;
        RECT -368.605 -84.675 -368.205 -84.325 ;
        RECT -296.925 -84.675 -296.525 -84.325 ;
        RECT -225.245 -84.675 -224.845 -84.325 ;
        RECT -152.445 -84.675 -152.045 -84.325 ;
        RECT -80.765 -84.675 -80.365 -84.325 ;
        RECT -9.085 -84.675 -8.685 -84.325 ;
        RECT 62.595 -84.675 62.995 -84.325 ;
        RECT -404.445 -87.185 -404.045 -86.835 ;
        RECT -261.085 -87.185 -260.685 -86.835 ;
        RECT -116.605 -87.185 -116.205 -86.835 ;
        RECT 26.755 -87.185 27.155 -86.835 ;
        RECT -404.445 -87.685 121.925 -87.185 ;
        RECT -404.445 -88.035 -404.045 -87.685 ;
        RECT -261.085 -88.035 -260.685 -87.685 ;
        RECT -116.605 -88.035 -116.205 -87.685 ;
        RECT 26.755 -88.035 27.155 -87.685 ;
        RECT -332.765 -90.545 -332.365 -90.195 ;
        RECT -44.925 -90.545 -44.525 -90.195 ;
        RECT -332.765 -91.045 121.925 -90.545 ;
        RECT -332.765 -91.395 -332.365 -91.045 ;
        RECT -44.925 -91.395 -44.525 -91.045 ;
        RECT -188.285 -93.905 -187.885 -93.555 ;
        RECT -188.285 -94.405 121.925 -93.905 ;
        RECT -188.285 -94.755 -187.885 -94.405 ;
        RECT -189.405 -97.265 -189.005 -96.915 ;
        RECT -189.405 -97.765 121.925 -97.265 ;
        RECT -189.405 -98.115 -189.005 -97.765 ;
        RECT 239.520 -117.620 243.520 -5.865 ;
        RECT 389.020 -14.510 389.300 -5.730 ;
        RECT 389.580 -13.950 389.860 0.990 ;
        RECT 385.660 -17.310 385.940 -14.690 ;
      LAYER Via4 ;
        RECT -497.475 83.425 -495.635 83.705 ;
        RECT -486.895 81.275 -486.615 83.115 ;
        RECT -496.915 70.260 -496.635 78.340 ;
        RECT -496.915 58.260 -496.635 66.340 ;
        RECT -496.915 46.260 -496.635 54.340 ;
        RECT -496.915 34.260 -496.635 42.340 ;
        RECT -496.915 22.260 -496.635 30.340 ;
        RECT -496.915 -30.340 -496.635 -22.260 ;
        RECT -496.915 -42.340 -496.635 -34.260 ;
        RECT -496.915 -54.340 -496.635 -46.260 ;
        RECT -496.915 -66.340 -496.635 -58.260 ;
        RECT -496.915 -78.340 -496.635 -70.260 ;
        RECT -486.895 -83.115 -486.615 -81.275 ;
        RECT -497.475 -83.705 -495.635 -83.425 ;
      LAYER Metal5 ;
        RECT -806.980 -450.000 -791.980 450.000 ;
        RECT -622.500 430.200 -607.500 976.200 ;
        RECT 607.500 430.200 622.500 976.200 ;
        RECT -497.595 83.315 -495.515 83.815 ;
        RECT -497.595 21.985 -496.555 83.315 ;
        RECT -487.105 78.615 -486.405 83.235 ;
        RECT -488.405 77.940 -486.405 78.615 ;
        RECT -495.145 70.660 -486.405 77.940 ;
        RECT -488.405 65.940 -486.405 70.660 ;
        RECT -495.145 58.660 -486.405 65.940 ;
        RECT -488.405 53.940 -486.405 58.660 ;
        RECT -495.145 46.660 -486.405 53.940 ;
        RECT -488.405 41.940 -486.405 46.660 ;
        RECT -495.145 34.660 -486.405 41.940 ;
        RECT -488.405 29.940 -486.405 34.660 ;
        RECT -495.145 22.660 -486.405 29.940 ;
        RECT -488.405 21.985 -486.405 22.660 ;
        RECT -497.595 -83.315 -496.555 -21.985 ;
        RECT -488.405 -22.660 -486.405 -21.985 ;
        RECT -495.145 -29.940 -486.405 -22.660 ;
        RECT -488.405 -34.660 -486.405 -29.940 ;
        RECT -495.145 -41.940 -486.405 -34.660 ;
        RECT -488.405 -46.660 -486.405 -41.940 ;
        RECT -495.145 -53.940 -486.405 -46.660 ;
        RECT -488.405 -58.660 -486.405 -53.940 ;
        RECT -495.145 -65.940 -486.405 -58.660 ;
        RECT -488.405 -70.660 -486.405 -65.940 ;
        RECT -495.145 -77.940 -486.405 -70.660 ;
        RECT -488.405 -78.615 -486.405 -77.940 ;
        RECT -487.105 -83.235 -486.405 -78.615 ;
        RECT -497.595 -83.815 -495.515 -83.315 ;
        RECT -622.500 -976.200 -607.500 -430.200 ;
        RECT 607.500 -976.200 622.500 -430.200 ;
        RECT 794.820 -450.000 809.820 450.000 ;
  END
END saradc
END LIBRARY

