* NGSPICE file created from carray_3.ext - technology: gf180mcuD

.subckt carray_3 carray_out n9 n0 n8 n7 n6 n5 n4 n3 n2 n1 ndum
C0 carray_out ndum 1.65633f
C1 n3 n6 0.618871f
C2 n7 carray_out 0.21201p
C3 n7 n3 1.41554f
C4 n4 n2 0.351771f
C5 n4 n6 1.16683f
C6 n2 n6 0.349007f
C7 n4 n7 2.75193f
C8 n1 n0 8.760937f
C9 n7 n2 0.747257f
C10 n1 carray_out 3.31266f
C11 n7 n6 38.4269f
C12 n7 ndum 0.108702f
C13 n1 n3 0.203114f
C14 n0 n9 0.238827f
C15 carray_out n9 0.853823p
C16 n5 carray_out 53.002514f
C17 n3 n9 2.561274f
C18 n4 n1 0.201445f
C19 n5 n3 0.623459f
C20 n0 n8 0.153648f
C21 n1 n2 16.6626f
C22 n1 n6 0.20118f
C23 carray_out n8 0.424139p
C24 n1 ndum 8.453368f
C25 n1 n7 0.301117f
C26 n8 n3 2.12966f
C27 n4 n9 5.040546f
C28 n4 n5 28.0344f
C29 n2 n9 1.321566f
C30 n5 n2 0.349129f
C31 n6 n9 19.91684f
C32 ndum n9 0.181793f
C33 n5 n6 29.673302f
C34 n7 n9 39.81507f
C35 n4 n8 4.18035f
C36 n7 n5 5.44073f
C37 n2 n8 1.10439f
C38 n8 n6 16.515598f
C39 n8 ndum 0.153648f
C40 n7 n8 60.691196f
C41 n0 carray_out 1.65633f
C42 n1 n9 0.450074f
C43 n1 n5 0.201323f
C44 carray_out n3 13.250643f
C45 n1 n8 0.391009f
C46 n5 n9 9.999403f
C47 n0 n2 0.131408f
C48 n4 carray_out 26.501268f
C49 n8 n9 0.107528p
C50 carray_out n2 6.625319f
C51 n4 n3 26.1647f
C52 n5 n8 8.28156f
C53 carray_out n6 0.106005p
C54 n0 n7 0.108702f
C55 n2 n3 22.977001f
C56 ndum VSUBS 13.371039f
C57 n8 VSUBS 59.384502f
C58 n7 VSUBS 56.43133f
C59 n4 VSUBS 37.69574f
C60 carray_out VSUBS 81.95506f
C61 n5 VSUBS 44.915176f
C62 n6 VSUBS 52.011745f
C63 n9 VSUBS 81.5176f
C64 n3 VSUBS 32.19483f
C65 n0 VSUBS 16.058037f
C66 n2 VSUBS 29.061958f
C67 n1 VSUBS 16.015188f
.ends

