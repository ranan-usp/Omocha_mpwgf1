VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.920 ;
  SYMMETRY X Y ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.711500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.858000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.770 0.810 16.350 2.985 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 16.800 4.220 ;
        RECT 1.440 2.930 1.780 3.620 ;
        RECT 3.180 3.005 3.520 3.620 ;
        RECT 7.705 2.700 8.045 3.620 ;
        RECT 12.850 3.280 13.190 3.620 ;
        RECT 14.845 2.755 15.185 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 17.230 4.350 ;
        RECT -0.430 1.760 7.265 1.885 ;
        RECT 14.620 1.760 17.230 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 7.265 1.760 14.620 1.885 ;
        RECT -0.430 -0.430 17.230 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.300 1.780 0.915 ;
        RECT 3.280 0.300 3.620 1.075 ;
        RECT 7.700 0.300 8.040 0.810 ;
        RECT 12.720 0.300 13.060 0.950 ;
        RECT 15.000 0.300 15.230 0.690 ;
        RECT 0.000 -0.300 16.800 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.475 2.590 0.705 3.225 ;
        RECT 2.515 2.710 2.845 3.225 ;
        RECT 3.830 3.160 6.355 3.390 ;
        RECT 3.830 2.710 4.060 3.160 ;
        RECT 13.430 3.100 14.615 3.330 ;
        RECT 13.430 3.050 13.660 3.100 ;
        RECT 0.475 2.360 2.165 2.590 ;
        RECT 1.935 1.375 2.165 2.360 ;
        RECT 0.375 1.145 2.165 1.375 ;
        RECT 2.515 2.480 4.060 2.710 ;
        RECT 4.420 2.645 5.290 2.875 ;
        RECT 0.375 0.735 0.605 1.145 ;
        RECT 2.515 0.735 2.845 2.480 ;
        RECT 5.055 1.075 5.290 2.645 ;
        RECT 4.400 0.845 5.290 1.075 ;
        RECT 5.575 2.050 5.915 2.795 ;
        RECT 9.040 2.390 9.380 2.930 ;
        RECT 7.095 2.050 9.380 2.390 ;
        RECT 5.575 1.820 6.780 2.050 ;
        RECT 5.575 0.790 5.805 1.820 ;
        RECT 6.550 1.730 6.780 1.820 ;
        RECT 6.090 1.270 6.320 1.590 ;
        RECT 6.550 1.500 8.700 1.730 ;
        RECT 6.090 1.040 8.560 1.270 ;
        RECT 8.330 0.760 8.560 1.040 ;
        RECT 9.040 0.990 9.380 2.050 ;
        RECT 10.160 2.585 10.500 2.930 ;
        RECT 11.790 2.815 13.660 3.050 ;
        RECT 10.160 2.355 13.630 2.585 ;
        RECT 10.160 0.990 10.500 2.355 ;
        RECT 13.290 2.105 13.630 2.355 ;
        RECT 11.195 0.760 11.425 2.095 ;
        RECT 13.925 1.885 14.155 2.850 ;
        RECT 14.385 2.345 14.615 3.100 ;
        RECT 14.385 2.115 15.460 2.345 ;
        RECT 13.925 1.875 15.000 1.885 ;
        RECT 12.175 1.640 15.000 1.875 ;
        RECT 13.900 1.500 15.000 1.640 ;
        RECT 11.655 1.180 13.520 1.410 ;
        RECT 11.655 0.890 11.885 1.180 ;
        RECT 8.330 0.530 11.425 0.760 ;
        RECT 13.290 0.760 13.520 1.180 ;
        RECT 13.900 0.990 14.240 1.500 ;
        RECT 15.230 1.150 15.460 2.115 ;
        RECT 14.540 0.920 15.460 1.150 ;
        RECT 14.540 0.760 14.770 0.920 ;
        RECT 13.290 0.530 14.770 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_1
END LIBRARY