* NGSPICE file created from dac_in.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8$1 Z I VDD VSS VPW VNW VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS VPW VNW VSUBS
X0 a_4604_375# a_4516_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3 a_4156_375# a_4068_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 a_5500_375# a_5412_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 VDD a_5052_375# a_4964_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 VDD a_6844_375# a_6756_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 a_5052_375# a_4964_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X11 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_4604_375# a_4516_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X14 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X15 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X16 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X17 a_5948_375# a_5860_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X18 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X19 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X20 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X21 VDD a_5500_375# a_5412_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X22 a_6844_375# a_6756_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X23 a_6396_375# a_6308_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X24 VDD a_6396_375# a_6308_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X25 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X26 VDD a_4156_375# a_4068_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X27 VDD a_5948_375# a_5860_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X28 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X29 a_3708_375# a_3620_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X30 VDD a_3708_375# a_3620_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X31 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna$1 VSS I VDD VPW VNW VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1 VDD VSS VPW VNW VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1 VDD VSS VPW VNW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1$1 VSS ZN I VDD VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1 VSS Z I VDD VPW VNW VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1$1 VSS Z I VDD VPW VNW VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt phase_inverter input_signal[0] input_signal[1] input_signal[2] input_signal[3]
+ input_signal[4] input_signal[5] input_signal[9] output_signal_minus[0] output_signal_minus[1]
+ output_signal_minus[2] output_signal_minus[3] output_signal_minus[4] output_signal_minus[5]
+ output_signal_minus[6] output_signal_minus[7] output_signal_minus[8] output_signal_minus[9]
+ output_signal_plus[0] output_signal_plus[1] output_signal_plus[2] output_signal_plus[3]
+ output_signal_plus[4] output_signal_plus[5] output_signal_plus[6] output_signal_plus[7]
+ output_signal_plus[8] output_signal_plus[9] input_signal[7] input_signal[8] input_signal[6]
+ vdd vss
XFILLER_0_1_72 vdd vss FILLER_0_1_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput20 output_signal_minus[9] _00_/ZN vdd vss output20/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput21 output_signal_plus[0] _10_/Z vdd vss output21/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_9_2 vdd vss FILLER_0_9_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_72 vdd vss FILLER_0_7_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XANTENNA_input3_I vss input_signal[2] vdd ANTENNA_input3_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
Xoutput22 output_signal_plus[1] _11_/Z vdd vss output22/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput11 output_signal_minus[0] _01_/ZN vdd vss output11/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput23 output_signal_plus[2] _12_/Z vdd vss output23/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_12_101 vdd vss FILLER_0_12_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xoutput12 output_signal_minus[1] _02_/ZN vdd vss output12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_13_66 vdd vss FILLER_0_13_66/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_10_12 vdd vss FILLER_0_10_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_8_107 vdd vss FILLER_0_8_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
Xoutput24 output_signal_plus[3] _13_/Z vdd vss output24/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput13 output_signal_minus[2] _03_/ZN vdd vss output13/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_7_2 vdd vss FILLER_0_7_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I vss input_signal[0] vdd ANTENNA_input1_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_1_44 vdd vss FILLER_0_1_44/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput25 output_signal_plus[4] _14_/Z vdd vss output25/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput14 output_signal_minus[3] _04_/ZN vdd vss output14/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_1_12 vdd vss FILLER_0_1_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_09_ vss _09_/ZN _18_/I vdd _09_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xoutput26 output_signal_plus[5] _15_/Z vdd vss output26/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_4_101 vdd vss FILLER_0_4_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xoutput15 output_signal_minus[4] net15 vdd vss output15/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_7_66 vdd vss FILLER_0_7_66/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_10_37 vdd vss FILLER_0_10_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08_ vss _08_/ZN _17_/I vdd _08_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
XFILLER_0_16_36 vdd vss FILLER_0_16_36/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xoutput27 output_signal_plus[6] _16_/Z vdd vss output27/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput16 output_signal_minus[5] _06_/ZN vdd vss output16/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_07_ vss _07_/ZN _16_/I vdd _07_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xoutput28 output_signal_plus[7] _17_/Z vdd vss output28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput17 output_signal_minus[6] _07_/ZN vdd vss output17/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XFILLER_0_10_28 vdd vss FILLER_0_10_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_12_107 vdd vss FILLER_0_12_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xoutput29 output_signal_plus[8] _18_/Z vdd vss output29/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
Xoutput18 output_signal_minus[7] _08_/ZN vdd vss output18/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
X_06_ vdd vss _15_/I _06_/ZN _06_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
XFILLER_0_4_37 vdd vss FILLER_0_4_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_72 vdd vss FILLER_0_11_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05_ vdd vss _14_/I net15 _05_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
Xoutput19 output_signal_minus[8] _09_/ZN vdd vss output19/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XANTENNA__04__I vss _13_/I vdd ANTENNA__04__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_16_18 vdd vss FILLER_0_16_18/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XANTENNA__15__I vss _15_/I vdd ANTENNA__15__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XANTENNA_input8_I vss input_signal[7] vdd ANTENNA_input8_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
X_04_ vdd vss _13_/I _04_/ZN _04_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
XFILLER_0_0_142 vdd vss FILLER_0_0_142/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_5_60 vdd vss FILLER_0_5_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
Xinput1 vss _10_/I input_signal[0] vdd input1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_7_104 vdd vss FILLER_0_7_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_03_ vdd vss _12_/I _03_/ZN _03_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
XFILLER_0_4_107 vdd vss FILLER_0_4_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_5_72 vdd vss FILLER_0_5_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xinput2 vss _11_/I input_signal[1] vdd input2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
X_02_ vdd vss _11_/I _02_/ZN _02_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
X_01_ vdd vss _10_/I _01_/ZN _01_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1$1
Xinput3 vss _12_/I input_signal[2] vdd input3/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA_input6_I vss input_signal[5] vdd ANTENNA_input6_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_11_66 vdd vss FILLER_0_11_66/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xinput4 vss _13_/I input_signal[3] vdd input4/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
X_00_ vss _00_/ZN _19_/I vdd _00_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1$1
Xinput5 vss _14_/I input_signal[4] vdd input5/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_11_136 vdd vss FILLER_0_11_136/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_14_12 vdd vss FILLER_0_14_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_14_101 vdd vss FILLER_0_14_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xinput6 vss _15_/I input_signal[5] vdd input6/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_0_104 vdd vss FILLER_0_0_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA_input4_I vss input_signal[3] vdd ANTENNA_input4_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
Xinput7 vss _16_/I input_signal[6] vdd input7/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_5_44 vdd vss FILLER_0_5_44/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
Xinput10 vss _19_/I input_signal[9] vdd input10/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_5_12 vdd vss FILLER_0_5_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
Xinput8 vss _17_/I input_signal[7] vdd input8/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_8_12 vdd vss FILLER_0_8_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_14_37 vdd vss FILLER_0_14_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_115 vdd vss FILLER_0_14_115/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
Xinput9 vss _18_/I input_signal[8] vdd input9/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_3_104 vdd vss FILLER_0_3_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_6_101 vdd vss FILLER_0_6_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA_input10_I vss input_signal[9] vdd ANTENNA_input10_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XANTENNA_input2_I vss input_signal[1] vdd ANTENNA_input2_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_2_37 vdd vss FILLER_0_2_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_28 vdd vss FILLER_0_14_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA__02__I vss _11_/I vdd ANTENNA__02__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_0_70 vdd vss FILLER_0_0_70/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_8_37 vdd vss FILLER_0_8_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_19_ vss _19_/Z _19_/I vdd _19_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA__05__I vss _14_/I vdd ANTENNA__05__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_15_72 vdd vss FILLER_0_15_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XANTENNA__13__I vss _13_/I vdd ANTENNA__13__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_14_107 vdd vss FILLER_0_14_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_3_60 vdd vss FILLER_0_3_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_18_ vss _18_/Z _18_/I vdd _18_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_40 vdd vss FILLER_0_15_40/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_6_2 vdd vss FILLER_0_6_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_3_72 vdd vss FILLER_0_3_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_8_28 vdd vss FILLER_0_8_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_17_ vss _17_/Z _17_/I vdd _17_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_10_101 vdd vss FILLER_0_10_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_16_ vss _16_/Z _16_/I vdd _16_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_9_72 vdd vss FILLER_0_9_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_15_64 vdd vss FILLER_0_15_64/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_9_104 vdd vss FILLER_0_9_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XFILLER_0_6_107 vdd vss FILLER_0_6_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_15_ vss _15_/Z _15_/I vdd _15_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_2 vdd vss FILLER_0_15_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_4_2 vdd vss FILLER_0_4_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_14_ vss _14_/Z _14_/I vdd _14_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XANTENNA_input9_I vss input_signal[8] vdd ANTENNA_input9_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_12_12 vdd vss FILLER_0_12_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_2_101 vdd vss FILLER_0_2_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
X_13_ vss _13_/Z _13_/I vdd _13_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_15_56 vdd vss FILLER_0_15_56/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_12_ vss _12_/Z _12_/I vdd _12_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_3_44 vdd vss FILLER_0_3_44/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_0_12 vdd vss FILLER_0_0_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_13_2 vdd vss FILLER_0_13_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_12 vdd vss FILLER_0_3_12/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_2_2 vdd vss FILLER_0_2_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
X_11_ vss _11_/Z _11_/I vdd _11_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1$1
XFILLER_0_9_66 vdd vss FILLER_0_9_66/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XANTENNA_input7_I vss input_signal[6] vdd ANTENNA_input7_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_12_37 vdd vss FILLER_0_12_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_107 vdd vss FILLER_0_10_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_13_104 vdd vss FILLER_0_13_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
X_10_ vss _10_/Z _10_/I vdd _10_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1$1
XFILLER_0_0_36 vdd vss FILLER_0_0_36/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_15_8 vdd vss FILLER_0_15_8/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XFILLER_0_11_2 vdd vss FILLER_0_11_2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_70 vdd vss FILLER_0_16_70/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_12_28 vdd vss FILLER_0_12_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_6_37 vdd vss FILLER_0_6_37/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input5_I vss input_signal[4] vdd ANTENNA_input5_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_8_101 vdd vss FILLER_0_8_101/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_16_104 vdd vss FILLER_0_16_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_2_107 vdd vss FILLER_0_2_107/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16$1
XFILLER_0_5_104 vdd vss FILLER_0_5_104/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
XANTENNA__11__I vss _11_/I vdd ANTENNA__11__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_13_72 vdd vss FILLER_0_13_72/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32$1
XANTENNA__06__I vss _15_/I vdd ANTENNA__06__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
XFILLER_0_0_28 vdd vss FILLER_0_0_28/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4$1
XFILLER_0_1_60 vdd vss FILLER_0_1_60/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8$1
Xoutput30 output_signal_plus[9] _19_/Z vdd vss output30/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8$1
XANTENNA__14__I vss _14_/I vdd ANTENNA__14__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna$1
.ends

.subckt dac_in inputp inputm vss vdd input_signal[0] input_signal[1] input_signal[2]
+ input_signal[3] input_signal[4] input_signal[5] input_signal[6] input_signal[7]
+ input_signal[8] input_signal[9]
Xphase_inverter_0 input_signal[0] input_signal[1] input_signal[2] input_signal[3]
+ input_signal[4] input_signal[5] input_signal[9] carray_in_1/n0 carray_in_1/n1 carray_in_1/n2
+ carray_in_1/n3 carray_in_1/n4 carray_in_1/n5 carray_in_1/n6 carray_in_1/n7 carray_in_1/n8
+ carray_in_1/n9 carray_in_0/n0 carray_in_0/n1 carray_in_0/n2 carray_in_0/n3 carray_in_0/n4
+ carray_in_0/n5 carray_in_0/n6 carray_in_0/n7 carray_in_0/n8 carray_in_0/n9 input_signal[7]
+ input_signal[8] input_signal[6] vdd vss phase_inverter
.ends

