* NGSPICE file created from sarlogic.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VPW VNW a_36_472# a_572_375# VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VNW VDD 0.11314f
C1 a_572_375# VDD 0.129266f
C2 VSS a_484_472# 0.148682f
C3 VSS a_124_375# 0.136476f
C4 VSS a_36_472# 0.151218f
C5 a_572_375# a_484_472# 0.285629f
C6 a_124_375# a_36_472# 0.285629f
C7 a_124_375# VNW 0.180172f
C8 a_484_472# VDD 0.179463f
C9 a_572_375# VNW 0.18122f
C10 a_124_375# VDD 0.12673f
C11 VSS VSUBS 0.360066f
C12 VDD VSUBS 0.286281f
C13 VNW VSUBS 1.65967f
C14 a_484_472# VSUBS 0.345058f
C15 a_36_472# VSUBS 0.404746f
C16 a_572_375# VSUBS 0.232991f
C17 a_124_375# VSUBS 0.185089f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VPW VNW VSUBS
D0 VSUBS I diode_nd2ps_06v0 pj=1.86u area=0.2052p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.2052p
C0 VSS VSUBS 0.12617f
C1 I VSUBS 0.139667f
C2 VNW VSUBS 0.615384f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 ZN A2 0.378409f
C1 ZN A1 0.579732f
C2 VDD A2 0.255318f
C3 VNW A2 0.128798f
C4 VSS A1 0.168633f
C5 VNW A1 0.136915f
C6 VDD ZN 0.117921f
C7 VSS VSUBS 0.331491f
C8 VDD VSUBS 0.218051f
C9 A1 VSUBS 0.331856f
C10 A2 VSUBS 0.334514f
C11 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD VPW VNW a_2665_112# a_36_151#
+ VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2 Q a_2665_112# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X5 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X15 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X16 a_2665_112# RN VDD VNW pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X24 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X25 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X26 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 D a_448_472# 0.328788f
C1 a_2665_112# RN 0.336469f
C2 a_448_472# a_2248_156# 0.510371f
C3 a_36_151# a_448_472# 0.536965f
C4 VSS a_448_472# 1.20207f
C5 VDD a_1204_472# 0.282626f
C6 VNW CLK 0.137037f
C7 a_2560_156# a_448_472# 0.277491f
C8 VNW D 0.128231f
C9 VNW a_2248_156# 0.212431f
C10 VNW a_36_151# 1.28833f
C11 a_1308_423# a_1000_472# 0.934191f
C12 VDD Q 0.149344f
C13 a_1000_472# a_1204_472# 0.66083f
C14 VDD a_2248_156# 1.11667f
C15 VDD a_36_151# 0.417088f
C16 a_796_472# a_448_472# 0.401636f
C17 RN VSS 0.441968f
C18 VNW a_448_472# 0.341284f
C19 a_2665_112# Q 0.109436f
C20 VDD a_448_472# 0.456269f
C21 a_2665_112# a_2248_156# 0.633318f
C22 a_2665_112# VSS 0.184997f
C23 a_2665_112# a_2560_156# 0.116059f
C24 a_1000_472# a_448_472# 0.361958f
C25 VNW VDD 0.503557f
C26 VNW RN 0.329494f
C27 CLK a_36_151# 0.669598f
C28 a_1308_423# a_448_472# 0.882105f
C29 VNW a_1000_472# 0.241357f
C30 VSS Q 0.113401f
C31 a_2665_112# VNW 0.354715f
C32 VSS a_36_151# 0.291264f
C33 VDD a_1000_472# 0.119211f
C34 a_2560_156# a_2248_156# 0.119687f
C35 a_2665_112# VDD 0.102046f
C36 a_1308_423# VNW 0.149014f
C37 a_2560_156# VSS 0.128503f
C38 Q VSUBS 0.114762f
C39 VSS VSUBS 1.26186f
C40 RN VSUBS 1.36673f
C41 D VSUBS 0.253406f
C42 VDD VSUBS 0.79945f
C43 CLK VSUBS 0.291241f
C44 VNW VSUBS 6.1377f
C45 a_2665_112# VSUBS 0.62251f
C46 a_2248_156# VSUBS 0.371662f
C47 a_1000_472# VSUBS 0.291735f
C48 a_1308_423# VSUBS 0.279043f
C49 a_448_472# VSUBS 0.684413f
C50 a_36_151# VSUBS 1.43589f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VPW VNW a_36_68# VSUBS
X0 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 ZN a_36_68# 0.419486f
C1 a_36_68# A2 0.340509f
C2 a_36_68# VSS 0.392965f
C3 A1 VNW 0.115376f
C4 a_36_68# B2 0.369561f
C5 a_36_68# VDD 0.787847f
C6 ZN A2 0.390894f
C7 VNW B1 0.125926f
C8 VNW A2 0.125671f
C9 A1 a_36_68# 0.160084f
C10 VDD B2 0.246452f
C11 A1 B1 0.163724f
C12 VNW B2 0.133721f
C13 VNW VDD 0.139306f
C14 a_36_68# B1 0.437534f
C15 ZN A1 0.430191f
C16 VSS VSUBS 0.383233f
C17 VDD VSUBS 0.318857f
C18 A2 VSUBS 0.2826f
C19 A1 VSUBS 0.258579f
C20 B1 VSUBS 0.257485f
C21 B2 VSUBS 0.309037f
C22 VNW VSUBS 2.00777f
C23 a_36_68# VSUBS 0.150048f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VPW VNW a_49_472#
+ VSUBS
X0 ZN B1 a_257_69# VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VSUBS nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
C0 VDD VNW 0.112326f
C1 A2 ZN 0.102518f
C2 VNW A2 0.131727f
C3 B1 B2 0.18297f
C4 VDD a_49_472# 0.887006f
C5 A2 VSS 0.150463f
C6 a_49_472# ZN 0.239204f
C7 VNW B2 0.129409f
C8 B1 ZN 0.367665f
C9 VNW B1 0.109456f
C10 A1 ZN 0.447732f
C11 A1 A2 0.392541f
C12 VNW A1 0.10965f
C13 B2 a_49_472# 0.151151f
C14 VSS VSUBS 0.39457f
C15 VDD VSUBS 0.243433f
C16 A2 VSUBS 0.322629f
C17 A1 VSUBS 0.250967f
C18 B1 VSUBS 0.261124f
C19 B2 VSUBS 0.322244f
C20 VNW VSUBS 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VPW VNW a_36_160# VSUBS
X0 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VSS Z 0.146199f
C1 a_36_160# Z 0.281838f
C2 Z VDD 0.128274f
C3 I VSS 0.12329f
C4 I a_36_160# 0.545454f
C5 a_36_160# VDD 0.2736f
C6 a_36_160# VNW 0.170864f
C7 I VNW 0.2276f
C8 VSS VSUBS 0.28275f
C9 Z VSUBS 0.10469f
C10 VDD VSUBS 0.178615f
C11 I VSUBS 0.323491f
C12 VNW VSUBS 1.31158f
C13 a_36_160# VSUBS 0.386641f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 I VNW 0.135368f
C1 ZN I 0.47009f
C2 I VDD 0.157124f
C3 VSS VSUBS 0.242183f
C4 VDD VSUBS 0.182097f
C5 I VSUBS 0.355642f
C6 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 I VNW 0.137757f
C1 ZN VSS 0.115297f
C2 ZN VDD 0.137375f
C3 ZN I 0.262199f
C4 VSS VSUBS 0.2316f
C5 ZN VSUBS 0.113404f
C6 VDD VSUBS 0.181139f
C7 I VSUBS 0.341982f
C8 VNW VSUBS 0.96348f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VPW VNW a_36_472# a_124_375# VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
C0 VNW a_124_375# 0.179924f
C1 a_36_472# a_124_375# 0.285629f
C2 VSS a_36_472# 0.150876f
C3 VDD a_124_375# 0.126034f
C4 VSS VSUBS 0.218985f
C5 VDD VSUBS 0.182777f
C6 VNW VSUBS 0.96348f
C7 a_36_472# VSUBS 0.417394f
C8 a_124_375# VSUBS 0.246306f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VPW VNW a_224_472# VSUBS
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 I a_224_472# 0.796069f
C1 VNW a_224_472# 1.14633f
C2 VSS Z 0.70427f
C3 VDD Z 0.819024f
C4 VSS I 0.158668f
C5 VDD I 0.1311f
C6 VDD VNW 0.305516f
C7 VSS a_224_472# 0.659695f
C8 VDD a_224_472# 0.74621f
C9 Z a_224_472# 2.29481f
C10 VNW I 0.55539f
C11 VSS VSUBS 0.910368f
C12 Z VSUBS 0.18914f
C13 VDD VSUBS 0.724491f
C14 I VSUBS 1.16773f
C15 VNW VSUBS 4.79254f
C16 a_224_472# VSUBS 2.38465f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VPW VNW a_36_472# VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VSUBS nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
C0 VNW A1 0.122087f
C1 a_36_472# A1 0.104556f
C2 A2 ZN 0.248411f
C3 A1 ZN 0.245346f
C4 B A1 0.157699f
C5 VNW B 0.137038f
C6 VNW VDD 0.11216f
C7 VNW A2 0.128282f
C8 a_36_472# VDD 0.581285f
C9 ZN VSS 0.304078f
C10 a_36_472# A2 0.10395f
C11 VSS VSUBS 0.361309f
C12 VDD VSUBS 0.259458f
C13 B VSUBS 0.378232f
C14 A1 VSUBS 0.264815f
C15 A2 VSUBS 0.3189f
C16 VNW VSUBS 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VPW VNW a_36_113# VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 VNW I 0.152645f
C1 a_36_113# VSS 0.11114f
C2 a_36_113# Z 0.191876f
C3 a_36_113# I 0.476912f
C4 VSS Z 0.136942f
C5 VNW a_36_113# 0.160792f
C6 a_36_113# VDD 0.278283f
C7 VSS VSUBS 0.283681f
C8 Z VSUBS 0.117185f
C9 VDD VSUBS 0.180237f
C10 I VSUBS 0.336876f
C11 VNW VSUBS 1.31158f
C12 a_36_113# VSUBS 0.418095f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VPW VNW a_3260_375# a_36_472#
+ VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_1916_375# a_1828_472# 0.285629f
C1 a_484_472# a_572_375# 0.285629f
C2 a_1380_472# a_1468_375# 0.285629f
C3 a_3260_375# VNW 0.18122f
C4 a_2812_375# VDD 0.129962f
C5 a_1020_375# VNW 0.181468f
C6 VSS a_2276_472# 0.142721f
C7 VDD a_1380_472# 0.179463f
C8 a_1020_375# VSS 0.131736f
C9 a_36_472# a_124_375# 0.285629f
C10 VDD a_932_472# 0.179463f
C11 a_1916_375# VNW 0.181468f
C12 a_2364_375# VNW 0.181468f
C13 a_2364_375# a_2276_472# 0.285629f
C14 a_484_472# VDD 0.179463f
C15 a_1916_375# VSS 0.131736f
C16 VDD a_3172_472# 0.179463f
C17 VSS a_2724_472# 0.142721f
C18 VNW a_572_375# 0.181468f
C19 a_2364_375# VSS 0.131736f
C20 VDD a_1828_472# 0.179463f
C21 VSS a_572_375# 0.131736f
C22 VNW a_124_375# 0.180172f
C23 VNW a_1468_375# 0.181468f
C24 VSS a_124_375# 0.131736f
C25 VSS a_1468_375# 0.131736f
C26 VNW VDD 0.425768f
C27 a_2812_375# VNW 0.181468f
C28 VDD a_2276_472# 0.179463f
C29 a_3260_375# VDD 0.129266f
C30 a_2812_375# VSS 0.131736f
C31 a_1020_375# VDD 0.129962f
C32 VSS a_1380_472# 0.142721f
C33 VSS a_932_472# 0.142721f
C34 a_1916_375# VDD 0.129962f
C35 a_1020_375# a_932_472# 0.285629f
C36 VDD a_2724_472# 0.179463f
C37 a_2812_375# a_2724_472# 0.285629f
C38 a_2364_375# VDD 0.129962f
C39 a_3260_375# a_3172_472# 0.285629f
C40 a_484_472# VSS 0.142721f
C41 VSS a_3172_472# 0.139489f
C42 VDD a_572_375# 0.129962f
C43 a_36_472# VSS 0.142026f
C44 VSS a_1828_472# 0.142721f
C45 VDD a_124_375# 0.12673f
C46 VDD a_1468_375# 0.129962f
C47 VSS VSUBS 1.20585f
C48 VDD VSUBS 0.907304f
C49 VNW VSUBS 5.83682f
C50 a_3172_472# VSUBS 0.345058f
C51 a_2724_472# VSUBS 0.33241f
C52 a_2276_472# VSUBS 0.33241f
C53 a_1828_472# VSUBS 0.33241f
C54 a_1380_472# VSUBS 0.33241f
C55 a_932_472# VSUBS 0.33241f
C56 a_484_472# VSUBS 0.33241f
C57 a_36_472# VSUBS 0.404746f
C58 a_3260_375# VSUBS 0.233093f
C59 a_2812_375# VSUBS 0.17167f
C60 a_2364_375# VSUBS 0.17167f
C61 a_1916_375# VSUBS 0.17167f
C62 a_1468_375# VSUBS 0.17167f
C63 a_1020_375# VSUBS 0.17167f
C64 a_572_375# VSUBS 0.17167f
C65 a_124_375# VSUBS 0.185915f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_455_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 VDD ZN 0.33173f
C1 A1 ZN 0.384588f
C2 VNW A2 0.121191f
C3 VSS A2 0.104901f
C4 VNW A3 0.148237f
C5 VNW VDD 0.112537f
C6 VNW A1 0.12917f
C7 A3 A2 0.117566f
C8 A2 A1 0.133044f
C9 VSS VSUBS 0.307914f
C10 ZN VSUBS 0.133449f
C11 VDD VSUBS 0.241872f
C12 A1 VSUBS 0.287469f
C13 A2 VSUBS 0.25736f
C14 A3 VSUBS 0.326833f
C15 VNW VSUBS 1.48562f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
C0 A1 VNW 0.119756f
C1 A1 VSS 0.131667f
C2 A1 A2 0.226398f
C3 VDD ZN 0.240333f
C4 A1 ZN 0.351362f
C5 VNW A2 0.125396f
C6 VSS VSUBS 0.238729f
C7 ZN VSUBS 0.105772f
C8 VDD VSUBS 0.243067f
C9 A1 VSUBS 0.290957f
C10 A2 VSUBS 0.314823f
C11 VNW VSUBS 1.13753f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
C0 Z a_67_603# 0.181586f
C1 VDD a_67_603# 0.307039f
C2 Z VSS 0.158265f
C3 VNW A1 0.220003f
C4 A2 VDD 0.147628f
C5 VNW a_67_603# 0.157241f
C6 Z VDD 0.196046f
C7 A1 a_67_603# 0.540888f
C8 A2 VNW 0.216313f
C9 VNW VDD 0.11771f
C10 VSS a_67_603# 0.250493f
C11 A2 a_67_603# 0.505374f
C12 VSS VSUBS 0.359722f
C13 Z VSUBS 0.102754f
C14 VDD VSUBS 0.233025f
C15 A2 VSUBS 0.313441f
C16 A1 VSUBS 0.39469f
C17 VNW VSUBS 1.65967f
C18 a_67_603# VSUBS 0.345683f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 VSS C a_2960_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X20 VSS C a_2124_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X23 a_36_68# B a_2552_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X26 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
C0 ZN A1 1.37575f
C1 a_36_68# C 0.105844f
C2 VDD A2 0.15752f
C3 B VNW 0.600992f
C4 A2 A1 1.73987f
C5 ZN C 0.514613f
C6 a_36_68# ZN 1.98502f
C7 a_36_68# VSS 3.64719f
C8 B C 1.73339f
C9 A2 VNW 0.590323f
C10 a_36_68# B 1.37417f
C11 VDD VNW 0.366897f
C12 a_36_68# A2 0.108262f
C13 A1 VNW 0.51833f
C14 B ZN 0.426118f
C15 ZN A2 1.2828f
C16 VDD ZN 2.06829f
C17 C VNW 0.636287f
C18 B VDD 0.100578f
C19 VSS VSUBS 1.08055f
C20 VDD VSUBS 0.846798f
C21 C VSUBS 1.06351f
C22 B VSUBS 1.11555f
C23 A1 VSUBS 1.1956f
C24 A2 VSUBS 1.16629f
C25 VNW VSUBS 5.892971f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VPW VNW a_36_160# VSUBS
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VSUBS nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VSUBS nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
C0 VDD VNW 0.111398f
C1 a_36_160# VNW 0.302514f
C2 Z VSS 0.111496f
C3 a_36_160# VSS 0.114407f
C4 VDD Z 0.161733f
C5 a_36_160# VDD 0.31851f
C6 I VNW 0.1633f
C7 a_36_160# Z 0.426617f
C8 I VSS 0.178818f
C9 a_36_160# I 0.564508f
C10 VSS VSUBS 0.397291f
C11 VDD VSUBS 0.238155f
C12 I VSUBS 0.333888f
C13 VNW VSUBS 1.65967f
C14 a_36_160# VSUBS 0.696445f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VPW VNW a_36_472# a_1468_375#
+ VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
C0 a_124_375# VSS 0.134699f
C1 a_572_375# VNW 0.181468f
C2 a_1468_375# VNW 0.18122f
C3 VSS a_484_472# 0.148077f
C4 VSS a_932_472# 0.148077f
C5 a_1020_375# a_932_472# 0.285629f
C6 a_1020_375# VNW 0.181468f
C7 a_572_375# VSS 0.134699f
C8 a_124_375# VDD 0.12673f
C9 VSS a_36_472# 0.147381f
C10 a_1380_472# a_1468_375# 0.285629f
C11 VDD a_484_472# 0.179463f
C12 VDD a_932_472# 0.179463f
C13 a_1020_375# VSS 0.134699f
C14 a_1380_472# VSS 0.144845f
C15 VDD VNW 0.217349f
C16 a_572_375# VDD 0.129962f
C17 VDD a_1468_375# 0.129266f
C18 a_124_375# VNW 0.180172f
C19 a_124_375# a_36_472# 0.285629f
C20 a_1020_375# VDD 0.129962f
C21 a_572_375# a_484_472# 0.285629f
C22 a_1380_472# VDD 0.179463f
C23 VSS VSUBS 0.642184f
C24 VDD VSUBS 0.493288f
C25 VNW VSUBS 3.05206f
C26 a_1380_472# VSUBS 0.345058f
C27 a_932_472# VSUBS 0.33241f
C28 a_484_472# VSUBS 0.33241f
C29 a_36_472# VSUBS 0.404746f
C30 a_1468_375# VSUBS 0.233029f
C31 a_1020_375# VSUBS 0.171606f
C32 a_572_375# VSUBS 0.171606f
C33 a_124_375# VSUBS 0.185399f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VPW VNW a_36_68# VSUBS
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VSUBS nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 VNW VDD 0.114912f
C1 VSS a_36_68# 0.156367f
C2 a_36_68# Z 0.432914f
C3 I a_36_68# 0.731677f
C4 VSS Z 0.133443f
C5 VSS I 0.128735f
C6 VDD a_36_68# 0.271105f
C7 VNW a_36_68# 0.296832f
C8 VDD Z 0.172592f
C9 VNW I 0.133333f
C10 VSS VSUBS 0.338876f
C11 Z VSUBS 0.103236f
C12 VDD VSUBS 0.234026f
C13 I VSUBS 0.298844f
C14 VNW VSUBS 1.65967f
C15 a_36_68# VSUBS 0.69549f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VPW VNW a_848_380# VSUBS
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VSUBS nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VSUBS nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
C0 I1 VNW 0.127749f
C1 a_848_380# S 0.754833f
C2 a_124_24# I1 0.564972f
C3 VDD VNW 0.182986f
C4 a_124_24# VDD 0.309232f
C5 VSS a_848_380# 0.130064f
C6 I0 VNW 0.103064f
C7 VSS Z 0.129676f
C8 a_124_24# VNW 0.277682f
C9 a_848_380# VDD 0.319708f
C10 I0 S 0.533789f
C11 VDD Z 0.20273f
C12 VNW S 0.253706f
C13 a_124_24# S 0.245829f
C14 a_848_380# VNW 0.174516f
C15 a_124_24# a_848_380# 0.302602f
C16 VSS I0 0.124513f
C17 I1 VDD 0.227359f
C18 VSS a_124_24# 0.501844f
C19 a_124_24# Z 0.219295f
C20 VSS VSUBS 0.565512f
C21 VDD VSUBS 0.424967f
C22 I0 VSUBS 0.267152f
C23 S VSUBS 0.549493f
C24 I1 VSUBS 0.247562f
C25 VNW VSUBS 2.87801f
C26 a_848_380# VSUBS 0.40208f
C27 a_124_24# VSUBS 0.591898f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VPW VNW VSUBS
X0 VSS B a_36_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
C0 VNW VDD 0.117098f
C1 ZN a_36_68# 0.56857f
C2 a_36_68# VDD 0.753239f
C3 VSS a_36_68# 0.117681f
C4 VNW B 0.163023f
C5 a_36_68# B 0.389329f
C6 VSS B 0.198567f
C7 A1 VNW 0.117811f
C8 VNW A2 0.122386f
C9 A1 a_36_68# 0.292244f
C10 a_36_68# A2 0.489122f
C11 ZN A1 0.496662f
C12 ZN A2 0.400775f
C13 VSS VSUBS 0.342662f
C14 VDD VSUBS 0.256635f
C15 B VSUBS 0.339176f
C16 A1 VSUBS 0.256004f
C17 A2 VSUBS 0.28395f
C18 VNW VSUBS 1.65967f
C19 a_36_68# VSUBS 0.112263f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VPW VNW VSUBS
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
C0 I a_224_552# 0.421587f
C1 Z VSS 0.275062f
C2 VNW VDD 0.176912f
C3 VDD Z 0.356369f
C4 I VNW 0.376531f
C5 a_224_552# VSS 0.331404f
C6 a_224_552# VNW 0.5926f
C7 a_224_552# VDD 0.347549f
C8 a_224_552# Z 1.17071f
C9 VSS VSUBS 0.628617f
C10 Z VSUBS 0.102362f
C11 VDD VSUBS 0.415149f
C12 I VSUBS 0.471574f
C13 VNW VSUBS 2.70396f
C14 a_224_552# VSUBS 1.31114f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
C0 VDD A2 0.13595f
C1 VSS ZN 0.460527f
C2 VNW VDD 0.137685f
C3 A1 A2 0.636124f
C4 ZN VDD 0.517479f
C5 A1 VNW 0.25895f
C6 VNW A2 0.275679f
C7 A1 ZN 0.274601f
C8 ZN A2 0.509001f
C9 VSS VSUBS 0.451405f
C10 ZN VSUBS 0.138491f
C11 VDD VSUBS 0.322159f
C12 A1 VSUBS 0.557317f
C13 A2 VSUBS 0.617688f
C14 VNW VSUBS 2.00777f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
C0 VNW VDD 0.11801f
C1 A2 A1 0.145555f
C2 ZN VDD 0.116419f
C3 VNW A1 0.127941f
C4 ZN A1 0.499849f
C5 A3 A2 0.416588f
C6 ZN VSS 0.283414f
C7 VNW A3 0.136756f
C8 VNW A2 0.116878f
C9 A3 VDD 0.201466f
C10 VSS VSUBS 0.367618f
C11 ZN VSUBS 0.134331f
C12 VDD VSUBS 0.264623f
C13 A1 VSUBS 0.311038f
C14 A2 VSUBS 0.285534f
C15 A3 VSUBS 0.334053f
C16 VNW VSUBS 1.65967f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A1 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.2561p ps=1.505u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.1722p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
C0 VDD VNW 0.292073f
C1 VDD A3 0.107959f
C2 A1 a_36_68# 0.118844f
C3 ZN a_36_68# 0.885472f
C4 A1 ZN 1.266f
C5 a_36_68# VSS 2.77545f
C6 VDD A1 0.115489f
C7 VDD ZN 1.57207f
C8 A2 VNW 0.630933f
C9 A2 A3 1.65768f
C10 A3 VNW 0.599629f
C11 A2 a_36_68# 0.223434f
C12 A1 VNW 0.700258f
C13 A3 a_36_68# 1.03106f
C14 A2 ZN 1.77619f
C15 A3 ZN 0.150755f
C16 A2 VDD 0.124271f
C17 VSS VSUBS 0.861061f
C18 ZN VSUBS 0.103891f
C19 VDD VSUBS 0.701563f
C20 A1 VSUBS 1.27704f
C21 A3 VSUBS 1.11693f
C22 A2 VSUBS 1.08692f
C23 VNW VSUBS 4.73584f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VSUBS nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VSUBS nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
C0 VNW a_36_159# 0.162496f
C1 A2 VDD 0.184025f
C2 VSS Z 0.102819f
C3 a_36_159# VSS 0.244357f
C4 VNW VDD 0.125609f
C5 VNW A1 0.206765f
C6 VNW A2 0.20463f
C7 a_36_159# Z 0.215269f
C8 Z VDD 0.158212f
C9 a_36_159# VDD 0.130189f
C10 a_36_159# A1 0.377122f
C11 a_36_159# A2 0.472781f
C12 VSS VSUBS 0.35312f
C13 VDD VSUBS 0.251252f
C14 A2 VSUBS 0.262264f
C15 A1 VSUBS 0.321274f
C16 VNW VSUBS 1.65967f
C17 a_36_159# VSUBS 0.374116f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VPW VNW VSUBS
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VSUBS nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VSUBS nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VSUBS nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VSUBS nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VSUBS nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VSUBS nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VSUBS nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VSUBS nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
C0 B C 1.34577f
C1 ZN A1 1.40746f
C2 ZN B 0.231932f
C3 VSS B 0.119454f
C4 VNW A1 0.480244f
C5 a_170_472# B 2.12702f
C6 VNW B 0.617219f
C7 A2 ZN 1.83822f
C8 A2 VSS 0.104058f
C9 A2 a_170_472# 0.109943f
C10 A2 VNW 0.513788f
C11 A2 A1 1.72617f
C12 VDD a_170_472# 2.96356f
C13 VNW VDD 0.393677f
C14 VDD B 0.110239f
C15 ZN C 1.79111f
C16 VNW C 0.61926f
C17 ZN VSS 1.77446f
C18 ZN a_170_472# 0.818521f
C19 VSS VSUBS 1.33264f
C20 VDD VSUBS 0.809429f
C21 ZN VSUBS 0.171181f
C22 C VSUBS 1.26656f
C23 B VSUBS 1.19887f
C24 A1 VSUBS 1.12703f
C25 A2 VSUBS 1.09165f
C26 VNW VSUBS 6.53302f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
C0 VNW VDD 0.286001f
C1 a_36_472# A1 0.174868f
C2 VNW A1 0.520086f
C3 A3 a_36_472# 0.100976f
C4 a_36_472# A2 0.993181f
C5 ZN VSS 2.18568f
C6 A3 A2 1.6562f
C7 A3 VNW 0.478769f
C8 VNW A2 0.539636f
C9 ZN A1 1.56829f
C10 VSS A1 0.115774f
C11 ZN a_36_472# 0.362263f
C12 VDD a_36_472# 1.90933f
C13 ZN A3 1.42151f
C14 ZN A2 0.250963f
C15 A3 VSS 0.10353f
C16 VSS A2 0.128956f
C17 VSS VSUBS 0.918064f
C18 ZN VSUBS 0.159858f
C19 VDD VSUBS 0.61695f
C20 A1 VSUBS 1.35739f
C21 A3 VSUBS 1.33073f
C22 A2 VSUBS 1.29013f
C23 VNW VSUBS 4.79254f
C24 a_36_472# VSUBS 0.137725f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VSUBS nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VSUBS nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
C0 A2 VNW 0.241313f
C1 A3 A1 0.292395f
C2 A3 ZN 1.03634f
C3 ZN VSS 1.3936f
C4 A2 A1 0.570018f
C5 A2 A3 0.624599f
C6 VNW VDD 0.178574f
C7 A2 ZN 0.694728f
C8 A3 VDD 0.178286f
C9 VDD ZN 0.579119f
C10 VNW A1 0.254404f
C11 VNW A3 0.28584f
C12 VSS VSUBS 0.509614f
C13 ZN VSUBS 0.172636f
C14 VDD VSUBS 0.441158f
C15 A1 VSUBS 0.622214f
C16 A2 VSUBS 0.627317f
C17 A3 VSUBS 0.692739f
C18 VNW VSUBS 2.70396f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VSS B ZN VSUBS nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X1 VSS C ZN VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VSUBS nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VSUBS nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VSUBS nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
C0 A2 ZN 0.752866f
C1 VNW C 0.268332f
C2 B C 0.560408f
C3 VDD a_36_488# 1.67897f
C4 a_36_488# ZN 0.459425f
C5 B VNW 0.298561f
C6 VNW A1 0.25321f
C7 A2 VNW 0.280457f
C8 VSS ZN 0.708286f
C9 A2 A1 0.652956f
C10 ZN C 0.191881f
C11 VDD VNW 0.191798f
C12 B a_36_488# 0.80489f
C13 B ZN 0.413891f
C14 ZN A1 0.372797f
C15 VSS VSUBS 0.653933f
C16 VDD VSUBS 0.406726f
C17 C VSUBS 0.626227f
C18 B VSUBS 0.654892f
C19 A1 VSUBS 0.552174f
C20 A2 VSUBS 0.559992f
C21 VNW VSUBS 3.2261f
C22 a_36_488# VSUBS 0.101145f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.161025p ps=1.135u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161025p pd=1.135u as=0.194p ps=1.415u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.415u as=93.59999f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.35315p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.35315p ps=1.96u w=1.22u l=0.5u
C0 A3 Z 0.259021f
C1 VNW a_728_93# 0.346549f
C2 A2 VNW 0.369075f
C3 A3 a_728_93# 0.720358f
C4 A1 a_728_93# 0.12992f
C5 A2 A1 0.321942f
C6 VSS Z 0.277351f
C7 a_1336_472# a_728_93# 0.62718f
C8 a_1936_472# Z 0.337902f
C9 VSS a_728_93# 0.709567f
C10 a_1936_472# VDD 0.595117f
C11 a_1936_472# a_728_93# 0.105997f
C12 VNW A3 0.268193f
C13 VNW A1 0.293766f
C14 a_1336_472# VNW 0.144065f
C15 a_1336_472# A3 0.490376f
C16 VSS A1 0.139902f
C17 a_1336_472# VSS 0.326133f
C18 a_718_524# VDD 0.554575f
C19 a_718_524# a_728_93# 0.329834f
C20 A2 a_56_524# 0.908796f
C21 a_718_524# A2 0.107911f
C22 Z a_728_93# 0.402606f
C23 a_728_93# VDD 0.575073f
C24 A2 VDD 0.208821f
C25 VNW a_56_524# 0.188846f
C26 A2 a_728_93# 0.416172f
C27 a_56_524# A1 0.569057f
C28 VSS a_56_524# 0.214447f
C29 VNW VDD 0.360391f
C30 VSS VSUBS 0.861752f
C31 A1 VSUBS 0.602985f
C32 A2 VSUBS 0.640744f
C33 VDD VSUBS 0.543474f
C34 A3 VSUBS 0.593976f
C35 VNW VSUBS 4.270391f
C36 a_56_524# VSUBS 0.41096f
C37 a_728_93# VSUBS 0.654825f
C38 a_1336_472# VSUBS 0.316639f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
C0 VNW A2 0.277885f
C1 A1 VSS 0.115936f
C2 VNW A1 0.232646f
C3 ZN VDD 0.409997f
C4 A1 A2 0.708017f
C5 ZN VSS 0.2597f
C6 VNW VDD 0.123338f
C7 ZN A2 0.891023f
C8 A1 ZN 0.363066f
C9 VSS VSUBS 0.385688f
C10 ZN VSUBS 0.120217f
C11 VDD VSUBS 0.305683f
C12 A1 VSUBS 0.522064f
C13 A2 VSUBS 0.568932f
C14 VNW VSUBS 1.83372f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VPW VNW VSUBS
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
C0 VDD ZN 1.08837f
C1 A1 A3 0.206693f
C2 a_36_68# ZN 1.49222f
C3 A2 A1 0.703324f
C4 VDD A3 0.555327f
C5 VNW A1 0.279057f
C6 B VNW 0.309147f
C7 VDD VNW 0.248379f
C8 a_36_68# A1 0.158235f
C9 B VDD 0.119783f
C10 B a_36_68# 0.184521f
C11 ZN A3 1.02771f
C12 A2 ZN 0.152712f
C13 A2 A3 1.11591f
C14 VNW A3 0.297068f
C15 a_36_68# VSS 2.0408f
C16 A1 ZN 0.619225f
C17 A2 VNW 0.281901f
C18 B ZN 0.244028f
C19 VSS VSUBS 0.663038f
C20 VDD VSUBS 0.512998f
C21 A1 VSUBS 0.643779f
C22 A2 VSUBS 0.561227f
C23 A3 VSUBS 0.573818f
C24 B VSUBS 0.585725f
C25 VNW VSUBS 3.48825f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK VPW VNW a_36_151# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2665_112# VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 VSS RN a_1456_156# VSUBS nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VDD a_2665_112# Q VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_796_472# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5 VSS a_2665_112# a_2560_156# VSUBS nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 a_1000_472# a_448_472# a_796_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X7 a_2248_156# a_36_151# a_1308_423# VNW pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X8 a_2248_156# a_448_472# a_1308_423# VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 a_1456_156# a_1308_423# a_1288_156# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X11 a_1308_423# a_1000_472# VSS VSUBS nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X12 Q a_2665_112# VSS VSUBS nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X13 a_2665_112# a_2248_156# a_3041_156# VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X14 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X15 a_1204_472# a_36_151# a_1000_472# VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X16 a_1204_472# RN VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X17 a_2560_156# a_36_151# a_2248_156# VSUBS nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X18 a_1288_156# a_448_472# a_1000_472# VSUBS nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_2665_112# RN VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X20 VDD a_1308_423# a_1204_472# VNW pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X21 a_2560_156# a_448_472# a_2248_156# VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 VDD a_2248_156# a_2665_112# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X24 a_3041_156# RN VSS VSUBS nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X25 VSS a_2665_112# Q VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X26 VDD a_2665_112# a_2560_156# VNW pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X27 a_1308_423# a_1000_472# VDD VNW pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X28 a_1000_472# a_36_151# a_796_472# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X29 a_796_472# D VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
C0 VDD a_2665_112# 0.152571f
C1 a_36_151# VDD 0.417101f
C2 a_448_472# VSS 1.20207f
C3 a_36_151# a_448_472# 0.536965f
C4 a_2248_156# a_2665_112# 0.63615f
C5 VNW a_2665_112# 0.486803f
C6 VNW a_36_151# 1.28833f
C7 RN a_2665_112# 0.322698f
C8 VSS RN 0.436942f
C9 VDD a_448_472# 0.456269f
C10 D a_448_472# 0.328788f
C11 a_2248_156# VDD 1.12036f
C12 VNW CLK 0.137037f
C13 VDD a_1204_472# 0.282626f
C14 a_2248_156# a_448_472# 0.510371f
C15 VNW VDD 0.546785f
C16 a_1308_423# a_448_472# 0.882105f
C17 VNW D 0.128231f
C18 VNW a_448_472# 0.341284f
C19 a_2248_156# VNW 0.181292f
C20 VNW a_1308_423# 0.149014f
C21 VNW RN 0.304626f
C22 a_2560_156# a_2665_112# 0.116229f
C23 a_2560_156# VSS 0.128503f
C24 a_1000_472# VDD 0.119211f
C25 Q a_2665_112# 0.263315f
C26 VSS Q 0.170514f
C27 a_1000_472# a_448_472# 0.361958f
C28 VSS a_2665_112# 0.21484f
C29 a_36_151# VSS 0.291264f
C30 a_1000_472# a_1204_472# 0.66083f
C31 a_2560_156# a_448_472# 0.277491f
C32 a_1308_423# a_1000_472# 0.934191f
C33 VNW a_1000_472# 0.241357f
C34 a_448_472# a_796_472# 0.401636f
C35 a_2248_156# a_2560_156# 0.119687f
C36 VDD Q 0.260055f
C37 a_36_151# CLK 0.669598f
C38 VSS VSUBS 1.33519f
C39 RN VSUBS 1.37098f
C40 D VSUBS 0.253406f
C41 VDD VSUBS 0.859994f
C42 CLK VSUBS 0.291241f
C43 VNW VSUBS 6.48579f
C44 a_2665_112# VSUBS 0.91969f
C45 a_2248_156# VSUBS 0.30886f
C46 a_1000_472# VSUBS 0.291735f
C47 a_1308_423# VSUBS 0.279043f
C48 a_448_472# VSUBS 0.684413f
C49 a_36_151# VSUBS 1.43587f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_1458_68# A3 a_1254_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VSUBS nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
C0 VNW A1 0.345207f
C1 VNW VDD 0.1769f
C2 A3 A2 0.40854f
C3 A2 A4 0.762551f
C4 VNW A2 0.317841f
C5 A3 VSS 0.248503f
C6 ZN VDD 1.39778f
C7 A3 A4 0.297972f
C8 A3 VNW 0.300046f
C9 VNW A4 0.388525f
C10 A1 A2 0.516286f
C11 ZN VSS 0.89636f
C12 ZN A3 0.881941f
C13 ZN A4 1.94271f
C14 A3 A1 0.831807f
C15 A1 A4 0.451294f
C16 VSS VSUBS 0.597574f
C17 VDD VSUBS 0.397078f
C18 ZN VSUBS 0.12583f
C19 A1 VSUBS 0.558392f
C20 A2 VSUBS 0.513744f
C21 A3 VSUBS 0.547819f
C22 A4 VSUBS 0.580825f
C23 VNW VSUBS 3.05206f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VPW VNW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VSUBS nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
C0 ZN I 0.614595f
C1 VDD ZN 0.24022f
C2 VSS ZN 0.15979f
C3 VNW I 0.283715f
C4 VDD VNW 0.103267f
C5 VDD I 0.164681f
C6 VSS VSUBS 0.345063f
C7 VDD VSUBS 0.235951f
C8 I VSUBS 0.642286f
C9 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
C0 VNW A3 0.13805f
C1 a_244_68# ZN 0.2576f
C2 VNW A1 0.125824f
C3 B1 A1 0.13457f
C4 ZN B2 0.371232f
C5 B1 ZN 0.457921f
C6 VDD a_244_68# 0.520053f
C7 a_244_68# B2 0.29062f
C8 B1 a_244_68# 0.212448f
C9 VDD VNW 0.158216f
C10 VNW B2 0.125762f
C11 A2 A3 0.129823f
C12 B1 VNW 0.116377f
C13 A1 ZN 0.164807f
C14 VSS a_244_68# 0.329999f
C15 A2 a_244_68# 0.356992f
C16 A2 VNW 0.121626f
C17 VDD A3 0.236688f
C18 a_244_68# A1 0.480797f
C19 VSS VSUBS 0.474343f
C20 VDD VSUBS 0.363224f
C21 B2 VSUBS 0.282623f
C22 B1 VSUBS 0.257203f
C23 A1 VSUBS 0.255736f
C24 A2 VSUBS 0.254473f
C25 A3 VSUBS 0.308666f
C26 VNW VSUBS 2.35586f
C27 a_244_68# VSUBS 0.138666f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_952_93# A1 a_728_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 a_244_567# A2 a_56_567# VNW pfet_06v0 ad=0.1026p pd=0.93u as=0.1584p ps=1.6u w=0.36u l=0.5u
X2 a_728_93# A1 a_718_527# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.1596p ps=1.13u w=0.56u l=0.5u
X3 ZN A3 a_1948_68# VSUBS nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN a_1296_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.352075p ps=1.895u w=1.095u l=0.5u
X5 VDD a_728_93# a_2172_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
X6 a_718_527# a_56_567# VDD VNW pfet_06v0 ad=0.1596p pd=1.13u as=0.184p ps=1.36u w=0.56u l=0.5u
X7 a_718_527# A2 a_728_93# VNW pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X8 VSS A1 a_56_567# VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X9 VSS A3 a_1504_93# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X10 a_1948_68# a_728_93# ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_2172_497# A3 ZN VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X12 a_1504_93# a_728_93# a_1296_93# VSUBS nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X13 a_56_567# A2 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X14 a_1948_68# a_1296_93# VSS VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X15 a_1296_93# a_728_93# VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X16 a_728_93# a_56_567# VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 VDD A3 a_1296_93# VNW pfet_06v0 ad=0.352075p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X18 VDD A1 a_244_567# VNW pfet_06v0 ad=0.184p pd=1.36u as=0.1026p ps=0.93u w=0.36u l=0.5u
X19 VSS A2 a_952_93# VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=57.599995f ps=0.68u w=0.36u l=0.6u
C0 A1 a_728_93# 0.281966f
C1 A2 A1 0.757944f
C2 VDD VNW 0.370487f
C3 VDD ZN 0.47211f
C4 a_56_567# VNW 0.187311f
C5 a_728_93# VNW 0.385878f
C6 A2 VNW 0.388997f
C7 ZN a_728_93# 0.663929f
C8 A3 a_728_93# 0.721889f
C9 a_1296_93# VNW 0.155715f
C10 a_1296_93# A3 0.356198f
C11 a_56_567# VSS 0.400197f
C12 VSS a_728_93# 0.328386f
C13 VDD a_728_93# 0.78216f
C14 A2 VDD 0.210416f
C15 a_1296_93# VSS 0.379749f
C16 a_56_567# A2 0.174541f
C17 A2 a_728_93# 0.516752f
C18 a_1296_93# a_728_93# 0.624643f
C19 a_1948_68# ZN 0.381585f
C20 A1 VNW 0.342048f
C21 a_1948_68# VSS 0.719859f
C22 A3 VNW 0.298581f
C23 a_718_527# VDD 0.618394f
C24 a_718_527# a_728_93# 0.21558f
C25 A2 a_718_527# 0.141128f
C26 a_56_567# A1 0.368741f
C27 VSS VSUBS 0.875791f
C28 A1 VSUBS 0.604039f
C29 A2 VSUBS 0.633287f
C30 VDD VSUBS 0.584594f
C31 A3 VSUBS 0.573218f
C32 VNW VSUBS 4.42794f
C33 a_56_567# VSUBS 0.424713f
C34 a_728_93# VSUBS 0.65929f
C35 a_1296_93# VSUBS 0.317801f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VPW VNW VSUBS
X0 a_1229_68# B a_36_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.21525p ps=1.345u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VSUBS nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4 a_36_68# B a_1657_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.31215p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.37905p pd=1.82u as=0.4599p ps=1.935u w=1.095u l=0.5u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.31215p ps=1.685u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X9 a_36_68# A2 ZN VSUBS nfet_06v0 ad=0.21525p pd=1.345u as=0.30965p ps=1.685u w=0.82u l=0.6u
X10 a_1657_68# C VSS VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.37905p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X13 VSS C a_1229_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
C0 VDD VNW 0.219901f
C1 C VNW 0.309331f
C2 A1 A2 0.722847f
C3 VNW A2 0.30827f
C4 VNW B 0.311256f
C5 VDD ZN 0.761655f
C6 ZN C 0.501479f
C7 ZN a_36_68# 0.528658f
C8 A1 VNW 0.269127f
C9 VDD A2 0.147417f
C10 ZN A2 1.02528f
C11 C B 0.698524f
C12 ZN B 0.3603f
C13 a_36_68# B 0.587375f
C14 VSS a_36_68# 2.1107f
C15 A1 ZN 0.622246f
C16 VSS VSUBS 0.620026f
C17 VDD VSUBS 0.531064f
C18 C VSUBS 0.529789f
C19 B VSUBS 0.589191f
C20 A1 VSUBS 0.58772f
C21 A2 VSUBS 0.613706f
C22 VNW VSUBS 3.34705f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VPW VNW VSUBS
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VSUBS nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VSUBS nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VSUBS nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VSUBS nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
C0 Z a_36_148# 0.156534f
C1 VDD Z 0.164783f
C2 VSS a_36_148# 0.798993f
C3 VNW A2 0.189332f
C4 A2 A3 0.340591f
C5 A2 a_36_148# 0.141951f
C6 VNW A3 0.213241f
C7 VNW a_36_148# 0.194548f
C8 VNW VDD 0.134134f
C9 A1 A2 0.307806f
C10 VNW A1 0.214361f
C11 a_36_148# A3 0.477475f
C12 VDD a_36_148# 0.556761f
C13 A1 a_36_148# 0.205722f
C14 VSS VSUBS 0.415001f
C15 VDD VSUBS 0.277732f
C16 A3 VSUBS 0.275015f
C17 A2 VSUBS 0.257076f
C18 A1 VSUBS 0.330738f
C19 VNW VSUBS 2.00777f
C20 a_36_148# VSUBS 0.388358f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VSUBS nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VSUBS nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VSUBS nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VSUBS nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
C0 VNW A2 0.279783f
C1 ZN A3 1.24554f
C2 VNW VDD 0.172362f
C3 A1 A2 0.708241f
C4 A3 A2 1.13496f
C5 A1 VNW 0.280755f
C6 VSS ZN 0.476547f
C7 VNW A3 0.347673f
C8 VSS A2 0.130985f
C9 ZN VDD 0.550625f
C10 A1 ZN 0.430404f
C11 VSS VSUBS 0.511432f
C12 ZN VSUBS 0.112753f
C13 VDD VSUBS 0.407724f
C14 A1 VSUBS 0.540441f
C15 A2 VSUBS 0.524145f
C16 A3 VSUBS 0.582222f
C17 VNW VSUBS 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X1 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.455625p pd=1.965u as=0.486p ps=2.015u w=1.215u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.486p ps=2.015u w=1.215u l=0.5u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.455625p ps=1.965u w=1.215u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.346275p ps=1.785u w=1.215u l=0.5u
X12 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X16 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346275p pd=1.785u as=0.5346p ps=3.31u w=1.215u l=0.5u
X18 VSS A4 ZN VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X20 VSS A2 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X26 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.015u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VSUBS nfet_06v0 ad=0.1584p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.015u as=0.486p ps=2.015u w=1.215u l=0.5u
X31 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
C0 A4 a_66_473# 0.100571f
C1 A4 A3 1.96796f
C2 ZN a_66_473# 0.956309f
C3 ZN A3 0.417545f
C4 VNW A2 0.584134f
C5 VDD VNW 0.394018f
C6 A2 a_66_473# 0.182327f
C7 VDD a_66_473# 3.19476f
C8 ZN A1 1.60655f
C9 ZN A4 1.44735f
C10 A1 A2 2.13585f
C11 VDD A4 0.110338f
C12 ZN A2 2.14591f
C13 ZN VSS 4.39577f
C14 VNW A3 0.567739f
C15 A3 a_66_473# 1.66251f
C16 A1 VNW 0.553741f
C17 A4 VNW 0.513548f
C18 VSS VSUBS 1.3434f
C19 ZN VSUBS 0.240026f
C20 VDD VSUBS 0.844436f
C21 A1 VSUBS 1.40024f
C22 A2 VSUBS 1.30271f
C23 A4 VSUBS 1.33565f
C24 A3 VSUBS 1.29175f
C25 VNW VSUBS 6.70706f
C26 a_66_473# VSUBS 0.11665f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VPW VNW VSUBS
X0 VSS A2 a_1133_69# VSUBS nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VSUBS nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VSUBS nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VSUBS nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VSUBS nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
C0 B ZN 0.20884f
C1 VNW A1 0.241301f
C2 A2 ZN 0.800412f
C3 VNW VDD 0.151549f
C4 VDD a_49_472# 1.09818f
C5 A2 A1 0.809974f
C6 ZN VSS 0.784804f
C7 ZN A1 0.182845f
C8 VNW B 0.260678f
C9 B a_49_472# 0.234399f
C10 VNW A2 0.272677f
C11 A1 VSS 0.129775f
C12 ZN a_49_472# 0.475008f
C13 VSS VSUBS 0.510011f
C14 VDD VSUBS 0.327438f
C15 A1 VSUBS 0.556927f
C16 A2 VSUBS 0.56333f
C17 B VSUBS 0.662515f
C18 VNW VSUBS 2.52991f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VPW VNW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
C0 ZN I 0.58604f
C1 VDD ZN 0.266247f
C2 VSS ZN 0.179304f
C3 VNW I 0.285482f
C4 VSS VSUBS 0.308828f
C5 ZN VSUBS 0.100523f
C6 VDD VSUBS 0.240805f
C7 I VSUBS 0.610668f
C8 VNW VSUBS 1.31158f
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN VPW VNW a_36_151# VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 a_1353_112# SETN a_1697_156# VSUBS nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2 a_836_156# D VDD VNW pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3 a_1040_527# a_36_151# a_836_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_1040_527# a_448_472# a_836_156# VNW pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X5 a_2225_156# a_36_151# a_1353_112# VNW pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X6 VSS a_1353_112# a_1284_156# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X7 a_2225_156# a_448_472# a_1353_112# VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 a_2449_156# a_448_472# a_2225_156# VNW pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X10 VDD a_3129_107# a_2449_156# VNW pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X11 Q a_3129_107# VSS VSUBS nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X12 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X13 a_2449_156# SETN VDD VNW pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X14 VSS a_3129_107# a_3081_151# VSUBS nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X15 a_836_156# D VSS VSUBS nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_1353_112# a_1040_527# VDD VNW pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X18 a_3129_107# a_2225_156# VSS VSUBS nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X19 VDD SETN a_1353_112# VNW pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X20 a_1284_156# a_448_472# a_1040_527# VSUBS nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X21 VDD a_1353_112# a_1293_527# VNW pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X22 Q a_3129_107# VDD VNW pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X23 a_3129_107# a_2225_156# VDD VNW pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X24 a_2449_156# a_36_151# a_2225_156# VSUBS nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X25 a_1293_527# a_36_151# a_1040_527# VNW pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X26 a_1697_156# a_1040_527# VSS VSUBS nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X27 a_3081_151# SETN a_2449_156# VSUBS nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
C0 VDD a_448_472# 0.624585f
C1 D a_448_472# 0.400104f
C2 a_1040_527# a_448_472# 0.869605f
C3 VNW SETN 0.811046f
C4 a_2225_156# a_448_472# 0.153996f
C5 VSS a_36_151# 0.286331f
C6 a_1353_112# a_1040_527# 0.387423f
C7 a_2225_156# a_1353_112# 0.152869f
C8 a_836_156# a_448_472# 0.427756f
C9 VSS a_3129_107# 0.136769f
C10 Q a_3129_107# 0.179468f
C11 CLK a_36_151# 0.700974f
C12 VSS a_448_472# 1.07431f
C13 a_36_151# VNW 0.909435f
C14 a_836_156# D 0.108102f
C15 CLK VNW 0.136589f
C16 a_3129_107# VNW 0.323464f
C17 VDD SETN 0.127822f
C18 a_36_151# a_448_472# 0.473132f
C19 a_1353_112# a_36_151# 0.840879f
C20 VNW a_448_472# 0.400964f
C21 a_2225_156# VSS 1.18908f
C22 Q VDD 0.282179f
C23 a_1353_112# VNW 0.219511f
C24 a_2449_156# VDD 0.208631f
C25 a_2225_156# a_2449_156# 0.569174f
C26 VDD a_36_151# 1.41468f
C27 a_36_151# a_1040_527# 0.206392f
C28 a_2225_156# a_36_151# 0.153684f
C29 a_1353_112# a_448_472# 0.317251f
C30 VDD VNW 0.539099f
C31 VDD a_3129_107# 0.351307f
C32 VNW D 0.1615f
C33 VNW a_1040_527# 0.223863f
C34 a_2225_156# VNW 0.209033f
C35 a_2449_156# SETN 0.302222f
C36 a_2225_156# a_3129_107# 0.514036f
C37 Q VSS 0.131272f
C38 Q VSUBS 0.105566f
C39 VSS VSUBS 1.35707f
C40 SETN VSUBS 0.710246f
C41 D VSUBS 0.247102f
C42 VDD VSUBS 0.833181f
C43 CLK VSUBS 0.290467f
C44 VNW VSUBS 6.44257f
C45 a_2225_156# VSUBS 0.434082f
C46 a_3129_107# VSUBS 0.58406f
C47 a_1040_527# VSUBS 0.302082f
C48 a_1353_112# VSUBS 0.286513f
C49 a_448_472# VSUBS 1.21246f
C50 a_36_151# VSUBS 1.31409f
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctln[8] ctln[9] 
+ ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] ctlp[8] ctlp[9] 
+ result[0] result[1] result[2] result[3] result[4] result[5] result[6] result[7] result[8] result[9] 
+ trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4] rstn en cal clk comp clkc sample valid vdd vss 

XFILLER_0_17_200 vdd vss FILLER_0_17_200/VPW vdd FILLER_0_17_200/a_36_472# FILLER_0_17_200/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout56_I vss net57 vdd ANTENNA_fanout56_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_294_ vdd vss _008_ _104_ _106_ _294_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_432_ _021_ mask\[3\] net63 vss net80 vdd _432_/VPW vdd _432_/a_2665_112# _432_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_363_ _153_ _154_ _155_ vdd vss _028_ _151_ _363_/VPW vdd _363_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_346_ _144_ mask\[5\] vdd vss _145_ mask\[4\] _141_ _346_/VPW vdd _346_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_415_ _004_ net27 net58 vss net75 vdd _415_/VPW vdd _415_/a_2665_112# _415_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_277_ vss _094_ _093_ vdd _277_/VPW vdd _277_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_200_ vdd vss net20 net10 _200_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_329_ vss _133_ calibrate vdd _329_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_19_125 vdd vss FILLER_0_19_125/VPW vdd FILLER_0_19_125/a_36_472# FILLER_0_19_125/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 vss _077_ vdd ANTENNA__392__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_150 vdd vss FILLER_0_15_150/VPW vdd FILLER_0_15_150/a_36_472# FILLER_0_15_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vss FILLER_0_21_142/VPW vdd FILLER_0_21_142/a_36_472# FILLER_0_21_142/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_73 vdd vss FILLER_0_16_73/VPW vdd FILLER_0_16_73/a_36_472# FILLER_0_16_73/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 ctlp[3] net20 vdd vss output20/VPW vdd output20/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 result[4] net31 vdd vss output31/VPW vdd output31/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 trim[4] net42 vdd vss output42/VPW vdd output42/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 ctln[0] net7 vdd vss output7/VPW vdd output7/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_117 vdd vss FILLER_0_5_117/VPW vdd FILLER_0_5_117/a_36_472# FILLER_0_5_117/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_128 vdd vss FILLER_0_5_128/VPW vdd FILLER_0_5_128/a_36_472# FILLER_0_5_128/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_293_ net31 vdd vss _106_ mask\[4\] _105_ _293_/VPW vdd _293_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_431_ _020_ mask\[2\] net53 vss net70 vdd _431_/VPW vdd _431_/a_2665_112# _431_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_362_ vdd vss trim_mask\[1\] _155_ _362_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_345_ vss _144_ _132_ vdd _345_/VPW vdd _345_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_276_ vss _093_ _092_ vdd _276_/VPW vdd _276_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_414_ _003_ cal_itt\[3\] net59 vss net76 vdd _414_/VPW vdd _414_/a_2665_112# _414_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_328_ vss _132_ _114_ vdd _328_/VPW vdd _328_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_28 vdd vss FILLER_0_9_28/VPW vdd FILLER_0_9_28/a_3260_375# FILLER_0_9_28/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_204 vdd vss FILLER_0_3_204/VPW vdd FILLER_0_3_204/a_36_472# FILLER_0_3_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _078_ vdd vss _080_ _073_ _076_ _259_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_107 vdd vss FILLER_0_16_107/VPW vdd FILLER_0_16_107/a_36_472# FILLER_0_16_107/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout79_I vss net81 vdd ANTENNA_fanout79_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__I vss _053_ vdd ANTENNA__358__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 ctlp[4] net21 vdd vss output21/VPW vdd output21/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 trimb[0] net43 vdd vss output43/VPW vdd output43/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 result[5] net32 vdd vss output32/VPW vdd output32/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 ctln[3] net10 vdd vss output10/VPW vdd output10/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 ctln[1] net8 vdd vss output8/VPW vdd output8/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input3_I vss comp vdd ANTENNA_input3_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ vss _105_ _098_ vdd _292_/VPW vdd _292_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_430_ _019_ mask\[1\] net63 vss net80 vdd _430_/VPW vdd _430_/a_2665_112# _430_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_361_ vdd vss _154_ _086_ _119_ _361_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_72 vdd vss FILLER_0_7_72/VPW vdd FILLER_0_7_72/a_3260_375# FILLER_0_7_72/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_344_ vdd vss _143_ _021_ _344_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ vdd vss _092_ _069_ _091_ _275_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__191__I vss net17 vdd ANTENNA__191__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ _002_ cal_itt\[2\] net59 vss net76 vdd _413_/VPW vdd _413_/a_2665_112# _413_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_24_96 vdd vss FILLER_0_24_96/VPW vdd FILLER_0_24_96/a_36_472# FILLER_0_24_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vdd vss FILLER_0_24_63/VPW vdd FILLER_0_24_63/a_36_472# FILLER_0_24_63/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ vdd vss _043_ net27 mask\[0\] _189_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_327_ _131_ vdd vss _016_ _127_ _130_ _327_/VPW vdd _327_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ vss _079_ _078_ vdd _258_/VPW vdd _258_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_171 vdd vss FILLER_0_18_171/VPW vdd FILLER_0_18_171/a_36_472# FILLER_0_18_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_130 vdd vss FILLER_0_24_130/VPW vdd FILLER_0_24_130/a_36_472# FILLER_0_24_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__A1 vss _053_ vdd ANTENNA__377__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_133 vdd vss FILLER_0_21_133/VPW vdd FILLER_0_21_133/a_36_472# FILLER_0_21_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_138 vdd vss FILLER_0_8_138/VPW vdd FILLER_0_8_138/a_36_472# FILLER_0_8_138/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_127 vdd vss FILLER_0_8_127/VPW vdd FILLER_0_8_127/a_36_472# FILLER_0_8_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 ctlp[5] net22 vdd vss output22/VPW vdd output22/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 result[6] net33 vdd vss output33/VPW vdd output33/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 trimb[1] net44 vdd vss output44/VPW vdd output44/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 ctln[4] net11 vdd vss output11/VPW vdd output11/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 ctln[2] net9 vdd vss output9/VPW vdd output9/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__194__I vss net18 vdd ANTENNA__194__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ vss _104_ _092_ vdd _291_/VPW vdd _291_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_152 vdd vss FILLER_0_4_152/VPW vdd FILLER_0_4_152/a_36_472# FILLER_0_4_152/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vss FILLER_0_4_185/VPW vdd FILLER_0_4_185/a_36_472# FILLER_0_4_185/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ vss _153_ _152_ vdd _360_/VPW vdd _360_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_65 vdd vss FILLER_0_13_65/VPW vdd FILLER_0_13_65/a_36_472# FILLER_0_13_65/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_343_ _137_ mask\[4\] vdd vss _143_ mask\[3\] _141_ _343_/VPW vdd _343_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_274_ _072_ _090_ vdd vss _091_ net4 _060_ _274_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_412_ _001_ cal_itt\[1\] net58 vss net75 vdd _412_/VPW vdd _412_/a_2665_112# _412_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__292__I vss _098_ vdd ANTENNA__292__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_326_ _131_ vss vdd _125_ _326_/VPW vdd _326_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_257_ _077_ vdd vss _078_ _053_ _075_ _257_/VPW vdd _257_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_309_ vss _116_ net4 vdd _309_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__197__I vss net19 vdd ANTENNA__197__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__301__A2 vss _098_ vdd ANTENNA__301__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vss FILLER_0_15_142/VPW vdd FILLER_0_15_142/a_36_472# FILLER_0_15_142/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 ctlp[6] net23 vdd vss output23/VPW vdd output23/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 trimb[2] net45 vdd vss output45/VPW vdd output45/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput34 result[7] net34 vdd vss output34/VPW vdd output34/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput12 ctln[5] net12 vdd vss output12/VPW vdd output12/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_109 vdd vss FILLER_0_5_109/VPW vdd FILLER_0_5_109/a_36_472# FILLER_0_5_109/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_226 vdd vss FILLER_0_17_226/VPW vdd FILLER_0_17_226/a_36_472# FILLER_0_17_226/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_197 vdd vss FILLER_0_4_197/VPW vdd FILLER_0_4_197/a_36_472# FILLER_0_4_197/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_290_ vdd vss _007_ _094_ _103_ _290_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_223 vdd vss FILLER_0_9_223/VPW vdd FILLER_0_9_223/a_36_472# FILLER_0_9_223/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_342_ vdd vss _142_ _020_ _342_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_273_ vss _090_ state\[0\] vdd _273_/VPW vdd _273_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_411_ _000_ cal_itt\[0\] net58 vss net75 vdd _411_/VPW vdd _411_/a_2665_112# _411_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout80 vss net80 net81 vdd fanout80/VPW vdd fanout80/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_325_ vdd vss _130_ _118_ _129_ _325_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_78 vdd vss FILLER_0_10_78/VPW vdd FILLER_0_10_78/a_36_472# FILLER_0_10_78/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_256_ _056_ _068_ vdd vss _077_ net4 _076_ _256_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_308_ _058_ vdd vss _115_ trim_mask\[0\] _114_ _308_/VPW vdd _308_/a_848_380# vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_98 vdd vss FILLER_0_1_98/VPW vdd FILLER_0_1_98/a_36_472# FILLER_0_1_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ net41 vss vdd _065_ _239_/VPW vdd _239_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_124 vdd vss FILLER_0_12_124/VPW vdd FILLER_0_12_124/a_36_472# FILLER_0_12_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss FILLER_0_8_107/VPW vdd FILLER_0_8_107/a_36_472# FILLER_0_8_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 ctlp[7] net24 vdd vss output24/VPW vdd output24/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 result[8] net35 vdd vss output35/VPW vdd output35/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 trimb[3] net46 vdd vss output46/VPW vdd output46/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vss FILLER_0_18_2/VPW vdd FILLER_0_18_2/a_3260_375# FILLER_0_18_2/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 ctln[6] net13 vdd vss output13/VPW vdd output13/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_162 vdd vss FILLER_0_7_162/VPW vdd FILLER_0_7_162/a_36_472# FILLER_0_7_162/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_195 vdd vss FILLER_0_7_195/VPW vdd FILLER_0_7_195/a_36_472# FILLER_0_7_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I vss cal vdd ANTENNA_input1_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__RN vss net59 vdd ANTENNA__414__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_341_ _137_ mask\[3\] vdd vss _142_ mask\[2\] _141_ _341_/VPW vdd _341_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_410_ vdd _188_ _187_ _042_ _120_ vss _410_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_272_ _089_ vdd vss _003_ _079_ _087_ _272_/VPW vdd _272_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout70 vss net70 net73 vdd fanout70/VPW vdd fanout70/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ _076_ vss vdd _057_ _255_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_324_ vdd vss _129_ calibrate _062_ _324_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output40_I vss net40 vdd ANTENNA_output40_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 vss net81 net82 vdd fanout81/VPW vdd fanout81/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_55 vdd vss FILLER_0_19_55/VPW vdd FILLER_0_19_55/a_36_472# FILLER_0_19_55/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A1 vss _093_ vdd ANTENNA__304__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_307_ vdd vss _114_ _113_ _096_ _307_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_238_ vdd vss _065_ trim_mask\[3\] trim_val\[3\] _238_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_125 vdd vss FILLER_0_21_125/VPW vdd FILLER_0_21_125/a_36_472# FILLER_0_21_125/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_89 vdd vss FILLER_0_16_89/VPW vdd FILLER_0_16_89/a_36_472# FILLER_0_16_89/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_136 vdd vss FILLER_0_12_136/VPW vdd FILLER_0_12_136/a_36_472# FILLER_0_12_136/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 ctlp[8] net25 vdd vss output25/VPW vdd output25/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput47 trimb[4] net47 vdd vss output47/VPW vdd output47/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 result[9] net36 vdd vss output36/VPW vdd output36/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 ctln[7] net14 vdd vss output14/VPW vdd output14/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_144 vdd vss FILLER_0_4_144/VPW vdd FILLER_0_4_144/a_36_472# FILLER_0_4_144/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vss FILLER_0_4_177/VPW vdd FILLER_0_4_177/a_36_472# FILLER_0_4_177/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_340_ vss _141_ _140_ vdd _340_/VPW vdd _340_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_271_ vdd vss cal_itt\[3\] _089_ _271_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__356__B vss _093_ vdd ANTENNA__356__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_256 vdd vss FILLER_0_10_256/VPW vdd FILLER_0_10_256/a_36_472# FILLER_0_10_256/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__200__I vss net20 vdd ANTENNA__200__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I vss net57 vdd ANTENNA_fanout52_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_99 vdd vss FILLER_0_4_99/VPW vdd FILLER_0_4_99/a_36_472# FILLER_0_4_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vss FILLER_0_6_239/VPW vdd FILLER_0_6_239/a_36_472# FILLER_0_6_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout71 vss net71 net73 vdd fanout71/VPW vdd fanout71/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 net60 vss vdd net61 fanout60/VPW vdd fanout60/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_323_ vss _015_ _128_ vdd _323_/VPW vdd _323_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout82 vss net82 net2 vdd fanout82/VPW vdd fanout82/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_254_ _074_ vdd vss _075_ cal_itt\[3\] _072_ _254_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_237_ vdd vss net40 net45 _237_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_306_ vss _113_ _057_ vdd _306_/VPW vdd _306_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_57 vdd vss FILLER_0_16_57/VPW vdd FILLER_0_16_57/a_36_472# FILLER_0_16_57/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput26 ctlp[9] net26 vdd vss output26/VPW vdd output26/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput15 ctln[8] net15 vdd vss output15/VPW vdd output15/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput48 valid net48 vdd vss output48/VPW vdd output48/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput37 sample net37 vdd vss output37/VPW vdd output37/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_17_218 vdd vss FILLER_0_17_218/VPW vdd FILLER_0_17_218/a_36_472# FILLER_0_17_218/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_123 vdd vss FILLER_0_4_123/VPW vdd FILLER_0_4_123/a_36_472# FILLER_0_4_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I vss net21 vdd ANTENNA__203__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _088_ vdd vss _002_ _079_ _087_ _270_/VPW vdd _270_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ vdd vss _179_ cal_count\[1\] _178_ _399_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_322_ _127_ vdd vss _128_ _068_ _124_ _322_/VPW vdd _322_/a_848_380# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout61 vss net61 net62 vdd fanout61/VPW vdd fanout61/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 vss net72 net74 vdd fanout72/VPW vdd fanout72/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd vss FILLER_0_10_37/VPW vdd FILLER_0_10_37/a_36_472# FILLER_0_10_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net50 vss vdd net52 fanout50/VPW vdd fanout50/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_253_ cal_itt\[2\] vdd vss _074_ cal_itt\[0\] cal_itt\[1\] _253_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_305_ vdd vss _112_ net1 _081_ _305_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_236_ net40 vss vdd _064_ _236_/VPW vdd _236_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__206__I vss net22 vdd ANTENNA__206__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vss FILLER_0_20_193/VPW vdd FILLER_0_20_193/a_36_472# FILLER_0_20_193/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ vss _053_ trim_mask\[0\] vdd _219_/VPW vdd _219_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 result[0] net27 vdd vss output27/VPW vdd output27/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput16 ctln[9] net16 vdd vss output16/VPW vdd output16/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 trim[0] net38 vdd vss output38/VPW vdd output38/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_16_241 vdd vss FILLER_0_16_241/VPW vdd FILLER_0_16_241/a_36_472# FILLER_0_16_241/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_398_ vss _178_ net3 vdd _398_/VPW vdd _398_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_247 vdd vss FILLER_0_10_247/VPW vdd FILLER_0_10_247/a_36_472# FILLER_0_10_247/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_214 vdd vss FILLER_0_10_214/VPW vdd FILLER_0_10_214/a_36_472# FILLER_0_10_214/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_91 vdd vss FILLER_0_14_91/VPW vdd FILLER_0_14_91/a_36_472# FILLER_0_14_91/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__209__I vss net23 vdd ANTENNA__209__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I vss net19 vdd ANTENNA_output19_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_47 vdd vss FILLER_0_19_47/VPW vdd FILLER_0_19_47/a_36_472# FILLER_0_19_47/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout73 vss net73 net74 vdd fanout73/VPW vdd fanout73/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout62 net62 vss vdd net64 fanout62/VPW vdd fanout62/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout51 vss net51 net52 vdd fanout51/VPW vdd fanout51/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ _076_ _125_ _126_ vdd vss _127_ _069_ _321_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_252_ vdd vss cal_itt\[0\] _073_ _252_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_100 vdd vss FILLER_0_18_100/VPW vdd FILLER_0_18_100/a_36_472# FILLER_0_18_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss FILLER_0_18_177/VPW vdd FILLER_0_18_177/a_3260_375# FILLER_0_18_177/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_304_ vdd vss _013_ _093_ _111_ _304_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_235_ vdd vss _064_ trim_mask\[2\] trim_val\[2\] _235_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_218_ vss net16 net26 vdd _218_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_37 vdd vss FILLER_0_16_37/VPW vdd FILLER_0_16_37/a_36_472# FILLER_0_16_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput17 ctlp[0] net17 vdd vss output17/VPW vdd output17/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 result[1] net28 vdd vss output28/VPW vdd output28/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput39 trim[1] net39 vdd vss output39/VPW vdd output39/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_212 vdd vss FILLER_0_13_212/VPW vdd FILLER_0_13_212/a_36_472# FILLER_0_13_212/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_397_ _177_ vdd vss _040_ _131_ _175_ _397_/VPW vdd _397_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_81 vdd vss FILLER_0_14_81/VPW vdd FILLER_0_14_81/a_36_472# FILLER_0_14_81/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout63 net63 vss vdd net64 fanout63/VPW vdd fanout63/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_320_ _096_ vdd vss _126_ mask\[0\] _113_ _320_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_28 vdd vss FILLER_0_10_28/VPW vdd FILLER_0_10_28/a_36_472# FILLER_0_10_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout74 vss net74 net82 vdd fanout74/VPW vdd fanout74/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net52 vss vdd net57 fanout52/VPW vdd fanout52/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_251_ _072_ vdd vss net48 _068_ _070_ _251_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_449_ _038_ en_co_clk net55 vss net72 vdd _449_/VPW vdd _449_/a_2665_112# _449_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_303_ net36 vdd vss _111_ mask\[9\] _098_ _303_/VPW vdd _303_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ vss net44 net39 vdd _234_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_217_ vss net26 _052_ vdd _217_/VPW vdd _217_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_181 vdd vss FILLER_0_14_181/VPW vdd FILLER_0_14_181/a_36_472# FILLER_0_14_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 ctlp[1] net18 vdd vss output18/VPW vdd output18/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput29 result[2] net29 vdd vss output29/VPW vdd output29/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_fanout80_I vss net81 vdd ANTENNA_fanout80_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_396_ vdd vss _177_ cal_count\[1\] _176_ _396_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout53 net53 vss vdd net56 fanout53/VPW vdd fanout53/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_250_ vss _072_ _071_ vdd _250_/VPW vdd _250_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout75 vss net75 net76 vdd fanout75/VPW vdd fanout75/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout64 vss net64 net65 vdd fanout64/VPW vdd fanout64/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_448_ _037_ trim_val\[4\] net59 vss net76 vdd _448_/VPW vdd _448_/a_2665_112# _448_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ trim_val\[1\] vdd vss _166_ trim_mask\[1\] _164_ _379_/VPW vdd _379_/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_302_ vdd vss _012_ _093_ _110_ _302_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_28 vdd vss FILLER_0_21_28/VPW vdd FILLER_0_21_28/a_3260_375# FILLER_0_21_28/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__216__A2 vss net36 vdd ANTENNA__216__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ vss net39 _063_ vdd _233_/VPW vdd _233_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_116 vdd vss FILLER_0_15_116/VPW vdd FILLER_0_15_116/a_36_472# FILLER_0_15_116/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__373__A1 vss cal_count\[3\] vdd ANTENNA__373__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_216_ vdd vss _052_ mask\[9\] net36 _216_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_146 vdd vss FILLER_0_7_146/VPW vdd FILLER_0_7_146/a_36_472# FILLER_0_7_146/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 ctlp[2] net19 vdd vss output19/VPW vdd output19/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_59 vdd vss FILLER_0_7_59/VPW vdd FILLER_0_7_59/a_36_472# FILLER_0_7_59/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_255 vdd vss FILLER_0_16_255/VPW vdd FILLER_0_16_255/a_36_472# FILLER_0_16_255/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_130 vdd vss FILLER_0_0_130/VPW vdd FILLER_0_0_130/a_36_472# FILLER_0_0_130/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_263 vdd vss FILLER_0_8_263/VPW vdd FILLER_0_8_263/a_36_472# FILLER_0_8_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_50 vdd vss FILLER_0_14_50/VPW vdd FILLER_0_14_50/a_36_472# FILLER_0_14_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_395_ _070_ _085_ vdd vss _176_ _116_ _072_ _395_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_4_49 vdd vss FILLER_0_4_49/VPW vdd FILLER_0_4_49/a_36_472# FILLER_0_4_49/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout54 net54 vss vdd net56 fanout54/VPW vdd fanout54/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout76 vss net76 net81 vdd fanout76/VPW vdd fanout76/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout65 vss net65 net5 vdd fanout65/VPW vdd fanout65/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_28 vdd vss FILLER_0_19_28/VPW vdd FILLER_0_19_28/a_36_472# FILLER_0_19_28/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_447_ _036_ trim_val\[3\] net50 vss net68 vdd _447_/VPW vdd _447_/a_2665_112# _447_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_2 vdd vss FILLER_0_3_2/VPW vdd FILLER_0_3_2/a_36_472# FILLER_0_3_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_378_ vdd vss _033_ _160_ _165_ _378_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_301_ net35 vdd vss _110_ mask\[8\] _098_ _301_/VPW vdd _301_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output17_I vss net17 vdd ANTENNA_output17_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_232_ vdd vss _063_ trim_mask\[1\] trim_val\[1\] _232_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_215_ vss net15 net25 vdd _215_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_142 vdd vss FILLER_0_11_142/VPW vdd FILLER_0_11_142/a_36_472# FILLER_0_11_142/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_93 vdd vss FILLER_0_2_93/VPW vdd FILLER_0_2_93/a_36_472# FILLER_0_2_93/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_72 vdd vss FILLER_0_17_72/VPW vdd FILLER_0_17_72/a_3260_375# FILLER_0_17_72/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_172 vdd vss FILLER_0_3_172/VPW vdd FILLER_0_3_172/a_3260_375# FILLER_0_3_172/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output47_I vss net47 vdd ANTENNA_output47_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _095_ vdd vss _175_ _174_ cal_count\[1\] _394_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xfanout55 net55 vss vdd net57 fanout55/VPW vdd fanout55/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_212 vdd vss FILLER_0_5_212/VPW vdd FILLER_0_5_212/a_36_472# FILLER_0_5_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout77 vss net77 net78 vdd fanout77/VPW vdd fanout77/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_446_ _035_ trim_val\[2\] net49 vss net66 vdd _446_/VPW vdd _446_/a_2665_112# _446_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout66 vss net66 net68 vdd fanout66/VPW vdd fanout66/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_377_ trim_val\[0\] vdd vss _165_ _053_ _164_ _377_/VPW vdd _377_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_300_ vdd vss _011_ _104_ _109_ _300_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_231_ vdd vss net37 _059_ _062_ _231_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_429_ _018_ mask\[0\] net62 vss net79 vdd _429_/VPW vdd _429_/a_2665_112# _429_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput1 vss net1 cal vdd input1/VPW vdd input1/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ vss net25 _051_ vdd _214_/VPW vdd _214_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_104 vdd vss FILLER_0_7_104/VPW vdd FILLER_0_7_104/a_36_472# FILLER_0_7_104/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vdd vss FILLER_0_4_107/VPW vdd FILLER_0_4_107/a_36_472# FILLER_0_4_107/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_290 vdd vss FILLER_0_24_290/VPW vdd FILLER_0_24_290/a_36_472# FILLER_0_24_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_290 vdd vss FILLER_0_15_290/VPW vdd FILLER_0_15_290/a_36_472# FILLER_0_15_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_198 vdd vss FILLER_0_0_198/VPW vdd FILLER_0_0_198/a_36_472# FILLER_0_0_198/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_393_ vdd vss cal_count\[0\] _174_ _393_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout78 vss net78 net79 vdd fanout78/VPW vdd fanout78/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 vss net56 net57 vdd fanout56/VPW vdd fanout56/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout67 vss net67 net68 vdd fanout67/VPW vdd fanout67/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_445_ _034_ trim_val\[1\] net49 vss net66 vdd _445_/VPW vdd _445_/a_2665_112# _445_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_376_ vss _164_ _163_ vdd _376_/VPW vdd _376_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_230_ vdd vss _062_ _060_ _061_ _230_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vss FILLER_0_5_72/VPW vdd FILLER_0_5_72/a_36_472# FILLER_0_5_72/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_428_ _017_ state\[2\] net53 vss net70 vdd _428_/VPW vdd _428_/a_2665_112# _428_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_11_64 vdd vss FILLER_0_11_64/VPW vdd FILLER_0_11_64/a_36_472# FILLER_0_11_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_359_ _131_ _129_ vdd vss _152_ _059_ _062_ _359_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput2 vss net2 clk vdd input2/VPW vdd input2/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output22_I vss net22 vdd ANTENNA_output22_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_213_ vdd vss _051_ mask\[8\] net35 _213_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_177 vdd vss FILLER_0_20_177/VPW vdd FILLER_0_20_177/a_36_472# FILLER_0_20_177/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_206 vdd vss FILLER_0_13_206/VPW vdd FILLER_0_13_206/a_36_472# FILLER_0_13_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_228 vdd vss FILLER_0_13_228/VPW vdd FILLER_0_13_228/a_36_472# FILLER_0_13_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_392_ vdd _173_ _077_ _039_ cal_count\[0\] vss _392_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__282__I vss _098_ vdd ANTENNA__282__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 vss net79 net81 vdd fanout79/VPW vdd fanout79/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_2 vdd vss FILLER_0_12_2/VPW vdd FILLER_0_12_2/a_36_472# FILLER_0_12_2/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout68 vss net68 net69 vdd fanout68/VPW vdd fanout68/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout57 vss net57 net65 vdd fanout57/VPW vdd fanout57/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _033_ trim_val\[0\] net50 vss net67 vdd _444_/VPW vdd _444_/a_2665_112# _444_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_375_ _074_ _161_ _162_ vdd vss _163_ cal_itt\[3\] _375_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__277__I vss _093_ vdd ANTENNA__277__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_139 vdd vss FILLER_0_18_139/VPW vdd FILLER_0_18_139/a_36_472# FILLER_0_18_139/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_161 vdd vss FILLER_0_17_161/VPW vdd FILLER_0_17_161/a_36_472# FILLER_0_17_161/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ _016_ state\[1\] net53 vdd vss net70 _427_/VPW vdd _427_/a_36_151# vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_358_ vdd vss _053_ _151_ _358_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__385__A2 vss net47 vdd ANTENNA__385__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_289_ net30 vdd vss _103_ mask\[3\] _099_ _289_/VPW vdd _289_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput3 vss net3 comp vdd input3/VPW vdd input3/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_212_ vss net14 net24 vdd _212_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_output15_I vss net15 vdd ANTENNA_output15_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vss FILLER_0_22_86/VPW vdd FILLER_0_22_86/a_36_472# FILLER_0_22_86/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_101 vdd vss FILLER_0_11_101/VPW vdd FILLER_0_11_101/a_36_472# FILLER_0_11_101/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_64 vdd vss FILLER_0_17_64/VPW vdd FILLER_0_17_64/a_36_472# FILLER_0_17_64/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_142 vdd vss FILLER_0_3_142/VPW vdd FILLER_0_3_142/a_36_472# FILLER_0_3_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_391_ vdd vss _173_ cal_count\[0\] _120_ _391_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 vss net69 net74 vdd fanout69/VPW vdd fanout69/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net58 vss vdd net59 fanout58/VPW vdd fanout58/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_374_ vdd _061_ _056_ _162_ calibrate vss _374_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_443_ _032_ trim_mask\[4\] net52 vss net69 vdd _443_/VPW vdd _443_/a_2665_112# _443_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_107 vdd vss FILLER_0_18_107/VPW vdd FILLER_0_18_107/a_3260_375# FILLER_0_18_107/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__394__A3 vss _095_ vdd ANTENNA__394__A3/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ vdd vss _006_ _094_ _102_ _288_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_357_ vdd vss _150_ _027_ _357_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ _015_ state\[0\] net64 vss net81 vdd _426_/VPW vdd _426_/a_2665_112# _426_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput4 vss net4 en vdd input4/VPW vdd input4/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_211_ vss net24 _050_ vdd _211_/VPW vdd _211_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_409_ vdd vss _188_ cal_count\[3\] _077_ _409_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_135 vdd vss FILLER_0_11_135/VPW vdd FILLER_0_11_135/a_36_472# FILLER_0_11_135/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vss FILLER_0_11_124/VPW vdd FILLER_0_11_124/a_36_472# FILLER_0_11_124/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vss FILLER_0_15_282/VPW vdd FILLER_0_15_282/a_36_472# FILLER_0_15_282/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__RN vss net59 vdd ANTENNA__413__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ _136_ _172_ _067_ vdd vss _038_ _070_ _390_/VPW vdd _390_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_14_99 vdd vss FILLER_0_14_99/VPW vdd FILLER_0_14_99/a_36_472# FILLER_0_14_99/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout59 net59 vss vdd net64 fanout59/VPW vdd fanout59/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_373_ _056_ _113_ vdd vss _161_ cal_count\[3\] _090_ _373_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_442_ _031_ trim_mask\[3\] net52 vss net69 vdd _442_/VPW vdd _442_/a_2665_112# _442_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_356_ _093_ vdd vss _150_ mask\[9\] _136_ _356_/VPW vdd _356_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_287_ net29 vdd vss _102_ mask\[2\] _099_ _287_/VPW vdd _287_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_78 vdd vss FILLER_0_11_78/VPW vdd FILLER_0_11_78/a_36_472# FILLER_0_11_78/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 vss net5 rstn vdd input5/VPW vdd input5/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _014_ calibrate net58 vss net75 vdd _425_/VPW vdd _425_/a_2665_112# _425_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_210_ vdd vss _050_ mask\[7\] net34 _210_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_169 vdd vss FILLER_0_20_169/VPW vdd FILLER_0_20_169/a_36_472# FILLER_0_20_169/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _186_ vdd vss _187_ _095_ cal_count\[3\] _408_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_339_ vss _140_ _091_ vdd _339_/VPW vdd _339_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output20_I vss net20 vdd ANTENNA_output20_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_286 vdd vss FILLER_0_21_286/VPW vdd FILLER_0_21_286/a_36_472# FILLER_0_21_286/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_220 vdd vss FILLER_0_12_220/VPW vdd FILLER_0_12_220/a_36_472# FILLER_0_12_220/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_247 vdd vss FILLER_0_8_247/VPW vdd FILLER_0_8_247/a_36_472# FILLER_0_8_247/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 net49 vss vdd net50 fanout49/VPW vdd fanout49/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_206 vdd vss FILLER_0_5_206/VPW vdd FILLER_0_5_206/a_36_472# FILLER_0_5_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ _030_ trim_mask\[2\] net49 vss net66 vdd _441_/VPW vdd _441_/a_2665_112# _441_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_372_ _070_ _076_ _068_ vdd vss _160_ _133_ _372_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__303__A2 vss _098_ vdd ANTENNA__303__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vss FILLER_0_17_142/VPW vdd FILLER_0_17_142/a_36_472# FILLER_0_17_142/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_54 vdd vss FILLER_0_5_54/VPW vdd FILLER_0_5_54/a_36_472# FILLER_0_5_54/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_355_ vdd vss _149_ _026_ _355_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_424_ _013_ net36 net55 vss net72 vdd _424_/VPW vdd _424_/a_2665_112# _424_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_286_ vdd vss _005_ _094_ _101_ _286_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_123 vdd vss FILLER_0_14_123/VPW vdd FILLER_0_14_123/a_36_472# FILLER_0_14_123/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ vdd vss _139_ _019_ _338_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_407_ _185_ vdd vss _186_ _181_ _184_ _407_/VPW vdd _407_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_269_ cal_itt\[2\] vdd vss _088_ _083_ _078_ _269_/VPW vdd _269_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_56 vdd vss FILLER_0_17_56/VPW vdd FILLER_0_17_56/a_36_472# FILLER_0_17_56/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I vss en vdd ANTENNA_input4_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ vss _032_ _159_ vdd _371_/VPW vdd _371_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_440_ _029_ trim_mask\[1\] net49 vss net66 vdd _440_/VPW vdd _440_/a_2665_112# _440_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_5_88 vdd vss FILLER_0_5_88/VPW vdd FILLER_0_5_88/a_36_472# FILLER_0_5_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ _012_ net35 net55 vss net72 vdd _423_/VPW vdd _423_/a_2665_112# _423_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_354_ _132_ mask\[9\] vdd vss _149_ mask\[8\] _140_ _354_/VPW vdd _354_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_285_ net28 vdd vss _101_ mask\[1\] _099_ _285_/VPW vdd _285_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_199_ net20 vss vdd _046_ _199_/VPW vdd _199_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_337_ _137_ mask\[2\] vdd vss _139_ mask\[1\] _136_ _337_/VPW vdd _337_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_406_ vdd vss _185_ _178_ cal_count\[2\] _406_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_268_ vdd vss _087_ _086_ _074_ _268_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_274 vdd vss FILLER_0_24_274/VPW vdd FILLER_0_24_274/a_36_472# FILLER_0_24_274/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ _152_ vdd vss _159_ trim_mask\[4\] _081_ _370_/VPW vdd _370_/a_848_380# vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout55_I vss net57 vdd ANTENNA_fanout55_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_266 vdd vss FILLER_0_1_266/VPW vdd FILLER_0_1_266/a_36_472# FILLER_0_1_266/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_422_ _011_ net34 net61 vss net78 vdd _422_/VPW vdd _422_/a_2665_112# _422_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_353_ vdd vss _148_ _025_ _353_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_133 vdd vss FILLER_0_17_133/VPW vdd FILLER_0_17_133/a_36_472# FILLER_0_17_133/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output36_I vss net36 vdd ANTENNA_output36_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_284_ vdd vss _004_ _094_ _100_ _284_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_198_ vdd vss _046_ mask\[3\] net30 _198_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_336_ vdd vss _138_ _018_ _336_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_405_ vdd vss _184_ _178_ cal_count\[2\] _405_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _071_ vdd vss _086_ _085_ state\[1\] _267_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_6_177 vdd vss FILLER_0_6_177/VPW vdd FILLER_0_6_177/a_36_472# FILLER_0_6_177/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_319_ vdd vss _125_ _058_ _119_ _319_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_239 vdd vss FILLER_0_8_239/VPW vdd FILLER_0_8_239/a_36_472# FILLER_0_8_239/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss FILLER_0_1_212/VPW vdd FILLER_0_1_212/a_36_472# FILLER_0_1_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _010_ net33 net60 vss net77 vdd _421_/VPW vdd _421_/a_2665_112# _421_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_352_ _144_ mask\[8\] vdd vss _148_ mask\[7\] _140_ _352_/VPW vdd _352_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_283_ net27 vdd vss _100_ mask\[0\] _099_ _283_/VPW vdd _283_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vdd vss FILLER_0_9_142/VPW vdd FILLER_0_9_142/a_36_472# FILLER_0_9_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vss FILLER_0_20_107/VPW vdd FILLER_0_20_107/a_36_472# FILLER_0_20_107/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_404_ _183_ vdd vss _041_ _131_ _182_ _404_/VPW vdd _404_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_335_ _137_ mask\[1\] vdd vss _138_ mask\[0\] _136_ _335_/VPW vdd _335_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_266_ vdd vss _055_ _085_ _266_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_197_ vdd vss net19 net9 _197_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_249_ vss _071_ state\[2\] vdd _249_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__409__A1 vss cal_count\[3\] vdd ANTENNA__409__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_318_ vdd vss _124_ _115_ _118_ _318_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_24 vdd vss FILLER_0_8_24/VPW vdd FILLER_0_8_24/a_36_472# FILLER_0_8_24/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__251__A2 vss _070_ vdd ANTENNA__251__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss FILLER_0_8_2/VPW vdd FILLER_0_8_2/a_36_472# FILLER_0_8_2/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss clk vdd ANTENNA_input2_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _009_ net32 net60 vss net77 vdd _420_/VPW vdd _420_/a_2665_112# _420_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_351_ vdd vss _147_ _024_ _351_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_282_ vss _099_ _098_ vdd _282_/VPW vdd _282_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__390__A1 vss _070_ vdd ANTENNA__390__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_334_ vss _137_ _132_ vdd _334_/VPW vdd _334_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_403_ vdd vss _183_ cal_count\[2\] _176_ _403_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output41_I vss net41 vdd ANTENNA_output41_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vss FILLER_0_6_90/VPW vdd FILLER_0_6_90/a_36_472# FILLER_0_6_90/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net19 vss vdd _045_ _196_/VPW vdd _196_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_265_ _084_ _079_ _082_ vdd vss _001_ _081_ _083_ _265_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__395__B vss _070_ vdd ANTENNA__395__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd vss FILLER_0_17_38/VPW vdd FILLER_0_17_38/a_36_472# FILLER_0_17_38/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_248_ vss _070_ _069_ vdd _248_/VPW vdd _248_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__409__A2 vss _077_ vdd ANTENNA__409__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ vss _014_ _123_ vdd _317_/VPW vdd _317_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_171 vdd vss FILLER_0_2_171/VPW vdd FILLER_0_2_171/a_36_472# FILLER_0_2_171/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_236 vdd vss FILLER_0_12_236/VPW vdd FILLER_0_12_236/a_36_472# FILLER_0_12_236/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_350_ _144_ mask\[7\] vdd vss _147_ mask\[6\] _140_ _350_/VPW vdd _350_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_281_ vdd vss _098_ _091_ _097_ _281_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__237__I vss net40 vdd ANTENNA__237__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_333_ vss _136_ _091_ vdd _333_/VPW vdd _333_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_195_ vdd vss _045_ mask\[2\] net29 _195_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_402_ _181_ vdd vss _182_ _095_ cal_count\[2\] _402_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_11_109 vdd vss FILLER_0_11_109/VPW vdd FILLER_0_11_109/a_36_472# FILLER_0_11_109/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_264_ vdd vss _084_ cal_itt\[0\] cal_itt\[1\] _264_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__372__A2 vss _070_ vdd ANTENNA__372__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_50 vdd vss FILLER_0_12_50/VPW vdd FILLER_0_12_50/a_36_472# FILLER_0_12_50/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_247_ _069_ vss vdd _060_ _247_/VPW vdd _247_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_316_ _122_ vdd vss _123_ _112_ calibrate _316_/VPW vdd _316_/a_848_380# vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_60 vdd vss FILLER_0_23_60/VPW vdd FILLER_0_23_60/a_36_472# FILLER_0_23_60/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vss FILLER_0_15_212/VPW vdd FILLER_0_15_212/a_36_472# FILLER_0_15_212/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vss FILLER_0_8_37/VPW vdd FILLER_0_8_37/a_36_472# FILLER_0_8_37/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_104 vdd vss FILLER_0_17_104/VPW vdd FILLER_0_17_104/a_36_472# FILLER_0_17_104/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_72 vdd vss FILLER_0_15_72/VPW vdd FILLER_0_15_72/a_36_472# FILLER_0_15_72/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_204 vdd vss FILLER_0_1_204/VPW vdd FILLER_0_1_204/a_36_472# FILLER_0_1_204/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_280_ vdd vss _097_ _095_ _096_ _280_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_107 vdd vss FILLER_0_14_107/VPW vdd FILLER_0_14_107/a_36_472# FILLER_0_14_107/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_401_ vdd _180_ _179_ _181_ _174_ vss _401_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_332_ _126_ vdd vss _017_ _127_ _135_ _332_/VPW vdd _332_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_194_ vss net8 net18 vdd _194_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_263_ vdd vss _083_ _073_ _082_ _263_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_181 vdd vss FILLER_0_5_181/VPW vdd FILLER_0_5_181/a_36_472# FILLER_0_5_181/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_246_ vss _068_ _055_ vdd _246_/VPW vdd _246_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_315_ _118_ _122_ _115_ _120_ _121_ vdd vss _315_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_290 vdd vss FILLER_0_23_290/VPW vdd FILLER_0_23_290/a_36_472# FILLER_0_23_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_235 vdd vss FILLER_0_15_235/VPW vdd FILLER_0_15_235/a_36_472# FILLER_0_15_235/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_229_ vdd vss _061_ _055_ _057_ _229_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_61 vdd vss FILLER_0_18_61/VPW vdd FILLER_0_18_61/a_36_472# FILLER_0_18_61/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vss FILLER_0_11_282/VPW vdd FILLER_0_11_282/a_36_472# FILLER_0_11_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I vss net81 vdd ANTENNA_fanout76_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_213 vdd vss FILLER_0_4_213/VPW vdd FILLER_0_4_213/a_36_472# FILLER_0_4_213/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_400_ vdd vss _180_ cal_count\[1\] _178_ _400_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_193_ net18 vss vdd _044_ _193_/VPW vdd _193_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_331_ _134_ vdd vss _135_ _086_ _132_ _331_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_262_ vdd vss cal_itt\[1\] _082_ _262_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__303__B vss net36 vdd ANTENNA__303__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ vdd vss _121_ _085_ _069_ _314_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_245_ vdd vss net6 _067_ net67 _245_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_206 vdd vss FILLER_0_21_206/VPW vdd FILLER_0_21_206/a_36_472# FILLER_0_21_206/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_228_ vss _060_ state\[1\] vdd _228_/VPW vdd _228_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_233 vdd vss FILLER_0_7_233/VPW vdd FILLER_0_7_233/a_36_472# FILLER_0_7_233/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_60 vdd vss FILLER_0_9_60/VPW vdd FILLER_0_9_60/a_36_472# FILLER_0_9_60/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vss FILLER_0_13_142/VPW vdd FILLER_0_13_142/a_36_472# FILLER_0_13_142/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ vdd vss _044_ mask\[1\] net28 _192_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_261_ vss _081_ _059_ vdd _261_/VPW vdd _261_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_330_ vdd vss _134_ _133_ _062_ _330_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_20 vdd vss FILLER_0_12_20/VPW vdd FILLER_0_12_20/a_36_472# FILLER_0_12_20/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_172 vdd vss FILLER_0_5_172/VPW vdd FILLER_0_5_172/a_36_472# FILLER_0_5_172/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ vdd vss en_co_clk _067_ _244_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__190__I vss _043_ vdd ANTENNA__190__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_313_ vdd vss _120_ _059_ _119_ _313_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__257__A1 vss _053_ vdd ANTENNA__257__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_227_ vss _059_ _058_ vdd _227_/VPW vdd _227_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__402__A1 vss _095_ vdd ANTENNA__402__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vss FILLER_0_20_31/VPW vdd FILLER_0_20_31/a_36_472# FILLER_0_20_31/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vss FILLER_0_9_72/VPW vdd FILLER_0_9_72/a_36_472# FILLER_0_9_72/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_96 vdd vss FILLER_0_0_96/VPW vdd FILLER_0_0_96/a_36_472# FILLER_0_0_96/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_260_ vdd _080_ _079_ _000_ _073_ vss _260_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _171_ vdd vss _172_ _115_ _120_ _389_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_191_ vdd vss net17 net7 _191_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_312_ vdd vss _119_ cal_itt\[3\] _074_ _312_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_243_ vdd vss net47 net42 _243_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_282 vdd vss FILLER_0_23_282/VPW vdd FILLER_0_23_282/a_36_472# FILLER_0_23_282/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_205 vdd vss FILLER_0_15_205/VPW vdd FILLER_0_15_205/a_36_472# FILLER_0_15_205/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vss FILLER_0_2_165/VPW vdd FILLER_0_2_165/a_36_472# FILLER_0_2_165/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vss FILLER_0_18_53/VPW vdd FILLER_0_18_53/a_36_472# FILLER_0_18_53/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_226_ _057_ vdd vss _058_ _055_ _056_ _226_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__426__CLK vss net81 vdd ANTENNA__426__CLK/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_98 vdd vss FILLER_0_20_98/VPW vdd FILLER_0_20_98/a_36_472# FILLER_0_20_98/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_87 vdd vss FILLER_0_20_87/VPW vdd FILLER_0_20_87/a_36_472# FILLER_0_20_87/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ vdd vss net23 net13 _209_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_171 vdd vss FILLER_0_19_171/VPW vdd FILLER_0_19_171/a_36_472# FILLER_0_19_171/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__302__A1 vss _093_ vdd ANTENNA__302__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_10 vdd vss FILLER_0_15_10/VPW vdd FILLER_0_15_10/a_36_472# FILLER_0_15_10/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vdd vss FILLER_0_15_2/VPW vdd FILLER_0_15_2/a_36_472# FILLER_0_15_2/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vss FILLER_0_22_177/VPW vdd FILLER_0_22_177/a_36_472# FILLER_0_22_177/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_100 vdd vss FILLER_0_13_100/VPW vdd FILLER_0_13_100/a_36_472# FILLER_0_13_100/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_105 vdd vss FILLER_0_9_105/VPW vdd FILLER_0_9_105/a_36_472# FILLER_0_9_105/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ net17 vss vdd _043_ _190_/VPW vdd _190_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_388_ vdd vss _126_ _171_ _388_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output18_I vss net18 vdd ANTENNA_output18_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ _114_ _117_ vdd vss _118_ _116_ _086_ _311_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_242_ net47 vss vdd _066_ _242_/VPW vdd _242_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_228 vdd vss FILLER_0_15_228/VPW vdd FILLER_0_15_228/a_36_472# FILLER_0_15_228/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_111 vdd vss FILLER_0_2_111/VPW vdd FILLER_0_2_111/a_36_472# FILLER_0_2_111/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_177 vdd vss FILLER_0_2_177/VPW vdd FILLER_0_2_177/a_36_472# FILLER_0_2_177/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_225_ vss _057_ state\[2\] vdd _225_/VPW vdd _225_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_76 vdd vss FILLER_0_18_76/VPW vdd FILLER_0_18_76/a_36_472# FILLER_0_18_76/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_208_ net23 vss vdd _049_ _208_/VPW vdd _208_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_387_ vss _037_ _170_ vdd _387_/VPW vdd _387_/a_36_113# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_310_ _090_ vdd vss _117_ _060_ _113_ _310_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_164 vdd vss FILLER_0_5_164/VPW vdd FILLER_0_5_164/a_36_472# FILLER_0_5_164/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_88 vdd vss FILLER_0_23_88/VPW vdd FILLER_0_23_88/a_36_472# FILLER_0_23_88/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_44 vdd vss FILLER_0_23_44/VPW vdd FILLER_0_23_44/a_36_472# FILLER_0_23_44/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_241_ vdd vss _066_ trim_mask\[4\] trim_val\[4\] _241_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_439_ _028_ trim_mask\[0\] net50 vss net67 vdd _439_/VPW vdd _439_/a_2665_112# _439_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_2_101 vdd vss FILLER_0_2_101/VPW vdd FILLER_0_2_101/a_36_472# FILLER_0_2_101/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_54 vdd vss FILLER_0_3_54/VPW vdd FILLER_0_3_54/a_36_472# FILLER_0_3_54/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ vss _056_ state\[1\] vdd _224_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_207_ vdd vss _049_ mask\[6\] net33 _207_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_195 vdd vss FILLER_0_19_195/VPW vdd FILLER_0_19_195/a_36_472# FILLER_0_19_195/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_232 vdd vss FILLER_0_0_232/VPW vdd FILLER_0_0_232/a_36_472# FILLER_0_0_232/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_154 vdd vss FILLER_0_16_154/VPW vdd FILLER_0_16_154/a_36_472# FILLER_0_16_154/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__257__B vss _077_ vdd ANTENNA__257__B/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__220__A2 vss _053_ vdd ANTENNA__220__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vss FILLER_0_20_2/VPW vdd FILLER_0_20_2/a_36_472# FILLER_0_20_2/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_386_ _163_ vdd vss _170_ trim_val\[4\] _169_ _386_/VPW vdd _386_/a_848_380# vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_198 vdd vss FILLER_0_5_198/VPW vdd FILLER_0_5_198/a_36_472# FILLER_0_5_198/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_240_ vdd vss net41 net46 _240_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_282 vdd vss FILLER_0_17_282/VPW vdd FILLER_0_17_282/a_36_472# FILLER_0_17_282/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_274 vdd vss FILLER_0_23_274/VPW vdd FILLER_0_23_274/a_36_472# FILLER_0_23_274/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_438_ _027_ mask\[9\] net54 vss net71 vdd _438_/VPW vdd _438_/a_2665_112# _438_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_369_ _153_ _154_ _158_ vdd vss _031_ _157_ _369_/VPW vdd _369_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output23_I vss net23 vdd ANTENNA_output23_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_263 vdd vss FILLER_0_14_263/VPW vdd FILLER_0_14_263/a_36_472# FILLER_0_14_263/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _055_ vss vdd state\[0\] _223_/VPW vdd _223_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_290 vdd vss FILLER_0_9_290/VPW vdd FILLER_0_9_290/a_36_472# FILLER_0_9_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ vdd vss net22 net12 _206_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_266 vdd vss FILLER_0_0_266/VPW vdd FILLER_0_0_266/a_36_472# FILLER_0_0_266/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ vdd net37 net47 _169_ _081_ vss _385_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_299_ net34 vdd vss _109_ mask\[7\] _105_ _299_/VPW vdd _299_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_437_ _026_ mask\[8\] net54 vss net71 vdd _437_/VPW vdd _437_/a_2665_112# _437_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_3_78 vdd vss FILLER_0_3_78/VPW vdd FILLER_0_3_78/a_36_472# FILLER_0_3_78/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_368_ vdd vss trim_mask\[4\] _158_ _368_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_222_ vdd vss net38 net43 _222_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_205_ net22 vss vdd _048_ _205_/VPW vdd _205_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_142 vdd vss FILLER_0_19_142/VPW vdd FILLER_0_19_142/a_36_472# FILLER_0_19_142/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_453_ _042_ cal_count\[3\] net51 vss net68 vdd _453_/VPW vdd _453_/a_2665_112# _453_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_384_ vdd vss _036_ _160_ _168_ _384_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_107 vdd vss FILLER_0_10_107/VPW vdd FILLER_0_10_107/a_36_472# FILLER_0_10_107/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_298_ vdd vss _010_ _104_ _108_ _298_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_436_ _025_ mask\[7\] net54 vss net71 vdd _436_/VPW vdd _436_/a_2665_112# _436_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A1 vss _095_ vdd ANTENNA__408__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _153_ _154_ _157_ vdd vss _030_ _156_ _367_/VPW vdd _367_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_80 vdd vss FILLER_0_13_80/VPW vdd FILLER_0_13_80/a_36_472# FILLER_0_13_80/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_192 vdd vss FILLER_0_1_192/VPW vdd FILLER_0_1_192/a_36_472# FILLER_0_1_192/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_270 vdd vss FILLER_0_9_270/VPW vdd FILLER_0_9_270/a_36_472# FILLER_0_9_270/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_221_ vss net38 _054_ vdd _221_/VPW vdd _221_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_419_ _008_ net31 net60 vss net77 vdd _419_/VPW vdd _419_/a_2665_112# _419_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_204_ vdd vss _048_ mask\[5\] net32 _204_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_15 vdd vss FILLER_0_20_15/VPW vdd FILLER_0_20_15/a_36_472# FILLER_0_20_15/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_187 vdd vss FILLER_0_19_187/VPW vdd FILLER_0_19_187/a_36_472# FILLER_0_19_187/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_221 vdd vss FILLER_0_3_221/VPW vdd FILLER_0_3_221/a_36_472# FILLER_0_3_221/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_59 vdd vss FILLER_0_15_59/VPW vdd FILLER_0_15_59/a_36_472# FILLER_0_15_59/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I vss net59 vdd ANTENNA_fanout58_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_79 vdd vss FILLER_0_6_79/VPW vdd FILLER_0_6_79/a_36_472# FILLER_0_6_79/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ vss net72 vdd _041_ cal_count\[2\] net55 _452_/VPW vdd _452_/a_36_151# vss
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_383_ trim_val\[3\] vdd vss _168_ trim_mask\[3\] _164_ _383_/VPW vdd _383_/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_297_ net33 vdd vss _108_ mask\[6\] _105_ _297_/VPW vdd _297_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_435_ _024_ mask\[6\] net63 vss net80 vdd _435_/VPW vdd _435_/a_2665_112# _435_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__408__A2 vss cal_count\[3\] vdd ANTENNA__408__A2/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ vdd vss trim_mask\[3\] _157_ _366_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_127 vdd vss FILLER_0_2_127/VPW vdd FILLER_0_2_127/a_36_472# FILLER_0_2_127/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vss FILLER_0_18_37/VPW vdd FILLER_0_18_37/a_36_472# FILLER_0_18_37/a_1468_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_282 vdd vss FILLER_0_9_282/VPW vdd FILLER_0_9_282/a_36_472# FILLER_0_9_282/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_220_ vdd vss _054_ trim_val\[0\] _053_ _220_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_349_ vdd vss _146_ _023_ _349_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _007_ net30 net60 vss net77 vdd _418_/VPW vdd _418_/a_2665_112# _418_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output21_I vss net21 vdd ANTENNA_output21_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_203_ vdd vss net21 net11 _203_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_155 vdd vss FILLER_0_19_155/VPW vdd FILLER_0_19_155/a_36_472# FILLER_0_19_155/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_111 vdd vss FILLER_0_19_111/VPW vdd FILLER_0_19_111/a_36_472# FILLER_0_19_111/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_128 vdd vss FILLER_0_22_128/VPW vdd FILLER_0_22_128/a_3260_375# FILLER_0_22_128/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_180 vdd vss FILLER_0_15_180/VPW vdd FILLER_0_15_180/a_36_472# FILLER_0_15_180/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_150 vdd vss FILLER_0_21_150/VPW vdd FILLER_0_21_150/a_36_472# FILLER_0_21_150/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_47 vdd vss FILLER_0_6_47/VPW vdd FILLER_0_6_47/a_3260_375# FILLER_0_6_47/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_451_ vss net70 vdd _040_ cal_count\[1\] net53 _451_/VPW vdd _451_/a_36_151# vss
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_28 vdd vss FILLER_0_12_28/VPW vdd FILLER_0_12_28/a_36_472# FILLER_0_12_28/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ vdd vss _035_ _160_ _167_ _382_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_209 vdd vss FILLER_0_18_209/VPW vdd FILLER_0_18_209/a_36_472# FILLER_0_18_209/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vss FILLER_0_5_136/VPW vdd FILLER_0_5_136/a_36_472# FILLER_0_5_136/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_296_ vdd vss _009_ _104_ _107_ _296_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_434_ _023_ mask\[5\] net63 vss net80 vdd _434_/VPW vdd _434_/a_2665_112# _434_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_365_ _153_ _154_ _156_ vdd vss _029_ _155_ _365_/VPW vdd _365_/a_36_68# vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__280__A1 vss _095_ vdd ANTENNA__280__A1/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__240__I vss net41 vdd ANTENNA__240__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _144_ mask\[6\] vdd vss _146_ mask\[5\] _141_ _348_/VPW vdd _348_/a_49_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_417_ _006_ net29 net62 vss net79 vdd _417_/VPW vdd _417_/a_2665_112# _417_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_279_ vdd vss _096_ _090_ state\[1\] _279_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_231 vdd vss FILLER_0_6_231/VPW vdd FILLER_0_6_231/a_36_472# FILLER_0_6_231/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_202_ net21 vss vdd _047_ _202_/VPW vdd _202_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output14_I vss net14 vdd ANTENNA_output14_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_91 vdd vss FILLER_0_4_91/VPW vdd FILLER_0_4_91/a_36_472# FILLER_0_4_91/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_94 vdd vss FILLER_0_10_94/VPW vdd FILLER_0_10_94/a_36_472# FILLER_0_10_94/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vss FILLER_0_3_212/VPW vdd FILLER_0_3_212/a_36_472# FILLER_0_3_212/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_134 vdd vss FILLER_0_19_134/VPW vdd FILLER_0_19_134/a_36_472# FILLER_0_19_134/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_115 vdd vss FILLER_0_16_115/VPW vdd FILLER_0_16_115/a_36_472# FILLER_0_16_115/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vss FILLER_0_22_107/VPW vdd FILLER_0_22_107/a_36_472# FILLER_0_22_107/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_60 vdd vss FILLER_0_21_60/VPW vdd FILLER_0_21_60/a_36_472# FILLER_0_21_60/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vss FILLER_0_6_37/VPW vdd FILLER_0_6_37/a_36_472# FILLER_0_6_37/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_156 vdd vss FILLER_0_8_156/VPW vdd FILLER_0_8_156/a_36_472# FILLER_0_8_156/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I vss rstn vdd ANTENNA_input5_I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__243__I vss net47 vdd ANTENNA__243__I/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_450_ vss net67 vdd _039_ cal_count\[0\] net51 _450_/VPW vdd _450_/a_36_151# vss
+ gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xoutput40 trim[2] net40 vdd vss output40/VPW vdd output40/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_381_ trim_val\[2\] vdd vss _167_ trim_mask\[2\] _164_ _381_/VPW vdd _381_/a_36_472#
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_148 vdd vss FILLER_0_5_148/VPW vdd FILLER_0_5_148/a_36_472# FILLER_0_5_148/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_433_ _022_ mask\[4\] net54 vss net71 vdd _433_/VPW vdd _433_/a_2665_112# _433_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_295_ net32 vdd vss _107_ mask\[5\] _105_ _295_/VPW vdd _295_/a_36_472# vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_364_ vdd vss trim_mask\[2\] _156_ _364_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_235 vdd vss FILLER_0_14_235/VPW vdd FILLER_0_14_235/a_36_472# FILLER_0_14_235/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vss FILLER_0_13_72/VPW vdd FILLER_0_13_72/a_36_472# FILLER_0_13_72/a_572_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_347_ vdd vss _145_ _022_ _347_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_278_ _095_ vss vdd net3 _278_/VPW vdd _278_/a_36_160# vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_290 vdd vss FILLER_0_13_290/VPW vdd FILLER_0_13_290/a_36_472# FILLER_0_13_290/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ _005_ net28 net62 vss net79 vdd _416_/VPW vdd _416_/a_2665_112# _416_/a_36_151#
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_201_ vdd vss _047_ mask\[4\] net31 _201_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__448__RN vss net59 vdd ANTENNA__448__RN/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 result[3] net30 vdd vss output30/VPW vdd output30/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_196 vdd vss FILLER_0_12_196/VPW vdd FILLER_0_12_196/a_36_472# FILLER_0_12_196/a_124_375#
+ vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 clkc net6 vdd vss output6/VPW vdd output6/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 trim[3] net41 vdd vss output41/VPW vdd output41/a_224_472# vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_380_ vdd vss _034_ _160_ _166_ _380_/VPW vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
C0 net57 _163_ 0.759175f
C1 FILLER_0_17_282/a_36_472# vdd 0.107351f
C2 net4 net59 0.102012f
C3 trimb[1] vdd 0.225206f
C4 _448_/a_36_151# vdd 0.133302f
C5 _010_ vdd 0.121474f
C6 net35 _050_ 0.28822f
C7 FILLER_0_23_282/a_36_472# vdd 0.106034f
C8 _074_ net21 0.186175f
C9 FILLER_0_13_142/a_36_472# vdd 0.104785f
C10 net61 net62 0.874859f
C11 net52 trim_mask\[3\] 0.666362f
C12 net39 _033_ 0.607942f
C13 result[9] vdd 0.597071f
C14 net15 net50 0.177988f
C15 _031_ _157_ 0.104339f
C16 FILLER_0_21_125/a_36_472# _140_ 0.101284f
C17 _018_ net22 0.141743f
C18 net35 vss 0.434438f
C19 _072_ net22 0.147672f
C20 _178_ cal_count\[1\] 0.470244f
C21 _080_ vdd 0.123811f
C22 _070_ _172_ 0.237178f
C23 _127_ vss 0.343764f
C24 FILLER_0_14_107/a_36_472# vdd 0.114495f
C25 _056_ _055_ 0.155993f
C26 _072_ vdd 0.715894f
C27 _058_ _059_ 0.990213f
C28 _239_/a_36_160# _447_/a_36_151# 0.137659f
C29 _072_ _116_ 0.283323f
C30 _068_ _055_ 0.443477f
C31 _053_ net50 0.711279f
C32 _073_ _080_ 0.455535f
C33 _072_ _118_ 0.120452f
C34 mask\[7\] _108_ 0.785154f
C35 result[5] _103_ 0.425479f
C36 _106_ mask\[3\] 0.249479f
C37 net39 _444_/a_36_151# 0.14155f
C38 _115_ _068_ 0.889978f
C39 fanout76/a_36_160# vdd 0.108854f
C40 net20 ctlp[2] 0.254928f
C41 _056_ state\[1\] 0.219625f
C42 _053_ cal_itt\[3\] 0.471909f
C43 net61 net18 0.71051f
C44 _184_ vdd 0.202732f
C45 net31 _103_ 0.227588f
C46 trim_mask\[0\] net14 0.499565f
C47 _164_ _167_ 0.311625f
C48 _055_ _113_ 0.153988f
C49 _027_ vdd 0.146607f
C50 net63 _091_ 0.767908f
C51 _126_ _113_ 0.547055f
C52 _105_ output19/a_224_472# 0.107668f
C53 FILLER_0_2_177/a_36_472# vdd 0.110255f
C54 _069_ vss 0.323941f
C55 _095_ vdd 1.051346f
C56 net31 mask\[4\] 0.499009f
C57 _036_ vdd 0.364747f
C58 net35 net25 0.129685f
C59 vss rstn 0.149553f
C60 vdd net14 2.23064f
C61 _164_ vdd 0.711488f
C62 FILLER_0_19_125/a_36_472# _144_ 0.153815f
C63 net28 vss 0.185012f
C64 net15 vss 1.330044f
C65 _114_ _176_ 0.147182f
C66 net29 _006_ 0.135646f
C67 state\[1\] _113_ 0.107642f
C68 mask\[8\] _148_ 0.356546f
C69 net81 vss 0.766885f
C70 net15 mask\[9\] 0.128816f
C71 _178_ cal_count\[2\] 0.119443f
C72 _119_ _061_ 0.132725f
C73 net54 net14 0.121719f
C74 net38 vdd 0.906502f
C75 ctln[0] trim[3] 0.216084f
C76 _065_ net68 0.194392f
C77 _104_ vdd 0.662413f
C78 mask\[5\] net33 0.251971f
C79 _093_ _131_ 0.254316f
C80 _077_ _072_ 0.178678f
C81 _178_ _043_ 0.130207f
C82 _140_ vss 0.53195f
C83 _144_ vdd 0.40911f
C84 _171_ _172_ 0.104216f
C85 _153_ vdd 0.672318f
C86 net20 mask\[0\] 0.103301f
C87 _105_ _109_ 0.107328f
C88 _053_ vss 0.85895f
C89 net65 net18 0.879399f
C90 _053_ trim_mask\[1\] 0.110786f
C91 FILLER_0_5_72/a_36_472# vdd 0.107678f
C92 trimb[3] ctlp[0] 0.384753f
C93 valid vss 0.308766f
C94 trim_mask\[4\] FILLER_0_2_165/a_36_472# 0.265591f
C95 _057_ cal_count\[3\] 0.416063f
C96 ctlp[3] result[8] 0.278543f
C97 _412_/a_36_151# output48/a_224_472# 0.229574f
C98 _187_ _120_ 0.144679f
C99 _098_ net22 0.157058f
C100 _185_ vdd 0.325358f
C101 FILLER_0_22_86/a_36_472# _098_ 0.182093f
C102 ctlp[6] _050_ 0.100418f
C103 state\[0\] vss 0.126943f
C104 _151_ _163_ 0.501188f
C105 _133_ _152_ 0.124374f
C106 _074_ _084_ 0.110937f
C107 net80 _098_ 1.289178f
C108 _425_/a_36_151# _014_ 0.12681f
C109 ctlp[6] vss 0.115894f
C110 net34 output19/a_224_472# 0.122464f
C111 _119_ vss 0.22921f
C112 _086_ vdd 1.212255f
C113 _098_ vdd 2.272938f
C114 _069_ net23 0.418375f
C115 _345_/a_36_160# FILLER_0_19_111/a_572_375# 0.132282f
C116 FILLER_0_8_2/a_36_472# vdd 0.104141f
C117 _414_/a_36_151# vdd 0.166006f
C118 _053_ _155_ 0.122798f
C119 _095_ net47 0.508892f
C120 _086_ _116_ 1.316798f
C121 result[6] vdd 0.513079f
C122 _088_ net22 0.17798f
C123 net79 net4 0.386068f
C124 _070_ _060_ 0.822179f
C125 _086_ _118_ 0.166544f
C126 _070_ vdd 1.546772f
C127 net82 net22 1.960347f
C128 net47 _164_ 0.118311f
C129 _132_ _144_ 0.185339f
C130 _116_ _070_ 0.166494f
C131 net57 vdd 1.260693f
C132 _340_/a_36_160# FILLER_0_20_169/a_36_472# 0.195478f
C133 net9 cal_itt\[0\] 0.110446f
C134 net55 vdd 1.248648f
C135 ctln[2] vdd 0.245598f
C136 net54 _098_ 0.116416f
C137 _088_ vdd 0.140259f
C138 _079_ vss 0.124667f
C139 _070_ _118_ 0.302298f
C140 net17 vdd 2.139315f
C141 trim_val\[1\] vdd 0.173304f
C142 output21/a_224_472# result[8] 0.149245f
C143 FILLER_0_10_107/a_36_472# vdd 0.117291f
C144 _092_ vss 0.346097f
C145 _448_/a_36_151# net12 0.133216f
C146 _082_ vdd 0.191411f
C147 net82 vdd 1.014512f
C148 _137_ vss 0.343959f
C149 net38 net47 0.352245f
C150 cal_count\[3\] _120_ 4.687877f
C151 cal_count\[3\] _038_ 0.682941f
C152 _111_ vdd 0.3227f
C153 net52 trim_val\[4\] 0.21532f
C154 FILLER_0_16_107/a_36_472# vdd 0.110244f
C155 output36/a_224_472# net19 0.106928f
C156 net47 _153_ 0.755476f
C157 _015_ net27 0.103416f
C158 net1 net59 0.920133f
C159 ctlp[2] vdd 0.617599f
C160 _081_ _163_ 0.427672f
C161 FILLER_0_4_107/a_36_472# vdd 0.119007f
C162 _185_ net47 0.185634f
C163 _131_ _183_ 0.227229f
C164 _154_ _160_ 0.395185f
C165 net32 vss 0.824307f
C166 FILLER_0_10_247/a_36_472# vdd 0.111658f
C167 result[6] net77 0.111093f
C168 calibrate vdd 0.857987f
C169 net20 _076_ 0.228128f
C170 mask\[7\] net22 0.275179f
C171 _333_/a_36_160# vdd 0.107883f
C172 _257_/a_36_472# cal_itt\[3\] 0.136487f
C173 net16 _181_ 0.48682f
C174 _128_ vdd 0.217501f
C175 trim_mask\[2\] vdd 0.376424f
C176 net70 _095_ 0.222423f
C177 _127_ _176_ 0.319517f
C178 net82 net2 0.451147f
C179 _061_ _055_ 0.853642f
C180 net15 net36 0.265646f
C181 _128_ _118_ 0.58787f
C182 mask\[7\] vdd 1.098711f
C183 net70 net14 0.106631f
C184 net76 net59 3.439686f
C185 net57 trim_mask\[4\] 0.259381f
C186 _072_ _085_ 0.408915f
C187 net5 vss 0.326032f
C188 net57 net47 0.279638f
C189 net20 _093_ 0.398457f
C190 net20 net65 0.335083f
C191 FILLER_0_16_241/a_36_472# _099_ 0.158391f
C192 _032_ net69 0.347645f
C193 net74 _070_ 0.394108f
C194 net44 vss 0.477283f
C195 mask\[1\] vdd 0.741266f
C196 FILLER_0_15_72/a_572_375# cal_count\[1\] 0.135344f
C197 _328_/a_36_113# vdd 0.136098f
C198 _016_ net53 0.180698f
C199 net17 net47 2.009509f
C200 trim_val\[1\] net47 0.34878f
C201 _077_ _070_ 0.29321f
C202 net75 net76 0.106326f
C203 net57 net74 2.360287f
C204 _323_/a_36_113# _223_/a_36_160# 0.238626f
C205 net82 trim_mask\[4\] 0.21475f
C206 mask\[5\] _140_ 0.103728f
C207 trimb[0] trimb[3] 0.549457f
C208 result[6] ctlp[1] 0.677825f
C209 net54 mask\[7\] 0.262465f
C210 net23 _049_ 0.215528f
C211 _214_/a_36_160# _051_ 0.207388f
C212 _104_ output34/a_224_472# 0.112239f
C213 cal_count\[3\] _043_ 0.721078f
C214 net60 net18 0.949607f
C215 mask\[0\] vdd 0.181371f
C216 net20 _108_ 0.125627f
C217 net17 net43 0.144179f
C218 net3 vdd 0.118499f
C219 net46 vss 0.110452f
C220 net16 vdd 2.255325f
C221 _099_ vdd 0.326559f
C222 _055_ vss 0.365503f
C223 _085_ _071_ 0.127349f
C224 net55 _177_ 0.327874f
C225 net81 net21 0.185411f
C226 _126_ vss 0.399848f
C227 FILLER_0_21_142/a_36_472# vdd 0.111749f
C228 FILLER_0_1_212/a_36_472# vdd 0.10765f
C229 output42/a_224_472# output6/a_224_472# 0.292612f
C230 _069_ _176_ 0.766885f
C231 vdd net62 1.53102f
C232 net52 net69 0.372114f
C233 _115_ vss 0.372063f
C234 _414_/a_448_472# cal_itt\[3\] 0.109704f
C235 cal_itt\[1\] _082_ 0.921465f
C236 net29 net19 0.305661f
C237 net82 cal_itt\[1\] 0.396149f
C238 trim_mask\[3\] vss 0.156544f
C239 result[1] vss 0.311464f
C240 ctln[8] vss 0.351742f
C241 _091_ _072_ 0.162027f
C242 _129_ _068_ 0.104827f
C243 _142_ vss 0.121933f
C244 state\[1\] vss 0.294171f
C245 ctlp[3] _107_ 0.132316f
C246 _178_ _184_ 0.436202f
C247 _128_ net74 0.121254f
C248 result[9] net30 0.231442f
C249 trim[0] vdd 0.125774f
C250 _151_ vdd 0.157764f
C251 fanout58/a_36_160# vdd 0.101571f
C252 _056_ _068_ 0.127175f
C253 ctlp[5] vdd 0.293399f
C254 net61 vdd 0.46584f
C255 _178_ _095_ 0.839141f
C256 cal_itt\[2\] net4 0.333682f
C257 net65 net8 0.203388f
C258 _440_/a_36_151# vdd 0.117768f
C259 _078_ net59 0.168928f
C260 _161_ _113_ 0.201931f
C261 ctln[4] vdd 0.210384f
C262 net55 _040_ 0.107198f
C263 net68 net49 0.607379f
C264 _131_ vdd 1.344823f
C265 ctlp[8] vdd 0.115254f
C266 output33/a_224_472# net19 0.12997f
C267 _261_/a_36_160# FILLER_0_5_148/a_36_472# 0.195478f
C268 vdd net40 1.984115f
C269 net18 vdd 1.496006f
C270 net15 _030_ 0.355335f
C271 _196_/a_36_160# vdd 0.106963f
C272 net56 vdd 0.277166f
C273 net32 mask\[5\] 0.304094f
C274 net77 net62 0.122747f
C275 net38 _178_ 0.123812f
C276 _086_ _085_ 0.374127f
C277 _170_ vdd 0.18848f
C278 _015_ vdd 0.27747f
C279 _277_/a_36_160# vdd 0.115507f
C280 _133_ vss 0.18326f
C281 _076_ vdd 0.806117f
C282 _081_ net22 0.103561f
C283 _114_ _057_ 0.30288f
C284 mask\[3\] _099_ 0.10534f
C285 net65 net22 0.374917f
C286 en_co_clk vdd 0.245319f
C287 fanout69/a_36_113# _371_/a_36_113# 0.259508f
C288 en fanout59/a_36_160# 0.242369f
C289 net39 net40 0.279259f
C290 net57 _085_ 0.211414f
C291 net80 _093_ 0.818824f
C292 _178_ _185_ 0.979797f
C293 _081_ vdd 0.729534f
C294 _219_/a_36_160# trim_mask\[0\] 0.395762f
C295 _093_ vdd 1.439861f
C296 _164_ _160_ 1.863027f
C297 net65 vdd 1.430654f
C298 net61 net77 0.986569f
C299 _132_ _131_ 0.444097f
C300 _074_ net1 0.128466f
C301 _028_ net15 0.223301f
C302 net10 ctln[4] 0.1323f
C303 en net5 0.892091f
C304 _090_ _060_ 0.396493f
C305 _104_ _105_ 0.931514f
C306 _090_ vdd 0.751973f
C307 _116_ _090_ 0.122467f
C308 net50 trim_val\[3\] 0.111824f
C309 _073_ net65 0.775972f
C310 _029_ vdd 0.223076f
C311 net18 net77 0.378783f
C312 result[8] mask\[6\] 0.111221f
C313 _108_ vdd 0.298249f
C314 _103_ _094_ 0.280781f
C315 net79 _043_ 0.393702f
C316 _153_ _160_ 0.304792f
C317 net47 net40 0.635497f
C318 net50 trim_val\[0\] 0.390586f
C319 _141_ _140_ 0.131685f
C320 net31 _094_ 0.203395f
C321 result[5] vss 0.307366f
C322 _091_ _098_ 1.501073f
C323 _178_ net17 0.115251f
C324 _131_ net74 0.227843f
C325 _053_ _028_ 0.891578f
C326 _122_ vss 0.750387f
C327 _114_ _120_ 0.334426f
C328 net61 ctlp[1] 2.770871f
C329 net41 _446_/a_36_151# 0.143017f
C330 net64 vss 0.636644f
C331 _163_ vdd 0.418075f
C332 net26 _052_ 0.100927f
C333 _091_ _070_ 0.162632f
C334 _022_ _145_ 0.199016f
C335 _132_ _093_ 0.105039f
C336 _117_ _060_ 0.149558f
C337 net52 net50 0.702793f
C338 net31 vss 0.562041f
C339 _114_ state\[2\] 0.528838f
C340 net27 vdd 0.88294f
C341 calibrate _062_ 2.032477f
C342 FILLER_0_11_142/a_36_472# vdd 0.110248f
C343 trim_mask\[4\] _081_ 0.111668f
C344 mask\[4\] vss 0.426009f
C345 _077_ _076_ 1.895143f
C346 _081_ net47 1.302193f
C347 _174_ vss 0.188373f
C348 FILLER_0_18_2/a_36_472# vdd 0.104532f
C349 cal_count\[3\] _071_ 0.214649f
C350 _093_ _012_ 0.141641f
C351 net20 vdd 2.14128f
C352 mask\[2\] vss 0.536426f
C353 net34 _147_ 0.144404f
C354 _104_ net34 0.293336f
C355 output39/a_224_472# net39 0.129913f
C356 ctlp[2] _011_ 0.101324f
C357 output33/a_224_472# net33 0.151281f
C358 _339_/a_36_160# FILLER_0_19_171/a_36_472# 0.195478f
C359 _075_ net22 0.180274f
C360 cal_itt\[3\] _161_ 0.20195f
C361 trim_val\[4\] vss 0.192567f
C362 trimb[3] vss 0.161605f
C363 _183_ vdd 0.109252f
C364 _141_ _137_ 0.40175f
C365 ctln[9] vdd 0.221231f
C366 net27 result[0] 0.106157f
C367 mask\[3\] _093_ 2.443356f
C368 _029_ net47 2.210804f
C369 net72 cal_count\[1\] 0.13509f
C370 net20 _073_ 0.437482f
C371 _105_ ctlp[2] 0.223601f
C372 state\[1\] net21 0.210202f
C373 net70 _131_ 0.57653f
C374 net72 FILLER_0_17_38/a_36_472# 0.123542f
C375 trim_val\[3\] vss 0.249446f
C376 _075_ vdd 0.190898f
C377 _066_ _169_ 0.222791f
C378 _122_ net23 0.276617f
C379 net50 net69 0.634381f
C380 net52 _031_ 0.633473f
C381 output34/a_224_472# net18 0.126175f
C382 ctln[1] cal 0.123834f
C383 state\[0\] net4 0.13193f
C384 _144_ _146_ 0.333799f
C385 net47 _163_ 0.64626f
C386 _115_ _176_ 1.300336f
C387 trim_val\[0\] vss 0.11063f
C388 _131_ _040_ 0.211618f
C389 vdd _039_ 0.219985f
C390 net80 _139_ 0.178583f
C391 _178_ net3 0.257606f
C392 _136_ _137_ 0.417639f
C393 net41 _095_ 0.641184f
C394 output19/a_224_472# net33 0.126671f
C395 _056_ _061_ 0.445098f
C396 net16 _178_ 0.30147f
C397 _105_ mask\[7\] 0.486236f
C398 trim_mask\[2\] _160_ 0.367302f
C399 net4 _083_ 0.135165f
C400 net52 vss 1.608047f
C401 mask\[4\] net23 0.111873f
C402 _061_ _068_ 1.857322f
C403 net60 vdd 0.575502f
C404 FILLER_0_4_177/a_36_472# vdd 0.114788f
C405 _119_ _058_ 0.692466f
C406 mask\[2\] net23 0.431197f
C407 net28 net29 0.178557f
C408 _086_ cal_count\[3\] 0.259095f
C409 _161_ vss 0.134214f
C410 _129_ vss 0.141494f
C411 output38/a_224_472# _445_/a_36_151# 0.199812f
C412 _088_ net59 0.270902f
C413 vdd trim[2] 0.166648f
C414 net8 vdd 0.593788f
C415 net49 _164_ 0.428468f
C416 ctln[3] ctln[1] 0.926618f
C417 vdd FILLER_0_3_212/a_36_472# 0.110132f
C418 net69 _031_ 0.450281f
C419 net82 net59 0.102279f
C420 _181_ vdd 0.209604f
C421 net34 ctlp[2] 0.953441f
C422 net63 net35 0.126544f
C423 _024_ _435_/a_36_151# 0.10993f
C424 _127_ _120_ 0.198577f
C425 _056_ vss 0.193804f
C426 mask\[8\] net35 2.631701f
C427 net75 _082_ 0.417366f
C428 _131_ _062_ 0.120189f
C429 _037_ vdd 0.158731f
C430 net75 net82 0.214597f
C431 result[7] result[9] 1.21288f
C432 net81 net37 0.18149f
C433 net38 net49 0.117427f
C434 net16 _160_ 0.354736f
C435 _068_ vss 0.547532f
C436 _073_ net8 0.206839f
C437 mask\[6\] vss 0.348967f
C438 net69 vss 0.34555f
C439 _105_ output18/a_224_472# 0.105478f
C440 ctlp[4] result[8] 0.151286f
C441 _100_ vdd 0.212037f
C442 _152_ vss 0.140215f
C443 trim_mask\[0\] vdd 0.154098f
C444 _010_ net19 0.408364f
C445 mask\[5\] mask\[4\] 0.176881f
C446 _060_ net22 0.533421f
C447 net23 _208_/a_36_160# 0.112626f
C448 net22 vdd 1.920713f
C449 _076_ _062_ 0.978627f
C450 output12/a_224_472# vdd 0.106635f
C451 net34 mask\[7\] 0.901671f
C452 net62 net30 0.339141f
C453 _072_ _074_ 2.017168f
C454 FILLER_0_10_78/a_36_472# cal_count\[3\] 0.266339f
C455 _013_ vss 0.163674f
C456 _077_ _039_ 0.104126f
C457 _116_ net22 0.122052f
C458 ctln[1] vss 0.27233f
C459 net80 vdd 1.045288f
C460 net4 net5 0.104296f
C461 result[9] net19 0.540761f
C462 _142_ _141_ 0.200324f
C463 _060_ vdd 0.349556f
C464 _113_ vss 0.147905f
C465 _165_ _164_ 0.351097f
C466 net75 calibrate 0.101912f
C467 FILLER_0_17_72/a_36_472# vdd 0.111688f
C468 net36 mask\[2\] 0.871463f
C469 calibrate _059_ 0.506928f
C470 _187_ net16 0.161791f
C471 _116_ vdd 0.399137f
C472 net41 net17 0.911377f
C473 FILLER_0_16_73/a_572_375# _175_ 0.138524f
C474 net71 vss 0.335256f
C475 _005_ mask\[1\] 0.246517f
C476 _118_ vdd 0.292155f
C477 result[5] _008_ 0.165753f
C478 _063_ _033_ 0.250192f
C479 mask\[9\] net71 0.344312f
C480 _123_ vdd 0.214703f
C481 net54 vdd 0.877573f
C482 _073_ vdd 0.258125f
C483 _064_ vss 0.228443f
C484 net40 _160_ 0.152292f
C485 net4 _055_ 0.216844f
C486 _079_ net37 0.408392f
C487 net39 vdd 0.2282f
C488 _068_ net23 0.432092f
C489 result[4] vss 0.306116f
C490 _008_ net31 0.292444f
C491 net26 net72 0.868238f
C492 result[8] vss 0.235206f
C493 result[0] vdd 0.193436f
C494 FILLER_0_5_212/a_36_472# vdd 0.107657f
C495 net34 output18/a_224_472# 0.17524f
C496 _132_ vdd 0.960634f
C497 FILLER_0_18_107/a_36_472# vdd 0.116746f
C498 net2 vdd 0.434557f
C499 net10 vdd 0.227004f
C500 _045_ vdd 0.246567f
C501 _091_ _090_ 0.117348f
C502 net77 vdd 0.526632f
C503 _104_ result[7] 0.475003f
C504 FILLER_0_8_247/a_36_472# vdd 0.112197f
C505 trim_mask\[4\] vdd 0.20602f
C506 net47 vdd 2.422992f
C507 _012_ vdd 0.261844f
C508 _006_ net62 0.136418f
C509 FILLER_0_15_212/a_36_472# vdd 0.105575f
C510 _064_ net66 0.304028f
C511 net74 vdd 1.451847f
C512 _182_ cal_count\[1\] 0.166348f
C513 result[9] _009_ 0.19745f
C514 net58 net81 0.375649f
C515 net15 net51 0.191328f
C516 _077_ vdd 1.61568f
C517 _154_ _157_ 0.447829f
C518 net45 net17 0.192181f
C519 _105_ _108_ 0.548284f
C520 output22/a_224_472# _435_/a_36_151# 0.12978f
C521 net43 vdd 0.210686f
C522 mask\[3\] vdd 0.340612f
C523 _059_ FILLER_0_8_156/a_36_472# 0.18373f
C524 _104_ net19 0.159483f
C525 ctlp[1] vdd 0.942436f
C526 cal vss 0.424638f
C527 ctln[4] net59 0.10527f
C528 net81 net76 0.236554f
C529 mask\[5\] mask\[6\] 0.140269f
C530 net80 _019_ 0.265857f
C531 _065_ ctln[9] 0.123393f
C532 net41 net16 2.918931f
C533 net39 net47 0.13057f
C534 result[6] result[7] 0.119475f
C535 net15 net68 0.205016f
C536 _086_ _074_ 0.186795f
C537 _114_ net14 0.127764f
C538 _177_ vdd 0.111636f
C539 net18 net59 0.695067f
C540 net58 valid 0.149817f
C541 _163_ _160_ 0.120564f
C542 net50 _054_ 0.131493f
C543 cal_itt\[1\] vdd 0.410279f
C544 _431_/a_36_151# vdd 0.145005f
C545 net15 net67 0.109181f
C546 net50 vss 1.178736f
C547 _074_ _070_ 0.102481f
C548 net1 _083_ 0.30074f
C549 net50 trim_mask\[1\] 0.502622f
C550 _102_ _099_ 0.151018f
C551 net24 net14 0.172253f
C552 _119_ _125_ 0.11554f
C553 valid net76 0.285892f
C554 _056_ net21 0.484506f
C555 _063_ _164_ 0.326812f
C556 _053_ net68 0.239882f
C557 _074_ net82 0.123449f
C558 cal_itt\[3\] vss 0.15522f
C559 net38 _445_/a_36_151# 0.112205f
C560 result[6] net19 0.834308f
C561 _101_ _094_ 0.304499f
C562 ctlp[4] vss 0.102044f
C563 _089_ _079_ 0.126206f
C564 net32 output19/a_224_472# 0.101682f
C565 mask\[4\] _141_ 0.948091f
C566 trim_mask\[4\] net47 0.264421f
C567 _081_ net59 0.185504f
C568 net70 vdd 0.858299f
C569 _053_ net67 0.672744f
C570 _076_ _059_ 1.03702f
C571 net21 mask\[6\] 0.634881f
C572 net36 net71 0.148833f
C573 net65 net59 0.790496f
C574 net53 _427_/a_36_151# 0.13192f
C575 net74 trim_mask\[4\] 0.548293f
C576 _057_ _055_ 0.290639f
C577 ctln[3] vss 0.133697f
C578 net34 _108_ 0.297364f
C579 ctlp[1] net77 0.716304f
C580 net75 net65 0.135447f
C581 net82 net19 1.14585f
C582 FILLER_0_19_142/a_36_472# vdd 0.107105f
C583 _432_/a_36_151# vdd 0.173104f
C584 net2 cal_itt\[1\] 0.284695f
C585 _086_ _114_ 1.371271f
C586 _415_/a_36_151# vdd 0.115639f
C587 net41 net40 2.687418f
C588 _079_ net76 2.404004f
C589 net74 _159_ 0.129233f
C590 _031_ vss 0.18315f
C591 _053_ _154_ 0.41707f
C592 net63 output35/a_224_472# 0.148302f
C593 _035_ trim[0] 0.171633f
C594 _114_ _070_ 0.507391f
C595 _094_ vss 0.24519f
C596 net72 _095_ 0.136566f
C597 cal_count\[3\] _090_ 0.243462f
C598 _057_ state\[1\] 0.284428f
C599 _114_ net57 0.22998f
C600 _418_/a_36_151# vdd 0.155643f
C601 net7 vdd 0.321735f
C602 _104_ _009_ 0.284256f
C603 net62 result[3] 0.451989f
C604 _178_ _181_ 0.188669f
C605 net78 vss 0.167812f
C606 ctlp[7] _050_ 0.153673f
C607 _050_ vss 0.26237f
C608 _136_ mask\[2\] 1.822289f
C609 _020_ vdd 0.194776f
C610 _132_ net70 0.534228f
C611 _054_ vss 0.176655f
C612 net1 net5 0.266194f
C613 mask\[0\] net79 0.243338f
C614 trim_mask\[1\] vss 0.449335f
C615 _085_ vdd 0.227153f
C616 vss _107_ 0.186994f
C617 _437_/a_36_151# vdd 0.115376f
C618 mask\[4\] _145_ 0.340415f
C619 _028_ net52 0.150861f
C620 mask\[9\] vss 0.649041f
C621 _053_ _078_ 0.137388f
C622 result[8] net21 0.166555f
C623 net58 net5 0.387314f
C624 net79 net62 1.615103f
C625 net48 _070_ 0.264809f
C626 _062_ vdd 0.393862f
C627 net69 _030_ 0.49547f
C628 _346_/a_49_472# _141_ 0.104653f
C629 _065_ vdd 0.646511f
C630 _155_ vss 0.13648f
C631 _187_ _039_ 0.228074f
C632 _008_ result[4] 0.134001f
C633 net44 cal_count\[2\] 0.191151f
C634 _178_ vdd 0.440802f
C635 _072_ _069_ 0.265737f
C636 net18 result[3] 0.237732f
C637 _004_ vdd 0.448886f
C638 net66 vss 0.265973f
C639 _067_ vss 0.20904f
C640 state\[2\] state\[1\] 0.229832f
C641 cal en 0.482495f
C642 net61 net79 0.159f
C643 _091_ net80 0.23053f
C644 net44 clkc 0.184915f
C645 _007_ vdd 0.129966f
C646 _106_ _092_ 0.140596f
C647 _091_ vdd 1.011371f
C648 net72 net55 0.233515f
C649 _011_ vdd 0.182751f
C650 _167_ _160_ 0.157458f
C651 net39 trim[1] 0.115976f
C652 _428_/a_36_151# vdd 0.131612f
C653 result[6] net33 0.363421f
C654 net19 net62 0.352148f
C655 net25 vss 0.528437f
C656 net23 vss 1.922425f
C657 output14/a_224_472# _442_/a_36_151# 0.172111f
C658 ctlp[2] _009_ 0.220631f
C659 _087_ _079_ 0.251042f
C660 net79 net18 0.222939f
C661 FILLER_0_11_109/a_36_472# vdd 0.109453f
C662 _122_ net37 3.870625f
C663 net48 calibrate 0.482314f
C664 _114_ _171_ 0.203692f
C665 cal_itt\[2\] net82 0.663246f
C666 _105_ vdd 0.565719f
C667 net16 _186_ 0.225785f
C668 _126_ _043_ 0.128227f
C669 vdd _160_ 0.606139f
C670 output13/a_224_472# vss 0.108144f
C671 _074_ _162_ 0.112872f
C672 trim_mask\[1\] _166_ 0.124855f
C673 _030_ _156_ 0.153053f
C674 vdd net30 0.636147f
C675 net29 mask\[2\] 0.122202f
C676 net61 net19 0.132027f
C677 vss cal_count\[0\] 0.160743f
C678 output28/a_224_472# net62 0.206137f
C679 _417_/a_36_151# vdd 0.140703f
C680 _119_ _072_ 0.189217f
C681 state\[1\] _043_ 0.1587f
C682 _161_ _058_ 0.101968f
C683 _136_ _138_ 0.186242f
C684 cal_itt\[0\] vss 0.11965f
C685 cal_itt\[3\] net21 0.175781f
C686 _144_ _022_ 0.139742f
C687 FILLER_0_11_124/a_36_472# _135_ 0.110114f
C688 net75 net8 0.553872f
C689 net67 _439_/a_36_151# 0.136402f
C690 _037_ net59 0.799647f
C691 _187_ vdd 0.194575f
C692 mask\[5\] vss 0.528441f
C693 _056_ _058_ 0.988919f
C694 FILLER_0_6_177/a_36_472# vdd 0.109918f
C695 net36 vss 1.788802f
C696 _053_ net14 0.713784f
C697 output20/a_224_472# net61 0.177946f
C698 ctln[5] _037_ 0.19244f
C699 _017_ vdd 0.26981f
C700 net34 vdd 1.161282f
C701 _122_ _120_ 0.143427f
C702 net22 net59 0.195226f
C703 en vss 0.466499f
C704 mask\[9\] net36 1.116767f
C705 _067_ cal_count\[0\] 0.201595f
C706 _394_/a_56_524# _095_ 0.10007f
C707 _086_ _069_ 0.580351f
C708 trim_mask\[4\] _160_ 0.244284f
C709 net47 _160_ 0.2966f
C710 _005_ vdd 0.506158f
C711 net59 vdd 2.180407f
C712 _144_ _140_ 0.415736f
C713 net16 net72 0.367221f
C714 _069_ _070_ 0.257147f
C715 net74 _160_ 0.165289f
C716 _127_ _128_ 0.257374f
C717 net21 vss 1.123312f
C718 _105_ ctlp[1] 0.158795f
C719 net75 vdd 1.265616f
C720 net35 mask\[7\] 0.954332f
C721 _074_ _163_ 0.446493f
C722 _008_ _094_ 0.234346f
C723 _096_ _126_ 0.258912f
C724 cal_count\[3\] vdd 1.020669f
C725 _059_ vdd 0.161836f
C726 ctln[5] vdd 0.256793f
C727 _006_ vdd 0.632993f
C728 _116_ cal_count\[3\] 0.384121f
C729 net15 net55 1.200864f
C730 mask\[3\] net30 0.451388f
C731 _132_ _017_ 0.155924f
C732 net75 _123_ 0.173358f
C733 _140_ _098_ 0.647503f
C734 net63 mask\[2\] 0.553545f
C735 net75 _073_ 0.34505f
C736 _008_ vss 0.355468f
C737 net58 net64 0.590523f
C738 fanout71/a_36_113# _433_/a_36_151# 0.138322f
C739 _176_ vss 0.761803f
C740 ctln[6] net52 0.1064f
C741 net20 result[7] 0.134149f
C742 _057_ _161_ 1.09228f
C743 output18/a_224_472# net33 0.135766f
C744 _124_ vss 0.110847f
C745 _250_/a_36_68# state\[1\] 0.103037f
C746 _053_ _070_ 2.345795f
C747 net2 net59 0.334636f
C748 _149_ net71 0.827628f
C749 _119_ _086_ 0.419383f
C750 net41 vdd 1.983262f
C751 _132_ cal_count\[3\] 0.193553f
C752 net72 _131_ 0.186396f
C753 _057_ _056_ 0.167928f
C754 _144_ _049_ 0.100508f
C755 net48 _081_ 0.137029f
C756 net20 _000_ 0.159624f
C757 sample net18 0.103617f
C758 _119_ _070_ 1.949038f
C759 net20 net19 0.384932f
C760 _292_/a_36_160# _205_/a_36_160# 0.105676f
C761 _057_ _068_ 0.393271f
C762 FILLER_0_17_142/a_36_472# vdd 0.108843f
C763 net42 net6 0.166896f
C764 _119_ net57 0.30462f
C765 clk rstn 0.541051f
C766 net63 _434_/a_2665_112# 0.120476f
C767 net34 ctlp[1] 0.127025f
C768 _102_ vdd 0.211559f
C769 _030_ vss 0.117034f
C770 net49 vdd 0.872948f
C771 net60 net79 0.113281f
C772 _174_ _043_ 0.964645f
C773 net32 _104_ 0.342568f
C774 output39/a_224_472# _445_/a_36_151# 0.11862f
C775 _430_/a_36_151# vdd 0.112575f
C776 _072_ state\[1\] 0.267762f
C777 _035_ vdd 0.215473f
C778 net28 mask\[1\] 0.572459f
C779 _077_ cal_count\[3\] 0.176576f
C780 result[7] net60 0.778099f
C781 _057_ _113_ 0.339862f
C782 net81 mask\[1\] 2.509493f
C783 FILLER_0_14_50/a_36_472# _180_ 0.153222f
C784 sample net65 0.148853f
C785 _079_ _082_ 0.709481f
C786 cal_itt\[1\] net59 0.227495f
C787 cal_itt\[2\] net65 0.514538f
C788 _009_ _108_ 1.645945f
C789 _421_/a_36_151# _419_/a_36_151# 0.561555f
C790 net38 net44 0.523774f
C791 net39 net49 0.158007f
C792 _052_ vdd 0.264744f
C793 _025_ vdd 0.259346f
C794 _127_ _131_ 0.470047f
C795 vdd _034_ 0.424437f
C796 state\[0\] _128_ 0.228492f
C797 net75 cal_itt\[1\] 0.704169f
C798 _141_ vss 0.308762f
C799 _068_ _120_ 0.447243f
C800 _028_ vss 0.410396f
C801 net81 mask\[0\] 0.320022f
C802 vdd result[3] 0.181788f
C803 _028_ trim_mask\[1\] 0.148182f
C804 _126_ net14 0.238336f
C805 net41 net47 0.19549f
C806 state\[1\] _071_ 0.196063f
C807 net60 net19 0.102311f
C808 _165_ vdd 0.168803f
C809 net81 _099_ 0.140011f
C810 _078_ _122_ 0.185069f
C811 net63 mask\[6\] 0.146994f
C812 mask\[5\] net21 0.212814f
C813 net79 _100_ 0.170973f
C814 FILLER_0_24_274/a_36_472# vdd 0.107635f
C815 trim_mask\[3\] net14 0.142743f
C816 _453_/a_36_151# vdd 0.164654f
C817 _127_ _076_ 0.137964f
C818 FILLER_0_15_282/a_36_472# vdd 0.10628f
C819 net67 trim_val\[0\] 0.382079f
C820 net81 net62 0.245647f
C821 net49 net47 0.53353f
C822 _136_ vss 0.947188f
C823 net79 vdd 1.283563f
C824 _035_ net47 0.101683f
C825 mask\[3\] _102_ 0.142836f
C826 trimb[4] net44 0.127019f
C827 net53 vss 0.426484f
C828 _176_ net36 0.336675f
C829 result[7] vdd 0.500292f
C830 trim[4] vdd 0.198218f
C831 mask\[8\] net71 0.424276f
C832 mask\[7\] _049_ 0.234746f
C833 net55 _041_ 0.972122f
C834 _137_ mask\[1\] 0.782055f
C835 net4 vss 0.774455f
C836 _086_ _055_ 0.113385f
C837 net20 cal_itt\[2\] 0.715447f
C838 _074_ vdd 1.221102f
C839 _087_ FILLER_0_5_181/a_36_472# 0.154469f
C840 _174_ _180_ 0.102241f
C841 net10 _411_/a_36_151# 0.127193f
C842 vss _145_ 0.399701f
C843 FILLER_0_3_172/a_36_472# fanout57/a_36_113# 0.19419f
C844 _141_ net23 0.782974f
C845 _070_ _055_ 0.516713f
C846 _086_ _115_ 0.4112f
C847 _182_ _179_ 0.109377f
C848 _053_ _151_ 0.538643f
C849 net57 FILLER_0_16_154/a_1468_375# 0.217874f
C850 ctln[5] net12 0.41364f
C851 net81 net18 0.102876f
C852 _074_ _123_ 0.157299f
C853 net46 net17 0.791341f
C854 _058_ vss 0.19427f
C855 _000_ vdd 0.215988f
C856 _115_ _070_ 0.890903f
C857 net19 vdd 2.167778f
C858 _042_ vdd 0.261947f
C859 _085_ cal_count\[3\] 0.653405f
C860 net79 net77 0.431572f
C861 _420_/a_36_151# vdd 0.137919f
C862 trim_mask\[1\] FILLER_0_4_91/a_36_472# 0.26171f
C863 net57 state\[1\] 0.154183f
C864 _000_ _073_ 0.222349f
C865 _093_ net15 0.145303f
C866 net45 net43 0.131763f
C867 _069_ _090_ 1.067281f
C868 _059_ _062_ 0.161331f
C869 _053_ _076_ 0.108358f
C870 _114_ vdd 1.30767f
C871 net7 net41 0.243942f
C872 net29 _094_ 0.313846f
C873 net53 net23 0.501857f
C874 _026_ net71 0.406369f
C875 net15 _029_ 0.111797f
C876 mask\[5\] _141_ 0.241158f
C877 net80 _434_/a_448_472# 0.113898f
C878 _105_ net34 0.784678f
C879 _016_ vdd 0.114288f
C880 net48 _112_ 0.284235f
C881 _128_ _055_ 1.887595f
C882 _053_ _081_ 0.698311f
C883 FILLER_0_20_107/a_36_472# vdd 0.117841f
C884 net24 vdd 0.223761f
C885 _131_ _182_ 0.113302f
C886 FILLER_0_8_138/a_124_375# _120_ 0.12254f
C887 net29 vss 0.259409f
C888 trim_val\[2\] _036_ 0.279133f
C889 net44 net3 0.195171f
C890 _063_ vdd 0.201806f
C891 _115_ _128_ 0.263909f
C892 _077_ _074_ 0.148596f
C893 mask\[9\] FILLER_0_19_111/a_36_472# 0.285112f
C894 _070_ _133_ 0.436976f
C895 vss trim[3] 0.235724f
C896 net67 net42 0.101108f
C897 net37 vss 0.666835f
C898 cal net1 0.336092f
C899 _013_ net26 0.174966f
C900 net48 vdd 0.35704f
C901 _174_ _095_ 0.977766f
C902 ctlp[3] mask\[7\] 0.103955f
C903 output32/a_224_472# net60 0.191561f
C904 FILLER_0_3_2/a_36_472# vdd 0.106665f
C905 net81 net27 1.118985f
C906 _074_ cal_itt\[1\] 0.120296f
C907 _077_ _188_ 0.1656f
C908 _009_ vdd 0.693198f
C909 _136_ net36 1.151311f
C910 FILLER_0_9_282/a_36_472# vdd 0.106034f
C911 _053_ _163_ 0.763235f
C912 _070_ _121_ 0.285424f
C913 net31 _104_ 0.102776f
C914 _057_ vss 0.169369f
C915 net48 _123_ 0.153061f
C916 _079_ _081_ 1.441057f
C917 FILLER_0_15_142/a_36_472# vdd 0.106034f
C918 ctlp[9] vdd 0.17413f
C919 result[2] _044_ 0.393081f
C920 _006_ net30 0.284414f
C921 net53 net36 3.423337f
C922 _092_ _093_ 0.287983f
C923 _093_ _137_ 0.201779f
C924 ctln[6] vss 0.45431f
C925 comp vdd 0.108153f
C926 net72 vdd 1.425686f
C927 sample vdd 0.154389f
C928 _144_ mask\[4\] 0.268823f
C929 FILLER_0_18_37/a_36_472# vdd 0.136723f
C930 cal_itt\[2\] vdd 0.267121f
C931 _114_ net74 0.559239f
C932 _096_ _113_ 0.650985f
C933 net64 _098_ 0.281888f
C934 FILLER_0_5_54/a_36_472# trim_mask\[1\] 0.101342f
C935 FILLER_0_17_200/a_36_472# mask\[3\] 0.27914f
C936 vdd FILLER_0_22_107/a_36_472# 0.114332f
C937 en net4 0.125535f
C938 _070_ _122_ 0.153373f
C939 _024_ vss 0.132549f
C940 cal_count\[1\] vss 0.307993f
C941 _016_ net74 0.568682f
C942 _023_ vss 0.114191f
C943 net33 vdd 0.42212f
C944 _063_ net47 0.142088f
C945 trim_val\[0\] _164_ 0.133785f
C946 net1 _001_ 0.300335f
C947 cal_itt\[2\] _073_ 0.202415f
C948 _072_ _068_ 0.185471f
C949 net20 state\[0\] 0.396139f
C950 net50 net68 0.224698f
C951 _120_ vss 0.42505f
C952 _038_ vss 0.373776f
C953 net19 FILLER_0_14_263/a_36_472# 0.135429f
C954 _176_ _136_ 0.114837f
C955 net52 _164_ 0.313379f
C956 _053_ _075_ 0.634359f
C957 net63 vss 0.566021f
C958 FILLER_0_11_282/a_36_472# vdd 0.106843f
C959 net50 net67 0.518421f
C960 net49 _160_ 1.243817f
C961 net46 net40 0.254778f
C962 mask\[8\] vss 0.378558f
C963 net35 vdd 1.0365f
C964 _077_ net48 0.142015f
C965 _126_ _131_ 0.626666f
C966 net20 _083_ 0.230786f
C967 state\[2\] vss 0.185787f
C968 net57 _097_ 0.100409f
C969 _175_ vss 0.162988f
C970 _127_ vdd 0.155954f
C971 _115_ _131_ 0.410424f
C972 _035_ _160_ 0.120469f
C973 net21 net11 0.10869f
C974 net20 _079_ 0.177911f
C975 net1 vss 0.161208f
C976 net54 net35 0.114666f
C977 _127_ _118_ 0.141388f
C978 _157_ vdd 0.419501f
C979 net57 trim_val\[4\] 0.295336f
C980 _242_/a_36_160# FILLER_0_5_164/a_36_472# 0.193804f
C981 FILLER_0_2_165/a_124_375# net22 0.206491f
C982 _128_ net64 0.291788f
C983 result[4] result[9] 0.101112f
C984 result[8] result[9] 0.242998f
C985 ctln[7] vss 0.132613f
C986 _004_ net79 0.27387f
C987 _125_ vss 0.149512f
C988 net58 vss 0.589419f
C989 net82 trim_val\[4\] 0.511271f
C990 net29 net36 0.370099f
C991 trim_mask\[2\] trim_val\[2\] 0.21814f
C992 net9 vdd 0.190349f
C993 _038_ _067_ 0.503045f
C994 _308_/a_848_380# FILLER_0_9_105/a_36_472# 0.15783f
C995 _036_ net69 0.353233f
C996 _415_/a_36_151# output28/a_224_472# 0.229574f
C997 net51 vss 0.21065f
C998 _069_ net22 0.327999f
C999 cal_count\[2\] vss 0.361185f
C1000 net76 vss 0.436111f
C1001 _132_ _127_ 0.112364f
C1002 _120_ net23 0.147166f
C1003 _069_ _060_ 0.538161f
C1004 _043_ vss 1.362912f
C1005 net16 _408_/a_728_93# 0.107634f
C1006 _069_ vdd 0.985405f
C1007 net81 _100_ 0.24831f
C1008 _147_ mask\[6\] 0.103475f
C1009 _142_ _093_ 0.492191f
C1010 net68 vss 0.635359f
C1011 ctlp[1] net33 0.11288f
C1012 _150_ mask\[9\] 0.162185f
C1013 _069_ _116_ 0.390834f
C1014 mask\[0\] net64 0.45093f
C1015 vdd rstn 0.160093f
C1016 state\[2\] net23 0.331644f
C1017 net67 _054_ 0.391592f
C1018 _144_ mask\[6\] 0.230129f
C1019 net28 vdd 0.489756f
C1020 net15 vdd 2.073988f
C1021 net67 vss 0.435869f
C1022 net52 net82 0.108202f
C1023 net71 net14 0.147175f
C1024 _131_ _133_ 0.20118f
C1025 _004_ net19 0.112289f
C1026 net16 trim_val\[2\] 0.124462f
C1027 net81 vdd 1.658963f
C1028 _132_ _135_ 0.345161f
C1029 _055_ _117_ 0.242156f
C1030 result[2] vss 0.327009f
C1031 net80 _140_ 0.188514f
C1032 net73 vss 0.342554f
C1033 _140_ vdd 0.598538f
C1034 _098_ mask\[6\] 0.297837f
C1035 _154_ vss 0.200253f
C1036 _053_ vdd 1.467835f
C1037 net73 mask\[9\] 0.383862f
C1038 _133_ _076_ 0.11688f
C1039 _070_ _068_ 1.019801f
C1040 _057_ net21 0.143214f
C1041 _049_ FILLER_0_22_128/a_3260_375# 0.16381f
C1042 _067_ _043_ 0.189767f
C1043 net27 result[1] 0.187252f
C1044 valid vdd 0.148392f
C1045 net20 _055_ 0.203142f
C1046 _099_ mask\[2\] 0.776725f
C1047 net68 net66 0.81104f
C1048 mask\[2\] FILLER_0_16_154/a_36_472# 0.312123f
C1049 net14 _156_ 0.184287f
C1050 net32 net60 0.509175f
C1051 state\[0\] vdd 0.120171f
C1052 net54 _140_ 1.37516f
C1053 net26 vss 0.263774f
C1054 _070_ _152_ 0.114651f
C1055 mask\[5\] net63 0.112147f
C1056 net67 _067_ 0.151887f
C1057 net44 _039_ 0.15647f
C1058 mask\[7\] _208_/a_36_160# 0.105845f
C1059 ctlp[6] vdd 0.207209f
C1060 _119_ vdd 0.38257f
C1061 _155_ _154_ 0.18488f
C1062 net41 net49 0.392356f
C1063 net19 net30 0.311153f
C1064 _021_ vss 0.142648f
C1065 net81 net2 1.204674f
C1066 output31/a_224_472# net60 0.216716f
C1067 _106_ vss 0.180823f
C1068 result[5] net18 0.173673f
C1069 _013_ net55 0.239055f
C1070 _098_ net71 1.076897f
C1071 output38/a_224_472# net66 0.148811f
C1072 _083_ vdd 0.157549f
C1073 _078_ vss 0.367953f
C1074 FILLER_0_2_111/a_36_472# _157_ 0.104961f
C1075 net64 net18 1.557441f
C1076 output46/a_224_472# net43 0.10562f
C1077 net58 cal_itt\[0\] 0.229955f
C1078 _153_ _156_ 0.539362f
C1079 net79 _005_ 1.006306f
C1080 cal_itt\[3\] _072_ 2.019868f
C1081 _079_ vdd 0.476075f
C1082 net80 _137_ 0.260786f
C1083 _182_ vdd 0.161134f
C1084 _096_ vss 0.126096f
C1085 FILLER_0_21_286/a_36_472# net18 0.18097f
C1086 _103_ net18 0.11279f
C1087 FILLER_0_10_37/a_36_472# vdd 0.141896f
C1088 net31 net18 0.114197f
C1089 _452_/a_36_151# vdd 0.109842f
C1090 _092_ vdd 0.140213f
C1091 _015_ net64 1.212892f
C1092 _137_ vdd 0.945976f
C1093 _077_ net15 0.238832f
C1094 _068_ calibrate 0.110297f
C1095 _180_ vss 0.106022f
C1096 _049_ vdd 0.199608f
C1097 _176_ cal_count\[1\] 0.297763f
C1098 _128_ _068_ 0.863174f
C1099 net63 net21 0.278824f
C1100 _072_ _061_ 0.448032f
C1101 _079_ _073_ 0.234533f
C1102 _081_ _122_ 2.557248f
C1103 _081_ _169_ 0.260462f
C1104 _064_ net17 0.108825f
C1105 net65 net64 0.119915f
C1106 input5/a_36_113# net59 0.257143f
C1107 output25/a_224_472# net25 0.179738f
C1108 mask\[7\] mask\[6\] 0.227476f
C1109 net75 _074_ 1.343862f
C1110 net50 net14 0.192231f
C1111 _176_ _120_ 0.169846f
C1112 _053_ _077_ 0.123663f
C1113 vdd _416_/a_36_151# 0.142481f
C1114 result[9] vss 0.348416f
C1115 _093_ _103_ 0.124026f
C1116 net32 vdd 0.50705f
C1117 net81 cal_itt\[1\] 0.387207f
C1118 _150_ net36 0.108945f
C1119 net31 _093_ 0.274432f
C1120 ctln[1] clk 0.551557f
C1121 _035_ _034_ 1.26804f
C1122 _077_ FILLER_0_12_50/a_36_472# 0.177624f
C1123 trim_val\[4\] _170_ 0.281942f
C1124 mask\[4\] _093_ 0.469687f
C1125 _072_ vss 0.439154f
C1126 net75 net19 1.345314f
C1127 _119_ _077_ 2.584241f
C1128 net5 vdd 0.516129f
C1129 _446_/a_36_151# output41/a_224_472# 0.135198f
C1130 _122_ _163_ 0.156898f
C1131 net44 vdd 0.897202f
C1132 mask\[0\] _138_ 0.22533f
C1133 net20 _046_ 0.194455f
C1134 _041_ vdd 0.19154f
C1135 net27 net64 1.364577f
C1136 _105_ net33 0.202272f
C1137 output43/a_224_472# net43 0.11662f
C1138 _071_ vss 0.126519f
C1139 _055_ _060_ 0.181186f
C1140 net46 vdd 0.255965f
C1141 result[8] mask\[7\] 0.110637f
C1142 mask\[3\] _137_ 0.231419f
C1143 net52 _170_ 0.378738f
C1144 _055_ vdd 0.406945f
C1145 net20 net64 0.374636f
C1146 _116_ _055_ 0.72331f
C1147 _126_ vdd 0.682779f
C1148 _095_ vss 1.465527f
C1149 _036_ vss 0.161195f
C1150 trim_val\[3\] _168_ 0.271475f
C1151 _115_ vdd 0.455713f
C1152 net20 _103_ 0.261438f
C1153 vss net14 1.003274f
C1154 net2 net5 0.47659f
C1155 net34 _009_ 0.325819f
C1156 _126_ _118_ 0.215385f
C1157 net20 net31 0.238809f
C1158 trim_mask\[3\] vdd 0.233305f
C1159 _164_ vss 0.597051f
C1160 result[1] vdd 0.221634f
C1161 ctln[8] vdd 0.125219f
C1162 ctlp[3] vdd 0.251098f
C1163 trim_mask\[1\] _164_ 0.195956f
C1164 net16 _064_ 0.121797f
C1165 _115_ _118_ 1.045555f
C1166 net35 _148_ 0.114816f
C1167 net79 result[3] 0.138076f
C1168 state\[1\] vdd 0.544231f
C1169 net38 _054_ 0.640545f
C1170 _086_ _061_ 0.152228f
C1171 net75 net48 0.10167f
C1172 _116_ state\[1\] 0.693219f
C1173 net38 vss 0.633752f
C1174 _104_ vss 0.564464f
C1175 net52 _168_ 0.726039f
C1176 _056_ _076_ 0.938912f
C1177 _155_ net14 0.10433f
C1178 _144_ vss 0.411237f
C1179 _153_ vss 0.256017f
C1180 FILLER_0_8_37/a_572_375# _054_ 0.137749f
C1181 net57 _061_ 0.127011f
C1182 _076_ _068_ 0.35956f
C1183 FILLER_0_8_37/a_36_472# vdd 0.135405f
C1184 _132_ _126_ 0.247838f
C1185 _161_ _090_ 0.207838f
C1186 _044_ net62 0.101165f
C1187 net34 net33 0.509436f
C1188 result[5] net60 0.16275f
C1189 _001_ _082_ 0.46787f
C1190 net50 trim_mask\[2\] 0.267074f
C1191 net41 _063_ 0.105528f
C1192 _053_ _062_ 0.185944f
C1193 _091_ _069_ 0.741596f
C1194 cal_itt\[2\] net75 0.143064f
C1195 _004_ net81 0.993594f
C1196 _086_ vss 0.615299f
C1197 _098_ vss 0.958032f
C1198 _056_ _090_ 0.177189f
C1199 output10/a_224_472# vdd 0.107357f
C1200 cal_itt\[3\] calibrate 1.141592f
C1201 result[6] vss 0.310169f
C1202 _081_ _152_ 0.172002f
C1203 net33 _146_ 0.306187f
C1204 _133_ vdd 0.27652f
C1205 _070_ vss 1.363355f
C1206 mask\[9\] _098_ 0.256513f
C1207 net34 net35 2.497277f
C1208 _126_ net74 1.001749f
C1209 net46 net43 0.215092f
C1210 net58 _084_ 0.141836f
C1211 _064_ net40 0.141744f
C1212 _002_ net76 0.213703f
C1213 _161_ _117_ 0.25528f
C1214 net57 vss 0.818311f
C1215 net55 vss 0.947665f
C1216 ctln[2] vss 0.256543f
C1217 _020_ _137_ 0.228674f
C1218 _088_ vss 0.326434f
C1219 FILLER_0_18_177/a_36_472# vdd 0.110153f
C1220 net17 vss 0.940703f
C1221 _077_ _115_ 0.131611f
C1222 net82 vss 0.550252f
C1223 trim_val\[1\] trim_mask\[1\] 0.519723f
C1224 _128_ _061_ 0.76584f
C1225 _158_ vdd 0.131365f
C1226 _014_ calibrate 0.403103f
C1227 _121_ vdd 0.106437f
C1228 net22 _047_ 0.132529f
C1229 _112_ _122_ 0.120159f
C1230 net18 _044_ 0.174456f
C1231 _111_ vss 0.233815f
C1232 ctlp[2] net78 0.369805f
C1233 _093_ net71 0.133323f
C1234 output40/a_224_472# output41/a_224_472# 0.292611f
C1235 _090_ _113_ 0.263235f
C1236 _443_/a_36_151# vdd 0.175472f
C1237 net41 net72 0.319547f
C1238 _111_ mask\[9\] 0.127919f
C1239 ctlp[2] vss 0.131085f
C1240 _427_/a_36_151# vdd 0.107344f
C1241 vdd _047_ 0.175913f
C1242 net58 net4 0.858616f
C1243 _127_ cal_count\[3\] 0.306114f
C1244 result[5] vdd 0.142481f
C1245 _027_ net36 0.185347f
C1246 _028_ _154_ 0.174927f
C1247 output24/a_224_472# net54 0.177947f
C1248 calibrate vss 1.140031f
C1249 _122_ vdd 0.379907f
C1250 FILLER_0_16_37/a_36_472# vdd 0.142203f
C1251 net64 vdd 1.155692f
C1252 _094_ mask\[1\] 0.49634f
C1253 _095_ net36 0.127549f
C1254 _128_ vss 0.859962f
C1255 _050_ mask\[7\] 0.128172f
C1256 trim_val\[2\] vdd 0.160419f
C1257 trim_mask\[2\] vss 0.182675f
C1258 _067_ net17 0.17227f
C1259 clk vss 0.210484f
C1260 trim_val\[4\] _037_ 0.258184f
C1261 _419_/a_36_151# vdd -0.110366f
C1262 _103_ vdd 0.590261f
C1263 _377_/a_36_472# trim_val\[0\] 0.135527f
C1264 net31 vdd 0.542738f
C1265 mask\[7\] vss 0.85153f
C1266 _101_ _099_ 0.198807f
C1267 net57 net23 0.324262f
C1268 _122_ _123_ 0.242965f
C1269 _072_ _176_ 0.298077f
C1270 cal net18 0.123815f
C1271 mask\[7\] _107_ 0.13732f
C1272 net74 _133_ 0.696379f
C1273 mask\[1\] vss 0.46268f
C1274 _091_ _137_ 0.486022f
C1275 mask\[4\] vdd 0.794539f
C1276 ctln[1] net20 0.135151f
C1277 _174_ vdd 0.18623f
C1278 net82 net23 0.18994f
C1279 mask\[5\] _144_ 0.38642f
C1280 _094_ _099_ 0.193065f
C1281 _097_ vdd 0.191424f
C1282 net72 _052_ 0.138281f
C1283 trim_val\[4\] net22 0.144267f
C1284 mask\[2\] vdd 0.433058f
C1285 _064_ output39/a_224_472# 0.107406f
C1286 mask\[0\] vss 0.694674f
C1287 _032_ vdd 0.174834f
C1288 cal_itt\[3\] _162_ 0.141474f
C1289 trim_val\[4\] vdd 0.245329f
C1290 fanout63/a_36_160# _282_/a_36_160# 0.23939f
C1291 trimb[3] vdd 0.283005f
C1292 net16 vss 0.679042f
C1293 _099_ vss 0.255039f
C1294 output28/a_224_472# net19 0.101711f
C1295 net52 _037_ 0.103749f
C1296 net51 net6 0.142515f
C1297 result[5] net77 0.142532f
C1298 _085_ _055_ 0.240451f
C1299 net75 net81 0.420021f
C1300 mask\[5\] _098_ 1.316993f
C1301 output33/a_224_472# output19/a_224_472# 0.115114f
C1302 trim_val\[3\] vdd 0.211478f
C1303 net48 _074_ 1.192591f
C1304 vss net62 1.17087f
C1305 output43/a_224_472# output45/a_224_472# 0.246888f
C1306 FILLER_0_22_177/a_36_472# vdd 0.111906f
C1307 _053_ net59 0.145863f
C1308 _140_ _146_ 0.135012f
C1309 net36 _098_ 3.387566f
C1310 result[7] _009_ 0.697145f
C1311 _419_/a_36_151# net77 0.163616f
C1312 net32 _105_ 2.08459f
C1313 net47 _169_ 0.528536f
C1314 _062_ _055_ 0.29425f
C1315 _149_ _026_ 0.243704f
C1316 valid net59 0.577796f
C1317 _077_ _122_ 0.144611f
C1318 mask\[7\] net23 0.225177f
C1319 net58 net37 0.15273f
C1320 net67 net6 0.345681f
C1321 _085_ state\[1\] 0.182697f
C1322 net61 net78 1.588656f
C1323 net55 net36 0.273956f
C1324 trim[0] vss 0.132654f
C1325 net4 _078_ 0.487587f
C1326 _008_ _104_ 0.135471f
C1327 net52 vdd 1.32956f
C1328 net50 _168_ 0.306226f
C1329 net61 vss 0.254538f
C1330 _094_ net18 0.468109f
C1331 _065_ ctln[8] 0.193903f
C1332 net76 net37 0.549565f
C1333 FILLER_0_7_72/a_36_472# vdd 0.106377f
C1334 _098_ net21 0.133694f
C1335 _083_ net59 0.408831f
C1336 _111_ net36 0.102444f
C1337 _175_ cal_count\[1\] 0.203153f
C1338 net78 net18 1.351707f
C1339 mask\[5\] ctlp[2] 0.104304f
C1340 ctln[4] vss 0.244634f
C1341 output31/a_224_472# net30 0.149277f
C1342 _161_ vdd 0.262564f
C1343 ctln[1] net8 0.678616f
C1344 _036_ _030_ 0.430683f
C1345 _129_ vdd 0.314544f
C1346 _131_ vss 0.549133f
C1347 ctlp[8] vss 0.107975f
C1348 _079_ net59 0.102335f
C1349 vss net40 0.898805f
C1350 mask\[4\] mask\[3\] 1.118454f
C1351 trim_val\[4\] trim_mask\[4\] 0.152123f
C1352 net18 vss 1.110302f
C1353 net56 vss 0.367812f
C1354 _095_ _406_/a_36_159# 0.131137f
C1355 _155_ _151_ 0.10611f
C1356 _129_ _118_ 0.213736f
C1357 net74 _032_ 0.208799f
C1358 fanout70/a_36_113# net73 0.21211f
C1359 net22 mask\[6\] 0.612004f
C1360 _056_ vdd 0.423512f
C1361 _086_ _176_ 0.837546f
C1362 result[4] net60 0.244453f
C1363 _170_ vss 0.280383f
C1364 trim[0] net66 0.376153f
C1365 _116_ _056_ 0.30649f
C1366 net16 _166_ 0.146913f
C1367 _068_ vdd 0.793549f
C1368 _076_ vss 1.132839f
C1369 net32 net34 0.330134f
C1370 fanout61/a_36_113# vdd 0.108255f
C1371 trimb[3] net43 0.221036f
C1372 net19 net33 0.254336f
C1373 _176_ _070_ 0.467961f
C1374 mask\[6\] vdd 0.573103f
C1375 _019_ mask\[2\] 0.155325f
C1376 net69 vdd 1.102677f
C1377 _068_ _118_ 1.374452f
C1378 _070_ _124_ 0.114614f
C1379 net57 _176_ 0.192223f
C1380 net55 _176_ 0.300149f
C1381 net16 cal_count\[0\] 0.152321f
C1382 _152_ vdd 0.354509f
C1383 _081_ vss 0.733408f
C1384 trimb[0] vdd 0.10929f
C1385 _093_ vss 2.002012f
C1386 net65 vss 0.471168f
C1387 net31 output34/a_224_472# 0.165772f
C1388 _133_ _062_ 1.210949f
C1389 net36 mask\[1\] 0.28584f
C1390 _013_ vdd 0.372605f
C1391 net66 net40 0.124825f
C1392 ctln[1] vdd 0.825166f
C1393 _093_ mask\[9\] 0.460108f
C1394 _120_ net51 1.716752f
C1395 fanout51/a_36_113# FILLER_0_11_78/a_36_472# 0.193759f
C1396 _090_ vss 0.267577f
C1397 _113_ vdd 0.774039f
C1398 _116_ _113_ 0.179616f
C1399 _168_ vss 0.171346f
C1400 _029_ vss 0.11129f
C1401 net5 net59 0.923076f
C1402 net71 vdd 0.775031f
C1403 _029_ trim_mask\[1\] 1.002118f
C1404 _108_ vss 0.160825f
C1405 net58 net1 0.626432f
C1406 net56 net23 0.930833f
C1407 net36 _099_ 0.325141f
C1408 _078_ net37 0.459092f
C1409 _129_ net74 0.476969f
C1410 en_co_clk _067_ 0.272082f
C1411 result[8] net22 0.278936f
C1412 _136_ net14 0.417108f
C1413 _163_ vss 0.638066f
C1414 _075_ cal_itt\[3\] 0.731221f
C1415 _170_ _066_ 0.189122f
C1416 net28 net79 0.116857f
C1417 _064_ vdd 0.874293f
C1418 trim_mask\[1\] _163_ 0.166315f
C1419 _053_ _165_ 0.123461f
C1420 net54 net71 0.536043f
C1421 net23 _170_ 0.107532f
C1422 _087_ net37 0.23484f
C1423 net53 _095_ 0.431214f
C1424 net42 vdd 0.178782f
C1425 output44/a_224_472# net38 0.106923f
C1426 _128_ _176_ 0.180252f
C1427 _155_ _029_ 0.174512f
C1428 _076_ net23 0.105196f
C1429 result[4] vdd 0.205815f
C1430 net81 net79 0.178225f
C1431 net20 _094_ 0.677838f
C1432 result[8] vdd 0.590386f
C1433 net27 vss 0.534444f
C1434 _128_ _124_ 0.111918f
C1435 net19 net9 0.342451f
C1436 _122_ _062_ 0.190871f
C1437 cal net8 0.271166f
C1438 _077_ _056_ 1.777574f
C1439 trim_mask\[4\] net69 0.185121f
C1440 ctln[1] net2 0.126801f
C1441 vdd _156_ 0.178622f
C1442 _044_ vdd 0.406979f
C1443 net20 net78 1.100401f
C1444 trim_mask\[4\] _152_ 0.224909f
C1445 _077_ _068_ 0.601166f
C1446 net58 net76 0.700034f
C1447 _152_ net47 0.242864f
C1448 _155_ _163_ 0.296236f
C1449 net74 net69 0.143604f
C1450 net20 vss 1.402494f
C1451 _064_ net39 0.558387f
C1452 net74 _152_ 1.007413f
C1453 _126_ cal_count\[3\] 0.418508f
C1454 _058_ net14 0.40635f
C1455 _098_ FILLER_0_15_180/a_36_472# 0.101593f
C1456 trimb[0] net43 0.109028f
C1457 ctln[9] vss 0.167242f
C1458 net28 net19 0.115252f
C1459 trim_mask\[2\] _030_ 1.467465f
C1460 _053_ _074_ 0.503728f
C1461 FILLER_0_13_65/a_36_472# fanout72/a_36_113# 0.193651f
C1462 _144_ _145_ 0.671767f
C1463 net81 net19 0.786284f
C1464 FILLER_0_1_98/a_36_472# trim_mask\[3\] 0.106084f
C1465 net56 net36 0.772486f
C1466 cal_count\[3\] state\[1\] 0.236393f
C1467 net18 _193_/a_36_160# 0.114176f
C1468 cal_count\[1\] _180_ 0.300952f
C1469 output8/a_224_472# _411_/a_36_151# 0.12978f
C1470 en net18 0.32189f
C1471 _442_/a_36_151# vdd 0.102701f
C1472 net57 _136_ 0.168299f
C1473 _064_ net47 0.110169f
C1474 cal vdd 0.318671f
C1475 mask\[4\] _143_ 0.352305f
C1476 net60 _094_ 0.579872f
C1477 net42 net47 0.237866f
C1478 vss _039_ 0.180364f
C1479 _149_ net14 0.102004f
C1480 _119_ _074_ 0.153267f
C1481 net68 net67 0.147318f
C1482 FILLER_0_12_2/a_36_472# vdd 0.104425f
C1483 net67 clkc 0.102244f
C1484 net4 _070_ 0.169392f
C1485 _065_ trim_val\[3\] 1.235816f
C1486 output37/a_224_472# net64 0.110037f
C1487 net50 vdd 0.661261f
C1488 fanout68/a_36_113# _441_/a_36_151# 0.138322f
C1489 cal_itt\[3\] net22 0.134309f
C1490 net60 vss 0.382678f
C1491 FILLER_0_13_212/a_36_472# vdd 0.105926f
C1492 net25 FILLER_0_23_88/a_36_472# 0.192699f
C1493 _093_ net36 0.214976f
C1494 _091_ mask\[2\] 2.252217f
C1495 ctlp[4] net22 0.257841f
C1496 output29/a_224_472# net62 0.138536f
C1497 net35 net33 1.594925f
C1498 FILLER_0_20_2/a_36_472# vdd 0.102471f
C1499 _438_/a_36_151# vdd 0.111691f
C1500 net82 net4 1.982825f
C1501 net31 net30 0.130396f
C1502 cal_itt\[3\] vdd 0.571239f
C1503 ctlp[4] vdd 0.278868f
C1504 _061_ net22 0.123662f
C1505 _176_ _131_ 1.798819f
C1506 net8 vss 0.171128f
C1507 _008_ net18 0.113775f
C1508 _057_ _071_ 0.139904f
C1509 _067_ _039_ 0.221585f
C1510 ctln[3] vdd 0.167569f
C1511 _061_ vdd 0.295557f
C1512 _311_/a_66_473# vdd 0.106886f
C1513 _129_ _062_ 0.20212f
C1514 _001_ vdd 0.122898f
C1515 FILLER_0_13_228/a_124_375# _043_ 0.133079f
C1516 FILLER_0_8_107/a_36_472# vdd 0.117254f
C1517 _149_ _098_ 0.398643f
C1518 FILLER_0_4_185/a_36_472# vdd 0.122463f
C1519 net32 result[7] 0.103491f
C1520 _061_ _118_ 0.268815f
C1521 _112_ vss 0.145781f
C1522 output8/a_224_472# _000_ 0.182377f
C1523 _087_ net76 0.529571f
C1524 _031_ vdd 0.327674f
C1525 cal_count\[2\] _180_ 0.153207f
C1526 _136_ mask\[1\] 0.407932f
C1527 _094_ vdd 0.717159f
C1528 _056_ _062_ 0.320621f
C1529 _096_ _043_ 0.842762f
C1530 _008_ _093_ 0.252609f
C1531 net22 vss 1.28233f
C1532 net78 vdd 0.265913f
C1533 _050_ vdd 0.484554f
C1534 net15 net72 0.157843f
C1535 _095_ cal_count\[1\] 0.853949f
C1536 output40/a_224_472# trim[3] 0.122003f
C1537 net80 vss 0.347557f
C1538 trim[4] net44 0.188184f
C1539 _054_ vdd 0.360345f
C1540 _060_ vss 0.318005f
C1541 net32 net19 0.65591f
C1542 ctlp[7] vdd 0.481613f
C1543 _033_ net67 0.148585f
C1544 vdd vss 15.42941f
C1545 _077_ net50 0.312283f
C1546 _122_ _059_ 0.190023f
C1547 trim_mask\[1\] vdd 0.241393f
C1548 _116_ vss 0.235141f
C1549 net52 _160_ 0.133292f
C1550 _039_ cal_count\[0\] 0.219667f
C1551 _118_ vss 0.217218f
C1552 mask\[9\] vdd 0.940144f
C1553 ctln[3] net10 0.873575f
C1554 net54 vss 0.715177f
C1555 _073_ vss 0.216342f
C1556 net31 _006_ 0.307613f
C1557 output36/a_224_472# net62 0.317201f
C1558 result[1] net79 0.25261f
C1559 valid sample 0.103192f
C1560 _086_ _057_ 0.82902f
C1561 output38/a_224_472# _446_/a_36_151# 0.117966f
C1562 _155_ vdd 0.193832f
C1563 net39 vss 0.170972f
C1564 result[0] vss 0.291352f
C1565 _094_ _045_ 0.102437f
C1566 _450_/a_36_151# output6/a_224_472# 0.134892f
C1567 _057_ net57 0.873864f
C1568 _132_ vss 0.492496f
C1569 _424_/a_36_151# vdd 0.125156f
C1570 net66 vdd 0.646189f
C1571 _067_ vdd 0.853589f
C1572 net78 net77 0.252376f
C1573 net2 vss 0.213737f
C1574 net10 vss 0.324553f
C1575 _132_ mask\[9\] 0.203851f
C1576 _008_ net20 0.153014f
C1577 cal_itt\[2\] _083_ 0.10423f
C1578 _064_ trim[1] 0.166575f
C1579 net77 vss 0.327705f
C1580 net35 _140_ 0.12583f
C1581 _144_ mask\[8\] 0.131592f
C1582 net28 _192_/a_67_603# 0.119061f
C1583 ctln[7] net14 0.197449f
C1584 _066_ vdd 0.14893f
C1585 _131_ _136_ 1.42765f
C1586 net47 _054_ 0.171966f
C1587 _152_ _160_ 0.286108f
C1588 output47/a_224_472# net55 0.160037f
C1589 net25 vdd 0.195306f
C1590 net23 vdd 1.576398f
C1591 trim_mask\[4\] vss 0.641217f
C1592 net47 vss 0.919407f
C1593 _012_ vss 0.454371f
C1594 calibrate net37 0.101109f
C1595 _141_ _093_ 0.396041f
C1596 net56 _136_ 0.462275f
C1597 _095_ cal_count\[2\] 0.270066f
C1598 trim_mask\[1\] net47 0.306848f
C1599 net55 cal_count\[1\] 0.204733f
C1600 _118_ net23 0.108864f
C1601 _086_ _120_ 0.408014f
C1602 net74 vss 0.589483f
C1603 _103_ _102_ 0.392644f
C1604 _077_ vss 1.071923f
C1605 vdd _166_ 0.108744f
C1606 _095_ _043_ 2.807456f
C1607 _159_ vss 0.102545f
C1608 net43 vss 0.132286f
C1609 mask\[3\] vss 0.664467f
C1610 net22 _205_/a_36_160# 0.109939f
C1611 _070_ _120_ 0.838223f
C1612 FILLER_0_3_142/a_36_472# vdd 0.10948f
C1613 net68 _036_ 0.168017f
C1614 _114_ _126_ 3.341247f
C1615 ctlp[1] vss 0.32843f
C1616 net52 cal_count\[3\] 0.348542f
C1617 vdd cal_count\[0\] 0.491891f
C1618 net68 _164_ 0.189377f
C1619 _114_ _115_ 0.148291f
C1620 ctln[4] net11 0.194506f
C1621 _019_ vss 0.10954f
C1622 net57 fanout52/a_36_160# 0.122432f
C1623 net29 _099_ 0.358926f
C1624 cal_itt\[1\] vss 0.327626f
C1625 cal_itt\[0\] vdd 0.438996f
C1626 _093_ _136_ 0.226819f
C1627 net57 state\[2\] 1.25275f
C1628 net4 _076_ 1.140706f
C1629 _028_ _163_ 0.199021f
C1630 net38 _043_ 0.117134f
C1631 net55 _175_ 0.142124f
C1632 net34 mask\[6\] 0.231853f
C1633 net66 net47 0.238874f
C1634 _008_ net60 0.314106f
C1635 _086_ _125_ 0.490983f
C1636 net32 net33 0.467071f
C1637 _185_ cal_count\[2\] 0.205002f
C1638 mask\[5\] vdd 0.79138f
C1639 net74 _067_ 0.674895f
C1640 net38 net67 1.762405f
C1641 _156_ _160_ 0.299745f
C1642 _073_ cal_itt\[0\] 0.211566f
C1643 result[4] net30 0.298966f
C1644 sample net5 0.359975f
C1645 net65 net4 0.614946f
C1646 result[9] _010_ 0.121471f
C1647 trim_mask\[4\] _066_ 0.396509f
C1648 _056_ cal_count\[3\] 0.186969f
C1649 _070_ _125_ 0.125523f
C1650 _076_ _058_ 0.912225f
C1651 net36 vdd 0.939735f
C1652 trim_mask\[4\] net23 0.180803f
C1653 mask\[6\] _146_ 0.181681f
C1654 mask\[7\] _024_ 0.122185f
C1655 net70 vss 0.175272f
C1656 _065_ net50 0.123581f
C1657 _068_ _059_ 0.255081f
C1658 output35/a_224_472# net33 0.170613f
C1659 net72 _041_ 0.467856f
C1660 en vdd 0.282941f
C1661 FILLER_0_9_142/a_36_472# vdd 0.107619f
C1662 _131_ _134_ 0.887647f
C1663 net22 net21 1.937266f
C1664 net81 valid 0.11798f
C1665 _040_ vss 0.216709f
C1666 _026_ _098_ 0.197713f
C1667 FILLER_0_3_142/a_124_375# net23 0.25251f
C1668 trimb[4] cal_count\[2\] 0.146942f
C1669 ctln[1] net75 0.159105f
C1670 _088_ net76 0.214494f
C1671 _154_ _153_ 0.719561f
C1672 net57 _043_ 1.955053f
C1673 _074_ _122_ 0.300373f
C1674 _021_ FILLER_0_18_171/a_36_472# 0.103755f
C1675 net21 vdd 1.653552f
C1676 output43/a_224_472# output46/a_224_472# 0.292611f
C1677 _061_ _062_ 0.344031f
C1678 _250_/a_36_68# _071_ 0.199512f
C1679 output33/a_224_472# output18/a_224_472# 0.111946f
C1680 result[7] _103_ 0.298427f
C1681 net17 _043_ 0.571818f
C1682 net63 mask\[1\] 0.120872f
C1683 net31 result[7] 0.231528f
C1684 net7 vss 0.117948f
C1685 net68 net17 0.601273f
C1686 _120_ _171_ 0.414533f
C1687 _173_ cal_count\[0\] 0.517178f
C1688 _276_/a_36_160# _291_/a_36_160# 0.239422f
C1689 net58 calibrate 0.205792f
C1690 _104_ _106_ 0.17237f
C1691 _165_ trim_val\[0\] 0.164683f
C1692 _086_ _154_ 0.102849f
C1693 _008_ vdd 0.284571f
C1694 _093_ FILLER_0_18_76/a_36_472# 0.129892f
C1695 _085_ vss 0.132721f
C1696 _176_ vdd 0.874707f
C1697 _005_ _044_ 0.50767f
C1698 output16/a_224_472# _447_/a_36_151# 0.200384f
C1699 net20 net4 0.650415f
C1700 net58 output27/a_224_472# 0.121438f
C1701 _176_ _118_ 0.392531f
C1702 _413_/a_36_151# vdd 0.130213f
C1703 _062_ vss 0.58133f
C1704 result[4] _006_ 0.271278f
C1705 _118_ _124_ 0.652002f
C1706 _004_ _094_ 0.213913f
C1707 output33/a_224_472# net18 0.110644f
C1708 _065_ vss 0.230397f
C1709 _072_ _071_ 0.296543f
C1710 trimb[1] net38 0.161478f
C1711 _127_ _126_ 0.398279f
C1712 _081_ net37 1.274337f
C1713 output29/a_224_472# vdd 0.103437f
C1714 _178_ _278_/a_36_160# 0.269109f
C1715 output9/a_224_472# net18 0.114757f
C1716 _178_ vss 0.150839f
C1717 _104_ _010_ 0.252687f
C1718 _094_ _007_ 0.170362f
C1719 _136_ _139_ 0.394888f
C1720 net26 net17 0.132516f
C1721 _004_ vss 0.115789f
C1722 _110_ vss 0.131865f
C1723 _177_ net36 0.371814f
C1724 _030_ vdd 0.244909f
C1725 mask\[8\] _354_/a_49_472# 0.105272f
C1726 _019_ net36 0.309649f
C1727 _104_ result[9] 0.169685f
C1728 net5 rstn 0.101356f
C1729 net41 _064_ 0.301777f
C1730 cal_count\[2\] _179_ 0.404284f
C1731 _079_ _083_ 0.872842f
C1732 net3 cal_count\[2\] 0.119728f
C1733 _091_ vss 0.56693f
C1734 cal net59 0.297816f
C1735 _131_ _120_ 0.191602f
C1736 mask\[3\] net21 0.100738f
C1737 net13 vdd 0.264116f
C1738 mask\[0\] _043_ 0.929722f
C1739 _057_ _090_ 0.112325f
C1740 _013_ _052_ 0.284735f
C1741 fanout54/a_36_160# FILLER_0_19_155/a_36_472# 0.193804f
C1742 _095_ _184_ 0.265966f
C1743 net48 _122_ 0.110769f
C1744 _094_ net30 0.188507f
C1745 _064_ net49 0.377675f
C1746 _105_ vss 0.485198f
C1747 _069_ _055_ 0.741952f
C1748 net16 net68 0.275467f
C1749 vss _160_ 1.119894f
C1750 _074_ _161_ 0.191658f
C1751 _141_ vdd 0.439746f
C1752 _008_ mask\[3\] 0.799138f
C1753 net74 _124_ 0.180235f
C1754 net22 _048_ 0.268142f
C1755 _076_ _120_ 0.736844f
C1756 _028_ vdd 0.626868f
C1757 _002_ vdd 0.152662f
C1758 vss net30 0.17209f
C1759 net36 _040_ 0.429029f
C1760 _048_ vdd 0.270091f
C1761 _086_ _072_ 0.220767f
C1762 _057_ _117_ 0.120323f
C1763 _084_ vdd 0.134578f
C1764 fanout55/a_36_160# _067_ 0.126784f
C1765 _177_ _176_ 0.226424f
C1766 net15 ctln[8] 0.205163f
C1767 _064_ _034_ 1.397143f
C1768 sample net64 0.209777f
C1769 _039_ net6 0.104745f
C1770 net63 _093_ 0.109689f
C1771 _072_ _070_ 2.141346f
C1772 result[2] net62 0.311075f
C1773 net57 _072_ 0.108982f
C1774 _136_ vdd 1.020301f
C1775 cal_count\[2\] net40 0.313209f
C1776 net1 _081_ 0.111227f
C1777 FILLER_0_15_2/a_36_472# vdd 0.104741f
C1778 output36/a_224_472# vdd 0.145046f
C1779 result[9] ctlp[2] 0.105977f
C1780 _153_ net14 0.260217f
C1781 net16 net26 0.273031f
C1782 _005_ _094_ 0.162984f
C1783 _363_/a_36_68# _154_ 0.149319f
C1784 net72 _174_ 0.199504f
C1785 net75 _014_ 0.204357f
C1786 net53 vdd 0.78288f
C1787 net34 vss 0.481379f
C1788 net4 _060_ 0.327437f
C1789 net4 vdd 1.218939f
C1790 FILLER_0_9_72/a_36_472# vdd 0.109576f
C1791 net58 net65 1.468105f
C1792 net67 net40 0.886781f
C1793 net57 _071_ 0.12089f
C1794 _151_ _154_ 0.108571f
C1795 net59 vss 1.191297f
C1796 net50 net49 0.238748f
C1797 _176_ _040_ 0.272465f
C1798 _376_/a_36_160# FILLER_0_6_90/a_36_472# 0.195478f
C1799 ctln[1] _000_ 0.223573f
C1800 _422_/a_36_151# vdd 0.177717f
C1801 output32/a_224_472# _419_/a_36_151# 0.129117f
C1802 net76 _081_ 0.706096f
C1803 _058_ vdd 0.511536f
C1804 net11 vdd 0.330644f
C1805 _166_ _160_ 0.492224f
C1806 net75 vss 0.662689f
C1807 _072_ calibrate 0.539702f
C1808 _114_ _068_ 1.097353f
C1809 net76 net65 0.14935f
C1810 _070_ net14 0.536953f
C1811 cal_count\[3\] vss 1.35143f
C1812 _093_ _150_ 0.406318f
C1813 _059_ vss 0.714648f
C1814 result[7] result[8] 0.201281f
C1815 trimb[2] trimb[3] 0.369908f
C1816 mask\[3\] _141_ 0.361692f
C1817 _095_ net17 0.172789f
C1818 ctln[5] vss 0.132862f
C1819 _006_ vss 0.111492f
C1820 ctln[0] vss 0.125714f
C1821 _036_ net17 0.153479f
C1822 _069_ _121_ 0.137961f
C1823 trim_val\[1\] _164_ 0.100504f
C1824 _144_ _098_ 1.252524f
C1825 net2 net4 0.854661f
C1826 net38 net55 0.10956f
C1827 _142_ _137_ 1.401722f
C1828 net16 _447_/a_36_151# 0.133348f
C1829 mask\[5\] _105_ 0.706158f
C1830 _149_ vdd 0.379674f
C1831 trimb[4] net38 0.124219f
C1832 _114_ _113_ 0.201729f
C1833 mask\[0\] FILLER_0_14_235/a_36_472# 0.287093f
C1834 _053_ _133_ 0.288819f
C1835 _408_/a_56_524# _043_ 0.10151f
C1836 vdd net6 0.134918f
C1837 net38 net17 1.634286f
C1838 net58 net27 0.190417f
C1839 mask\[0\] _018_ 0.328328f
C1840 net73 _093_ 0.350073f
C1841 _134_ vdd 0.482157f
C1842 result[9] net62 0.339372f
C1843 cal_itt\[1\] _084_ 0.495918f
C1844 net19 _044_ 0.138869f
C1845 _102_ _094_ 0.727442f
C1846 net53 net74 0.164124f
C1847 net41 vss 0.810444f
C1848 net54 _149_ 0.212511f
C1849 _434_/a_36_151# vdd 0.104871f
C1850 cal_count\[3\] _067_ 0.478427f
C1851 _120_ _039_ 0.148356f
C1852 _187_ cal_count\[0\] 0.645851f
C1853 output7/a_224_472# trim[3] 0.103375f
C1854 net29 vdd 0.611195f
C1855 trim_mask\[2\] _036_ 0.466145f
C1856 _077_ net4 0.656292f
C1857 _086_ _070_ 0.123033f
C1858 _185_ net17 0.270086f
C1859 _104_ ctlp[2] 1.420577f
C1860 _033_ net40 0.298492f
C1861 _086_ net57 0.126563f
C1862 _345_/a_36_160# vdd 0.100094f
C1863 trim_mask\[2\] _164_ 1.859062f
C1864 net49 vss 0.689397f
C1865 vdd trim[3] 0.147228f
C1866 net81 net64 0.455159f
C1867 _029_ _154_ 0.116532f
C1868 _059_ net23 0.265909f
C1869 net37 vdd 0.544653f
C1870 _016_ _130_ 0.114514f
C1871 net57 _070_ 0.202843f
C1872 _181_ cal_count\[1\] 0.186904f
C1873 _057_ net22 0.163773f
C1874 FILLER_0_15_72/a_36_472# vdd 0.108844f
C1875 _077_ _058_ 3.018054f
C1876 _035_ vss 0.105648f
C1877 FILLER_0_5_128/a_36_472# _360_/a_36_160# 0.195479f
C1878 _078_ _081_ 0.445443f
C1879 _258_/a_36_160# _080_ 0.261387f
C1880 _053_ _122_ 0.368823f
C1881 _163_ _154_ 0.190662f
C1882 net57 net82 0.91473f
C1883 _057_ vdd 0.801978f
C1884 mask\[7\] _147_ 0.295801f
C1885 _088_ net82 0.160444f
C1886 net33 mask\[6\] 0.881813f
C1887 _144_ mask\[7\] 0.111088f
C1888 net47 net6 0.23883f
C1889 net16 _036_ 0.637538f
C1890 net82 _082_ 0.286003f
C1891 _127_ _129_ 0.716384f
C1892 ctln[6] vdd 0.116327f
C1893 net70 net53 1.170795f
C1894 net51 _039_ 0.398642f
C1895 cal_itt\[3\] _074_ 0.584958f
C1896 _136_ _040_ 0.788826f
C1897 output9/a_224_472# vdd 0.102412f
C1898 _119_ _122_ 0.155432f
C1899 _429_/a_36_151# _018_ 0.118135f
C1900 _008_ net30 1.112351f
C1901 vss result[3] 0.28152f
C1902 net29 _045_ 0.344478f
C1903 net66 net49 0.657679f
C1904 net80 _023_ 0.261119f
C1905 net38 net3 0.103189f
C1906 _070_ calibrate 0.675125f
C1907 cal_count\[1\] vdd 0.516859f
C1908 trim_mask\[2\] fanout49/a_36_160# 0.12844f
C1909 net79 _094_ 0.301878f
C1910 _126_ state\[1\] 1.191746f
C1911 _128_ _070_ 1.279188f
C1912 _035_ net66 1.624557f
C1913 en net59 0.490893f
C1914 net58 net8 0.175026f
C1915 net63 net22 0.223664f
C1916 _098_ mask\[1\] 1.476748f
C1917 _425_/a_448_472# calibrate 0.105581f
C1918 vdd FILLER_0_13_72/a_36_472# 0.108152f
C1919 net67 _039_ 0.302826f
C1920 net63 net80 0.337396f
C1921 _120_ vdd 0.750809f
C1922 net79 vss 0.770834f
C1923 _184_ net40 0.122833f
C1924 net69 _157_ 0.112249f
C1925 net15 net52 0.166073f
C1926 net63 vdd 1.002883f
C1927 net66 _034_ 0.139638f
C1928 mask\[8\] vdd 0.423606f
C1929 _181_ cal_count\[2\] 0.375819f
C1930 _118_ _120_ 0.339442f
C1931 _143_ _141_ 0.192528f
C1932 net59 net21 0.157689f
C1933 output23/a_224_472# net23 0.122379f
C1934 state\[2\] vdd 0.392508f
C1935 net20 _078_ 0.105266f
C1936 _053_ trim_val\[0\] 0.446477f
C1937 _175_ vdd 0.147794f
C1938 result[7] vss 0.49466f
C1939 result[8] net33 0.474056f
C1940 _095_ net40 0.674445f
C1941 _036_ net40 0.599505f
C1942 _074_ vss 0.404343f
C1943 net1 vdd 0.63891f
C1944 vdd FILLER_0_6_37/a_36_472# 0.138008f
C1945 _185_ _402_/a_56_567# 0.107713f
C1946 net54 mask\[8\] 0.162104f
C1947 _104_ net61 1.149805f
C1948 _077_ _057_ 0.584179f
C1949 _137_ mask\[2\] 0.440828f
C1950 FILLER_0_20_177/a_36_472# vdd 0.114932f
C1951 net60 _421_/a_36_151# 0.224039f
C1952 net78 net19 0.507249f
C1953 _114_ _061_ 0.123371f
C1954 ctln[7] vdd 0.359832f
C1955 trim_mask\[2\] FILLER_0_2_93/a_36_472# 0.281054f
C1956 _125_ vdd 0.218505f
C1957 net16 trim_val\[1\] 0.164715f
C1958 net38 net40 1.103743f
C1959 _000_ vss 0.205593f
C1960 net58 vdd 0.929215f
C1961 _130_ _127_ 0.195571f
C1962 net19 vss 1.140787f
C1963 net76 net22 0.118787f
C1964 FILLER_0_21_206/a_36_472# net21 0.132984f
C1965 _125_ _118_ 0.239695f
C1966 net51 vdd 0.692054f
C1967 cal_count\[2\] vdd 0.932907f
C1968 input3/a_36_113# vdd 0.117445f
C1969 net20 result[9] 1.593573f
C1970 net76 vdd 1.272072f
C1971 _058_ _062_ 1.676625f
C1972 _093_ net14 0.11038f
C1973 result[6] net61 0.120359f
C1974 ctln[1] rstn 0.62944f
C1975 _043_ vdd 0.827689f
C1976 net1 net2 0.624657f
C1977 net15 _013_ 0.152142f
C1978 _086_ _162_ 0.107276f
C1979 net68 vdd 1.026897f
C1980 _026_ vdd 0.15542f
C1981 _086_ _131_ 0.886615f
C1982 vdd clkc 0.190259f
C1983 _114_ vss 0.365613f
C1984 fanout53/a_36_160# net56 0.196684f
C1985 net58 result[0] 0.443436f
C1986 _140_ mask\[6\] 0.605898f
C1987 _091_ net4 0.125608f
C1988 _077_ _120_ 0.205715f
C1989 fanout65/a_36_113# vdd 0.10473f
C1990 net67 vdd 0.638702f
C1991 _104_ _093_ 0.109158f
C1992 _131_ _070_ 0.161861f
C1993 net48 _014_ 0.276733f
C1994 output42/a_224_472# net42 0.117956f
C1995 net63 mask\[3\] 0.37365f
C1996 net55 _131_ 0.314732f
C1997 net24 vss 0.172755f
C1998 result[2] vdd 0.18482f
C1999 net73 vdd 0.44835f
C2000 ctln[2] net18 0.106494f
C2001 _086_ _076_ 0.79237f
C2002 _063_ vss 0.157186f
C2003 net17 net40 1.095167f
C2004 output22/a_224_472# vdd 0.111234f
C2005 _099_ mask\[1\] 0.19135f
C2006 _063_ trim_mask\[1\] 0.127216f
C2007 net60 _010_ 0.108311f
C2008 _154_ vdd 0.639978f
C2009 _070_ _076_ 0.198272f
C2010 FILLER_0_4_144/a_36_472# _370_/a_848_380# 0.15783f
C2011 net48 vss 0.161385f
C2012 _181_ _180_ 0.216908f
C2013 result[9] net60 0.251903f
C2014 mask\[1\] net62 0.227329f
C2015 _093_ _098_ 0.556613f
C2016 FILLER_0_4_185/a_124_375# _087_ 0.120668f
C2017 net57 en_co_clk 0.195533f
C2018 cal_count\[2\] net47 0.274891f
C2019 net28 _044_ 0.481924f
C2020 fanout64/a_36_160# net65 0.214347f
C2021 net26 vdd 0.487733f
C2022 net1 cal_itt\[1\] 0.229522f
C2023 _009_ vss 0.105833f
C2024 _163_ _153_ 0.243815f
C2025 _021_ net80 0.254353f
C2026 _077_ net51 0.76967f
C2027 _093_ net55 0.182194f
C2028 ctln[2] net65 0.113266f
C2029 _162_ calibrate 0.228839f
C2030 mask\[0\] net62 0.552008f
C2031 _057_ _085_ 0.543871f
C2032 ctlp[5] mask\[7\] 0.131468f
C2033 mask\[3\] FILLER_0_17_161/a_36_472# 0.13873f
C2034 _106_ vdd 0.232973f
C2035 _070_ _090_ 0.369847f
C2036 _132_ net73 0.460325f
C2037 net74 _043_ 0.65119f
C2038 _078_ vdd 0.181583f
C2039 net82 net65 0.630327f
C2040 net58 cal_itt\[1\] 0.79493f
C2041 trim_mask\[2\] net40 0.401672f
C2042 net67 net47 0.126281f
C2043 comp vss 0.148428f
C2044 net19 cal_itt\[0\] 0.111163f
C2045 sample vss 0.276162f
C2046 net72 vss 0.472104f
C2047 cal_itt\[2\] vss 0.249871f
C2048 _093_ _111_ 0.555171f
C2049 _087_ vdd 0.281159f
C2050 net20 _104_ 0.482229f
C2051 _086_ _163_ 0.413768f
C2052 _096_ vdd 0.557569f
C2053 _033_ vdd 0.509957f
C2054 _015_ calibrate 0.105287f
C2055 trim_val\[3\] trim_mask\[3\] 0.48462f
C2056 _076_ calibrate 1.005804f
C2057 _180_ vdd 0.176915f
C2058 net79 net21 0.645949f
C2059 trimb[2] vss 0.102375f
C2060 _070_ _163_ 1.884485f
C2061 net33 vss 0.674927f
C2062 _034_ 0 0.304805f
C2063 _160_ 0 1.542665f
C2064 _166_ 0 0.299751f
C2065 trim[3] 0 1.777626f
C2066 output41/a_224_472# 0 2.38465f
C2067 clkc 0 0.763769f
C2068 net6 0 1.112469f
C2069 output6/a_224_472# 0 2.38465f
C2070 FILLER_0_12_196/a_36_472# 0 0.417394f
C2071 FILLER_0_12_196/a_124_375# 0 0.246306f
C2072 result[3] 0 0.50376f
C2073 net30 0 1.81422f
C2074 output30/a_224_472# 0 2.38465f
C2075 _047_ 0 0.374694f
C2077 net62 0 4.932099f
C2078 _416_/a_2665_112# 0 0.62251f
C2083 _416_/a_36_151# 0 1.43589f
C2084 FILLER_0_13_290/a_36_472# 0 0.417394f
C2085 FILLER_0_13_290/a_124_375# 0 0.246306f
C2086 _278_/a_36_160# 0 0.696445f
C2087 _145_ 0 0.546455f
C2089 FILLER_0_13_72/a_36_472# 0 0.404746f
C2090 FILLER_0_13_72/a_572_375# 0 0.232991f
C2093 FILLER_0_14_235/a_36_472# 0 0.404746f
C2094 FILLER_0_14_235/a_572_375# 0 0.232991f
C2096 _156_ 0 0.593796f
C2097 _107_ 0 0.391583f
C2098 _022_ 0 0.387773f
C2099 _433_/a_2665_112# 0 0.62251f
C2104 _433_/a_36_151# 0 1.43589f
C2106 FILLER_0_5_148/a_36_472# 0 0.404746f
C2107 FILLER_0_5_148/a_572_375# 0 0.232991f
C2109 _167_ 0 0.285904f
C2110 trim[2] 0 0.79181f
C2111 net40 0 1.845219f
C2112 output40/a_224_472# 0 2.38465f
C2113 cal_count\[0\] 0 0.893784f
C2114 _039_ 0 0.412301f
C2120 _450_/a_36_151# 0 1.31409f
C2121 rstn 0 1.86494f
C2123 FILLER_0_8_156/a_36_472# 0 0.404746f
C2124 FILLER_0_8_156/a_572_375# 0 0.232991f
C2126 FILLER_0_6_37/a_36_472# 0 0.417394f
C2127 FILLER_0_6_37/a_124_375# 0 0.246306f
C2129 FILLER_0_21_60/a_36_472# 0 0.404746f
C2130 FILLER_0_21_60/a_572_375# 0 0.232991f
C2133 FILLER_0_22_107/a_36_472# 0 0.404746f
C2134 FILLER_0_22_107/a_572_375# 0 0.232991f
C2136 FILLER_0_16_115/a_36_472# 0 0.417394f
C2137 FILLER_0_16_115/a_124_375# 0 0.246306f
C2138 FILLER_0_19_134/a_36_472# 0 0.417394f
C2139 FILLER_0_19_134/a_124_375# 0 0.246306f
C2140 FILLER_0_3_212/a_36_472# 0 0.417394f
C2141 FILLER_0_3_212/a_124_375# 0 0.246306f
C2143 FILLER_0_10_94/a_36_472# 0 0.404746f
C2144 FILLER_0_10_94/a_572_375# 0 0.232991f
C2147 FILLER_0_4_91/a_36_472# 0 0.404746f
C2148 FILLER_0_4_91/a_572_375# 0 0.232991f
C2150 net14 0 1.508711f
C2151 _202_/a_36_160# 0 0.696445f
C2153 FILLER_0_6_231/a_36_472# 0 0.404746f
C2154 FILLER_0_6_231/a_572_375# 0 0.232991f
C2156 vss 0 65.60368f
C2157 vdd 0 1.086009p
C2158 _006_ 0 0.41456f
C2159 _417_/a_2665_112# 0 0.62251f
C2164 _417_/a_36_151# 0 1.43589f
C2165 _146_ 0 0.35443f
C2166 mask\[6\] 0 1.246962f
C2167 _365_/a_36_68# 0 0.150048f
C2168 _023_ 0 0.345812f
C2169 _434_/a_2665_112# 0 0.62251f
C2174 _434_/a_36_151# 0 1.43589f
C2175 FILLER_0_5_136/a_36_472# 0 0.417394f
C2176 FILLER_0_5_136/a_124_375# 0 0.246306f
C2178 FILLER_0_18_209/a_36_472# 0 0.404746f
C2179 FILLER_0_18_209/a_572_375# 0 0.232991f
C2181 FILLER_0_12_28/a_36_472# 0 0.417394f
C2182 FILLER_0_12_28/a_124_375# 0 0.246306f
C2183 _040_ 0 0.355703f
C2189 _451_/a_36_151# 0 1.31409f
C2197 FILLER_0_6_47/a_36_472# 0 0.404746f
C2198 FILLER_0_6_47/a_3260_375# 0 0.233093f
C2206 FILLER_0_21_150/a_36_472# 0 0.417394f
C2207 FILLER_0_21_150/a_124_375# 0 0.246306f
C2209 FILLER_0_15_180/a_36_472# 0 0.404746f
C2210 FILLER_0_15_180/a_572_375# 0 0.232991f
C2219 FILLER_0_22_128/a_36_472# 0 0.404746f
C2220 FILLER_0_22_128/a_3260_375# 0 0.233093f
C2229 FILLER_0_19_111/a_36_472# 0 0.404746f
C2230 FILLER_0_19_111/a_572_375# 0 0.232991f
C2233 FILLER_0_19_155/a_36_472# 0 0.404746f
C2234 FILLER_0_19_155/a_572_375# 0 0.232991f
C2236 net11 0 1.328455f
C2237 net21 0 1.922829f
C2238 _007_ 0 0.309495f
C2239 net77 0 1.39077f
C2240 _418_/a_2665_112# 0 0.62251f
C2245 _418_/a_36_151# 0 1.43589f
C2248 FILLER_0_9_282/a_36_472# 0 0.404746f
C2249 FILLER_0_9_282/a_572_375# 0 0.232991f
C2254 FILLER_0_18_37/a_36_472# 0 0.404746f
C2255 FILLER_0_18_37/a_1468_375# 0 0.233029f
C2259 FILLER_0_2_127/a_36_472# 0 0.417394f
C2260 FILLER_0_2_127/a_124_375# 0 0.246306f
C2261 _157_ 0 0.531763f
C2262 _435_/a_2665_112# 0 0.62251f
C2267 _435_/a_36_151# 0 1.43589f
C2268 _108_ 0 0.411979f
C2269 trim_mask\[3\] 0 1.081535f
C2270 _164_ 0 1.3268f
C2271 _041_ 0 0.299289f
C2277 _452_/a_36_151# 0 1.31409f
C2278 FILLER_0_6_79/a_36_472# 0 0.417394f
C2279 FILLER_0_6_79/a_124_375# 0 0.246306f
C2280 net59 0 5.044369f
C2282 FILLER_0_15_59/a_36_472# 0 0.404746f
C2283 FILLER_0_15_59/a_572_375# 0 0.232991f
C2288 FILLER_0_3_221/a_36_472# 0 0.404746f
C2289 FILLER_0_3_221/a_1468_375# 0 0.233029f
C2294 FILLER_0_19_187/a_36_472# 0 0.404746f
C2295 FILLER_0_19_187/a_572_375# 0 0.232991f
C2300 FILLER_0_20_15/a_36_472# 0 0.404746f
C2301 FILLER_0_20_15/a_1468_375# 0 0.233029f
C2306 _419_/a_2665_112# 0 0.62251f
C2311 _419_/a_36_151# 0 1.43589f
C2312 _054_ 0 0.522819f
C2313 _221_/a_36_160# 0 0.386641f
C2315 FILLER_0_9_270/a_36_472# 0 0.404746f
C2316 FILLER_0_9_270/a_572_375# 0 0.232991f
C2318 FILLER_0_1_192/a_36_472# 0 0.417394f
C2319 FILLER_0_1_192/a_124_375# 0 0.246306f
C2320 FILLER_0_13_80/a_36_472# 0 0.417394f
C2321 FILLER_0_13_80/a_124_375# 0 0.246306f
C2322 _153_ 0 1.165862f
C2323 _154_ 0 1.167112f
C2324 _367_/a_36_68# 0 0.150048f
C2325 _436_/a_2665_112# 0 0.62251f
C2330 _436_/a_36_151# 0 1.43589f
C2332 FILLER_0_10_107/a_36_472# 0 0.404746f
C2333 FILLER_0_10_107/a_572_375# 0 0.232991f
C2335 _168_ 0 0.336537f
C2336 net51 0 2.105066f
C2337 _042_ 0 0.323587f
C2338 _453_/a_2665_112# 0 0.62251f
C2343 _453_/a_36_151# 0 1.43589f
C2344 FILLER_0_19_142/a_36_472# 0 0.417394f
C2345 FILLER_0_19_142/a_124_375# 0 0.246306f
C2346 _048_ 0 0.358805f
C2347 _205_/a_36_160# 0 0.696445f
C2348 net43 0 1.236377f
C2350 FILLER_0_3_78/a_36_472# 0 0.404746f
C2351 FILLER_0_3_78/a_572_375# 0 0.232991f
C2353 _437_/a_2665_112# 0 0.62251f
C2358 _437_/a_36_151# 0 1.43589f
C2359 _109_ 0 0.319326f
C2360 net37 0 1.529713f
C2362 FILLER_0_0_266/a_36_472# 0 0.417394f
C2363 FILLER_0_0_266/a_124_375# 0 0.246306f
C2364 net12 0 1.263595f
C2365 net22 0 2.108509f
C2366 FILLER_0_9_290/a_36_472# 0 0.417394f
C2367 FILLER_0_9_290/a_124_375# 0 0.246306f
C2368 _223_/a_36_160# 0 0.696445f
C2369 FILLER_0_14_263/a_36_472# 0 0.417394f
C2370 FILLER_0_14_263/a_124_375# 0 0.246306f
C2371 _158_ 0 0.309522f
C2372 _369_/a_36_68# 0 0.150048f
C2373 net71 0 1.420869f
C2374 _438_/a_2665_112# 0 0.62251f
C2379 _438_/a_36_151# 0 1.43589f
C2380 FILLER_0_23_274/a_36_472# 0 0.417394f
C2381 FILLER_0_23_274/a_124_375# 0 0.246306f
C2382 FILLER_0_17_282/a_36_472# 0 0.417394f
C2383 FILLER_0_17_282/a_124_375# 0 0.246306f
C2385 FILLER_0_5_198/a_36_472# 0 0.404746f
C2386 FILLER_0_5_198/a_572_375# 0 0.232991f
C2388 _163_ 0 1.03762f
C2389 _169_ 0 0.245383f
C2390 _386_/a_848_380# 0 0.40208f
C2393 FILLER_0_20_2/a_36_472# 0 0.404746f
C2394 FILLER_0_20_2/a_572_375# 0 0.232991f
C2399 FILLER_0_16_154/a_36_472# 0 0.404746f
C2400 FILLER_0_16_154/a_1468_375# 0 0.233029f
C2404 FILLER_0_0_232/a_36_472# 0 0.417394f
C2405 FILLER_0_0_232/a_124_375# 0 0.246306f
C2406 FILLER_0_19_195/a_36_472# 0 0.417394f
C2407 FILLER_0_19_195/a_124_375# 0 0.246306f
C2408 _049_ 0 0.329957f
C2409 net33 0 1.934915f
C2411 FILLER_0_3_54/a_36_472# 0 0.417394f
C2412 FILLER_0_3_54/a_124_375# 0 0.246306f
C2413 FILLER_0_2_101/a_36_472# 0 0.417394f
C2414 FILLER_0_2_101/a_124_375# 0 0.246306f
C2415 trim_mask\[0\] 0 0.605753f
C2416 _439_/a_2665_112# 0 0.62251f
C2421 _439_/a_36_151# 0 1.43589f
C2422 _066_ 0 0.333041f
C2426 FILLER_0_23_44/a_36_472# 0 0.404746f
C2427 FILLER_0_23_44/a_1468_375# 0 0.233029f
C2431 FILLER_0_23_88/a_36_472# 0 0.417394f
C2432 FILLER_0_23_88/a_124_375# 0 0.246306f
C2434 FILLER_0_5_164/a_36_472# 0 0.404746f
C2435 FILLER_0_5_164/a_572_375# 0 0.232991f
C2437 _060_ 0 2.485177f
C2438 _113_ 0 2.833205f
C2439 _090_ 0 2.629271f
C2440 _037_ 0 0.467089f
C2441 _170_ 0 0.413995f
C2442 _387_/a_36_113# 0 0.418095f
C2443 _208_/a_36_160# 0 0.696445f
C2445 FILLER_0_18_76/a_36_472# 0 0.404746f
C2446 FILLER_0_18_76/a_572_375# 0 0.232991f
C2448 _225_/a_36_160# 0 0.386641f
C2450 FILLER_0_2_177/a_36_472# 0 0.404746f
C2451 FILLER_0_2_177/a_572_375# 0 0.232991f
C2456 FILLER_0_2_111/a_36_472# 0 0.404746f
C2457 FILLER_0_2_111/a_1468_375# 0 0.233029f
C2461 FILLER_0_15_228/a_36_472# 0 0.417394f
C2462 FILLER_0_15_228/a_124_375# 0 0.246306f
C2463 net47 0 2.314376f
C2464 _242_/a_36_160# 0 0.696445f
C2465 _117_ 0 1.266251f
C2467 _043_ 0 0.487279f
C2468 _190_/a_36_160# 0 0.696445f
C2470 FILLER_0_9_105/a_36_472# 0 0.404746f
C2471 FILLER_0_9_105/a_572_375# 0 0.232991f
C2473 FILLER_0_13_100/a_36_472# 0 0.417394f
C2474 FILLER_0_13_100/a_124_375# 0 0.246306f
C2478 FILLER_0_22_177/a_36_472# 0 0.404746f
C2479 FILLER_0_22_177/a_1468_375# 0 0.233029f
C2484 FILLER_0_15_2/a_36_472# 0 0.404746f
C2485 FILLER_0_15_2/a_572_375# 0 0.232991f
C2487 FILLER_0_15_10/a_36_472# 0 0.417394f
C2488 FILLER_0_15_10/a_124_375# 0 0.246306f
C2492 FILLER_0_19_171/a_36_472# 0 0.404746f
C2493 FILLER_0_19_171/a_1468_375# 0 0.233029f
C2497 net13 0 1.176306f
C2498 net23 0 2.091399f
C2499 FILLER_0_20_87/a_36_472# 0 0.417394f
C2500 FILLER_0_20_87/a_124_375# 0 0.246306f
C2501 FILLER_0_20_98/a_36_472# 0 0.417394f
C2502 FILLER_0_20_98/a_124_375# 0 0.246306f
C2503 _055_ 0 1.782885f
C2505 FILLER_0_18_53/a_36_472# 0 0.404746f
C2506 FILLER_0_18_53/a_572_375# 0 0.232991f
C2508 FILLER_0_2_165/a_36_472# 0 0.417394f
C2509 FILLER_0_2_165/a_124_375# 0 0.246306f
C2510 FILLER_0_15_205/a_36_472# 0 0.417394f
C2511 FILLER_0_15_205/a_124_375# 0 0.246306f
C2513 FILLER_0_23_282/a_36_472# 0 0.404746f
C2514 FILLER_0_23_282/a_572_375# 0 0.232991f
C2516 net42 0 1.067446f
C2517 net17 0 2.210219f
C2518 _172_ 0 0.265782f
C2519 _171_ 0 0.300355f
C2521 _080_ 0 0.328202f
C2523 FILLER_0_0_96/a_36_472# 0 0.417394f
C2524 FILLER_0_0_96/a_124_375# 0 0.246306f
C2528 FILLER_0_9_72/a_36_472# 0 0.404746f
C2529 FILLER_0_9_72/a_1468_375# 0 0.233029f
C2533 FILLER_0_20_31/a_36_472# 0 0.417394f
C2534 FILLER_0_20_31/a_124_375# 0 0.246306f
C2535 _227_/a_36_160# 0 0.386641f
C2536 _120_ 0 1.533088f
C2538 FILLER_0_5_172/a_36_472# 0 0.417394f
C2539 FILLER_0_5_172/a_124_375# 0 0.246306f
C2541 FILLER_0_12_20/a_36_472# 0 0.404746f
C2542 FILLER_0_12_20/a_572_375# 0 0.232991f
C2544 _134_ 0 0.365972f
C2545 _062_ 0 1.717773f
C2546 _059_ 0 1.686761f
C2547 _261_/a_36_160# 0 0.386641f
C2548 _044_ 0 0.388801f
C2549 mask\[1\] 0 1.295078f
C2554 FILLER_0_13_142/a_36_472# 0 0.404746f
C2555 FILLER_0_13_142/a_1468_375# 0 0.233029f
C2560 FILLER_0_9_60/a_36_472# 0 0.404746f
C2561 FILLER_0_9_60/a_572_375# 0 0.232991f
C2563 FILLER_0_7_233/a_36_472# 0 0.417394f
C2564 FILLER_0_7_233/a_124_375# 0 0.246306f
C2565 _228_/a_36_68# 0 0.69549f
C2566 FILLER_0_21_206/a_36_472# 0 0.417394f
C2567 FILLER_0_21_206/a_124_375# 0 0.246306f
C2568 _067_ 0 0.851951f
C2569 _135_ 0 0.339478f
C2570 _193_/a_36_160# 0 0.696445f
C2571 _180_ 0 0.390598f
C2572 cal_count\[1\] 0 1.568289f
C2574 FILLER_0_4_213/a_36_472# 0 0.404746f
C2575 FILLER_0_4_213/a_572_375# 0 0.232991f
C2577 FILLER_0_11_282/a_36_472# 0 0.417394f
C2578 FILLER_0_11_282/a_124_375# 0 0.246306f
C2579 FILLER_0_18_61/a_36_472# 0 0.417394f
C2580 FILLER_0_18_61/a_124_375# 0 0.246306f
C2582 FILLER_0_15_235/a_36_472# 0 0.404746f
C2583 FILLER_0_15_235/a_572_375# 0 0.232991f
C2585 FILLER_0_23_290/a_36_472# 0 0.417394f
C2586 FILLER_0_23_290/a_124_375# 0 0.246306f
C2587 _121_ 0 0.532847f
C2588 _246_/a_36_68# 0 0.69549f
C2589 FILLER_0_5_181/a_36_472# 0 0.417394f
C2590 FILLER_0_5_181/a_124_375# 0 0.246306f
C2591 _082_ 0 0.619901f
C2592 net8 0 1.163723f
C2593 net18 0 2.032159f
C2594 _179_ 0 0.336984f
C2599 FILLER_0_14_107/a_36_472# 0 0.404746f
C2600 FILLER_0_14_107/a_1468_375# 0 0.233029f
C2604 _097_ 0 0.592554f
C2605 FILLER_0_1_204/a_36_472# 0 0.417394f
C2606 FILLER_0_1_204/a_124_375# 0 0.246306f
C2608 FILLER_0_15_72/a_36_472# 0 0.404746f
C2609 FILLER_0_15_72/a_572_375# 0 0.232991f
C2614 FILLER_0_17_104/a_36_472# 0 0.404746f
C2615 FILLER_0_17_104/a_1468_375# 0 0.233029f
C2620 FILLER_0_8_37/a_36_472# 0 0.404746f
C2621 FILLER_0_8_37/a_572_375# 0 0.232991f
C2626 FILLER_0_15_212/a_36_472# 0 0.404746f
C2627 FILLER_0_15_212/a_1468_375# 0 0.233029f
C2631 FILLER_0_23_60/a_36_472# 0 0.417394f
C2632 FILLER_0_23_60/a_124_375# 0 0.246306f
C2633 _123_ 0 0.344874f
C2634 _122_ 0 0.600118f
C2635 calibrate 0 1.343796f
C2636 _316_/a_848_380# 0 0.40208f
C2638 _247_/a_36_160# 0 0.696445f
C2639 FILLER_0_12_50/a_36_472# 0 0.417394f
C2640 FILLER_0_12_50/a_124_375# 0 0.246306f
C2641 _084_ 0 0.296163f
C2642 cal_itt\[0\] 0 1.831055f
C2643 cal_itt\[1\] 0 1.705665f
C2644 FILLER_0_11_109/a_36_472# 0 0.417394f
C2645 FILLER_0_11_109/a_124_375# 0 0.246306f
C2646 _182_ 0 0.34197f
C2650 _045_ 0 0.349338f
C2651 mask\[2\] 0 1.335688f
C2653 _333_/a_36_160# 0 0.386641f
C2654 _098_ 0 1.816151f
C2655 _147_ 0 0.322539f
C2657 FILLER_0_12_236/a_36_472# 0 0.404746f
C2658 FILLER_0_12_236/a_572_375# 0 0.232991f
C2660 FILLER_0_2_171/a_36_472# 0 0.417394f
C2661 FILLER_0_2_171/a_124_375# 0 0.246306f
C2662 _014_ 0 0.363432f
C2663 _317_/a_36_113# 0 0.418095f
C2664 _248_/a_36_68# 0 0.69549f
C2666 FILLER_0_17_38/a_36_472# 0 0.404746f
C2667 FILLER_0_17_38/a_572_375# 0 0.232991f
C2669 _001_ 0 0.285216f
C2671 _196_/a_36_160# 0 0.696445f
C2673 FILLER_0_6_90/a_36_472# 0 0.404746f
C2674 FILLER_0_6_90/a_572_375# 0 0.232991f
C2676 _183_ 0 0.356629f
C2677 _334_/a_36_160# 0 0.386641f
C2678 _282_/a_36_160# 0 0.386641f
C2679 _024_ 0 0.451815f
C2680 _009_ 0 0.397943f
C2681 _420_/a_2665_112# 0 0.62251f
C2686 _420_/a_36_151# 0 1.43589f
C2687 clk 0 1.162312f
C2688 FILLER_0_8_2/a_36_472# 0 0.417394f
C2689 FILLER_0_8_2/a_124_375# 0 0.246306f
C2691 FILLER_0_8_24/a_36_472# 0 0.404746f
C2692 FILLER_0_8_24/a_572_375# 0 0.232991f
C2694 _124_ 0 0.294081f
C2695 _118_ 0 1.378735f
C2696 _071_ 0 1.600488f
C2697 net9 0 1.13171f
C2698 net19 0 1.889339f
C2699 _138_ 0 0.33132f
C2700 _137_ 0 1.178616f
C2701 FILLER_0_20_107/a_36_472# 0 0.417394f
C2702 FILLER_0_20_107/a_124_375# 0 0.246306f
C2703 FILLER_0_9_142/a_36_472# 0 0.417394f
C2704 FILLER_0_9_142/a_124_375# 0 0.246306f
C2705 _099_ 0 1.152785f
C2706 mask\[7\] 0 1.477838f
C2707 _010_ 0 0.377779f
C2708 _421_/a_2665_112# 0 0.62251f
C2713 _421_/a_36_151# 0 1.43589f
C2714 FILLER_0_1_212/a_36_472# 0 0.417394f
C2715 FILLER_0_1_212/a_124_375# 0 0.246306f
C2716 FILLER_0_8_239/a_36_472# 0 0.417394f
C2717 FILLER_0_8_239/a_124_375# 0 0.246306f
C2718 _125_ 0 1.526603f
C2719 _058_ 0 1.483584f
C2721 FILLER_0_6_177/a_36_472# 0 0.404746f
C2722 FILLER_0_6_177/a_572_375# 0 0.232991f
C2724 state\[1\] 0 2.652405f
C2726 _184_ 0 0.350066f
C2727 cal_count\[2\] 0 1.971854f
C2729 _018_ 0 0.358633f
C2730 _046_ 0 0.361963f
C2732 _094_ 0 1.263877f
C2733 _100_ 0 0.333135f
C2734 net36 0 2.262756f
C2735 FILLER_0_17_133/a_36_472# 0 0.417394f
C2736 FILLER_0_17_133/a_124_375# 0 0.246306f
C2737 _025_ 0 0.350324f
C2738 _148_ 0 0.325709f
C2739 _422_/a_2665_112# 0 0.62251f
C2744 _422_/a_36_151# 0 1.43589f
C2746 FILLER_0_1_266/a_36_472# 0 0.404746f
C2747 FILLER_0_1_266/a_572_375# 0 0.232991f
C2749 _152_ 0 0.918583f
C2750 _081_ 0 1.140656f
C2751 _370_/a_848_380# 0 0.40208f
C2756 FILLER_0_24_274/a_36_472# 0 0.404746f
C2757 FILLER_0_24_274/a_1468_375# 0 0.233029f
C2761 _185_ 0 0.386917f
C2763 _199_/a_36_160# 0 0.696445f
C2764 _012_ 0 0.75195f
C2765 _423_/a_2665_112# 0 0.62251f
C2770 _423_/a_36_151# 0 1.43589f
C2771 FILLER_0_5_88/a_36_472# 0 0.417394f
C2772 FILLER_0_5_88/a_124_375# 0 0.246306f
C2773 trim_mask\[1\] 0 1.020743f
C2774 _029_ 0 0.308904f
C2775 _440_/a_2665_112# 0 0.62251f
C2780 _440_/a_36_151# 0 1.43589f
C2781 _159_ 0 0.351814f
C2782 _371_/a_36_113# 0 0.418095f
C2784 FILLER_0_17_56/a_36_472# 0 0.404746f
C2785 FILLER_0_17_56/a_572_375# 0 0.232991f
C2787 _083_ 0 0.527882f
C2788 _078_ 0 0.904554f
C2789 _181_ 0 0.829168f
C2790 _019_ 0 0.32907f
C2791 _139_ 0 0.346404f
C2792 FILLER_0_14_123/a_36_472# 0 0.417394f
C2793 FILLER_0_14_123/a_124_375# 0 0.246306f
C2794 _005_ 0 0.340993f
C2795 _101_ 0 0.280497f
C2796 _424_/a_2665_112# 0 0.62251f
C2801 _424_/a_36_151# 0 1.43589f
C2802 _026_ 0 0.320379f
C2803 _149_ 0 0.305496f
C2807 FILLER_0_5_54/a_36_472# 0 0.404746f
C2808 FILLER_0_5_54/a_1468_375# 0 0.233029f
C2813 FILLER_0_17_142/a_36_472# 0 0.404746f
C2814 FILLER_0_17_142/a_572_375# 0 0.232991f
C2816 _068_ 0 3.162692f
C2817 _076_ 0 3.812442f
C2818 _133_ 0 1.430901f
C2819 _070_ 0 3.115722f
C2820 net49 0 5.140563f
C2821 _030_ 0 0.307083f
C2822 net66 0 1.472669f
C2823 _441_/a_2665_112# 0 0.62251f
C2828 _441_/a_36_151# 0 1.43589f
C2829 FILLER_0_5_206/a_36_472# 0 0.417394f
C2830 FILLER_0_5_206/a_124_375# 0 0.246306f
C2831 fanout49/a_36_160# 0 0.696445f
C2835 FILLER_0_8_247/a_36_472# 0 0.404746f
C2836 FILLER_0_8_247/a_1468_375# 0 0.233029f
C2843 FILLER_0_12_220/a_36_472# 0 0.404746f
C2844 FILLER_0_12_220/a_1468_375# 0 0.233029f
C2849 FILLER_0_21_286/a_36_472# 0 0.404746f
C2850 FILLER_0_21_286/a_572_375# 0 0.232991f
C2852 _140_ 0 1.276518f
C2853 _339_/a_36_160# 0 0.386641f
C2854 _095_ 0 2.689027f
C2855 _186_ 0 0.580923f
C2859 FILLER_0_20_169/a_36_472# 0 0.417394f
C2860 FILLER_0_20_169/a_124_375# 0 0.246306f
C2862 _425_/a_2665_112# 0 0.62251f
C2867 _425_/a_36_151# 0 1.43589f
C2868 net5 0 0.610761f
C2869 input5/a_36_113# 0 0.418095f
C2871 FILLER_0_11_78/a_36_472# 0 0.404746f
C2872 FILLER_0_11_78/a_572_375# 0 0.232991f
C2874 _102_ 0 0.335308f
C2875 mask\[9\] 0 1.383606f
C2876 _031_ 0 0.417351f
C2877 net69 0 1.020293f
C2878 _442_/a_2665_112# 0 0.62251f
C2883 _442_/a_36_151# 0 1.43589f
C2884 net64 0 2.598514f
C2885 fanout59/a_36_160# 0 0.696445f
C2886 FILLER_0_14_99/a_36_472# 0 0.417394f
C2887 FILLER_0_14_99/a_124_375# 0 0.246306f
C2888 _038_ 0 0.362839f
C2889 _136_ 0 1.345638f
C2890 _390_/a_36_68# 0 0.150048f
C2892 FILLER_0_15_282/a_36_472# 0 0.404746f
C2893 FILLER_0_15_282/a_572_375# 0 0.232991f
C2895 FILLER_0_11_124/a_36_472# 0 0.417394f
C2896 FILLER_0_11_124/a_124_375# 0 0.246306f
C2897 FILLER_0_11_135/a_36_472# 0 0.417394f
C2898 FILLER_0_11_135/a_124_375# 0 0.246306f
C2899 _188_ 0 0.349407f
C2900 cal_count\[3\] 0 1.862896f
C2901 _050_ 0 0.622354f
C2902 _211_/a_36_160# 0 0.386641f
C2903 net4 0 2.711508f
C2904 en 0 0.833743f
C2905 input4/a_36_68# 0 0.69549f
C2906 _426_/a_2665_112# 0 0.62251f
C2911 _426_/a_36_151# 0 1.43589f
C2912 _027_ 0 0.302949f
C2913 _150_ 0 0.320497f
C2921 FILLER_0_18_107/a_36_472# 0 0.404746f
C2922 FILLER_0_18_107/a_3260_375# 0 0.233093f
C2930 trim_mask\[4\] 0 0.987791f
C2931 _032_ 0 0.34876f
C2932 _443_/a_2665_112# 0 0.62251f
C2937 _443_/a_36_151# 0 1.43589f
C2938 _061_ 0 0.84986f
C2939 _056_ 0 2.393362f
C2941 fanout58/a_36_160# 0 0.696445f
C2942 net74 0 1.237373f
C2943 fanout69/a_36_113# 0 0.418095f
C2944 _173_ 0 0.339446f
C2945 FILLER_0_3_142/a_36_472# 0 0.417394f
C2946 FILLER_0_3_142/a_124_375# 0 0.246306f
C2947 FILLER_0_17_64/a_36_472# 0 0.417394f
C2948 FILLER_0_17_64/a_124_375# 0 0.246306f
C2950 FILLER_0_11_101/a_36_472# 0 0.404746f
C2951 FILLER_0_11_101/a_572_375# 0 0.232991f
C2956 FILLER_0_22_86/a_36_472# 0 0.404746f
C2957 FILLER_0_22_86/a_1468_375# 0 0.233029f
C2961 net24 0 1.61895f
C2962 net3 0 0.740676f
C2963 input3/a_36_113# 0 0.418095f
C2964 _103_ 0 0.350464f
C2965 _151_ 0 0.300777f
C2971 _427_/a_36_151# 0 1.43587f
C2972 FILLER_0_17_161/a_36_472# 0 0.417394f
C2973 FILLER_0_17_161/a_124_375# 0 0.246306f
C2977 FILLER_0_18_139/a_36_472# 0 0.404746f
C2978 FILLER_0_18_139/a_1468_375# 0 0.233029f
C2982 _161_ 0 0.592909f
C2983 _162_ 0 0.597238f
C2984 trim_val\[0\] 0 0.742779f
C2985 net67 0 1.662327f
C2986 _444_/a_2665_112# 0 0.62251f
C2991 _444_/a_36_151# 0 1.43589f
C2992 net65 0 0.804072f
C2993 fanout57/a_36_113# 0 0.418095f
C2994 fanout68/a_36_113# 0 0.418095f
C2996 FILLER_0_12_2/a_36_472# 0 0.404746f
C2997 FILLER_0_12_2/a_572_375# 0 0.232991f
C2999 net79 0 1.584979f
C3000 fanout79/a_36_160# 0 0.386641f
C3002 FILLER_0_13_228/a_36_472# 0 0.417394f
C3003 FILLER_0_13_228/a_124_375# 0 0.246306f
C3004 FILLER_0_13_206/a_36_472# 0 0.417394f
C3005 FILLER_0_13_206/a_124_375# 0 0.246306f
C3009 FILLER_0_20_177/a_36_472# 0 0.404746f
C3010 FILLER_0_20_177/a_1468_375# 0 0.233029f
C3014 _051_ 0 0.349381f
C3016 net2 0 0.461658f
C3017 input2/a_36_113# 0 0.418095f
C3018 _129_ 0 0.926508f
C3019 _131_ 0 1.734297f
C3021 FILLER_0_11_64/a_36_472# 0 0.417394f
C3022 FILLER_0_11_64/a_124_375# 0 0.246306f
C3023 state\[2\] 0 0.607433f
C3024 net53 0 4.483899f
C3025 _017_ 0 0.334329f
C3026 net70 0 1.238296f
C3027 _428_/a_2665_112# 0 0.62251f
C3032 _428_/a_36_151# 0 1.43589f
C3036 FILLER_0_5_72/a_36_472# 0 0.404746f
C3037 FILLER_0_5_72/a_1468_375# 0 0.233029f
C3041 _376_/a_36_160# 0 0.386641f
C3042 trim_val\[1\] 0 0.683578f
C3043 _445_/a_2665_112# 0 0.62251f
C3048 _445_/a_36_151# 0 1.43589f
C3049 fanout67/a_36_160# 0 0.386641f
C3050 fanout56/a_36_113# 0 0.418095f
C3051 net78 0 0.686263f
C3052 fanout78/a_36_113# 0 0.418095f
C3053 _174_ 0 0.979741f
C3054 FILLER_0_0_198/a_36_472# 0 0.417394f
C3055 FILLER_0_0_198/a_124_375# 0 0.246306f
C3056 FILLER_0_15_290/a_36_472# 0 0.417394f
C3057 FILLER_0_15_290/a_124_375# 0 0.246306f
C3058 FILLER_0_24_290/a_36_472# 0 0.417394f
C3059 FILLER_0_24_290/a_124_375# 0 0.246306f
C3063 FILLER_0_4_107/a_36_472# 0 0.404746f
C3064 FILLER_0_4_107/a_1468_375# 0 0.233029f
C3071 FILLER_0_7_104/a_36_472# 0 0.404746f
C3072 FILLER_0_7_104/a_1468_375# 0 0.233029f
C3076 _214_/a_36_160# 0 0.386641f
C3077 net1 0 0.364811f
C3078 input1/a_36_113# 0 0.418095f
C3079 _429_/a_2665_112# 0 0.62251f
C3084 _429_/a_36_151# 0 1.43589f
C3085 _011_ 0 0.278979f
C3086 fanout66/a_36_113# 0 0.418095f
C3087 _035_ 0 0.327801f
C3088 _446_/a_2665_112# 0 0.62251f
C3093 _446_/a_36_151# 0 1.43589f
C3094 fanout77/a_36_113# 0 0.418095f
C3095 FILLER_0_5_212/a_36_472# 0 0.417394f
C3096 FILLER_0_5_212/a_124_375# 0 0.246306f
C3097 fanout55/a_36_160# 0 0.696445f
C3098 _175_ 0 0.344159f
C3109 FILLER_0_3_172/a_36_472# 0 0.404746f
C3110 FILLER_0_3_172/a_3260_375# 0 0.233093f
C3125 FILLER_0_17_72/a_36_472# 0 0.404746f
C3126 FILLER_0_17_72/a_3260_375# 0 0.233093f
C3135 FILLER_0_2_93/a_36_472# 0 0.404746f
C3136 FILLER_0_2_93/a_572_375# 0 0.232991f
C3139 FILLER_0_11_142/a_36_472# 0 0.404746f
C3140 FILLER_0_11_142/a_572_375# 0 0.232991f
C3142 net25 0 1.803174f
C3144 net35 0 1.844415f
C3145 mask\[8\] 0 1.276111f
C3146 _033_ 0 0.323682f
C3147 _165_ 0 0.331995f
C3148 FILLER_0_3_2/a_36_472# 0 0.417394f
C3149 FILLER_0_3_2/a_124_375# 0 0.246306f
C3150 trim_val\[3\] 0 0.719615f
C3151 _036_ 0 0.369206f
C3152 net68 0 1.735004f
C3153 _447_/a_2665_112# 0 0.62251f
C3158 _447_/a_36_151# 0 1.43589f
C3160 FILLER_0_19_28/a_36_472# 0 0.404746f
C3161 FILLER_0_19_28/a_572_375# 0 0.232991f
C3163 fanout65/a_36_113# 0 0.418095f
C3164 fanout76/a_36_160# 0 0.386641f
C3165 net54 0 5.456963f
C3166 fanout54/a_36_160# 0 0.696445f
C3168 FILLER_0_4_49/a_36_472# 0 0.404746f
C3169 FILLER_0_4_49/a_572_375# 0 0.232991f
C3171 _176_ 0 0.804011f
C3172 _085_ 0 2.280803f
C3173 _116_ 0 1.959915f
C3175 FILLER_0_14_50/a_36_472# 0 0.417394f
C3176 FILLER_0_14_50/a_124_375# 0 0.246306f
C3177 FILLER_0_8_263/a_36_472# 0 0.417394f
C3178 FILLER_0_8_263/a_124_375# 0 0.246306f
C3179 FILLER_0_0_130/a_36_472# 0 0.417394f
C3180 FILLER_0_0_130/a_124_375# 0 0.246306f
C3181 FILLER_0_16_255/a_36_472# 0 0.417394f
C3182 FILLER_0_16_255/a_124_375# 0 0.246306f
C3184 FILLER_0_7_59/a_36_472# 0 0.404746f
C3185 FILLER_0_7_59/a_572_375# 0 0.232991f
C3187 ctlp[2] 0 0.17528f
C3188 output19/a_224_472# 0 2.38465f
C3189 FILLER_0_7_146/a_36_472# 0 0.417394f
C3190 FILLER_0_7_146/a_124_375# 0 0.246306f
C3193 FILLER_0_15_116/a_36_472# 0 0.404746f
C3194 FILLER_0_15_116/a_572_375# 0 0.232991f
C3196 _063_ 0 0.370155f
C3197 _233_/a_36_160# 0 0.386641f
C3205 FILLER_0_21_28/a_36_472# 0 0.404746f
C3206 FILLER_0_21_28/a_3260_375# 0 0.233093f
C3214 _110_ 0 0.323912f
C3215 trim_val\[4\] 0 0.662409f
C3216 net76 0 1.454269f
C3217 _448_/a_2665_112# 0 0.62251f
C3222 _448_/a_36_151# 0 1.43589f
C3223 fanout64/a_36_160# 0 0.386641f
C3224 fanout75/a_36_113# 0 0.418095f
C3225 _250_/a_36_68# 0 0.69549f
C3226 net56 0 0.843396f
C3227 fanout53/a_36_160# 0 0.696445f
C3228 _177_ 0 0.358286f
C3229 result[2] 0 0.230851f
C3230 net29 0 1.802718f
C3231 output29/a_224_472# 0 2.38465f
C3232 ctlp[1] 0 0.17418f
C3233 output18/a_224_472# 0 2.38465f
C3234 FILLER_0_14_181/a_36_472# 0 0.417394f
C3235 FILLER_0_14_181/a_124_375# 0 0.246306f
C3236 _052_ 0 0.569133f
C3237 _217_/a_36_160# 0 0.386641f
C3238 net44 0 1.407054f
C3239 en_co_clk 0 0.346872f
C3240 net55 0 5.119958f
C3241 net72 0 1.366255f
C3242 _449_/a_2665_112# 0 0.62251f
C3247 _449_/a_36_151# 0 1.43589f
C3248 fanout52/a_36_160# 0 0.696445f
C3249 net82 0 0.706042f
C3250 fanout74/a_36_113# 0 0.418095f
C3251 FILLER_0_10_28/a_36_472# 0 0.417394f
C3252 FILLER_0_10_28/a_124_375# 0 0.246306f
C3253 mask\[0\] 0 2.242948f
C3255 fanout63/a_36_160# 0 0.696445f
C3256 FILLER_0_14_81/a_36_472# 0 0.417394f
C3257 FILLER_0_14_81/a_124_375# 0 0.246306f
C3261 FILLER_0_13_212/a_36_472# 0 0.404746f
C3262 FILLER_0_13_212/a_1468_375# 0 0.233029f
C3266 trim[1] 0 0.793787f
C3267 net39 0 1.445128f
C3268 output39/a_224_472# 0 2.38465f
C3269 result[1] 0 0.229507f
C3270 net28 0 1.759728f
C3271 output28/a_224_472# 0 2.38465f
C3272 ctlp[0] 0 1.002286f
C3273 output17/a_224_472# 0 2.38465f
C3274 FILLER_0_16_37/a_36_472# 0 0.417394f
C3275 FILLER_0_16_37/a_124_375# 0 0.246306f
C3276 net26 0 1.671545f
C3277 _064_ 0 0.581481f
C3278 trim_val\[2\] 0 0.65354f
C3279 trim_mask\[2\] 0 0.92551f
C3281 _013_ 0 0.48783f
C3282 _111_ 0 0.369652f
C3290 FILLER_0_18_177/a_36_472# 0 0.404746f
C3291 FILLER_0_18_177/a_3260_375# 0 0.233093f
C3299 FILLER_0_18_100/a_36_472# 0 0.417394f
C3300 FILLER_0_18_100/a_124_375# 0 0.246306f
C3301 _073_ 0 0.953711f
C3302 _126_ 0 2.036767f
C3303 _069_ 0 2.034557f
C3304 fanout51/a_36_113# 0 0.418095f
C3305 fanout62/a_36_160# 0 0.696445f
C3306 fanout73/a_36_113# 0 0.418095f
C3308 FILLER_0_19_47/a_36_472# 0 0.404746f
C3309 FILLER_0_19_47/a_572_375# 0 0.232991f
C3312 FILLER_0_14_91/a_36_472# 0 0.404746f
C3313 FILLER_0_14_91/a_572_375# 0 0.232991f
C3315 FILLER_0_10_214/a_36_472# 0 0.417394f
C3316 FILLER_0_10_214/a_124_375# 0 0.246306f
C3317 FILLER_0_10_247/a_36_472# 0 0.417394f
C3318 FILLER_0_10_247/a_124_375# 0 0.246306f
C3319 _178_ 0 1.252435f
C3320 _398_/a_36_113# 0 0.418095f
C3321 FILLER_0_16_241/a_36_472# 0 0.417394f
C3322 FILLER_0_16_241/a_124_375# 0 0.246306f
C3323 trim[0] 0 0.796081f
C3324 net38 0 1.529392f
C3325 output38/a_224_472# 0 2.38465f
C3326 ctln[9] 0 0.904836f
C3327 net16 0 1.295744f
C3328 output16/a_224_472# 0 2.38465f
C3329 result[0] 0 0.56622f
C3330 net27 0 2.023744f
C3331 output27/a_224_472# 0 2.38465f
C3332 _219_/a_36_160# 0 0.386641f
C3334 FILLER_0_20_193/a_36_472# 0 0.404746f
C3335 FILLER_0_20_193/a_572_375# 0 0.232991f
C3337 _236_/a_36_160# 0 0.696445f
C3338 _112_ 0 0.308886f
C3340 _074_ 0 1.813232f
C3341 net50 0 4.486121f
C3342 net52 0 3.536016f
C3343 fanout50/a_36_160# 0 0.696445f
C3344 FILLER_0_10_37/a_36_472# 0 0.417394f
C3345 FILLER_0_10_37/a_124_375# 0 0.246306f
C3346 fanout72/a_36_113# 0 0.418095f
C3347 fanout61/a_36_113# 0 0.418095f
C3348 _128_ 0 0.447252f
C3349 _127_ 0 1.291729f
C3350 _322_/a_848_380# 0 0.40208f
C3352 _088_ 0 0.457961f
C3353 _079_ 0 1.114894f
C3354 _087_ 0 0.601674f
C3355 FILLER_0_4_123/a_36_472# 0 0.417394f
C3356 FILLER_0_4_123/a_124_375# 0 0.246306f
C3358 FILLER_0_17_218/a_36_472# 0 0.404746f
C3359 FILLER_0_17_218/a_572_375# 0 0.232991f
C3361 sample 0 0.508149f
C3362 output37/a_224_472# 0 2.38465f
C3363 valid 0 0.272072f
C3364 net48 0 1.219262f
C3365 output48/a_224_472# 0 2.38465f
C3366 ctln[8] 0 1.547984f
C3367 net15 0 1.440851f
C3368 output15/a_224_472# 0 2.38465f
C3369 ctlp[9] 0 0.73349f
C3370 output26/a_224_472# 0 2.38465f
C3374 FILLER_0_16_57/a_36_472# 0 0.404746f
C3375 FILLER_0_16_57/a_1468_375# 0 0.233029f
C3379 _306_/a_36_68# 0 0.69549f
C3380 _072_ 0 2.604301f
C3381 fanout82/a_36_113# 0 0.418095f
C3382 _015_ 0 0.406653f
C3383 _323_/a_36_113# 0 0.418095f
C3384 net60 0 5.024503f
C3385 net61 0 1.666523f
C3386 fanout60/a_36_160# 0 0.696445f
C3387 fanout71/a_36_113# 0 0.418095f
C3388 FILLER_0_6_239/a_36_472# 0 0.417394f
C3389 FILLER_0_6_239/a_124_375# 0 0.246306f
C3390 FILLER_0_4_99/a_36_472# 0 0.417394f
C3391 FILLER_0_4_99/a_124_375# 0 0.246306f
C3392 net57 0 1.383718f
C3393 FILLER_0_10_256/a_36_472# 0 0.417394f
C3394 FILLER_0_10_256/a_124_375# 0 0.246306f
C3395 cal_itt\[3\] 0 1.854962f
C3396 _340_/a_36_160# 0 0.386641f
C3398 FILLER_0_4_177/a_36_472# 0 0.404746f
C3399 FILLER_0_4_177/a_572_375# 0 0.232991f
C3402 FILLER_0_4_144/a_36_472# 0 0.404746f
C3403 FILLER_0_4_144/a_572_375# 0 0.232991f
C3405 ctln[7] 0 1.265946f
C3406 output14/a_224_472# 0 2.38465f
C3407 result[9] 0 0.8197f
C3408 output36/a_224_472# 0 2.38465f
C3409 trimb[4] 0 0.752332f
C3410 output47/a_224_472# 0 2.38465f
C3411 ctlp[8] 0 1.136333f
C3412 output25/a_224_472# 0 2.38465f
C3416 FILLER_0_12_136/a_36_472# 0 0.404746f
C3417 FILLER_0_12_136/a_1468_375# 0 0.233029f
C3424 FILLER_0_16_89/a_36_472# 0 0.404746f
C3425 FILLER_0_16_89/a_1468_375# 0 0.233029f
C3430 FILLER_0_21_125/a_36_472# 0 0.404746f
C3431 FILLER_0_21_125/a_572_375# 0 0.232991f
C3434 _096_ 0 2.205532f
C3435 _093_ 0 1.893313f
C3436 FILLER_0_19_55/a_36_472# 0 0.417394f
C3437 FILLER_0_19_55/a_124_375# 0 0.246306f
C3438 net81 0 1.738987f
C3439 fanout81/a_36_160# 0 0.386641f
C3440 _057_ 0 1.600886f
C3442 net73 0 1.058857f
C3443 fanout70/a_36_113# 0 0.418095f
C3444 _003_ 0 0.3064f
C3445 _089_ 0 0.36777f
C3446 _187_ 0 0.311229f
C3448 _141_ 0 1.249289f
C3449 mask\[3\] 0 1.26722f
C3450 cal 0 0.793393f
C3451 FILLER_0_7_195/a_36_472# 0 0.417394f
C3452 FILLER_0_7_195/a_124_375# 0 0.246306f
C3453 FILLER_0_7_162/a_36_472# 0 0.417394f
C3454 FILLER_0_7_162/a_124_375# 0 0.246306f
C3455 ctln[6] 0 1.451644f
C3456 output13/a_224_472# 0 2.38465f
C3464 FILLER_0_18_2/a_36_472# 0 0.404746f
C3465 FILLER_0_18_2/a_3260_375# 0 0.233093f
C3473 trimb[3] 0 0.34698f
C3474 net46 0 1.13395f
C3475 output46/a_224_472# 0 2.38465f
C3476 result[8] 0 0.68837f
C3477 output35/a_224_472# 0 2.38465f
C3478 ctlp[7] 0 0.83567f
C3479 output24/a_224_472# 0 2.38465f
C3480 FILLER_0_8_107/a_36_472# 0 0.417394f
C3481 FILLER_0_8_107/a_124_375# 0 0.246306f
C3482 FILLER_0_12_124/a_36_472# 0 0.417394f
C3483 FILLER_0_12_124/a_124_375# 0 0.246306f
C3484 net41 0 1.746759f
C3485 _065_ 0 0.523724f
C3486 _239_/a_36_160# 0 0.696445f
C3487 FILLER_0_1_98/a_36_472# 0 0.417394f
C3488 FILLER_0_1_98/a_124_375# 0 0.246306f
C3489 _115_ 0 1.281516f
C3490 _114_ 0 2.293579f
C3491 _308_/a_848_380# 0 0.40208f
C3496 FILLER_0_10_78/a_36_472# 0 0.404746f
C3497 FILLER_0_10_78/a_1468_375# 0 0.233029f
C3501 _130_ 0 0.304085f
C3502 net80 0 1.375599f
C3503 fanout80/a_36_113# 0 0.418095f
C3504 net58 0 5.308423f
C3505 _000_ 0 0.382358f
C3506 net75 0 1.474299f
C3507 _411_/a_2665_112# 0 0.62251f
C3512 _411_/a_36_151# 0 1.43589f
C3513 state\[0\] 0 0.680109f
C3514 _273_/a_36_68# 0 0.69549f
C3515 _142_ 0 0.324372f
C3517 FILLER_0_9_223/a_36_472# 0 0.404746f
C3518 FILLER_0_9_223/a_572_375# 0 0.232991f
C3523 FILLER_0_4_197/a_36_472# 0 0.404746f
C3524 FILLER_0_4_197/a_1468_375# 0 0.233029f
C3528 FILLER_0_17_226/a_36_472# 0 0.417394f
C3529 FILLER_0_17_226/a_124_375# 0 0.246306f
C3531 FILLER_0_5_109/a_36_472# 0 0.404746f
C3532 FILLER_0_5_109/a_572_375# 0 0.232991f
C3534 ctln[5] 0 1.585113f
C3535 output12/a_224_472# 0 2.38465f
C3536 result[7] 0 0.24756f
C3537 net34 0 1.724665f
C3538 output34/a_224_472# 0 2.38465f
C3539 trimb[2] 0 0.839614f
C3540 net45 0 1.12041f
C3541 output45/a_224_472# 0 2.38465f
C3542 ctlp[6] 0 1.243017f
C3543 output23/a_224_472# 0 2.38465f
C3545 FILLER_0_15_142/a_36_472# 0 0.404746f
C3546 FILLER_0_15_142/a_572_375# 0 0.232991f
C3548 _077_ 0 1.645892f
C3549 _075_ 0 0.374516f
C3550 _326_/a_36_160# 0 0.696445f
C3551 _412_/a_2665_112# 0 0.62251f
C3556 _412_/a_36_151# 0 1.43589f
C3557 _091_ 0 1.841339f
C3558 _143_ 0 0.329289f
C3559 mask\[4\] 0 1.300438f
C3560 FILLER_0_13_65/a_36_472# 0 0.417394f
C3561 FILLER_0_13_65/a_124_375# 0 0.246306f
C3562 _360_/a_36_160# 0 0.386641f
C3563 FILLER_0_4_185/a_36_472# 0 0.417394f
C3564 FILLER_0_4_185/a_124_375# 0 0.246306f
C3565 FILLER_0_4_152/a_36_472# 0 0.417394f
C3566 FILLER_0_4_152/a_124_375# 0 0.246306f
C3567 _291_/a_36_160# 0 0.386641f
C3568 ctln[2] 0 1.833091f
C3569 output9/a_224_472# 0 2.38465f
C3570 ctln[4] 0 1.461847f
C3571 output11/a_224_472# 0 2.38465f
C3572 trimb[1] 0 0.378532f
C3573 output44/a_224_472# 0 2.38465f
C3574 result[6] 0 0.19512f
C3575 output33/a_224_472# 0 2.38465f
C3576 ctlp[5] 0 1.282822f
C3577 output22/a_224_472# 0 2.38465f
C3578 FILLER_0_8_127/a_36_472# 0 0.417394f
C3579 FILLER_0_8_127/a_124_375# 0 0.246306f
C3580 FILLER_0_8_138/a_36_472# 0 0.417394f
C3581 FILLER_0_8_138/a_124_375# 0 0.246306f
C3582 FILLER_0_21_133/a_36_472# 0 0.417394f
C3583 FILLER_0_21_133/a_124_375# 0 0.246306f
C3584 FILLER_0_24_130/a_36_472# 0 0.417394f
C3585 FILLER_0_24_130/a_124_375# 0 0.246306f
C3586 FILLER_0_18_171/a_36_472# 0 0.417394f
C3587 FILLER_0_18_171/a_124_375# 0 0.246306f
C3588 _258_/a_36_160# 0 0.386641f
C3589 _016_ 0 0.314121f
C3591 FILLER_0_24_63/a_36_472# 0 0.417394f
C3592 FILLER_0_24_63/a_124_375# 0 0.246306f
C3593 FILLER_0_24_96/a_36_472# 0 0.417394f
C3594 FILLER_0_24_96/a_124_375# 0 0.246306f
C3595 cal_itt\[2\] 0 1.473514f
C3596 _002_ 0 0.289553f
C3597 _413_/a_2665_112# 0 0.62251f
C3602 _413_/a_36_151# 0 1.43589f
C3603 _092_ 0 0.680239f
C3611 FILLER_0_7_72/a_36_472# 0 0.404746f
C3612 FILLER_0_7_72/a_3260_375# 0 0.233093f
C3620 _086_ 0 2.45259f
C3621 _119_ 0 1.237181f
C3622 net63 0 5.362473f
C3623 _430_/a_2665_112# 0 0.62251f
C3628 _430_/a_36_151# 0 1.43589f
C3629 _292_/a_36_160# 0 0.386641f
C3630 comp 0 1.022965f
C3631 ctln[1] 0 1.11973f
C3632 output8/a_224_472# 0 2.38465f
C3633 ctln[3] 0 0.835391f
C3634 output10/a_224_472# 0 2.38465f
C3635 result[5] 0 0.206867f
C3636 net32 0 1.78884f
C3637 output32/a_224_472# 0 2.38465f
C3638 trimb[0] 0 0.847787f
C3639 output43/a_224_472# 0 2.38465f
C3640 ctlp[4] 0 0.37565f
C3641 output21/a_224_472# 0 2.38465f
C3642 _053_ 0 1.705161f
C3644 FILLER_0_16_107/a_36_472# 0 0.404746f
C3645 FILLER_0_16_107/a_572_375# 0 0.232991f
C3647 FILLER_0_3_204/a_36_472# 0 0.417394f
C3648 FILLER_0_3_204/a_124_375# 0 0.246306f
C3656 FILLER_0_9_28/a_36_472# 0 0.404746f
C3657 FILLER_0_9_28/a_3260_375# 0 0.233093f
C3665 _132_ 0 1.491425f
C3666 _328_/a_36_113# 0 0.418095f
C3667 _414_/a_2665_112# 0 0.62251f
C3672 _414_/a_36_151# 0 1.43589f
C3673 _276_/a_36_160# 0 0.386641f
C3674 _144_ 0 1.173846f
C3675 _345_/a_36_160# 0 0.386641f
C3676 _155_ 0 0.638535f
C3677 _020_ 0 0.316793f
C3678 _431_/a_2665_112# 0 0.62251f
C3683 _431_/a_36_151# 0 1.43589f
C3684 _105_ 0 1.21281f
C3686 FILLER_0_5_128/a_36_472# 0 0.404746f
C3687 FILLER_0_5_128/a_572_375# 0 0.232991f
C3689 FILLER_0_5_117/a_36_472# 0 0.417394f
C3690 FILLER_0_5_117/a_124_375# 0 0.246306f
C3691 ctln[0] 0 1.423102f
C3692 net7 0 1.174913f
C3693 output7/a_224_472# 0 2.38465f
C3694 trim[4] 0 0.763069f
C3695 output42/a_224_472# 0 2.38465f
C3696 net31 0 1.912935f
C3697 output31/a_224_472# 0 2.38465f
C3698 ctlp[3] 0 1.14968f
C3699 output20/a_224_472# 0 2.38465f
C3701 FILLER_0_16_73/a_36_472# 0 0.404746f
C3702 FILLER_0_16_73/a_572_375# 0 0.232991f
C3705 FILLER_0_21_142/a_36_472# 0 0.404746f
C3706 FILLER_0_21_142/a_572_375# 0 0.232991f
C3708 FILLER_0_15_150/a_36_472# 0 0.417394f
C3709 FILLER_0_15_150/a_124_375# 0 0.246306f
C3710 FILLER_0_19_125/a_36_472# 0 0.417394f
C3711 FILLER_0_19_125/a_124_375# 0 0.246306f
C3712 net10 0 1.480101f
C3713 net20 0 2.034189f
C3714 _277_/a_36_160# 0 0.386641f
C3715 _004_ 0 0.390107f
C3716 _415_/a_2665_112# 0 0.62251f
C3721 _415_/a_36_151# 0 1.43589f
C3722 mask\[5\] 0 1.334568f
C3723 _028_ 0 0.386029f
C3724 _363_/a_36_68# 0 0.150048f
C3725 _021_ 0 0.316776f
C3726 _432_/a_2665_112# 0 0.62251f
C3731 _432_/a_36_151# 0 1.43589f
C3732 _008_ 0 0.423631f
C3733 _104_ 0 1.435764f
C3734 _106_ 0 0.378703f
C3736 FILLER_0_17_200/a_36_472# 0 0.404746f
C3737 FILLER_0_17_200/a_572_375# 0 0.232991f
.ends


