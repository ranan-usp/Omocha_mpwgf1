magic
tech gf180mcuD
magscale 1 10
timestamp 1701229121
<< metal1 >>
rect 1344 22762 34608 22796
rect 1344 22710 5372 22762
rect 5424 22710 5476 22762
rect 5528 22710 5580 22762
rect 5632 22710 13688 22762
rect 13740 22710 13792 22762
rect 13844 22710 13896 22762
rect 13948 22710 22004 22762
rect 22056 22710 22108 22762
rect 22160 22710 22212 22762
rect 22264 22710 30320 22762
rect 30372 22710 30424 22762
rect 30476 22710 30528 22762
rect 30580 22710 34608 22762
rect 1344 22676 34608 22710
rect 2270 22594 2322 22606
rect 2270 22530 2322 22542
rect 6638 22594 6690 22606
rect 6638 22530 6690 22542
rect 9550 22594 9602 22606
rect 9550 22530 9602 22542
rect 14142 22594 14194 22606
rect 14142 22530 14194 22542
rect 17166 22594 17218 22606
rect 17166 22530 17218 22542
rect 20974 22594 21026 22606
rect 20974 22530 21026 22542
rect 25566 22594 25618 22606
rect 25566 22530 25618 22542
rect 28590 22594 28642 22606
rect 28590 22530 28642 22542
rect 4162 22318 4174 22370
rect 4226 22318 4238 22370
rect 5954 22318 5966 22370
rect 6018 22318 6030 22370
rect 11442 22318 11454 22370
rect 11506 22318 11518 22370
rect 13122 22318 13134 22370
rect 13186 22318 13198 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 23314 22318 23326 22370
rect 23378 22318 23390 22370
rect 24546 22318 24558 22370
rect 24610 22318 24622 22370
rect 27794 22318 27806 22370
rect 27858 22318 27870 22370
rect 30930 22318 30942 22370
rect 30994 22318 31006 22370
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 19966 22146 20018 22158
rect 19966 22082 20018 22094
rect 23774 22146 23826 22158
rect 23774 22082 23826 22094
rect 27582 22146 27634 22158
rect 27582 22082 27634 22094
rect 31390 22146 31442 22158
rect 31390 22082 31442 22094
rect 1344 21978 34768 22012
rect 1344 21926 9530 21978
rect 9582 21926 9634 21978
rect 9686 21926 9738 21978
rect 9790 21926 17846 21978
rect 17898 21926 17950 21978
rect 18002 21926 18054 21978
rect 18106 21926 26162 21978
rect 26214 21926 26266 21978
rect 26318 21926 26370 21978
rect 26422 21926 34478 21978
rect 34530 21926 34582 21978
rect 34634 21926 34686 21978
rect 34738 21926 34768 21978
rect 1344 21892 34768 21926
rect 10670 21810 10722 21822
rect 12910 21810 12962 21822
rect 20638 21810 20690 21822
rect 10322 21758 10334 21810
rect 10386 21758 10398 21810
rect 10994 21758 11006 21810
rect 11058 21758 11070 21810
rect 12562 21758 12574 21810
rect 12626 21758 12638 21810
rect 17378 21758 17390 21810
rect 17442 21758 17454 21810
rect 10670 21746 10722 21758
rect 12910 21746 12962 21758
rect 20638 21746 20690 21758
rect 26574 21810 26626 21822
rect 26574 21746 26626 21758
rect 8990 21698 9042 21710
rect 8990 21634 9042 21646
rect 12126 21698 12178 21710
rect 12126 21634 12178 21646
rect 16158 21698 16210 21710
rect 16158 21634 16210 21646
rect 23886 21698 23938 21710
rect 23886 21634 23938 21646
rect 27918 21698 27970 21710
rect 27918 21634 27970 21646
rect 31278 21698 31330 21710
rect 31278 21634 31330 21646
rect 4622 21586 4674 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 4622 21522 4674 21534
rect 13246 21586 13298 21598
rect 18958 21586 19010 21598
rect 19518 21586 19570 21598
rect 13906 21534 13918 21586
rect 13970 21534 13982 21586
rect 19282 21534 19294 21586
rect 19346 21534 19358 21586
rect 13246 21522 13298 21534
rect 18958 21522 19010 21534
rect 19518 21522 19570 21534
rect 19742 21586 19794 21598
rect 20974 21586 21026 21598
rect 25230 21586 25282 21598
rect 19954 21534 19966 21586
rect 20018 21534 20030 21586
rect 21522 21534 21534 21586
rect 21586 21534 21598 21586
rect 19742 21522 19794 21534
rect 20974 21522 21026 21534
rect 25230 21522 25282 21534
rect 25454 21586 25506 21598
rect 25454 21522 25506 21534
rect 25902 21586 25954 21598
rect 25902 21522 25954 21534
rect 26126 21586 26178 21598
rect 26126 21522 26178 21534
rect 26350 21586 26402 21598
rect 26350 21522 26402 21534
rect 26798 21586 26850 21598
rect 30830 21586 30882 21598
rect 30146 21534 30158 21586
rect 30210 21534 30222 21586
rect 26798 21522 26850 21534
rect 30830 21522 30882 21534
rect 1934 21474 1986 21486
rect 1934 21410 1986 21422
rect 4734 21474 4786 21486
rect 4734 21410 4786 21422
rect 5182 21474 5234 21486
rect 5182 21410 5234 21422
rect 5630 21474 5682 21486
rect 5630 21410 5682 21422
rect 6078 21474 6130 21486
rect 6078 21410 6130 21422
rect 9774 21474 9826 21486
rect 9774 21410 9826 21422
rect 17950 21474 18002 21486
rect 19630 21474 19682 21486
rect 18498 21422 18510 21474
rect 18562 21422 18574 21474
rect 17950 21410 18002 21422
rect 19630 21410 19682 21422
rect 20526 21474 20578 21486
rect 20526 21410 20578 21422
rect 25678 21474 25730 21486
rect 25678 21410 25730 21422
rect 31054 21474 31106 21486
rect 31054 21410 31106 21422
rect 31838 21474 31890 21486
rect 31838 21410 31890 21422
rect 5070 21362 5122 21374
rect 5070 21298 5122 21310
rect 8878 21362 8930 21374
rect 8878 21298 8930 21310
rect 9998 21362 10050 21374
rect 9998 21298 10050 21310
rect 12238 21362 12290 21374
rect 12238 21298 12290 21310
rect 16942 21362 16994 21374
rect 16942 21298 16994 21310
rect 17726 21362 17778 21374
rect 17726 21298 17778 21310
rect 24670 21362 24722 21374
rect 24670 21298 24722 21310
rect 27134 21362 27186 21374
rect 27134 21298 27186 21310
rect 31390 21362 31442 21374
rect 31390 21298 31442 21310
rect 1344 21194 34608 21228
rect 1344 21142 5372 21194
rect 5424 21142 5476 21194
rect 5528 21142 5580 21194
rect 5632 21142 13688 21194
rect 13740 21142 13792 21194
rect 13844 21142 13896 21194
rect 13948 21142 22004 21194
rect 22056 21142 22108 21194
rect 22160 21142 22212 21194
rect 22264 21142 30320 21194
rect 30372 21142 30424 21194
rect 30476 21142 30528 21194
rect 30580 21142 34608 21194
rect 1344 21108 34608 21142
rect 14366 21026 14418 21038
rect 14366 20962 14418 20974
rect 19406 21026 19458 21038
rect 19406 20962 19458 20974
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 4734 20914 4786 20926
rect 4734 20850 4786 20862
rect 9550 20914 9602 20926
rect 9550 20850 9602 20862
rect 19966 20914 20018 20926
rect 27582 20914 27634 20926
rect 25106 20862 25118 20914
rect 25170 20862 25182 20914
rect 19966 20850 20018 20862
rect 27582 20850 27634 20862
rect 29598 20914 29650 20926
rect 29598 20850 29650 20862
rect 30046 20914 30098 20926
rect 30046 20850 30098 20862
rect 30158 20914 30210 20926
rect 30158 20850 30210 20862
rect 5854 20802 5906 20814
rect 9774 20802 9826 20814
rect 3826 20750 3838 20802
rect 3890 20750 3902 20802
rect 6514 20750 6526 20802
rect 6578 20750 6590 20802
rect 5854 20738 5906 20750
rect 9774 20738 9826 20750
rect 9998 20802 10050 20814
rect 9998 20738 10050 20750
rect 10446 20802 10498 20814
rect 15262 20802 15314 20814
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 10446 20738 10498 20750
rect 15262 20738 15314 20750
rect 19742 20802 19794 20814
rect 29150 20802 29202 20814
rect 23090 20750 23102 20802
rect 23154 20750 23166 20802
rect 28466 20750 28478 20802
rect 28530 20750 28542 20802
rect 19742 20738 19794 20750
rect 29150 20738 29202 20750
rect 29374 20802 29426 20814
rect 34078 20802 34130 20814
rect 30370 20750 30382 20802
rect 30434 20750 30446 20802
rect 33618 20750 33630 20802
rect 33682 20750 33694 20802
rect 29374 20738 29426 20750
rect 34078 20738 34130 20750
rect 14478 20690 14530 20702
rect 14478 20626 14530 20638
rect 15150 20690 15202 20702
rect 15150 20626 15202 20638
rect 20302 20690 20354 20702
rect 20302 20626 20354 20638
rect 29710 20690 29762 20702
rect 29710 20626 29762 20638
rect 10110 20578 10162 20590
rect 8754 20526 8766 20578
rect 8818 20526 8830 20578
rect 10110 20514 10162 20526
rect 10894 20578 10946 20590
rect 10894 20514 10946 20526
rect 15038 20578 15090 20590
rect 15038 20514 15090 20526
rect 15374 20578 15426 20590
rect 15374 20514 15426 20526
rect 20414 20578 20466 20590
rect 20414 20514 20466 20526
rect 30606 20578 30658 20590
rect 31378 20526 31390 20578
rect 31442 20526 31454 20578
rect 30606 20514 30658 20526
rect 1344 20410 34768 20444
rect 1344 20358 9530 20410
rect 9582 20358 9634 20410
rect 9686 20358 9738 20410
rect 9790 20358 17846 20410
rect 17898 20358 17950 20410
rect 18002 20358 18054 20410
rect 18106 20358 26162 20410
rect 26214 20358 26266 20410
rect 26318 20358 26370 20410
rect 26422 20358 34478 20410
rect 34530 20358 34582 20410
rect 34634 20358 34686 20410
rect 34738 20358 34768 20410
rect 1344 20324 34768 20358
rect 14254 20242 14306 20254
rect 14254 20178 14306 20190
rect 14926 20242 14978 20254
rect 23090 20190 23102 20242
rect 23154 20190 23166 20242
rect 14926 20178 14978 20190
rect 9662 20130 9714 20142
rect 9662 20066 9714 20078
rect 9774 20130 9826 20142
rect 9774 20066 9826 20078
rect 9886 20130 9938 20142
rect 9886 20066 9938 20078
rect 13470 20130 13522 20142
rect 13470 20066 13522 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 19742 20130 19794 20142
rect 19742 20066 19794 20078
rect 28926 20130 28978 20142
rect 28926 20066 28978 20078
rect 29710 20130 29762 20142
rect 29710 20066 29762 20078
rect 10558 20018 10610 20030
rect 14702 20018 14754 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 11218 19966 11230 20018
rect 11282 19966 11294 20018
rect 14466 19966 14478 20018
rect 14530 19966 14542 20018
rect 10558 19954 10610 19966
rect 14702 19954 14754 19966
rect 15038 20018 15090 20030
rect 19294 20018 19346 20030
rect 19058 19966 19070 20018
rect 19122 19966 19134 20018
rect 15038 19954 15090 19966
rect 19294 19954 19346 19966
rect 19518 20018 19570 20030
rect 19518 19954 19570 19966
rect 20414 20018 20466 20030
rect 25566 20018 25618 20030
rect 32622 20018 32674 20030
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 26562 19966 26574 20018
rect 26626 19966 26638 20018
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 20414 19954 20466 19966
rect 25566 19954 25618 19966
rect 32622 19954 32674 19966
rect 10334 19906 10386 19918
rect 2034 19854 2046 19906
rect 2098 19854 2110 19906
rect 10334 19842 10386 19854
rect 14814 19906 14866 19918
rect 14814 19842 14866 19854
rect 24222 19906 24274 19918
rect 24222 19842 24274 19854
rect 25790 19906 25842 19918
rect 25790 19842 25842 19854
rect 28478 19906 28530 19918
rect 28478 19842 28530 19854
rect 33294 19906 33346 19918
rect 33294 19842 33346 19854
rect 23886 19794 23938 19806
rect 23886 19730 23938 19742
rect 25230 19794 25282 19806
rect 25230 19730 25282 19742
rect 1344 19626 34608 19660
rect 1344 19574 5372 19626
rect 5424 19574 5476 19626
rect 5528 19574 5580 19626
rect 5632 19574 13688 19626
rect 13740 19574 13792 19626
rect 13844 19574 13896 19626
rect 13948 19574 22004 19626
rect 22056 19574 22108 19626
rect 22160 19574 22212 19626
rect 22264 19574 30320 19626
rect 30372 19574 30424 19626
rect 30476 19574 30528 19626
rect 30580 19574 34608 19626
rect 1344 19540 34608 19574
rect 2718 19458 2770 19470
rect 2718 19394 2770 19406
rect 12014 19458 12066 19470
rect 12014 19394 12066 19406
rect 27582 19458 27634 19470
rect 27582 19394 27634 19406
rect 10446 19346 10498 19358
rect 10446 19282 10498 19294
rect 12126 19346 12178 19358
rect 12126 19282 12178 19294
rect 23998 19346 24050 19358
rect 24434 19294 24446 19346
rect 24498 19294 24510 19346
rect 23998 19282 24050 19294
rect 9662 19234 9714 19246
rect 5618 19182 5630 19234
rect 5682 19182 5694 19234
rect 6178 19182 6190 19234
rect 6242 19182 6254 19234
rect 9662 19170 9714 19182
rect 10110 19234 10162 19246
rect 10110 19170 10162 19182
rect 14814 19234 14866 19246
rect 19182 19234 19234 19246
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 14814 19170 14866 19182
rect 19182 19170 19234 19182
rect 20078 19234 20130 19246
rect 20078 19170 20130 19182
rect 24894 19234 24946 19246
rect 24894 19170 24946 19182
rect 25342 19234 25394 19246
rect 32734 19234 32786 19246
rect 28466 19182 28478 19234
rect 28530 19182 28542 19234
rect 32050 19182 32062 19234
rect 32114 19182 32126 19234
rect 33170 19182 33182 19234
rect 33234 19182 33246 19234
rect 25342 19170 25394 19182
rect 32734 19170 32786 19182
rect 2830 19122 2882 19134
rect 2830 19058 2882 19070
rect 9214 19122 9266 19134
rect 9214 19058 9266 19070
rect 9438 19122 9490 19134
rect 9438 19058 9490 19070
rect 14254 19122 14306 19134
rect 14254 19058 14306 19070
rect 14590 19122 14642 19134
rect 14590 19058 14642 19070
rect 17726 19122 17778 19134
rect 17726 19058 17778 19070
rect 18510 19122 18562 19134
rect 18510 19058 18562 19070
rect 19406 19122 19458 19134
rect 33854 19122 33906 19134
rect 25666 19070 25678 19122
rect 25730 19070 25742 19122
rect 19406 19058 19458 19070
rect 33854 19058 33906 19070
rect 34190 19122 34242 19134
rect 34190 19058 34242 19070
rect 9886 19010 9938 19022
rect 8642 18958 8654 19010
rect 8706 18958 8718 19010
rect 9886 18946 9938 18958
rect 10894 19010 10946 19022
rect 10894 18946 10946 18958
rect 18846 19010 18898 19022
rect 18846 18946 18898 18958
rect 18958 19010 19010 19022
rect 18958 18946 19010 18958
rect 19070 19010 19122 19022
rect 29038 19010 29090 19022
rect 32958 19010 33010 19022
rect 19730 18958 19742 19010
rect 19794 18958 19806 19010
rect 29810 18958 29822 19010
rect 29874 18958 29886 19010
rect 19070 18946 19122 18958
rect 29038 18946 29090 18958
rect 32958 18946 33010 18958
rect 1344 18842 34768 18876
rect 1344 18790 9530 18842
rect 9582 18790 9634 18842
rect 9686 18790 9738 18842
rect 9790 18790 17846 18842
rect 17898 18790 17950 18842
rect 18002 18790 18054 18842
rect 18106 18790 26162 18842
rect 26214 18790 26266 18842
rect 26318 18790 26370 18842
rect 26422 18790 34478 18842
rect 34530 18790 34582 18842
rect 34634 18790 34686 18842
rect 34738 18790 34768 18842
rect 1344 18756 34768 18790
rect 9662 18674 9714 18686
rect 14814 18674 14866 18686
rect 16046 18674 16098 18686
rect 33742 18674 33794 18686
rect 5954 18622 5966 18674
rect 6018 18622 6030 18674
rect 13122 18622 13134 18674
rect 13186 18622 13198 18674
rect 15138 18622 15150 18674
rect 15202 18622 15214 18674
rect 19954 18622 19966 18674
rect 20018 18622 20030 18674
rect 9662 18610 9714 18622
rect 14814 18610 14866 18622
rect 16046 18610 16098 18622
rect 33742 18610 33794 18622
rect 8990 18562 9042 18574
rect 8990 18498 9042 18510
rect 6414 18450 6466 18462
rect 2146 18398 2158 18450
rect 2210 18398 2222 18450
rect 5730 18398 5742 18450
rect 5794 18398 5806 18450
rect 6414 18386 6466 18398
rect 8766 18450 8818 18462
rect 8766 18386 8818 18398
rect 10222 18450 10274 18462
rect 13694 18450 13746 18462
rect 10658 18398 10670 18450
rect 10722 18398 10734 18450
rect 10222 18386 10274 18398
rect 13694 18386 13746 18398
rect 16158 18450 16210 18462
rect 16158 18386 16210 18398
rect 17950 18450 18002 18462
rect 20302 18450 20354 18462
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 17950 18386 18002 18398
rect 20302 18386 20354 18398
rect 24446 18450 24498 18462
rect 24446 18386 24498 18398
rect 25566 18450 25618 18462
rect 25566 18386 25618 18398
rect 26238 18450 26290 18462
rect 26238 18386 26290 18398
rect 26462 18450 26514 18462
rect 26462 18386 26514 18398
rect 26798 18450 26850 18462
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 29922 18398 29934 18450
rect 29986 18398 29998 18450
rect 33394 18398 33406 18450
rect 33458 18398 33470 18450
rect 33954 18398 33966 18450
rect 34018 18398 34030 18450
rect 26798 18386 26850 18398
rect 8430 18338 8482 18350
rect 25230 18338 25282 18350
rect 23986 18286 23998 18338
rect 24050 18286 24062 18338
rect 8430 18274 8482 18286
rect 25230 18274 25282 18286
rect 25790 18338 25842 18350
rect 25790 18274 25842 18286
rect 26574 18338 26626 18350
rect 26574 18274 26626 18286
rect 29374 18338 29426 18350
rect 31826 18286 31838 18338
rect 31890 18286 31902 18338
rect 29374 18274 29426 18286
rect 2718 18226 2770 18238
rect 2718 18162 2770 18174
rect 6302 18226 6354 18238
rect 6302 18162 6354 18174
rect 33070 18226 33122 18238
rect 33070 18162 33122 18174
rect 33406 18226 33458 18238
rect 33406 18162 33458 18174
rect 1344 18058 34608 18092
rect 1344 18006 5372 18058
rect 5424 18006 5476 18058
rect 5528 18006 5580 18058
rect 5632 18006 13688 18058
rect 13740 18006 13792 18058
rect 13844 18006 13896 18058
rect 13948 18006 22004 18058
rect 22056 18006 22108 18058
rect 22160 18006 22212 18058
rect 22264 18006 30320 18058
rect 30372 18006 30424 18058
rect 30476 18006 30528 18058
rect 30580 18006 34608 18058
rect 1344 17972 34608 18006
rect 9214 17890 9266 17902
rect 9214 17826 9266 17838
rect 10894 17890 10946 17902
rect 10894 17826 10946 17838
rect 29934 17890 29986 17902
rect 29934 17826 29986 17838
rect 8978 17726 8990 17778
rect 9042 17726 9054 17778
rect 27570 17726 27582 17778
rect 27634 17726 27646 17778
rect 11006 17666 11058 17678
rect 11006 17602 11058 17614
rect 11454 17666 11506 17678
rect 11454 17602 11506 17614
rect 11678 17666 11730 17678
rect 11678 17602 11730 17614
rect 11790 17666 11842 17678
rect 11790 17602 11842 17614
rect 12014 17666 12066 17678
rect 12014 17602 12066 17614
rect 19294 17666 19346 17678
rect 19294 17602 19346 17614
rect 19518 17666 19570 17678
rect 19518 17602 19570 17614
rect 20190 17666 20242 17678
rect 26574 17666 26626 17678
rect 34078 17666 34130 17678
rect 26114 17614 26126 17666
rect 26178 17614 26190 17666
rect 30258 17614 30270 17666
rect 30322 17614 30334 17666
rect 33618 17614 33630 17666
rect 33682 17614 33694 17666
rect 20190 17602 20242 17614
rect 26574 17602 26626 17614
rect 34078 17602 34130 17614
rect 8990 17554 9042 17566
rect 8990 17490 9042 17502
rect 9662 17554 9714 17566
rect 29474 17502 29486 17554
rect 29538 17502 29550 17554
rect 9662 17490 9714 17502
rect 12350 17442 12402 17454
rect 12350 17378 12402 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 19630 17442 19682 17454
rect 19630 17378 19682 17390
rect 19742 17442 19794 17454
rect 19742 17378 19794 17390
rect 20302 17442 20354 17454
rect 28030 17442 28082 17454
rect 25890 17390 25902 17442
rect 25954 17390 25966 17442
rect 26898 17390 26910 17442
rect 26962 17390 26974 17442
rect 20302 17378 20354 17390
rect 28030 17378 28082 17390
rect 28590 17442 28642 17454
rect 28590 17378 28642 17390
rect 29150 17442 29202 17454
rect 29150 17378 29202 17390
rect 30046 17442 30098 17454
rect 30046 17378 30098 17390
rect 30606 17442 30658 17454
rect 31378 17390 31390 17442
rect 31442 17390 31454 17442
rect 30606 17378 30658 17390
rect 1344 17274 34768 17308
rect 1344 17222 9530 17274
rect 9582 17222 9634 17274
rect 9686 17222 9738 17274
rect 9790 17222 17846 17274
rect 17898 17222 17950 17274
rect 18002 17222 18054 17274
rect 18106 17222 26162 17274
rect 26214 17222 26266 17274
rect 26318 17222 26370 17274
rect 26422 17222 34478 17274
rect 34530 17222 34582 17274
rect 34634 17222 34686 17274
rect 34738 17222 34768 17274
rect 1344 17188 34768 17222
rect 15262 17106 15314 17118
rect 23662 17106 23714 17118
rect 23090 17054 23102 17106
rect 23154 17054 23166 17106
rect 15262 17042 15314 17054
rect 23662 17042 23714 17054
rect 25454 17106 25506 17118
rect 25454 17042 25506 17054
rect 27582 17106 27634 17118
rect 29150 17106 29202 17118
rect 28130 17054 28142 17106
rect 28194 17054 28206 17106
rect 27582 17042 27634 17054
rect 29150 17042 29202 17054
rect 34190 17106 34242 17118
rect 34190 17042 34242 17054
rect 19182 16994 19234 17006
rect 15586 16942 15598 16994
rect 15650 16942 15662 16994
rect 19182 16930 19234 16942
rect 28702 16994 28754 17006
rect 28702 16930 28754 16942
rect 29598 16994 29650 17006
rect 29598 16930 29650 16942
rect 6862 16882 6914 16894
rect 2706 16830 2718 16882
rect 2770 16830 2782 16882
rect 4946 16830 4958 16882
rect 5010 16830 5022 16882
rect 5506 16830 5518 16882
rect 5570 16830 5582 16882
rect 6862 16818 6914 16830
rect 6974 16882 7026 16894
rect 6974 16818 7026 16830
rect 7198 16882 7250 16894
rect 7198 16818 7250 16830
rect 7422 16882 7474 16894
rect 7422 16818 7474 16830
rect 16046 16882 16098 16894
rect 16046 16818 16098 16830
rect 18622 16882 18674 16894
rect 18622 16818 18674 16830
rect 18734 16882 18786 16894
rect 18734 16818 18786 16830
rect 18958 16882 19010 16894
rect 29038 16882 29090 16894
rect 20066 16830 20078 16882
rect 20130 16830 20142 16882
rect 20514 16830 20526 16882
rect 20578 16830 20590 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 18958 16818 19010 16830
rect 29038 16818 29090 16830
rect 29262 16882 29314 16894
rect 33630 16882 33682 16894
rect 29922 16830 29934 16882
rect 29986 16830 29998 16882
rect 31602 16830 31614 16882
rect 31666 16830 31678 16882
rect 29262 16818 29314 16830
rect 33630 16818 33682 16830
rect 18846 16770 18898 16782
rect 18846 16706 18898 16718
rect 27358 16770 27410 16782
rect 28478 16770 28530 16782
rect 27682 16718 27694 16770
rect 27746 16718 27758 16770
rect 27358 16706 27410 16718
rect 28478 16706 28530 16718
rect 15934 16658 15986 16670
rect 1698 16606 1710 16658
rect 1762 16606 1774 16658
rect 15934 16594 15986 16606
rect 25566 16658 25618 16670
rect 25566 16594 25618 16606
rect 1344 16490 34608 16524
rect 1344 16438 5372 16490
rect 5424 16438 5476 16490
rect 5528 16438 5580 16490
rect 5632 16438 13688 16490
rect 13740 16438 13792 16490
rect 13844 16438 13896 16490
rect 13948 16438 22004 16490
rect 22056 16438 22108 16490
rect 22160 16438 22212 16490
rect 22264 16438 30320 16490
rect 30372 16438 30424 16490
rect 30476 16438 30528 16490
rect 30580 16438 34608 16490
rect 1344 16404 34608 16438
rect 1934 16210 1986 16222
rect 1934 16146 1986 16158
rect 7422 16210 7474 16222
rect 29262 16210 29314 16222
rect 22530 16158 22542 16210
rect 22594 16158 22606 16210
rect 7422 16146 7474 16158
rect 29262 16146 29314 16158
rect 4734 16098 4786 16110
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 4734 16034 4786 16046
rect 10446 16098 10498 16110
rect 10446 16034 10498 16046
rect 10782 16098 10834 16110
rect 10782 16034 10834 16046
rect 11006 16098 11058 16110
rect 11006 16034 11058 16046
rect 14814 16098 14866 16110
rect 22206 16098 22258 16110
rect 15474 16046 15486 16098
rect 15538 16046 15550 16098
rect 21410 16046 21422 16098
rect 21474 16046 21486 16098
rect 14814 16034 14866 16046
rect 22206 16034 22258 16046
rect 22990 16098 23042 16110
rect 26910 16098 26962 16110
rect 23538 16046 23550 16098
rect 23602 16046 23614 16098
rect 22990 16034 23042 16046
rect 26910 16034 26962 16046
rect 29374 16098 29426 16110
rect 34078 16098 34130 16110
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 29374 16034 29426 16046
rect 34078 16034 34130 16046
rect 6190 15986 6242 15998
rect 6190 15922 6242 15934
rect 7534 15986 7586 15998
rect 7534 15922 7586 15934
rect 21982 15986 22034 15998
rect 21982 15922 22034 15934
rect 29150 15986 29202 15998
rect 29150 15922 29202 15934
rect 29710 15986 29762 15998
rect 29710 15922 29762 15934
rect 30606 15986 30658 15998
rect 30606 15922 30658 15934
rect 6302 15874 6354 15886
rect 6302 15810 6354 15822
rect 6414 15874 6466 15886
rect 6414 15810 6466 15822
rect 7310 15874 7362 15886
rect 7310 15810 7362 15822
rect 10782 15874 10834 15886
rect 18510 15874 18562 15886
rect 17714 15822 17726 15874
rect 17778 15822 17790 15874
rect 10782 15810 10834 15822
rect 18510 15810 18562 15822
rect 20414 15874 20466 15886
rect 22430 15874 22482 15886
rect 21634 15822 21646 15874
rect 21698 15822 21710 15874
rect 20414 15810 20466 15822
rect 22430 15810 22482 15822
rect 22542 15874 22594 15886
rect 26686 15874 26738 15886
rect 26114 15822 26126 15874
rect 26178 15822 26190 15874
rect 22542 15810 22594 15822
rect 26686 15810 26738 15822
rect 27470 15874 27522 15886
rect 27470 15810 27522 15822
rect 27806 15874 27858 15886
rect 28130 15822 28142 15874
rect 28194 15822 28206 15874
rect 31378 15822 31390 15874
rect 31442 15822 31454 15874
rect 27806 15810 27858 15822
rect 1344 15706 34768 15740
rect 1344 15654 9530 15706
rect 9582 15654 9634 15706
rect 9686 15654 9738 15706
rect 9790 15654 17846 15706
rect 17898 15654 17950 15706
rect 18002 15654 18054 15706
rect 18106 15654 26162 15706
rect 26214 15654 26266 15706
rect 26318 15654 26370 15706
rect 26422 15654 34478 15706
rect 34530 15654 34582 15706
rect 34634 15654 34686 15706
rect 34738 15654 34768 15706
rect 1344 15620 34768 15654
rect 7198 15538 7250 15550
rect 7198 15474 7250 15486
rect 19854 15538 19906 15550
rect 19854 15474 19906 15486
rect 20638 15538 20690 15550
rect 20638 15474 20690 15486
rect 22990 15538 23042 15550
rect 22990 15474 23042 15486
rect 23326 15538 23378 15550
rect 23326 15474 23378 15486
rect 27470 15538 27522 15550
rect 27470 15474 27522 15486
rect 28702 15538 28754 15550
rect 28702 15474 28754 15486
rect 3390 15426 3442 15438
rect 3390 15362 3442 15374
rect 6862 15426 6914 15438
rect 6862 15362 6914 15374
rect 7646 15426 7698 15438
rect 7646 15362 7698 15374
rect 15598 15426 15650 15438
rect 15598 15362 15650 15374
rect 15934 15426 15986 15438
rect 15934 15362 15986 15374
rect 16270 15426 16322 15438
rect 16270 15362 16322 15374
rect 22878 15426 22930 15438
rect 22878 15362 22930 15374
rect 29038 15426 29090 15438
rect 29038 15362 29090 15374
rect 3838 15314 3890 15326
rect 7310 15314 7362 15326
rect 4946 15262 4958 15314
rect 5010 15262 5022 15314
rect 6402 15262 6414 15314
rect 6466 15262 6478 15314
rect 3838 15250 3890 15262
rect 7310 15250 7362 15262
rect 7422 15314 7474 15326
rect 20526 15314 20578 15326
rect 23662 15314 23714 15326
rect 11442 15262 11454 15314
rect 11506 15262 11518 15314
rect 13570 15262 13582 15314
rect 13634 15262 13646 15314
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 19394 15262 19406 15314
rect 19458 15262 19470 15314
rect 20066 15262 20078 15314
rect 20130 15262 20142 15314
rect 20850 15262 20862 15314
rect 20914 15262 20926 15314
rect 7422 15250 7474 15262
rect 20526 15250 20578 15262
rect 23662 15250 23714 15262
rect 29262 15314 29314 15326
rect 29922 15262 29934 15314
rect 29986 15262 29998 15314
rect 29262 15250 29314 15262
rect 3614 15202 3666 15214
rect 18958 15202 19010 15214
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 3614 15138 3666 15150
rect 18958 15138 19010 15150
rect 24110 15202 24162 15214
rect 31042 15150 31054 15202
rect 31106 15150 31118 15202
rect 24110 15138 24162 15150
rect 29598 15090 29650 15102
rect 4162 15038 4174 15090
rect 4226 15038 4238 15090
rect 10434 15038 10446 15090
rect 10498 15038 10510 15090
rect 29598 15026 29650 15038
rect 1344 14922 34608 14956
rect 1344 14870 5372 14922
rect 5424 14870 5476 14922
rect 5528 14870 5580 14922
rect 5632 14870 13688 14922
rect 13740 14870 13792 14922
rect 13844 14870 13896 14922
rect 13948 14870 22004 14922
rect 22056 14870 22108 14922
rect 22160 14870 22212 14922
rect 22264 14870 30320 14922
rect 30372 14870 30424 14922
rect 30476 14870 30528 14922
rect 30580 14870 34608 14922
rect 1344 14836 34608 14870
rect 4398 14754 4450 14766
rect 4398 14690 4450 14702
rect 11006 14754 11058 14766
rect 33506 14702 33518 14754
rect 33570 14702 33582 14754
rect 11006 14690 11058 14702
rect 10222 14642 10274 14654
rect 8082 14590 8094 14642
rect 8146 14590 8158 14642
rect 10222 14578 10274 14590
rect 20526 14642 20578 14654
rect 22866 14590 22878 14642
rect 22930 14590 22942 14642
rect 20526 14578 20578 14590
rect 2606 14530 2658 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 2606 14466 2658 14478
rect 3278 14530 3330 14542
rect 3278 14466 3330 14478
rect 3838 14530 3890 14542
rect 3838 14466 3890 14478
rect 5518 14530 5570 14542
rect 5518 14466 5570 14478
rect 5854 14530 5906 14542
rect 5854 14466 5906 14478
rect 6078 14530 6130 14542
rect 6078 14466 6130 14478
rect 6526 14530 6578 14542
rect 6526 14466 6578 14478
rect 6862 14530 6914 14542
rect 6862 14466 6914 14478
rect 15822 14530 15874 14542
rect 22430 14530 22482 14542
rect 16370 14478 16382 14530
rect 16434 14478 16446 14530
rect 15822 14466 15874 14478
rect 22430 14466 22482 14478
rect 22542 14530 22594 14542
rect 23550 14530 23602 14542
rect 29038 14530 29090 14542
rect 22978 14478 22990 14530
rect 23042 14478 23054 14530
rect 23986 14478 23998 14530
rect 24050 14478 24062 14530
rect 24434 14478 24446 14530
rect 24498 14478 24510 14530
rect 22542 14466 22594 14478
rect 23550 14466 23602 14478
rect 29038 14466 29090 14478
rect 30046 14530 30098 14542
rect 30046 14466 30098 14478
rect 30606 14530 30658 14542
rect 31714 14478 31726 14530
rect 31778 14478 31790 14530
rect 30606 14466 30658 14478
rect 2046 14418 2098 14430
rect 2046 14354 2098 14366
rect 2942 14418 2994 14430
rect 2942 14354 2994 14366
rect 4174 14418 4226 14430
rect 4174 14354 4226 14366
rect 6638 14418 6690 14430
rect 11118 14418 11170 14430
rect 8530 14366 8542 14418
rect 8594 14366 8606 14418
rect 9986 14366 9998 14418
rect 10050 14366 10062 14418
rect 6638 14354 6690 14366
rect 11118 14354 11170 14366
rect 11342 14418 11394 14430
rect 11342 14354 11394 14366
rect 18734 14418 18786 14430
rect 18734 14354 18786 14366
rect 20638 14418 20690 14430
rect 20638 14354 20690 14366
rect 23662 14418 23714 14430
rect 23662 14354 23714 14366
rect 26798 14418 26850 14430
rect 26798 14354 26850 14366
rect 29486 14418 29538 14430
rect 29486 14354 29538 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 5742 14306 5794 14318
rect 4722 14254 4734 14306
rect 4786 14254 4798 14306
rect 5742 14242 5794 14254
rect 7646 14306 7698 14318
rect 7646 14242 7698 14254
rect 19518 14306 19570 14318
rect 19518 14242 19570 14254
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 22766 14306 22818 14318
rect 22766 14242 22818 14254
rect 27582 14306 27634 14318
rect 27582 14242 27634 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 1344 14138 34768 14172
rect 1344 14086 9530 14138
rect 9582 14086 9634 14138
rect 9686 14086 9738 14138
rect 9790 14086 17846 14138
rect 17898 14086 17950 14138
rect 18002 14086 18054 14138
rect 18106 14086 26162 14138
rect 26214 14086 26266 14138
rect 26318 14086 26370 14138
rect 26422 14086 34478 14138
rect 34530 14086 34582 14138
rect 34634 14086 34686 14138
rect 34738 14086 34768 14138
rect 1344 14052 34768 14086
rect 1822 13970 1874 13982
rect 1822 13906 1874 13918
rect 2942 13970 2994 13982
rect 2942 13906 2994 13918
rect 6526 13970 6578 13982
rect 6526 13906 6578 13918
rect 7534 13970 7586 13982
rect 7534 13906 7586 13918
rect 8094 13970 8146 13982
rect 21758 13970 21810 13982
rect 29486 13970 29538 13982
rect 16146 13918 16158 13970
rect 16210 13918 16222 13970
rect 27458 13918 27470 13970
rect 27522 13918 27534 13970
rect 8094 13906 8146 13918
rect 21758 13906 21810 13918
rect 29486 13906 29538 13918
rect 3390 13858 3442 13870
rect 22206 13858 22258 13870
rect 4386 13806 4398 13858
rect 4450 13806 4462 13858
rect 5730 13806 5742 13858
rect 5794 13806 5806 13858
rect 19842 13806 19854 13858
rect 19906 13806 19918 13858
rect 3390 13794 3442 13806
rect 22206 13794 22258 13806
rect 28590 13858 28642 13870
rect 28590 13794 28642 13806
rect 29262 13858 29314 13870
rect 29262 13794 29314 13806
rect 10894 13746 10946 13758
rect 4610 13694 4622 13746
rect 4674 13694 4686 13746
rect 8306 13694 8318 13746
rect 8370 13694 8382 13746
rect 10894 13682 10946 13694
rect 11454 13746 11506 13758
rect 11454 13682 11506 13694
rect 11902 13746 11954 13758
rect 19518 13746 19570 13758
rect 21758 13746 21810 13758
rect 13346 13694 13358 13746
rect 13410 13694 13422 13746
rect 13906 13694 13918 13746
rect 13970 13694 13982 13746
rect 20626 13694 20638 13746
rect 20690 13694 20702 13746
rect 21074 13694 21086 13746
rect 21138 13694 21150 13746
rect 11902 13682 11954 13694
rect 19518 13682 19570 13694
rect 21758 13682 21810 13694
rect 23438 13746 23490 13758
rect 23438 13682 23490 13694
rect 27806 13746 27858 13758
rect 27806 13682 27858 13694
rect 28478 13746 28530 13758
rect 28478 13682 28530 13694
rect 29038 13746 29090 13758
rect 33070 13746 33122 13758
rect 30146 13694 30158 13746
rect 30210 13694 30222 13746
rect 29038 13682 29090 13694
rect 33070 13682 33122 13694
rect 5966 13634 6018 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 5966 13570 6018 13582
rect 6414 13634 6466 13646
rect 6414 13570 6466 13582
rect 7086 13634 7138 13646
rect 7086 13570 7138 13582
rect 12350 13634 12402 13646
rect 12350 13570 12402 13582
rect 20526 13634 20578 13646
rect 20526 13570 20578 13582
rect 28030 13634 28082 13646
rect 28030 13570 28082 13582
rect 28814 13634 28866 13646
rect 31826 13582 31838 13634
rect 31890 13582 31902 13634
rect 33506 13582 33518 13634
rect 33570 13582 33582 13634
rect 28814 13570 28866 13582
rect 11790 13522 11842 13534
rect 11790 13458 11842 13470
rect 16942 13522 16994 13534
rect 16942 13458 16994 13470
rect 29598 13522 29650 13534
rect 29598 13458 29650 13470
rect 1344 13354 34608 13388
rect 1344 13302 5372 13354
rect 5424 13302 5476 13354
rect 5528 13302 5580 13354
rect 5632 13302 13688 13354
rect 13740 13302 13792 13354
rect 13844 13302 13896 13354
rect 13948 13302 22004 13354
rect 22056 13302 22108 13354
rect 22160 13302 22212 13354
rect 22264 13302 30320 13354
rect 30372 13302 30424 13354
rect 30476 13302 30528 13354
rect 30580 13302 34608 13354
rect 1344 13268 34608 13302
rect 11454 13186 11506 13198
rect 11454 13122 11506 13134
rect 11678 13186 11730 13198
rect 11678 13122 11730 13134
rect 29150 13186 29202 13198
rect 29150 13122 29202 13134
rect 30046 13186 30098 13198
rect 30046 13122 30098 13134
rect 30382 13186 30434 13198
rect 30382 13122 30434 13134
rect 14590 13074 14642 13086
rect 3042 13022 3054 13074
rect 3106 13022 3118 13074
rect 14590 13010 14642 13022
rect 16270 13074 16322 13086
rect 16270 13010 16322 13022
rect 20750 13074 20802 13086
rect 29822 13074 29874 13086
rect 22418 13022 22430 13074
rect 22482 13022 22494 13074
rect 29474 13022 29486 13074
rect 29538 13022 29550 13074
rect 20750 13010 20802 13022
rect 29822 13010 29874 13022
rect 5630 12962 5682 12974
rect 3154 12910 3166 12962
rect 3218 12910 3230 12962
rect 5630 12898 5682 12910
rect 6078 12962 6130 12974
rect 6078 12898 6130 12910
rect 7982 12962 8034 12974
rect 12350 12962 12402 12974
rect 8418 12910 8430 12962
rect 8482 12910 8494 12962
rect 12002 12910 12014 12962
rect 12066 12910 12078 12962
rect 7982 12898 8034 12910
rect 12350 12898 12402 12910
rect 14926 12962 14978 12974
rect 14926 12898 14978 12910
rect 15822 12962 15874 12974
rect 15822 12898 15874 12910
rect 18622 12962 18674 12974
rect 30606 12962 30658 12974
rect 34078 12962 34130 12974
rect 21522 12910 21534 12962
rect 21586 12910 21598 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 23874 12910 23886 12962
rect 23938 12910 23950 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 18622 12898 18674 12910
rect 30606 12898 30658 12910
rect 34078 12898 34130 12910
rect 13470 12850 13522 12862
rect 13470 12786 13522 12798
rect 13806 12850 13858 12862
rect 13806 12786 13858 12798
rect 14478 12850 14530 12862
rect 14478 12786 14530 12798
rect 14814 12850 14866 12862
rect 14814 12786 14866 12798
rect 16046 12850 16098 12862
rect 16046 12786 16098 12798
rect 16382 12850 16434 12862
rect 16382 12786 16434 12798
rect 19630 12850 19682 12862
rect 24670 12850 24722 12862
rect 21298 12798 21310 12850
rect 21362 12798 21374 12850
rect 22642 12798 22654 12850
rect 22706 12798 22718 12850
rect 19630 12786 19682 12798
rect 24670 12786 24722 12798
rect 25790 12850 25842 12862
rect 25790 12786 25842 12798
rect 29374 12850 29426 12862
rect 29374 12786 29426 12798
rect 31390 12850 31442 12862
rect 31390 12786 31442 12798
rect 3278 12738 3330 12750
rect 3278 12674 3330 12686
rect 6190 12738 6242 12750
rect 6190 12674 6242 12686
rect 6302 12738 6354 12750
rect 6302 12674 6354 12686
rect 6862 12738 6914 12750
rect 12126 12738 12178 12750
rect 10882 12686 10894 12738
rect 10946 12686 10958 12738
rect 6862 12674 6914 12686
rect 12126 12674 12178 12686
rect 12238 12738 12290 12750
rect 12238 12674 12290 12686
rect 12910 12738 12962 12750
rect 12910 12674 12962 12686
rect 18734 12738 18786 12750
rect 18734 12674 18786 12686
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 20190 12738 20242 12750
rect 20190 12674 20242 12686
rect 23102 12738 23154 12750
rect 23102 12674 23154 12686
rect 23998 12738 24050 12750
rect 23998 12674 24050 12686
rect 24558 12738 24610 12750
rect 24558 12674 24610 12686
rect 25230 12738 25282 12750
rect 25230 12674 25282 12686
rect 1344 12570 34768 12604
rect 1344 12518 9530 12570
rect 9582 12518 9634 12570
rect 9686 12518 9738 12570
rect 9790 12518 17846 12570
rect 17898 12518 17950 12570
rect 18002 12518 18054 12570
rect 18106 12518 26162 12570
rect 26214 12518 26266 12570
rect 26318 12518 26370 12570
rect 26422 12518 34478 12570
rect 34530 12518 34582 12570
rect 34634 12518 34686 12570
rect 34738 12518 34768 12570
rect 1344 12484 34768 12518
rect 5406 12402 5458 12414
rect 5406 12338 5458 12350
rect 5630 12402 5682 12414
rect 5630 12338 5682 12350
rect 5854 12402 5906 12414
rect 5854 12338 5906 12350
rect 7310 12402 7362 12414
rect 7310 12338 7362 12350
rect 7870 12402 7922 12414
rect 14590 12402 14642 12414
rect 12002 12350 12014 12402
rect 12066 12350 12078 12402
rect 7870 12338 7922 12350
rect 14590 12338 14642 12350
rect 16158 12402 16210 12414
rect 16158 12338 16210 12350
rect 23998 12402 24050 12414
rect 29250 12350 29262 12402
rect 29314 12350 29326 12402
rect 23998 12338 24050 12350
rect 5966 12290 6018 12302
rect 5966 12226 6018 12238
rect 6526 12290 6578 12302
rect 6526 12226 6578 12238
rect 7086 12290 7138 12302
rect 7086 12226 7138 12238
rect 9550 12290 9602 12302
rect 9550 12226 9602 12238
rect 11454 12290 11506 12302
rect 11454 12226 11506 12238
rect 12462 12290 12514 12302
rect 12462 12226 12514 12238
rect 16046 12290 16098 12302
rect 16046 12226 16098 12238
rect 19854 12290 19906 12302
rect 23650 12238 23662 12290
rect 23714 12238 23726 12290
rect 25778 12238 25790 12290
rect 25842 12238 25854 12290
rect 19854 12226 19906 12238
rect 6302 12178 6354 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 2258 12126 2270 12178
rect 2322 12126 2334 12178
rect 4498 12126 4510 12178
rect 4562 12126 4574 12178
rect 6302 12114 6354 12126
rect 6974 12178 7026 12190
rect 6974 12114 7026 12126
rect 7422 12178 7474 12190
rect 7422 12114 7474 12126
rect 9886 12178 9938 12190
rect 9886 12114 9938 12126
rect 11342 12178 11394 12190
rect 11342 12114 11394 12126
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 12350 12178 12402 12190
rect 14702 12178 14754 12190
rect 19406 12178 19458 12190
rect 14466 12126 14478 12178
rect 14530 12126 14542 12178
rect 18946 12126 18958 12178
rect 19010 12126 19022 12178
rect 12350 12114 12402 12126
rect 14702 12114 14754 12126
rect 19406 12114 19458 12126
rect 21086 12178 21138 12190
rect 24558 12178 24610 12190
rect 26910 12178 26962 12190
rect 29598 12178 29650 12190
rect 33630 12178 33682 12190
rect 22306 12126 22318 12178
rect 22370 12126 22382 12178
rect 22866 12126 22878 12178
rect 22930 12126 22942 12178
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 26114 12126 26126 12178
rect 26178 12126 26190 12178
rect 27122 12126 27134 12178
rect 27186 12126 27198 12178
rect 30258 12126 30270 12178
rect 30322 12126 30334 12178
rect 21086 12114 21138 12126
rect 24558 12114 24610 12126
rect 26910 12114 26962 12126
rect 29598 12114 29650 12126
rect 33630 12114 33682 12126
rect 34190 12178 34242 12190
rect 34190 12114 34242 12126
rect 6414 12066 6466 12078
rect 6414 12002 6466 12014
rect 8318 12066 8370 12078
rect 8318 12002 8370 12014
rect 21646 12066 21698 12078
rect 31826 12014 31838 12066
rect 31890 12014 31902 12066
rect 21646 12002 21698 12014
rect 14926 11954 14978 11966
rect 14926 11890 14978 11902
rect 16270 11954 16322 11966
rect 16270 11890 16322 11902
rect 18622 11954 18674 11966
rect 18622 11890 18674 11902
rect 18958 11954 19010 11966
rect 25678 11954 25730 11966
rect 22530 11902 22542 11954
rect 22594 11902 22606 11954
rect 18958 11890 19010 11902
rect 25678 11890 25730 11902
rect 1344 11786 34608 11820
rect 1344 11734 5372 11786
rect 5424 11734 5476 11786
rect 5528 11734 5580 11786
rect 5632 11734 13688 11786
rect 13740 11734 13792 11786
rect 13844 11734 13896 11786
rect 13948 11734 22004 11786
rect 22056 11734 22108 11786
rect 22160 11734 22212 11786
rect 22264 11734 30320 11786
rect 30372 11734 30424 11786
rect 30476 11734 30528 11786
rect 30580 11734 34608 11786
rect 1344 11700 34608 11734
rect 1934 11618 1986 11630
rect 1934 11554 1986 11566
rect 9998 11618 10050 11630
rect 9998 11554 10050 11566
rect 20078 11506 20130 11518
rect 26126 11506 26178 11518
rect 22866 11454 22878 11506
rect 22930 11454 22942 11506
rect 24994 11454 25006 11506
rect 25058 11454 25070 11506
rect 20078 11442 20130 11454
rect 26126 11442 26178 11454
rect 29822 11506 29874 11518
rect 29822 11442 29874 11454
rect 6526 11394 6578 11406
rect 24558 11394 24610 11406
rect 3826 11342 3838 11394
rect 3890 11342 3902 11394
rect 6850 11342 6862 11394
rect 6914 11342 6926 11394
rect 15138 11342 15150 11394
rect 15202 11342 15214 11394
rect 15698 11342 15710 11394
rect 15762 11342 15774 11394
rect 17266 11342 17278 11394
rect 17330 11342 17342 11394
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 19730 11342 19742 11394
rect 19794 11342 19806 11394
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 22082 11342 22094 11394
rect 22146 11342 22158 11394
rect 22418 11342 22430 11394
rect 22482 11342 22494 11394
rect 23538 11342 23550 11394
rect 23602 11342 23614 11394
rect 6526 11330 6578 11342
rect 24558 11330 24610 11342
rect 26686 11394 26738 11406
rect 26686 11330 26738 11342
rect 27022 11394 27074 11406
rect 27022 11330 27074 11342
rect 27582 11394 27634 11406
rect 30706 11342 30718 11394
rect 30770 11342 30782 11394
rect 31154 11342 31166 11394
rect 31218 11342 31230 11394
rect 27582 11330 27634 11342
rect 9214 11282 9266 11294
rect 9214 11218 9266 11230
rect 14590 11282 14642 11294
rect 14590 11218 14642 11230
rect 14814 11282 14866 11294
rect 27918 11282 27970 11294
rect 18610 11230 18622 11282
rect 18674 11230 18686 11282
rect 20402 11230 20414 11282
rect 20466 11230 20478 11282
rect 22978 11230 22990 11282
rect 23042 11230 23054 11282
rect 23874 11230 23886 11282
rect 23938 11230 23950 11282
rect 14814 11218 14866 11230
rect 27918 11218 27970 11230
rect 14702 11170 14754 11182
rect 21422 11170 21474 11182
rect 28254 11170 28306 11182
rect 34302 11170 34354 11182
rect 17602 11118 17614 11170
rect 17666 11118 17678 11170
rect 23426 11118 23438 11170
rect 23490 11118 23502 11170
rect 33506 11118 33518 11170
rect 33570 11118 33582 11170
rect 14702 11106 14754 11118
rect 21422 11106 21474 11118
rect 28254 11106 28306 11118
rect 34302 11106 34354 11118
rect 1344 11002 34768 11036
rect 1344 10950 9530 11002
rect 9582 10950 9634 11002
rect 9686 10950 9738 11002
rect 9790 10950 17846 11002
rect 17898 10950 17950 11002
rect 18002 10950 18054 11002
rect 18106 10950 26162 11002
rect 26214 10950 26266 11002
rect 26318 10950 26370 11002
rect 26422 10950 34478 11002
rect 34530 10950 34582 11002
rect 34634 10950 34686 11002
rect 34738 10950 34768 11002
rect 1344 10916 34768 10950
rect 11678 10834 11730 10846
rect 11678 10770 11730 10782
rect 14814 10834 14866 10846
rect 14814 10770 14866 10782
rect 15486 10834 15538 10846
rect 15486 10770 15538 10782
rect 27358 10834 27410 10846
rect 31390 10834 31442 10846
rect 28018 10782 28030 10834
rect 28082 10782 28094 10834
rect 27358 10770 27410 10782
rect 31390 10770 31442 10782
rect 21422 10722 21474 10734
rect 12562 10670 12574 10722
rect 12626 10670 12638 10722
rect 16370 10670 16382 10722
rect 16434 10670 16446 10722
rect 21422 10658 21474 10670
rect 22878 10722 22930 10734
rect 22878 10658 22930 10670
rect 24558 10722 24610 10734
rect 24558 10658 24610 10670
rect 25566 10722 25618 10734
rect 25566 10658 25618 10670
rect 12014 10610 12066 10622
rect 15822 10610 15874 10622
rect 18846 10610 18898 10622
rect 21870 10610 21922 10622
rect 3826 10558 3838 10610
rect 3890 10558 3902 10610
rect 12786 10558 12798 10610
rect 12850 10558 12862 10610
rect 16594 10558 16606 10610
rect 16658 10558 16670 10610
rect 18050 10558 18062 10610
rect 18114 10558 18126 10610
rect 19058 10558 19070 10610
rect 19122 10558 19134 10610
rect 12014 10546 12066 10558
rect 15822 10546 15874 10558
rect 18846 10546 18898 10558
rect 21870 10546 21922 10558
rect 22318 10610 22370 10622
rect 30830 10610 30882 10622
rect 30370 10558 30382 10610
rect 30434 10558 30446 10610
rect 22318 10546 22370 10558
rect 30830 10546 30882 10558
rect 14254 10498 14306 10510
rect 18386 10446 18398 10498
rect 18450 10446 18462 10498
rect 20626 10446 20638 10498
rect 20690 10446 20702 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 26002 10446 26014 10498
rect 26066 10446 26078 10498
rect 14254 10434 14306 10446
rect 1934 10386 1986 10398
rect 24334 10386 24386 10398
rect 18946 10334 18958 10386
rect 19010 10334 19022 10386
rect 1934 10322 1986 10334
rect 24334 10322 24386 10334
rect 1344 10218 34608 10252
rect 1344 10166 5372 10218
rect 5424 10166 5476 10218
rect 5528 10166 5580 10218
rect 5632 10166 13688 10218
rect 13740 10166 13792 10218
rect 13844 10166 13896 10218
rect 13948 10166 22004 10218
rect 22056 10166 22108 10218
rect 22160 10166 22212 10218
rect 22264 10166 30320 10218
rect 30372 10166 30424 10218
rect 30476 10166 30528 10218
rect 30580 10166 34608 10218
rect 1344 10132 34608 10166
rect 2158 10050 2210 10062
rect 2158 9986 2210 9998
rect 3390 10050 3442 10062
rect 17390 10050 17442 10062
rect 14690 9998 14702 10050
rect 14754 9998 14766 10050
rect 3390 9986 3442 9998
rect 17390 9986 17442 9998
rect 17726 10050 17778 10062
rect 25554 9998 25566 10050
rect 25618 9998 25630 10050
rect 33506 9998 33518 10050
rect 33570 9998 33582 10050
rect 17726 9986 17778 9998
rect 3278 9938 3330 9950
rect 3278 9874 3330 9886
rect 3838 9938 3890 9950
rect 3838 9874 3890 9886
rect 12238 9938 12290 9950
rect 12238 9874 12290 9886
rect 14142 9938 14194 9950
rect 16482 9886 16494 9938
rect 16546 9886 16558 9938
rect 21746 9886 21758 9938
rect 21810 9886 21822 9938
rect 14142 9874 14194 9886
rect 6862 9826 6914 9838
rect 2706 9774 2718 9826
rect 2770 9774 2782 9826
rect 6862 9762 6914 9774
rect 7982 9826 8034 9838
rect 7982 9762 8034 9774
rect 8542 9826 8594 9838
rect 14814 9826 14866 9838
rect 9202 9774 9214 9826
rect 9266 9774 9278 9826
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 8542 9762 8594 9774
rect 14814 9762 14866 9774
rect 14926 9826 14978 9838
rect 18286 9826 18338 9838
rect 16594 9774 16606 9826
rect 16658 9774 16670 9826
rect 14926 9762 14978 9774
rect 18286 9762 18338 9774
rect 20750 9826 20802 9838
rect 22990 9826 23042 9838
rect 26350 9826 26402 9838
rect 22530 9774 22542 9826
rect 22594 9774 22606 9826
rect 25218 9774 25230 9826
rect 25282 9774 25294 9826
rect 26674 9774 26686 9826
rect 26738 9774 26750 9826
rect 31826 9774 31838 9826
rect 31890 9774 31902 9826
rect 20750 9762 20802 9774
rect 22990 9762 23042 9774
rect 26350 9762 26402 9774
rect 2270 9714 2322 9726
rect 7086 9714 7138 9726
rect 2930 9662 2942 9714
rect 2994 9662 3006 9714
rect 2270 9650 2322 9662
rect 7086 9650 7138 9662
rect 14254 9714 14306 9726
rect 14254 9650 14306 9662
rect 16270 9714 16322 9726
rect 16270 9650 16322 9662
rect 17950 9714 18002 9726
rect 20302 9714 20354 9726
rect 18610 9662 18622 9714
rect 18674 9662 18686 9714
rect 17950 9650 18002 9662
rect 20302 9650 20354 9662
rect 22766 9714 22818 9726
rect 23090 9662 23102 9714
rect 23154 9662 23166 9714
rect 23874 9662 23886 9714
rect 23938 9662 23950 9714
rect 25106 9662 25118 9714
rect 25170 9662 25182 9714
rect 22766 9650 22818 9662
rect 7534 9602 7586 9614
rect 14030 9602 14082 9614
rect 6514 9550 6526 9602
rect 6578 9550 6590 9602
rect 8306 9550 8318 9602
rect 8370 9550 8382 9602
rect 11442 9550 11454 9602
rect 11506 9550 11518 9602
rect 12786 9550 12798 9602
rect 12850 9550 12862 9602
rect 7534 9538 7586 9550
rect 14030 9538 14082 9550
rect 20526 9602 20578 9614
rect 20526 9538 20578 9550
rect 20638 9602 20690 9614
rect 20638 9538 20690 9550
rect 1344 9434 34768 9468
rect 1344 9382 9530 9434
rect 9582 9382 9634 9434
rect 9686 9382 9738 9434
rect 9790 9382 17846 9434
rect 17898 9382 17950 9434
rect 18002 9382 18054 9434
rect 18106 9382 26162 9434
rect 26214 9382 26266 9434
rect 26318 9382 26370 9434
rect 26422 9382 34478 9434
rect 34530 9382 34582 9434
rect 34634 9382 34686 9434
rect 34738 9382 34768 9434
rect 1344 9348 34768 9382
rect 6862 9266 6914 9278
rect 5954 9214 5966 9266
rect 6018 9214 6030 9266
rect 6862 9202 6914 9214
rect 28702 9266 28754 9278
rect 32622 9266 32674 9278
rect 32050 9214 32062 9266
rect 32114 9214 32126 9266
rect 33170 9214 33182 9266
rect 33234 9214 33246 9266
rect 28702 9202 28754 9214
rect 32622 9202 32674 9214
rect 6526 9154 6578 9166
rect 17502 9154 17554 9166
rect 27246 9154 27298 9166
rect 16706 9102 16718 9154
rect 16770 9102 16782 9154
rect 18722 9102 18734 9154
rect 18786 9102 18798 9154
rect 22866 9102 22878 9154
rect 22930 9102 22942 9154
rect 6526 9090 6578 9102
rect 17502 9090 17554 9102
rect 27246 9090 27298 9102
rect 33854 9154 33906 9166
rect 33854 9090 33906 9102
rect 2270 9042 2322 9054
rect 2270 8978 2322 8990
rect 3054 9042 3106 9054
rect 6750 9042 6802 9054
rect 3490 8990 3502 9042
rect 3554 8990 3566 9042
rect 3054 8978 3106 8990
rect 6750 8978 6802 8990
rect 7086 9042 7138 9054
rect 7086 8978 7138 8990
rect 7198 9042 7250 9054
rect 21086 9042 21138 9054
rect 15250 8990 15262 9042
rect 15314 8990 15326 9042
rect 15810 8990 15822 9042
rect 15874 8990 15886 9042
rect 16482 8990 16494 9042
rect 16546 8990 16558 9042
rect 19170 8990 19182 9042
rect 19234 8990 19246 9042
rect 20514 8990 20526 9042
rect 20578 8990 20590 9042
rect 7198 8978 7250 8990
rect 21086 8978 21138 8990
rect 24558 9042 24610 9054
rect 28926 9042 28978 9054
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 26114 8990 26126 9042
rect 26178 8990 26190 9042
rect 28466 8990 28478 9042
rect 28530 8990 28542 9042
rect 29474 8990 29486 9042
rect 29538 8990 29550 9042
rect 33394 8990 33406 9042
rect 33458 8990 33470 9042
rect 34066 8990 34078 9042
rect 34130 8990 34142 9042
rect 24558 8978 24610 8990
rect 28926 8978 28978 8990
rect 7758 8930 7810 8942
rect 17390 8930 17442 8942
rect 20302 8930 20354 8942
rect 24334 8930 24386 8942
rect 1810 8878 1822 8930
rect 1874 8878 1886 8930
rect 16594 8878 16606 8930
rect 16658 8878 16670 8930
rect 19282 8878 19294 8930
rect 19346 8878 19358 8930
rect 22530 8878 22542 8930
rect 22594 8878 22606 8930
rect 25778 8878 25790 8930
rect 25842 8878 25854 8930
rect 7758 8866 7810 8878
rect 17390 8866 17442 8878
rect 20302 8866 20354 8878
rect 24334 8866 24386 8878
rect 21310 8818 21362 8830
rect 24222 8818 24274 8830
rect 20178 8766 20190 8818
rect 20242 8766 20254 8818
rect 22642 8766 22654 8818
rect 22706 8766 22718 8818
rect 21310 8754 21362 8766
rect 24222 8754 24274 8766
rect 24670 8818 24722 8830
rect 26450 8766 26462 8818
rect 26514 8766 26526 8818
rect 24670 8754 24722 8766
rect 1344 8650 34608 8684
rect 1344 8598 5372 8650
rect 5424 8598 5476 8650
rect 5528 8598 5580 8650
rect 5632 8598 13688 8650
rect 13740 8598 13792 8650
rect 13844 8598 13896 8650
rect 13948 8598 22004 8650
rect 22056 8598 22108 8650
rect 22160 8598 22212 8650
rect 22264 8598 30320 8650
rect 30372 8598 30424 8650
rect 30476 8598 30528 8650
rect 30580 8598 34608 8650
rect 1344 8564 34608 8598
rect 33966 8482 34018 8494
rect 33966 8418 34018 8430
rect 1934 8370 1986 8382
rect 6414 8370 6466 8382
rect 6066 8318 6078 8370
rect 6130 8318 6142 8370
rect 1934 8306 1986 8318
rect 6414 8306 6466 8318
rect 14030 8370 14082 8382
rect 14030 8306 14082 8318
rect 25790 8370 25842 8382
rect 25790 8306 25842 8318
rect 27022 8370 27074 8382
rect 27022 8306 27074 8318
rect 29262 8370 29314 8382
rect 29262 8306 29314 8318
rect 29598 8370 29650 8382
rect 29598 8306 29650 8318
rect 13470 8258 13522 8270
rect 14478 8258 14530 8270
rect 3826 8206 3838 8258
rect 3890 8206 3902 8258
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 13470 8194 13522 8206
rect 14478 8194 14530 8206
rect 14814 8258 14866 8270
rect 20302 8258 20354 8270
rect 16706 8206 16718 8258
rect 16770 8206 16782 8258
rect 17042 8206 17054 8258
rect 17106 8206 17118 8258
rect 18274 8206 18286 8258
rect 18338 8206 18350 8258
rect 14814 8194 14866 8206
rect 20302 8194 20354 8206
rect 22094 8258 22146 8270
rect 25902 8258 25954 8270
rect 22642 8206 22654 8258
rect 22706 8206 22718 8258
rect 22094 8194 22146 8206
rect 25902 8194 25954 8206
rect 26238 8258 26290 8270
rect 26238 8194 26290 8206
rect 26462 8258 26514 8270
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 26462 8194 26514 8206
rect 12462 8146 12514 8158
rect 4610 8094 4622 8146
rect 4674 8094 4686 8146
rect 12462 8082 12514 8094
rect 12798 8146 12850 8158
rect 12798 8082 12850 8094
rect 14702 8146 14754 8158
rect 31278 8146 31330 8158
rect 15586 8094 15598 8146
rect 15650 8094 15662 8146
rect 29810 8094 29822 8146
rect 29874 8094 29886 8146
rect 30146 8094 30158 8146
rect 30210 8094 30222 8146
rect 14702 8082 14754 8094
rect 31278 8082 31330 8094
rect 4958 8034 5010 8046
rect 4958 7970 5010 7982
rect 6190 8034 6242 8046
rect 11230 8034 11282 8046
rect 10882 7982 10894 8034
rect 10946 7982 10958 8034
rect 6190 7970 6242 7982
rect 11230 7970 11282 7982
rect 12910 8034 12962 8046
rect 12910 7970 12962 7982
rect 13918 8034 13970 8046
rect 13918 7970 13970 7982
rect 14142 8034 14194 8046
rect 14142 7970 14194 7982
rect 15262 8034 15314 8046
rect 15262 7970 15314 7982
rect 19294 8034 19346 8046
rect 19294 7970 19346 7982
rect 19518 8034 19570 8046
rect 19518 7970 19570 7982
rect 19630 8034 19682 8046
rect 19630 7970 19682 7982
rect 19742 8034 19794 8046
rect 19742 7970 19794 7982
rect 20638 8034 20690 8046
rect 26238 8034 26290 8046
rect 25218 7982 25230 8034
rect 25282 7982 25294 8034
rect 20638 7970 20690 7982
rect 26238 7970 26290 7982
rect 30942 8034 30994 8046
rect 30942 7970 30994 7982
rect 1344 7866 34768 7900
rect 1344 7814 9530 7866
rect 9582 7814 9634 7866
rect 9686 7814 9738 7866
rect 9790 7814 17846 7866
rect 17898 7814 17950 7866
rect 18002 7814 18054 7866
rect 18106 7814 26162 7866
rect 26214 7814 26266 7866
rect 26318 7814 26370 7866
rect 26422 7814 34478 7866
rect 34530 7814 34582 7866
rect 34634 7814 34686 7866
rect 34738 7814 34768 7866
rect 1344 7780 34768 7814
rect 6078 7698 6130 7710
rect 12126 7698 12178 7710
rect 4834 7646 4846 7698
rect 4898 7646 4910 7698
rect 6626 7646 6638 7698
rect 6690 7646 6702 7698
rect 6078 7634 6130 7646
rect 12126 7634 12178 7646
rect 13022 7698 13074 7710
rect 13022 7634 13074 7646
rect 17726 7698 17778 7710
rect 17726 7634 17778 7646
rect 21310 7698 21362 7710
rect 21310 7634 21362 7646
rect 22542 7698 22594 7710
rect 22542 7634 22594 7646
rect 25790 7698 25842 7710
rect 25790 7634 25842 7646
rect 26798 7698 26850 7710
rect 33630 7698 33682 7710
rect 29586 7646 29598 7698
rect 29650 7646 29662 7698
rect 26798 7634 26850 7646
rect 33630 7634 33682 7646
rect 5966 7586 6018 7598
rect 5966 7522 6018 7534
rect 7198 7586 7250 7598
rect 7198 7522 7250 7534
rect 12014 7586 12066 7598
rect 21198 7586 21250 7598
rect 15138 7534 15150 7586
rect 15202 7534 15214 7586
rect 17378 7534 17390 7586
rect 17442 7534 17454 7586
rect 12014 7522 12066 7534
rect 21198 7522 21250 7534
rect 23326 7586 23378 7598
rect 23326 7522 23378 7534
rect 26574 7586 26626 7598
rect 26574 7522 26626 7534
rect 27022 7586 27074 7598
rect 27022 7522 27074 7534
rect 27358 7586 27410 7598
rect 28702 7586 28754 7598
rect 27682 7534 27694 7586
rect 27746 7534 27758 7586
rect 27358 7522 27410 7534
rect 28702 7522 28754 7534
rect 2046 7474 2098 7486
rect 5518 7474 5570 7486
rect 2482 7422 2494 7474
rect 2546 7422 2558 7474
rect 2046 7410 2098 7422
rect 5518 7410 5570 7422
rect 5854 7474 5906 7486
rect 5854 7410 5906 7422
rect 6414 7474 6466 7486
rect 6414 7410 6466 7422
rect 6974 7474 7026 7486
rect 13246 7474 13298 7486
rect 12898 7422 12910 7474
rect 12962 7422 12974 7474
rect 6974 7410 7026 7422
rect 13246 7410 13298 7422
rect 15486 7474 15538 7486
rect 21534 7474 21586 7486
rect 19394 7422 19406 7474
rect 19458 7422 19470 7474
rect 15486 7410 15538 7422
rect 21534 7410 21586 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 22654 7474 22706 7486
rect 22654 7410 22706 7422
rect 22878 7474 22930 7486
rect 22878 7410 22930 7422
rect 23214 7474 23266 7486
rect 29262 7474 29314 7486
rect 28466 7422 28478 7474
rect 28530 7422 28542 7474
rect 29922 7422 29934 7474
rect 29986 7422 29998 7474
rect 23214 7410 23266 7422
rect 29262 7410 29314 7422
rect 13134 7362 13186 7374
rect 13134 7298 13186 7310
rect 18958 7362 19010 7374
rect 18958 7298 19010 7310
rect 26126 7362 26178 7374
rect 26126 7298 26178 7310
rect 29038 7362 29090 7374
rect 33406 7362 33458 7374
rect 31826 7310 31838 7362
rect 31890 7310 31902 7362
rect 29038 7298 29090 7310
rect 33406 7298 33458 7310
rect 34190 7362 34242 7374
rect 34190 7298 34242 7310
rect 12574 7250 12626 7262
rect 12574 7186 12626 7198
rect 27134 7250 27186 7262
rect 27134 7186 27186 7198
rect 1344 7082 34608 7116
rect 1344 7030 5372 7082
rect 5424 7030 5476 7082
rect 5528 7030 5580 7082
rect 5632 7030 13688 7082
rect 13740 7030 13792 7082
rect 13844 7030 13896 7082
rect 13948 7030 22004 7082
rect 22056 7030 22108 7082
rect 22160 7030 22212 7082
rect 22264 7030 30320 7082
rect 30372 7030 30424 7082
rect 30476 7030 30528 7082
rect 30580 7030 34608 7082
rect 1344 6996 34608 7030
rect 5630 6914 5682 6926
rect 4834 6862 4846 6914
rect 4898 6911 4910 6914
rect 4898 6865 5007 6911
rect 4898 6862 4910 6865
rect 4734 6690 4786 6702
rect 4050 6638 4062 6690
rect 4114 6638 4126 6690
rect 4961 6687 5007 6865
rect 5630 6850 5682 6862
rect 5966 6914 6018 6926
rect 5966 6850 6018 6862
rect 16382 6914 16434 6926
rect 16382 6850 16434 6862
rect 19518 6914 19570 6926
rect 19518 6850 19570 6862
rect 29598 6802 29650 6814
rect 6290 6750 6302 6802
rect 6354 6750 6366 6802
rect 28242 6750 28254 6802
rect 28306 6750 28318 6802
rect 29598 6738 29650 6750
rect 29822 6802 29874 6814
rect 29822 6738 29874 6750
rect 7758 6690 7810 6702
rect 11454 6690 11506 6702
rect 22542 6690 22594 6702
rect 5170 6687 5182 6690
rect 4961 6641 5182 6687
rect 5170 6638 5182 6641
rect 5234 6638 5246 6690
rect 8418 6638 8430 6690
rect 8482 6638 8494 6690
rect 20066 6638 20078 6690
rect 20130 6638 20142 6690
rect 4734 6626 4786 6638
rect 7758 6626 7810 6638
rect 11454 6626 11506 6638
rect 22542 6626 22594 6638
rect 22878 6690 22930 6702
rect 22878 6626 22930 6638
rect 26462 6690 26514 6702
rect 26462 6626 26514 6638
rect 26798 6690 26850 6702
rect 26798 6626 26850 6638
rect 26910 6690 26962 6702
rect 26910 6626 26962 6638
rect 27246 6690 27298 6702
rect 27246 6626 27298 6638
rect 27918 6690 27970 6702
rect 27918 6626 27970 6638
rect 29374 6690 29426 6702
rect 29374 6626 29426 6638
rect 30158 6690 30210 6702
rect 30158 6626 30210 6638
rect 30606 6690 30658 6702
rect 31154 6638 31166 6690
rect 31218 6638 31230 6690
rect 30606 6626 30658 6638
rect 6638 6578 6690 6590
rect 23214 6578 23266 6590
rect 2482 6526 2494 6578
rect 2546 6526 2558 6578
rect 16594 6526 16606 6578
rect 16658 6526 16670 6578
rect 16930 6526 16942 6578
rect 16994 6526 17006 6578
rect 20178 6526 20190 6578
rect 20242 6526 20254 6578
rect 6638 6514 6690 6526
rect 23214 6514 23266 6526
rect 26574 6578 26626 6590
rect 26574 6514 26626 6526
rect 28590 6578 28642 6590
rect 28590 6514 28642 6526
rect 30046 6578 30098 6590
rect 30046 6514 30098 6526
rect 30270 6578 30322 6590
rect 30270 6514 30322 6526
rect 33518 6578 33570 6590
rect 33518 6514 33570 6526
rect 5742 6466 5794 6478
rect 5742 6402 5794 6414
rect 6414 6466 6466 6478
rect 16046 6466 16098 6478
rect 10658 6414 10670 6466
rect 10722 6414 10734 6466
rect 6414 6402 6466 6414
rect 16046 6402 16098 6414
rect 19182 6466 19234 6478
rect 19182 6402 19234 6414
rect 22766 6466 22818 6478
rect 22766 6402 22818 6414
rect 27694 6466 27746 6478
rect 27694 6402 27746 6414
rect 27806 6466 27858 6478
rect 27806 6402 27858 6414
rect 28366 6466 28418 6478
rect 28366 6402 28418 6414
rect 34302 6466 34354 6478
rect 34302 6402 34354 6414
rect 1344 6298 34768 6332
rect 1344 6246 9530 6298
rect 9582 6246 9634 6298
rect 9686 6246 9738 6298
rect 9790 6246 17846 6298
rect 17898 6246 17950 6298
rect 18002 6246 18054 6298
rect 18106 6246 26162 6298
rect 26214 6246 26266 6298
rect 26318 6246 26370 6298
rect 26422 6246 34478 6298
rect 34530 6246 34582 6298
rect 34634 6246 34686 6298
rect 34738 6246 34768 6298
rect 1344 6212 34768 6246
rect 6638 6130 6690 6142
rect 5170 6078 5182 6130
rect 5234 6078 5246 6130
rect 6638 6066 6690 6078
rect 8318 6130 8370 6142
rect 8318 6066 8370 6078
rect 9662 6130 9714 6142
rect 9662 6066 9714 6078
rect 12798 6130 12850 6142
rect 12798 6066 12850 6078
rect 13694 6130 13746 6142
rect 13694 6066 13746 6078
rect 16494 6130 16546 6142
rect 16494 6066 16546 6078
rect 17726 6130 17778 6142
rect 17726 6066 17778 6078
rect 19518 6130 19570 6142
rect 19518 6066 19570 6078
rect 20078 6130 20130 6142
rect 20078 6066 20130 6078
rect 25902 6130 25954 6142
rect 25902 6066 25954 6078
rect 31054 6130 31106 6142
rect 33182 6130 33234 6142
rect 31826 6078 31838 6130
rect 31890 6078 31902 6130
rect 32162 6078 32174 6130
rect 32226 6078 32238 6130
rect 31054 6066 31106 6078
rect 33182 6066 33234 6078
rect 34190 6130 34242 6142
rect 34190 6066 34242 6078
rect 12126 6018 12178 6030
rect 12126 5954 12178 5966
rect 14814 6018 14866 6030
rect 14814 5954 14866 5966
rect 15150 6018 15202 6030
rect 15150 5954 15202 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 18174 6018 18226 6030
rect 31166 6018 31218 6030
rect 28690 5966 28702 6018
rect 28754 5966 28766 6018
rect 18174 5954 18226 5966
rect 31166 5954 31218 5966
rect 2270 5906 2322 5918
rect 5966 5906 6018 5918
rect 2930 5854 2942 5906
rect 2994 5854 3006 5906
rect 2270 5842 2322 5854
rect 5966 5842 6018 5854
rect 6190 5906 6242 5918
rect 6190 5842 6242 5854
rect 6526 5906 6578 5918
rect 6526 5842 6578 5854
rect 6862 5906 6914 5918
rect 11118 5906 11170 5918
rect 12574 5906 12626 5918
rect 8530 5854 8542 5906
rect 8594 5854 8606 5906
rect 11554 5854 11566 5906
rect 11618 5854 11630 5906
rect 6862 5842 6914 5854
rect 11118 5842 11170 5854
rect 12574 5842 12626 5854
rect 13022 5906 13074 5918
rect 13022 5842 13074 5854
rect 13246 5906 13298 5918
rect 13246 5842 13298 5854
rect 13918 5906 13970 5918
rect 15486 5906 15538 5918
rect 20414 5906 20466 5918
rect 31502 5906 31554 5918
rect 33630 5906 33682 5918
rect 14018 5854 14030 5906
rect 14082 5854 14094 5906
rect 15922 5854 15934 5906
rect 15986 5854 15998 5906
rect 16706 5854 16718 5906
rect 16770 5854 16782 5906
rect 18610 5854 18622 5906
rect 18674 5854 18686 5906
rect 29586 5854 29598 5906
rect 29650 5854 29662 5906
rect 30034 5854 30046 5906
rect 30098 5854 30110 5906
rect 32386 5854 32398 5906
rect 32450 5854 32462 5906
rect 13918 5842 13970 5854
rect 15486 5842 15538 5854
rect 20414 5842 20466 5854
rect 31502 5842 31554 5854
rect 33630 5842 33682 5854
rect 7198 5794 7250 5806
rect 7198 5730 7250 5742
rect 12014 5794 12066 5806
rect 12014 5730 12066 5742
rect 12686 5794 12738 5806
rect 12686 5730 12738 5742
rect 13806 5794 13858 5806
rect 18946 5742 18958 5794
rect 19010 5742 19022 5794
rect 19394 5742 19406 5794
rect 19458 5742 19470 5794
rect 28802 5742 28814 5794
rect 28866 5742 28878 5794
rect 13806 5730 13858 5742
rect 9550 5682 9602 5694
rect 9550 5618 9602 5630
rect 9886 5682 9938 5694
rect 9886 5618 9938 5630
rect 14366 5682 14418 5694
rect 14366 5618 14418 5630
rect 14702 5682 14754 5694
rect 14702 5618 14754 5630
rect 19742 5682 19794 5694
rect 19742 5618 19794 5630
rect 1344 5514 34608 5548
rect 1344 5462 5372 5514
rect 5424 5462 5476 5514
rect 5528 5462 5580 5514
rect 5632 5462 13688 5514
rect 13740 5462 13792 5514
rect 13844 5462 13896 5514
rect 13948 5462 22004 5514
rect 22056 5462 22108 5514
rect 22160 5462 22212 5514
rect 22264 5462 30320 5514
rect 30372 5462 30424 5514
rect 30476 5462 30528 5514
rect 30580 5462 34608 5514
rect 1344 5428 34608 5462
rect 5742 5346 5794 5358
rect 5742 5282 5794 5294
rect 6078 5346 6130 5358
rect 6078 5282 6130 5294
rect 11678 5346 11730 5358
rect 11678 5282 11730 5294
rect 13582 5346 13634 5358
rect 13582 5282 13634 5294
rect 19742 5346 19794 5358
rect 19742 5282 19794 5294
rect 25790 5346 25842 5358
rect 25790 5282 25842 5294
rect 29262 5346 29314 5358
rect 29262 5282 29314 5294
rect 4734 5234 4786 5246
rect 4734 5170 4786 5182
rect 6302 5234 6354 5246
rect 6302 5170 6354 5182
rect 6750 5234 6802 5246
rect 6750 5170 6802 5182
rect 20302 5234 20354 5246
rect 20302 5170 20354 5182
rect 29374 5234 29426 5246
rect 29374 5170 29426 5182
rect 30046 5234 30098 5246
rect 30046 5170 30098 5182
rect 33630 5234 33682 5246
rect 33630 5170 33682 5182
rect 7758 5122 7810 5134
rect 4274 5070 4286 5122
rect 4338 5070 4350 5122
rect 7758 5058 7810 5070
rect 8206 5122 8258 5134
rect 16046 5122 16098 5134
rect 22318 5122 22370 5134
rect 34190 5122 34242 5134
rect 8642 5070 8654 5122
rect 8706 5070 8718 5122
rect 16594 5070 16606 5122
rect 16658 5070 16670 5122
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 29586 5070 29598 5122
rect 29650 5070 29662 5122
rect 30706 5070 30718 5122
rect 30770 5070 30782 5122
rect 8206 5058 8258 5070
rect 16046 5058 16098 5070
rect 22318 5058 22370 5070
rect 34190 5058 34242 5070
rect 7422 5010 7474 5022
rect 7422 4946 7474 4958
rect 13470 5010 13522 5022
rect 13470 4946 13522 4958
rect 29934 5010 29986 5022
rect 29934 4946 29986 4958
rect 3278 4898 3330 4910
rect 3278 4834 3330 4846
rect 4622 4898 4674 4910
rect 27582 4898 27634 4910
rect 11106 4846 11118 4898
rect 11170 4846 11182 4898
rect 18946 4846 18958 4898
rect 19010 4846 19022 4898
rect 25106 4846 25118 4898
rect 25170 4846 25182 4898
rect 4622 4834 4674 4846
rect 27582 4834 27634 4846
rect 31726 4898 31778 4910
rect 31726 4834 31778 4846
rect 1344 4730 34768 4764
rect 1344 4678 9530 4730
rect 9582 4678 9634 4730
rect 9686 4678 9738 4730
rect 9790 4678 17846 4730
rect 17898 4678 17950 4730
rect 18002 4678 18054 4730
rect 18106 4678 26162 4730
rect 26214 4678 26266 4730
rect 26318 4678 26370 4730
rect 26422 4678 34478 4730
rect 34530 4678 34582 4730
rect 34634 4678 34686 4730
rect 34738 4678 34768 4730
rect 1344 4644 34768 4678
rect 10782 4562 10834 4574
rect 8530 4510 8542 4562
rect 8594 4510 8606 4562
rect 10782 4498 10834 4510
rect 13134 4562 13186 4574
rect 18622 4562 18674 4574
rect 22654 4562 22706 4574
rect 13682 4510 13694 4562
rect 13746 4510 13758 4562
rect 19394 4510 19406 4562
rect 19458 4510 19470 4562
rect 13134 4498 13186 4510
rect 18622 4498 18674 4510
rect 22654 4498 22706 4510
rect 23998 4562 24050 4574
rect 23998 4498 24050 4510
rect 25678 4562 25730 4574
rect 29934 4562 29986 4574
rect 29362 4510 29374 4562
rect 29426 4510 29438 4562
rect 25678 4498 25730 4510
rect 29934 4498 29986 4510
rect 30494 4562 30546 4574
rect 30494 4498 30546 4510
rect 30942 4562 30994 4574
rect 30942 4498 30994 4510
rect 32174 4562 32226 4574
rect 32174 4498 32226 4510
rect 33854 4562 33906 4574
rect 33854 4498 33906 4510
rect 10670 4450 10722 4462
rect 10670 4386 10722 4398
rect 11006 4450 11058 4462
rect 11006 4386 11058 4398
rect 12126 4450 12178 4462
rect 12126 4386 12178 4398
rect 17502 4450 17554 4462
rect 17502 4386 17554 4398
rect 18398 4450 18450 4462
rect 18398 4386 18450 4398
rect 23438 4450 23490 4462
rect 23438 4386 23490 4398
rect 25902 4450 25954 4462
rect 25902 4386 25954 4398
rect 33182 4450 33234 4462
rect 33182 4386 33234 4398
rect 4622 4338 4674 4350
rect 3938 4286 3950 4338
rect 4002 4286 4014 4338
rect 4622 4274 4674 4286
rect 5182 4338 5234 4350
rect 5182 4274 5234 4286
rect 5630 4338 5682 4350
rect 9102 4338 9154 4350
rect 11118 4338 11170 4350
rect 5954 4286 5966 4338
rect 6018 4286 6030 4338
rect 10210 4286 10222 4338
rect 10274 4286 10286 4338
rect 5630 4274 5682 4286
rect 9102 4274 9154 4286
rect 11118 4274 11170 4286
rect 11902 4338 11954 4350
rect 22318 4338 22370 4350
rect 16146 4286 16158 4338
rect 16210 4286 16222 4338
rect 16706 4286 16718 4338
rect 16770 4286 16782 4338
rect 18162 4286 18174 4338
rect 18226 4286 18238 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 11902 4274 11954 4286
rect 22318 4274 22370 4286
rect 26462 4338 26514 4350
rect 30382 4338 30434 4350
rect 26898 4286 26910 4338
rect 26962 4286 26974 4338
rect 26462 4274 26514 4286
rect 30382 4274 30434 4286
rect 32622 4338 32674 4350
rect 34066 4286 34078 4338
rect 34130 4286 34142 4338
rect 32622 4274 32674 4286
rect 11566 4226 11618 4238
rect 9874 4174 9886 4226
rect 9938 4174 9950 4226
rect 11566 4162 11618 4174
rect 33070 4226 33122 4238
rect 33070 4162 33122 4174
rect 1934 4114 1986 4126
rect 1934 4050 1986 4062
rect 17390 4114 17442 4126
rect 17390 4050 17442 4062
rect 23550 4114 23602 4126
rect 23550 4050 23602 4062
rect 26014 4114 26066 4126
rect 26014 4050 26066 4062
rect 1344 3946 34608 3980
rect 1344 3894 5372 3946
rect 5424 3894 5476 3946
rect 5528 3894 5580 3946
rect 5632 3894 13688 3946
rect 13740 3894 13792 3946
rect 13844 3894 13896 3946
rect 13948 3894 22004 3946
rect 22056 3894 22108 3946
rect 22160 3894 22212 3946
rect 22264 3894 30320 3946
rect 30372 3894 30424 3946
rect 30476 3894 30528 3946
rect 30580 3894 34608 3946
rect 1344 3860 34608 3894
rect 2270 3666 2322 3678
rect 2270 3602 2322 3614
rect 8878 3666 8930 3678
rect 8878 3602 8930 3614
rect 10334 3666 10386 3678
rect 10334 3602 10386 3614
rect 12686 3666 12738 3678
rect 12686 3602 12738 3614
rect 14142 3666 14194 3678
rect 14142 3602 14194 3614
rect 19966 3666 20018 3678
rect 25566 3666 25618 3678
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 19966 3602 20018 3614
rect 25566 3602 25618 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 32958 3666 33010 3678
rect 32958 3602 33010 3614
rect 20078 3554 20130 3566
rect 31726 3554 31778 3566
rect 4610 3502 4622 3554
rect 4674 3502 4686 3554
rect 5954 3502 5966 3554
rect 6018 3502 6030 3554
rect 9314 3502 9326 3554
rect 9378 3502 9390 3554
rect 13122 3502 13134 3554
rect 13186 3502 13198 3554
rect 17378 3502 17390 3554
rect 17442 3502 17454 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 33282 3502 33294 3554
rect 33346 3502 33358 3554
rect 20078 3490 20130 3502
rect 31726 3490 31778 3502
rect 32510 3442 32562 3454
rect 18498 3390 18510 3442
rect 18562 3390 18574 3442
rect 32510 3378 32562 3390
rect 33518 3442 33570 3454
rect 33518 3378 33570 3390
rect 33854 3442 33906 3454
rect 33854 3378 33906 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 6638 3330 6690 3342
rect 6638 3266 6690 3278
rect 1344 3162 34768 3196
rect 1344 3110 9530 3162
rect 9582 3110 9634 3162
rect 9686 3110 9738 3162
rect 9790 3110 17846 3162
rect 17898 3110 17950 3162
rect 18002 3110 18054 3162
rect 18106 3110 26162 3162
rect 26214 3110 26266 3162
rect 26318 3110 26370 3162
rect 26422 3110 34478 3162
rect 34530 3110 34582 3162
rect 34634 3110 34686 3162
rect 34738 3110 34768 3162
rect 1344 3076 34768 3110
<< via1 >>
rect 5372 22710 5424 22762
rect 5476 22710 5528 22762
rect 5580 22710 5632 22762
rect 13688 22710 13740 22762
rect 13792 22710 13844 22762
rect 13896 22710 13948 22762
rect 22004 22710 22056 22762
rect 22108 22710 22160 22762
rect 22212 22710 22264 22762
rect 30320 22710 30372 22762
rect 30424 22710 30476 22762
rect 30528 22710 30580 22762
rect 2270 22542 2322 22594
rect 6638 22542 6690 22594
rect 9550 22542 9602 22594
rect 14142 22542 14194 22594
rect 17166 22542 17218 22594
rect 20974 22542 21026 22594
rect 25566 22542 25618 22594
rect 28590 22542 28642 22594
rect 4174 22318 4226 22370
rect 5966 22318 6018 22370
rect 11454 22318 11506 22370
rect 13134 22318 13186 22370
rect 19070 22318 19122 22370
rect 23326 22318 23378 22370
rect 24558 22318 24610 22370
rect 27806 22318 27858 22370
rect 30942 22318 30994 22370
rect 27470 22206 27522 22258
rect 19966 22094 20018 22146
rect 23774 22094 23826 22146
rect 27582 22094 27634 22146
rect 31390 22094 31442 22146
rect 9530 21926 9582 21978
rect 9634 21926 9686 21978
rect 9738 21926 9790 21978
rect 17846 21926 17898 21978
rect 17950 21926 18002 21978
rect 18054 21926 18106 21978
rect 26162 21926 26214 21978
rect 26266 21926 26318 21978
rect 26370 21926 26422 21978
rect 34478 21926 34530 21978
rect 34582 21926 34634 21978
rect 34686 21926 34738 21978
rect 10334 21758 10386 21810
rect 10670 21758 10722 21810
rect 11006 21758 11058 21810
rect 12574 21758 12626 21810
rect 12910 21758 12962 21810
rect 17390 21758 17442 21810
rect 20638 21758 20690 21810
rect 26574 21758 26626 21810
rect 8990 21646 9042 21698
rect 12126 21646 12178 21698
rect 16158 21646 16210 21698
rect 23886 21646 23938 21698
rect 27918 21646 27970 21698
rect 31278 21646 31330 21698
rect 4286 21534 4338 21586
rect 4622 21534 4674 21586
rect 13246 21534 13298 21586
rect 13918 21534 13970 21586
rect 18958 21534 19010 21586
rect 19294 21534 19346 21586
rect 19518 21534 19570 21586
rect 19742 21534 19794 21586
rect 19966 21534 20018 21586
rect 20974 21534 21026 21586
rect 21534 21534 21586 21586
rect 25230 21534 25282 21586
rect 25454 21534 25506 21586
rect 25902 21534 25954 21586
rect 26126 21534 26178 21586
rect 26350 21534 26402 21586
rect 26798 21534 26850 21586
rect 30158 21534 30210 21586
rect 30830 21534 30882 21586
rect 1934 21422 1986 21474
rect 4734 21422 4786 21474
rect 5182 21422 5234 21474
rect 5630 21422 5682 21474
rect 6078 21422 6130 21474
rect 9774 21422 9826 21474
rect 17950 21422 18002 21474
rect 18510 21422 18562 21474
rect 19630 21422 19682 21474
rect 20526 21422 20578 21474
rect 25678 21422 25730 21474
rect 31054 21422 31106 21474
rect 31838 21422 31890 21474
rect 5070 21310 5122 21362
rect 8878 21310 8930 21362
rect 9998 21310 10050 21362
rect 12238 21310 12290 21362
rect 16942 21310 16994 21362
rect 17726 21310 17778 21362
rect 24670 21310 24722 21362
rect 27134 21310 27186 21362
rect 31390 21310 31442 21362
rect 5372 21142 5424 21194
rect 5476 21142 5528 21194
rect 5580 21142 5632 21194
rect 13688 21142 13740 21194
rect 13792 21142 13844 21194
rect 13896 21142 13948 21194
rect 22004 21142 22056 21194
rect 22108 21142 22160 21194
rect 22212 21142 22264 21194
rect 30320 21142 30372 21194
rect 30424 21142 30476 21194
rect 30528 21142 30580 21194
rect 14366 20974 14418 21026
rect 19406 20974 19458 21026
rect 1934 20862 1986 20914
rect 4734 20862 4786 20914
rect 9550 20862 9602 20914
rect 19966 20862 20018 20914
rect 25118 20862 25170 20914
rect 27582 20862 27634 20914
rect 29598 20862 29650 20914
rect 30046 20862 30098 20914
rect 30158 20862 30210 20914
rect 3838 20750 3890 20802
rect 5854 20750 5906 20802
rect 6526 20750 6578 20802
rect 9774 20750 9826 20802
rect 9998 20750 10050 20802
rect 10446 20750 10498 20802
rect 14814 20750 14866 20802
rect 15262 20750 15314 20802
rect 19742 20750 19794 20802
rect 23102 20750 23154 20802
rect 28478 20750 28530 20802
rect 29150 20750 29202 20802
rect 29374 20750 29426 20802
rect 30382 20750 30434 20802
rect 33630 20750 33682 20802
rect 34078 20750 34130 20802
rect 14478 20638 14530 20690
rect 15150 20638 15202 20690
rect 20302 20638 20354 20690
rect 29710 20638 29762 20690
rect 8766 20526 8818 20578
rect 10110 20526 10162 20578
rect 10894 20526 10946 20578
rect 15038 20526 15090 20578
rect 15374 20526 15426 20578
rect 20414 20526 20466 20578
rect 30606 20526 30658 20578
rect 31390 20526 31442 20578
rect 9530 20358 9582 20410
rect 9634 20358 9686 20410
rect 9738 20358 9790 20410
rect 17846 20358 17898 20410
rect 17950 20358 18002 20410
rect 18054 20358 18106 20410
rect 26162 20358 26214 20410
rect 26266 20358 26318 20410
rect 26370 20358 26422 20410
rect 34478 20358 34530 20410
rect 34582 20358 34634 20410
rect 34686 20358 34738 20410
rect 14254 20190 14306 20242
rect 14926 20190 14978 20242
rect 23102 20190 23154 20242
rect 9662 20078 9714 20130
rect 9774 20078 9826 20130
rect 9886 20078 9938 20130
rect 13470 20078 13522 20130
rect 19406 20078 19458 20130
rect 19742 20078 19794 20130
rect 28926 20078 28978 20130
rect 29710 20078 29762 20130
rect 4286 19966 4338 20018
rect 10558 19966 10610 20018
rect 11230 19966 11282 20018
rect 14478 19966 14530 20018
rect 14702 19966 14754 20018
rect 15038 19966 15090 20018
rect 19070 19966 19122 20018
rect 19294 19966 19346 20018
rect 19518 19966 19570 20018
rect 20414 19966 20466 20018
rect 20750 19966 20802 20018
rect 25566 19966 25618 20018
rect 26574 19966 26626 20018
rect 31950 19966 32002 20018
rect 32622 19966 32674 20018
rect 2046 19854 2098 19906
rect 10334 19854 10386 19906
rect 14814 19854 14866 19906
rect 24222 19854 24274 19906
rect 25790 19854 25842 19906
rect 28478 19854 28530 19906
rect 33294 19854 33346 19906
rect 23886 19742 23938 19794
rect 25230 19742 25282 19794
rect 5372 19574 5424 19626
rect 5476 19574 5528 19626
rect 5580 19574 5632 19626
rect 13688 19574 13740 19626
rect 13792 19574 13844 19626
rect 13896 19574 13948 19626
rect 22004 19574 22056 19626
rect 22108 19574 22160 19626
rect 22212 19574 22264 19626
rect 30320 19574 30372 19626
rect 30424 19574 30476 19626
rect 30528 19574 30580 19626
rect 2718 19406 2770 19458
rect 12014 19406 12066 19458
rect 27582 19406 27634 19458
rect 10446 19294 10498 19346
rect 12126 19294 12178 19346
rect 23998 19294 24050 19346
rect 24446 19294 24498 19346
rect 5630 19182 5682 19234
rect 6190 19182 6242 19234
rect 9662 19182 9714 19234
rect 10110 19182 10162 19234
rect 14814 19182 14866 19234
rect 15486 19182 15538 19234
rect 19182 19182 19234 19234
rect 20078 19182 20130 19234
rect 24894 19182 24946 19234
rect 25342 19182 25394 19234
rect 28478 19182 28530 19234
rect 32062 19182 32114 19234
rect 32734 19182 32786 19234
rect 33182 19182 33234 19234
rect 2830 19070 2882 19122
rect 9214 19070 9266 19122
rect 9438 19070 9490 19122
rect 14254 19070 14306 19122
rect 14590 19070 14642 19122
rect 17726 19070 17778 19122
rect 18510 19070 18562 19122
rect 19406 19070 19458 19122
rect 25678 19070 25730 19122
rect 33854 19070 33906 19122
rect 34190 19070 34242 19122
rect 8654 18958 8706 19010
rect 9886 18958 9938 19010
rect 10894 18958 10946 19010
rect 18846 18958 18898 19010
rect 18958 18958 19010 19010
rect 19070 18958 19122 19010
rect 19742 18958 19794 19010
rect 29038 18958 29090 19010
rect 29822 18958 29874 19010
rect 32958 18958 33010 19010
rect 9530 18790 9582 18842
rect 9634 18790 9686 18842
rect 9738 18790 9790 18842
rect 17846 18790 17898 18842
rect 17950 18790 18002 18842
rect 18054 18790 18106 18842
rect 26162 18790 26214 18842
rect 26266 18790 26318 18842
rect 26370 18790 26422 18842
rect 34478 18790 34530 18842
rect 34582 18790 34634 18842
rect 34686 18790 34738 18842
rect 5966 18622 6018 18674
rect 9662 18622 9714 18674
rect 13134 18622 13186 18674
rect 14814 18622 14866 18674
rect 15150 18622 15202 18674
rect 16046 18622 16098 18674
rect 19966 18622 20018 18674
rect 33742 18622 33794 18674
rect 8990 18510 9042 18562
rect 2158 18398 2210 18450
rect 5742 18398 5794 18450
rect 6414 18398 6466 18450
rect 8766 18398 8818 18450
rect 10222 18398 10274 18450
rect 10670 18398 10722 18450
rect 13694 18398 13746 18450
rect 16158 18398 16210 18450
rect 17950 18398 18002 18450
rect 18398 18398 18450 18450
rect 20302 18398 20354 18450
rect 24446 18398 24498 18450
rect 25566 18398 25618 18450
rect 26238 18398 26290 18450
rect 26462 18398 26514 18450
rect 26798 18398 26850 18450
rect 27134 18398 27186 18450
rect 29934 18398 29986 18450
rect 33406 18398 33458 18450
rect 33966 18398 34018 18450
rect 8430 18286 8482 18338
rect 23998 18286 24050 18338
rect 25230 18286 25282 18338
rect 25790 18286 25842 18338
rect 26574 18286 26626 18338
rect 29374 18286 29426 18338
rect 31838 18286 31890 18338
rect 2718 18174 2770 18226
rect 6302 18174 6354 18226
rect 33070 18174 33122 18226
rect 33406 18174 33458 18226
rect 5372 18006 5424 18058
rect 5476 18006 5528 18058
rect 5580 18006 5632 18058
rect 13688 18006 13740 18058
rect 13792 18006 13844 18058
rect 13896 18006 13948 18058
rect 22004 18006 22056 18058
rect 22108 18006 22160 18058
rect 22212 18006 22264 18058
rect 30320 18006 30372 18058
rect 30424 18006 30476 18058
rect 30528 18006 30580 18058
rect 9214 17838 9266 17890
rect 10894 17838 10946 17890
rect 29934 17838 29986 17890
rect 8990 17726 9042 17778
rect 27582 17726 27634 17778
rect 11006 17614 11058 17666
rect 11454 17614 11506 17666
rect 11678 17614 11730 17666
rect 11790 17614 11842 17666
rect 12014 17614 12066 17666
rect 19294 17614 19346 17666
rect 19518 17614 19570 17666
rect 20190 17614 20242 17666
rect 26126 17614 26178 17666
rect 26574 17614 26626 17666
rect 30270 17614 30322 17666
rect 33630 17614 33682 17666
rect 34078 17614 34130 17666
rect 8990 17502 9042 17554
rect 9662 17502 9714 17554
rect 29486 17502 29538 17554
rect 12350 17390 12402 17442
rect 19406 17390 19458 17442
rect 19630 17390 19682 17442
rect 19742 17390 19794 17442
rect 20302 17390 20354 17442
rect 25902 17390 25954 17442
rect 26910 17390 26962 17442
rect 28030 17390 28082 17442
rect 28590 17390 28642 17442
rect 29150 17390 29202 17442
rect 30046 17390 30098 17442
rect 30606 17390 30658 17442
rect 31390 17390 31442 17442
rect 9530 17222 9582 17274
rect 9634 17222 9686 17274
rect 9738 17222 9790 17274
rect 17846 17222 17898 17274
rect 17950 17222 18002 17274
rect 18054 17222 18106 17274
rect 26162 17222 26214 17274
rect 26266 17222 26318 17274
rect 26370 17222 26422 17274
rect 34478 17222 34530 17274
rect 34582 17222 34634 17274
rect 34686 17222 34738 17274
rect 15262 17054 15314 17106
rect 23102 17054 23154 17106
rect 23662 17054 23714 17106
rect 25454 17054 25506 17106
rect 27582 17054 27634 17106
rect 28142 17054 28194 17106
rect 29150 17054 29202 17106
rect 34190 17054 34242 17106
rect 15598 16942 15650 16994
rect 19182 16942 19234 16994
rect 28702 16942 28754 16994
rect 29598 16942 29650 16994
rect 2718 16830 2770 16882
rect 4958 16830 5010 16882
rect 5518 16830 5570 16882
rect 6862 16830 6914 16882
rect 6974 16830 7026 16882
rect 7198 16830 7250 16882
rect 7422 16830 7474 16882
rect 16046 16830 16098 16882
rect 18622 16830 18674 16882
rect 18734 16830 18786 16882
rect 18958 16830 19010 16882
rect 20078 16830 20130 16882
rect 20526 16830 20578 16882
rect 25230 16830 25282 16882
rect 29038 16830 29090 16882
rect 29262 16830 29314 16882
rect 29934 16830 29986 16882
rect 31614 16830 31666 16882
rect 33630 16830 33682 16882
rect 18846 16718 18898 16770
rect 27358 16718 27410 16770
rect 27694 16718 27746 16770
rect 28478 16718 28530 16770
rect 1710 16606 1762 16658
rect 15934 16606 15986 16658
rect 25566 16606 25618 16658
rect 5372 16438 5424 16490
rect 5476 16438 5528 16490
rect 5580 16438 5632 16490
rect 13688 16438 13740 16490
rect 13792 16438 13844 16490
rect 13896 16438 13948 16490
rect 22004 16438 22056 16490
rect 22108 16438 22160 16490
rect 22212 16438 22264 16490
rect 30320 16438 30372 16490
rect 30424 16438 30476 16490
rect 30528 16438 30580 16490
rect 1934 16158 1986 16210
rect 7422 16158 7474 16210
rect 22542 16158 22594 16210
rect 29262 16158 29314 16210
rect 4286 16046 4338 16098
rect 4734 16046 4786 16098
rect 10446 16046 10498 16098
rect 10782 16046 10834 16098
rect 11006 16046 11058 16098
rect 14814 16046 14866 16098
rect 15486 16046 15538 16098
rect 21422 16046 21474 16098
rect 22206 16046 22258 16098
rect 22990 16046 23042 16098
rect 23550 16046 23602 16098
rect 26910 16046 26962 16098
rect 29374 16046 29426 16098
rect 33630 16046 33682 16098
rect 34078 16046 34130 16098
rect 6190 15934 6242 15986
rect 7534 15934 7586 15986
rect 21982 15934 22034 15986
rect 29150 15934 29202 15986
rect 29710 15934 29762 15986
rect 30606 15934 30658 15986
rect 6302 15822 6354 15874
rect 6414 15822 6466 15874
rect 7310 15822 7362 15874
rect 10782 15822 10834 15874
rect 17726 15822 17778 15874
rect 18510 15822 18562 15874
rect 20414 15822 20466 15874
rect 21646 15822 21698 15874
rect 22430 15822 22482 15874
rect 22542 15822 22594 15874
rect 26126 15822 26178 15874
rect 26686 15822 26738 15874
rect 27470 15822 27522 15874
rect 27806 15822 27858 15874
rect 28142 15822 28194 15874
rect 31390 15822 31442 15874
rect 9530 15654 9582 15706
rect 9634 15654 9686 15706
rect 9738 15654 9790 15706
rect 17846 15654 17898 15706
rect 17950 15654 18002 15706
rect 18054 15654 18106 15706
rect 26162 15654 26214 15706
rect 26266 15654 26318 15706
rect 26370 15654 26422 15706
rect 34478 15654 34530 15706
rect 34582 15654 34634 15706
rect 34686 15654 34738 15706
rect 7198 15486 7250 15538
rect 19854 15486 19906 15538
rect 20638 15486 20690 15538
rect 22990 15486 23042 15538
rect 23326 15486 23378 15538
rect 27470 15486 27522 15538
rect 28702 15486 28754 15538
rect 3390 15374 3442 15426
rect 6862 15374 6914 15426
rect 7646 15374 7698 15426
rect 15598 15374 15650 15426
rect 15934 15374 15986 15426
rect 16270 15374 16322 15426
rect 22878 15374 22930 15426
rect 29038 15374 29090 15426
rect 3838 15262 3890 15314
rect 4958 15262 5010 15314
rect 6414 15262 6466 15314
rect 7310 15262 7362 15314
rect 7422 15262 7474 15314
rect 11454 15262 11506 15314
rect 13582 15262 13634 15314
rect 14030 15262 14082 15314
rect 16494 15262 16546 15314
rect 19406 15262 19458 15314
rect 20078 15262 20130 15314
rect 20526 15262 20578 15314
rect 20862 15262 20914 15314
rect 23662 15262 23714 15314
rect 29262 15262 29314 15314
rect 29934 15262 29986 15314
rect 3614 15150 3666 15202
rect 4622 15150 4674 15202
rect 18958 15150 19010 15202
rect 24110 15150 24162 15202
rect 31054 15150 31106 15202
rect 4174 15038 4226 15090
rect 10446 15038 10498 15090
rect 29598 15038 29650 15090
rect 5372 14870 5424 14922
rect 5476 14870 5528 14922
rect 5580 14870 5632 14922
rect 13688 14870 13740 14922
rect 13792 14870 13844 14922
rect 13896 14870 13948 14922
rect 22004 14870 22056 14922
rect 22108 14870 22160 14922
rect 22212 14870 22264 14922
rect 30320 14870 30372 14922
rect 30424 14870 30476 14922
rect 30528 14870 30580 14922
rect 4398 14702 4450 14754
rect 11006 14702 11058 14754
rect 33518 14702 33570 14754
rect 8094 14590 8146 14642
rect 10222 14590 10274 14642
rect 20526 14590 20578 14642
rect 22878 14590 22930 14642
rect 1822 14478 1874 14530
rect 2606 14478 2658 14530
rect 3278 14478 3330 14530
rect 3838 14478 3890 14530
rect 5518 14478 5570 14530
rect 5854 14478 5906 14530
rect 6078 14478 6130 14530
rect 6526 14478 6578 14530
rect 6862 14478 6914 14530
rect 15822 14478 15874 14530
rect 16382 14478 16434 14530
rect 22430 14478 22482 14530
rect 22542 14478 22594 14530
rect 22990 14478 23042 14530
rect 23550 14478 23602 14530
rect 23998 14478 24050 14530
rect 24446 14478 24498 14530
rect 29038 14478 29090 14530
rect 30046 14478 30098 14530
rect 30606 14478 30658 14530
rect 31726 14478 31778 14530
rect 2046 14366 2098 14418
rect 2942 14366 2994 14418
rect 4174 14366 4226 14418
rect 6638 14366 6690 14418
rect 8542 14366 8594 14418
rect 9998 14366 10050 14418
rect 11118 14366 11170 14418
rect 11342 14366 11394 14418
rect 18734 14366 18786 14418
rect 20638 14366 20690 14418
rect 23662 14366 23714 14418
rect 26798 14366 26850 14418
rect 29486 14366 29538 14418
rect 29710 14366 29762 14418
rect 4734 14254 4786 14306
rect 5742 14254 5794 14306
rect 7646 14254 7698 14306
rect 19518 14254 19570 14306
rect 20414 14254 20466 14306
rect 21422 14254 21474 14306
rect 22766 14254 22818 14306
rect 27582 14254 27634 14306
rect 29262 14254 29314 14306
rect 9530 14086 9582 14138
rect 9634 14086 9686 14138
rect 9738 14086 9790 14138
rect 17846 14086 17898 14138
rect 17950 14086 18002 14138
rect 18054 14086 18106 14138
rect 26162 14086 26214 14138
rect 26266 14086 26318 14138
rect 26370 14086 26422 14138
rect 34478 14086 34530 14138
rect 34582 14086 34634 14138
rect 34686 14086 34738 14138
rect 1822 13918 1874 13970
rect 2942 13918 2994 13970
rect 6526 13918 6578 13970
rect 7534 13918 7586 13970
rect 8094 13918 8146 13970
rect 16158 13918 16210 13970
rect 21758 13918 21810 13970
rect 27470 13918 27522 13970
rect 29486 13918 29538 13970
rect 3390 13806 3442 13858
rect 4398 13806 4450 13858
rect 5742 13806 5794 13858
rect 19854 13806 19906 13858
rect 22206 13806 22258 13858
rect 28590 13806 28642 13858
rect 29262 13806 29314 13858
rect 4622 13694 4674 13746
rect 8318 13694 8370 13746
rect 10894 13694 10946 13746
rect 11454 13694 11506 13746
rect 11902 13694 11954 13746
rect 13358 13694 13410 13746
rect 13918 13694 13970 13746
rect 19518 13694 19570 13746
rect 20638 13694 20690 13746
rect 21086 13694 21138 13746
rect 21758 13694 21810 13746
rect 23438 13694 23490 13746
rect 27806 13694 27858 13746
rect 28478 13694 28530 13746
rect 29038 13694 29090 13746
rect 30158 13694 30210 13746
rect 33070 13694 33122 13746
rect 2494 13582 2546 13634
rect 5966 13582 6018 13634
rect 6414 13582 6466 13634
rect 7086 13582 7138 13634
rect 12350 13582 12402 13634
rect 20526 13582 20578 13634
rect 28030 13582 28082 13634
rect 28814 13582 28866 13634
rect 31838 13582 31890 13634
rect 33518 13582 33570 13634
rect 11790 13470 11842 13522
rect 16942 13470 16994 13522
rect 29598 13470 29650 13522
rect 5372 13302 5424 13354
rect 5476 13302 5528 13354
rect 5580 13302 5632 13354
rect 13688 13302 13740 13354
rect 13792 13302 13844 13354
rect 13896 13302 13948 13354
rect 22004 13302 22056 13354
rect 22108 13302 22160 13354
rect 22212 13302 22264 13354
rect 30320 13302 30372 13354
rect 30424 13302 30476 13354
rect 30528 13302 30580 13354
rect 11454 13134 11506 13186
rect 11678 13134 11730 13186
rect 29150 13134 29202 13186
rect 30046 13134 30098 13186
rect 30382 13134 30434 13186
rect 3054 13022 3106 13074
rect 14590 13022 14642 13074
rect 16270 13022 16322 13074
rect 20750 13022 20802 13074
rect 22430 13022 22482 13074
rect 29486 13022 29538 13074
rect 29822 13022 29874 13074
rect 3166 12910 3218 12962
rect 5630 12910 5682 12962
rect 6078 12910 6130 12962
rect 7982 12910 8034 12962
rect 8430 12910 8482 12962
rect 12014 12910 12066 12962
rect 12350 12910 12402 12962
rect 14926 12910 14978 12962
rect 15822 12910 15874 12962
rect 18622 12910 18674 12962
rect 21534 12910 21586 12962
rect 22094 12910 22146 12962
rect 23886 12910 23938 12962
rect 30606 12910 30658 12962
rect 33630 12910 33682 12962
rect 34078 12910 34130 12962
rect 13470 12798 13522 12850
rect 13806 12798 13858 12850
rect 14478 12798 14530 12850
rect 14814 12798 14866 12850
rect 16046 12798 16098 12850
rect 16382 12798 16434 12850
rect 19630 12798 19682 12850
rect 21310 12798 21362 12850
rect 22654 12798 22706 12850
rect 24670 12798 24722 12850
rect 25790 12798 25842 12850
rect 29374 12798 29426 12850
rect 31390 12798 31442 12850
rect 3278 12686 3330 12738
rect 6190 12686 6242 12738
rect 6302 12686 6354 12738
rect 6862 12686 6914 12738
rect 10894 12686 10946 12738
rect 12126 12686 12178 12738
rect 12238 12686 12290 12738
rect 12910 12686 12962 12738
rect 18734 12686 18786 12738
rect 19070 12686 19122 12738
rect 20190 12686 20242 12738
rect 23102 12686 23154 12738
rect 23998 12686 24050 12738
rect 24558 12686 24610 12738
rect 25230 12686 25282 12738
rect 9530 12518 9582 12570
rect 9634 12518 9686 12570
rect 9738 12518 9790 12570
rect 17846 12518 17898 12570
rect 17950 12518 18002 12570
rect 18054 12518 18106 12570
rect 26162 12518 26214 12570
rect 26266 12518 26318 12570
rect 26370 12518 26422 12570
rect 34478 12518 34530 12570
rect 34582 12518 34634 12570
rect 34686 12518 34738 12570
rect 5406 12350 5458 12402
rect 5630 12350 5682 12402
rect 5854 12350 5906 12402
rect 7310 12350 7362 12402
rect 7870 12350 7922 12402
rect 12014 12350 12066 12402
rect 14590 12350 14642 12402
rect 16158 12350 16210 12402
rect 23998 12350 24050 12402
rect 29262 12350 29314 12402
rect 5966 12238 6018 12290
rect 6526 12238 6578 12290
rect 7086 12238 7138 12290
rect 9550 12238 9602 12290
rect 11454 12238 11506 12290
rect 12462 12238 12514 12290
rect 16046 12238 16098 12290
rect 19854 12238 19906 12290
rect 23662 12238 23714 12290
rect 25790 12238 25842 12290
rect 1822 12126 1874 12178
rect 2270 12126 2322 12178
rect 4510 12126 4562 12178
rect 6302 12126 6354 12178
rect 6974 12126 7026 12178
rect 7422 12126 7474 12178
rect 9886 12126 9938 12178
rect 11342 12126 11394 12178
rect 11566 12126 11618 12178
rect 12350 12126 12402 12178
rect 14478 12126 14530 12178
rect 14702 12126 14754 12178
rect 18958 12126 19010 12178
rect 19406 12126 19458 12178
rect 21086 12126 21138 12178
rect 22318 12126 22370 12178
rect 22878 12126 22930 12178
rect 23438 12126 23490 12178
rect 24558 12126 24610 12178
rect 26126 12126 26178 12178
rect 26910 12126 26962 12178
rect 27134 12126 27186 12178
rect 29598 12126 29650 12178
rect 30270 12126 30322 12178
rect 33630 12126 33682 12178
rect 34190 12126 34242 12178
rect 6414 12014 6466 12066
rect 8318 12014 8370 12066
rect 21646 12014 21698 12066
rect 31838 12014 31890 12066
rect 14926 11902 14978 11954
rect 16270 11902 16322 11954
rect 18622 11902 18674 11954
rect 18958 11902 19010 11954
rect 22542 11902 22594 11954
rect 25678 11902 25730 11954
rect 5372 11734 5424 11786
rect 5476 11734 5528 11786
rect 5580 11734 5632 11786
rect 13688 11734 13740 11786
rect 13792 11734 13844 11786
rect 13896 11734 13948 11786
rect 22004 11734 22056 11786
rect 22108 11734 22160 11786
rect 22212 11734 22264 11786
rect 30320 11734 30372 11786
rect 30424 11734 30476 11786
rect 30528 11734 30580 11786
rect 1934 11566 1986 11618
rect 9998 11566 10050 11618
rect 20078 11454 20130 11506
rect 22878 11454 22930 11506
rect 25006 11454 25058 11506
rect 26126 11454 26178 11506
rect 29822 11454 29874 11506
rect 3838 11342 3890 11394
rect 6526 11342 6578 11394
rect 6862 11342 6914 11394
rect 15150 11342 15202 11394
rect 15710 11342 15762 11394
rect 17278 11342 17330 11394
rect 19182 11342 19234 11394
rect 19742 11342 19794 11394
rect 20526 11342 20578 11394
rect 22094 11342 22146 11394
rect 22430 11342 22482 11394
rect 23550 11342 23602 11394
rect 24558 11342 24610 11394
rect 26686 11342 26738 11394
rect 27022 11342 27074 11394
rect 27582 11342 27634 11394
rect 30718 11342 30770 11394
rect 31166 11342 31218 11394
rect 9214 11230 9266 11282
rect 14590 11230 14642 11282
rect 14814 11230 14866 11282
rect 18622 11230 18674 11282
rect 20414 11230 20466 11282
rect 22990 11230 23042 11282
rect 23886 11230 23938 11282
rect 27918 11230 27970 11282
rect 14702 11118 14754 11170
rect 17614 11118 17666 11170
rect 21422 11118 21474 11170
rect 23438 11118 23490 11170
rect 28254 11118 28306 11170
rect 33518 11118 33570 11170
rect 34302 11118 34354 11170
rect 9530 10950 9582 11002
rect 9634 10950 9686 11002
rect 9738 10950 9790 11002
rect 17846 10950 17898 11002
rect 17950 10950 18002 11002
rect 18054 10950 18106 11002
rect 26162 10950 26214 11002
rect 26266 10950 26318 11002
rect 26370 10950 26422 11002
rect 34478 10950 34530 11002
rect 34582 10950 34634 11002
rect 34686 10950 34738 11002
rect 11678 10782 11730 10834
rect 14814 10782 14866 10834
rect 15486 10782 15538 10834
rect 27358 10782 27410 10834
rect 28030 10782 28082 10834
rect 31390 10782 31442 10834
rect 12574 10670 12626 10722
rect 16382 10670 16434 10722
rect 21422 10670 21474 10722
rect 22878 10670 22930 10722
rect 24558 10670 24610 10722
rect 25566 10670 25618 10722
rect 3838 10558 3890 10610
rect 12014 10558 12066 10610
rect 12798 10558 12850 10610
rect 15822 10558 15874 10610
rect 16606 10558 16658 10610
rect 18062 10558 18114 10610
rect 18846 10558 18898 10610
rect 19070 10558 19122 10610
rect 21870 10558 21922 10610
rect 22318 10558 22370 10610
rect 30382 10558 30434 10610
rect 30830 10558 30882 10610
rect 14254 10446 14306 10498
rect 18398 10446 18450 10498
rect 20638 10446 20690 10498
rect 24670 10446 24722 10498
rect 26014 10446 26066 10498
rect 1934 10334 1986 10386
rect 18958 10334 19010 10386
rect 24334 10334 24386 10386
rect 5372 10166 5424 10218
rect 5476 10166 5528 10218
rect 5580 10166 5632 10218
rect 13688 10166 13740 10218
rect 13792 10166 13844 10218
rect 13896 10166 13948 10218
rect 22004 10166 22056 10218
rect 22108 10166 22160 10218
rect 22212 10166 22264 10218
rect 30320 10166 30372 10218
rect 30424 10166 30476 10218
rect 30528 10166 30580 10218
rect 2158 9998 2210 10050
rect 3390 9998 3442 10050
rect 14702 9998 14754 10050
rect 17390 9998 17442 10050
rect 17726 9998 17778 10050
rect 25566 9998 25618 10050
rect 33518 9998 33570 10050
rect 3278 9886 3330 9938
rect 3838 9886 3890 9938
rect 12238 9886 12290 9938
rect 14142 9886 14194 9938
rect 16494 9886 16546 9938
rect 21758 9886 21810 9938
rect 2718 9774 2770 9826
rect 6862 9774 6914 9826
rect 7982 9774 8034 9826
rect 8542 9774 8594 9826
rect 9214 9774 9266 9826
rect 12574 9774 12626 9826
rect 14814 9774 14866 9826
rect 14926 9774 14978 9826
rect 16606 9774 16658 9826
rect 18286 9774 18338 9826
rect 20750 9774 20802 9826
rect 22542 9774 22594 9826
rect 22990 9774 23042 9826
rect 25230 9774 25282 9826
rect 26350 9774 26402 9826
rect 26686 9774 26738 9826
rect 31838 9774 31890 9826
rect 2270 9662 2322 9714
rect 2942 9662 2994 9714
rect 7086 9662 7138 9714
rect 14254 9662 14306 9714
rect 16270 9662 16322 9714
rect 17950 9662 18002 9714
rect 18622 9662 18674 9714
rect 20302 9662 20354 9714
rect 22766 9662 22818 9714
rect 23102 9662 23154 9714
rect 23886 9662 23938 9714
rect 25118 9662 25170 9714
rect 6526 9550 6578 9602
rect 7534 9550 7586 9602
rect 8318 9550 8370 9602
rect 11454 9550 11506 9602
rect 12798 9550 12850 9602
rect 14030 9550 14082 9602
rect 20526 9550 20578 9602
rect 20638 9550 20690 9602
rect 9530 9382 9582 9434
rect 9634 9382 9686 9434
rect 9738 9382 9790 9434
rect 17846 9382 17898 9434
rect 17950 9382 18002 9434
rect 18054 9382 18106 9434
rect 26162 9382 26214 9434
rect 26266 9382 26318 9434
rect 26370 9382 26422 9434
rect 34478 9382 34530 9434
rect 34582 9382 34634 9434
rect 34686 9382 34738 9434
rect 5966 9214 6018 9266
rect 6862 9214 6914 9266
rect 28702 9214 28754 9266
rect 32062 9214 32114 9266
rect 32622 9214 32674 9266
rect 33182 9214 33234 9266
rect 6526 9102 6578 9154
rect 16718 9102 16770 9154
rect 17502 9102 17554 9154
rect 18734 9102 18786 9154
rect 22878 9102 22930 9154
rect 27246 9102 27298 9154
rect 33854 9102 33906 9154
rect 2270 8990 2322 9042
rect 3054 8990 3106 9042
rect 3502 8990 3554 9042
rect 6750 8990 6802 9042
rect 7086 8990 7138 9042
rect 7198 8990 7250 9042
rect 15262 8990 15314 9042
rect 15822 8990 15874 9042
rect 16494 8990 16546 9042
rect 19182 8990 19234 9042
rect 20526 8990 20578 9042
rect 21086 8990 21138 9042
rect 24558 8990 24610 9042
rect 25902 8990 25954 9042
rect 26126 8990 26178 9042
rect 28478 8990 28530 9042
rect 28926 8990 28978 9042
rect 29486 8990 29538 9042
rect 33406 8990 33458 9042
rect 34078 8990 34130 9042
rect 1822 8878 1874 8930
rect 7758 8878 7810 8930
rect 16606 8878 16658 8930
rect 17390 8878 17442 8930
rect 19294 8878 19346 8930
rect 20302 8878 20354 8930
rect 22542 8878 22594 8930
rect 24334 8878 24386 8930
rect 25790 8878 25842 8930
rect 20190 8766 20242 8818
rect 21310 8766 21362 8818
rect 22654 8766 22706 8818
rect 24222 8766 24274 8818
rect 24670 8766 24722 8818
rect 26462 8766 26514 8818
rect 5372 8598 5424 8650
rect 5476 8598 5528 8650
rect 5580 8598 5632 8650
rect 13688 8598 13740 8650
rect 13792 8598 13844 8650
rect 13896 8598 13948 8650
rect 22004 8598 22056 8650
rect 22108 8598 22160 8650
rect 22212 8598 22264 8650
rect 30320 8598 30372 8650
rect 30424 8598 30476 8650
rect 30528 8598 30580 8650
rect 33966 8430 34018 8482
rect 1934 8318 1986 8370
rect 6078 8318 6130 8370
rect 6414 8318 6466 8370
rect 14030 8318 14082 8370
rect 25790 8318 25842 8370
rect 27022 8318 27074 8370
rect 29262 8318 29314 8370
rect 29598 8318 29650 8370
rect 3838 8206 3890 8258
rect 13470 8206 13522 8258
rect 13806 8206 13858 8258
rect 14478 8206 14530 8258
rect 14814 8206 14866 8258
rect 16718 8206 16770 8258
rect 17054 8206 17106 8258
rect 18286 8206 18338 8258
rect 20302 8206 20354 8258
rect 22094 8206 22146 8258
rect 22654 8206 22706 8258
rect 25902 8206 25954 8258
rect 26238 8206 26290 8258
rect 26462 8206 26514 8258
rect 31614 8206 31666 8258
rect 4622 8094 4674 8146
rect 12462 8094 12514 8146
rect 12798 8094 12850 8146
rect 14702 8094 14754 8146
rect 15598 8094 15650 8146
rect 29822 8094 29874 8146
rect 30158 8094 30210 8146
rect 31278 8094 31330 8146
rect 4958 7982 5010 8034
rect 6190 7982 6242 8034
rect 10894 7982 10946 8034
rect 11230 7982 11282 8034
rect 12910 7982 12962 8034
rect 13918 7982 13970 8034
rect 14142 7982 14194 8034
rect 15262 7982 15314 8034
rect 19294 7982 19346 8034
rect 19518 7982 19570 8034
rect 19630 7982 19682 8034
rect 19742 7982 19794 8034
rect 20638 7982 20690 8034
rect 25230 7982 25282 8034
rect 26238 7982 26290 8034
rect 30942 7982 30994 8034
rect 9530 7814 9582 7866
rect 9634 7814 9686 7866
rect 9738 7814 9790 7866
rect 17846 7814 17898 7866
rect 17950 7814 18002 7866
rect 18054 7814 18106 7866
rect 26162 7814 26214 7866
rect 26266 7814 26318 7866
rect 26370 7814 26422 7866
rect 34478 7814 34530 7866
rect 34582 7814 34634 7866
rect 34686 7814 34738 7866
rect 4846 7646 4898 7698
rect 6078 7646 6130 7698
rect 6638 7646 6690 7698
rect 12126 7646 12178 7698
rect 13022 7646 13074 7698
rect 17726 7646 17778 7698
rect 21310 7646 21362 7698
rect 22542 7646 22594 7698
rect 25790 7646 25842 7698
rect 26798 7646 26850 7698
rect 29598 7646 29650 7698
rect 33630 7646 33682 7698
rect 5966 7534 6018 7586
rect 7198 7534 7250 7586
rect 12014 7534 12066 7586
rect 15150 7534 15202 7586
rect 17390 7534 17442 7586
rect 21198 7534 21250 7586
rect 23326 7534 23378 7586
rect 26574 7534 26626 7586
rect 27022 7534 27074 7586
rect 27358 7534 27410 7586
rect 27694 7534 27746 7586
rect 28702 7534 28754 7586
rect 2046 7422 2098 7474
rect 2494 7422 2546 7474
rect 5518 7422 5570 7474
rect 5854 7422 5906 7474
rect 6414 7422 6466 7474
rect 6974 7422 7026 7474
rect 12910 7422 12962 7474
rect 13246 7422 13298 7474
rect 15486 7422 15538 7474
rect 19406 7422 19458 7474
rect 21534 7422 21586 7474
rect 22206 7422 22258 7474
rect 22654 7422 22706 7474
rect 22878 7422 22930 7474
rect 23214 7422 23266 7474
rect 28478 7422 28530 7474
rect 29262 7422 29314 7474
rect 29934 7422 29986 7474
rect 13134 7310 13186 7362
rect 18958 7310 19010 7362
rect 26126 7310 26178 7362
rect 29038 7310 29090 7362
rect 31838 7310 31890 7362
rect 33406 7310 33458 7362
rect 34190 7310 34242 7362
rect 12574 7198 12626 7250
rect 27134 7198 27186 7250
rect 5372 7030 5424 7082
rect 5476 7030 5528 7082
rect 5580 7030 5632 7082
rect 13688 7030 13740 7082
rect 13792 7030 13844 7082
rect 13896 7030 13948 7082
rect 22004 7030 22056 7082
rect 22108 7030 22160 7082
rect 22212 7030 22264 7082
rect 30320 7030 30372 7082
rect 30424 7030 30476 7082
rect 30528 7030 30580 7082
rect 4846 6862 4898 6914
rect 4062 6638 4114 6690
rect 4734 6638 4786 6690
rect 5630 6862 5682 6914
rect 5966 6862 6018 6914
rect 16382 6862 16434 6914
rect 19518 6862 19570 6914
rect 6302 6750 6354 6802
rect 28254 6750 28306 6802
rect 29598 6750 29650 6802
rect 29822 6750 29874 6802
rect 5182 6638 5234 6690
rect 7758 6638 7810 6690
rect 8430 6638 8482 6690
rect 11454 6638 11506 6690
rect 20078 6638 20130 6690
rect 22542 6638 22594 6690
rect 22878 6638 22930 6690
rect 26462 6638 26514 6690
rect 26798 6638 26850 6690
rect 26910 6638 26962 6690
rect 27246 6638 27298 6690
rect 27918 6638 27970 6690
rect 29374 6638 29426 6690
rect 30158 6638 30210 6690
rect 30606 6638 30658 6690
rect 31166 6638 31218 6690
rect 2494 6526 2546 6578
rect 6638 6526 6690 6578
rect 16606 6526 16658 6578
rect 16942 6526 16994 6578
rect 20190 6526 20242 6578
rect 23214 6526 23266 6578
rect 26574 6526 26626 6578
rect 28590 6526 28642 6578
rect 30046 6526 30098 6578
rect 30270 6526 30322 6578
rect 33518 6526 33570 6578
rect 5742 6414 5794 6466
rect 6414 6414 6466 6466
rect 10670 6414 10722 6466
rect 16046 6414 16098 6466
rect 19182 6414 19234 6466
rect 22766 6414 22818 6466
rect 27694 6414 27746 6466
rect 27806 6414 27858 6466
rect 28366 6414 28418 6466
rect 34302 6414 34354 6466
rect 9530 6246 9582 6298
rect 9634 6246 9686 6298
rect 9738 6246 9790 6298
rect 17846 6246 17898 6298
rect 17950 6246 18002 6298
rect 18054 6246 18106 6298
rect 26162 6246 26214 6298
rect 26266 6246 26318 6298
rect 26370 6246 26422 6298
rect 34478 6246 34530 6298
rect 34582 6246 34634 6298
rect 34686 6246 34738 6298
rect 5182 6078 5234 6130
rect 6638 6078 6690 6130
rect 8318 6078 8370 6130
rect 9662 6078 9714 6130
rect 12798 6078 12850 6130
rect 13694 6078 13746 6130
rect 16494 6078 16546 6130
rect 17726 6078 17778 6130
rect 19518 6078 19570 6130
rect 20078 6078 20130 6130
rect 25902 6078 25954 6130
rect 31054 6078 31106 6130
rect 31838 6078 31890 6130
rect 32174 6078 32226 6130
rect 33182 6078 33234 6130
rect 34190 6078 34242 6130
rect 12126 5966 12178 6018
rect 14814 5966 14866 6018
rect 15150 5966 15202 6018
rect 16158 5966 16210 6018
rect 18174 5966 18226 6018
rect 28702 5966 28754 6018
rect 31166 5966 31218 6018
rect 2270 5854 2322 5906
rect 2942 5854 2994 5906
rect 5966 5854 6018 5906
rect 6190 5854 6242 5906
rect 6526 5854 6578 5906
rect 6862 5854 6914 5906
rect 8542 5854 8594 5906
rect 11118 5854 11170 5906
rect 11566 5854 11618 5906
rect 12574 5854 12626 5906
rect 13022 5854 13074 5906
rect 13246 5854 13298 5906
rect 13918 5854 13970 5906
rect 14030 5854 14082 5906
rect 15486 5854 15538 5906
rect 15934 5854 15986 5906
rect 16718 5854 16770 5906
rect 18622 5854 18674 5906
rect 20414 5854 20466 5906
rect 29598 5854 29650 5906
rect 30046 5854 30098 5906
rect 31502 5854 31554 5906
rect 32398 5854 32450 5906
rect 33630 5854 33682 5906
rect 7198 5742 7250 5794
rect 12014 5742 12066 5794
rect 12686 5742 12738 5794
rect 13806 5742 13858 5794
rect 18958 5742 19010 5794
rect 19406 5742 19458 5794
rect 28814 5742 28866 5794
rect 9550 5630 9602 5682
rect 9886 5630 9938 5682
rect 14366 5630 14418 5682
rect 14702 5630 14754 5682
rect 19742 5630 19794 5682
rect 5372 5462 5424 5514
rect 5476 5462 5528 5514
rect 5580 5462 5632 5514
rect 13688 5462 13740 5514
rect 13792 5462 13844 5514
rect 13896 5462 13948 5514
rect 22004 5462 22056 5514
rect 22108 5462 22160 5514
rect 22212 5462 22264 5514
rect 30320 5462 30372 5514
rect 30424 5462 30476 5514
rect 30528 5462 30580 5514
rect 5742 5294 5794 5346
rect 6078 5294 6130 5346
rect 11678 5294 11730 5346
rect 13582 5294 13634 5346
rect 19742 5294 19794 5346
rect 25790 5294 25842 5346
rect 29262 5294 29314 5346
rect 4734 5182 4786 5234
rect 6302 5182 6354 5234
rect 6750 5182 6802 5234
rect 20302 5182 20354 5234
rect 29374 5182 29426 5234
rect 30046 5182 30098 5234
rect 33630 5182 33682 5234
rect 4286 5070 4338 5122
rect 7758 5070 7810 5122
rect 8206 5070 8258 5122
rect 8654 5070 8706 5122
rect 16046 5070 16098 5122
rect 16606 5070 16658 5122
rect 22318 5070 22370 5122
rect 22766 5070 22818 5122
rect 28478 5070 28530 5122
rect 29598 5070 29650 5122
rect 30718 5070 30770 5122
rect 34190 5070 34242 5122
rect 7422 4958 7474 5010
rect 13470 4958 13522 5010
rect 29934 4958 29986 5010
rect 3278 4846 3330 4898
rect 4622 4846 4674 4898
rect 11118 4846 11170 4898
rect 18958 4846 19010 4898
rect 25118 4846 25170 4898
rect 27582 4846 27634 4898
rect 31726 4846 31778 4898
rect 9530 4678 9582 4730
rect 9634 4678 9686 4730
rect 9738 4678 9790 4730
rect 17846 4678 17898 4730
rect 17950 4678 18002 4730
rect 18054 4678 18106 4730
rect 26162 4678 26214 4730
rect 26266 4678 26318 4730
rect 26370 4678 26422 4730
rect 34478 4678 34530 4730
rect 34582 4678 34634 4730
rect 34686 4678 34738 4730
rect 8542 4510 8594 4562
rect 10782 4510 10834 4562
rect 13134 4510 13186 4562
rect 13694 4510 13746 4562
rect 18622 4510 18674 4562
rect 19406 4510 19458 4562
rect 22654 4510 22706 4562
rect 23998 4510 24050 4562
rect 25678 4510 25730 4562
rect 29374 4510 29426 4562
rect 29934 4510 29986 4562
rect 30494 4510 30546 4562
rect 30942 4510 30994 4562
rect 32174 4510 32226 4562
rect 33854 4510 33906 4562
rect 10670 4398 10722 4450
rect 11006 4398 11058 4450
rect 12126 4398 12178 4450
rect 17502 4398 17554 4450
rect 18398 4398 18450 4450
rect 23438 4398 23490 4450
rect 25902 4398 25954 4450
rect 33182 4398 33234 4450
rect 3950 4286 4002 4338
rect 4622 4286 4674 4338
rect 5182 4286 5234 4338
rect 5630 4286 5682 4338
rect 5966 4286 6018 4338
rect 9102 4286 9154 4338
rect 10222 4286 10274 4338
rect 11118 4286 11170 4338
rect 11902 4286 11954 4338
rect 16158 4286 16210 4338
rect 16718 4286 16770 4338
rect 18174 4286 18226 4338
rect 21646 4286 21698 4338
rect 22318 4286 22370 4338
rect 26462 4286 26514 4338
rect 26910 4286 26962 4338
rect 30382 4286 30434 4338
rect 32622 4286 32674 4338
rect 34078 4286 34130 4338
rect 9886 4174 9938 4226
rect 11566 4174 11618 4226
rect 33070 4174 33122 4226
rect 1934 4062 1986 4114
rect 17390 4062 17442 4114
rect 23550 4062 23602 4114
rect 26014 4062 26066 4114
rect 5372 3894 5424 3946
rect 5476 3894 5528 3946
rect 5580 3894 5632 3946
rect 13688 3894 13740 3946
rect 13792 3894 13844 3946
rect 13896 3894 13948 3946
rect 22004 3894 22056 3946
rect 22108 3894 22160 3946
rect 22212 3894 22264 3946
rect 30320 3894 30372 3946
rect 30424 3894 30476 3946
rect 30528 3894 30580 3946
rect 2270 3614 2322 3666
rect 8878 3614 8930 3666
rect 10334 3614 10386 3666
rect 12686 3614 12738 3666
rect 14142 3614 14194 3666
rect 19966 3614 20018 3666
rect 21870 3614 21922 3666
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 32958 3614 33010 3666
rect 4622 3502 4674 3554
rect 5966 3502 6018 3554
rect 9326 3502 9378 3554
rect 13134 3502 13186 3554
rect 17390 3502 17442 3554
rect 20078 3502 20130 3554
rect 20750 3502 20802 3554
rect 24558 3502 24610 3554
rect 28590 3502 28642 3554
rect 31726 3502 31778 3554
rect 33294 3502 33346 3554
rect 18510 3390 18562 3442
rect 32510 3390 32562 3442
rect 33518 3390 33570 3442
rect 33854 3390 33906 3442
rect 34190 3390 34242 3442
rect 6638 3278 6690 3330
rect 9530 3110 9582 3162
rect 9634 3110 9686 3162
rect 9738 3110 9790 3162
rect 17846 3110 17898 3162
rect 17950 3110 18002 3162
rect 18054 3110 18106 3162
rect 26162 3110 26214 3162
rect 26266 3110 26318 3162
rect 26370 3110 26422 3162
rect 34478 3110 34530 3162
rect 34582 3110 34634 3162
rect 34686 3110 34738 3162
<< metal2 >>
rect 1792 25200 1904 26000
rect 5376 25200 5488 26000
rect 8960 25200 9072 26000
rect 9212 25228 9604 25284
rect 1820 24276 1876 25200
rect 1820 24220 2324 24276
rect 2044 24052 2100 24062
rect 1932 22036 1988 22046
rect 1932 21474 1988 21980
rect 1932 21422 1934 21474
rect 1986 21422 1988 21474
rect 1932 21410 1988 21422
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20020 1988 20862
rect 1932 19954 1988 19964
rect 2044 19906 2100 23996
rect 2268 22594 2324 24220
rect 5404 23492 5460 25200
rect 8988 25060 9044 25200
rect 9212 25060 9268 25228
rect 8988 25004 9268 25060
rect 5404 23426 5460 23436
rect 6636 23492 6692 23502
rect 5370 22764 5634 22774
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5370 22698 5634 22708
rect 2268 22542 2270 22594
rect 2322 22542 2324 22594
rect 2268 22530 2324 22542
rect 6636 22594 6692 23436
rect 6636 22542 6638 22594
rect 6690 22542 6692 22594
rect 6636 22530 6692 22542
rect 9548 22594 9604 25228
rect 12544 25200 12656 26000
rect 16128 25200 16240 26000
rect 19712 25200 19824 26000
rect 23296 25200 23408 26000
rect 26880 25200 26992 26000
rect 30464 25200 30576 26000
rect 34048 25200 34160 26000
rect 9548 22542 9550 22594
rect 9602 22542 9604 22594
rect 9548 22530 9604 22542
rect 12572 22596 12628 25200
rect 13686 22764 13950 22774
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13686 22698 13950 22708
rect 12572 22530 12628 22540
rect 14140 22596 14196 22606
rect 14140 22502 14196 22540
rect 16156 22596 16212 25200
rect 16156 22530 16212 22540
rect 17164 22596 17220 22606
rect 17164 22502 17220 22540
rect 19740 22596 19796 25200
rect 22002 22764 22266 22774
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22002 22698 22266 22708
rect 19740 22530 19796 22540
rect 20972 22596 21028 22606
rect 20972 22502 21028 22540
rect 23324 22596 23380 25200
rect 23324 22530 23380 22540
rect 25116 23156 25172 23166
rect 4172 22372 4228 22382
rect 4060 22370 4228 22372
rect 4060 22318 4174 22370
rect 4226 22318 4228 22370
rect 4060 22316 4228 22318
rect 4060 21476 4116 22316
rect 4172 22306 4228 22316
rect 5964 22370 6020 22382
rect 11452 22372 11508 22382
rect 13132 22372 13188 22382
rect 5964 22318 5966 22370
rect 6018 22318 6020 22370
rect 4284 21588 4340 21598
rect 4620 21588 4676 21598
rect 4284 21586 4676 21588
rect 4284 21534 4286 21586
rect 4338 21534 4622 21586
rect 4674 21534 4676 21586
rect 4284 21532 4676 21534
rect 4284 21522 4340 21532
rect 4620 21522 4676 21532
rect 2044 19854 2046 19906
rect 2098 19854 2100 19906
rect 2044 19842 2100 19854
rect 2716 20804 2772 20814
rect 2716 19458 2772 20748
rect 3836 20804 3892 20814
rect 3836 20710 3892 20748
rect 2716 19406 2718 19458
rect 2770 19406 2772 19458
rect 2716 19394 2772 19406
rect 2828 19122 2884 19134
rect 2828 19070 2830 19122
rect 2882 19070 2884 19122
rect 2156 18450 2212 18462
rect 2156 18398 2158 18450
rect 2210 18398 2212 18450
rect 1708 16658 1764 16670
rect 1708 16606 1710 16658
rect 1762 16606 1764 16658
rect 1708 15316 1764 16606
rect 1932 16212 1988 16222
rect 1932 16118 1988 16156
rect 1708 15250 1764 15260
rect 1820 14530 1876 14542
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 13972 1876 14478
rect 2044 14532 2100 14542
rect 2044 14418 2100 14476
rect 2044 14366 2046 14418
rect 2098 14366 2100 14418
rect 2044 14354 2100 14366
rect 1820 13878 1876 13916
rect 1820 12180 1876 12190
rect 2044 12180 2100 12190
rect 1820 12178 2044 12180
rect 1820 12126 1822 12178
rect 1874 12126 2044 12178
rect 1820 12124 2044 12126
rect 1820 12114 1876 12124
rect 2044 12114 2100 12124
rect 1932 11956 1988 11966
rect 1932 11618 1988 11900
rect 1932 11566 1934 11618
rect 1986 11566 1988 11618
rect 1932 11554 1988 11566
rect 1932 10386 1988 10398
rect 1932 10334 1934 10386
rect 1986 10334 1988 10386
rect 1932 9940 1988 10334
rect 2156 10050 2212 18398
rect 2716 18228 2772 18238
rect 2716 18134 2772 18172
rect 2716 16884 2772 16894
rect 2716 16790 2772 16828
rect 2604 14532 2660 14542
rect 2604 14438 2660 14476
rect 2492 13748 2548 13758
rect 2492 13634 2548 13692
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13570 2548 13582
rect 2828 13188 2884 19070
rect 3388 15428 3444 15438
rect 3388 15426 3780 15428
rect 3388 15374 3390 15426
rect 3442 15374 3780 15426
rect 3388 15372 3780 15374
rect 3388 15362 3444 15372
rect 3612 15202 3668 15214
rect 3612 15150 3614 15202
rect 3666 15150 3668 15202
rect 3276 14532 3332 14542
rect 3276 14438 3332 14476
rect 2940 14420 2996 14430
rect 2940 14326 2996 14364
rect 3612 14420 3668 15150
rect 3724 15148 3780 15372
rect 3836 15316 3892 15326
rect 3836 15222 3892 15260
rect 3724 15092 3892 15148
rect 3612 14354 3668 14364
rect 3836 14530 3892 15092
rect 3836 14478 3838 14530
rect 3890 14478 3892 14530
rect 3836 14084 3892 14478
rect 3836 14018 3892 14028
rect 3948 14980 4004 14990
rect 2940 13972 2996 13982
rect 2940 13878 2996 13916
rect 3388 13860 3444 13870
rect 3388 13766 3444 13804
rect 3164 13188 3220 13198
rect 2828 13132 2996 13188
rect 2268 12404 2324 12414
rect 2268 12178 2324 12348
rect 2268 12126 2270 12178
rect 2322 12126 2324 12178
rect 2268 12114 2324 12126
rect 2156 9998 2158 10050
rect 2210 9998 2212 10050
rect 2156 9986 2212 9998
rect 1932 9874 1988 9884
rect 2716 9826 2772 9838
rect 2716 9774 2718 9826
rect 2770 9774 2772 9826
rect 2268 9716 2324 9726
rect 2268 9714 2436 9716
rect 2268 9662 2270 9714
rect 2322 9662 2436 9714
rect 2268 9660 2436 9662
rect 2268 9650 2324 9660
rect 2268 9042 2324 9054
rect 2268 8990 2270 9042
rect 2322 8990 2324 9042
rect 1820 8932 1876 8942
rect 1820 8838 1876 8876
rect 1932 8370 1988 8382
rect 1932 8318 1934 8370
rect 1986 8318 1988 8370
rect 1932 7924 1988 8318
rect 1932 7858 1988 7868
rect 2044 7476 2100 7486
rect 2044 7474 2212 7476
rect 2044 7422 2046 7474
rect 2098 7422 2212 7474
rect 2044 7420 2212 7422
rect 2044 7410 2100 7420
rect 2156 6692 2212 7420
rect 2268 7028 2324 8990
rect 2380 8260 2436 9660
rect 2716 9604 2772 9774
rect 2940 9716 2996 13132
rect 2940 9622 2996 9660
rect 3052 13074 3108 13086
rect 3052 13022 3054 13074
rect 3106 13022 3108 13074
rect 3052 12180 3108 13022
rect 3164 12962 3220 13132
rect 3164 12910 3166 12962
rect 3218 12910 3220 12962
rect 3164 12898 3220 12910
rect 2716 9538 2772 9548
rect 3052 9044 3108 12124
rect 3276 12738 3332 12750
rect 3276 12686 3278 12738
rect 3330 12686 3332 12738
rect 3276 11396 3332 12686
rect 3276 11330 3332 11340
rect 3836 11396 3892 11406
rect 3836 11302 3892 11340
rect 3836 10612 3892 10622
rect 3388 10610 3892 10612
rect 3388 10558 3838 10610
rect 3890 10558 3892 10610
rect 3388 10556 3892 10558
rect 3388 10050 3444 10556
rect 3836 10546 3892 10556
rect 3388 9998 3390 10050
rect 3442 9998 3444 10050
rect 3388 9986 3444 9998
rect 3276 9940 3332 9950
rect 3276 9846 3332 9884
rect 3836 9940 3892 9950
rect 3948 9940 4004 14924
rect 4060 13748 4116 21420
rect 4732 21474 4788 21486
rect 4732 21422 4734 21474
rect 4786 21422 4788 21474
rect 4284 21364 4340 21374
rect 4284 20018 4340 21308
rect 4732 20914 4788 21422
rect 5180 21476 5236 21486
rect 5628 21476 5684 21486
rect 5180 21474 5684 21476
rect 5180 21422 5182 21474
rect 5234 21422 5630 21474
rect 5682 21422 5684 21474
rect 5180 21420 5684 21422
rect 5068 21364 5124 21374
rect 5068 21270 5124 21308
rect 4732 20862 4734 20914
rect 4786 20862 4788 20914
rect 4732 20188 4788 20862
rect 5180 20188 5236 21420
rect 5628 21410 5684 21420
rect 5370 21196 5634 21206
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5370 21130 5634 21140
rect 4732 20132 4900 20188
rect 4284 19966 4286 20018
rect 4338 19966 4340 20018
rect 4284 19954 4340 19966
rect 4284 16100 4340 16110
rect 4732 16100 4788 16110
rect 4284 16098 4788 16100
rect 4284 16046 4286 16098
rect 4338 16046 4734 16098
rect 4786 16046 4788 16098
rect 4284 16044 4788 16046
rect 4172 15090 4228 15102
rect 4172 15038 4174 15090
rect 4226 15038 4228 15090
rect 4172 14756 4228 15038
rect 4284 14980 4340 16044
rect 4732 16034 4788 16044
rect 4620 15316 4676 15326
rect 4620 15204 4676 15260
rect 4396 15202 4676 15204
rect 4396 15150 4622 15202
rect 4674 15150 4676 15202
rect 4396 15148 4676 15150
rect 4396 15092 4788 15148
rect 4284 14914 4340 14924
rect 4396 14756 4452 14766
rect 4732 14756 4788 15092
rect 4172 14700 4340 14756
rect 4284 14532 4340 14700
rect 4396 14754 4788 14756
rect 4396 14702 4398 14754
rect 4450 14702 4788 14754
rect 4396 14700 4788 14702
rect 4396 14690 4452 14700
rect 4284 14466 4340 14476
rect 4172 14420 4228 14430
rect 4172 14326 4228 14364
rect 4732 14308 4788 14318
rect 4732 14214 4788 14252
rect 4396 14084 4452 14094
rect 4396 13858 4452 14028
rect 4396 13806 4398 13858
rect 4450 13806 4452 13858
rect 4396 13794 4452 13806
rect 4172 13748 4228 13758
rect 4060 13692 4172 13748
rect 3892 9884 4004 9940
rect 3836 9846 3892 9884
rect 4060 9716 4116 9726
rect 3052 8950 3108 8988
rect 3500 9042 3556 9054
rect 3500 8990 3502 9042
rect 3554 8990 3556 9042
rect 3500 8372 3556 8990
rect 3500 8306 3556 8316
rect 3948 8932 4004 8942
rect 2380 8194 2436 8204
rect 3836 8260 3892 8270
rect 3836 8166 3892 8204
rect 2268 6962 2324 6972
rect 2492 7474 2548 7486
rect 2492 7422 2494 7474
rect 2546 7422 2548 7474
rect 2492 6916 2548 7422
rect 2492 6850 2548 6860
rect 2156 5908 2212 6636
rect 2940 6804 2996 6814
rect 2492 6578 2548 6590
rect 2492 6526 2494 6578
rect 2546 6526 2548 6578
rect 2268 5908 2324 5918
rect 2156 5906 2324 5908
rect 2156 5854 2270 5906
rect 2322 5854 2324 5906
rect 2156 5852 2324 5854
rect 2268 5842 2324 5852
rect 2492 5908 2548 6526
rect 2492 5842 2548 5852
rect 2940 5906 2996 6748
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 2940 5842 2996 5854
rect 3948 5796 4004 8876
rect 4060 6690 4116 9660
rect 4060 6638 4062 6690
rect 4114 6638 4116 6690
rect 4060 6626 4116 6638
rect 3276 4900 3332 4910
rect 3276 4898 3444 4900
rect 3276 4846 3278 4898
rect 3330 4846 3444 4898
rect 3276 4844 3444 4846
rect 3276 4834 3332 4844
rect 1932 4116 1988 4126
rect 1932 4022 1988 4060
rect 2268 3666 2324 3678
rect 2268 3614 2270 3666
rect 2322 3614 2324 3666
rect 2268 3388 2324 3614
rect 1820 3332 2324 3388
rect 1820 800 1876 3332
rect 3388 1876 3444 4844
rect 3948 4338 4004 5740
rect 4172 5236 4228 13692
rect 4620 13746 4676 13758
rect 4620 13694 4622 13746
rect 4674 13694 4676 13746
rect 4620 13636 4676 13694
rect 4620 13570 4676 13580
rect 4508 12180 4564 12190
rect 4508 12086 4564 12124
rect 4732 9940 4788 9950
rect 4620 8260 4676 8270
rect 4620 8146 4676 8204
rect 4620 8094 4622 8146
rect 4674 8094 4676 8146
rect 4620 8082 4676 8094
rect 4732 7252 4788 9884
rect 4844 8932 4900 20132
rect 5068 20132 5236 20188
rect 5852 20802 5908 20814
rect 5852 20750 5854 20802
rect 5906 20750 5908 20802
rect 4956 16884 5012 16894
rect 4956 16790 5012 16828
rect 4956 15314 5012 15326
rect 4956 15262 4958 15314
rect 5010 15262 5012 15314
rect 4956 14084 5012 15262
rect 4956 14018 5012 14028
rect 4844 8866 4900 8876
rect 4956 8036 5012 8046
rect 4956 7942 5012 7980
rect 4732 7186 4788 7196
rect 4844 7698 4900 7710
rect 4844 7646 4846 7698
rect 4898 7646 4900 7698
rect 4844 6914 4900 7646
rect 5068 7252 5124 20132
rect 5370 19628 5634 19638
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5370 19562 5634 19572
rect 5628 19236 5684 19246
rect 5852 19236 5908 20750
rect 5628 19234 5908 19236
rect 5628 19182 5630 19234
rect 5682 19182 5908 19234
rect 5628 19180 5908 19182
rect 5628 18228 5684 19180
rect 5964 18674 6020 22318
rect 11004 22370 11508 22372
rect 11004 22318 11454 22370
rect 11506 22318 11508 22370
rect 11004 22316 11508 22318
rect 9528 21980 9792 21990
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9528 21914 9792 21924
rect 8988 21812 9044 21822
rect 8988 21698 9044 21756
rect 10332 21812 10388 21822
rect 10668 21812 10724 21822
rect 10332 21810 10724 21812
rect 10332 21758 10334 21810
rect 10386 21758 10670 21810
rect 10722 21758 10724 21810
rect 10332 21756 10724 21758
rect 10332 21746 10388 21756
rect 10668 21746 10724 21756
rect 11004 21812 11060 22316
rect 11452 22306 11508 22316
rect 12572 22370 13188 22372
rect 12572 22318 13134 22370
rect 13186 22318 13188 22370
rect 12572 22316 13188 22318
rect 12572 21812 12628 22316
rect 13132 22306 13188 22316
rect 19068 22370 19124 22382
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 19068 22148 19124 22318
rect 23324 22370 23380 22382
rect 23324 22318 23326 22370
rect 23378 22318 23380 22370
rect 19964 22148 20020 22158
rect 19068 22146 20020 22148
rect 19068 22094 19966 22146
rect 20018 22094 20020 22146
rect 19068 22092 20020 22094
rect 17844 21980 18108 21990
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 17844 21914 18108 21924
rect 11004 21718 11060 21756
rect 12124 21810 12628 21812
rect 12124 21758 12574 21810
rect 12626 21758 12628 21810
rect 12124 21756 12628 21758
rect 8988 21646 8990 21698
rect 9042 21646 9044 21698
rect 8988 21634 9044 21646
rect 12124 21698 12180 21756
rect 12572 21746 12628 21756
rect 12908 21812 12964 21822
rect 12908 21718 12964 21756
rect 17388 21812 17444 21822
rect 19068 21812 19124 22092
rect 19964 22082 20020 22092
rect 23324 22148 23380 22318
rect 24556 22370 24612 22382
rect 24556 22318 24558 22370
rect 24610 22318 24612 22370
rect 23324 22082 23380 22092
rect 23772 22148 23828 22158
rect 23772 22054 23828 22092
rect 17388 21718 17444 21756
rect 18844 21756 19124 21812
rect 20636 21812 20692 21822
rect 20636 21810 21588 21812
rect 20636 21758 20638 21810
rect 20690 21758 21588 21810
rect 20636 21756 21588 21758
rect 12124 21646 12126 21698
rect 12178 21646 12180 21698
rect 12124 21634 12180 21646
rect 16156 21698 16212 21710
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 13244 21586 13300 21598
rect 13244 21534 13246 21586
rect 13298 21534 13300 21586
rect 6076 21476 6132 21486
rect 6076 21382 6132 21420
rect 9772 21476 9828 21486
rect 9772 21474 9940 21476
rect 9772 21422 9774 21474
rect 9826 21422 9940 21474
rect 9772 21420 9940 21422
rect 9772 21410 9828 21420
rect 8876 21362 8932 21374
rect 8876 21310 8878 21362
rect 8930 21310 8932 21362
rect 6524 20802 6580 20814
rect 6524 20750 6526 20802
rect 6578 20750 6580 20802
rect 6524 20132 6580 20750
rect 6524 20066 6580 20076
rect 8764 20578 8820 20590
rect 8764 20526 8766 20578
rect 8818 20526 8820 20578
rect 6188 19236 6244 19246
rect 6188 19234 6580 19236
rect 6188 19182 6190 19234
rect 6242 19182 6580 19234
rect 6188 19180 6580 19182
rect 6188 19170 6244 19180
rect 5964 18622 5966 18674
rect 6018 18622 6020 18674
rect 5740 18452 5796 18462
rect 5964 18452 6020 18622
rect 6412 18452 6468 18462
rect 5964 18450 6468 18452
rect 5964 18398 6414 18450
rect 6466 18398 6468 18450
rect 5964 18396 6468 18398
rect 5740 18358 5796 18396
rect 6412 18386 6468 18396
rect 6300 18228 6356 18238
rect 5628 18172 5796 18228
rect 5370 18060 5634 18070
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5370 17994 5634 18004
rect 5516 16884 5572 16894
rect 5740 16884 5796 18172
rect 5516 16882 5796 16884
rect 5516 16830 5518 16882
rect 5570 16830 5796 16882
rect 5516 16828 5796 16830
rect 5964 18226 6356 18228
rect 5964 18174 6302 18226
rect 6354 18174 6356 18226
rect 5964 18172 6356 18174
rect 5516 16660 5572 16828
rect 5516 16594 5572 16604
rect 5370 16492 5634 16502
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5370 16426 5634 16436
rect 5852 15316 5908 15326
rect 5370 14924 5634 14934
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5370 14858 5634 14868
rect 5516 14530 5572 14542
rect 5516 14478 5518 14530
rect 5570 14478 5572 14530
rect 5516 14308 5572 14478
rect 5852 14530 5908 15260
rect 5852 14478 5854 14530
rect 5906 14478 5908 14530
rect 5852 14466 5908 14478
rect 5516 14242 5572 14252
rect 5740 14306 5796 14318
rect 5740 14254 5742 14306
rect 5794 14254 5796 14306
rect 5740 13858 5796 14254
rect 5964 13860 6020 18172
rect 6300 18162 6356 18172
rect 6524 17892 6580 19180
rect 8652 19012 8708 19022
rect 8764 19012 8820 20526
rect 8652 19010 8820 19012
rect 8652 18958 8654 19010
rect 8706 18958 8820 19010
rect 8652 18956 8820 18958
rect 8428 18340 8484 18350
rect 8428 18246 8484 18284
rect 6524 17826 6580 17836
rect 8652 16996 8708 18956
rect 8764 18676 8820 18686
rect 8764 18450 8820 18620
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8764 18386 8820 18398
rect 8652 16930 8708 16940
rect 6860 16882 6916 16894
rect 6860 16830 6862 16882
rect 6914 16830 6916 16882
rect 6188 15986 6244 15998
rect 6188 15934 6190 15986
rect 6242 15934 6244 15986
rect 6188 15148 6244 15934
rect 6300 15876 6356 15886
rect 6300 15782 6356 15820
rect 6412 15874 6468 15886
rect 6412 15822 6414 15874
rect 6466 15822 6468 15874
rect 6412 15540 6468 15822
rect 6412 15484 6692 15540
rect 6412 15316 6468 15326
rect 6412 15222 6468 15260
rect 6188 15092 6580 15148
rect 6076 14532 6132 14542
rect 6076 14438 6132 14476
rect 6524 14530 6580 15092
rect 6524 14478 6526 14530
rect 6578 14478 6580 14530
rect 6524 14420 6580 14478
rect 6524 14354 6580 14364
rect 6636 14644 6692 15484
rect 6860 15426 6916 16830
rect 6972 16884 7028 16894
rect 6972 16790 7028 16828
rect 7196 16882 7252 16894
rect 7196 16830 7198 16882
rect 7250 16830 7252 16882
rect 7196 16100 7252 16830
rect 7420 16882 7476 16894
rect 7420 16830 7422 16882
rect 7474 16830 7476 16882
rect 7420 16210 7476 16830
rect 7420 16158 7422 16210
rect 7474 16158 7476 16210
rect 7420 16146 7476 16158
rect 7980 16660 8036 16670
rect 7196 16034 7252 16044
rect 7532 15988 7588 15998
rect 7532 15894 7588 15932
rect 7196 15876 7252 15886
rect 7196 15538 7252 15820
rect 7196 15486 7198 15538
rect 7250 15486 7252 15538
rect 7196 15474 7252 15486
rect 7308 15874 7364 15886
rect 7308 15822 7310 15874
rect 7362 15822 7364 15874
rect 7308 15540 7364 15822
rect 7308 15474 7364 15484
rect 7084 15428 7140 15438
rect 6860 15374 6862 15426
rect 6914 15374 6916 15426
rect 6860 15362 6916 15374
rect 6972 15372 7084 15428
rect 6972 15148 7028 15372
rect 7084 15362 7140 15372
rect 7644 15428 7700 15438
rect 7644 15334 7700 15372
rect 7308 15316 7364 15326
rect 7308 15222 7364 15260
rect 7420 15314 7476 15326
rect 7420 15262 7422 15314
rect 7474 15262 7476 15314
rect 6636 14418 6692 14588
rect 6860 15092 7028 15148
rect 6860 14530 6916 15092
rect 6860 14478 6862 14530
rect 6914 14478 6916 14530
rect 6860 14466 6916 14478
rect 6636 14366 6638 14418
rect 6690 14366 6692 14418
rect 6636 14354 6692 14366
rect 6524 13972 6580 13982
rect 6524 13878 6580 13916
rect 7420 13972 7476 15262
rect 7644 14308 7700 14318
rect 7420 13906 7476 13916
rect 7532 14252 7644 14308
rect 7532 14084 7588 14252
rect 7644 14214 7700 14252
rect 7532 13970 7588 14028
rect 7532 13918 7534 13970
rect 7586 13918 7588 13970
rect 7532 13906 7588 13918
rect 7980 13972 8036 16604
rect 8092 14644 8148 14654
rect 8092 14550 8148 14588
rect 8540 14418 8596 14430
rect 8540 14366 8542 14418
rect 8594 14366 8596 14418
rect 8092 13972 8148 13982
rect 7980 13970 8148 13972
rect 7980 13918 8094 13970
rect 8146 13918 8148 13970
rect 7980 13916 8148 13918
rect 5740 13806 5742 13858
rect 5794 13806 5796 13858
rect 5740 13794 5796 13806
rect 5852 13804 6020 13860
rect 5852 13636 5908 13804
rect 4844 6862 4846 6914
rect 4898 6862 4900 6914
rect 4844 6850 4900 6862
rect 4956 7196 5124 7252
rect 5180 13580 5908 13636
rect 5964 13634 6020 13646
rect 6412 13636 6468 13646
rect 5964 13582 5966 13634
rect 6018 13582 6020 13634
rect 5180 7252 5236 13580
rect 5370 13356 5634 13366
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5370 13290 5634 13300
rect 5628 12962 5684 12974
rect 5628 12910 5630 12962
rect 5682 12910 5684 12962
rect 5404 12852 5460 12862
rect 5404 12402 5460 12796
rect 5404 12350 5406 12402
rect 5458 12350 5460 12402
rect 5404 12338 5460 12350
rect 5628 12402 5684 12910
rect 5628 12350 5630 12402
rect 5682 12350 5684 12402
rect 5628 12338 5684 12350
rect 5852 12852 5908 12862
rect 5852 12402 5908 12796
rect 5964 12628 6020 13582
rect 6076 13634 6468 13636
rect 6076 13582 6414 13634
rect 6466 13582 6468 13634
rect 6076 13580 6468 13582
rect 6076 12964 6132 13580
rect 6412 13570 6468 13580
rect 7084 13636 7140 13646
rect 7140 13580 7252 13636
rect 7084 13542 7140 13580
rect 6076 12870 6132 12908
rect 6188 12738 6244 12750
rect 6188 12686 6190 12738
rect 6242 12686 6244 12738
rect 5964 12572 6132 12628
rect 5852 12350 5854 12402
rect 5906 12350 5908 12402
rect 5852 12338 5908 12350
rect 5964 12292 6020 12302
rect 5964 12198 6020 12236
rect 6076 12180 6132 12572
rect 6188 12404 6244 12686
rect 6300 12738 6356 12750
rect 6300 12686 6302 12738
rect 6354 12686 6356 12738
rect 6300 12628 6356 12686
rect 6300 12562 6356 12572
rect 6860 12738 6916 12750
rect 6860 12686 6862 12738
rect 6914 12686 6916 12738
rect 6860 12628 6916 12686
rect 6188 12338 6244 12348
rect 6524 12292 6580 12302
rect 6524 12198 6580 12236
rect 6300 12180 6356 12190
rect 6076 12178 6356 12180
rect 6076 12126 6302 12178
rect 6354 12126 6356 12178
rect 6076 12124 6356 12126
rect 6300 12114 6356 12124
rect 6412 12066 6468 12078
rect 6412 12014 6414 12066
rect 6466 12014 6468 12066
rect 5370 11788 5634 11798
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5370 11722 5634 11732
rect 6412 11732 6468 12014
rect 6860 12068 6916 12572
rect 7196 12404 7252 13580
rect 7980 12962 8036 13916
rect 8092 13906 8148 13916
rect 8540 13972 8596 14366
rect 8540 13906 8596 13916
rect 8316 13748 8372 13758
rect 8316 13654 8372 13692
rect 7980 12910 7982 12962
rect 8034 12910 8036 12962
rect 7980 12898 8036 12910
rect 8428 12962 8484 12974
rect 8428 12910 8430 12962
rect 8482 12910 8484 12962
rect 8428 12740 8484 12910
rect 8428 12674 8484 12684
rect 7308 12404 7364 12414
rect 7196 12348 7308 12404
rect 7308 12310 7364 12348
rect 7868 12404 7924 12414
rect 7868 12310 7924 12348
rect 7084 12290 7140 12302
rect 7084 12238 7086 12290
rect 7138 12238 7140 12290
rect 6972 12180 7028 12190
rect 7084 12180 7140 12238
rect 6972 12178 7140 12180
rect 6972 12126 6974 12178
rect 7026 12126 7140 12178
rect 6972 12124 7140 12126
rect 7420 12178 7476 12190
rect 7420 12126 7422 12178
rect 7474 12126 7476 12178
rect 6972 12114 7028 12124
rect 6860 12002 6916 12012
rect 7420 12068 7476 12126
rect 7420 12002 7476 12012
rect 8316 12068 8372 12078
rect 6412 11676 6916 11732
rect 6524 11394 6580 11406
rect 6524 11342 6526 11394
rect 6578 11342 6580 11394
rect 5370 10220 5634 10230
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5370 10154 5634 10164
rect 6524 9828 6580 11342
rect 6860 11394 6916 11676
rect 6860 11342 6862 11394
rect 6914 11342 6916 11394
rect 6860 11330 6916 11342
rect 8316 9940 8372 12012
rect 8316 9874 8372 9884
rect 6524 9762 6580 9772
rect 6860 9828 6916 9838
rect 7980 9828 8036 9838
rect 6860 9826 7028 9828
rect 6860 9774 6862 9826
rect 6914 9774 7028 9826
rect 6860 9772 7028 9774
rect 6860 9762 6916 9772
rect 6524 9604 6580 9614
rect 6524 9510 6580 9548
rect 5964 9268 6020 9278
rect 6860 9268 6916 9278
rect 5964 9174 6020 9212
rect 6636 9266 6916 9268
rect 6636 9214 6862 9266
rect 6914 9214 6916 9266
rect 6636 9212 6916 9214
rect 6524 9156 6580 9166
rect 6524 9062 6580 9100
rect 5370 8652 5634 8662
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 6636 8596 6692 9212
rect 6860 9202 6916 9212
rect 5370 8586 5634 8596
rect 6412 8540 6692 8596
rect 6748 9042 6804 9054
rect 6748 8990 6750 9042
rect 6802 8990 6804 9042
rect 6076 8372 6132 8382
rect 6076 8278 6132 8316
rect 6412 8370 6468 8540
rect 6412 8318 6414 8370
rect 6466 8318 6468 8370
rect 6412 8306 6468 8318
rect 6188 8034 6244 8046
rect 6188 7982 6190 8034
rect 6242 7982 6244 8034
rect 6076 7698 6132 7710
rect 6076 7646 6078 7698
rect 6130 7646 6132 7698
rect 5964 7588 6020 7598
rect 5964 7494 6020 7532
rect 5516 7476 5572 7486
rect 5852 7476 5908 7486
rect 5516 7474 5852 7476
rect 5516 7422 5518 7474
rect 5570 7422 5852 7474
rect 5516 7420 5852 7422
rect 5516 7410 5572 7420
rect 5852 7382 5908 7420
rect 5180 7196 5908 7252
rect 4732 6692 4788 6702
rect 4956 6692 5012 7196
rect 5370 7084 5634 7094
rect 4172 5170 4228 5180
rect 4284 6690 5012 6692
rect 4284 6638 4734 6690
rect 4786 6638 5012 6690
rect 4284 6636 5012 6638
rect 5068 7028 5124 7038
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5370 7018 5634 7028
rect 4284 5124 4340 6636
rect 4732 6626 4788 6636
rect 5068 5348 5124 6972
rect 5628 6916 5684 6926
rect 5628 6822 5684 6860
rect 5180 6690 5236 6702
rect 5180 6638 5182 6690
rect 5234 6638 5236 6690
rect 5180 6468 5236 6638
rect 5180 6130 5236 6412
rect 5180 6078 5182 6130
rect 5234 6078 5236 6130
rect 5180 6066 5236 6078
rect 5740 6466 5796 6478
rect 5740 6414 5742 6466
rect 5794 6414 5796 6466
rect 5740 6132 5796 6414
rect 5740 6066 5796 6076
rect 5370 5516 5634 5526
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5370 5450 5634 5460
rect 5740 5348 5796 5358
rect 5068 5346 5796 5348
rect 5068 5294 5742 5346
rect 5794 5294 5796 5346
rect 5068 5292 5796 5294
rect 5740 5282 5796 5292
rect 4732 5236 4788 5246
rect 4732 5142 4788 5180
rect 5628 5124 5684 5134
rect 4284 5122 4452 5124
rect 4284 5070 4286 5122
rect 4338 5070 4452 5122
rect 4284 5068 4452 5070
rect 4284 5058 4340 5068
rect 3948 4286 3950 4338
rect 4002 4286 4004 4338
rect 3948 4274 4004 4286
rect 4396 4340 4452 5068
rect 4620 4900 4676 4910
rect 4620 4898 4788 4900
rect 4620 4846 4622 4898
rect 4674 4846 4788 4898
rect 4620 4844 4788 4846
rect 4620 4834 4676 4844
rect 4620 4340 4676 4350
rect 4396 4338 4676 4340
rect 4396 4286 4622 4338
rect 4674 4286 4676 4338
rect 4396 4284 4676 4286
rect 4620 4274 4676 4284
rect 4620 3556 4676 3566
rect 4732 3556 4788 4844
rect 5180 4338 5236 4350
rect 5180 4286 5182 4338
rect 5234 4286 5236 4338
rect 5180 4228 5236 4286
rect 5628 4338 5684 5068
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 5628 4274 5684 4286
rect 5180 4162 5236 4172
rect 5370 3948 5634 3958
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5370 3882 5634 3892
rect 4620 3554 4788 3556
rect 4620 3502 4622 3554
rect 4674 3502 4788 3554
rect 4620 3500 4788 3502
rect 5852 3556 5908 7196
rect 5964 6916 6020 6926
rect 6076 6916 6132 7646
rect 5964 6914 6132 6916
rect 5964 6862 5966 6914
rect 6018 6862 6132 6914
rect 5964 6860 6132 6862
rect 5964 6850 6020 6860
rect 6188 6468 6244 7982
rect 6636 8036 6692 8046
rect 6636 7698 6692 7980
rect 6636 7646 6638 7698
rect 6690 7646 6692 7698
rect 6636 7634 6692 7646
rect 6412 7474 6468 7486
rect 6412 7422 6414 7474
rect 6466 7422 6468 7474
rect 6412 6916 6468 7422
rect 6748 6916 6804 8990
rect 6972 9044 7028 9772
rect 7084 9716 7140 9726
rect 7084 9714 7252 9716
rect 7084 9662 7086 9714
rect 7138 9662 7252 9714
rect 7084 9660 7252 9662
rect 7084 9650 7140 9660
rect 7196 9156 7252 9660
rect 7084 9044 7140 9054
rect 6972 9042 7140 9044
rect 6972 8990 7086 9042
rect 7138 8990 7140 9042
rect 6972 8988 7140 8990
rect 7084 8932 7140 8988
rect 7196 9042 7252 9100
rect 7196 8990 7198 9042
rect 7250 8990 7252 9042
rect 7196 8978 7252 8990
rect 7532 9602 7588 9614
rect 7532 9550 7534 9602
rect 7586 9550 7588 9602
rect 7532 8932 7588 9550
rect 7756 8932 7812 8942
rect 7532 8876 7756 8932
rect 7084 8866 7140 8876
rect 7756 8838 7812 8876
rect 7196 7588 7252 7598
rect 7196 7494 7252 7532
rect 6972 7476 7028 7486
rect 6972 7382 7028 7420
rect 6412 6860 6804 6916
rect 6300 6804 6356 6814
rect 6300 6710 6356 6748
rect 6636 6578 6692 6590
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 6412 6468 6468 6478
rect 6188 6466 6468 6468
rect 6188 6414 6414 6466
rect 6466 6414 6468 6466
rect 6188 6412 6468 6414
rect 6412 6132 6468 6412
rect 6412 6066 6468 6076
rect 6636 6130 6692 6526
rect 6636 6078 6638 6130
rect 6690 6078 6692 6130
rect 6636 6066 6692 6078
rect 6748 6020 6804 6860
rect 7756 6692 7812 6702
rect 7756 6598 7812 6636
rect 7420 6580 7476 6590
rect 6860 6020 6916 6030
rect 6748 5964 6860 6020
rect 5964 5908 6020 5918
rect 6188 5908 6244 5918
rect 6524 5908 6580 5918
rect 5964 5906 6244 5908
rect 5964 5854 5966 5906
rect 6018 5854 6190 5906
rect 6242 5854 6244 5906
rect 5964 5852 6244 5854
rect 5964 5842 6020 5852
rect 5964 5684 6020 5694
rect 5964 4338 6020 5628
rect 6076 5346 6132 5852
rect 6188 5842 6244 5852
rect 6300 5852 6524 5908
rect 6076 5294 6078 5346
rect 6130 5294 6132 5346
rect 6076 5282 6132 5294
rect 6300 5234 6356 5852
rect 6524 5814 6580 5852
rect 6860 5906 6916 5964
rect 6860 5854 6862 5906
rect 6914 5854 6916 5906
rect 6860 5842 6916 5854
rect 7196 5796 7252 5806
rect 7196 5702 7252 5740
rect 6300 5182 6302 5234
rect 6354 5182 6356 5234
rect 6300 5170 6356 5182
rect 6748 5236 6804 5246
rect 6748 5142 6804 5180
rect 7420 5124 7476 6524
rect 7980 6580 8036 9772
rect 8540 9826 8596 9838
rect 8540 9774 8542 9826
rect 8594 9774 8596 9826
rect 8316 9604 8372 9614
rect 8540 9604 8596 9774
rect 8316 9602 8596 9604
rect 8316 9550 8318 9602
rect 8370 9550 8596 9602
rect 8316 9548 8596 9550
rect 8316 9044 8372 9548
rect 8316 8978 8372 8988
rect 8428 7364 8484 7374
rect 7980 6514 8036 6524
rect 8316 6692 8372 6702
rect 8316 6130 8372 6636
rect 8428 6690 8484 7308
rect 8428 6638 8430 6690
rect 8482 6638 8484 6690
rect 8428 6626 8484 6638
rect 8316 6078 8318 6130
rect 8370 6078 8372 6130
rect 7420 5010 7476 5068
rect 7756 5348 7812 5358
rect 7756 5122 7812 5292
rect 7756 5070 7758 5122
rect 7810 5070 7812 5122
rect 7756 5058 7812 5070
rect 8204 5124 8260 5134
rect 8316 5124 8372 6078
rect 8540 6580 8596 6590
rect 8540 5906 8596 6524
rect 8540 5854 8542 5906
rect 8594 5854 8596 5906
rect 8540 5842 8596 5854
rect 8764 5796 8820 5806
rect 8204 5122 8372 5124
rect 8204 5070 8206 5122
rect 8258 5070 8372 5122
rect 8204 5068 8372 5070
rect 8652 5124 8708 5134
rect 8764 5124 8820 5740
rect 8652 5122 8820 5124
rect 8652 5070 8654 5122
rect 8706 5070 8820 5122
rect 8652 5068 8820 5070
rect 8204 5058 8260 5068
rect 8652 5058 8708 5068
rect 7420 4958 7422 5010
rect 7474 4958 7476 5010
rect 7420 4946 7476 4958
rect 8540 5012 8596 5022
rect 8540 4562 8596 4956
rect 8540 4510 8542 4562
rect 8594 4510 8596 4562
rect 8540 4498 8596 4510
rect 5964 4286 5966 4338
rect 6018 4286 6020 4338
rect 5964 4274 6020 4286
rect 8876 3892 8932 21310
rect 9548 20916 9604 20926
rect 9772 20916 9828 20926
rect 9548 20914 9772 20916
rect 9548 20862 9550 20914
rect 9602 20862 9772 20914
rect 9548 20860 9772 20862
rect 9548 20850 9604 20860
rect 9772 20802 9828 20860
rect 9772 20750 9774 20802
rect 9826 20750 9828 20802
rect 9772 20738 9828 20750
rect 9884 20804 9940 21420
rect 9996 21362 10052 21374
rect 9996 21310 9998 21362
rect 10050 21310 10052 21362
rect 9996 21028 10052 21310
rect 9996 20962 10052 20972
rect 12236 21362 12292 21374
rect 12236 21310 12238 21362
rect 12290 21310 12292 21362
rect 9996 20804 10052 20814
rect 9884 20748 9996 20804
rect 9996 20710 10052 20748
rect 10444 20802 10500 20814
rect 10444 20750 10446 20802
rect 10498 20750 10500 20802
rect 10108 20578 10164 20590
rect 10108 20526 10110 20578
rect 10162 20526 10164 20578
rect 9528 20412 9792 20422
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9528 20346 9792 20356
rect 10108 20188 10164 20526
rect 9660 20130 9716 20142
rect 9660 20078 9662 20130
rect 9714 20078 9716 20130
rect 9660 19460 9716 20078
rect 9772 20132 9828 20142
rect 9772 20038 9828 20076
rect 9884 20132 10164 20188
rect 9884 20130 9940 20132
rect 9884 20078 9886 20130
rect 9938 20078 9940 20130
rect 9884 20066 9940 20078
rect 10444 20020 10500 20750
rect 10892 20578 10948 20590
rect 10892 20526 10894 20578
rect 10946 20526 10948 20578
rect 10332 19906 10388 19918
rect 10332 19854 10334 19906
rect 10386 19854 10388 19906
rect 10332 19460 10388 19854
rect 9660 19404 10388 19460
rect 9324 19292 9716 19348
rect 9212 19124 9268 19134
rect 9212 18788 9268 19068
rect 9212 18722 9268 18732
rect 8988 18564 9044 18574
rect 9324 18564 9380 19292
rect 9660 19234 9716 19292
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 9660 19170 9716 19182
rect 9436 19124 9492 19134
rect 9436 19030 9492 19068
rect 9884 19010 9940 19022
rect 9884 18958 9886 19010
rect 9938 18958 9940 19010
rect 9528 18844 9792 18854
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9528 18778 9792 18788
rect 9660 18676 9716 18686
rect 9660 18582 9716 18620
rect 8988 18562 9380 18564
rect 8988 18510 8990 18562
rect 9042 18510 9380 18562
rect 8988 18508 9380 18510
rect 8988 18498 9044 18508
rect 9100 18452 9156 18508
rect 9100 18386 9156 18396
rect 9884 18116 9940 18958
rect 9212 18060 9940 18116
rect 8988 17892 9044 17902
rect 8988 17778 9044 17836
rect 9212 17890 9268 18060
rect 9212 17838 9214 17890
rect 9266 17838 9268 17890
rect 9212 17826 9268 17838
rect 8988 17726 8990 17778
rect 9042 17726 9044 17778
rect 8988 17714 9044 17726
rect 8988 17556 9044 17566
rect 8988 17462 9044 17500
rect 9660 17556 9716 17566
rect 9996 17556 10052 19404
rect 10444 19348 10500 19964
rect 10108 19346 10500 19348
rect 10108 19294 10446 19346
rect 10498 19294 10500 19346
rect 10108 19292 10500 19294
rect 10108 19234 10164 19292
rect 10444 19282 10500 19292
rect 10556 20132 10612 20142
rect 10556 20018 10612 20076
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 19170 10164 19182
rect 10220 18452 10276 18462
rect 10556 18452 10612 19966
rect 10892 20020 10948 20526
rect 12236 20188 12292 21310
rect 12236 20132 12740 20188
rect 10892 19460 10948 19964
rect 11228 20020 11284 20030
rect 11228 19926 11284 19964
rect 12012 20020 12068 20030
rect 10892 19394 10948 19404
rect 12012 19458 12068 19964
rect 12012 19406 12014 19458
rect 12066 19406 12068 19458
rect 12012 19394 12068 19406
rect 12124 19908 12180 19918
rect 12124 19346 12180 19852
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 10892 19010 10948 19022
rect 10892 18958 10894 19010
rect 10946 18958 10948 19010
rect 10892 18676 10948 18958
rect 10892 18564 10948 18620
rect 10892 18508 11172 18564
rect 10220 18450 10612 18452
rect 10220 18398 10222 18450
rect 10274 18398 10612 18450
rect 10220 18396 10612 18398
rect 10668 18452 10724 18462
rect 10668 18450 10948 18452
rect 10668 18398 10670 18450
rect 10722 18398 10948 18450
rect 10668 18396 10948 18398
rect 10220 18386 10276 18396
rect 10668 18386 10724 18396
rect 10892 17890 10948 18396
rect 10892 17838 10894 17890
rect 10946 17838 10948 17890
rect 10892 17826 10948 17838
rect 11004 17668 11060 17678
rect 11004 17574 11060 17612
rect 10108 17556 10164 17566
rect 9996 17500 10108 17556
rect 9660 17462 9716 17500
rect 10108 17490 10164 17500
rect 9528 17276 9792 17286
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9528 17210 9792 17220
rect 10668 16996 10724 17006
rect 10444 16100 10500 16110
rect 10220 16098 10500 16100
rect 10220 16046 10446 16098
rect 10498 16046 10500 16098
rect 10220 16044 10500 16046
rect 9528 15708 9792 15718
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9528 15642 9792 15652
rect 10220 14642 10276 16044
rect 10444 16034 10500 16044
rect 10668 15148 10724 16940
rect 10780 16100 10836 16138
rect 10780 16034 10836 16044
rect 11004 16098 11060 16110
rect 11004 16046 11006 16098
rect 11058 16046 11060 16098
rect 10780 15876 10836 15886
rect 10780 15782 10836 15820
rect 10220 14590 10222 14642
rect 10274 14590 10276 14642
rect 10220 14578 10276 14590
rect 10444 15090 10500 15102
rect 10668 15092 10948 15148
rect 10444 15038 10446 15090
rect 10498 15038 10500 15090
rect 10444 14644 10500 15038
rect 10444 14578 10500 14588
rect 9996 14418 10052 14430
rect 9996 14366 9998 14418
rect 10050 14366 10052 14418
rect 9996 14308 10052 14366
rect 9996 14242 10052 14252
rect 9528 14140 9792 14150
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9528 14074 9792 14084
rect 10892 13746 10948 15092
rect 11004 14754 11060 16046
rect 11116 15428 11172 18508
rect 11676 18452 11732 18462
rect 11452 17666 11508 17678
rect 11452 17614 11454 17666
rect 11506 17614 11508 17666
rect 11452 17556 11508 17614
rect 11676 17666 11732 18396
rect 11676 17614 11678 17666
rect 11730 17614 11732 17666
rect 11676 17602 11732 17614
rect 11788 17668 11844 17678
rect 11788 17574 11844 17612
rect 12012 17666 12068 17678
rect 12012 17614 12014 17666
rect 12066 17614 12068 17666
rect 11452 17108 11508 17500
rect 11452 17042 11508 17052
rect 11116 15362 11172 15372
rect 11228 15988 11284 15998
rect 11004 14702 11006 14754
rect 11058 14702 11060 14754
rect 11004 14690 11060 14702
rect 11116 14644 11172 14654
rect 11116 14418 11172 14588
rect 11116 14366 11118 14418
rect 11170 14366 11172 14418
rect 11116 14354 11172 14366
rect 11228 14420 11284 15932
rect 12012 15988 12068 17614
rect 12348 17442 12404 17454
rect 12348 17390 12350 17442
rect 12402 17390 12404 17442
rect 12348 17108 12404 17390
rect 12348 17042 12404 17052
rect 12068 15932 12292 15988
rect 12012 15922 12068 15932
rect 11452 15316 11508 15326
rect 11452 15222 11508 15260
rect 11340 14420 11396 14430
rect 11228 14418 11396 14420
rect 11228 14366 11342 14418
rect 11394 14366 11396 14418
rect 11228 14364 11396 14366
rect 10892 13694 10894 13746
rect 10946 13694 10948 13746
rect 10892 12738 10948 13694
rect 10892 12686 10894 12738
rect 10946 12686 10948 12738
rect 10892 12674 10948 12686
rect 9528 12572 9792 12582
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9528 12506 9792 12516
rect 9996 12404 10052 12414
rect 9548 12290 9604 12302
rect 9548 12238 9550 12290
rect 9602 12238 9604 12290
rect 9212 12180 9268 12190
rect 9212 11282 9268 12124
rect 9548 12180 9604 12238
rect 9548 12114 9604 12124
rect 9884 12178 9940 12190
rect 9884 12126 9886 12178
rect 9938 12126 9940 12178
rect 9212 11230 9214 11282
rect 9266 11230 9268 11282
rect 9212 11218 9268 11230
rect 9528 11004 9792 11014
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9528 10938 9792 10948
rect 9212 9826 9268 9838
rect 9212 9774 9214 9826
rect 9266 9774 9268 9826
rect 9212 8372 9268 9774
rect 9528 9436 9792 9446
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9528 9370 9792 9380
rect 9212 8306 9268 8316
rect 9528 7868 9792 7878
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9528 7802 9792 7812
rect 9884 6468 9940 12126
rect 9996 11618 10052 12348
rect 9996 11566 9998 11618
rect 10050 11566 10052 11618
rect 9996 11554 10052 11566
rect 11228 11508 11284 14364
rect 11340 14354 11396 14364
rect 11452 13746 11508 13758
rect 11900 13748 11956 13758
rect 11452 13694 11454 13746
rect 11506 13694 11508 13746
rect 11452 13636 11508 13694
rect 11452 13570 11508 13580
rect 11564 13746 11956 13748
rect 11564 13694 11902 13746
rect 11954 13694 11956 13746
rect 11564 13692 11956 13694
rect 11452 13188 11508 13198
rect 11564 13188 11620 13692
rect 11900 13682 11956 13692
rect 11788 13522 11844 13534
rect 11788 13470 11790 13522
rect 11842 13470 11844 13522
rect 11452 13186 11620 13188
rect 11452 13134 11454 13186
rect 11506 13134 11620 13186
rect 11452 13132 11620 13134
rect 11676 13188 11732 13198
rect 11788 13188 11844 13470
rect 11732 13132 11844 13188
rect 11452 13122 11508 13132
rect 11676 13094 11732 13132
rect 12012 12962 12068 12974
rect 12012 12910 12014 12962
rect 12066 12910 12068 12962
rect 12012 12402 12068 12910
rect 12236 12964 12292 15932
rect 12348 13636 12404 13646
rect 12348 13542 12404 13580
rect 12460 13076 12516 13086
rect 12348 12964 12404 12974
rect 12236 12962 12404 12964
rect 12236 12910 12350 12962
rect 12402 12910 12404 12962
rect 12236 12908 12404 12910
rect 12348 12898 12404 12908
rect 12012 12350 12014 12402
rect 12066 12350 12068 12402
rect 12012 12338 12068 12350
rect 12124 12738 12180 12750
rect 12124 12686 12126 12738
rect 12178 12686 12180 12738
rect 11452 12292 11508 12302
rect 11452 12198 11508 12236
rect 11228 11442 11284 11452
rect 11340 12178 11396 12190
rect 11340 12126 11342 12178
rect 11394 12126 11396 12178
rect 11340 11284 11396 12126
rect 11564 12180 11620 12190
rect 11564 12086 11620 12124
rect 11340 10836 11396 11228
rect 12012 12068 12068 12078
rect 11676 10836 11732 10846
rect 11340 10834 11732 10836
rect 11340 10782 11678 10834
rect 11730 10782 11732 10834
rect 11340 10780 11732 10782
rect 11676 10770 11732 10780
rect 12012 10610 12068 12012
rect 12124 11732 12180 12686
rect 12236 12740 12292 12750
rect 12236 12646 12292 12684
rect 12460 12290 12516 13020
rect 12460 12238 12462 12290
rect 12514 12238 12516 12290
rect 12460 12226 12516 12238
rect 12348 12180 12404 12190
rect 12348 12086 12404 12124
rect 12124 11666 12180 11676
rect 12012 10558 12014 10610
rect 12066 10558 12068 10610
rect 12012 10546 12068 10558
rect 12572 10722 12628 10734
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12236 9940 12292 9950
rect 12572 9940 12628 10670
rect 12236 9938 12628 9940
rect 12236 9886 12238 9938
rect 12290 9886 12628 9938
rect 12236 9884 12628 9886
rect 12236 9874 12292 9884
rect 12572 9826 12628 9884
rect 12572 9774 12574 9826
rect 12626 9774 12628 9826
rect 12572 9762 12628 9774
rect 11452 9602 11508 9614
rect 11452 9550 11454 9602
rect 11506 9550 11508 9602
rect 11452 9268 11508 9550
rect 11508 9212 11620 9268
rect 11452 9202 11508 9212
rect 10892 8034 10948 8046
rect 10892 7982 10894 8034
rect 10946 7982 10948 8034
rect 10668 6468 10724 6478
rect 9884 6412 10052 6468
rect 9528 6300 9792 6310
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9528 6234 9792 6244
rect 9884 6244 9940 6254
rect 9660 6132 9716 6142
rect 9884 6132 9940 6188
rect 9716 6076 9940 6132
rect 9660 6038 9716 6076
rect 9548 5684 9604 5694
rect 9548 5590 9604 5628
rect 9884 5682 9940 5694
rect 9884 5630 9886 5682
rect 9938 5630 9940 5682
rect 9528 4732 9792 4742
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9528 4666 9792 4676
rect 9884 4564 9940 5630
rect 9996 5124 10052 6412
rect 10668 6374 10724 6412
rect 10892 6244 10948 7982
rect 11228 8036 11284 8046
rect 11228 7942 11284 7980
rect 11452 7588 11508 7598
rect 11452 6690 11508 7532
rect 11452 6638 11454 6690
rect 11506 6638 11508 6690
rect 11452 6626 11508 6638
rect 10668 6188 10948 6244
rect 11116 6468 11172 6478
rect 10668 6020 10724 6188
rect 9996 5068 10164 5124
rect 9884 4498 9940 4508
rect 9996 4900 10052 4910
rect 9100 4340 9156 4350
rect 9100 4246 9156 4284
rect 9884 4228 9940 4238
rect 9996 4228 10052 4844
rect 10108 4676 10164 5068
rect 10108 4340 10164 4620
rect 10668 4450 10724 5964
rect 11116 5906 11172 6412
rect 11116 5854 11118 5906
rect 11170 5854 11172 5906
rect 11116 4898 11172 5854
rect 11564 5906 11620 9212
rect 12684 8484 12740 20132
rect 13244 20132 13300 21534
rect 13916 21588 13972 21598
rect 13916 21586 14420 21588
rect 13916 21534 13918 21586
rect 13970 21534 14420 21586
rect 13916 21532 14420 21534
rect 13916 21522 13972 21532
rect 13686 21196 13950 21206
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13686 21130 13950 21140
rect 14364 21026 14420 21532
rect 14364 20974 14366 21026
rect 14418 20974 14420 21026
rect 14364 20962 14420 20974
rect 14252 20804 14308 20814
rect 14252 20242 14308 20748
rect 14812 20804 14868 20814
rect 14476 20692 14532 20702
rect 14476 20598 14532 20636
rect 14252 20190 14254 20242
rect 14306 20190 14308 20242
rect 14252 20178 14308 20190
rect 14812 20244 14868 20748
rect 15260 20804 15316 20814
rect 15260 20710 15316 20748
rect 15148 20692 15204 20702
rect 15148 20598 15204 20636
rect 15036 20578 15092 20590
rect 15036 20526 15038 20578
rect 15090 20526 15092 20578
rect 14924 20244 14980 20254
rect 14812 20242 14980 20244
rect 14812 20190 14926 20242
rect 14978 20190 14980 20242
rect 14812 20188 14980 20190
rect 14924 20178 14980 20188
rect 15036 20188 15092 20526
rect 15372 20578 15428 20590
rect 15372 20526 15374 20578
rect 15426 20526 15428 20578
rect 13244 20066 13300 20076
rect 13468 20132 13524 20142
rect 15036 20132 15204 20188
rect 13132 18676 13188 18686
rect 13468 18676 13524 20076
rect 14252 20020 14308 20030
rect 13686 19628 13950 19638
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13686 19562 13950 19572
rect 14252 19236 14308 19964
rect 14252 19122 14308 19180
rect 14252 19070 14254 19122
rect 14306 19070 14308 19122
rect 14252 19058 14308 19070
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 13132 18674 13524 18676
rect 13132 18622 13134 18674
rect 13186 18622 13524 18674
rect 13132 18620 13524 18622
rect 13132 18610 13188 18620
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 14476 18452 14532 19966
rect 14700 20018 14756 20030
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14476 18386 14532 18396
rect 14588 19122 14644 19134
rect 14588 19070 14590 19122
rect 14642 19070 14644 19122
rect 13686 18060 13950 18070
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13686 17994 13950 18004
rect 14588 17444 14644 19070
rect 14700 18676 14756 19966
rect 15036 20020 15092 20030
rect 15036 19926 15092 19964
rect 14812 19908 14868 19918
rect 14812 19814 14868 19852
rect 14812 19236 14868 19246
rect 14812 19142 14868 19180
rect 15148 19236 15204 20132
rect 15372 20020 15428 20526
rect 16156 20132 16212 21646
rect 17948 21474 18004 21486
rect 17948 21422 17950 21474
rect 18002 21422 18004 21474
rect 16940 21364 16996 21374
rect 16940 20804 16996 21308
rect 17724 21362 17780 21374
rect 17724 21310 17726 21362
rect 17778 21310 17780 21362
rect 17724 21028 17780 21310
rect 17948 21364 18004 21422
rect 17948 21298 18004 21308
rect 18508 21476 18564 21486
rect 18844 21476 18900 21756
rect 20636 21746 20692 21756
rect 18956 21588 19012 21598
rect 18956 21586 19236 21588
rect 18956 21534 18958 21586
rect 19010 21534 19236 21586
rect 18956 21532 19236 21534
rect 18956 21522 19012 21532
rect 18508 21474 18900 21476
rect 18508 21422 18510 21474
rect 18562 21422 18900 21474
rect 18508 21420 18900 21422
rect 17724 20962 17780 20972
rect 16940 20738 16996 20748
rect 17844 20412 18108 20422
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 17844 20346 18108 20356
rect 18508 20188 18564 21420
rect 19180 21028 19236 21532
rect 19292 21586 19348 21598
rect 19292 21534 19294 21586
rect 19346 21534 19348 21586
rect 19292 21364 19348 21534
rect 19292 21298 19348 21308
rect 19516 21586 19572 21598
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19404 21028 19460 21038
rect 19180 21026 19460 21028
rect 19180 20974 19406 21026
rect 19458 20974 19460 21026
rect 19180 20972 19460 20974
rect 19404 20962 19460 20972
rect 19404 20692 19460 20702
rect 16156 20066 16212 20076
rect 17724 20132 17780 20142
rect 18508 20132 18676 20188
rect 15372 19954 15428 19964
rect 14812 18676 14868 18686
rect 14700 18674 15092 18676
rect 14700 18622 14814 18674
rect 14866 18622 15092 18674
rect 14700 18620 15092 18622
rect 14812 18610 14868 18620
rect 14588 17378 14644 17388
rect 15036 17108 15092 18620
rect 15148 18674 15204 19180
rect 15484 19236 15540 19246
rect 15484 19234 16100 19236
rect 15484 19182 15486 19234
rect 15538 19182 16100 19234
rect 15484 19180 16100 19182
rect 15484 19170 15540 19180
rect 15148 18622 15150 18674
rect 15202 18622 15204 18674
rect 15148 18610 15204 18622
rect 16044 18674 16100 19180
rect 17724 19122 17780 20076
rect 17724 19070 17726 19122
rect 17778 19070 17780 19122
rect 16044 18622 16046 18674
rect 16098 18622 16100 18674
rect 16044 18610 16100 18622
rect 16156 19012 16212 19022
rect 16156 18450 16212 18956
rect 16156 18398 16158 18450
rect 16210 18398 16212 18450
rect 16156 18386 16212 18398
rect 17724 18452 17780 19070
rect 18508 19124 18564 19134
rect 18508 19030 18564 19068
rect 17844 18844 18108 18854
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 17844 18778 18108 18788
rect 17948 18452 18004 18462
rect 17724 18450 18004 18452
rect 17724 18398 17950 18450
rect 18002 18398 18004 18450
rect 17724 18396 18004 18398
rect 17948 18386 18004 18396
rect 18396 18450 18452 18462
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 16156 17444 16212 17454
rect 16212 17388 16324 17444
rect 16156 17378 16212 17388
rect 15260 17108 15316 17118
rect 14700 17106 15316 17108
rect 14700 17054 15262 17106
rect 15314 17054 15316 17106
rect 14700 17052 15316 17054
rect 13686 16492 13950 16502
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13686 16426 13950 16436
rect 13580 15876 13636 15886
rect 13580 15314 13636 15820
rect 13580 15262 13582 15314
rect 13634 15262 13636 15314
rect 13580 15250 13636 15262
rect 14028 15314 14084 15326
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 15204 14084 15262
rect 14028 15138 14084 15148
rect 13356 15092 13412 15102
rect 13356 13746 13412 15036
rect 13686 14924 13950 14934
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13686 14858 13950 14868
rect 13356 13694 13358 13746
rect 13410 13694 13412 13746
rect 13356 13682 13412 13694
rect 13916 13748 13972 13758
rect 13916 13746 14084 13748
rect 13916 13694 13918 13746
rect 13970 13694 14084 13746
rect 13916 13692 14084 13694
rect 13916 13682 13972 13692
rect 13686 13356 13950 13366
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13686 13290 13950 13300
rect 13468 13188 13524 13198
rect 13468 12850 13524 13132
rect 14028 13076 14084 13692
rect 14588 13076 14644 13086
rect 14028 13074 14644 13076
rect 14028 13022 14590 13074
rect 14642 13022 14644 13074
rect 14028 13020 14644 13022
rect 14588 13010 14644 13020
rect 13468 12798 13470 12850
rect 13522 12798 13524 12850
rect 12908 12738 12964 12750
rect 12908 12686 12910 12738
rect 12962 12686 12964 12738
rect 12908 11732 12964 12686
rect 13468 12068 13524 12798
rect 13804 12850 13860 12862
rect 13804 12798 13806 12850
rect 13858 12798 13860 12850
rect 13804 12740 13860 12798
rect 14476 12852 14532 12862
rect 14476 12850 14644 12852
rect 14476 12798 14478 12850
rect 14530 12798 14644 12850
rect 14476 12796 14644 12798
rect 14476 12786 14532 12796
rect 13916 12740 13972 12750
rect 13804 12684 13916 12740
rect 13916 12674 13972 12684
rect 14588 12402 14644 12796
rect 14588 12350 14590 12402
rect 14642 12350 14644 12402
rect 14588 12338 14644 12350
rect 14700 12740 14756 17052
rect 15260 17042 15316 17052
rect 15596 16994 15652 17006
rect 15596 16942 15598 16994
rect 15650 16942 15652 16994
rect 15596 16884 15652 16942
rect 15596 16818 15652 16828
rect 16044 16882 16100 16894
rect 16044 16830 16046 16882
rect 16098 16830 16100 16882
rect 16044 16772 16100 16830
rect 16044 16706 16100 16716
rect 15932 16660 15988 16670
rect 15484 16658 15988 16660
rect 15484 16606 15934 16658
rect 15986 16606 15988 16658
rect 15484 16604 15988 16606
rect 14812 16098 14868 16110
rect 14812 16046 14814 16098
rect 14866 16046 14868 16098
rect 14812 15204 14868 16046
rect 14812 15138 14868 15148
rect 14924 16100 14980 16110
rect 14924 15148 14980 16044
rect 15484 16098 15540 16604
rect 15932 16594 15988 16604
rect 15484 16046 15486 16098
rect 15538 16046 15540 16098
rect 15484 16034 15540 16046
rect 15596 15426 15652 15438
rect 15596 15374 15598 15426
rect 15650 15374 15652 15426
rect 15596 15204 15652 15374
rect 15932 15428 15988 15438
rect 16268 15428 16324 17388
rect 17844 17276 18108 17286
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 17844 17210 18108 17220
rect 15932 15426 16324 15428
rect 15932 15374 15934 15426
rect 15986 15374 16270 15426
rect 16322 15374 16324 15426
rect 15932 15372 16324 15374
rect 15932 15362 15988 15372
rect 16268 15362 16324 15372
rect 17724 15874 17780 15886
rect 17724 15822 17726 15874
rect 17778 15822 17780 15874
rect 16492 15314 16548 15326
rect 16492 15262 16494 15314
rect 16546 15262 16548 15314
rect 15652 15148 15876 15204
rect 14924 15092 15092 15148
rect 15596 15138 15652 15148
rect 14924 13076 14980 13086
rect 14924 12962 14980 13020
rect 14924 12910 14926 12962
rect 14978 12910 14980 12962
rect 14924 12898 14980 12910
rect 15036 12964 15092 15092
rect 15820 14530 15876 15148
rect 15820 14478 15822 14530
rect 15874 14478 15876 14530
rect 15820 14466 15876 14478
rect 16156 15092 16212 15102
rect 16156 13970 16212 15036
rect 16156 13918 16158 13970
rect 16210 13918 16212 13970
rect 16156 13906 16212 13918
rect 16380 14530 16436 14542
rect 16380 14478 16382 14530
rect 16434 14478 16436 14530
rect 14812 12852 14868 12862
rect 14812 12758 14868 12796
rect 14476 12180 14532 12190
rect 13468 12002 13524 12012
rect 14140 12178 14532 12180
rect 14140 12126 14478 12178
rect 14530 12126 14532 12178
rect 14140 12124 14532 12126
rect 13686 11788 13950 11798
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13686 11722 13950 11732
rect 12908 10724 12964 11676
rect 12908 10658 12964 10668
rect 12796 10610 12852 10622
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12796 9828 12852 10558
rect 13686 10220 13950 10230
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13686 10154 13950 10164
rect 14140 9938 14196 12124
rect 14476 12114 14532 12124
rect 14700 12178 14756 12684
rect 14700 12126 14702 12178
rect 14754 12126 14756 12178
rect 14700 12114 14756 12126
rect 14252 11956 14308 11966
rect 14252 10498 14308 11900
rect 14924 11954 14980 11966
rect 14924 11902 14926 11954
rect 14978 11902 14980 11954
rect 14476 11844 14532 11854
rect 14364 11284 14420 11294
rect 14364 10612 14420 11228
rect 14476 10948 14532 11788
rect 14924 11844 14980 11902
rect 15036 11956 15092 12908
rect 15036 11890 15092 11900
rect 15596 13524 15652 13534
rect 14924 11778 14980 11788
rect 15148 11396 15204 11406
rect 14924 11394 15204 11396
rect 14924 11342 15150 11394
rect 15202 11342 15204 11394
rect 14924 11340 15204 11342
rect 14588 11284 14644 11294
rect 14588 11190 14644 11228
rect 14812 11284 14868 11294
rect 14812 11190 14868 11228
rect 14700 11172 14756 11182
rect 14700 11078 14756 11116
rect 14476 10892 14644 10948
rect 14364 10546 14420 10556
rect 14252 10446 14254 10498
rect 14306 10446 14308 10498
rect 14252 10388 14308 10446
rect 14252 10332 14420 10388
rect 14140 9886 14142 9938
rect 14194 9886 14196 9938
rect 14140 9874 14196 9886
rect 12796 9762 12852 9772
rect 14252 9716 14308 9726
rect 14252 9622 14308 9660
rect 12348 8428 12740 8484
rect 12796 9602 12852 9614
rect 12796 9550 12798 9602
rect 12850 9550 12852 9602
rect 12796 8932 12852 9550
rect 14028 9604 14084 9614
rect 14028 9510 14084 9548
rect 14364 9044 14420 10332
rect 14364 8978 14420 8988
rect 12124 7700 12180 7710
rect 12124 7606 12180 7644
rect 12012 7588 12068 7598
rect 12012 7494 12068 7532
rect 12236 6132 12292 6142
rect 12124 6076 12236 6132
rect 12124 6018 12180 6076
rect 12236 6066 12292 6076
rect 12124 5966 12126 6018
rect 12178 5966 12180 6018
rect 12124 5954 12180 5966
rect 11564 5854 11566 5906
rect 11618 5854 11620 5906
rect 11564 5012 11620 5854
rect 11788 5908 11844 5918
rect 11788 5796 11844 5852
rect 12012 5796 12068 5806
rect 11788 5794 12068 5796
rect 11788 5742 12014 5794
rect 12066 5742 12068 5794
rect 11788 5740 12068 5742
rect 11676 5348 11732 5358
rect 11788 5348 11844 5740
rect 12012 5730 12068 5740
rect 12348 5572 12404 8428
rect 12460 8148 12516 8158
rect 12460 8054 12516 8092
rect 12796 8148 12852 8876
rect 13686 8652 13950 8662
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13686 8586 13950 8596
rect 14028 8372 14084 8382
rect 14028 8278 14084 8316
rect 13468 8260 13524 8270
rect 12796 8054 12852 8092
rect 13020 8258 13524 8260
rect 13020 8206 13470 8258
rect 13522 8206 13524 8258
rect 13020 8204 13524 8206
rect 12908 8036 12964 8046
rect 12908 7942 12964 7980
rect 13020 7700 13076 8204
rect 13468 8194 13524 8204
rect 13804 8260 13860 8270
rect 13020 7606 13076 7644
rect 12908 7588 12964 7598
rect 12908 7474 12964 7532
rect 13804 7588 13860 8204
rect 14476 8260 14532 8270
rect 14476 8166 14532 8204
rect 14588 8148 14644 10892
rect 14812 10836 14868 10846
rect 14924 10836 14980 11340
rect 15148 11330 15204 11340
rect 14700 10834 14980 10836
rect 14700 10782 14814 10834
rect 14866 10782 14980 10834
rect 14700 10780 14980 10782
rect 15484 10836 15540 10846
rect 14700 10050 14756 10780
rect 14812 10770 14868 10780
rect 15484 10742 15540 10780
rect 15372 10724 15428 10734
rect 15372 10164 15428 10668
rect 14700 9998 14702 10050
rect 14754 9998 14756 10050
rect 14700 9986 14756 9998
rect 14812 10052 14868 10062
rect 14812 9826 14868 9996
rect 14812 9774 14814 9826
rect 14866 9774 14868 9826
rect 14812 8258 14868 9774
rect 14924 9828 14980 9838
rect 14924 9734 14980 9772
rect 15260 9044 15316 9054
rect 15260 8950 15316 8988
rect 14812 8206 14814 8258
rect 14866 8206 14868 8258
rect 14812 8194 14868 8206
rect 15372 8260 15428 10108
rect 15596 9828 15652 13468
rect 15708 13076 15764 13086
rect 15708 11394 15764 13020
rect 16268 13076 16324 13086
rect 16380 13076 16436 14478
rect 16492 13524 16548 15262
rect 17724 15316 17780 15822
rect 17844 15708 18108 15718
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 17844 15642 18108 15652
rect 18396 15540 18452 18398
rect 18620 17108 18676 20132
rect 19404 20130 19460 20636
rect 19404 20078 19406 20130
rect 19458 20078 19460 20130
rect 19404 20066 19460 20078
rect 19068 20018 19124 20030
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 19068 19572 19124 19966
rect 18508 17052 18676 17108
rect 18844 19516 19124 19572
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 18844 19010 18900 19516
rect 19180 19236 19236 19246
rect 19180 19142 19236 19180
rect 18844 18958 18846 19010
rect 18898 18958 18900 19010
rect 18508 16100 18564 17052
rect 18844 16996 18900 18958
rect 18956 19124 19012 19134
rect 19292 19124 19348 19966
rect 19516 20018 19572 21534
rect 19740 21588 19796 21598
rect 19964 21588 20020 21598
rect 19740 21586 19908 21588
rect 19740 21534 19742 21586
rect 19794 21534 19908 21586
rect 19740 21532 19908 21534
rect 19740 21522 19796 21532
rect 19628 21476 19684 21486
rect 19628 21382 19684 21420
rect 19852 20916 19908 21532
rect 19964 21586 20132 21588
rect 19964 21534 19966 21586
rect 20018 21534 20132 21586
rect 19964 21532 20132 21534
rect 19964 21522 20020 21532
rect 19964 20916 20020 20926
rect 19852 20914 20020 20916
rect 19852 20862 19966 20914
rect 20018 20862 20020 20914
rect 19852 20860 20020 20862
rect 19740 20804 19796 20814
rect 19740 20710 19796 20748
rect 19852 20244 19908 20860
rect 19964 20850 20020 20860
rect 19740 20132 19908 20188
rect 19740 20130 19796 20132
rect 19740 20078 19742 20130
rect 19794 20078 19796 20130
rect 19740 20066 19796 20078
rect 19516 19966 19518 20018
rect 19570 19966 19572 20018
rect 19516 19236 19572 19966
rect 19516 19170 19572 19180
rect 20076 20020 20132 21532
rect 20972 21586 21028 21598
rect 20972 21534 20974 21586
rect 21026 21534 21028 21586
rect 20524 21476 20580 21486
rect 20524 21382 20580 21420
rect 20300 20692 20356 20702
rect 20300 20598 20356 20636
rect 20412 20578 20468 20590
rect 20412 20526 20414 20578
rect 20466 20526 20468 20578
rect 20412 20188 20468 20526
rect 20412 20132 20804 20188
rect 20076 19234 20132 19964
rect 20412 20020 20468 20030
rect 20412 20018 20692 20020
rect 20412 19966 20414 20018
rect 20466 19966 20692 20018
rect 20412 19964 20692 19966
rect 20412 19954 20468 19964
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 19404 19124 19460 19134
rect 19292 19068 19404 19124
rect 18956 19010 19012 19068
rect 19404 19030 19460 19068
rect 18956 18958 18958 19010
rect 19010 18958 19012 19010
rect 18956 17668 19012 18958
rect 19068 19012 19124 19022
rect 19740 19012 19796 19022
rect 19068 18918 19124 18956
rect 19628 19010 19796 19012
rect 19628 18958 19742 19010
rect 19794 18958 19796 19010
rect 19628 18956 19796 18958
rect 19292 17668 19348 17678
rect 18956 17666 19348 17668
rect 18956 17614 19294 17666
rect 19346 17614 19348 17666
rect 18956 17612 19348 17614
rect 19292 17556 19348 17612
rect 19516 17668 19572 17678
rect 19628 17668 19684 18956
rect 19740 18946 19796 18956
rect 19964 18676 20020 18686
rect 20076 18676 20132 19182
rect 19964 18674 20132 18676
rect 19964 18622 19966 18674
rect 20018 18622 20132 18674
rect 19964 18620 20132 18622
rect 20636 19796 20692 19964
rect 20748 20018 20804 20132
rect 20748 19966 20750 20018
rect 20802 19966 20804 20018
rect 20748 19954 20804 19966
rect 20972 19796 21028 21534
rect 21532 21586 21588 21756
rect 23884 21700 23940 21710
rect 21532 21534 21534 21586
rect 21586 21534 21588 21586
rect 21532 21522 21588 21534
rect 23772 21698 23940 21700
rect 23772 21646 23886 21698
rect 23938 21646 23940 21698
rect 23772 21644 23940 21646
rect 22002 21196 22266 21206
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22002 21130 22266 21140
rect 23100 20804 23156 20814
rect 23100 20710 23156 20748
rect 20636 19740 21028 19796
rect 23100 20242 23156 20254
rect 23100 20190 23102 20242
rect 23154 20190 23156 20242
rect 23100 20188 23156 20190
rect 23772 20188 23828 21644
rect 23884 21634 23940 21644
rect 23100 20132 23828 20188
rect 19964 18610 20020 18620
rect 20300 18452 20356 18462
rect 20524 18452 20580 18462
rect 20300 18450 20524 18452
rect 20300 18398 20302 18450
rect 20354 18398 20524 18450
rect 20300 18396 20524 18398
rect 20300 18386 20356 18396
rect 20524 18386 20580 18396
rect 20076 17668 20132 17678
rect 20188 17668 20244 17678
rect 19628 17612 19796 17668
rect 19516 17574 19572 17612
rect 19292 17490 19348 17500
rect 19404 17442 19460 17454
rect 19404 17390 19406 17442
rect 19458 17390 19460 17442
rect 19404 17220 19460 17390
rect 18844 16930 18900 16940
rect 19068 17164 19460 17220
rect 19628 17442 19684 17454
rect 19628 17390 19630 17442
rect 19682 17390 19684 17442
rect 19628 17332 19684 17390
rect 18620 16884 18676 16894
rect 18620 16790 18676 16828
rect 18732 16882 18788 16894
rect 18732 16830 18734 16882
rect 18786 16830 18788 16882
rect 18508 16044 18676 16100
rect 18508 15876 18564 15886
rect 18508 15782 18564 15820
rect 18396 15474 18452 15484
rect 17724 15250 17780 15260
rect 18620 14308 18676 16044
rect 18732 15876 18788 16830
rect 18956 16884 19012 16894
rect 19068 16884 19124 17164
rect 19180 16996 19236 17006
rect 19628 16996 19684 17276
rect 19180 16994 19684 16996
rect 19180 16942 19182 16994
rect 19234 16942 19684 16994
rect 19180 16940 19684 16942
rect 19740 17442 19796 17612
rect 20132 17666 20244 17668
rect 20132 17614 20190 17666
rect 20242 17614 20244 17666
rect 20132 17612 20244 17614
rect 20076 17602 20132 17612
rect 20188 17602 20244 17612
rect 19740 17390 19742 17442
rect 19794 17390 19796 17442
rect 19180 16930 19236 16940
rect 18956 16882 19124 16884
rect 18956 16830 18958 16882
rect 19010 16830 19124 16882
rect 18956 16828 19124 16830
rect 19740 16884 19796 17390
rect 20300 17442 20356 17454
rect 20300 17390 20302 17442
rect 20354 17390 20356 17442
rect 20300 17108 20356 17390
rect 20300 17052 20580 17108
rect 18844 16772 18900 16782
rect 18844 16678 18900 16716
rect 18956 16660 19012 16828
rect 19740 16818 19796 16828
rect 20076 16884 20132 16894
rect 20076 16790 20132 16828
rect 20524 16882 20580 17052
rect 20524 16830 20526 16882
rect 20578 16830 20580 16882
rect 20524 16818 20580 16830
rect 20636 16884 20692 19740
rect 22002 19628 22266 19638
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22002 19562 22266 19572
rect 20860 19460 20916 19470
rect 20636 16818 20692 16828
rect 20748 19404 20860 19460
rect 18956 16594 19012 16604
rect 20412 15876 20468 15886
rect 18732 15810 18788 15820
rect 20188 15874 20468 15876
rect 20188 15822 20414 15874
rect 20466 15822 20468 15874
rect 20188 15820 20468 15822
rect 19404 15540 19460 15550
rect 18732 15316 18788 15326
rect 18732 15204 18788 15260
rect 19404 15314 19460 15484
rect 19852 15540 19908 15550
rect 19852 15446 19908 15484
rect 20076 15316 20132 15326
rect 20188 15316 20244 15820
rect 20412 15810 20468 15820
rect 20636 15540 20692 15550
rect 20748 15540 20804 19404
rect 20860 19394 20916 19404
rect 20636 15538 20804 15540
rect 20636 15486 20638 15538
rect 20690 15486 20804 15538
rect 20636 15484 20804 15486
rect 20860 18452 20916 18462
rect 20860 16100 20916 18396
rect 22002 18060 22266 18070
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22002 17994 22266 18004
rect 23100 17106 23156 20132
rect 24220 19908 24276 19918
rect 24556 19908 24612 22318
rect 24780 22148 24836 22158
rect 24668 21364 24724 21374
rect 24668 20244 24724 21308
rect 24668 20178 24724 20188
rect 24220 19906 24612 19908
rect 24220 19854 24222 19906
rect 24274 19854 24612 19906
rect 24220 19852 24612 19854
rect 23884 19796 23940 19806
rect 23884 19124 23940 19740
rect 23996 19460 24052 19470
rect 23996 19346 24052 19404
rect 23996 19294 23998 19346
rect 24050 19294 24052 19346
rect 23996 19282 24052 19294
rect 23884 19058 23940 19068
rect 23996 18340 24052 18350
rect 24220 18340 24276 19852
rect 24444 19348 24500 19358
rect 24780 19348 24836 22092
rect 25116 20914 25172 23100
rect 25564 22596 25620 22606
rect 25564 22502 25620 22540
rect 26908 22596 26964 25200
rect 30492 22932 30548 25200
rect 31612 24724 31668 24734
rect 30492 22876 30772 22932
rect 30318 22764 30582 22774
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30318 22698 30582 22708
rect 26908 22530 26964 22540
rect 28588 22596 28644 22606
rect 28588 22502 28644 22540
rect 27804 22370 27860 22382
rect 27804 22318 27806 22370
rect 27858 22318 27860 22370
rect 26572 22260 26628 22270
rect 26160 21980 26424 21990
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26160 21914 26424 21924
rect 26572 21810 26628 22204
rect 27468 22260 27524 22270
rect 27468 22166 27524 22204
rect 26572 21758 26574 21810
rect 26626 21758 26628 21810
rect 26572 21746 26628 21758
rect 27580 22146 27636 22158
rect 27580 22094 27582 22146
rect 27634 22094 27636 22146
rect 25116 20862 25118 20914
rect 25170 20862 25172 20914
rect 25116 20850 25172 20862
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 20692 25284 21534
rect 25452 21586 25508 21598
rect 25452 21534 25454 21586
rect 25506 21534 25508 21586
rect 25452 21364 25508 21534
rect 25900 21588 25956 21598
rect 25676 21476 25732 21486
rect 25676 21382 25732 21420
rect 25452 21298 25508 21308
rect 25228 20626 25284 20636
rect 25564 20804 25620 20814
rect 25564 20018 25620 20748
rect 25900 20692 25956 21532
rect 26124 21586 26180 21598
rect 26124 21534 26126 21586
rect 26178 21534 26180 21586
rect 26124 20804 26180 21534
rect 26124 20738 26180 20748
rect 26348 21586 26404 21598
rect 26348 21534 26350 21586
rect 26402 21534 26404 21586
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25564 19954 25620 19966
rect 25676 20636 25956 20692
rect 25228 19796 25284 19806
rect 24444 19346 24836 19348
rect 24444 19294 24446 19346
rect 24498 19294 24836 19346
rect 24444 19292 24836 19294
rect 24892 19794 25284 19796
rect 24892 19742 25230 19794
rect 25282 19742 25284 19794
rect 24892 19740 25284 19742
rect 24444 19282 24500 19292
rect 24444 18452 24500 18462
rect 24444 18358 24500 18396
rect 23996 18338 24276 18340
rect 23996 18286 23998 18338
rect 24050 18286 24276 18338
rect 23996 18284 24276 18286
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 22988 16884 23044 16894
rect 22002 16492 22266 16502
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22002 16426 22266 16436
rect 22204 16324 22260 16334
rect 20636 15428 20692 15484
rect 20636 15362 20692 15372
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19404 15250 19460 15262
rect 19964 15314 20244 15316
rect 19964 15262 20078 15314
rect 20130 15262 20244 15314
rect 19964 15260 20244 15262
rect 20524 15314 20580 15326
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 18956 15204 19012 15214
rect 18732 15202 19012 15204
rect 18732 15150 18958 15202
rect 19010 15150 19012 15202
rect 18732 15148 19012 15150
rect 18732 14418 18788 15148
rect 18956 15138 19012 15148
rect 18732 14366 18734 14418
rect 18786 14366 18788 14418
rect 18732 14354 18788 14366
rect 19516 14308 19572 14318
rect 18508 14252 18676 14308
rect 19404 14306 19572 14308
rect 19404 14254 19518 14306
rect 19570 14254 19572 14306
rect 19404 14252 19572 14254
rect 17844 14140 18108 14150
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 17844 14074 18108 14084
rect 16492 13458 16548 13468
rect 16940 13524 16996 13534
rect 16940 13430 16996 13468
rect 16268 13074 16436 13076
rect 16268 13022 16270 13074
rect 16322 13022 16436 13074
rect 16268 13020 16436 13022
rect 16268 13010 16324 13020
rect 15820 12964 15876 12974
rect 15820 12870 15876 12908
rect 16044 12852 16100 12862
rect 16380 12852 16436 12862
rect 16044 12758 16100 12796
rect 16156 12850 16436 12852
rect 16156 12798 16382 12850
rect 16434 12798 16436 12850
rect 16156 12796 16436 12798
rect 16156 12402 16212 12796
rect 16380 12786 16436 12796
rect 16604 12852 16660 12862
rect 16156 12350 16158 12402
rect 16210 12350 16212 12402
rect 16156 12338 16212 12350
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 15708 11330 15764 11342
rect 16044 12290 16100 12302
rect 16044 12238 16046 12290
rect 16098 12238 16100 12290
rect 16044 11284 16100 12238
rect 16268 11956 16324 11966
rect 16268 11954 16548 11956
rect 16268 11902 16270 11954
rect 16322 11902 16548 11954
rect 16268 11900 16548 11902
rect 16268 11890 16324 11900
rect 15820 11172 15876 11182
rect 15820 10610 15876 11116
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15820 10546 15876 10558
rect 16044 10500 16100 11228
rect 16380 10724 16436 10734
rect 16380 10630 16436 10668
rect 16044 10434 16100 10444
rect 16492 9940 16548 11900
rect 16604 11172 16660 12796
rect 17844 12572 18108 12582
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 17844 12506 18108 12516
rect 17388 12292 17444 12302
rect 16604 10610 16660 11116
rect 16604 10558 16606 10610
rect 16658 10558 16660 10610
rect 16604 10546 16660 10558
rect 17276 11394 17332 11406
rect 17276 11342 17278 11394
rect 17330 11342 17332 11394
rect 15820 9938 16548 9940
rect 15820 9886 16494 9938
rect 16546 9886 16548 9938
rect 15820 9884 16548 9886
rect 15596 9772 15764 9828
rect 15372 8194 15428 8204
rect 15596 9604 15652 9614
rect 15596 8932 15652 9548
rect 14700 8148 14756 8158
rect 14588 8146 14756 8148
rect 14588 8094 14702 8146
rect 14754 8094 14756 8146
rect 14588 8092 14756 8094
rect 14700 8082 14756 8092
rect 15596 8146 15652 8876
rect 15708 8428 15764 9772
rect 15820 9042 15876 9884
rect 16492 9874 16548 9884
rect 16604 9826 16660 9838
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 15820 8990 15822 9042
rect 15874 8990 15876 9042
rect 15820 8978 15876 8990
rect 16268 9716 16324 9726
rect 16268 9044 16324 9660
rect 16604 9268 16660 9774
rect 16604 9202 16660 9212
rect 16716 9716 16772 9726
rect 16716 9154 16772 9660
rect 16716 9102 16718 9154
rect 16770 9102 16772 9154
rect 16716 9090 16772 9102
rect 17276 9604 17332 11342
rect 17388 10276 17444 12236
rect 17612 11172 17668 11182
rect 17612 11078 17668 11116
rect 17844 11004 18108 11014
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 17844 10938 18108 10948
rect 18172 10724 18228 10734
rect 18060 10612 18116 10622
rect 18060 10518 18116 10556
rect 17388 10050 17444 10220
rect 18172 10388 18228 10668
rect 18396 10500 18452 10510
rect 18396 10406 18452 10444
rect 17388 9998 17390 10050
rect 17442 9998 17444 10050
rect 17388 9986 17444 9998
rect 17724 10052 17780 10062
rect 17724 9958 17780 9996
rect 17948 9716 18004 9726
rect 17948 9604 18004 9660
rect 16492 9044 16548 9054
rect 16268 8988 16492 9044
rect 16492 8950 16548 8988
rect 16604 8930 16660 8942
rect 16604 8878 16606 8930
rect 16658 8878 16660 8930
rect 15708 8372 16548 8428
rect 15596 8094 15598 8146
rect 15650 8094 15652 8146
rect 15596 8082 15652 8094
rect 13916 8036 13972 8046
rect 13916 7942 13972 7980
rect 14140 8034 14196 8046
rect 14140 7982 14142 8034
rect 14194 7982 14196 8034
rect 13860 7532 14084 7588
rect 13804 7522 13860 7532
rect 12908 7422 12910 7474
rect 12962 7422 12964 7474
rect 12908 7410 12964 7422
rect 13244 7476 13300 7486
rect 13300 7420 13524 7476
rect 13244 7382 13300 7420
rect 13132 7364 13188 7374
rect 13132 7270 13188 7308
rect 12572 7252 12628 7262
rect 12572 7250 12740 7252
rect 12572 7198 12574 7250
rect 12626 7198 12740 7250
rect 12572 7196 12740 7198
rect 12572 7186 12628 7196
rect 12572 6916 12628 6926
rect 12572 5906 12628 6860
rect 12684 6132 12740 7196
rect 13468 6916 13524 7420
rect 13686 7084 13950 7094
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13686 7018 13950 7028
rect 13524 6860 13748 6916
rect 13468 6822 13524 6860
rect 12796 6132 12852 6142
rect 12740 6130 12852 6132
rect 12740 6078 12798 6130
rect 12850 6078 12852 6130
rect 12740 6076 12852 6078
rect 12684 6038 12740 6076
rect 12796 6066 12852 6076
rect 13692 6130 13748 6860
rect 13692 6078 13694 6130
rect 13746 6078 13748 6130
rect 13692 6066 13748 6078
rect 12572 5854 12574 5906
rect 12626 5854 12628 5906
rect 12572 5842 12628 5854
rect 13020 6020 13076 6030
rect 13020 5906 13076 5964
rect 14028 6020 14084 7532
rect 14140 7476 14196 7982
rect 15260 8034 15316 8046
rect 15260 7982 15262 8034
rect 15314 7982 15316 8034
rect 14140 7410 14196 7420
rect 15148 7586 15204 7598
rect 15148 7534 15150 7586
rect 15202 7534 15204 7586
rect 15148 7476 15204 7534
rect 15148 7410 15204 7420
rect 15260 6244 15316 7982
rect 15484 7474 15540 7486
rect 15484 7422 15486 7474
rect 15538 7422 15540 7474
rect 15484 6580 15540 7422
rect 16380 6916 16436 6926
rect 16380 6822 16436 6860
rect 15484 6514 15540 6524
rect 16044 6468 16100 6478
rect 15260 6178 15316 6188
rect 15932 6466 16100 6468
rect 15932 6414 16046 6466
rect 16098 6414 16100 6466
rect 15932 6412 16100 6414
rect 13020 5854 13022 5906
rect 13074 5854 13076 5906
rect 13020 5842 13076 5854
rect 13244 5908 13300 5918
rect 13916 5908 13972 5918
rect 13300 5852 13524 5908
rect 13244 5814 13300 5852
rect 12684 5796 12740 5806
rect 12684 5702 12740 5740
rect 12348 5516 12740 5572
rect 11676 5346 11844 5348
rect 11676 5294 11678 5346
rect 11730 5294 11844 5346
rect 11676 5292 11844 5294
rect 11676 5282 11732 5292
rect 11564 4946 11620 4956
rect 11116 4846 11118 4898
rect 11170 4846 11172 4898
rect 11116 4834 11172 4846
rect 10780 4564 10836 4574
rect 10780 4470 10836 4508
rect 10668 4398 10670 4450
rect 10722 4398 10724 4450
rect 10668 4386 10724 4398
rect 11004 4452 11060 4462
rect 11004 4358 11060 4396
rect 12124 4452 12180 4462
rect 12124 4358 12180 4396
rect 10220 4340 10276 4350
rect 10108 4338 10276 4340
rect 10108 4286 10222 4338
rect 10274 4286 10276 4338
rect 10108 4284 10276 4286
rect 10220 4274 10276 4284
rect 11116 4340 11172 4350
rect 11116 4246 11172 4284
rect 11900 4340 11956 4350
rect 11900 4246 11956 4284
rect 9884 4226 10052 4228
rect 9884 4174 9886 4226
rect 9938 4174 10052 4226
rect 9884 4172 10052 4174
rect 11564 4228 11620 4238
rect 9884 4162 9940 4172
rect 11564 4134 11620 4172
rect 8876 3836 9380 3892
rect 8876 3666 8932 3836
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 8876 3602 8932 3614
rect 8988 3668 9044 3678
rect 5964 3556 6020 3566
rect 5852 3554 6020 3556
rect 5852 3502 5966 3554
rect 6018 3502 6020 3554
rect 5852 3500 6020 3502
rect 4620 3490 4676 3500
rect 5964 3490 6020 3500
rect 3388 1810 3444 1820
rect 5404 3444 5460 3454
rect 5404 800 5460 3388
rect 6636 3444 6692 3454
rect 6636 3330 6692 3388
rect 6636 3278 6638 3330
rect 6690 3278 6692 3330
rect 6636 3266 6692 3278
rect 8988 800 9044 3612
rect 9324 3554 9380 3836
rect 10332 3668 10388 3678
rect 10332 3574 10388 3612
rect 12572 3668 12628 3678
rect 9324 3502 9326 3554
rect 9378 3502 9380 3554
rect 9324 3490 9380 3502
rect 9528 3164 9792 3174
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9528 3098 9792 3108
rect 12572 800 12628 3612
rect 12684 3668 12740 5516
rect 13468 5348 13524 5852
rect 13916 5814 13972 5852
rect 14028 5906 14084 5964
rect 14812 6132 14868 6142
rect 14812 6018 14868 6076
rect 14812 5966 14814 6018
rect 14866 5966 14868 6018
rect 14812 5954 14868 5966
rect 15148 6018 15204 6030
rect 15596 6020 15652 6030
rect 15148 5966 15150 6018
rect 15202 5966 15204 6018
rect 14028 5854 14030 5906
rect 14082 5854 14084 5906
rect 14028 5842 14084 5854
rect 13804 5794 13860 5806
rect 13804 5742 13806 5794
rect 13858 5742 13860 5794
rect 13804 5684 13860 5742
rect 14364 5684 14420 5694
rect 14700 5684 14756 5694
rect 13804 5628 14084 5684
rect 13686 5516 13950 5526
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13686 5450 13950 5460
rect 13580 5348 13636 5358
rect 13468 5346 13636 5348
rect 13468 5294 13582 5346
rect 13634 5294 13636 5346
rect 13468 5292 13636 5294
rect 13580 5282 13636 5292
rect 13468 5012 13524 5022
rect 13132 5010 13524 5012
rect 13132 4958 13470 5010
rect 13522 4958 13524 5010
rect 13132 4956 13524 4958
rect 13132 4562 13188 4956
rect 13468 4946 13524 4956
rect 14028 4900 14084 5628
rect 14364 5682 14756 5684
rect 14364 5630 14366 5682
rect 14418 5630 14702 5682
rect 14754 5630 14756 5682
rect 14364 5628 14756 5630
rect 14364 5618 14420 5628
rect 14700 5618 14756 5628
rect 15148 5348 15204 5966
rect 15484 5964 15596 6020
rect 15484 5906 15540 5964
rect 15596 5954 15652 5964
rect 15484 5854 15486 5906
rect 15538 5854 15540 5906
rect 15484 5842 15540 5854
rect 15932 5906 15988 6412
rect 16044 6402 16100 6412
rect 16492 6130 16548 8372
rect 16604 6580 16660 8878
rect 17276 8428 17332 9548
rect 17724 9548 18004 9604
rect 17500 9268 17556 9278
rect 17500 9154 17556 9212
rect 17500 9102 17502 9154
rect 17554 9102 17556 9154
rect 17500 9090 17556 9102
rect 17388 8932 17444 8942
rect 17388 8838 17444 8876
rect 17052 8372 17332 8428
rect 16716 8260 16772 8270
rect 16716 8166 16772 8204
rect 17052 8258 17108 8372
rect 17052 8206 17054 8258
rect 17106 8206 17108 8258
rect 17052 8194 17108 8206
rect 17724 7698 17780 9548
rect 17844 9436 18108 9446
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 17844 9370 18108 9380
rect 18172 8428 18228 10332
rect 18284 9828 18340 9838
rect 18284 9734 18340 9772
rect 18172 8372 18340 8428
rect 18284 8258 18340 8372
rect 18284 8206 18286 8258
rect 18338 8206 18340 8258
rect 18284 8194 18340 8206
rect 17844 7868 18108 7878
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 17844 7802 18108 7812
rect 17724 7646 17726 7698
rect 17778 7646 17780 7698
rect 17724 7634 17780 7646
rect 17388 7588 17444 7598
rect 17388 6916 17444 7532
rect 17388 6850 17444 6860
rect 16604 6486 16660 6524
rect 16940 6578 16996 6590
rect 16940 6526 16942 6578
rect 16994 6526 16996 6578
rect 16492 6078 16494 6130
rect 16546 6078 16548 6130
rect 15932 5854 15934 5906
rect 15986 5854 15988 5906
rect 15932 5842 15988 5854
rect 16156 6018 16212 6030
rect 16156 5966 16158 6018
rect 16210 5966 16212 6018
rect 15148 5282 15204 5292
rect 16044 5348 16100 5358
rect 16044 5122 16100 5292
rect 16044 5070 16046 5122
rect 16098 5070 16100 5122
rect 16044 5058 16100 5070
rect 16156 5124 16212 5966
rect 16492 6020 16548 6078
rect 16940 6468 16996 6526
rect 16940 6132 16996 6412
rect 17844 6300 18108 6310
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 17844 6234 18108 6244
rect 17724 6132 17780 6142
rect 16940 6066 16996 6076
rect 17500 6076 17724 6132
rect 16492 5954 16548 5964
rect 16716 5908 16772 5918
rect 16716 5814 16772 5852
rect 16604 5348 16660 5358
rect 16660 5292 16772 5348
rect 16604 5282 16660 5292
rect 16604 5124 16660 5134
rect 16156 5122 16660 5124
rect 16156 5070 16606 5122
rect 16658 5070 16660 5122
rect 16156 5068 16660 5070
rect 16604 5058 16660 5068
rect 14028 4834 14084 4844
rect 16156 4900 16212 4910
rect 13132 4510 13134 4562
rect 13186 4510 13188 4562
rect 13132 4452 13188 4510
rect 13692 4676 13748 4686
rect 13692 4562 13748 4620
rect 13692 4510 13694 4562
rect 13746 4510 13748 4562
rect 13692 4498 13748 4510
rect 13132 4386 13188 4396
rect 16156 4338 16212 4844
rect 16156 4286 16158 4338
rect 16210 4286 16212 4338
rect 16156 4274 16212 4286
rect 16716 4338 16772 5292
rect 17500 4450 17556 6076
rect 17724 6038 17780 6076
rect 18508 6132 18564 14252
rect 18620 13524 18676 13534
rect 18620 12962 18676 13468
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18620 12898 18676 12910
rect 19404 12964 19460 14252
rect 19516 14242 19572 14252
rect 19852 13858 19908 13870
rect 19852 13806 19854 13858
rect 19906 13806 19908 13858
rect 19516 13746 19572 13758
rect 19516 13694 19518 13746
rect 19570 13694 19572 13746
rect 19516 13524 19572 13694
rect 19516 13458 19572 13468
rect 18732 12740 18788 12750
rect 19068 12740 19124 12750
rect 18732 12738 19068 12740
rect 18732 12686 18734 12738
rect 18786 12686 19068 12738
rect 18732 12684 19068 12686
rect 18732 12674 18788 12684
rect 19068 12646 19124 12684
rect 18956 12180 19012 12218
rect 18956 12114 19012 12124
rect 19404 12178 19460 12908
rect 19404 12126 19406 12178
rect 19458 12126 19460 12178
rect 19404 12114 19460 12126
rect 19628 12850 19684 12862
rect 19628 12798 19630 12850
rect 19682 12798 19684 12850
rect 18620 11954 18676 11966
rect 18620 11902 18622 11954
rect 18674 11902 18676 11954
rect 18620 11620 18676 11902
rect 18620 11282 18676 11564
rect 18620 11230 18622 11282
rect 18674 11230 18676 11282
rect 18620 11218 18676 11230
rect 18956 11954 19012 11966
rect 18956 11902 18958 11954
rect 19010 11902 19012 11954
rect 18844 10610 18900 10622
rect 18844 10558 18846 10610
rect 18898 10558 18900 10610
rect 18844 10276 18900 10558
rect 18956 10612 19012 11902
rect 19180 11394 19236 11406
rect 19180 11342 19182 11394
rect 19234 11342 19236 11394
rect 19180 11284 19236 11342
rect 19628 11396 19684 12798
rect 19740 12740 19796 12750
rect 19740 12292 19796 12684
rect 19852 12628 19908 13806
rect 19852 12562 19908 12572
rect 19964 13636 20020 15260
rect 20076 15222 20132 15260
rect 20524 14642 20580 15262
rect 20860 15314 20916 16044
rect 21420 16100 21476 16110
rect 21420 16006 21476 16044
rect 22204 16100 22260 16268
rect 22540 16212 22596 16222
rect 22540 16210 22932 16212
rect 22540 16158 22542 16210
rect 22594 16158 22932 16210
rect 22540 16156 22932 16158
rect 22540 16146 22596 16156
rect 22204 16098 22372 16100
rect 22204 16046 22206 16098
rect 22258 16046 22372 16098
rect 22204 16044 22372 16046
rect 22204 16034 22260 16044
rect 21980 15988 22036 15998
rect 21980 15894 22036 15932
rect 21644 15876 21700 15886
rect 21644 15782 21700 15820
rect 22316 15540 22372 16044
rect 22428 15874 22484 15886
rect 22428 15822 22430 15874
rect 22482 15822 22484 15874
rect 22428 15652 22484 15822
rect 22540 15876 22596 15886
rect 22596 15820 22820 15876
rect 22540 15782 22596 15820
rect 22428 15596 22708 15652
rect 22316 15484 22596 15540
rect 20860 15262 20862 15314
rect 20914 15262 20916 15314
rect 20860 15250 20916 15262
rect 22428 15204 22484 15214
rect 22002 14924 22266 14934
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22002 14858 22266 14868
rect 20524 14590 20526 14642
rect 20578 14590 20580 14642
rect 20524 14578 20580 14590
rect 22428 14530 22484 15148
rect 22428 14478 22430 14530
rect 22482 14478 22484 14530
rect 22428 14466 22484 14478
rect 22540 14530 22596 15484
rect 22652 15204 22708 15596
rect 22764 15204 22820 15820
rect 22876 15426 22932 16156
rect 22988 16098 23044 16828
rect 23100 16324 23156 17054
rect 23660 17332 23716 17342
rect 23660 17106 23716 17276
rect 23660 17054 23662 17106
rect 23714 17054 23716 17106
rect 23660 16996 23716 17054
rect 23660 16930 23716 16940
rect 23100 16258 23156 16268
rect 22988 16046 22990 16098
rect 23042 16046 23044 16098
rect 22988 15988 23044 16046
rect 23548 16098 23604 16110
rect 23548 16046 23550 16098
rect 23602 16046 23604 16098
rect 22988 15932 23268 15988
rect 22988 15652 23044 15662
rect 22988 15538 23044 15596
rect 22988 15486 22990 15538
rect 23042 15486 23044 15538
rect 22988 15474 23044 15486
rect 23212 15540 23268 15932
rect 23548 15652 23604 16046
rect 23548 15586 23604 15596
rect 23324 15540 23380 15550
rect 23212 15538 23380 15540
rect 23212 15486 23326 15538
rect 23378 15486 23380 15538
rect 23212 15484 23380 15486
rect 23324 15474 23380 15484
rect 22876 15374 22878 15426
rect 22930 15374 22932 15426
rect 22876 15362 22932 15374
rect 23660 15314 23716 15326
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 22764 15148 23044 15204
rect 22652 15138 22708 15148
rect 22540 14478 22542 14530
rect 22594 14478 22596 14530
rect 22540 14466 22596 14478
rect 22876 14642 22932 14654
rect 22876 14590 22878 14642
rect 22930 14590 22932 14642
rect 22876 14532 22932 14590
rect 22876 14466 22932 14476
rect 22988 14530 23044 15148
rect 23660 15092 23716 15262
rect 23660 15026 23716 15036
rect 23996 14980 24052 18284
rect 24108 15204 24164 15214
rect 24108 15202 24276 15204
rect 24108 15150 24110 15202
rect 24162 15150 24276 15202
rect 24108 15148 24276 15150
rect 24108 15138 24164 15148
rect 24220 15092 24276 15148
rect 24220 15026 24276 15036
rect 23996 14924 24164 14980
rect 22988 14478 22990 14530
rect 23042 14478 23044 14530
rect 22988 14466 23044 14478
rect 23548 14532 23604 14542
rect 23548 14438 23604 14476
rect 23996 14530 24052 14542
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 20636 14418 20692 14430
rect 20636 14366 20638 14418
rect 20690 14366 20692 14418
rect 20412 14308 20468 14318
rect 20412 14214 20468 14252
rect 20636 13860 20692 14366
rect 23660 14420 23716 14430
rect 23660 14326 23716 14364
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 22764 14308 22820 14318
rect 22764 14214 22820 14252
rect 23436 14308 23492 14318
rect 21756 13972 21812 13982
rect 21756 13970 21924 13972
rect 21756 13918 21758 13970
rect 21810 13918 21924 13970
rect 21756 13916 21924 13918
rect 21756 13906 21812 13916
rect 20636 13746 20692 13804
rect 21084 13748 21140 13758
rect 20636 13694 20638 13746
rect 20690 13694 20692 13746
rect 20636 13682 20692 13694
rect 20748 13692 21084 13748
rect 19852 12292 19908 12302
rect 19740 12290 19908 12292
rect 19740 12238 19854 12290
rect 19906 12238 19908 12290
rect 19740 12236 19908 12238
rect 19852 12226 19908 12236
rect 19628 11330 19684 11340
rect 19740 12068 19796 12078
rect 19740 11394 19796 12012
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19740 11330 19796 11342
rect 19068 10612 19124 10622
rect 18956 10610 19124 10612
rect 18956 10558 19070 10610
rect 19122 10558 19124 10610
rect 18956 10556 19124 10558
rect 19068 10546 19124 10556
rect 18844 10210 18900 10220
rect 18956 10386 19012 10398
rect 18956 10334 18958 10386
rect 19010 10334 19012 10386
rect 18620 9716 18676 9726
rect 18676 9660 18788 9716
rect 18620 9622 18676 9660
rect 18732 9154 18788 9660
rect 18732 9102 18734 9154
rect 18786 9102 18788 9154
rect 18732 9090 18788 9102
rect 18956 7812 19012 10334
rect 19180 10164 19236 11228
rect 19180 10098 19236 10108
rect 19068 10052 19124 10062
rect 19068 9828 19124 9996
rect 19068 9762 19124 9772
rect 19180 9492 19236 9502
rect 19180 9044 19236 9436
rect 19180 8950 19236 8988
rect 18956 7746 19012 7756
rect 19292 8930 19348 8942
rect 19292 8878 19294 8930
rect 19346 8878 19348 8930
rect 19292 8034 19348 8878
rect 19292 7982 19294 8034
rect 19346 7982 19348 8034
rect 19292 7700 19348 7982
rect 19292 7634 19348 7644
rect 19516 8034 19572 8046
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19516 7924 19572 7982
rect 19516 7588 19572 7868
rect 19516 7522 19572 7532
rect 19628 8034 19684 8046
rect 19628 7982 19630 8034
rect 19682 7982 19684 8034
rect 19404 7474 19460 7486
rect 19404 7422 19406 7474
rect 19458 7422 19460 7474
rect 18956 7362 19012 7374
rect 18956 7310 18958 7362
rect 19010 7310 19012 7362
rect 18956 7028 19012 7310
rect 18956 6962 19012 6972
rect 18508 6066 18564 6076
rect 19180 6466 19236 6478
rect 19180 6414 19182 6466
rect 19234 6414 19236 6466
rect 18172 6020 18228 6030
rect 18172 5926 18228 5964
rect 18620 6020 18676 6030
rect 18620 5906 18676 5964
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5842 18676 5854
rect 18956 5794 19012 5806
rect 18956 5742 18958 5794
rect 19010 5742 19012 5794
rect 18620 5684 18676 5694
rect 18172 5348 18228 5358
rect 17844 4732 18108 4742
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 17844 4666 18108 4676
rect 17500 4398 17502 4450
rect 17554 4398 17556 4450
rect 17500 4386 17556 4398
rect 16716 4286 16718 4338
rect 16770 4286 16772 4338
rect 16716 4274 16772 4286
rect 18172 4338 18228 5292
rect 18620 4562 18676 5628
rect 18956 4900 19012 5742
rect 19180 5348 19236 6414
rect 19404 5794 19460 7422
rect 19516 6916 19572 6926
rect 19628 6916 19684 7982
rect 19740 8036 19796 8046
rect 19740 7028 19796 7980
rect 19740 6962 19796 6972
rect 19516 6914 19684 6916
rect 19516 6862 19518 6914
rect 19570 6862 19684 6914
rect 19516 6860 19684 6862
rect 19516 6850 19572 6860
rect 19516 6468 19572 6478
rect 19516 6132 19572 6412
rect 19964 6132 20020 13580
rect 20524 13634 20580 13646
rect 20524 13582 20526 13634
rect 20578 13582 20580 13634
rect 20524 13188 20580 13582
rect 20524 13122 20580 13132
rect 20748 13074 20804 13692
rect 21084 13654 21140 13692
rect 21756 13748 21812 13758
rect 20748 13022 20750 13074
rect 20802 13022 20804 13074
rect 20748 13010 20804 13022
rect 21532 12964 21588 12974
rect 21420 12962 21588 12964
rect 21420 12910 21534 12962
rect 21586 12910 21588 12962
rect 21420 12908 21588 12910
rect 21308 12852 21364 12862
rect 21084 12850 21364 12852
rect 21084 12798 21310 12850
rect 21362 12798 21364 12850
rect 21084 12796 21364 12798
rect 20188 12738 20244 12750
rect 20188 12686 20190 12738
rect 20242 12686 20244 12738
rect 20188 12628 20244 12686
rect 20188 12068 20244 12572
rect 21084 12180 21140 12796
rect 21308 12786 21364 12796
rect 21084 12086 21140 12124
rect 20188 12002 20244 12012
rect 20412 11844 20468 11854
rect 20076 11508 20132 11518
rect 20076 11414 20132 11452
rect 20412 11282 20468 11788
rect 20412 11230 20414 11282
rect 20466 11230 20468 11282
rect 20412 11218 20468 11230
rect 20524 11396 20580 11406
rect 20300 10612 20356 10622
rect 20188 9828 20244 9838
rect 20188 8818 20244 9772
rect 20300 9714 20356 10556
rect 20524 10500 20580 11340
rect 21420 11396 21476 12908
rect 21532 12898 21588 12908
rect 21420 11330 21476 11340
rect 21532 12740 21588 12750
rect 21532 11844 21588 12684
rect 21756 12180 21812 13692
rect 21868 13076 21924 13916
rect 22204 13860 22260 13870
rect 22260 13804 22484 13860
rect 22204 13766 22260 13804
rect 22002 13356 22266 13366
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22002 13290 22266 13300
rect 21868 13010 21924 13020
rect 22428 13074 22484 13804
rect 23436 13746 23492 14252
rect 23436 13694 23438 13746
rect 23490 13694 23492 13746
rect 23436 13682 23492 13694
rect 23996 13300 24052 14478
rect 23996 13234 24052 13244
rect 22428 13022 22430 13074
rect 22482 13022 22484 13074
rect 22428 13010 22484 13022
rect 22092 12964 22148 12974
rect 22092 12870 22148 12908
rect 23884 12964 23940 12974
rect 22652 12850 22708 12862
rect 22652 12798 22654 12850
rect 22706 12798 22708 12850
rect 22316 12180 22372 12190
rect 21756 12178 22372 12180
rect 21756 12126 22318 12178
rect 22370 12126 22372 12178
rect 21756 12124 22372 12126
rect 22652 12180 22708 12798
rect 23100 12738 23156 12750
rect 23100 12686 23102 12738
rect 23154 12686 23156 12738
rect 23100 12404 23156 12686
rect 23660 12628 23716 12638
rect 23156 12348 23492 12404
rect 23100 12338 23156 12348
rect 22876 12180 22932 12190
rect 22652 12178 22932 12180
rect 22652 12126 22878 12178
rect 22930 12126 22932 12178
rect 22652 12124 22932 12126
rect 21308 11284 21364 11294
rect 21308 11172 21364 11228
rect 21420 11172 21476 11182
rect 21308 11116 21420 11172
rect 21420 11078 21476 11116
rect 21420 10724 21476 10734
rect 21532 10724 21588 11788
rect 21420 10722 21588 10724
rect 21420 10670 21422 10722
rect 21474 10670 21588 10722
rect 21420 10668 21588 10670
rect 21644 12066 21700 12078
rect 21644 12014 21646 12066
rect 21698 12014 21700 12066
rect 21644 11956 21700 12014
rect 22316 12068 22372 12124
rect 22316 12012 22484 12068
rect 21420 10658 21476 10668
rect 21644 10612 21700 11900
rect 22002 11788 22266 11798
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22002 11722 22266 11732
rect 22092 11620 22148 11630
rect 22092 11394 22148 11564
rect 22092 11342 22094 11394
rect 22146 11342 22148 11394
rect 22092 11330 22148 11342
rect 22428 11394 22484 12012
rect 22540 11956 22596 11966
rect 22540 11954 22708 11956
rect 22540 11902 22542 11954
rect 22594 11902 22708 11954
rect 22540 11900 22708 11902
rect 22540 11890 22596 11900
rect 22428 11342 22430 11394
rect 22482 11342 22484 11394
rect 22428 11330 22484 11342
rect 22540 11732 22596 11742
rect 21868 10612 21924 10622
rect 21644 10610 21924 10612
rect 21644 10558 21870 10610
rect 21922 10558 21924 10610
rect 21644 10556 21924 10558
rect 21868 10546 21924 10556
rect 22316 10610 22372 10622
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 20300 9662 20302 9714
rect 20354 9662 20356 9714
rect 20300 9650 20356 9662
rect 20412 10444 20580 10500
rect 20636 10500 20692 10510
rect 20188 8766 20190 8818
rect 20242 8766 20244 8818
rect 20188 8754 20244 8766
rect 20300 8930 20356 8942
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 20300 8820 20356 8878
rect 20412 8932 20468 10444
rect 20636 10406 20692 10444
rect 22316 10388 22372 10558
rect 22316 10322 22372 10332
rect 22002 10220 22266 10230
rect 21308 10164 21364 10174
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22002 10154 22266 10164
rect 22540 10164 22596 11676
rect 20748 9828 20804 9838
rect 20748 9734 20804 9772
rect 20524 9602 20580 9614
rect 20524 9550 20526 9602
rect 20578 9550 20580 9602
rect 20524 9268 20580 9550
rect 20524 9202 20580 9212
rect 20636 9602 20692 9614
rect 20636 9550 20638 9602
rect 20690 9550 20692 9602
rect 20524 9044 20580 9054
rect 20636 9044 20692 9550
rect 21308 9492 21364 10108
rect 21756 10052 21812 10062
rect 21756 9938 21812 9996
rect 21756 9886 21758 9938
rect 21810 9886 21812 9938
rect 21756 9604 21812 9886
rect 22540 9826 22596 10108
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 22540 9762 22596 9774
rect 21756 9538 21812 9548
rect 21308 9436 21476 9492
rect 21084 9044 21140 9054
rect 20636 9042 21140 9044
rect 20636 8990 21086 9042
rect 21138 8990 21140 9042
rect 20636 8988 21140 8990
rect 20524 8950 20580 8988
rect 21084 8978 21140 8988
rect 20412 8866 20468 8876
rect 20300 8754 20356 8764
rect 21196 8820 21252 8830
rect 20300 8260 20356 8270
rect 20300 8166 20356 8204
rect 20076 8148 20132 8158
rect 20076 6690 20132 8092
rect 20636 8036 20692 8046
rect 20636 7942 20692 7980
rect 21196 7586 21252 8764
rect 21308 8818 21364 8830
rect 21308 8766 21310 8818
rect 21362 8766 21364 8818
rect 21308 8148 21364 8766
rect 21308 8082 21364 8092
rect 21308 7700 21364 7710
rect 21420 7700 21476 9436
rect 22540 8930 22596 8942
rect 22540 8878 22542 8930
rect 22594 8878 22596 8930
rect 22540 8708 22596 8878
rect 22652 8818 22708 11900
rect 22876 11732 22932 12124
rect 23436 12178 23492 12348
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23436 12114 23492 12126
rect 23660 12290 23716 12572
rect 23884 12404 23940 12908
rect 23996 12738 24052 12750
rect 23996 12686 23998 12738
rect 24050 12686 24052 12738
rect 23996 12628 24052 12686
rect 23996 12562 24052 12572
rect 23996 12404 24052 12414
rect 23884 12402 24052 12404
rect 23884 12350 23998 12402
rect 24050 12350 24052 12402
rect 23884 12348 24052 12350
rect 23996 12338 24052 12348
rect 23660 12238 23662 12290
rect 23714 12238 23716 12290
rect 22876 11666 22932 11676
rect 22876 11506 22932 11518
rect 22876 11454 22878 11506
rect 22930 11454 22932 11506
rect 22876 10722 22932 11454
rect 23100 11396 23156 11406
rect 22988 11284 23044 11294
rect 22988 11190 23044 11228
rect 22876 10670 22878 10722
rect 22930 10670 22932 10722
rect 22876 10658 22932 10670
rect 23100 10724 23156 11340
rect 23548 11394 23604 11406
rect 23548 11342 23550 11394
rect 23602 11342 23604 11394
rect 22876 10164 22932 10174
rect 22932 10108 23044 10164
rect 22876 10098 22932 10108
rect 22988 9826 23044 10108
rect 22988 9774 22990 9826
rect 23042 9774 23044 9826
rect 22988 9762 23044 9774
rect 22764 9716 22820 9726
rect 22764 9622 22820 9660
rect 23100 9714 23156 10668
rect 23100 9662 23102 9714
rect 23154 9662 23156 9714
rect 23100 9650 23156 9662
rect 23436 11170 23492 11182
rect 23436 11118 23438 11170
rect 23490 11118 23492 11170
rect 23436 9492 23492 11118
rect 23548 10612 23604 11342
rect 23548 10546 23604 10556
rect 23660 9828 23716 12238
rect 23884 11284 23940 11294
rect 23884 11190 23940 11228
rect 23660 9716 23716 9772
rect 23884 9716 23940 9726
rect 23660 9660 23884 9716
rect 23884 9622 23940 9660
rect 23436 9426 23492 9436
rect 22652 8766 22654 8818
rect 22706 8766 22708 8818
rect 22652 8754 22708 8766
rect 22876 9154 22932 9166
rect 22876 9102 22878 9154
rect 22930 9102 22932 9154
rect 22876 9044 22932 9102
rect 22002 8652 22266 8662
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22540 8642 22596 8652
rect 22002 8586 22266 8596
rect 22876 8428 22932 8988
rect 24108 8428 24164 14924
rect 24444 14530 24500 14542
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 24220 14420 24276 14430
rect 24444 14420 24500 14478
rect 24276 14364 24500 14420
rect 24220 14354 24276 14364
rect 24556 14308 24612 19292
rect 24892 19234 24948 19740
rect 25228 19730 25284 19740
rect 24892 19182 24894 19234
rect 24946 19182 24948 19234
rect 24892 19170 24948 19182
rect 25340 19460 25396 19470
rect 25340 19234 25396 19404
rect 25340 19182 25342 19234
rect 25394 19182 25396 19234
rect 25340 19170 25396 19182
rect 25676 19122 25732 20636
rect 26348 20580 26404 21534
rect 25788 20524 26404 20580
rect 26796 21588 26852 21598
rect 26796 20692 26852 21532
rect 25788 19906 25844 20524
rect 26160 20412 26424 20422
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26160 20346 26424 20356
rect 26572 20132 26628 20142
rect 26572 20018 26628 20076
rect 26572 19966 26574 20018
rect 26626 19966 26628 20018
rect 26572 19954 26628 19966
rect 25788 19854 25790 19906
rect 25842 19854 25844 19906
rect 25788 19796 25844 19854
rect 25788 19730 25844 19740
rect 25676 19070 25678 19122
rect 25730 19070 25732 19122
rect 25676 19058 25732 19070
rect 26160 18844 26424 18854
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26160 18778 26424 18788
rect 25228 18452 25284 18462
rect 25228 18338 25284 18396
rect 25564 18452 25620 18462
rect 25564 18358 25620 18396
rect 26236 18452 26292 18462
rect 26236 18358 26292 18396
rect 26460 18450 26516 18462
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 25228 18286 25230 18338
rect 25282 18286 25284 18338
rect 25228 18274 25284 18286
rect 25788 18340 25844 18350
rect 25788 17556 25844 18284
rect 26460 18340 26516 18398
rect 26796 18450 26852 20636
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 18386 26852 18398
rect 27132 21362 27188 21374
rect 27132 21310 27134 21362
rect 27186 21310 27188 21362
rect 27132 21028 27188 21310
rect 27580 21364 27636 22094
rect 27580 21298 27636 21308
rect 27132 18450 27188 20972
rect 27580 20916 27636 20926
rect 27580 20822 27636 20860
rect 27804 20804 27860 22318
rect 27580 19460 27636 19470
rect 27580 19366 27636 19404
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18386 27188 18398
rect 26460 18274 26516 18284
rect 26572 18340 26628 18350
rect 26572 18338 26740 18340
rect 26572 18286 26574 18338
rect 26626 18286 26740 18338
rect 26572 18284 26740 18286
rect 26572 18274 26628 18284
rect 26124 17668 26180 17678
rect 26572 17668 26628 17678
rect 25788 17490 25844 17500
rect 26012 17666 26628 17668
rect 26012 17614 26126 17666
rect 26178 17614 26574 17666
rect 26626 17614 26628 17666
rect 26012 17612 26628 17614
rect 25900 17442 25956 17454
rect 25900 17390 25902 17442
rect 25954 17390 25956 17442
rect 25900 17332 25956 17390
rect 25900 17266 25956 17276
rect 25452 17108 25508 17118
rect 26012 17108 26068 17612
rect 26124 17602 26180 17612
rect 26572 17602 26628 17612
rect 26160 17276 26424 17286
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26160 17210 26424 17220
rect 25452 17106 26068 17108
rect 25452 17054 25454 17106
rect 25506 17054 26068 17106
rect 25452 17052 26068 17054
rect 25452 17042 25508 17052
rect 24444 14252 24612 14308
rect 25228 16882 25284 16894
rect 25228 16830 25230 16882
rect 25282 16830 25284 16882
rect 24332 10386 24388 10398
rect 24332 10334 24334 10386
rect 24386 10334 24388 10386
rect 24332 10164 24388 10334
rect 24332 10098 24388 10108
rect 24332 8932 24388 8942
rect 24332 8838 24388 8876
rect 24220 8818 24276 8830
rect 24220 8766 24222 8818
rect 24274 8766 24276 8818
rect 24220 8708 24276 8766
rect 24220 8642 24276 8652
rect 22876 8372 23604 8428
rect 21308 7698 21476 7700
rect 21308 7646 21310 7698
rect 21362 7646 21476 7698
rect 21308 7644 21476 7646
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 21308 7634 21364 7644
rect 21196 7534 21198 7586
rect 21250 7534 21252 7586
rect 21196 7522 21252 7534
rect 21532 7476 21588 7486
rect 21532 7382 21588 7420
rect 22092 7252 22148 8206
rect 22652 8258 22708 8270
rect 22652 8206 22654 8258
rect 22706 8206 22708 8258
rect 22540 7700 22596 7710
rect 22652 7700 22708 8206
rect 22540 7698 22708 7700
rect 22540 7646 22542 7698
rect 22594 7646 22708 7698
rect 22540 7644 22708 7646
rect 22540 7634 22596 7644
rect 23324 7586 23380 8372
rect 23548 8306 23604 8316
rect 23996 8372 24164 8428
rect 23324 7534 23326 7586
rect 23378 7534 23380 7586
rect 23324 7522 23380 7534
rect 22204 7476 22260 7486
rect 22652 7476 22708 7486
rect 22876 7476 22932 7486
rect 23212 7476 23268 7486
rect 22260 7420 22596 7476
rect 22204 7382 22260 7420
rect 22092 7186 22148 7196
rect 22428 7252 22484 7262
rect 22002 7084 22266 7094
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22002 7018 22266 7028
rect 20076 6638 20078 6690
rect 20130 6638 20132 6690
rect 20076 6626 20132 6638
rect 20188 6578 20244 6590
rect 20188 6526 20190 6578
rect 20242 6526 20244 6578
rect 20076 6132 20132 6142
rect 19516 6130 19684 6132
rect 19516 6078 19518 6130
rect 19570 6078 19684 6130
rect 19516 6076 19684 6078
rect 19516 6066 19572 6076
rect 19404 5742 19406 5794
rect 19458 5742 19460 5794
rect 19404 5730 19460 5742
rect 19628 5348 19684 6076
rect 19964 6130 20132 6132
rect 19964 6078 20078 6130
rect 20130 6078 20132 6130
rect 19964 6076 20132 6078
rect 19964 6020 20020 6076
rect 20076 6066 20132 6076
rect 19964 5954 20020 5964
rect 19740 5684 19796 5694
rect 19740 5590 19796 5628
rect 20188 5684 20244 6526
rect 20188 5618 20244 5628
rect 20300 5908 20356 5918
rect 19740 5348 19796 5358
rect 19628 5346 19796 5348
rect 19628 5294 19742 5346
rect 19794 5294 19796 5346
rect 19628 5292 19796 5294
rect 19180 5282 19236 5292
rect 19740 5282 19796 5292
rect 18956 4806 19012 4844
rect 20300 5234 20356 5852
rect 20300 5182 20302 5234
rect 20354 5182 20356 5234
rect 18620 4510 18622 4562
rect 18674 4510 18676 4562
rect 18620 4498 18676 4510
rect 19404 4564 19460 4574
rect 19404 4470 19460 4508
rect 18396 4452 18452 4462
rect 20300 4452 20356 5182
rect 20412 5906 20468 5918
rect 20412 5854 20414 5906
rect 20466 5854 20468 5906
rect 20412 5236 20468 5854
rect 22002 5516 22266 5526
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22002 5450 22266 5460
rect 20412 5170 20468 5180
rect 18396 4358 18452 4396
rect 19964 4396 20356 4452
rect 22316 5124 22372 5134
rect 22428 5124 22484 7196
rect 22540 6690 22596 7420
rect 22652 7474 22820 7476
rect 22652 7422 22654 7474
rect 22706 7422 22820 7474
rect 22652 7420 22820 7422
rect 22652 7410 22708 7420
rect 22540 6638 22542 6690
rect 22594 6638 22596 6690
rect 22540 6626 22596 6638
rect 22764 7364 22820 7420
rect 22876 7474 23268 7476
rect 22876 7422 22878 7474
rect 22930 7422 23214 7474
rect 23266 7422 23268 7474
rect 22876 7420 23268 7422
rect 22876 7410 22932 7420
rect 23212 7410 23268 7420
rect 22764 6692 22820 7308
rect 22876 6692 22932 6702
rect 22764 6690 22932 6692
rect 22764 6638 22878 6690
rect 22930 6638 22932 6690
rect 22764 6636 22932 6638
rect 22876 6626 22932 6636
rect 23212 6580 23268 6590
rect 23212 6486 23268 6524
rect 22316 5122 22484 5124
rect 22316 5070 22318 5122
rect 22370 5070 22484 5122
rect 22316 5068 22484 5070
rect 22764 6466 22820 6478
rect 22764 6414 22766 6466
rect 22818 6414 22820 6466
rect 22764 5122 22820 6414
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 18172 4286 18174 4338
rect 18226 4286 18228 4338
rect 18172 4274 18228 4286
rect 17388 4114 17444 4126
rect 17388 4062 17390 4114
rect 17442 4062 17444 4114
rect 13686 3948 13950 3958
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13686 3882 13950 3892
rect 14140 3668 14196 3678
rect 12684 3666 13188 3668
rect 12684 3614 12686 3666
rect 12738 3614 13188 3666
rect 12684 3612 13188 3614
rect 12684 3602 12740 3612
rect 13132 3554 13188 3612
rect 14140 3574 14196 3612
rect 13132 3502 13134 3554
rect 13186 3502 13188 3554
rect 13132 3490 13188 3502
rect 17388 3554 17444 4062
rect 17388 3502 17390 3554
rect 17442 3502 17444 3554
rect 17388 3490 17444 3502
rect 19740 3668 19796 3678
rect 16156 3444 16212 3454
rect 16156 800 16212 3388
rect 18508 3444 18564 3454
rect 18508 3350 18564 3388
rect 17844 3164 18108 3174
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 17844 3098 18108 3108
rect 19740 800 19796 3612
rect 19964 3666 20020 4396
rect 21644 4340 21700 4350
rect 21644 4246 21700 4284
rect 22316 4338 22372 5068
rect 22764 5058 22820 5070
rect 22652 4900 22708 4910
rect 22652 4564 22708 4844
rect 23996 4564 24052 8372
rect 24444 5908 24500 14252
rect 24668 12852 24724 12862
rect 24668 12758 24724 12796
rect 24556 12740 24612 12750
rect 24556 12646 24612 12684
rect 25228 12738 25284 16830
rect 26684 16772 26740 18284
rect 27580 17778 27636 17790
rect 27580 17726 27582 17778
rect 27634 17726 27636 17778
rect 27580 17668 27636 17726
rect 27580 17602 27636 17612
rect 26908 17442 26964 17454
rect 26908 17390 26910 17442
rect 26962 17390 26964 17442
rect 26908 17108 26964 17390
rect 27804 17332 27860 20748
rect 27916 21698 27972 21710
rect 27916 21646 27918 21698
rect 27970 21646 27972 21698
rect 27916 19348 27972 21646
rect 29372 21700 29428 21710
rect 29148 21028 29204 21038
rect 28476 20802 28532 20814
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28476 20244 28532 20750
rect 29148 20802 29204 20972
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20738 29204 20750
rect 29372 20802 29428 21644
rect 30156 21586 30212 21598
rect 30156 21534 30158 21586
rect 30210 21534 30212 21586
rect 29596 20916 29652 20926
rect 30044 20916 30100 20926
rect 29596 20914 30100 20916
rect 29596 20862 29598 20914
rect 29650 20862 30046 20914
rect 30098 20862 30100 20914
rect 29596 20860 30100 20862
rect 29596 20850 29652 20860
rect 30044 20850 30100 20860
rect 30156 20914 30212 21534
rect 30318 21196 30582 21206
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30318 21130 30582 21140
rect 30156 20862 30158 20914
rect 30210 20862 30212 20914
rect 30156 20850 30212 20862
rect 30716 20916 30772 22876
rect 30940 22370 30996 22382
rect 30940 22318 30942 22370
rect 30994 22318 30996 22370
rect 30940 22148 30996 22318
rect 31388 22148 31444 22158
rect 30940 22146 31444 22148
rect 30940 22094 31390 22146
rect 31442 22094 31444 22146
rect 30940 22092 31444 22094
rect 30716 20850 30772 20860
rect 30828 21586 30884 21598
rect 30828 21534 30830 21586
rect 30882 21534 30884 21586
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 29372 20738 29428 20750
rect 30380 20804 30436 20814
rect 30380 20710 30436 20748
rect 29708 20692 29764 20702
rect 29708 20598 29764 20636
rect 28476 20178 28532 20188
rect 29932 20580 29988 20590
rect 28924 20132 28980 20142
rect 28924 20038 28980 20076
rect 29708 20130 29764 20142
rect 29708 20078 29710 20130
rect 29762 20078 29764 20130
rect 28476 20020 28532 20030
rect 28476 19906 28532 19964
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28476 19842 28532 19854
rect 27916 19282 27972 19292
rect 28476 19234 28532 19246
rect 28476 19182 28478 19234
rect 28530 19182 28532 19234
rect 28476 19124 28532 19182
rect 28476 19058 28532 19068
rect 29036 19010 29092 19022
rect 29036 18958 29038 19010
rect 29090 18958 29092 19010
rect 29036 18452 29092 18958
rect 29708 19012 29764 20078
rect 29820 19012 29876 19022
rect 29708 18956 29820 19012
rect 29820 18918 29876 18956
rect 27580 17276 27860 17332
rect 27916 17668 27972 17678
rect 27580 17108 27636 17276
rect 26908 17106 27636 17108
rect 26908 17054 27582 17106
rect 27634 17054 27636 17106
rect 26908 17052 27636 17054
rect 27580 17042 27636 17052
rect 27692 17108 27748 17118
rect 26684 16706 26740 16716
rect 27356 16772 27412 16782
rect 27356 16678 27412 16716
rect 27692 16770 27748 17052
rect 27692 16718 27694 16770
rect 27746 16718 27748 16770
rect 27692 16706 27748 16718
rect 25228 12686 25230 12738
rect 25282 12686 25284 12738
rect 24556 12180 24612 12190
rect 24556 11394 24612 12124
rect 25004 11508 25060 11518
rect 25228 11508 25284 12686
rect 25564 16658 25620 16670
rect 25564 16606 25566 16658
rect 25618 16606 25620 16658
rect 25564 16100 25620 16606
rect 27916 16548 27972 17612
rect 28028 17444 28084 17454
rect 28588 17444 28644 17454
rect 28028 17442 28196 17444
rect 28028 17390 28030 17442
rect 28082 17390 28196 17442
rect 28028 17388 28196 17390
rect 28028 17378 28084 17388
rect 28140 17106 28196 17388
rect 28588 17350 28644 17388
rect 29036 17332 29092 18396
rect 29372 18676 29428 18686
rect 29372 18338 29428 18620
rect 29932 18450 29988 20524
rect 30604 20580 30660 20590
rect 30604 20486 30660 20524
rect 30716 20244 30772 20254
rect 30318 19628 30582 19638
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30318 19562 30582 19572
rect 29932 18398 29934 18450
rect 29986 18398 29988 18450
rect 29932 18386 29988 18398
rect 29372 18286 29374 18338
rect 29426 18286 29428 18338
rect 29372 18274 29428 18286
rect 29260 18228 29316 18238
rect 29148 17444 29204 17454
rect 29148 17350 29204 17388
rect 29036 17266 29092 17276
rect 29260 17220 29316 18172
rect 30318 18060 30582 18070
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30318 17994 30582 18004
rect 29932 17892 29988 17902
rect 28140 17054 28142 17106
rect 28194 17054 28196 17106
rect 28140 17042 28196 17054
rect 29148 17164 29316 17220
rect 29372 17890 29988 17892
rect 29372 17838 29934 17890
rect 29986 17838 29988 17890
rect 29372 17836 29988 17838
rect 29148 17106 29204 17164
rect 29148 17054 29150 17106
rect 29202 17054 29204 17106
rect 29148 17042 29204 17054
rect 28700 16996 28756 17006
rect 28700 16902 28756 16940
rect 29260 16996 29316 17006
rect 28476 16884 28532 16894
rect 28476 16770 28532 16828
rect 28476 16718 28478 16770
rect 28530 16718 28532 16770
rect 28476 16706 28532 16718
rect 29036 16882 29092 16894
rect 29036 16830 29038 16882
rect 29090 16830 29092 16882
rect 27244 16492 27972 16548
rect 25564 11956 25620 16044
rect 26124 16100 26180 16110
rect 26124 15874 26180 16044
rect 26908 16100 26964 16110
rect 26908 16006 26964 16044
rect 26124 15822 26126 15874
rect 26178 15822 26180 15874
rect 26124 15810 26180 15822
rect 26684 15874 26740 15886
rect 26684 15822 26686 15874
rect 26738 15822 26740 15874
rect 26160 15708 26424 15718
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26160 15642 26424 15652
rect 26684 15204 26740 15822
rect 26684 15138 26740 15148
rect 26796 14420 26852 14430
rect 26796 14326 26852 14364
rect 26160 14140 26424 14150
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26160 14074 26424 14084
rect 25788 12852 25844 12862
rect 27132 12852 27188 12862
rect 25788 12850 25956 12852
rect 25788 12798 25790 12850
rect 25842 12798 25956 12850
rect 25788 12796 25956 12798
rect 25788 12786 25844 12796
rect 25788 12290 25844 12302
rect 25788 12238 25790 12290
rect 25842 12238 25844 12290
rect 25676 11956 25732 11966
rect 25564 11954 25732 11956
rect 25564 11902 25678 11954
rect 25730 11902 25732 11954
rect 25564 11900 25732 11902
rect 25676 11890 25732 11900
rect 25060 11452 25284 11508
rect 25004 11414 25060 11452
rect 24556 11342 24558 11394
rect 24610 11342 24612 11394
rect 24556 11284 24612 11342
rect 24556 11218 24612 11228
rect 24556 10724 24612 10734
rect 24556 10630 24612 10668
rect 25564 10724 25620 10734
rect 25564 10630 25620 10668
rect 24668 10612 24724 10622
rect 24668 10498 24724 10556
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10434 24724 10446
rect 25228 10500 25284 10510
rect 25228 9826 25284 10444
rect 25564 10050 25620 10062
rect 25564 9998 25566 10050
rect 25618 9998 25620 10050
rect 25564 9940 25620 9998
rect 25564 9874 25620 9884
rect 25228 9774 25230 9826
rect 25282 9774 25284 9826
rect 25228 9762 25284 9774
rect 25116 9716 25172 9726
rect 25116 9622 25172 9660
rect 24556 9044 24612 9054
rect 24556 8950 24612 8988
rect 25788 8932 25844 12238
rect 25900 11172 25956 12796
rect 26160 12572 26424 12582
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26160 12506 26424 12516
rect 26124 12178 26180 12190
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 26124 11732 26180 12126
rect 26908 12180 26964 12190
rect 27132 12180 27188 12796
rect 26908 12086 26964 12124
rect 27020 12178 27188 12180
rect 27020 12126 27134 12178
rect 27186 12126 27188 12178
rect 27020 12124 27188 12126
rect 27020 11844 27076 12124
rect 27132 12114 27188 12124
rect 26124 11506 26180 11676
rect 26124 11454 26126 11506
rect 26178 11454 26180 11506
rect 26124 11442 26180 11454
rect 26796 11788 27076 11844
rect 26684 11396 26740 11406
rect 26684 11302 26740 11340
rect 25900 9156 25956 11116
rect 26160 11004 26424 11014
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26160 10938 26424 10948
rect 26012 10500 26068 10510
rect 26012 9268 26068 10444
rect 26460 9940 26516 9950
rect 26516 9884 26628 9940
rect 26460 9874 26516 9884
rect 26348 9828 26404 9838
rect 26348 9734 26404 9772
rect 26160 9436 26424 9446
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26160 9370 26424 9380
rect 26012 9212 26180 9268
rect 25900 9042 25956 9100
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25900 8978 25956 8990
rect 26124 9042 26180 9212
rect 26124 8990 26126 9042
rect 26178 8990 26180 9042
rect 26124 8978 26180 8990
rect 25788 8838 25844 8876
rect 24668 8818 24724 8830
rect 24668 8766 24670 8818
rect 24722 8766 24724 8818
rect 24668 8260 24724 8766
rect 26460 8820 26516 8830
rect 26460 8726 26516 8764
rect 26572 8484 26628 9884
rect 26684 9828 26740 9838
rect 26796 9828 26852 11788
rect 27020 11394 27076 11406
rect 27020 11342 27022 11394
rect 27074 11342 27076 11394
rect 27020 10724 27076 11342
rect 27020 10658 27076 10668
rect 27244 10612 27300 16492
rect 28924 16100 28980 16110
rect 27468 15876 27524 15886
rect 27468 15874 27748 15876
rect 27468 15822 27470 15874
rect 27522 15822 27748 15874
rect 27468 15820 27748 15822
rect 27468 15810 27524 15820
rect 27468 15540 27524 15550
rect 27468 15446 27524 15484
rect 27692 14420 27748 15820
rect 27804 15874 27860 15886
rect 27804 15822 27806 15874
rect 27858 15822 27860 15874
rect 27804 15540 27860 15822
rect 28140 15876 28196 15886
rect 28140 15782 28196 15820
rect 27804 15474 27860 15484
rect 28700 15652 28756 15662
rect 28700 15538 28756 15596
rect 28700 15486 28702 15538
rect 28754 15486 28756 15538
rect 28700 15474 28756 15486
rect 28924 15428 28980 16044
rect 29036 15988 29092 16830
rect 29260 16882 29316 16940
rect 29260 16830 29262 16882
rect 29314 16830 29316 16882
rect 29260 16818 29316 16830
rect 29372 16660 29428 17836
rect 29932 17826 29988 17836
rect 29260 16604 29428 16660
rect 29484 17668 29540 17678
rect 29484 17554 29540 17612
rect 30268 17668 30324 17678
rect 30268 17574 30324 17612
rect 29484 17502 29486 17554
rect 29538 17502 29540 17554
rect 29260 16210 29316 16604
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 29372 16100 29428 16110
rect 29372 16006 29428 16044
rect 29148 15988 29204 15998
rect 29036 15986 29204 15988
rect 29036 15934 29150 15986
rect 29202 15934 29204 15986
rect 29036 15932 29204 15934
rect 29148 15876 29204 15932
rect 29036 15428 29092 15438
rect 28924 15426 29092 15428
rect 28924 15374 29038 15426
rect 29090 15374 29092 15426
rect 28924 15372 29092 15374
rect 29036 15362 29092 15372
rect 28924 15204 28980 15214
rect 28700 15092 28756 15102
rect 27692 14364 27972 14420
rect 27580 14308 27636 14318
rect 27636 14252 27860 14308
rect 27580 14214 27636 14252
rect 27468 13972 27524 13982
rect 27468 13878 27524 13916
rect 27804 13860 27860 14252
rect 27804 13746 27860 13804
rect 27804 13694 27806 13746
rect 27858 13694 27860 13746
rect 27804 13682 27860 13694
rect 27916 12404 27972 14364
rect 28588 13860 28644 13870
rect 28588 13766 28644 13804
rect 28476 13746 28532 13758
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28028 13636 28084 13646
rect 28476 13636 28532 13694
rect 28028 13634 28532 13636
rect 28028 13582 28030 13634
rect 28082 13582 28532 13634
rect 28028 13580 28532 13582
rect 28028 13570 28084 13580
rect 27916 12348 28084 12404
rect 27580 11396 27636 11406
rect 27356 11340 27580 11396
rect 27356 10834 27412 11340
rect 27580 11302 27636 11340
rect 27356 10782 27358 10834
rect 27410 10782 27412 10834
rect 27356 10770 27412 10782
rect 27916 11282 27972 11294
rect 27916 11230 27918 11282
rect 27970 11230 27972 11282
rect 27916 10836 27972 11230
rect 27916 10770 27972 10780
rect 28028 10834 28084 12348
rect 28028 10782 28030 10834
rect 28082 10782 28084 10834
rect 28028 10724 28084 10782
rect 28028 10658 28084 10668
rect 28252 11170 28308 11182
rect 28252 11118 28254 11170
rect 28306 11118 28308 11170
rect 28252 10612 28308 11118
rect 28476 10948 28532 13580
rect 28700 11732 28756 15036
rect 28924 14644 28980 15148
rect 28924 14578 28980 14588
rect 29036 14532 29092 14542
rect 29148 14532 29204 15820
rect 29260 15988 29316 15998
rect 29260 15314 29316 15932
rect 29260 15262 29262 15314
rect 29314 15262 29316 15314
rect 29260 15250 29316 15262
rect 29484 14868 29540 17502
rect 30044 17442 30100 17454
rect 30044 17390 30046 17442
rect 30098 17390 30100 17442
rect 29932 17332 29988 17342
rect 29596 16996 29652 17006
rect 29596 16902 29652 16940
rect 29932 16882 29988 17276
rect 29932 16830 29934 16882
rect 29986 16830 29988 16882
rect 29932 16818 29988 16830
rect 30044 16324 30100 17390
rect 30604 17442 30660 17454
rect 30604 17390 30606 17442
rect 30658 17390 30660 17442
rect 30604 16996 30660 17390
rect 30604 16930 30660 16940
rect 30318 16492 30582 16502
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30318 16426 30582 16436
rect 30044 16258 30100 16268
rect 29708 15988 29764 15998
rect 29708 15894 29764 15932
rect 30156 15988 30212 15998
rect 29932 15652 29988 15662
rect 29932 15314 29988 15596
rect 29932 15262 29934 15314
rect 29986 15262 29988 15314
rect 29932 15250 29988 15262
rect 29596 15092 29652 15102
rect 29596 15090 30100 15092
rect 29596 15038 29598 15090
rect 29650 15038 30100 15090
rect 29596 15036 30100 15038
rect 29596 15026 29652 15036
rect 29036 14530 29204 14532
rect 29036 14478 29038 14530
rect 29090 14478 29204 14530
rect 29036 14476 29204 14478
rect 29372 14812 29540 14868
rect 29036 13746 29092 14476
rect 29260 14306 29316 14318
rect 29260 14254 29262 14306
rect 29314 14254 29316 14306
rect 29260 13858 29316 14254
rect 29260 13806 29262 13858
rect 29314 13806 29316 13858
rect 29260 13794 29316 13806
rect 29372 13972 29428 14812
rect 29484 14644 29540 14654
rect 29484 14418 29540 14588
rect 30044 14530 30100 15036
rect 30044 14478 30046 14530
rect 30098 14478 30100 14530
rect 30044 14466 30100 14478
rect 29484 14366 29486 14418
rect 29538 14366 29540 14418
rect 29484 14196 29540 14366
rect 29708 14420 29764 14430
rect 29708 14418 29876 14420
rect 29708 14366 29710 14418
rect 29762 14366 29876 14418
rect 29708 14364 29876 14366
rect 29708 14354 29764 14364
rect 29484 14140 29764 14196
rect 29484 13972 29540 13982
rect 29372 13970 29540 13972
rect 29372 13918 29486 13970
rect 29538 13918 29540 13970
rect 29372 13916 29540 13918
rect 29036 13694 29038 13746
rect 29090 13694 29092 13746
rect 29036 13682 29092 13694
rect 28812 13634 28868 13646
rect 28812 13582 28814 13634
rect 28866 13582 28868 13634
rect 28812 13300 28868 13582
rect 29260 13300 29316 13310
rect 28812 13244 29204 13300
rect 29148 13186 29204 13244
rect 29148 13134 29150 13186
rect 29202 13134 29204 13186
rect 29148 13122 29204 13134
rect 29260 12964 29316 13244
rect 29260 12402 29316 12908
rect 29372 12850 29428 13916
rect 29484 13906 29540 13916
rect 29596 13522 29652 13534
rect 29596 13470 29598 13522
rect 29650 13470 29652 13522
rect 29596 13188 29652 13470
rect 29596 13122 29652 13132
rect 29372 12798 29374 12850
rect 29426 12798 29428 12850
rect 29372 12786 29428 12798
rect 29484 13074 29540 13086
rect 29484 13022 29486 13074
rect 29538 13022 29540 13074
rect 29260 12350 29262 12402
rect 29314 12350 29316 12402
rect 29260 12338 29316 12350
rect 28700 11666 28756 11676
rect 29484 11620 29540 13022
rect 29708 13076 29764 14140
rect 29820 13300 29876 14364
rect 30156 13746 30212 15932
rect 30604 15988 30660 15998
rect 30604 15894 30660 15932
rect 30716 15148 30772 20188
rect 30828 19236 30884 21534
rect 30828 19170 30884 19180
rect 30828 17780 30884 17790
rect 30940 17780 30996 22092
rect 31388 22082 31444 22092
rect 31276 21698 31332 21710
rect 31276 21646 31278 21698
rect 31330 21646 31332 21698
rect 31164 21588 31220 21598
rect 31052 21476 31108 21486
rect 31052 21382 31108 21420
rect 30884 17724 30996 17780
rect 31052 21140 31108 21150
rect 30828 17714 30884 17724
rect 31052 15202 31108 21084
rect 31164 18676 31220 21532
rect 31276 20804 31332 21646
rect 31388 21362 31444 21374
rect 31388 21310 31390 21362
rect 31442 21310 31444 21362
rect 31388 21028 31444 21310
rect 31612 21140 31668 24668
rect 31612 21074 31668 21084
rect 31836 21474 31892 21486
rect 31836 21422 31838 21474
rect 31890 21422 31892 21474
rect 31388 20972 31556 21028
rect 31500 20916 31556 20972
rect 31500 20860 31780 20916
rect 31276 20738 31332 20748
rect 31164 18610 31220 18620
rect 31388 20578 31444 20590
rect 31388 20526 31390 20578
rect 31442 20526 31444 20578
rect 31388 19012 31444 20526
rect 31724 20020 31780 20860
rect 31836 20244 31892 21422
rect 33628 21364 33684 21374
rect 33628 20802 33684 21308
rect 34076 21028 34132 25200
rect 34476 21980 34740 21990
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34476 21914 34740 21924
rect 33628 20750 33630 20802
rect 33682 20750 33684 20802
rect 33628 20738 33684 20750
rect 33964 20972 34132 21028
rect 31836 20178 31892 20188
rect 31948 20020 32004 20030
rect 31724 20018 32004 20020
rect 31724 19966 31950 20018
rect 32002 19966 32004 20018
rect 31724 19964 32004 19966
rect 31948 19954 32004 19964
rect 32620 20020 32676 20030
rect 32620 20018 32788 20020
rect 32620 19966 32622 20018
rect 32674 19966 32788 20018
rect 32620 19964 32788 19966
rect 32620 19954 32676 19964
rect 31388 17444 31444 18956
rect 32060 19234 32116 19246
rect 32060 19182 32062 19234
rect 32114 19182 32116 19234
rect 31836 18452 31892 18462
rect 31836 18338 31892 18396
rect 31836 18286 31838 18338
rect 31890 18286 31892 18338
rect 31836 18274 31892 18286
rect 31388 17350 31444 17388
rect 32060 17108 32116 19182
rect 32732 19234 32788 19964
rect 33292 19906 33348 19918
rect 33292 19854 33294 19906
rect 33346 19854 33348 19906
rect 32732 19182 32734 19234
rect 32786 19182 32788 19234
rect 32732 19012 32788 19182
rect 33180 19236 33236 19246
rect 33180 19142 33236 19180
rect 33292 19124 33348 19854
rect 33964 19460 34020 20972
rect 33964 19394 34020 19404
rect 34076 20802 34132 20814
rect 34076 20750 34078 20802
rect 34130 20750 34132 20802
rect 33852 19348 33908 19358
rect 32956 19012 33012 19022
rect 32732 18956 32956 19012
rect 32956 18918 33012 18956
rect 33292 18564 33348 19068
rect 33740 19236 33796 19246
rect 33740 18674 33796 19180
rect 33852 19122 33908 19292
rect 33852 19070 33854 19122
rect 33906 19070 33908 19122
rect 33852 18900 33908 19070
rect 33852 18834 33908 18844
rect 34076 19012 34132 20750
rect 34476 20412 34740 20422
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34476 20346 34740 20356
rect 34188 19124 34244 19134
rect 34188 19122 34356 19124
rect 34188 19070 34190 19122
rect 34242 19070 34356 19122
rect 34188 19068 34356 19070
rect 34188 19058 34244 19068
rect 33740 18622 33742 18674
rect 33794 18622 33796 18674
rect 33740 18610 33796 18622
rect 33180 18508 33348 18564
rect 33068 18228 33124 18238
rect 33068 18134 33124 18172
rect 32060 17042 32116 17052
rect 31724 16996 31780 17006
rect 31612 16884 31668 16894
rect 31612 16790 31668 16828
rect 31052 15150 31054 15202
rect 31106 15150 31108 15202
rect 30716 15092 30884 15148
rect 31052 15138 31108 15150
rect 31388 15874 31444 15886
rect 31388 15822 31390 15874
rect 31442 15822 31444 15874
rect 31388 15148 31444 15822
rect 31612 15204 31668 15214
rect 30318 14924 30582 14934
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30318 14858 30582 14868
rect 30604 14530 30660 14542
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14308 30660 14478
rect 30828 14308 30884 15092
rect 31388 15092 31668 15148
rect 31388 14420 31444 15092
rect 31724 14530 31780 16940
rect 31724 14478 31726 14530
rect 31778 14478 31780 14530
rect 31724 14466 31780 14478
rect 30604 14252 30996 14308
rect 30156 13694 30158 13746
rect 30210 13694 30212 13746
rect 30156 13682 30212 13694
rect 30716 13524 30772 13534
rect 30318 13356 30582 13366
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 29820 13244 30100 13300
rect 30318 13290 30582 13300
rect 30044 13188 30100 13244
rect 30380 13188 30436 13198
rect 30716 13188 30772 13468
rect 30044 13186 30324 13188
rect 30044 13134 30046 13186
rect 30098 13134 30324 13186
rect 30044 13132 30324 13134
rect 30044 13122 30100 13132
rect 29820 13076 29876 13086
rect 29708 13074 29876 13076
rect 29708 13022 29822 13074
rect 29874 13022 29876 13074
rect 29708 13020 29876 13022
rect 29820 13010 29876 13020
rect 30268 12964 30324 13132
rect 30380 13186 30772 13188
rect 30380 13134 30382 13186
rect 30434 13134 30772 13186
rect 30380 13132 30772 13134
rect 30380 13122 30436 13132
rect 30604 12964 30660 12974
rect 30268 12962 30660 12964
rect 30268 12910 30606 12962
rect 30658 12910 30660 12962
rect 30268 12908 30660 12910
rect 29596 12178 29652 12190
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29596 11732 29652 12126
rect 30268 12178 30324 12908
rect 30604 12898 30660 12908
rect 30268 12126 30270 12178
rect 30322 12126 30324 12178
rect 30268 12114 30324 12126
rect 30318 11788 30582 11798
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 29652 11676 29876 11732
rect 30318 11722 30582 11732
rect 29596 11666 29652 11676
rect 29484 11554 29540 11564
rect 29820 11508 29876 11676
rect 29820 11414 29876 11452
rect 30828 11508 30884 11518
rect 28476 10882 28532 10892
rect 30716 11394 30772 11406
rect 30716 11342 30718 11394
rect 30770 11342 30772 11394
rect 27244 10556 27412 10612
rect 26684 9826 26852 9828
rect 26684 9774 26686 9826
rect 26738 9774 26852 9826
rect 26684 9772 26852 9774
rect 26684 9762 26740 9772
rect 26796 8820 26852 9772
rect 25788 8372 25844 8382
rect 25788 8278 25844 8316
rect 26460 8372 26628 8428
rect 26684 8764 26852 8820
rect 26908 9828 26964 9838
rect 24668 8194 24724 8204
rect 25900 8260 25956 8270
rect 26236 8260 26292 8270
rect 25900 8166 25956 8204
rect 26124 8258 26292 8260
rect 26124 8206 26238 8258
rect 26290 8206 26292 8258
rect 26124 8204 26292 8206
rect 25788 8148 25844 8158
rect 25228 8034 25284 8046
rect 25228 7982 25230 8034
rect 25282 7982 25284 8034
rect 24780 7924 24836 7934
rect 24780 7476 24836 7868
rect 24780 7410 24836 7420
rect 25228 7140 25284 7982
rect 25788 8036 25844 8092
rect 26124 8036 26180 8204
rect 26236 8194 26292 8204
rect 26460 8258 26516 8372
rect 26460 8206 26462 8258
rect 26514 8206 26516 8258
rect 26460 8194 26516 8206
rect 25788 7980 26180 8036
rect 26236 8036 26292 8074
rect 25788 7698 25844 7980
rect 26236 7970 26292 7980
rect 26460 8036 26516 8046
rect 26516 7980 26628 8036
rect 26460 7970 26516 7980
rect 26160 7868 26424 7878
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26160 7802 26424 7812
rect 25788 7646 25790 7698
rect 25842 7646 25844 7698
rect 25788 7634 25844 7646
rect 26572 7588 26628 7980
rect 26460 7532 26572 7588
rect 26124 7362 26180 7374
rect 26124 7310 26126 7362
rect 26178 7310 26180 7362
rect 26124 7140 26180 7310
rect 24444 5842 24500 5852
rect 25116 7084 25228 7140
rect 25116 4900 25172 7084
rect 25228 7074 25284 7084
rect 25900 7084 26124 7140
rect 25900 6130 25956 7084
rect 26124 7074 26180 7084
rect 26460 6690 26516 7532
rect 26572 7494 26628 7532
rect 26460 6638 26462 6690
rect 26514 6638 26516 6690
rect 26460 6626 26516 6638
rect 26572 6580 26628 6590
rect 26572 6486 26628 6524
rect 26160 6300 26424 6310
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26160 6234 26424 6244
rect 25900 6078 25902 6130
rect 25954 6078 25956 6130
rect 25900 6066 25956 6078
rect 26684 5684 26740 8764
rect 26908 8708 26964 9772
rect 27244 9156 27300 9166
rect 27244 9062 27300 9100
rect 26796 8652 26964 8708
rect 26796 7698 26852 8652
rect 26908 8484 26964 8494
rect 27356 8428 27412 10556
rect 28252 10546 28308 10556
rect 30380 10612 30436 10622
rect 30380 10518 30436 10556
rect 30318 10220 30582 10230
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30318 10154 30582 10164
rect 28700 9268 28756 9278
rect 28588 9266 28756 9268
rect 28588 9214 28702 9266
rect 28754 9214 28756 9266
rect 28588 9212 28756 9214
rect 28476 9042 28532 9054
rect 28476 8990 28478 9042
rect 28530 8990 28532 9042
rect 26908 8372 27076 8428
rect 27356 8372 27524 8428
rect 27020 8370 27076 8372
rect 27020 8318 27022 8370
rect 27074 8318 27076 8370
rect 27020 8306 27076 8318
rect 26796 7646 26798 7698
rect 26850 7646 26852 7698
rect 26796 7634 26852 7646
rect 27020 7586 27076 7598
rect 27020 7534 27022 7586
rect 27074 7534 27076 7586
rect 27020 7476 27076 7534
rect 27356 7588 27412 7598
rect 27356 7494 27412 7532
rect 27020 7420 27300 7476
rect 27244 7364 27300 7420
rect 27244 7308 27412 7364
rect 27132 7252 27188 7262
rect 27132 7250 27300 7252
rect 27132 7198 27134 7250
rect 27186 7198 27300 7250
rect 27132 7196 27300 7198
rect 27132 7186 27188 7196
rect 26796 6804 26852 6814
rect 26796 6690 26852 6748
rect 26796 6638 26798 6690
rect 26850 6638 26852 6690
rect 26796 6626 26852 6638
rect 26908 6690 26964 6702
rect 27132 6692 27188 6702
rect 26908 6638 26910 6690
rect 26962 6638 26964 6690
rect 26908 6020 26964 6638
rect 26908 5796 26964 5964
rect 26684 5618 26740 5628
rect 26796 5740 26964 5796
rect 27020 6636 27132 6692
rect 25788 5348 25844 5358
rect 25788 5254 25844 5292
rect 26796 5348 26852 5740
rect 27020 5460 27076 6636
rect 27132 6626 27188 6636
rect 27244 6690 27300 7196
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 27244 6626 27300 6638
rect 27356 6468 27412 7308
rect 27468 6692 27524 8372
rect 28476 8372 28532 8990
rect 28588 9044 28644 9212
rect 28700 9202 28756 9212
rect 29596 9268 29652 9278
rect 28924 9044 28980 9054
rect 28588 8978 28644 8988
rect 28700 9042 28980 9044
rect 28700 8990 28926 9042
rect 28978 8990 28980 9042
rect 28700 8988 28980 8990
rect 28476 8306 28532 8316
rect 27692 7586 27748 7598
rect 27692 7534 27694 7586
rect 27746 7534 27748 7586
rect 27692 7364 27748 7534
rect 28700 7586 28756 8988
rect 28924 8978 28980 8988
rect 29484 9044 29540 9082
rect 29484 8978 29540 8988
rect 29484 8820 29540 8830
rect 28700 7534 28702 7586
rect 28754 7534 28756 7586
rect 28476 7474 28532 7486
rect 28476 7422 28478 7474
rect 28530 7422 28532 7474
rect 28476 7364 28532 7422
rect 27748 7308 27972 7364
rect 27692 7298 27748 7308
rect 27468 6626 27524 6636
rect 27916 6692 27972 7308
rect 28476 7298 28532 7308
rect 28252 6804 28308 6814
rect 28252 6710 28308 6748
rect 27916 6598 27972 6636
rect 28588 6580 28644 6590
rect 28588 6486 28644 6524
rect 27692 6468 27748 6478
rect 27356 6412 27692 6468
rect 27692 6374 27748 6412
rect 27804 6466 27860 6478
rect 27804 6414 27806 6466
rect 27858 6414 27860 6466
rect 26796 5282 26852 5292
rect 26908 5404 27076 5460
rect 25116 4806 25172 4844
rect 25900 5012 25956 5022
rect 22652 4470 22708 4508
rect 23436 4562 24052 4564
rect 23436 4510 23998 4562
rect 24050 4510 24052 4562
rect 23436 4508 24052 4510
rect 23436 4450 23492 4508
rect 23996 4498 24052 4508
rect 25676 4564 25732 4574
rect 25900 4564 25956 4956
rect 26908 5012 26964 5404
rect 27804 5124 27860 6414
rect 26908 4946 26964 4956
rect 27132 5068 27860 5124
rect 28364 6468 28420 6478
rect 28364 5124 28420 6412
rect 28700 6356 28756 7534
rect 28588 6300 28700 6356
rect 26160 4732 26424 4742
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26160 4666 26424 4676
rect 25676 4562 25956 4564
rect 25676 4510 25678 4562
rect 25730 4510 25956 4562
rect 25676 4508 25956 4510
rect 25676 4498 25732 4508
rect 23436 4398 23438 4450
rect 23490 4398 23492 4450
rect 23436 4386 23492 4398
rect 25900 4450 25956 4508
rect 25900 4398 25902 4450
rect 25954 4398 25956 4450
rect 25900 4386 25956 4398
rect 22316 4286 22318 4338
rect 22370 4286 22372 4338
rect 22316 4274 22372 4286
rect 26460 4340 26516 4350
rect 26460 4246 26516 4284
rect 26908 4338 26964 4350
rect 26908 4286 26910 4338
rect 26962 4286 26964 4338
rect 26908 4228 26964 4286
rect 27132 4228 27188 5068
rect 28364 5058 28420 5068
rect 28476 5122 28532 5134
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 26908 4172 27188 4228
rect 27580 4898 27636 4910
rect 27580 4846 27582 4898
rect 27634 4846 27636 4898
rect 23548 4114 23604 4126
rect 23548 4062 23550 4114
rect 23602 4062 23604 4114
rect 22002 3948 22266 3958
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22002 3882 22266 3892
rect 19964 3614 19966 3666
rect 20018 3614 20020 3666
rect 19964 3602 20020 3614
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 23324 3668 23380 3678
rect 20076 3556 20132 3566
rect 20076 3462 20132 3500
rect 20748 3556 20804 3566
rect 20748 3462 20804 3500
rect 23324 800 23380 3612
rect 23548 3556 23604 4062
rect 26012 4114 26068 4126
rect 26012 4062 26014 4114
rect 26066 4062 26068 4114
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3556 24612 3566
rect 23548 3554 24612 3556
rect 23548 3502 24558 3554
rect 24610 3502 24612 3554
rect 23548 3500 24612 3502
rect 24556 3490 24612 3500
rect 26012 3556 26068 4062
rect 27580 3780 27636 4846
rect 28476 4228 28532 5070
rect 28588 4340 28644 6300
rect 28700 6262 28756 6300
rect 28812 8708 28868 8718
rect 28700 6020 28756 6030
rect 28700 5926 28756 5964
rect 28812 5794 28868 8652
rect 29260 8372 29316 8382
rect 29260 8278 29316 8316
rect 29260 7476 29316 7486
rect 29484 7476 29540 8764
rect 29596 8370 29652 9212
rect 30318 8652 30582 8662
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30318 8586 30582 8596
rect 29596 8318 29598 8370
rect 29650 8318 29652 8370
rect 29596 8306 29652 8318
rect 29820 8148 29876 8158
rect 30156 8148 30212 8158
rect 29820 8054 29876 8092
rect 29932 8146 30212 8148
rect 29932 8094 30158 8146
rect 30210 8094 30212 8146
rect 29932 8092 30212 8094
rect 29932 7812 29988 8092
rect 30156 8082 30212 8092
rect 29596 7756 29988 7812
rect 29596 7698 29652 7756
rect 29596 7646 29598 7698
rect 29650 7646 29652 7698
rect 29596 7634 29652 7646
rect 29932 7476 29988 7486
rect 29316 7420 29428 7476
rect 29484 7474 29988 7476
rect 29484 7422 29934 7474
rect 29986 7422 29988 7474
rect 29484 7420 29988 7422
rect 29260 7382 29316 7420
rect 29036 7362 29092 7374
rect 29036 7310 29038 7362
rect 29090 7310 29092 7362
rect 29036 6916 29092 7310
rect 29372 7252 29428 7420
rect 29932 7410 29988 7420
rect 29372 7196 29876 7252
rect 29036 6850 29092 6860
rect 29596 6804 29652 6814
rect 29596 6710 29652 6748
rect 29820 6802 29876 7196
rect 30318 7084 30582 7094
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30318 7018 30582 7028
rect 29820 6750 29822 6802
rect 29874 6750 29876 6802
rect 29820 6738 29876 6750
rect 29372 6690 29428 6702
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 28812 5742 28814 5794
rect 28866 5742 28868 5794
rect 28812 5730 28868 5742
rect 29260 5908 29316 5918
rect 29260 5346 29316 5852
rect 29260 5294 29262 5346
rect 29314 5294 29316 5346
rect 29260 5282 29316 5294
rect 29372 5234 29428 6638
rect 29932 6692 29988 6702
rect 30156 6692 30212 6702
rect 29988 6636 30100 6692
rect 29932 6626 29988 6636
rect 30044 6578 30100 6636
rect 30156 6598 30212 6636
rect 30604 6692 30660 6702
rect 30716 6692 30772 11342
rect 30828 10836 30884 11452
rect 30828 10610 30884 10780
rect 30828 10558 30830 10610
rect 30882 10558 30884 10610
rect 30828 10546 30884 10558
rect 30940 8428 30996 14252
rect 31388 12850 31444 14364
rect 33068 13748 33124 13758
rect 33068 13654 33124 13692
rect 31836 13636 31892 13646
rect 31836 13542 31892 13580
rect 33180 13524 33236 18508
rect 33404 18452 33460 18462
rect 33292 18450 33460 18452
rect 33292 18398 33406 18450
rect 33458 18398 33460 18450
rect 33292 18396 33460 18398
rect 33292 17668 33348 18396
rect 33404 18386 33460 18396
rect 33964 18450 34020 18462
rect 33964 18398 33966 18450
rect 34018 18398 34020 18450
rect 33404 18228 33460 18238
rect 33404 18226 33684 18228
rect 33404 18174 33406 18226
rect 33458 18174 33684 18226
rect 33404 18172 33684 18174
rect 33404 18162 33460 18172
rect 33292 17602 33348 17612
rect 33628 17666 33684 18172
rect 33628 17614 33630 17666
rect 33682 17614 33684 17666
rect 33628 17602 33684 17614
rect 33628 17444 33684 17454
rect 33628 16882 33684 17388
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33628 16818 33684 16830
rect 33628 16324 33684 16334
rect 33628 16098 33684 16268
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 16034 33684 16046
rect 33964 16100 34020 18398
rect 34076 17666 34132 18956
rect 34076 17614 34078 17666
rect 34130 17614 34132 17666
rect 34076 17602 34132 17614
rect 34188 18900 34244 18910
rect 34188 17106 34244 18844
rect 34188 17054 34190 17106
rect 34242 17054 34244 17106
rect 34188 17042 34244 17054
rect 34076 16100 34132 16110
rect 33964 16098 34132 16100
rect 33964 16046 34078 16098
rect 34130 16046 34132 16098
rect 33964 16044 34132 16046
rect 33516 15316 33572 15326
rect 33516 14754 33572 15260
rect 33516 14702 33518 14754
rect 33570 14702 33572 14754
rect 33516 14690 33572 14702
rect 33516 13634 33572 13646
rect 33516 13582 33518 13634
rect 33570 13582 33572 13634
rect 33516 13524 33572 13582
rect 31388 12798 31390 12850
rect 31442 12798 31444 12850
rect 31388 12786 31444 12798
rect 33068 13468 33572 13524
rect 31836 12068 31892 12078
rect 31836 11974 31892 12012
rect 31164 11620 31220 11630
rect 31164 11394 31220 11564
rect 31164 11342 31166 11394
rect 31218 11342 31220 11394
rect 31164 11330 31220 11342
rect 31836 10948 31892 10958
rect 30604 6690 30772 6692
rect 30604 6638 30606 6690
rect 30658 6638 30772 6690
rect 30604 6636 30772 6638
rect 30828 8372 30996 8428
rect 31388 10836 31444 10846
rect 30044 6526 30046 6578
rect 30098 6526 30100 6578
rect 30044 6514 30100 6526
rect 30268 6580 30324 6590
rect 30268 6486 30324 6524
rect 29596 6468 29652 6478
rect 29596 5908 29652 6412
rect 30604 6356 30660 6636
rect 30604 6290 30660 6300
rect 29596 5814 29652 5852
rect 30044 5906 30100 5918
rect 30044 5854 30046 5906
rect 30098 5854 30100 5906
rect 29372 5182 29374 5234
rect 29426 5182 29428 5234
rect 29372 5170 29428 5182
rect 29484 5348 29540 5358
rect 29372 4564 29428 4574
rect 29484 4564 29540 5292
rect 30044 5236 30100 5854
rect 30318 5516 30582 5526
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30318 5450 30582 5460
rect 29596 5234 30100 5236
rect 29596 5182 30046 5234
rect 30098 5182 30100 5234
rect 29596 5180 30100 5182
rect 29596 5122 29652 5180
rect 29596 5070 29598 5122
rect 29650 5070 29652 5122
rect 29596 5058 29652 5070
rect 29932 5012 29988 5022
rect 29932 4918 29988 4956
rect 29372 4562 29540 4564
rect 29372 4510 29374 4562
rect 29426 4510 29540 4562
rect 29372 4508 29540 4510
rect 29932 4564 29988 4574
rect 30044 4564 30100 5180
rect 30716 5124 30772 5134
rect 29932 4562 30100 4564
rect 29932 4510 29934 4562
rect 29986 4510 30100 4562
rect 29932 4508 30100 4510
rect 30492 5122 30772 5124
rect 30492 5070 30718 5122
rect 30770 5070 30772 5122
rect 30492 5068 30772 5070
rect 30492 4562 30548 5068
rect 30716 5058 30772 5068
rect 30828 4564 30884 8372
rect 31276 8146 31332 8158
rect 31276 8094 31278 8146
rect 31330 8094 31332 8146
rect 30940 8034 30996 8046
rect 30940 7982 30942 8034
rect 30994 7982 30996 8034
rect 30940 5796 30996 7982
rect 31164 6692 31220 6702
rect 31164 6598 31220 6636
rect 31052 6580 31108 6590
rect 31052 6130 31108 6524
rect 31052 6078 31054 6130
rect 31106 6078 31108 6130
rect 31052 6066 31108 6078
rect 31164 6468 31220 6478
rect 31164 6018 31220 6412
rect 31164 5966 31166 6018
rect 31218 5966 31220 6018
rect 31164 5954 31220 5966
rect 30940 5730 30996 5740
rect 31276 5684 31332 8094
rect 31388 6132 31444 10780
rect 31836 9826 31892 10892
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31836 9762 31892 9774
rect 32060 9604 32116 9614
rect 32060 9266 32116 9548
rect 32060 9214 32062 9266
rect 32114 9214 32116 9266
rect 31612 8258 31668 8270
rect 31612 8206 31614 8258
rect 31666 8206 31668 8258
rect 31612 7700 31668 8206
rect 31612 7634 31668 7644
rect 31836 7476 31892 7486
rect 31836 7362 31892 7420
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31836 7298 31892 7310
rect 32060 6580 32116 9214
rect 32620 9268 32676 9278
rect 32620 9174 32676 9212
rect 32844 9044 32900 9054
rect 31388 6066 31444 6076
rect 31836 6132 31892 6142
rect 31836 6038 31892 6076
rect 31500 5906 31556 5918
rect 31500 5854 31502 5906
rect 31554 5854 31556 5906
rect 31500 5796 31556 5854
rect 31500 5730 31556 5740
rect 31276 5618 31332 5628
rect 32060 5348 32116 6524
rect 32172 7364 32228 7374
rect 32172 6130 32228 7308
rect 32172 6078 32174 6130
rect 32226 6078 32228 6130
rect 32172 6066 32228 6078
rect 32396 6132 32452 6142
rect 32396 5906 32452 6076
rect 32396 5854 32398 5906
rect 32450 5854 32452 5906
rect 32396 5842 32452 5854
rect 32060 5282 32116 5292
rect 32844 5236 32900 8988
rect 32844 5170 32900 5180
rect 31724 4900 31780 4910
rect 31276 4898 31780 4900
rect 31276 4846 31726 4898
rect 31778 4846 31780 4898
rect 31276 4844 31780 4846
rect 30940 4564 30996 4574
rect 30492 4510 30494 4562
rect 30546 4510 30548 4562
rect 29372 4498 29428 4508
rect 29932 4498 29988 4508
rect 30492 4498 30548 4510
rect 30604 4562 30996 4564
rect 30604 4510 30942 4562
rect 30994 4510 30996 4562
rect 30604 4508 30996 4510
rect 28588 4274 28644 4284
rect 30380 4340 30436 4350
rect 30604 4340 30660 4508
rect 30940 4498 30996 4508
rect 30380 4338 30660 4340
rect 30380 4286 30382 4338
rect 30434 4286 30660 4338
rect 30380 4284 30660 4286
rect 30380 4274 30436 4284
rect 28476 4162 28532 4172
rect 30318 3948 30582 3958
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30318 3882 30582 3892
rect 27580 3714 27636 3724
rect 26012 3490 26068 3500
rect 26908 3668 26964 3678
rect 26160 3164 26424 3174
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26160 3098 26424 3108
rect 26908 800 26964 3612
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3556 28644 3566
rect 28588 3462 28644 3500
rect 30492 924 30884 980
rect 30492 800 30548 924
rect 1792 0 1904 800
rect 5376 0 5488 800
rect 8960 0 9072 800
rect 12544 0 12656 800
rect 16128 0 16240 800
rect 19712 0 19824 800
rect 23296 0 23408 800
rect 26880 0 26992 800
rect 30464 0 30576 800
rect 30828 756 30884 924
rect 31276 756 31332 4844
rect 31724 4834 31780 4844
rect 32172 4564 32228 4574
rect 33068 4564 33124 13468
rect 33628 12964 33684 12974
rect 33628 12870 33684 12908
rect 34076 12962 34132 16044
rect 34076 12910 34078 12962
rect 34130 12910 34132 12962
rect 34076 12852 34132 12910
rect 34076 12786 34132 12796
rect 34188 15204 34244 15214
rect 34300 15148 34356 19068
rect 34476 18844 34740 18854
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34476 18778 34740 18788
rect 34476 17276 34740 17286
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34476 17210 34740 17220
rect 34476 15708 34740 15718
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34476 15642 34740 15652
rect 34188 15092 34356 15148
rect 33628 12178 33684 12190
rect 33628 12126 33630 12178
rect 33682 12126 33684 12178
rect 33628 11396 33684 12126
rect 34188 12178 34244 15092
rect 34476 14140 34740 14150
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34476 14074 34740 14084
rect 34476 12572 34740 12582
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34476 12506 34740 12516
rect 34188 12126 34190 12178
rect 34242 12126 34244 12178
rect 34188 12114 34244 12126
rect 33180 11340 33684 11396
rect 33180 10724 33236 11340
rect 33516 11172 33572 11182
rect 33180 9266 33236 10668
rect 33404 11170 33572 11172
rect 33404 11118 33518 11170
rect 33570 11118 33572 11170
rect 33404 11116 33572 11118
rect 33404 9604 33460 11116
rect 33516 11106 33572 11116
rect 34300 11172 34356 11182
rect 34300 11078 34356 11116
rect 34476 11004 34740 11014
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34476 10938 34740 10948
rect 33516 10612 33572 10622
rect 33516 10050 33572 10556
rect 33516 9998 33518 10050
rect 33570 9998 33572 10050
rect 33516 9986 33572 9998
rect 33404 9538 33460 9548
rect 34476 9436 34740 9446
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34476 9370 34740 9380
rect 33180 9214 33182 9266
rect 33234 9214 33236 9266
rect 33180 8428 33236 9214
rect 33852 9154 33908 9166
rect 33852 9102 33854 9154
rect 33906 9102 33908 9154
rect 33404 9044 33460 9054
rect 33852 9044 33908 9102
rect 33460 8988 33908 9044
rect 33964 9044 34020 9054
rect 33404 8950 33460 8988
rect 33964 8482 34020 8988
rect 33964 8430 33966 8482
rect 34018 8430 34020 8482
rect 33180 8372 33684 8428
rect 33964 8418 34020 8430
rect 34076 9042 34132 9054
rect 34076 8990 34078 9042
rect 34130 8990 34132 9042
rect 33628 7698 33684 8372
rect 33628 7646 33630 7698
rect 33682 7646 33684 7698
rect 33628 7634 33684 7646
rect 33404 7364 33460 7374
rect 33292 7362 33460 7364
rect 33292 7310 33406 7362
rect 33458 7310 33460 7362
rect 33292 7308 33460 7310
rect 33180 6132 33236 6142
rect 33180 6038 33236 6076
rect 33180 5796 33236 5806
rect 33180 4676 33236 5740
rect 33292 5124 33348 7308
rect 33404 7298 33460 7308
rect 33516 6916 33572 6926
rect 33292 5058 33348 5068
rect 33404 6860 33516 6916
rect 33180 4620 33348 4676
rect 32172 4562 33124 4564
rect 32172 4510 32174 4562
rect 32226 4510 33124 4562
rect 32172 4508 33124 4510
rect 32172 4498 32228 4508
rect 33068 4452 33124 4508
rect 33180 4452 33236 4462
rect 33068 4450 33236 4452
rect 33068 4398 33182 4450
rect 33234 4398 33236 4450
rect 33068 4396 33236 4398
rect 33180 4386 33236 4396
rect 32620 4340 32676 4350
rect 32620 4246 32676 4284
rect 33068 4228 33124 4238
rect 33068 4134 33124 4172
rect 33292 4004 33348 4620
rect 32956 3948 33348 4004
rect 32956 3666 33012 3948
rect 32956 3614 32958 3666
rect 33010 3614 33012 3666
rect 32956 3602 33012 3614
rect 31724 3556 31780 3566
rect 31724 3462 31780 3500
rect 33292 3556 33348 3566
rect 32508 3444 32564 3454
rect 32508 3350 32564 3388
rect 33292 1204 33348 3500
rect 33404 3444 33460 6860
rect 33516 6850 33572 6860
rect 34076 6916 34132 8990
rect 34476 7868 34740 7878
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34476 7802 34740 7812
rect 34076 6850 34132 6860
rect 34188 7362 34244 7374
rect 34188 7310 34190 7362
rect 34242 7310 34244 7362
rect 34188 7252 34244 7310
rect 33852 6804 33908 6814
rect 33516 6580 33572 6590
rect 33516 5908 33572 6524
rect 33628 5908 33684 5918
rect 33516 5906 33684 5908
rect 33516 5854 33630 5906
rect 33682 5854 33684 5906
rect 33516 5852 33684 5854
rect 33628 5842 33684 5852
rect 33740 5684 33796 5694
rect 33628 5460 33684 5470
rect 33628 5234 33684 5404
rect 33628 5182 33630 5234
rect 33682 5182 33684 5234
rect 33628 5170 33684 5182
rect 33516 3444 33572 3454
rect 33404 3442 33572 3444
rect 33404 3390 33518 3442
rect 33570 3390 33572 3442
rect 33404 3388 33572 3390
rect 33740 3444 33796 5628
rect 33852 4562 33908 6748
rect 34188 6130 34244 7196
rect 34300 6468 34356 6478
rect 34300 6374 34356 6412
rect 34476 6300 34740 6310
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34476 6234 34740 6244
rect 34188 6078 34190 6130
rect 34242 6078 34244 6130
rect 33852 4510 33854 4562
rect 33906 4510 33908 4562
rect 33852 4498 33908 4510
rect 34076 5908 34132 5918
rect 34076 4340 34132 5852
rect 34188 5796 34244 6078
rect 34188 5730 34244 5740
rect 34188 5124 34244 5134
rect 34244 5068 34356 5124
rect 34188 5030 34244 5068
rect 34076 4246 34132 4284
rect 34300 4340 34356 5068
rect 34476 4732 34740 4742
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34476 4666 34740 4676
rect 34300 4274 34356 4284
rect 34076 3780 34132 3790
rect 33852 3444 33908 3454
rect 33740 3442 33908 3444
rect 33740 3390 33854 3442
rect 33906 3390 33908 3442
rect 33740 3388 33908 3390
rect 33516 3378 33572 3388
rect 33852 3378 33908 3388
rect 33292 1138 33348 1148
rect 34076 800 34132 3724
rect 34188 3444 34244 3454
rect 34188 2772 34244 3388
rect 34476 3164 34740 3174
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34476 3098 34740 3108
rect 34188 2706 34244 2716
rect 30828 700 31332 756
rect 34048 0 34160 800
<< via2 >>
rect 2044 23996 2100 24052
rect 1932 21980 1988 22036
rect 1932 19964 1988 20020
rect 5404 23436 5460 23492
rect 6636 23436 6692 23492
rect 5370 22762 5426 22764
rect 5370 22710 5372 22762
rect 5372 22710 5424 22762
rect 5424 22710 5426 22762
rect 5370 22708 5426 22710
rect 5474 22762 5530 22764
rect 5474 22710 5476 22762
rect 5476 22710 5528 22762
rect 5528 22710 5530 22762
rect 5474 22708 5530 22710
rect 5578 22762 5634 22764
rect 5578 22710 5580 22762
rect 5580 22710 5632 22762
rect 5632 22710 5634 22762
rect 5578 22708 5634 22710
rect 13686 22762 13742 22764
rect 13686 22710 13688 22762
rect 13688 22710 13740 22762
rect 13740 22710 13742 22762
rect 13686 22708 13742 22710
rect 13790 22762 13846 22764
rect 13790 22710 13792 22762
rect 13792 22710 13844 22762
rect 13844 22710 13846 22762
rect 13790 22708 13846 22710
rect 13894 22762 13950 22764
rect 13894 22710 13896 22762
rect 13896 22710 13948 22762
rect 13948 22710 13950 22762
rect 13894 22708 13950 22710
rect 12572 22540 12628 22596
rect 14140 22594 14196 22596
rect 14140 22542 14142 22594
rect 14142 22542 14194 22594
rect 14194 22542 14196 22594
rect 14140 22540 14196 22542
rect 16156 22540 16212 22596
rect 17164 22594 17220 22596
rect 17164 22542 17166 22594
rect 17166 22542 17218 22594
rect 17218 22542 17220 22594
rect 17164 22540 17220 22542
rect 22002 22762 22058 22764
rect 22002 22710 22004 22762
rect 22004 22710 22056 22762
rect 22056 22710 22058 22762
rect 22002 22708 22058 22710
rect 22106 22762 22162 22764
rect 22106 22710 22108 22762
rect 22108 22710 22160 22762
rect 22160 22710 22162 22762
rect 22106 22708 22162 22710
rect 22210 22762 22266 22764
rect 22210 22710 22212 22762
rect 22212 22710 22264 22762
rect 22264 22710 22266 22762
rect 22210 22708 22266 22710
rect 19740 22540 19796 22596
rect 20972 22594 21028 22596
rect 20972 22542 20974 22594
rect 20974 22542 21026 22594
rect 21026 22542 21028 22594
rect 20972 22540 21028 22542
rect 23324 22540 23380 22596
rect 25116 23100 25172 23156
rect 4060 21420 4116 21476
rect 2716 20748 2772 20804
rect 3836 20802 3892 20804
rect 3836 20750 3838 20802
rect 3838 20750 3890 20802
rect 3890 20750 3892 20802
rect 3836 20748 3892 20750
rect 1932 16210 1988 16212
rect 1932 16158 1934 16210
rect 1934 16158 1986 16210
rect 1986 16158 1988 16210
rect 1932 16156 1988 16158
rect 1708 15260 1764 15316
rect 2044 14476 2100 14532
rect 1820 13970 1876 13972
rect 1820 13918 1822 13970
rect 1822 13918 1874 13970
rect 1874 13918 1876 13970
rect 1820 13916 1876 13918
rect 2044 12124 2100 12180
rect 1932 11900 1988 11956
rect 2716 18226 2772 18228
rect 2716 18174 2718 18226
rect 2718 18174 2770 18226
rect 2770 18174 2772 18226
rect 2716 18172 2772 18174
rect 2716 16882 2772 16884
rect 2716 16830 2718 16882
rect 2718 16830 2770 16882
rect 2770 16830 2772 16882
rect 2716 16828 2772 16830
rect 2604 14530 2660 14532
rect 2604 14478 2606 14530
rect 2606 14478 2658 14530
rect 2658 14478 2660 14530
rect 2604 14476 2660 14478
rect 2492 13692 2548 13748
rect 3276 14530 3332 14532
rect 3276 14478 3278 14530
rect 3278 14478 3330 14530
rect 3330 14478 3332 14530
rect 3276 14476 3332 14478
rect 2940 14418 2996 14420
rect 2940 14366 2942 14418
rect 2942 14366 2994 14418
rect 2994 14366 2996 14418
rect 2940 14364 2996 14366
rect 3836 15314 3892 15316
rect 3836 15262 3838 15314
rect 3838 15262 3890 15314
rect 3890 15262 3892 15314
rect 3836 15260 3892 15262
rect 3612 14364 3668 14420
rect 3836 14028 3892 14084
rect 3948 14924 4004 14980
rect 2940 13970 2996 13972
rect 2940 13918 2942 13970
rect 2942 13918 2994 13970
rect 2994 13918 2996 13970
rect 2940 13916 2996 13918
rect 3388 13858 3444 13860
rect 3388 13806 3390 13858
rect 3390 13806 3442 13858
rect 3442 13806 3444 13858
rect 3388 13804 3444 13806
rect 2268 12348 2324 12404
rect 1932 9884 1988 9940
rect 1820 8930 1876 8932
rect 1820 8878 1822 8930
rect 1822 8878 1874 8930
rect 1874 8878 1876 8930
rect 1820 8876 1876 8878
rect 1932 7868 1988 7924
rect 3164 13132 3220 13188
rect 2940 9714 2996 9716
rect 2940 9662 2942 9714
rect 2942 9662 2994 9714
rect 2994 9662 2996 9714
rect 2940 9660 2996 9662
rect 3052 12124 3108 12180
rect 2716 9548 2772 9604
rect 3276 11340 3332 11396
rect 3836 11394 3892 11396
rect 3836 11342 3838 11394
rect 3838 11342 3890 11394
rect 3890 11342 3892 11394
rect 3836 11340 3892 11342
rect 3276 9938 3332 9940
rect 3276 9886 3278 9938
rect 3278 9886 3330 9938
rect 3330 9886 3332 9938
rect 3276 9884 3332 9886
rect 4284 21308 4340 21364
rect 5068 21362 5124 21364
rect 5068 21310 5070 21362
rect 5070 21310 5122 21362
rect 5122 21310 5124 21362
rect 5068 21308 5124 21310
rect 5370 21194 5426 21196
rect 5370 21142 5372 21194
rect 5372 21142 5424 21194
rect 5424 21142 5426 21194
rect 5370 21140 5426 21142
rect 5474 21194 5530 21196
rect 5474 21142 5476 21194
rect 5476 21142 5528 21194
rect 5528 21142 5530 21194
rect 5474 21140 5530 21142
rect 5578 21194 5634 21196
rect 5578 21142 5580 21194
rect 5580 21142 5632 21194
rect 5632 21142 5634 21194
rect 5578 21140 5634 21142
rect 4620 15260 4676 15316
rect 4284 14924 4340 14980
rect 4284 14476 4340 14532
rect 4172 14418 4228 14420
rect 4172 14366 4174 14418
rect 4174 14366 4226 14418
rect 4226 14366 4228 14418
rect 4172 14364 4228 14366
rect 4732 14306 4788 14308
rect 4732 14254 4734 14306
rect 4734 14254 4786 14306
rect 4786 14254 4788 14306
rect 4732 14252 4788 14254
rect 4396 14028 4452 14084
rect 4172 13692 4228 13748
rect 3836 9938 3892 9940
rect 3836 9886 3838 9938
rect 3838 9886 3890 9938
rect 3890 9886 3892 9938
rect 3836 9884 3892 9886
rect 4060 9660 4116 9716
rect 3052 9042 3108 9044
rect 3052 8990 3054 9042
rect 3054 8990 3106 9042
rect 3106 8990 3108 9042
rect 3052 8988 3108 8990
rect 3500 8316 3556 8372
rect 3948 8876 4004 8932
rect 2380 8204 2436 8260
rect 3836 8258 3892 8260
rect 3836 8206 3838 8258
rect 3838 8206 3890 8258
rect 3890 8206 3892 8258
rect 3836 8204 3892 8206
rect 2268 6972 2324 7028
rect 2492 6860 2548 6916
rect 2156 6636 2212 6692
rect 2940 6748 2996 6804
rect 2492 5852 2548 5908
rect 3948 5740 4004 5796
rect 1932 4114 1988 4116
rect 1932 4062 1934 4114
rect 1934 4062 1986 4114
rect 1986 4062 1988 4114
rect 1932 4060 1988 4062
rect 4620 13580 4676 13636
rect 4508 12178 4564 12180
rect 4508 12126 4510 12178
rect 4510 12126 4562 12178
rect 4562 12126 4564 12178
rect 4508 12124 4564 12126
rect 4732 9884 4788 9940
rect 4620 8204 4676 8260
rect 4956 16882 5012 16884
rect 4956 16830 4958 16882
rect 4958 16830 5010 16882
rect 5010 16830 5012 16882
rect 4956 16828 5012 16830
rect 4956 14028 5012 14084
rect 4844 8876 4900 8932
rect 4956 8034 5012 8036
rect 4956 7982 4958 8034
rect 4958 7982 5010 8034
rect 5010 7982 5012 8034
rect 4956 7980 5012 7982
rect 4732 7196 4788 7252
rect 5370 19626 5426 19628
rect 5370 19574 5372 19626
rect 5372 19574 5424 19626
rect 5424 19574 5426 19626
rect 5370 19572 5426 19574
rect 5474 19626 5530 19628
rect 5474 19574 5476 19626
rect 5476 19574 5528 19626
rect 5528 19574 5530 19626
rect 5474 19572 5530 19574
rect 5578 19626 5634 19628
rect 5578 19574 5580 19626
rect 5580 19574 5632 19626
rect 5632 19574 5634 19626
rect 5578 19572 5634 19574
rect 9528 21978 9584 21980
rect 9528 21926 9530 21978
rect 9530 21926 9582 21978
rect 9582 21926 9584 21978
rect 9528 21924 9584 21926
rect 9632 21978 9688 21980
rect 9632 21926 9634 21978
rect 9634 21926 9686 21978
rect 9686 21926 9688 21978
rect 9632 21924 9688 21926
rect 9736 21978 9792 21980
rect 9736 21926 9738 21978
rect 9738 21926 9790 21978
rect 9790 21926 9792 21978
rect 9736 21924 9792 21926
rect 8988 21756 9044 21812
rect 17844 21978 17900 21980
rect 17844 21926 17846 21978
rect 17846 21926 17898 21978
rect 17898 21926 17900 21978
rect 17844 21924 17900 21926
rect 17948 21978 18004 21980
rect 17948 21926 17950 21978
rect 17950 21926 18002 21978
rect 18002 21926 18004 21978
rect 17948 21924 18004 21926
rect 18052 21978 18108 21980
rect 18052 21926 18054 21978
rect 18054 21926 18106 21978
rect 18106 21926 18108 21978
rect 18052 21924 18108 21926
rect 11004 21810 11060 21812
rect 11004 21758 11006 21810
rect 11006 21758 11058 21810
rect 11058 21758 11060 21810
rect 11004 21756 11060 21758
rect 12908 21810 12964 21812
rect 12908 21758 12910 21810
rect 12910 21758 12962 21810
rect 12962 21758 12964 21810
rect 12908 21756 12964 21758
rect 23324 22092 23380 22148
rect 23772 22146 23828 22148
rect 23772 22094 23774 22146
rect 23774 22094 23826 22146
rect 23826 22094 23828 22146
rect 23772 22092 23828 22094
rect 17388 21810 17444 21812
rect 17388 21758 17390 21810
rect 17390 21758 17442 21810
rect 17442 21758 17444 21810
rect 17388 21756 17444 21758
rect 6076 21474 6132 21476
rect 6076 21422 6078 21474
rect 6078 21422 6130 21474
rect 6130 21422 6132 21474
rect 6076 21420 6132 21422
rect 6524 20076 6580 20132
rect 5740 18450 5796 18452
rect 5740 18398 5742 18450
rect 5742 18398 5794 18450
rect 5794 18398 5796 18450
rect 5740 18396 5796 18398
rect 5370 18058 5426 18060
rect 5370 18006 5372 18058
rect 5372 18006 5424 18058
rect 5424 18006 5426 18058
rect 5370 18004 5426 18006
rect 5474 18058 5530 18060
rect 5474 18006 5476 18058
rect 5476 18006 5528 18058
rect 5528 18006 5530 18058
rect 5474 18004 5530 18006
rect 5578 18058 5634 18060
rect 5578 18006 5580 18058
rect 5580 18006 5632 18058
rect 5632 18006 5634 18058
rect 5578 18004 5634 18006
rect 5516 16604 5572 16660
rect 5370 16490 5426 16492
rect 5370 16438 5372 16490
rect 5372 16438 5424 16490
rect 5424 16438 5426 16490
rect 5370 16436 5426 16438
rect 5474 16490 5530 16492
rect 5474 16438 5476 16490
rect 5476 16438 5528 16490
rect 5528 16438 5530 16490
rect 5474 16436 5530 16438
rect 5578 16490 5634 16492
rect 5578 16438 5580 16490
rect 5580 16438 5632 16490
rect 5632 16438 5634 16490
rect 5578 16436 5634 16438
rect 5852 15260 5908 15316
rect 5370 14922 5426 14924
rect 5370 14870 5372 14922
rect 5372 14870 5424 14922
rect 5424 14870 5426 14922
rect 5370 14868 5426 14870
rect 5474 14922 5530 14924
rect 5474 14870 5476 14922
rect 5476 14870 5528 14922
rect 5528 14870 5530 14922
rect 5474 14868 5530 14870
rect 5578 14922 5634 14924
rect 5578 14870 5580 14922
rect 5580 14870 5632 14922
rect 5632 14870 5634 14922
rect 5578 14868 5634 14870
rect 5516 14252 5572 14308
rect 8428 18338 8484 18340
rect 8428 18286 8430 18338
rect 8430 18286 8482 18338
rect 8482 18286 8484 18338
rect 8428 18284 8484 18286
rect 6524 17836 6580 17892
rect 8764 18620 8820 18676
rect 8652 16940 8708 16996
rect 6300 15874 6356 15876
rect 6300 15822 6302 15874
rect 6302 15822 6354 15874
rect 6354 15822 6356 15874
rect 6300 15820 6356 15822
rect 6412 15314 6468 15316
rect 6412 15262 6414 15314
rect 6414 15262 6466 15314
rect 6466 15262 6468 15314
rect 6412 15260 6468 15262
rect 6076 14530 6132 14532
rect 6076 14478 6078 14530
rect 6078 14478 6130 14530
rect 6130 14478 6132 14530
rect 6076 14476 6132 14478
rect 6524 14364 6580 14420
rect 6972 16882 7028 16884
rect 6972 16830 6974 16882
rect 6974 16830 7026 16882
rect 7026 16830 7028 16882
rect 6972 16828 7028 16830
rect 7980 16604 8036 16660
rect 7196 16044 7252 16100
rect 7532 15986 7588 15988
rect 7532 15934 7534 15986
rect 7534 15934 7586 15986
rect 7586 15934 7588 15986
rect 7532 15932 7588 15934
rect 7196 15820 7252 15876
rect 7308 15484 7364 15540
rect 7084 15372 7140 15428
rect 7644 15426 7700 15428
rect 7644 15374 7646 15426
rect 7646 15374 7698 15426
rect 7698 15374 7700 15426
rect 7644 15372 7700 15374
rect 7308 15314 7364 15316
rect 7308 15262 7310 15314
rect 7310 15262 7362 15314
rect 7362 15262 7364 15314
rect 7308 15260 7364 15262
rect 6636 14588 6692 14644
rect 6524 13970 6580 13972
rect 6524 13918 6526 13970
rect 6526 13918 6578 13970
rect 6578 13918 6580 13970
rect 6524 13916 6580 13918
rect 7420 13916 7476 13972
rect 7644 14306 7700 14308
rect 7644 14254 7646 14306
rect 7646 14254 7698 14306
rect 7698 14254 7700 14306
rect 7644 14252 7700 14254
rect 7532 14028 7588 14084
rect 8092 14642 8148 14644
rect 8092 14590 8094 14642
rect 8094 14590 8146 14642
rect 8146 14590 8148 14642
rect 8092 14588 8148 14590
rect 5370 13354 5426 13356
rect 5370 13302 5372 13354
rect 5372 13302 5424 13354
rect 5424 13302 5426 13354
rect 5370 13300 5426 13302
rect 5474 13354 5530 13356
rect 5474 13302 5476 13354
rect 5476 13302 5528 13354
rect 5528 13302 5530 13354
rect 5474 13300 5530 13302
rect 5578 13354 5634 13356
rect 5578 13302 5580 13354
rect 5580 13302 5632 13354
rect 5632 13302 5634 13354
rect 5578 13300 5634 13302
rect 5404 12796 5460 12852
rect 5852 12796 5908 12852
rect 7084 13634 7140 13636
rect 7084 13582 7086 13634
rect 7086 13582 7138 13634
rect 7138 13582 7140 13634
rect 7084 13580 7140 13582
rect 6076 12962 6132 12964
rect 6076 12910 6078 12962
rect 6078 12910 6130 12962
rect 6130 12910 6132 12962
rect 6076 12908 6132 12910
rect 5964 12290 6020 12292
rect 5964 12238 5966 12290
rect 5966 12238 6018 12290
rect 6018 12238 6020 12290
rect 5964 12236 6020 12238
rect 6300 12572 6356 12628
rect 6860 12572 6916 12628
rect 6188 12348 6244 12404
rect 6524 12290 6580 12292
rect 6524 12238 6526 12290
rect 6526 12238 6578 12290
rect 6578 12238 6580 12290
rect 6524 12236 6580 12238
rect 5370 11786 5426 11788
rect 5370 11734 5372 11786
rect 5372 11734 5424 11786
rect 5424 11734 5426 11786
rect 5370 11732 5426 11734
rect 5474 11786 5530 11788
rect 5474 11734 5476 11786
rect 5476 11734 5528 11786
rect 5528 11734 5530 11786
rect 5474 11732 5530 11734
rect 5578 11786 5634 11788
rect 5578 11734 5580 11786
rect 5580 11734 5632 11786
rect 5632 11734 5634 11786
rect 5578 11732 5634 11734
rect 8540 13916 8596 13972
rect 8316 13746 8372 13748
rect 8316 13694 8318 13746
rect 8318 13694 8370 13746
rect 8370 13694 8372 13746
rect 8316 13692 8372 13694
rect 8428 12684 8484 12740
rect 7308 12402 7364 12404
rect 7308 12350 7310 12402
rect 7310 12350 7362 12402
rect 7362 12350 7364 12402
rect 7308 12348 7364 12350
rect 7868 12402 7924 12404
rect 7868 12350 7870 12402
rect 7870 12350 7922 12402
rect 7922 12350 7924 12402
rect 7868 12348 7924 12350
rect 6860 12012 6916 12068
rect 7420 12012 7476 12068
rect 8316 12066 8372 12068
rect 8316 12014 8318 12066
rect 8318 12014 8370 12066
rect 8370 12014 8372 12066
rect 8316 12012 8372 12014
rect 5370 10218 5426 10220
rect 5370 10166 5372 10218
rect 5372 10166 5424 10218
rect 5424 10166 5426 10218
rect 5370 10164 5426 10166
rect 5474 10218 5530 10220
rect 5474 10166 5476 10218
rect 5476 10166 5528 10218
rect 5528 10166 5530 10218
rect 5474 10164 5530 10166
rect 5578 10218 5634 10220
rect 5578 10166 5580 10218
rect 5580 10166 5632 10218
rect 5632 10166 5634 10218
rect 5578 10164 5634 10166
rect 8316 9884 8372 9940
rect 6524 9772 6580 9828
rect 6524 9602 6580 9604
rect 6524 9550 6526 9602
rect 6526 9550 6578 9602
rect 6578 9550 6580 9602
rect 6524 9548 6580 9550
rect 5964 9266 6020 9268
rect 5964 9214 5966 9266
rect 5966 9214 6018 9266
rect 6018 9214 6020 9266
rect 5964 9212 6020 9214
rect 6524 9154 6580 9156
rect 6524 9102 6526 9154
rect 6526 9102 6578 9154
rect 6578 9102 6580 9154
rect 6524 9100 6580 9102
rect 5370 8650 5426 8652
rect 5370 8598 5372 8650
rect 5372 8598 5424 8650
rect 5424 8598 5426 8650
rect 5370 8596 5426 8598
rect 5474 8650 5530 8652
rect 5474 8598 5476 8650
rect 5476 8598 5528 8650
rect 5528 8598 5530 8650
rect 5474 8596 5530 8598
rect 5578 8650 5634 8652
rect 5578 8598 5580 8650
rect 5580 8598 5632 8650
rect 5632 8598 5634 8650
rect 5578 8596 5634 8598
rect 6076 8370 6132 8372
rect 6076 8318 6078 8370
rect 6078 8318 6130 8370
rect 6130 8318 6132 8370
rect 6076 8316 6132 8318
rect 5964 7586 6020 7588
rect 5964 7534 5966 7586
rect 5966 7534 6018 7586
rect 6018 7534 6020 7586
rect 5964 7532 6020 7534
rect 5852 7474 5908 7476
rect 5852 7422 5854 7474
rect 5854 7422 5906 7474
rect 5906 7422 5908 7474
rect 5852 7420 5908 7422
rect 5370 7082 5426 7084
rect 4172 5180 4228 5236
rect 5068 6972 5124 7028
rect 5370 7030 5372 7082
rect 5372 7030 5424 7082
rect 5424 7030 5426 7082
rect 5370 7028 5426 7030
rect 5474 7082 5530 7084
rect 5474 7030 5476 7082
rect 5476 7030 5528 7082
rect 5528 7030 5530 7082
rect 5474 7028 5530 7030
rect 5578 7082 5634 7084
rect 5578 7030 5580 7082
rect 5580 7030 5632 7082
rect 5632 7030 5634 7082
rect 5578 7028 5634 7030
rect 5628 6914 5684 6916
rect 5628 6862 5630 6914
rect 5630 6862 5682 6914
rect 5682 6862 5684 6914
rect 5628 6860 5684 6862
rect 5180 6412 5236 6468
rect 5740 6076 5796 6132
rect 5370 5514 5426 5516
rect 5370 5462 5372 5514
rect 5372 5462 5424 5514
rect 5424 5462 5426 5514
rect 5370 5460 5426 5462
rect 5474 5514 5530 5516
rect 5474 5462 5476 5514
rect 5476 5462 5528 5514
rect 5528 5462 5530 5514
rect 5474 5460 5530 5462
rect 5578 5514 5634 5516
rect 5578 5462 5580 5514
rect 5580 5462 5632 5514
rect 5632 5462 5634 5514
rect 5578 5460 5634 5462
rect 4732 5234 4788 5236
rect 4732 5182 4734 5234
rect 4734 5182 4786 5234
rect 4786 5182 4788 5234
rect 4732 5180 4788 5182
rect 5628 5068 5684 5124
rect 5180 4172 5236 4228
rect 5370 3946 5426 3948
rect 5370 3894 5372 3946
rect 5372 3894 5424 3946
rect 5424 3894 5426 3946
rect 5370 3892 5426 3894
rect 5474 3946 5530 3948
rect 5474 3894 5476 3946
rect 5476 3894 5528 3946
rect 5528 3894 5530 3946
rect 5474 3892 5530 3894
rect 5578 3946 5634 3948
rect 5578 3894 5580 3946
rect 5580 3894 5632 3946
rect 5632 3894 5634 3946
rect 5578 3892 5634 3894
rect 6636 7980 6692 8036
rect 7980 9826 8036 9828
rect 7980 9774 7982 9826
rect 7982 9774 8034 9826
rect 8034 9774 8036 9826
rect 7980 9772 8036 9774
rect 7196 9100 7252 9156
rect 7084 8876 7140 8932
rect 7756 8930 7812 8932
rect 7756 8878 7758 8930
rect 7758 8878 7810 8930
rect 7810 8878 7812 8930
rect 7756 8876 7812 8878
rect 7196 7586 7252 7588
rect 7196 7534 7198 7586
rect 7198 7534 7250 7586
rect 7250 7534 7252 7586
rect 7196 7532 7252 7534
rect 6972 7474 7028 7476
rect 6972 7422 6974 7474
rect 6974 7422 7026 7474
rect 7026 7422 7028 7474
rect 6972 7420 7028 7422
rect 6300 6802 6356 6804
rect 6300 6750 6302 6802
rect 6302 6750 6354 6802
rect 6354 6750 6356 6802
rect 6300 6748 6356 6750
rect 6412 6076 6468 6132
rect 7756 6690 7812 6692
rect 7756 6638 7758 6690
rect 7758 6638 7810 6690
rect 7810 6638 7812 6690
rect 7756 6636 7812 6638
rect 7420 6524 7476 6580
rect 6860 5964 6916 6020
rect 5964 5628 6020 5684
rect 6524 5906 6580 5908
rect 6524 5854 6526 5906
rect 6526 5854 6578 5906
rect 6578 5854 6580 5906
rect 6524 5852 6580 5854
rect 7196 5794 7252 5796
rect 7196 5742 7198 5794
rect 7198 5742 7250 5794
rect 7250 5742 7252 5794
rect 7196 5740 7252 5742
rect 6748 5234 6804 5236
rect 6748 5182 6750 5234
rect 6750 5182 6802 5234
rect 6802 5182 6804 5234
rect 6748 5180 6804 5182
rect 8316 8988 8372 9044
rect 8428 7308 8484 7364
rect 7980 6524 8036 6580
rect 8316 6636 8372 6692
rect 7420 5068 7476 5124
rect 7756 5292 7812 5348
rect 8540 6524 8596 6580
rect 8764 5740 8820 5796
rect 8540 4956 8596 5012
rect 9772 20860 9828 20916
rect 9996 20972 10052 21028
rect 9996 20802 10052 20804
rect 9996 20750 9998 20802
rect 9998 20750 10050 20802
rect 10050 20750 10052 20802
rect 9996 20748 10052 20750
rect 9528 20410 9584 20412
rect 9528 20358 9530 20410
rect 9530 20358 9582 20410
rect 9582 20358 9584 20410
rect 9528 20356 9584 20358
rect 9632 20410 9688 20412
rect 9632 20358 9634 20410
rect 9634 20358 9686 20410
rect 9686 20358 9688 20410
rect 9632 20356 9688 20358
rect 9736 20410 9792 20412
rect 9736 20358 9738 20410
rect 9738 20358 9790 20410
rect 9790 20358 9792 20410
rect 9736 20356 9792 20358
rect 9772 20130 9828 20132
rect 9772 20078 9774 20130
rect 9774 20078 9826 20130
rect 9826 20078 9828 20130
rect 9772 20076 9828 20078
rect 10444 19964 10500 20020
rect 9212 19122 9268 19124
rect 9212 19070 9214 19122
rect 9214 19070 9266 19122
rect 9266 19070 9268 19122
rect 9212 19068 9268 19070
rect 9212 18732 9268 18788
rect 9436 19122 9492 19124
rect 9436 19070 9438 19122
rect 9438 19070 9490 19122
rect 9490 19070 9492 19122
rect 9436 19068 9492 19070
rect 9528 18842 9584 18844
rect 9528 18790 9530 18842
rect 9530 18790 9582 18842
rect 9582 18790 9584 18842
rect 9528 18788 9584 18790
rect 9632 18842 9688 18844
rect 9632 18790 9634 18842
rect 9634 18790 9686 18842
rect 9686 18790 9688 18842
rect 9632 18788 9688 18790
rect 9736 18842 9792 18844
rect 9736 18790 9738 18842
rect 9738 18790 9790 18842
rect 9790 18790 9792 18842
rect 9736 18788 9792 18790
rect 9660 18674 9716 18676
rect 9660 18622 9662 18674
rect 9662 18622 9714 18674
rect 9714 18622 9716 18674
rect 9660 18620 9716 18622
rect 9100 18396 9156 18452
rect 8988 17836 9044 17892
rect 8988 17554 9044 17556
rect 8988 17502 8990 17554
rect 8990 17502 9042 17554
rect 9042 17502 9044 17554
rect 8988 17500 9044 17502
rect 9660 17554 9716 17556
rect 9660 17502 9662 17554
rect 9662 17502 9714 17554
rect 9714 17502 9716 17554
rect 9660 17500 9716 17502
rect 10556 20076 10612 20132
rect 10892 19964 10948 20020
rect 11228 20018 11284 20020
rect 11228 19966 11230 20018
rect 11230 19966 11282 20018
rect 11282 19966 11284 20018
rect 11228 19964 11284 19966
rect 12012 19964 12068 20020
rect 10892 19404 10948 19460
rect 12124 19852 12180 19908
rect 10892 18620 10948 18676
rect 11004 17666 11060 17668
rect 11004 17614 11006 17666
rect 11006 17614 11058 17666
rect 11058 17614 11060 17666
rect 11004 17612 11060 17614
rect 10108 17500 10164 17556
rect 9528 17274 9584 17276
rect 9528 17222 9530 17274
rect 9530 17222 9582 17274
rect 9582 17222 9584 17274
rect 9528 17220 9584 17222
rect 9632 17274 9688 17276
rect 9632 17222 9634 17274
rect 9634 17222 9686 17274
rect 9686 17222 9688 17274
rect 9632 17220 9688 17222
rect 9736 17274 9792 17276
rect 9736 17222 9738 17274
rect 9738 17222 9790 17274
rect 9790 17222 9792 17274
rect 9736 17220 9792 17222
rect 10668 16940 10724 16996
rect 9528 15706 9584 15708
rect 9528 15654 9530 15706
rect 9530 15654 9582 15706
rect 9582 15654 9584 15706
rect 9528 15652 9584 15654
rect 9632 15706 9688 15708
rect 9632 15654 9634 15706
rect 9634 15654 9686 15706
rect 9686 15654 9688 15706
rect 9632 15652 9688 15654
rect 9736 15706 9792 15708
rect 9736 15654 9738 15706
rect 9738 15654 9790 15706
rect 9790 15654 9792 15706
rect 9736 15652 9792 15654
rect 10780 16098 10836 16100
rect 10780 16046 10782 16098
rect 10782 16046 10834 16098
rect 10834 16046 10836 16098
rect 10780 16044 10836 16046
rect 10780 15874 10836 15876
rect 10780 15822 10782 15874
rect 10782 15822 10834 15874
rect 10834 15822 10836 15874
rect 10780 15820 10836 15822
rect 10444 14588 10500 14644
rect 9996 14252 10052 14308
rect 9528 14138 9584 14140
rect 9528 14086 9530 14138
rect 9530 14086 9582 14138
rect 9582 14086 9584 14138
rect 9528 14084 9584 14086
rect 9632 14138 9688 14140
rect 9632 14086 9634 14138
rect 9634 14086 9686 14138
rect 9686 14086 9688 14138
rect 9632 14084 9688 14086
rect 9736 14138 9792 14140
rect 9736 14086 9738 14138
rect 9738 14086 9790 14138
rect 9790 14086 9792 14138
rect 9736 14084 9792 14086
rect 11676 18396 11732 18452
rect 11788 17666 11844 17668
rect 11788 17614 11790 17666
rect 11790 17614 11842 17666
rect 11842 17614 11844 17666
rect 11788 17612 11844 17614
rect 11452 17500 11508 17556
rect 11452 17052 11508 17108
rect 11116 15372 11172 15428
rect 11228 15932 11284 15988
rect 11116 14588 11172 14644
rect 12348 17052 12404 17108
rect 12012 15932 12068 15988
rect 11452 15314 11508 15316
rect 11452 15262 11454 15314
rect 11454 15262 11506 15314
rect 11506 15262 11508 15314
rect 11452 15260 11508 15262
rect 9528 12570 9584 12572
rect 9528 12518 9530 12570
rect 9530 12518 9582 12570
rect 9582 12518 9584 12570
rect 9528 12516 9584 12518
rect 9632 12570 9688 12572
rect 9632 12518 9634 12570
rect 9634 12518 9686 12570
rect 9686 12518 9688 12570
rect 9632 12516 9688 12518
rect 9736 12570 9792 12572
rect 9736 12518 9738 12570
rect 9738 12518 9790 12570
rect 9790 12518 9792 12570
rect 9736 12516 9792 12518
rect 9996 12348 10052 12404
rect 9212 12124 9268 12180
rect 9548 12124 9604 12180
rect 9528 11002 9584 11004
rect 9528 10950 9530 11002
rect 9530 10950 9582 11002
rect 9582 10950 9584 11002
rect 9528 10948 9584 10950
rect 9632 11002 9688 11004
rect 9632 10950 9634 11002
rect 9634 10950 9686 11002
rect 9686 10950 9688 11002
rect 9632 10948 9688 10950
rect 9736 11002 9792 11004
rect 9736 10950 9738 11002
rect 9738 10950 9790 11002
rect 9790 10950 9792 11002
rect 9736 10948 9792 10950
rect 9528 9434 9584 9436
rect 9528 9382 9530 9434
rect 9530 9382 9582 9434
rect 9582 9382 9584 9434
rect 9528 9380 9584 9382
rect 9632 9434 9688 9436
rect 9632 9382 9634 9434
rect 9634 9382 9686 9434
rect 9686 9382 9688 9434
rect 9632 9380 9688 9382
rect 9736 9434 9792 9436
rect 9736 9382 9738 9434
rect 9738 9382 9790 9434
rect 9790 9382 9792 9434
rect 9736 9380 9792 9382
rect 9212 8316 9268 8372
rect 9528 7866 9584 7868
rect 9528 7814 9530 7866
rect 9530 7814 9582 7866
rect 9582 7814 9584 7866
rect 9528 7812 9584 7814
rect 9632 7866 9688 7868
rect 9632 7814 9634 7866
rect 9634 7814 9686 7866
rect 9686 7814 9688 7866
rect 9632 7812 9688 7814
rect 9736 7866 9792 7868
rect 9736 7814 9738 7866
rect 9738 7814 9790 7866
rect 9790 7814 9792 7866
rect 9736 7812 9792 7814
rect 11452 13580 11508 13636
rect 11676 13186 11732 13188
rect 11676 13134 11678 13186
rect 11678 13134 11730 13186
rect 11730 13134 11732 13186
rect 11676 13132 11732 13134
rect 12348 13634 12404 13636
rect 12348 13582 12350 13634
rect 12350 13582 12402 13634
rect 12402 13582 12404 13634
rect 12348 13580 12404 13582
rect 12460 13020 12516 13076
rect 11452 12290 11508 12292
rect 11452 12238 11454 12290
rect 11454 12238 11506 12290
rect 11506 12238 11508 12290
rect 11452 12236 11508 12238
rect 11228 11452 11284 11508
rect 11564 12178 11620 12180
rect 11564 12126 11566 12178
rect 11566 12126 11618 12178
rect 11618 12126 11620 12178
rect 11564 12124 11620 12126
rect 11340 11228 11396 11284
rect 12012 12012 12068 12068
rect 12236 12738 12292 12740
rect 12236 12686 12238 12738
rect 12238 12686 12290 12738
rect 12290 12686 12292 12738
rect 12236 12684 12292 12686
rect 12348 12178 12404 12180
rect 12348 12126 12350 12178
rect 12350 12126 12402 12178
rect 12402 12126 12404 12178
rect 12348 12124 12404 12126
rect 12124 11676 12180 11732
rect 11452 9212 11508 9268
rect 9528 6298 9584 6300
rect 9528 6246 9530 6298
rect 9530 6246 9582 6298
rect 9582 6246 9584 6298
rect 9528 6244 9584 6246
rect 9632 6298 9688 6300
rect 9632 6246 9634 6298
rect 9634 6246 9686 6298
rect 9686 6246 9688 6298
rect 9632 6244 9688 6246
rect 9736 6298 9792 6300
rect 9736 6246 9738 6298
rect 9738 6246 9790 6298
rect 9790 6246 9792 6298
rect 9736 6244 9792 6246
rect 9884 6188 9940 6244
rect 9660 6130 9716 6132
rect 9660 6078 9662 6130
rect 9662 6078 9714 6130
rect 9714 6078 9716 6130
rect 9660 6076 9716 6078
rect 9548 5682 9604 5684
rect 9548 5630 9550 5682
rect 9550 5630 9602 5682
rect 9602 5630 9604 5682
rect 9548 5628 9604 5630
rect 9528 4730 9584 4732
rect 9528 4678 9530 4730
rect 9530 4678 9582 4730
rect 9582 4678 9584 4730
rect 9528 4676 9584 4678
rect 9632 4730 9688 4732
rect 9632 4678 9634 4730
rect 9634 4678 9686 4730
rect 9686 4678 9688 4730
rect 9632 4676 9688 4678
rect 9736 4730 9792 4732
rect 9736 4678 9738 4730
rect 9738 4678 9790 4730
rect 9790 4678 9792 4730
rect 9736 4676 9792 4678
rect 10668 6466 10724 6468
rect 10668 6414 10670 6466
rect 10670 6414 10722 6466
rect 10722 6414 10724 6466
rect 10668 6412 10724 6414
rect 11228 8034 11284 8036
rect 11228 7982 11230 8034
rect 11230 7982 11282 8034
rect 11282 7982 11284 8034
rect 11228 7980 11284 7982
rect 11452 7532 11508 7588
rect 11116 6412 11172 6468
rect 10668 5964 10724 6020
rect 9884 4508 9940 4564
rect 9996 4844 10052 4900
rect 9100 4338 9156 4340
rect 9100 4286 9102 4338
rect 9102 4286 9154 4338
rect 9154 4286 9156 4338
rect 9100 4284 9156 4286
rect 10108 4620 10164 4676
rect 13686 21194 13742 21196
rect 13686 21142 13688 21194
rect 13688 21142 13740 21194
rect 13740 21142 13742 21194
rect 13686 21140 13742 21142
rect 13790 21194 13846 21196
rect 13790 21142 13792 21194
rect 13792 21142 13844 21194
rect 13844 21142 13846 21194
rect 13790 21140 13846 21142
rect 13894 21194 13950 21196
rect 13894 21142 13896 21194
rect 13896 21142 13948 21194
rect 13948 21142 13950 21194
rect 13894 21140 13950 21142
rect 14252 20748 14308 20804
rect 14812 20802 14868 20804
rect 14812 20750 14814 20802
rect 14814 20750 14866 20802
rect 14866 20750 14868 20802
rect 14812 20748 14868 20750
rect 14476 20690 14532 20692
rect 14476 20638 14478 20690
rect 14478 20638 14530 20690
rect 14530 20638 14532 20690
rect 14476 20636 14532 20638
rect 15260 20802 15316 20804
rect 15260 20750 15262 20802
rect 15262 20750 15314 20802
rect 15314 20750 15316 20802
rect 15260 20748 15316 20750
rect 15148 20690 15204 20692
rect 15148 20638 15150 20690
rect 15150 20638 15202 20690
rect 15202 20638 15204 20690
rect 15148 20636 15204 20638
rect 13244 20076 13300 20132
rect 13468 20130 13524 20132
rect 13468 20078 13470 20130
rect 13470 20078 13522 20130
rect 13522 20078 13524 20130
rect 13468 20076 13524 20078
rect 14252 19964 14308 20020
rect 13686 19626 13742 19628
rect 13686 19574 13688 19626
rect 13688 19574 13740 19626
rect 13740 19574 13742 19626
rect 13686 19572 13742 19574
rect 13790 19626 13846 19628
rect 13790 19574 13792 19626
rect 13792 19574 13844 19626
rect 13844 19574 13846 19626
rect 13790 19572 13846 19574
rect 13894 19626 13950 19628
rect 13894 19574 13896 19626
rect 13896 19574 13948 19626
rect 13948 19574 13950 19626
rect 13894 19572 13950 19574
rect 14252 19180 14308 19236
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 14476 18396 14532 18452
rect 13686 18058 13742 18060
rect 13686 18006 13688 18058
rect 13688 18006 13740 18058
rect 13740 18006 13742 18058
rect 13686 18004 13742 18006
rect 13790 18058 13846 18060
rect 13790 18006 13792 18058
rect 13792 18006 13844 18058
rect 13844 18006 13846 18058
rect 13790 18004 13846 18006
rect 13894 18058 13950 18060
rect 13894 18006 13896 18058
rect 13896 18006 13948 18058
rect 13948 18006 13950 18058
rect 13894 18004 13950 18006
rect 15036 20018 15092 20020
rect 15036 19966 15038 20018
rect 15038 19966 15090 20018
rect 15090 19966 15092 20018
rect 15036 19964 15092 19966
rect 14812 19906 14868 19908
rect 14812 19854 14814 19906
rect 14814 19854 14866 19906
rect 14866 19854 14868 19906
rect 14812 19852 14868 19854
rect 14812 19234 14868 19236
rect 14812 19182 14814 19234
rect 14814 19182 14866 19234
rect 14866 19182 14868 19234
rect 14812 19180 14868 19182
rect 16940 21362 16996 21364
rect 16940 21310 16942 21362
rect 16942 21310 16994 21362
rect 16994 21310 16996 21362
rect 16940 21308 16996 21310
rect 17948 21308 18004 21364
rect 17724 20972 17780 21028
rect 16940 20748 16996 20804
rect 17844 20410 17900 20412
rect 17844 20358 17846 20410
rect 17846 20358 17898 20410
rect 17898 20358 17900 20410
rect 17844 20356 17900 20358
rect 17948 20410 18004 20412
rect 17948 20358 17950 20410
rect 17950 20358 18002 20410
rect 18002 20358 18004 20410
rect 17948 20356 18004 20358
rect 18052 20410 18108 20412
rect 18052 20358 18054 20410
rect 18054 20358 18106 20410
rect 18106 20358 18108 20410
rect 18052 20356 18108 20358
rect 19292 21308 19348 21364
rect 19404 20636 19460 20692
rect 16156 20076 16212 20132
rect 17724 20076 17780 20132
rect 15372 19964 15428 20020
rect 15148 19180 15204 19236
rect 14588 17388 14644 17444
rect 16156 18956 16212 19012
rect 18508 19122 18564 19124
rect 18508 19070 18510 19122
rect 18510 19070 18562 19122
rect 18562 19070 18564 19122
rect 18508 19068 18564 19070
rect 17844 18842 17900 18844
rect 17844 18790 17846 18842
rect 17846 18790 17898 18842
rect 17898 18790 17900 18842
rect 17844 18788 17900 18790
rect 17948 18842 18004 18844
rect 17948 18790 17950 18842
rect 17950 18790 18002 18842
rect 18002 18790 18004 18842
rect 17948 18788 18004 18790
rect 18052 18842 18108 18844
rect 18052 18790 18054 18842
rect 18054 18790 18106 18842
rect 18106 18790 18108 18842
rect 18052 18788 18108 18790
rect 16156 17388 16212 17444
rect 13686 16490 13742 16492
rect 13686 16438 13688 16490
rect 13688 16438 13740 16490
rect 13740 16438 13742 16490
rect 13686 16436 13742 16438
rect 13790 16490 13846 16492
rect 13790 16438 13792 16490
rect 13792 16438 13844 16490
rect 13844 16438 13846 16490
rect 13790 16436 13846 16438
rect 13894 16490 13950 16492
rect 13894 16438 13896 16490
rect 13896 16438 13948 16490
rect 13948 16438 13950 16490
rect 13894 16436 13950 16438
rect 13580 15820 13636 15876
rect 14028 15148 14084 15204
rect 13356 15036 13412 15092
rect 13686 14922 13742 14924
rect 13686 14870 13688 14922
rect 13688 14870 13740 14922
rect 13740 14870 13742 14922
rect 13686 14868 13742 14870
rect 13790 14922 13846 14924
rect 13790 14870 13792 14922
rect 13792 14870 13844 14922
rect 13844 14870 13846 14922
rect 13790 14868 13846 14870
rect 13894 14922 13950 14924
rect 13894 14870 13896 14922
rect 13896 14870 13948 14922
rect 13948 14870 13950 14922
rect 13894 14868 13950 14870
rect 13686 13354 13742 13356
rect 13686 13302 13688 13354
rect 13688 13302 13740 13354
rect 13740 13302 13742 13354
rect 13686 13300 13742 13302
rect 13790 13354 13846 13356
rect 13790 13302 13792 13354
rect 13792 13302 13844 13354
rect 13844 13302 13846 13354
rect 13790 13300 13846 13302
rect 13894 13354 13950 13356
rect 13894 13302 13896 13354
rect 13896 13302 13948 13354
rect 13948 13302 13950 13354
rect 13894 13300 13950 13302
rect 13468 13132 13524 13188
rect 13916 12684 13972 12740
rect 15596 16828 15652 16884
rect 16044 16716 16100 16772
rect 14812 15148 14868 15204
rect 14924 16044 14980 16100
rect 17844 17274 17900 17276
rect 17844 17222 17846 17274
rect 17846 17222 17898 17274
rect 17898 17222 17900 17274
rect 17844 17220 17900 17222
rect 17948 17274 18004 17276
rect 17948 17222 17950 17274
rect 17950 17222 18002 17274
rect 18002 17222 18004 17274
rect 17948 17220 18004 17222
rect 18052 17274 18108 17276
rect 18052 17222 18054 17274
rect 18054 17222 18106 17274
rect 18106 17222 18108 17274
rect 18052 17220 18108 17222
rect 15596 15148 15652 15204
rect 14924 13020 14980 13076
rect 16156 15036 16212 15092
rect 15036 12908 15092 12964
rect 14812 12850 14868 12852
rect 14812 12798 14814 12850
rect 14814 12798 14866 12850
rect 14866 12798 14868 12850
rect 14812 12796 14868 12798
rect 14700 12684 14756 12740
rect 13468 12012 13524 12068
rect 12908 11676 12964 11732
rect 13686 11786 13742 11788
rect 13686 11734 13688 11786
rect 13688 11734 13740 11786
rect 13740 11734 13742 11786
rect 13686 11732 13742 11734
rect 13790 11786 13846 11788
rect 13790 11734 13792 11786
rect 13792 11734 13844 11786
rect 13844 11734 13846 11786
rect 13790 11732 13846 11734
rect 13894 11786 13950 11788
rect 13894 11734 13896 11786
rect 13896 11734 13948 11786
rect 13948 11734 13950 11786
rect 13894 11732 13950 11734
rect 12908 10668 12964 10724
rect 13686 10218 13742 10220
rect 13686 10166 13688 10218
rect 13688 10166 13740 10218
rect 13740 10166 13742 10218
rect 13686 10164 13742 10166
rect 13790 10218 13846 10220
rect 13790 10166 13792 10218
rect 13792 10166 13844 10218
rect 13844 10166 13846 10218
rect 13790 10164 13846 10166
rect 13894 10218 13950 10220
rect 13894 10166 13896 10218
rect 13896 10166 13948 10218
rect 13948 10166 13950 10218
rect 13894 10164 13950 10166
rect 14252 11900 14308 11956
rect 14476 11788 14532 11844
rect 14364 11228 14420 11284
rect 15036 11900 15092 11956
rect 15596 13468 15652 13524
rect 14924 11788 14980 11844
rect 14588 11282 14644 11284
rect 14588 11230 14590 11282
rect 14590 11230 14642 11282
rect 14642 11230 14644 11282
rect 14588 11228 14644 11230
rect 14812 11282 14868 11284
rect 14812 11230 14814 11282
rect 14814 11230 14866 11282
rect 14866 11230 14868 11282
rect 14812 11228 14868 11230
rect 14700 11170 14756 11172
rect 14700 11118 14702 11170
rect 14702 11118 14754 11170
rect 14754 11118 14756 11170
rect 14700 11116 14756 11118
rect 14364 10556 14420 10612
rect 12796 9772 12852 9828
rect 14252 9714 14308 9716
rect 14252 9662 14254 9714
rect 14254 9662 14306 9714
rect 14306 9662 14308 9714
rect 14252 9660 14308 9662
rect 14028 9602 14084 9604
rect 14028 9550 14030 9602
rect 14030 9550 14082 9602
rect 14082 9550 14084 9602
rect 14028 9548 14084 9550
rect 14364 8988 14420 9044
rect 12796 8876 12852 8932
rect 12124 7698 12180 7700
rect 12124 7646 12126 7698
rect 12126 7646 12178 7698
rect 12178 7646 12180 7698
rect 12124 7644 12180 7646
rect 12012 7586 12068 7588
rect 12012 7534 12014 7586
rect 12014 7534 12066 7586
rect 12066 7534 12068 7586
rect 12012 7532 12068 7534
rect 12236 6076 12292 6132
rect 11788 5852 11844 5908
rect 12460 8146 12516 8148
rect 12460 8094 12462 8146
rect 12462 8094 12514 8146
rect 12514 8094 12516 8146
rect 12460 8092 12516 8094
rect 13686 8650 13742 8652
rect 13686 8598 13688 8650
rect 13688 8598 13740 8650
rect 13740 8598 13742 8650
rect 13686 8596 13742 8598
rect 13790 8650 13846 8652
rect 13790 8598 13792 8650
rect 13792 8598 13844 8650
rect 13844 8598 13846 8650
rect 13790 8596 13846 8598
rect 13894 8650 13950 8652
rect 13894 8598 13896 8650
rect 13896 8598 13948 8650
rect 13948 8598 13950 8650
rect 13894 8596 13950 8598
rect 14028 8370 14084 8372
rect 14028 8318 14030 8370
rect 14030 8318 14082 8370
rect 14082 8318 14084 8370
rect 14028 8316 14084 8318
rect 12796 8146 12852 8148
rect 12796 8094 12798 8146
rect 12798 8094 12850 8146
rect 12850 8094 12852 8146
rect 12796 8092 12852 8094
rect 12908 8034 12964 8036
rect 12908 7982 12910 8034
rect 12910 7982 12962 8034
rect 12962 7982 12964 8034
rect 12908 7980 12964 7982
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 13020 7698 13076 7700
rect 13020 7646 13022 7698
rect 13022 7646 13074 7698
rect 13074 7646 13076 7698
rect 13020 7644 13076 7646
rect 12908 7532 12964 7588
rect 14476 8258 14532 8260
rect 14476 8206 14478 8258
rect 14478 8206 14530 8258
rect 14530 8206 14532 8258
rect 14476 8204 14532 8206
rect 15484 10834 15540 10836
rect 15484 10782 15486 10834
rect 15486 10782 15538 10834
rect 15538 10782 15540 10834
rect 15484 10780 15540 10782
rect 15372 10668 15428 10724
rect 15372 10108 15428 10164
rect 14812 9996 14868 10052
rect 14924 9826 14980 9828
rect 14924 9774 14926 9826
rect 14926 9774 14978 9826
rect 14978 9774 14980 9826
rect 14924 9772 14980 9774
rect 15260 9042 15316 9044
rect 15260 8990 15262 9042
rect 15262 8990 15314 9042
rect 15314 8990 15316 9042
rect 15260 8988 15316 8990
rect 15708 13020 15764 13076
rect 17844 15706 17900 15708
rect 17844 15654 17846 15706
rect 17846 15654 17898 15706
rect 17898 15654 17900 15706
rect 17844 15652 17900 15654
rect 17948 15706 18004 15708
rect 17948 15654 17950 15706
rect 17950 15654 18002 15706
rect 18002 15654 18004 15706
rect 17948 15652 18004 15654
rect 18052 15706 18108 15708
rect 18052 15654 18054 15706
rect 18054 15654 18106 15706
rect 18106 15654 18108 15706
rect 18052 15652 18108 15654
rect 19180 19234 19236 19236
rect 19180 19182 19182 19234
rect 19182 19182 19234 19234
rect 19234 19182 19236 19234
rect 19180 19180 19236 19182
rect 18956 19068 19012 19124
rect 19628 21474 19684 21476
rect 19628 21422 19630 21474
rect 19630 21422 19682 21474
rect 19682 21422 19684 21474
rect 19628 21420 19684 21422
rect 19740 20802 19796 20804
rect 19740 20750 19742 20802
rect 19742 20750 19794 20802
rect 19794 20750 19796 20802
rect 19740 20748 19796 20750
rect 19852 20188 19908 20244
rect 19516 19180 19572 19236
rect 20524 21474 20580 21476
rect 20524 21422 20526 21474
rect 20526 21422 20578 21474
rect 20578 21422 20580 21474
rect 20524 21420 20580 21422
rect 20300 20690 20356 20692
rect 20300 20638 20302 20690
rect 20302 20638 20354 20690
rect 20354 20638 20356 20690
rect 20300 20636 20356 20638
rect 20076 19964 20132 20020
rect 19404 19122 19460 19124
rect 19404 19070 19406 19122
rect 19406 19070 19458 19122
rect 19458 19070 19460 19122
rect 19404 19068 19460 19070
rect 19068 19010 19124 19012
rect 19068 18958 19070 19010
rect 19070 18958 19122 19010
rect 19122 18958 19124 19010
rect 19068 18956 19124 18958
rect 19516 17666 19572 17668
rect 19516 17614 19518 17666
rect 19518 17614 19570 17666
rect 19570 17614 19572 17666
rect 19516 17612 19572 17614
rect 22002 21194 22058 21196
rect 22002 21142 22004 21194
rect 22004 21142 22056 21194
rect 22056 21142 22058 21194
rect 22002 21140 22058 21142
rect 22106 21194 22162 21196
rect 22106 21142 22108 21194
rect 22108 21142 22160 21194
rect 22160 21142 22162 21194
rect 22106 21140 22162 21142
rect 22210 21194 22266 21196
rect 22210 21142 22212 21194
rect 22212 21142 22264 21194
rect 22264 21142 22266 21194
rect 22210 21140 22266 21142
rect 23100 20802 23156 20804
rect 23100 20750 23102 20802
rect 23102 20750 23154 20802
rect 23154 20750 23156 20802
rect 23100 20748 23156 20750
rect 20524 18396 20580 18452
rect 19292 17500 19348 17556
rect 18844 16940 18900 16996
rect 19628 17276 19684 17332
rect 18620 16882 18676 16884
rect 18620 16830 18622 16882
rect 18622 16830 18674 16882
rect 18674 16830 18676 16882
rect 18620 16828 18676 16830
rect 18508 15874 18564 15876
rect 18508 15822 18510 15874
rect 18510 15822 18562 15874
rect 18562 15822 18564 15874
rect 18508 15820 18564 15822
rect 18396 15484 18452 15540
rect 17724 15260 17780 15316
rect 20076 17612 20132 17668
rect 19740 16828 19796 16884
rect 18844 16770 18900 16772
rect 18844 16718 18846 16770
rect 18846 16718 18898 16770
rect 18898 16718 18900 16770
rect 18844 16716 18900 16718
rect 20076 16882 20132 16884
rect 20076 16830 20078 16882
rect 20078 16830 20130 16882
rect 20130 16830 20132 16882
rect 20076 16828 20132 16830
rect 22002 19626 22058 19628
rect 22002 19574 22004 19626
rect 22004 19574 22056 19626
rect 22056 19574 22058 19626
rect 22002 19572 22058 19574
rect 22106 19626 22162 19628
rect 22106 19574 22108 19626
rect 22108 19574 22160 19626
rect 22160 19574 22162 19626
rect 22106 19572 22162 19574
rect 22210 19626 22266 19628
rect 22210 19574 22212 19626
rect 22212 19574 22264 19626
rect 22264 19574 22266 19626
rect 22210 19572 22266 19574
rect 20636 16828 20692 16884
rect 20860 19404 20916 19460
rect 18956 16604 19012 16660
rect 18732 15820 18788 15876
rect 19404 15484 19460 15540
rect 18732 15260 18788 15316
rect 19852 15538 19908 15540
rect 19852 15486 19854 15538
rect 19854 15486 19906 15538
rect 19906 15486 19908 15538
rect 19852 15484 19908 15486
rect 20860 18396 20916 18452
rect 22002 18058 22058 18060
rect 22002 18006 22004 18058
rect 22004 18006 22056 18058
rect 22056 18006 22058 18058
rect 22002 18004 22058 18006
rect 22106 18058 22162 18060
rect 22106 18006 22108 18058
rect 22108 18006 22160 18058
rect 22160 18006 22162 18058
rect 22106 18004 22162 18006
rect 22210 18058 22266 18060
rect 22210 18006 22212 18058
rect 22212 18006 22264 18058
rect 22264 18006 22266 18058
rect 22210 18004 22266 18006
rect 24780 22092 24836 22148
rect 24668 21362 24724 21364
rect 24668 21310 24670 21362
rect 24670 21310 24722 21362
rect 24722 21310 24724 21362
rect 24668 21308 24724 21310
rect 24668 20188 24724 20244
rect 23884 19794 23940 19796
rect 23884 19742 23886 19794
rect 23886 19742 23938 19794
rect 23938 19742 23940 19794
rect 23884 19740 23940 19742
rect 23996 19404 24052 19460
rect 23884 19068 23940 19124
rect 25564 22594 25620 22596
rect 25564 22542 25566 22594
rect 25566 22542 25618 22594
rect 25618 22542 25620 22594
rect 25564 22540 25620 22542
rect 31612 24668 31668 24724
rect 30318 22762 30374 22764
rect 30318 22710 30320 22762
rect 30320 22710 30372 22762
rect 30372 22710 30374 22762
rect 30318 22708 30374 22710
rect 30422 22762 30478 22764
rect 30422 22710 30424 22762
rect 30424 22710 30476 22762
rect 30476 22710 30478 22762
rect 30422 22708 30478 22710
rect 30526 22762 30582 22764
rect 30526 22710 30528 22762
rect 30528 22710 30580 22762
rect 30580 22710 30582 22762
rect 30526 22708 30582 22710
rect 26908 22540 26964 22596
rect 28588 22594 28644 22596
rect 28588 22542 28590 22594
rect 28590 22542 28642 22594
rect 28642 22542 28644 22594
rect 28588 22540 28644 22542
rect 26572 22204 26628 22260
rect 26160 21978 26216 21980
rect 26160 21926 26162 21978
rect 26162 21926 26214 21978
rect 26214 21926 26216 21978
rect 26160 21924 26216 21926
rect 26264 21978 26320 21980
rect 26264 21926 26266 21978
rect 26266 21926 26318 21978
rect 26318 21926 26320 21978
rect 26264 21924 26320 21926
rect 26368 21978 26424 21980
rect 26368 21926 26370 21978
rect 26370 21926 26422 21978
rect 26422 21926 26424 21978
rect 26368 21924 26424 21926
rect 27468 22258 27524 22260
rect 27468 22206 27470 22258
rect 27470 22206 27522 22258
rect 27522 22206 27524 22258
rect 27468 22204 27524 22206
rect 25900 21586 25956 21588
rect 25900 21534 25902 21586
rect 25902 21534 25954 21586
rect 25954 21534 25956 21586
rect 25900 21532 25956 21534
rect 25676 21474 25732 21476
rect 25676 21422 25678 21474
rect 25678 21422 25730 21474
rect 25730 21422 25732 21474
rect 25676 21420 25732 21422
rect 25452 21308 25508 21364
rect 25228 20636 25284 20692
rect 25564 20748 25620 20804
rect 26124 20748 26180 20804
rect 24444 18450 24500 18452
rect 24444 18398 24446 18450
rect 24446 18398 24498 18450
rect 24498 18398 24500 18450
rect 24444 18396 24500 18398
rect 22988 16828 23044 16884
rect 22002 16490 22058 16492
rect 22002 16438 22004 16490
rect 22004 16438 22056 16490
rect 22056 16438 22058 16490
rect 22002 16436 22058 16438
rect 22106 16490 22162 16492
rect 22106 16438 22108 16490
rect 22108 16438 22160 16490
rect 22160 16438 22162 16490
rect 22106 16436 22162 16438
rect 22210 16490 22266 16492
rect 22210 16438 22212 16490
rect 22212 16438 22264 16490
rect 22264 16438 22266 16490
rect 22210 16436 22266 16438
rect 22204 16268 22260 16324
rect 20860 16044 20916 16100
rect 20636 15372 20692 15428
rect 17844 14138 17900 14140
rect 17844 14086 17846 14138
rect 17846 14086 17898 14138
rect 17898 14086 17900 14138
rect 17844 14084 17900 14086
rect 17948 14138 18004 14140
rect 17948 14086 17950 14138
rect 17950 14086 18002 14138
rect 18002 14086 18004 14138
rect 17948 14084 18004 14086
rect 18052 14138 18108 14140
rect 18052 14086 18054 14138
rect 18054 14086 18106 14138
rect 18106 14086 18108 14138
rect 18052 14084 18108 14086
rect 16492 13468 16548 13524
rect 16940 13522 16996 13524
rect 16940 13470 16942 13522
rect 16942 13470 16994 13522
rect 16994 13470 16996 13522
rect 16940 13468 16996 13470
rect 15820 12962 15876 12964
rect 15820 12910 15822 12962
rect 15822 12910 15874 12962
rect 15874 12910 15876 12962
rect 15820 12908 15876 12910
rect 16044 12850 16100 12852
rect 16044 12798 16046 12850
rect 16046 12798 16098 12850
rect 16098 12798 16100 12850
rect 16044 12796 16100 12798
rect 16604 12796 16660 12852
rect 16044 11228 16100 11284
rect 15820 11116 15876 11172
rect 16380 10722 16436 10724
rect 16380 10670 16382 10722
rect 16382 10670 16434 10722
rect 16434 10670 16436 10722
rect 16380 10668 16436 10670
rect 16044 10444 16100 10500
rect 17844 12570 17900 12572
rect 17844 12518 17846 12570
rect 17846 12518 17898 12570
rect 17898 12518 17900 12570
rect 17844 12516 17900 12518
rect 17948 12570 18004 12572
rect 17948 12518 17950 12570
rect 17950 12518 18002 12570
rect 18002 12518 18004 12570
rect 17948 12516 18004 12518
rect 18052 12570 18108 12572
rect 18052 12518 18054 12570
rect 18054 12518 18106 12570
rect 18106 12518 18108 12570
rect 18052 12516 18108 12518
rect 17388 12236 17444 12292
rect 16604 11116 16660 11172
rect 15372 8204 15428 8260
rect 15596 9548 15652 9604
rect 15596 8876 15652 8932
rect 16268 9714 16324 9716
rect 16268 9662 16270 9714
rect 16270 9662 16322 9714
rect 16322 9662 16324 9714
rect 16268 9660 16324 9662
rect 16604 9212 16660 9268
rect 16716 9660 16772 9716
rect 17612 11170 17668 11172
rect 17612 11118 17614 11170
rect 17614 11118 17666 11170
rect 17666 11118 17668 11170
rect 17612 11116 17668 11118
rect 17844 11002 17900 11004
rect 17844 10950 17846 11002
rect 17846 10950 17898 11002
rect 17898 10950 17900 11002
rect 17844 10948 17900 10950
rect 17948 11002 18004 11004
rect 17948 10950 17950 11002
rect 17950 10950 18002 11002
rect 18002 10950 18004 11002
rect 17948 10948 18004 10950
rect 18052 11002 18108 11004
rect 18052 10950 18054 11002
rect 18054 10950 18106 11002
rect 18106 10950 18108 11002
rect 18052 10948 18108 10950
rect 18172 10668 18228 10724
rect 18060 10610 18116 10612
rect 18060 10558 18062 10610
rect 18062 10558 18114 10610
rect 18114 10558 18116 10610
rect 18060 10556 18116 10558
rect 17388 10220 17444 10276
rect 18396 10498 18452 10500
rect 18396 10446 18398 10498
rect 18398 10446 18450 10498
rect 18450 10446 18452 10498
rect 18396 10444 18452 10446
rect 18172 10332 18228 10388
rect 17724 10050 17780 10052
rect 17724 9998 17726 10050
rect 17726 9998 17778 10050
rect 17778 9998 17780 10050
rect 17724 9996 17780 9998
rect 17948 9714 18004 9716
rect 17948 9662 17950 9714
rect 17950 9662 18002 9714
rect 18002 9662 18004 9714
rect 17948 9660 18004 9662
rect 17276 9548 17332 9604
rect 16492 9042 16548 9044
rect 16492 8990 16494 9042
rect 16494 8990 16546 9042
rect 16546 8990 16548 9042
rect 16492 8988 16548 8990
rect 13916 8034 13972 8036
rect 13916 7982 13918 8034
rect 13918 7982 13970 8034
rect 13970 7982 13972 8034
rect 13916 7980 13972 7982
rect 13804 7532 13860 7588
rect 13244 7474 13300 7476
rect 13244 7422 13246 7474
rect 13246 7422 13298 7474
rect 13298 7422 13300 7474
rect 13244 7420 13300 7422
rect 13132 7362 13188 7364
rect 13132 7310 13134 7362
rect 13134 7310 13186 7362
rect 13186 7310 13188 7362
rect 13132 7308 13188 7310
rect 12572 6860 12628 6916
rect 13686 7082 13742 7084
rect 13686 7030 13688 7082
rect 13688 7030 13740 7082
rect 13740 7030 13742 7082
rect 13686 7028 13742 7030
rect 13790 7082 13846 7084
rect 13790 7030 13792 7082
rect 13792 7030 13844 7082
rect 13844 7030 13846 7082
rect 13790 7028 13846 7030
rect 13894 7082 13950 7084
rect 13894 7030 13896 7082
rect 13896 7030 13948 7082
rect 13948 7030 13950 7082
rect 13894 7028 13950 7030
rect 13468 6860 13524 6916
rect 12684 6076 12740 6132
rect 13020 5964 13076 6020
rect 14140 7420 14196 7476
rect 15148 7420 15204 7476
rect 16380 6914 16436 6916
rect 16380 6862 16382 6914
rect 16382 6862 16434 6914
rect 16434 6862 16436 6914
rect 16380 6860 16436 6862
rect 15484 6524 15540 6580
rect 15260 6188 15316 6244
rect 14028 5964 14084 6020
rect 13244 5906 13300 5908
rect 13244 5854 13246 5906
rect 13246 5854 13298 5906
rect 13298 5854 13300 5906
rect 13244 5852 13300 5854
rect 12684 5794 12740 5796
rect 12684 5742 12686 5794
rect 12686 5742 12738 5794
rect 12738 5742 12740 5794
rect 12684 5740 12740 5742
rect 11564 4956 11620 5012
rect 10780 4562 10836 4564
rect 10780 4510 10782 4562
rect 10782 4510 10834 4562
rect 10834 4510 10836 4562
rect 10780 4508 10836 4510
rect 11004 4450 11060 4452
rect 11004 4398 11006 4450
rect 11006 4398 11058 4450
rect 11058 4398 11060 4450
rect 11004 4396 11060 4398
rect 12124 4450 12180 4452
rect 12124 4398 12126 4450
rect 12126 4398 12178 4450
rect 12178 4398 12180 4450
rect 12124 4396 12180 4398
rect 11116 4338 11172 4340
rect 11116 4286 11118 4338
rect 11118 4286 11170 4338
rect 11170 4286 11172 4338
rect 11116 4284 11172 4286
rect 11900 4338 11956 4340
rect 11900 4286 11902 4338
rect 11902 4286 11954 4338
rect 11954 4286 11956 4338
rect 11900 4284 11956 4286
rect 11564 4226 11620 4228
rect 11564 4174 11566 4226
rect 11566 4174 11618 4226
rect 11618 4174 11620 4226
rect 11564 4172 11620 4174
rect 8988 3612 9044 3668
rect 3388 1820 3444 1876
rect 5404 3388 5460 3444
rect 6636 3388 6692 3444
rect 10332 3666 10388 3668
rect 10332 3614 10334 3666
rect 10334 3614 10386 3666
rect 10386 3614 10388 3666
rect 10332 3612 10388 3614
rect 12572 3612 12628 3668
rect 9528 3162 9584 3164
rect 9528 3110 9530 3162
rect 9530 3110 9582 3162
rect 9582 3110 9584 3162
rect 9528 3108 9584 3110
rect 9632 3162 9688 3164
rect 9632 3110 9634 3162
rect 9634 3110 9686 3162
rect 9686 3110 9688 3162
rect 9632 3108 9688 3110
rect 9736 3162 9792 3164
rect 9736 3110 9738 3162
rect 9738 3110 9790 3162
rect 9790 3110 9792 3162
rect 9736 3108 9792 3110
rect 13916 5906 13972 5908
rect 13916 5854 13918 5906
rect 13918 5854 13970 5906
rect 13970 5854 13972 5906
rect 13916 5852 13972 5854
rect 14812 6076 14868 6132
rect 13686 5514 13742 5516
rect 13686 5462 13688 5514
rect 13688 5462 13740 5514
rect 13740 5462 13742 5514
rect 13686 5460 13742 5462
rect 13790 5514 13846 5516
rect 13790 5462 13792 5514
rect 13792 5462 13844 5514
rect 13844 5462 13846 5514
rect 13790 5460 13846 5462
rect 13894 5514 13950 5516
rect 13894 5462 13896 5514
rect 13896 5462 13948 5514
rect 13948 5462 13950 5514
rect 13894 5460 13950 5462
rect 15596 5964 15652 6020
rect 17500 9212 17556 9268
rect 17388 8930 17444 8932
rect 17388 8878 17390 8930
rect 17390 8878 17442 8930
rect 17442 8878 17444 8930
rect 17388 8876 17444 8878
rect 16716 8258 16772 8260
rect 16716 8206 16718 8258
rect 16718 8206 16770 8258
rect 16770 8206 16772 8258
rect 16716 8204 16772 8206
rect 17844 9434 17900 9436
rect 17844 9382 17846 9434
rect 17846 9382 17898 9434
rect 17898 9382 17900 9434
rect 17844 9380 17900 9382
rect 17948 9434 18004 9436
rect 17948 9382 17950 9434
rect 17950 9382 18002 9434
rect 18002 9382 18004 9434
rect 17948 9380 18004 9382
rect 18052 9434 18108 9436
rect 18052 9382 18054 9434
rect 18054 9382 18106 9434
rect 18106 9382 18108 9434
rect 18052 9380 18108 9382
rect 18284 9826 18340 9828
rect 18284 9774 18286 9826
rect 18286 9774 18338 9826
rect 18338 9774 18340 9826
rect 18284 9772 18340 9774
rect 17844 7866 17900 7868
rect 17844 7814 17846 7866
rect 17846 7814 17898 7866
rect 17898 7814 17900 7866
rect 17844 7812 17900 7814
rect 17948 7866 18004 7868
rect 17948 7814 17950 7866
rect 17950 7814 18002 7866
rect 18002 7814 18004 7866
rect 17948 7812 18004 7814
rect 18052 7866 18108 7868
rect 18052 7814 18054 7866
rect 18054 7814 18106 7866
rect 18106 7814 18108 7866
rect 18052 7812 18108 7814
rect 17388 7586 17444 7588
rect 17388 7534 17390 7586
rect 17390 7534 17442 7586
rect 17442 7534 17444 7586
rect 17388 7532 17444 7534
rect 17388 6860 17444 6916
rect 16604 6578 16660 6580
rect 16604 6526 16606 6578
rect 16606 6526 16658 6578
rect 16658 6526 16660 6578
rect 16604 6524 16660 6526
rect 15148 5292 15204 5348
rect 16044 5292 16100 5348
rect 16940 6412 16996 6468
rect 17844 6298 17900 6300
rect 17844 6246 17846 6298
rect 17846 6246 17898 6298
rect 17898 6246 17900 6298
rect 17844 6244 17900 6246
rect 17948 6298 18004 6300
rect 17948 6246 17950 6298
rect 17950 6246 18002 6298
rect 18002 6246 18004 6298
rect 17948 6244 18004 6246
rect 18052 6298 18108 6300
rect 18052 6246 18054 6298
rect 18054 6246 18106 6298
rect 18106 6246 18108 6298
rect 18052 6244 18108 6246
rect 16940 6076 16996 6132
rect 17724 6130 17780 6132
rect 17724 6078 17726 6130
rect 17726 6078 17778 6130
rect 17778 6078 17780 6130
rect 17724 6076 17780 6078
rect 16492 5964 16548 6020
rect 16716 5906 16772 5908
rect 16716 5854 16718 5906
rect 16718 5854 16770 5906
rect 16770 5854 16772 5906
rect 16716 5852 16772 5854
rect 16604 5292 16660 5348
rect 14028 4844 14084 4900
rect 16156 4844 16212 4900
rect 13692 4620 13748 4676
rect 13132 4396 13188 4452
rect 18620 13468 18676 13524
rect 19516 13468 19572 13524
rect 19404 12908 19460 12964
rect 19068 12738 19124 12740
rect 19068 12686 19070 12738
rect 19070 12686 19122 12738
rect 19122 12686 19124 12738
rect 19068 12684 19124 12686
rect 18956 12178 19012 12180
rect 18956 12126 18958 12178
rect 18958 12126 19010 12178
rect 19010 12126 19012 12178
rect 18956 12124 19012 12126
rect 18620 11564 18676 11620
rect 19740 12684 19796 12740
rect 19852 12572 19908 12628
rect 21420 16098 21476 16100
rect 21420 16046 21422 16098
rect 21422 16046 21474 16098
rect 21474 16046 21476 16098
rect 21420 16044 21476 16046
rect 21980 15986 22036 15988
rect 21980 15934 21982 15986
rect 21982 15934 22034 15986
rect 22034 15934 22036 15986
rect 21980 15932 22036 15934
rect 21644 15874 21700 15876
rect 21644 15822 21646 15874
rect 21646 15822 21698 15874
rect 21698 15822 21700 15874
rect 21644 15820 21700 15822
rect 22540 15874 22596 15876
rect 22540 15822 22542 15874
rect 22542 15822 22594 15874
rect 22594 15822 22596 15874
rect 22540 15820 22596 15822
rect 22428 15148 22484 15204
rect 22002 14922 22058 14924
rect 22002 14870 22004 14922
rect 22004 14870 22056 14922
rect 22056 14870 22058 14922
rect 22002 14868 22058 14870
rect 22106 14922 22162 14924
rect 22106 14870 22108 14922
rect 22108 14870 22160 14922
rect 22160 14870 22162 14922
rect 22106 14868 22162 14870
rect 22210 14922 22266 14924
rect 22210 14870 22212 14922
rect 22212 14870 22264 14922
rect 22264 14870 22266 14922
rect 22210 14868 22266 14870
rect 22652 15148 22708 15204
rect 23660 17276 23716 17332
rect 23660 16940 23716 16996
rect 23100 16268 23156 16324
rect 22988 15596 23044 15652
rect 23548 15596 23604 15652
rect 22876 14476 22932 14532
rect 23660 15036 23716 15092
rect 24220 15036 24276 15092
rect 23548 14530 23604 14532
rect 23548 14478 23550 14530
rect 23550 14478 23602 14530
rect 23602 14478 23604 14530
rect 23548 14476 23604 14478
rect 20412 14306 20468 14308
rect 20412 14254 20414 14306
rect 20414 14254 20466 14306
rect 20466 14254 20468 14306
rect 20412 14252 20468 14254
rect 23660 14418 23716 14420
rect 23660 14366 23662 14418
rect 23662 14366 23714 14418
rect 23714 14366 23716 14418
rect 23660 14364 23716 14366
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 22764 14306 22820 14308
rect 22764 14254 22766 14306
rect 22766 14254 22818 14306
rect 22818 14254 22820 14306
rect 22764 14252 22820 14254
rect 23436 14252 23492 14308
rect 20636 13804 20692 13860
rect 21084 13746 21140 13748
rect 21084 13694 21086 13746
rect 21086 13694 21138 13746
rect 21138 13694 21140 13746
rect 21084 13692 21140 13694
rect 19964 13580 20020 13636
rect 19628 11340 19684 11396
rect 19740 12012 19796 12068
rect 19180 11228 19236 11284
rect 18844 10220 18900 10276
rect 18620 9714 18676 9716
rect 18620 9662 18622 9714
rect 18622 9662 18674 9714
rect 18674 9662 18676 9714
rect 18620 9660 18676 9662
rect 19180 10108 19236 10164
rect 19068 9996 19124 10052
rect 19068 9772 19124 9828
rect 19180 9436 19236 9492
rect 19180 9042 19236 9044
rect 19180 8990 19182 9042
rect 19182 8990 19234 9042
rect 19234 8990 19236 9042
rect 19180 8988 19236 8990
rect 18956 7756 19012 7812
rect 19292 7644 19348 7700
rect 19516 7868 19572 7924
rect 19516 7532 19572 7588
rect 18956 6972 19012 7028
rect 18508 6076 18564 6132
rect 18172 6018 18228 6020
rect 18172 5966 18174 6018
rect 18174 5966 18226 6018
rect 18226 5966 18228 6018
rect 18172 5964 18228 5966
rect 18620 5964 18676 6020
rect 18620 5628 18676 5684
rect 18172 5292 18228 5348
rect 17844 4730 17900 4732
rect 17844 4678 17846 4730
rect 17846 4678 17898 4730
rect 17898 4678 17900 4730
rect 17844 4676 17900 4678
rect 17948 4730 18004 4732
rect 17948 4678 17950 4730
rect 17950 4678 18002 4730
rect 18002 4678 18004 4730
rect 17948 4676 18004 4678
rect 18052 4730 18108 4732
rect 18052 4678 18054 4730
rect 18054 4678 18106 4730
rect 18106 4678 18108 4730
rect 18052 4676 18108 4678
rect 19740 8034 19796 8036
rect 19740 7982 19742 8034
rect 19742 7982 19794 8034
rect 19794 7982 19796 8034
rect 19740 7980 19796 7982
rect 19740 6972 19796 7028
rect 19516 6412 19572 6468
rect 20524 13132 20580 13188
rect 21756 13746 21812 13748
rect 21756 13694 21758 13746
rect 21758 13694 21810 13746
rect 21810 13694 21812 13746
rect 21756 13692 21812 13694
rect 20188 12572 20244 12628
rect 21084 12178 21140 12180
rect 21084 12126 21086 12178
rect 21086 12126 21138 12178
rect 21138 12126 21140 12178
rect 21084 12124 21140 12126
rect 20188 12012 20244 12068
rect 20412 11788 20468 11844
rect 20076 11506 20132 11508
rect 20076 11454 20078 11506
rect 20078 11454 20130 11506
rect 20130 11454 20132 11506
rect 20076 11452 20132 11454
rect 20524 11394 20580 11396
rect 20524 11342 20526 11394
rect 20526 11342 20578 11394
rect 20578 11342 20580 11394
rect 20524 11340 20580 11342
rect 20300 10556 20356 10612
rect 20188 9772 20244 9828
rect 21420 11340 21476 11396
rect 21532 12684 21588 12740
rect 22204 13858 22260 13860
rect 22204 13806 22206 13858
rect 22206 13806 22258 13858
rect 22258 13806 22260 13858
rect 22204 13804 22260 13806
rect 22002 13354 22058 13356
rect 22002 13302 22004 13354
rect 22004 13302 22056 13354
rect 22056 13302 22058 13354
rect 22002 13300 22058 13302
rect 22106 13354 22162 13356
rect 22106 13302 22108 13354
rect 22108 13302 22160 13354
rect 22160 13302 22162 13354
rect 22106 13300 22162 13302
rect 22210 13354 22266 13356
rect 22210 13302 22212 13354
rect 22212 13302 22264 13354
rect 22264 13302 22266 13354
rect 22210 13300 22266 13302
rect 21868 13020 21924 13076
rect 23996 13244 24052 13300
rect 22092 12962 22148 12964
rect 22092 12910 22094 12962
rect 22094 12910 22146 12962
rect 22146 12910 22148 12962
rect 22092 12908 22148 12910
rect 23884 12962 23940 12964
rect 23884 12910 23886 12962
rect 23886 12910 23938 12962
rect 23938 12910 23940 12962
rect 23884 12908 23940 12910
rect 23660 12572 23716 12628
rect 23100 12348 23156 12404
rect 21532 11788 21588 11844
rect 21308 11228 21364 11284
rect 21420 11170 21476 11172
rect 21420 11118 21422 11170
rect 21422 11118 21474 11170
rect 21474 11118 21476 11170
rect 21420 11116 21476 11118
rect 21644 11900 21700 11956
rect 22002 11786 22058 11788
rect 22002 11734 22004 11786
rect 22004 11734 22056 11786
rect 22056 11734 22058 11786
rect 22002 11732 22058 11734
rect 22106 11786 22162 11788
rect 22106 11734 22108 11786
rect 22108 11734 22160 11786
rect 22160 11734 22162 11786
rect 22106 11732 22162 11734
rect 22210 11786 22266 11788
rect 22210 11734 22212 11786
rect 22212 11734 22264 11786
rect 22264 11734 22266 11786
rect 22210 11732 22266 11734
rect 22092 11564 22148 11620
rect 22540 11676 22596 11732
rect 20636 10498 20692 10500
rect 20636 10446 20638 10498
rect 20638 10446 20690 10498
rect 20690 10446 20692 10498
rect 20636 10444 20692 10446
rect 22316 10332 22372 10388
rect 22002 10218 22058 10220
rect 21308 10108 21364 10164
rect 22002 10166 22004 10218
rect 22004 10166 22056 10218
rect 22056 10166 22058 10218
rect 22002 10164 22058 10166
rect 22106 10218 22162 10220
rect 22106 10166 22108 10218
rect 22108 10166 22160 10218
rect 22160 10166 22162 10218
rect 22106 10164 22162 10166
rect 22210 10218 22266 10220
rect 22210 10166 22212 10218
rect 22212 10166 22264 10218
rect 22264 10166 22266 10218
rect 22210 10164 22266 10166
rect 20748 9826 20804 9828
rect 20748 9774 20750 9826
rect 20750 9774 20802 9826
rect 20802 9774 20804 9826
rect 20748 9772 20804 9774
rect 20524 9212 20580 9268
rect 20524 9042 20580 9044
rect 20524 8990 20526 9042
rect 20526 8990 20578 9042
rect 20578 8990 20580 9042
rect 20524 8988 20580 8990
rect 22540 10108 22596 10164
rect 21756 9996 21812 10052
rect 21756 9548 21812 9604
rect 20412 8876 20468 8932
rect 20300 8764 20356 8820
rect 21196 8764 21252 8820
rect 20300 8258 20356 8260
rect 20300 8206 20302 8258
rect 20302 8206 20354 8258
rect 20354 8206 20356 8258
rect 20300 8204 20356 8206
rect 20076 8092 20132 8148
rect 20636 8034 20692 8036
rect 20636 7982 20638 8034
rect 20638 7982 20690 8034
rect 20690 7982 20692 8034
rect 20636 7980 20692 7982
rect 21308 8092 21364 8148
rect 23996 12572 24052 12628
rect 22876 11676 22932 11732
rect 23100 11340 23156 11396
rect 22988 11282 23044 11284
rect 22988 11230 22990 11282
rect 22990 11230 23042 11282
rect 23042 11230 23044 11282
rect 22988 11228 23044 11230
rect 23100 10668 23156 10724
rect 22876 10108 22932 10164
rect 22764 9714 22820 9716
rect 22764 9662 22766 9714
rect 22766 9662 22818 9714
rect 22818 9662 22820 9714
rect 22764 9660 22820 9662
rect 23548 10556 23604 10612
rect 23884 11282 23940 11284
rect 23884 11230 23886 11282
rect 23886 11230 23938 11282
rect 23938 11230 23940 11282
rect 23884 11228 23940 11230
rect 23660 9772 23716 9828
rect 23884 9714 23940 9716
rect 23884 9662 23886 9714
rect 23886 9662 23938 9714
rect 23938 9662 23940 9714
rect 23884 9660 23940 9662
rect 23436 9436 23492 9492
rect 22876 8988 22932 9044
rect 22002 8650 22058 8652
rect 22002 8598 22004 8650
rect 22004 8598 22056 8650
rect 22056 8598 22058 8650
rect 22002 8596 22058 8598
rect 22106 8650 22162 8652
rect 22106 8598 22108 8650
rect 22108 8598 22160 8650
rect 22160 8598 22162 8650
rect 22106 8596 22162 8598
rect 22210 8650 22266 8652
rect 22210 8598 22212 8650
rect 22212 8598 22264 8650
rect 22264 8598 22266 8650
rect 22540 8652 22596 8708
rect 22210 8596 22266 8598
rect 24220 14364 24276 14420
rect 25340 19404 25396 19460
rect 26796 21586 26852 21588
rect 26796 21534 26798 21586
rect 26798 21534 26850 21586
rect 26850 21534 26852 21586
rect 26796 21532 26852 21534
rect 26796 20636 26852 20692
rect 26160 20410 26216 20412
rect 26160 20358 26162 20410
rect 26162 20358 26214 20410
rect 26214 20358 26216 20410
rect 26160 20356 26216 20358
rect 26264 20410 26320 20412
rect 26264 20358 26266 20410
rect 26266 20358 26318 20410
rect 26318 20358 26320 20410
rect 26264 20356 26320 20358
rect 26368 20410 26424 20412
rect 26368 20358 26370 20410
rect 26370 20358 26422 20410
rect 26422 20358 26424 20410
rect 26368 20356 26424 20358
rect 26572 20076 26628 20132
rect 25788 19740 25844 19796
rect 26160 18842 26216 18844
rect 26160 18790 26162 18842
rect 26162 18790 26214 18842
rect 26214 18790 26216 18842
rect 26160 18788 26216 18790
rect 26264 18842 26320 18844
rect 26264 18790 26266 18842
rect 26266 18790 26318 18842
rect 26318 18790 26320 18842
rect 26264 18788 26320 18790
rect 26368 18842 26424 18844
rect 26368 18790 26370 18842
rect 26370 18790 26422 18842
rect 26422 18790 26424 18842
rect 26368 18788 26424 18790
rect 25228 18396 25284 18452
rect 25564 18450 25620 18452
rect 25564 18398 25566 18450
rect 25566 18398 25618 18450
rect 25618 18398 25620 18450
rect 25564 18396 25620 18398
rect 26236 18450 26292 18452
rect 26236 18398 26238 18450
rect 26238 18398 26290 18450
rect 26290 18398 26292 18450
rect 26236 18396 26292 18398
rect 25788 18338 25844 18340
rect 25788 18286 25790 18338
rect 25790 18286 25842 18338
rect 25842 18286 25844 18338
rect 25788 18284 25844 18286
rect 27580 21308 27636 21364
rect 27132 20972 27188 21028
rect 27580 20914 27636 20916
rect 27580 20862 27582 20914
rect 27582 20862 27634 20914
rect 27634 20862 27636 20914
rect 27580 20860 27636 20862
rect 27804 20748 27860 20804
rect 27580 19458 27636 19460
rect 27580 19406 27582 19458
rect 27582 19406 27634 19458
rect 27634 19406 27636 19458
rect 27580 19404 27636 19406
rect 26460 18284 26516 18340
rect 25788 17500 25844 17556
rect 25900 17276 25956 17332
rect 26160 17274 26216 17276
rect 26160 17222 26162 17274
rect 26162 17222 26214 17274
rect 26214 17222 26216 17274
rect 26160 17220 26216 17222
rect 26264 17274 26320 17276
rect 26264 17222 26266 17274
rect 26266 17222 26318 17274
rect 26318 17222 26320 17274
rect 26264 17220 26320 17222
rect 26368 17274 26424 17276
rect 26368 17222 26370 17274
rect 26370 17222 26422 17274
rect 26422 17222 26424 17274
rect 26368 17220 26424 17222
rect 24332 10108 24388 10164
rect 24332 8930 24388 8932
rect 24332 8878 24334 8930
rect 24334 8878 24386 8930
rect 24386 8878 24388 8930
rect 24332 8876 24388 8878
rect 24220 8652 24276 8708
rect 21532 7474 21588 7476
rect 21532 7422 21534 7474
rect 21534 7422 21586 7474
rect 21586 7422 21588 7474
rect 21532 7420 21588 7422
rect 23548 8316 23604 8372
rect 22204 7474 22260 7476
rect 22204 7422 22206 7474
rect 22206 7422 22258 7474
rect 22258 7422 22260 7474
rect 22204 7420 22260 7422
rect 22092 7196 22148 7252
rect 22428 7196 22484 7252
rect 22002 7082 22058 7084
rect 22002 7030 22004 7082
rect 22004 7030 22056 7082
rect 22056 7030 22058 7082
rect 22002 7028 22058 7030
rect 22106 7082 22162 7084
rect 22106 7030 22108 7082
rect 22108 7030 22160 7082
rect 22160 7030 22162 7082
rect 22106 7028 22162 7030
rect 22210 7082 22266 7084
rect 22210 7030 22212 7082
rect 22212 7030 22264 7082
rect 22264 7030 22266 7082
rect 22210 7028 22266 7030
rect 19180 5292 19236 5348
rect 19964 5964 20020 6020
rect 19740 5682 19796 5684
rect 19740 5630 19742 5682
rect 19742 5630 19794 5682
rect 19794 5630 19796 5682
rect 19740 5628 19796 5630
rect 20188 5628 20244 5684
rect 20300 5852 20356 5908
rect 18956 4898 19012 4900
rect 18956 4846 18958 4898
rect 18958 4846 19010 4898
rect 19010 4846 19012 4898
rect 18956 4844 19012 4846
rect 19404 4562 19460 4564
rect 19404 4510 19406 4562
rect 19406 4510 19458 4562
rect 19458 4510 19460 4562
rect 19404 4508 19460 4510
rect 22002 5514 22058 5516
rect 22002 5462 22004 5514
rect 22004 5462 22056 5514
rect 22056 5462 22058 5514
rect 22002 5460 22058 5462
rect 22106 5514 22162 5516
rect 22106 5462 22108 5514
rect 22108 5462 22160 5514
rect 22160 5462 22162 5514
rect 22106 5460 22162 5462
rect 22210 5514 22266 5516
rect 22210 5462 22212 5514
rect 22212 5462 22264 5514
rect 22264 5462 22266 5514
rect 22210 5460 22266 5462
rect 20412 5180 20468 5236
rect 18396 4450 18452 4452
rect 18396 4398 18398 4450
rect 18398 4398 18450 4450
rect 18450 4398 18452 4450
rect 18396 4396 18452 4398
rect 22764 7308 22820 7364
rect 23212 6578 23268 6580
rect 23212 6526 23214 6578
rect 23214 6526 23266 6578
rect 23266 6526 23268 6578
rect 23212 6524 23268 6526
rect 13686 3946 13742 3948
rect 13686 3894 13688 3946
rect 13688 3894 13740 3946
rect 13740 3894 13742 3946
rect 13686 3892 13742 3894
rect 13790 3946 13846 3948
rect 13790 3894 13792 3946
rect 13792 3894 13844 3946
rect 13844 3894 13846 3946
rect 13790 3892 13846 3894
rect 13894 3946 13950 3948
rect 13894 3894 13896 3946
rect 13896 3894 13948 3946
rect 13948 3894 13950 3946
rect 13894 3892 13950 3894
rect 14140 3666 14196 3668
rect 14140 3614 14142 3666
rect 14142 3614 14194 3666
rect 14194 3614 14196 3666
rect 14140 3612 14196 3614
rect 19740 3612 19796 3668
rect 16156 3388 16212 3444
rect 18508 3442 18564 3444
rect 18508 3390 18510 3442
rect 18510 3390 18562 3442
rect 18562 3390 18564 3442
rect 18508 3388 18564 3390
rect 17844 3162 17900 3164
rect 17844 3110 17846 3162
rect 17846 3110 17898 3162
rect 17898 3110 17900 3162
rect 17844 3108 17900 3110
rect 17948 3162 18004 3164
rect 17948 3110 17950 3162
rect 17950 3110 18002 3162
rect 18002 3110 18004 3162
rect 17948 3108 18004 3110
rect 18052 3162 18108 3164
rect 18052 3110 18054 3162
rect 18054 3110 18106 3162
rect 18106 3110 18108 3162
rect 18052 3108 18108 3110
rect 21644 4338 21700 4340
rect 21644 4286 21646 4338
rect 21646 4286 21698 4338
rect 21698 4286 21700 4338
rect 21644 4284 21700 4286
rect 22652 4844 22708 4900
rect 24668 12850 24724 12852
rect 24668 12798 24670 12850
rect 24670 12798 24722 12850
rect 24722 12798 24724 12850
rect 24668 12796 24724 12798
rect 24556 12738 24612 12740
rect 24556 12686 24558 12738
rect 24558 12686 24610 12738
rect 24610 12686 24612 12738
rect 24556 12684 24612 12686
rect 27580 17612 27636 17668
rect 29372 21644 29428 21700
rect 29148 20972 29204 21028
rect 30318 21194 30374 21196
rect 30318 21142 30320 21194
rect 30320 21142 30372 21194
rect 30372 21142 30374 21194
rect 30318 21140 30374 21142
rect 30422 21194 30478 21196
rect 30422 21142 30424 21194
rect 30424 21142 30476 21194
rect 30476 21142 30478 21194
rect 30422 21140 30478 21142
rect 30526 21194 30582 21196
rect 30526 21142 30528 21194
rect 30528 21142 30580 21194
rect 30580 21142 30582 21194
rect 30526 21140 30582 21142
rect 30716 20860 30772 20916
rect 30380 20802 30436 20804
rect 30380 20750 30382 20802
rect 30382 20750 30434 20802
rect 30434 20750 30436 20802
rect 30380 20748 30436 20750
rect 29708 20690 29764 20692
rect 29708 20638 29710 20690
rect 29710 20638 29762 20690
rect 29762 20638 29764 20690
rect 29708 20636 29764 20638
rect 28476 20188 28532 20244
rect 29932 20524 29988 20580
rect 28924 20130 28980 20132
rect 28924 20078 28926 20130
rect 28926 20078 28978 20130
rect 28978 20078 28980 20130
rect 28924 20076 28980 20078
rect 28476 19964 28532 20020
rect 27916 19292 27972 19348
rect 28476 19068 28532 19124
rect 29820 19010 29876 19012
rect 29820 18958 29822 19010
rect 29822 18958 29874 19010
rect 29874 18958 29876 19010
rect 29820 18956 29876 18958
rect 29036 18396 29092 18452
rect 27916 17612 27972 17668
rect 27692 17052 27748 17108
rect 26684 16716 26740 16772
rect 27356 16770 27412 16772
rect 27356 16718 27358 16770
rect 27358 16718 27410 16770
rect 27410 16718 27412 16770
rect 27356 16716 27412 16718
rect 24556 12178 24612 12180
rect 24556 12126 24558 12178
rect 24558 12126 24610 12178
rect 24610 12126 24612 12178
rect 24556 12124 24612 12126
rect 28588 17442 28644 17444
rect 28588 17390 28590 17442
rect 28590 17390 28642 17442
rect 28642 17390 28644 17442
rect 28588 17388 28644 17390
rect 29372 18620 29428 18676
rect 30604 20578 30660 20580
rect 30604 20526 30606 20578
rect 30606 20526 30658 20578
rect 30658 20526 30660 20578
rect 30604 20524 30660 20526
rect 30716 20188 30772 20244
rect 30318 19626 30374 19628
rect 30318 19574 30320 19626
rect 30320 19574 30372 19626
rect 30372 19574 30374 19626
rect 30318 19572 30374 19574
rect 30422 19626 30478 19628
rect 30422 19574 30424 19626
rect 30424 19574 30476 19626
rect 30476 19574 30478 19626
rect 30422 19572 30478 19574
rect 30526 19626 30582 19628
rect 30526 19574 30528 19626
rect 30528 19574 30580 19626
rect 30580 19574 30582 19626
rect 30526 19572 30582 19574
rect 29260 18172 29316 18228
rect 29148 17442 29204 17444
rect 29148 17390 29150 17442
rect 29150 17390 29202 17442
rect 29202 17390 29204 17442
rect 29148 17388 29204 17390
rect 29036 17276 29092 17332
rect 30318 18058 30374 18060
rect 30318 18006 30320 18058
rect 30320 18006 30372 18058
rect 30372 18006 30374 18058
rect 30318 18004 30374 18006
rect 30422 18058 30478 18060
rect 30422 18006 30424 18058
rect 30424 18006 30476 18058
rect 30476 18006 30478 18058
rect 30422 18004 30478 18006
rect 30526 18058 30582 18060
rect 30526 18006 30528 18058
rect 30528 18006 30580 18058
rect 30580 18006 30582 18058
rect 30526 18004 30582 18006
rect 28700 16994 28756 16996
rect 28700 16942 28702 16994
rect 28702 16942 28754 16994
rect 28754 16942 28756 16994
rect 28700 16940 28756 16942
rect 29260 16940 29316 16996
rect 28476 16828 28532 16884
rect 25564 16044 25620 16100
rect 26124 16044 26180 16100
rect 26908 16098 26964 16100
rect 26908 16046 26910 16098
rect 26910 16046 26962 16098
rect 26962 16046 26964 16098
rect 26908 16044 26964 16046
rect 26160 15706 26216 15708
rect 26160 15654 26162 15706
rect 26162 15654 26214 15706
rect 26214 15654 26216 15706
rect 26160 15652 26216 15654
rect 26264 15706 26320 15708
rect 26264 15654 26266 15706
rect 26266 15654 26318 15706
rect 26318 15654 26320 15706
rect 26264 15652 26320 15654
rect 26368 15706 26424 15708
rect 26368 15654 26370 15706
rect 26370 15654 26422 15706
rect 26422 15654 26424 15706
rect 26368 15652 26424 15654
rect 26684 15148 26740 15204
rect 26796 14418 26852 14420
rect 26796 14366 26798 14418
rect 26798 14366 26850 14418
rect 26850 14366 26852 14418
rect 26796 14364 26852 14366
rect 26160 14138 26216 14140
rect 26160 14086 26162 14138
rect 26162 14086 26214 14138
rect 26214 14086 26216 14138
rect 26160 14084 26216 14086
rect 26264 14138 26320 14140
rect 26264 14086 26266 14138
rect 26266 14086 26318 14138
rect 26318 14086 26320 14138
rect 26264 14084 26320 14086
rect 26368 14138 26424 14140
rect 26368 14086 26370 14138
rect 26370 14086 26422 14138
rect 26422 14086 26424 14138
rect 26368 14084 26424 14086
rect 25004 11506 25060 11508
rect 25004 11454 25006 11506
rect 25006 11454 25058 11506
rect 25058 11454 25060 11506
rect 25004 11452 25060 11454
rect 24556 11228 24612 11284
rect 24556 10722 24612 10724
rect 24556 10670 24558 10722
rect 24558 10670 24610 10722
rect 24610 10670 24612 10722
rect 24556 10668 24612 10670
rect 25564 10722 25620 10724
rect 25564 10670 25566 10722
rect 25566 10670 25618 10722
rect 25618 10670 25620 10722
rect 25564 10668 25620 10670
rect 24668 10556 24724 10612
rect 25228 10444 25284 10500
rect 25564 9884 25620 9940
rect 25116 9714 25172 9716
rect 25116 9662 25118 9714
rect 25118 9662 25170 9714
rect 25170 9662 25172 9714
rect 25116 9660 25172 9662
rect 24556 9042 24612 9044
rect 24556 8990 24558 9042
rect 24558 8990 24610 9042
rect 24610 8990 24612 9042
rect 24556 8988 24612 8990
rect 27132 12796 27188 12852
rect 26160 12570 26216 12572
rect 26160 12518 26162 12570
rect 26162 12518 26214 12570
rect 26214 12518 26216 12570
rect 26160 12516 26216 12518
rect 26264 12570 26320 12572
rect 26264 12518 26266 12570
rect 26266 12518 26318 12570
rect 26318 12518 26320 12570
rect 26264 12516 26320 12518
rect 26368 12570 26424 12572
rect 26368 12518 26370 12570
rect 26370 12518 26422 12570
rect 26422 12518 26424 12570
rect 26368 12516 26424 12518
rect 26908 12178 26964 12180
rect 26908 12126 26910 12178
rect 26910 12126 26962 12178
rect 26962 12126 26964 12178
rect 26908 12124 26964 12126
rect 26124 11676 26180 11732
rect 26684 11394 26740 11396
rect 26684 11342 26686 11394
rect 26686 11342 26738 11394
rect 26738 11342 26740 11394
rect 26684 11340 26740 11342
rect 25900 11116 25956 11172
rect 26160 11002 26216 11004
rect 26160 10950 26162 11002
rect 26162 10950 26214 11002
rect 26214 10950 26216 11002
rect 26160 10948 26216 10950
rect 26264 11002 26320 11004
rect 26264 10950 26266 11002
rect 26266 10950 26318 11002
rect 26318 10950 26320 11002
rect 26264 10948 26320 10950
rect 26368 11002 26424 11004
rect 26368 10950 26370 11002
rect 26370 10950 26422 11002
rect 26422 10950 26424 11002
rect 26368 10948 26424 10950
rect 26012 10498 26068 10500
rect 26012 10446 26014 10498
rect 26014 10446 26066 10498
rect 26066 10446 26068 10498
rect 26012 10444 26068 10446
rect 26460 9884 26516 9940
rect 26348 9826 26404 9828
rect 26348 9774 26350 9826
rect 26350 9774 26402 9826
rect 26402 9774 26404 9826
rect 26348 9772 26404 9774
rect 26160 9434 26216 9436
rect 26160 9382 26162 9434
rect 26162 9382 26214 9434
rect 26214 9382 26216 9434
rect 26160 9380 26216 9382
rect 26264 9434 26320 9436
rect 26264 9382 26266 9434
rect 26266 9382 26318 9434
rect 26318 9382 26320 9434
rect 26264 9380 26320 9382
rect 26368 9434 26424 9436
rect 26368 9382 26370 9434
rect 26370 9382 26422 9434
rect 26422 9382 26424 9434
rect 26368 9380 26424 9382
rect 25900 9100 25956 9156
rect 25788 8930 25844 8932
rect 25788 8878 25790 8930
rect 25790 8878 25842 8930
rect 25842 8878 25844 8930
rect 25788 8876 25844 8878
rect 26460 8818 26516 8820
rect 26460 8766 26462 8818
rect 26462 8766 26514 8818
rect 26514 8766 26516 8818
rect 26460 8764 26516 8766
rect 27020 10668 27076 10724
rect 28924 16044 28980 16100
rect 27468 15538 27524 15540
rect 27468 15486 27470 15538
rect 27470 15486 27522 15538
rect 27522 15486 27524 15538
rect 27468 15484 27524 15486
rect 28140 15874 28196 15876
rect 28140 15822 28142 15874
rect 28142 15822 28194 15874
rect 28194 15822 28196 15874
rect 28140 15820 28196 15822
rect 27804 15484 27860 15540
rect 28700 15596 28756 15652
rect 29484 17612 29540 17668
rect 30268 17666 30324 17668
rect 30268 17614 30270 17666
rect 30270 17614 30322 17666
rect 30322 17614 30324 17666
rect 30268 17612 30324 17614
rect 29372 16098 29428 16100
rect 29372 16046 29374 16098
rect 29374 16046 29426 16098
rect 29426 16046 29428 16098
rect 29372 16044 29428 16046
rect 29148 15820 29204 15876
rect 28924 15148 28980 15204
rect 28700 15036 28756 15092
rect 27580 14306 27636 14308
rect 27580 14254 27582 14306
rect 27582 14254 27634 14306
rect 27634 14254 27636 14306
rect 27580 14252 27636 14254
rect 27468 13970 27524 13972
rect 27468 13918 27470 13970
rect 27470 13918 27522 13970
rect 27522 13918 27524 13970
rect 27468 13916 27524 13918
rect 27804 13804 27860 13860
rect 28588 13858 28644 13860
rect 28588 13806 28590 13858
rect 28590 13806 28642 13858
rect 28642 13806 28644 13858
rect 28588 13804 28644 13806
rect 27580 11394 27636 11396
rect 27580 11342 27582 11394
rect 27582 11342 27634 11394
rect 27634 11342 27636 11394
rect 27580 11340 27636 11342
rect 27916 10780 27972 10836
rect 28028 10668 28084 10724
rect 28924 14588 28980 14644
rect 29260 15932 29316 15988
rect 29932 17276 29988 17332
rect 29596 16994 29652 16996
rect 29596 16942 29598 16994
rect 29598 16942 29650 16994
rect 29650 16942 29652 16994
rect 29596 16940 29652 16942
rect 30604 16940 30660 16996
rect 30318 16490 30374 16492
rect 30318 16438 30320 16490
rect 30320 16438 30372 16490
rect 30372 16438 30374 16490
rect 30318 16436 30374 16438
rect 30422 16490 30478 16492
rect 30422 16438 30424 16490
rect 30424 16438 30476 16490
rect 30476 16438 30478 16490
rect 30422 16436 30478 16438
rect 30526 16490 30582 16492
rect 30526 16438 30528 16490
rect 30528 16438 30580 16490
rect 30580 16438 30582 16490
rect 30526 16436 30582 16438
rect 30044 16268 30100 16324
rect 29708 15986 29764 15988
rect 29708 15934 29710 15986
rect 29710 15934 29762 15986
rect 29762 15934 29764 15986
rect 29708 15932 29764 15934
rect 30156 15932 30212 15988
rect 29932 15596 29988 15652
rect 29484 14588 29540 14644
rect 29260 13244 29316 13300
rect 29260 12908 29316 12964
rect 29596 13132 29652 13188
rect 28700 11676 28756 11732
rect 30604 15986 30660 15988
rect 30604 15934 30606 15986
rect 30606 15934 30658 15986
rect 30658 15934 30660 15986
rect 30604 15932 30660 15934
rect 30828 19180 30884 19236
rect 31164 21532 31220 21588
rect 31052 21474 31108 21476
rect 31052 21422 31054 21474
rect 31054 21422 31106 21474
rect 31106 21422 31108 21474
rect 31052 21420 31108 21422
rect 30828 17724 30884 17780
rect 31052 21084 31108 21140
rect 31612 21084 31668 21140
rect 31276 20748 31332 20804
rect 31164 18620 31220 18676
rect 33628 21308 33684 21364
rect 34476 21978 34532 21980
rect 34476 21926 34478 21978
rect 34478 21926 34530 21978
rect 34530 21926 34532 21978
rect 34476 21924 34532 21926
rect 34580 21978 34636 21980
rect 34580 21926 34582 21978
rect 34582 21926 34634 21978
rect 34634 21926 34636 21978
rect 34580 21924 34636 21926
rect 34684 21978 34740 21980
rect 34684 21926 34686 21978
rect 34686 21926 34738 21978
rect 34738 21926 34740 21978
rect 34684 21924 34740 21926
rect 31836 20188 31892 20244
rect 31388 18956 31444 19012
rect 31836 18396 31892 18452
rect 31388 17442 31444 17444
rect 31388 17390 31390 17442
rect 31390 17390 31442 17442
rect 31442 17390 31444 17442
rect 31388 17388 31444 17390
rect 33180 19234 33236 19236
rect 33180 19182 33182 19234
rect 33182 19182 33234 19234
rect 33234 19182 33236 19234
rect 33180 19180 33236 19182
rect 33964 19404 34020 19460
rect 33852 19292 33908 19348
rect 33292 19068 33348 19124
rect 32956 19010 33012 19012
rect 32956 18958 32958 19010
rect 32958 18958 33010 19010
rect 33010 18958 33012 19010
rect 32956 18956 33012 18958
rect 33740 19180 33796 19236
rect 33852 18844 33908 18900
rect 34476 20410 34532 20412
rect 34476 20358 34478 20410
rect 34478 20358 34530 20410
rect 34530 20358 34532 20410
rect 34476 20356 34532 20358
rect 34580 20410 34636 20412
rect 34580 20358 34582 20410
rect 34582 20358 34634 20410
rect 34634 20358 34636 20410
rect 34580 20356 34636 20358
rect 34684 20410 34740 20412
rect 34684 20358 34686 20410
rect 34686 20358 34738 20410
rect 34738 20358 34740 20410
rect 34684 20356 34740 20358
rect 34076 18956 34132 19012
rect 33068 18226 33124 18228
rect 33068 18174 33070 18226
rect 33070 18174 33122 18226
rect 33122 18174 33124 18226
rect 33068 18172 33124 18174
rect 32060 17052 32116 17108
rect 31724 16940 31780 16996
rect 31612 16882 31668 16884
rect 31612 16830 31614 16882
rect 31614 16830 31666 16882
rect 31666 16830 31668 16882
rect 31612 16828 31668 16830
rect 31612 15148 31668 15204
rect 30318 14922 30374 14924
rect 30318 14870 30320 14922
rect 30320 14870 30372 14922
rect 30372 14870 30374 14922
rect 30318 14868 30374 14870
rect 30422 14922 30478 14924
rect 30422 14870 30424 14922
rect 30424 14870 30476 14922
rect 30476 14870 30478 14922
rect 30422 14868 30478 14870
rect 30526 14922 30582 14924
rect 30526 14870 30528 14922
rect 30528 14870 30580 14922
rect 30580 14870 30582 14922
rect 30526 14868 30582 14870
rect 31388 14364 31444 14420
rect 30716 13468 30772 13524
rect 30318 13354 30374 13356
rect 30318 13302 30320 13354
rect 30320 13302 30372 13354
rect 30372 13302 30374 13354
rect 30318 13300 30374 13302
rect 30422 13354 30478 13356
rect 30422 13302 30424 13354
rect 30424 13302 30476 13354
rect 30476 13302 30478 13354
rect 30422 13300 30478 13302
rect 30526 13354 30582 13356
rect 30526 13302 30528 13354
rect 30528 13302 30580 13354
rect 30580 13302 30582 13354
rect 30526 13300 30582 13302
rect 30318 11786 30374 11788
rect 30318 11734 30320 11786
rect 30320 11734 30372 11786
rect 30372 11734 30374 11786
rect 30318 11732 30374 11734
rect 30422 11786 30478 11788
rect 30422 11734 30424 11786
rect 30424 11734 30476 11786
rect 30476 11734 30478 11786
rect 30422 11732 30478 11734
rect 30526 11786 30582 11788
rect 30526 11734 30528 11786
rect 30528 11734 30580 11786
rect 30580 11734 30582 11786
rect 30526 11732 30582 11734
rect 29596 11676 29652 11732
rect 29484 11564 29540 11620
rect 29820 11506 29876 11508
rect 29820 11454 29822 11506
rect 29822 11454 29874 11506
rect 29874 11454 29876 11506
rect 29820 11452 29876 11454
rect 30828 11452 30884 11508
rect 28476 10892 28532 10948
rect 26572 8428 26628 8484
rect 25788 8370 25844 8372
rect 25788 8318 25790 8370
rect 25790 8318 25842 8370
rect 25842 8318 25844 8370
rect 25788 8316 25844 8318
rect 26908 9772 26964 9828
rect 24668 8204 24724 8260
rect 25900 8258 25956 8260
rect 25900 8206 25902 8258
rect 25902 8206 25954 8258
rect 25954 8206 25956 8258
rect 25900 8204 25956 8206
rect 25788 8092 25844 8148
rect 24780 7868 24836 7924
rect 24780 7420 24836 7476
rect 26236 8034 26292 8036
rect 26236 7982 26238 8034
rect 26238 7982 26290 8034
rect 26290 7982 26292 8034
rect 26236 7980 26292 7982
rect 26460 7980 26516 8036
rect 26160 7866 26216 7868
rect 26160 7814 26162 7866
rect 26162 7814 26214 7866
rect 26214 7814 26216 7866
rect 26160 7812 26216 7814
rect 26264 7866 26320 7868
rect 26264 7814 26266 7866
rect 26266 7814 26318 7866
rect 26318 7814 26320 7866
rect 26264 7812 26320 7814
rect 26368 7866 26424 7868
rect 26368 7814 26370 7866
rect 26370 7814 26422 7866
rect 26422 7814 26424 7866
rect 26368 7812 26424 7814
rect 26572 7586 26628 7588
rect 26572 7534 26574 7586
rect 26574 7534 26626 7586
rect 26626 7534 26628 7586
rect 26572 7532 26628 7534
rect 24444 5852 24500 5908
rect 25228 7084 25284 7140
rect 26124 7084 26180 7140
rect 26572 6578 26628 6580
rect 26572 6526 26574 6578
rect 26574 6526 26626 6578
rect 26626 6526 26628 6578
rect 26572 6524 26628 6526
rect 26160 6298 26216 6300
rect 26160 6246 26162 6298
rect 26162 6246 26214 6298
rect 26214 6246 26216 6298
rect 26160 6244 26216 6246
rect 26264 6298 26320 6300
rect 26264 6246 26266 6298
rect 26266 6246 26318 6298
rect 26318 6246 26320 6298
rect 26264 6244 26320 6246
rect 26368 6298 26424 6300
rect 26368 6246 26370 6298
rect 26370 6246 26422 6298
rect 26422 6246 26424 6298
rect 26368 6244 26424 6246
rect 27244 9154 27300 9156
rect 27244 9102 27246 9154
rect 27246 9102 27298 9154
rect 27298 9102 27300 9154
rect 27244 9100 27300 9102
rect 26908 8428 26964 8484
rect 28252 10556 28308 10612
rect 30380 10610 30436 10612
rect 30380 10558 30382 10610
rect 30382 10558 30434 10610
rect 30434 10558 30436 10610
rect 30380 10556 30436 10558
rect 30318 10218 30374 10220
rect 30318 10166 30320 10218
rect 30320 10166 30372 10218
rect 30372 10166 30374 10218
rect 30318 10164 30374 10166
rect 30422 10218 30478 10220
rect 30422 10166 30424 10218
rect 30424 10166 30476 10218
rect 30476 10166 30478 10218
rect 30422 10164 30478 10166
rect 30526 10218 30582 10220
rect 30526 10166 30528 10218
rect 30528 10166 30580 10218
rect 30580 10166 30582 10218
rect 30526 10164 30582 10166
rect 27356 7586 27412 7588
rect 27356 7534 27358 7586
rect 27358 7534 27410 7586
rect 27410 7534 27412 7586
rect 27356 7532 27412 7534
rect 26796 6748 26852 6804
rect 26908 5964 26964 6020
rect 26684 5628 26740 5684
rect 27132 6636 27188 6692
rect 25788 5346 25844 5348
rect 25788 5294 25790 5346
rect 25790 5294 25842 5346
rect 25842 5294 25844 5346
rect 25788 5292 25844 5294
rect 29596 9212 29652 9268
rect 28588 8988 28644 9044
rect 28476 8316 28532 8372
rect 29484 9042 29540 9044
rect 29484 8990 29486 9042
rect 29486 8990 29538 9042
rect 29538 8990 29540 9042
rect 29484 8988 29540 8990
rect 29484 8764 29540 8820
rect 27692 7308 27748 7364
rect 27468 6636 27524 6692
rect 28476 7308 28532 7364
rect 28252 6802 28308 6804
rect 28252 6750 28254 6802
rect 28254 6750 28306 6802
rect 28306 6750 28308 6802
rect 28252 6748 28308 6750
rect 27916 6690 27972 6692
rect 27916 6638 27918 6690
rect 27918 6638 27970 6690
rect 27970 6638 27972 6690
rect 27916 6636 27972 6638
rect 28588 6578 28644 6580
rect 28588 6526 28590 6578
rect 28590 6526 28642 6578
rect 28642 6526 28644 6578
rect 28588 6524 28644 6526
rect 27692 6466 27748 6468
rect 27692 6414 27694 6466
rect 27694 6414 27746 6466
rect 27746 6414 27748 6466
rect 27692 6412 27748 6414
rect 26796 5292 26852 5348
rect 25116 4898 25172 4900
rect 25116 4846 25118 4898
rect 25118 4846 25170 4898
rect 25170 4846 25172 4898
rect 25116 4844 25172 4846
rect 25900 4956 25956 5012
rect 22652 4562 22708 4564
rect 22652 4510 22654 4562
rect 22654 4510 22706 4562
rect 22706 4510 22708 4562
rect 22652 4508 22708 4510
rect 26908 4956 26964 5012
rect 28364 6466 28420 6468
rect 28364 6414 28366 6466
rect 28366 6414 28418 6466
rect 28418 6414 28420 6466
rect 28364 6412 28420 6414
rect 28700 6300 28756 6356
rect 28364 5068 28420 5124
rect 26160 4730 26216 4732
rect 26160 4678 26162 4730
rect 26162 4678 26214 4730
rect 26214 4678 26216 4730
rect 26160 4676 26216 4678
rect 26264 4730 26320 4732
rect 26264 4678 26266 4730
rect 26266 4678 26318 4730
rect 26318 4678 26320 4730
rect 26264 4676 26320 4678
rect 26368 4730 26424 4732
rect 26368 4678 26370 4730
rect 26370 4678 26422 4730
rect 26422 4678 26424 4730
rect 26368 4676 26424 4678
rect 26460 4338 26516 4340
rect 26460 4286 26462 4338
rect 26462 4286 26514 4338
rect 26514 4286 26516 4338
rect 26460 4284 26516 4286
rect 22002 3946 22058 3948
rect 22002 3894 22004 3946
rect 22004 3894 22056 3946
rect 22056 3894 22058 3946
rect 22002 3892 22058 3894
rect 22106 3946 22162 3948
rect 22106 3894 22108 3946
rect 22108 3894 22160 3946
rect 22160 3894 22162 3946
rect 22106 3892 22162 3894
rect 22210 3946 22266 3948
rect 22210 3894 22212 3946
rect 22212 3894 22264 3946
rect 22264 3894 22266 3946
rect 22210 3892 22266 3894
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 23324 3612 23380 3668
rect 20076 3554 20132 3556
rect 20076 3502 20078 3554
rect 20078 3502 20130 3554
rect 20130 3502 20132 3554
rect 20076 3500 20132 3502
rect 20748 3554 20804 3556
rect 20748 3502 20750 3554
rect 20750 3502 20802 3554
rect 20802 3502 20804 3554
rect 20748 3500 20804 3502
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 28812 8652 28868 8708
rect 28700 6018 28756 6020
rect 28700 5966 28702 6018
rect 28702 5966 28754 6018
rect 28754 5966 28756 6018
rect 28700 5964 28756 5966
rect 29260 8370 29316 8372
rect 29260 8318 29262 8370
rect 29262 8318 29314 8370
rect 29314 8318 29316 8370
rect 29260 8316 29316 8318
rect 30318 8650 30374 8652
rect 30318 8598 30320 8650
rect 30320 8598 30372 8650
rect 30372 8598 30374 8650
rect 30318 8596 30374 8598
rect 30422 8650 30478 8652
rect 30422 8598 30424 8650
rect 30424 8598 30476 8650
rect 30476 8598 30478 8650
rect 30422 8596 30478 8598
rect 30526 8650 30582 8652
rect 30526 8598 30528 8650
rect 30528 8598 30580 8650
rect 30580 8598 30582 8650
rect 30526 8596 30582 8598
rect 29820 8146 29876 8148
rect 29820 8094 29822 8146
rect 29822 8094 29874 8146
rect 29874 8094 29876 8146
rect 29820 8092 29876 8094
rect 29260 7474 29316 7476
rect 29260 7422 29262 7474
rect 29262 7422 29314 7474
rect 29314 7422 29316 7474
rect 29260 7420 29316 7422
rect 29036 6860 29092 6916
rect 29596 6802 29652 6804
rect 29596 6750 29598 6802
rect 29598 6750 29650 6802
rect 29650 6750 29652 6802
rect 29596 6748 29652 6750
rect 30318 7082 30374 7084
rect 30318 7030 30320 7082
rect 30320 7030 30372 7082
rect 30372 7030 30374 7082
rect 30318 7028 30374 7030
rect 30422 7082 30478 7084
rect 30422 7030 30424 7082
rect 30424 7030 30476 7082
rect 30476 7030 30478 7082
rect 30422 7028 30478 7030
rect 30526 7082 30582 7084
rect 30526 7030 30528 7082
rect 30528 7030 30580 7082
rect 30580 7030 30582 7082
rect 30526 7028 30582 7030
rect 29260 5852 29316 5908
rect 29932 6636 29988 6692
rect 30156 6690 30212 6692
rect 30156 6638 30158 6690
rect 30158 6638 30210 6690
rect 30210 6638 30212 6690
rect 30156 6636 30212 6638
rect 30828 10780 30884 10836
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 31836 13634 31892 13636
rect 31836 13582 31838 13634
rect 31838 13582 31890 13634
rect 31890 13582 31892 13634
rect 31836 13580 31892 13582
rect 33292 17612 33348 17668
rect 33628 17388 33684 17444
rect 33628 16268 33684 16324
rect 34188 18844 34244 18900
rect 33516 15260 33572 15316
rect 31836 12066 31892 12068
rect 31836 12014 31838 12066
rect 31838 12014 31890 12066
rect 31890 12014 31892 12066
rect 31836 12012 31892 12014
rect 31164 11564 31220 11620
rect 31836 10892 31892 10948
rect 31388 10834 31444 10836
rect 31388 10782 31390 10834
rect 31390 10782 31442 10834
rect 31442 10782 31444 10834
rect 31388 10780 31444 10782
rect 30268 6578 30324 6580
rect 30268 6526 30270 6578
rect 30270 6526 30322 6578
rect 30322 6526 30324 6578
rect 30268 6524 30324 6526
rect 29596 6412 29652 6468
rect 30604 6300 30660 6356
rect 29596 5906 29652 5908
rect 29596 5854 29598 5906
rect 29598 5854 29650 5906
rect 29650 5854 29652 5906
rect 29596 5852 29652 5854
rect 29484 5292 29540 5348
rect 30318 5514 30374 5516
rect 30318 5462 30320 5514
rect 30320 5462 30372 5514
rect 30372 5462 30374 5514
rect 30318 5460 30374 5462
rect 30422 5514 30478 5516
rect 30422 5462 30424 5514
rect 30424 5462 30476 5514
rect 30476 5462 30478 5514
rect 30422 5460 30478 5462
rect 30526 5514 30582 5516
rect 30526 5462 30528 5514
rect 30528 5462 30580 5514
rect 30580 5462 30582 5514
rect 30526 5460 30582 5462
rect 29932 5010 29988 5012
rect 29932 4958 29934 5010
rect 29934 4958 29986 5010
rect 29986 4958 29988 5010
rect 29932 4956 29988 4958
rect 31164 6690 31220 6692
rect 31164 6638 31166 6690
rect 31166 6638 31218 6690
rect 31218 6638 31220 6690
rect 31164 6636 31220 6638
rect 31052 6524 31108 6580
rect 31164 6412 31220 6468
rect 30940 5740 30996 5796
rect 32060 9548 32116 9604
rect 31612 7644 31668 7700
rect 31836 7420 31892 7476
rect 32620 9266 32676 9268
rect 32620 9214 32622 9266
rect 32622 9214 32674 9266
rect 32674 9214 32676 9266
rect 32620 9212 32676 9214
rect 32844 8988 32900 9044
rect 32060 6524 32116 6580
rect 31388 6076 31444 6132
rect 31836 6130 31892 6132
rect 31836 6078 31838 6130
rect 31838 6078 31890 6130
rect 31890 6078 31892 6130
rect 31836 6076 31892 6078
rect 31500 5740 31556 5796
rect 31276 5628 31332 5684
rect 32172 7308 32228 7364
rect 32396 6076 32452 6132
rect 32060 5292 32116 5348
rect 32844 5180 32900 5236
rect 28588 4284 28644 4340
rect 28476 4172 28532 4228
rect 30318 3946 30374 3948
rect 30318 3894 30320 3946
rect 30320 3894 30372 3946
rect 30372 3894 30374 3946
rect 30318 3892 30374 3894
rect 30422 3946 30478 3948
rect 30422 3894 30424 3946
rect 30424 3894 30476 3946
rect 30476 3894 30478 3946
rect 30422 3892 30478 3894
rect 30526 3946 30582 3948
rect 30526 3894 30528 3946
rect 30528 3894 30580 3946
rect 30580 3894 30582 3946
rect 30526 3892 30582 3894
rect 27580 3724 27636 3780
rect 26012 3500 26068 3556
rect 26908 3612 26964 3668
rect 26160 3162 26216 3164
rect 26160 3110 26162 3162
rect 26162 3110 26214 3162
rect 26214 3110 26216 3162
rect 26160 3108 26216 3110
rect 26264 3162 26320 3164
rect 26264 3110 26266 3162
rect 26266 3110 26318 3162
rect 26318 3110 26320 3162
rect 26264 3108 26320 3110
rect 26368 3162 26424 3164
rect 26368 3110 26370 3162
rect 26370 3110 26422 3162
rect 26422 3110 26424 3162
rect 26368 3108 26424 3110
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 28588 3554 28644 3556
rect 28588 3502 28590 3554
rect 28590 3502 28642 3554
rect 28642 3502 28644 3554
rect 28588 3500 28644 3502
rect 33628 12962 33684 12964
rect 33628 12910 33630 12962
rect 33630 12910 33682 12962
rect 33682 12910 33684 12962
rect 33628 12908 33684 12910
rect 34076 12796 34132 12852
rect 34188 15148 34244 15204
rect 34476 18842 34532 18844
rect 34476 18790 34478 18842
rect 34478 18790 34530 18842
rect 34530 18790 34532 18842
rect 34476 18788 34532 18790
rect 34580 18842 34636 18844
rect 34580 18790 34582 18842
rect 34582 18790 34634 18842
rect 34634 18790 34636 18842
rect 34580 18788 34636 18790
rect 34684 18842 34740 18844
rect 34684 18790 34686 18842
rect 34686 18790 34738 18842
rect 34738 18790 34740 18842
rect 34684 18788 34740 18790
rect 34476 17274 34532 17276
rect 34476 17222 34478 17274
rect 34478 17222 34530 17274
rect 34530 17222 34532 17274
rect 34476 17220 34532 17222
rect 34580 17274 34636 17276
rect 34580 17222 34582 17274
rect 34582 17222 34634 17274
rect 34634 17222 34636 17274
rect 34580 17220 34636 17222
rect 34684 17274 34740 17276
rect 34684 17222 34686 17274
rect 34686 17222 34738 17274
rect 34738 17222 34740 17274
rect 34684 17220 34740 17222
rect 34476 15706 34532 15708
rect 34476 15654 34478 15706
rect 34478 15654 34530 15706
rect 34530 15654 34532 15706
rect 34476 15652 34532 15654
rect 34580 15706 34636 15708
rect 34580 15654 34582 15706
rect 34582 15654 34634 15706
rect 34634 15654 34636 15706
rect 34580 15652 34636 15654
rect 34684 15706 34740 15708
rect 34684 15654 34686 15706
rect 34686 15654 34738 15706
rect 34738 15654 34740 15706
rect 34684 15652 34740 15654
rect 34476 14138 34532 14140
rect 34476 14086 34478 14138
rect 34478 14086 34530 14138
rect 34530 14086 34532 14138
rect 34476 14084 34532 14086
rect 34580 14138 34636 14140
rect 34580 14086 34582 14138
rect 34582 14086 34634 14138
rect 34634 14086 34636 14138
rect 34580 14084 34636 14086
rect 34684 14138 34740 14140
rect 34684 14086 34686 14138
rect 34686 14086 34738 14138
rect 34738 14086 34740 14138
rect 34684 14084 34740 14086
rect 34476 12570 34532 12572
rect 34476 12518 34478 12570
rect 34478 12518 34530 12570
rect 34530 12518 34532 12570
rect 34476 12516 34532 12518
rect 34580 12570 34636 12572
rect 34580 12518 34582 12570
rect 34582 12518 34634 12570
rect 34634 12518 34636 12570
rect 34580 12516 34636 12518
rect 34684 12570 34740 12572
rect 34684 12518 34686 12570
rect 34686 12518 34738 12570
rect 34738 12518 34740 12570
rect 34684 12516 34740 12518
rect 33180 10668 33236 10724
rect 34300 11170 34356 11172
rect 34300 11118 34302 11170
rect 34302 11118 34354 11170
rect 34354 11118 34356 11170
rect 34300 11116 34356 11118
rect 34476 11002 34532 11004
rect 34476 10950 34478 11002
rect 34478 10950 34530 11002
rect 34530 10950 34532 11002
rect 34476 10948 34532 10950
rect 34580 11002 34636 11004
rect 34580 10950 34582 11002
rect 34582 10950 34634 11002
rect 34634 10950 34636 11002
rect 34580 10948 34636 10950
rect 34684 11002 34740 11004
rect 34684 10950 34686 11002
rect 34686 10950 34738 11002
rect 34738 10950 34740 11002
rect 34684 10948 34740 10950
rect 33516 10556 33572 10612
rect 33404 9548 33460 9604
rect 34476 9434 34532 9436
rect 34476 9382 34478 9434
rect 34478 9382 34530 9434
rect 34530 9382 34532 9434
rect 34476 9380 34532 9382
rect 34580 9434 34636 9436
rect 34580 9382 34582 9434
rect 34582 9382 34634 9434
rect 34634 9382 34636 9434
rect 34580 9380 34636 9382
rect 34684 9434 34740 9436
rect 34684 9382 34686 9434
rect 34686 9382 34738 9434
rect 34738 9382 34740 9434
rect 34684 9380 34740 9382
rect 33404 9042 33460 9044
rect 33404 8990 33406 9042
rect 33406 8990 33458 9042
rect 33458 8990 33460 9042
rect 33404 8988 33460 8990
rect 33964 8988 34020 9044
rect 33180 6130 33236 6132
rect 33180 6078 33182 6130
rect 33182 6078 33234 6130
rect 33234 6078 33236 6130
rect 33180 6076 33236 6078
rect 33180 5740 33236 5796
rect 33292 5068 33348 5124
rect 33516 6860 33572 6916
rect 32620 4338 32676 4340
rect 32620 4286 32622 4338
rect 32622 4286 32674 4338
rect 32674 4286 32676 4338
rect 32620 4284 32676 4286
rect 33068 4226 33124 4228
rect 33068 4174 33070 4226
rect 33070 4174 33122 4226
rect 33122 4174 33124 4226
rect 33068 4172 33124 4174
rect 31724 3554 31780 3556
rect 31724 3502 31726 3554
rect 31726 3502 31778 3554
rect 31778 3502 31780 3554
rect 31724 3500 31780 3502
rect 33292 3554 33348 3556
rect 33292 3502 33294 3554
rect 33294 3502 33346 3554
rect 33346 3502 33348 3554
rect 33292 3500 33348 3502
rect 32508 3442 32564 3444
rect 32508 3390 32510 3442
rect 32510 3390 32562 3442
rect 32562 3390 32564 3442
rect 32508 3388 32564 3390
rect 34476 7866 34532 7868
rect 34476 7814 34478 7866
rect 34478 7814 34530 7866
rect 34530 7814 34532 7866
rect 34476 7812 34532 7814
rect 34580 7866 34636 7868
rect 34580 7814 34582 7866
rect 34582 7814 34634 7866
rect 34634 7814 34636 7866
rect 34580 7812 34636 7814
rect 34684 7866 34740 7868
rect 34684 7814 34686 7866
rect 34686 7814 34738 7866
rect 34738 7814 34740 7866
rect 34684 7812 34740 7814
rect 34076 6860 34132 6916
rect 34188 7196 34244 7252
rect 33852 6748 33908 6804
rect 33516 6578 33572 6580
rect 33516 6526 33518 6578
rect 33518 6526 33570 6578
rect 33570 6526 33572 6578
rect 33516 6524 33572 6526
rect 33740 5628 33796 5684
rect 33628 5404 33684 5460
rect 34300 6466 34356 6468
rect 34300 6414 34302 6466
rect 34302 6414 34354 6466
rect 34354 6414 34356 6466
rect 34300 6412 34356 6414
rect 34476 6298 34532 6300
rect 34476 6246 34478 6298
rect 34478 6246 34530 6298
rect 34530 6246 34532 6298
rect 34476 6244 34532 6246
rect 34580 6298 34636 6300
rect 34580 6246 34582 6298
rect 34582 6246 34634 6298
rect 34634 6246 34636 6298
rect 34580 6244 34636 6246
rect 34684 6298 34740 6300
rect 34684 6246 34686 6298
rect 34686 6246 34738 6298
rect 34738 6246 34740 6298
rect 34684 6244 34740 6246
rect 34076 5852 34132 5908
rect 34188 5740 34244 5796
rect 34188 5122 34244 5124
rect 34188 5070 34190 5122
rect 34190 5070 34242 5122
rect 34242 5070 34244 5122
rect 34188 5068 34244 5070
rect 34076 4338 34132 4340
rect 34076 4286 34078 4338
rect 34078 4286 34130 4338
rect 34130 4286 34132 4338
rect 34076 4284 34132 4286
rect 34476 4730 34532 4732
rect 34476 4678 34478 4730
rect 34478 4678 34530 4730
rect 34530 4678 34532 4730
rect 34476 4676 34532 4678
rect 34580 4730 34636 4732
rect 34580 4678 34582 4730
rect 34582 4678 34634 4730
rect 34634 4678 34636 4730
rect 34580 4676 34636 4678
rect 34684 4730 34740 4732
rect 34684 4678 34686 4730
rect 34686 4678 34738 4730
rect 34738 4678 34740 4730
rect 34684 4676 34740 4678
rect 34300 4284 34356 4340
rect 34076 3724 34132 3780
rect 33292 1148 33348 1204
rect 34188 3442 34244 3444
rect 34188 3390 34190 3442
rect 34190 3390 34242 3442
rect 34242 3390 34244 3442
rect 34188 3388 34244 3390
rect 34476 3162 34532 3164
rect 34476 3110 34478 3162
rect 34478 3110 34530 3162
rect 34530 3110 34532 3162
rect 34476 3108 34532 3110
rect 34580 3162 34636 3164
rect 34580 3110 34582 3162
rect 34582 3110 34634 3162
rect 34634 3110 34636 3162
rect 34580 3108 34636 3110
rect 34684 3162 34740 3164
rect 34684 3110 34686 3162
rect 34686 3110 34738 3162
rect 34738 3110 34740 3162
rect 34684 3108 34740 3110
rect 34188 2716 34244 2772
<< metal3 >>
rect 35200 24724 36000 24752
rect 31602 24668 31612 24724
rect 31668 24668 36000 24724
rect 35200 24640 36000 24668
rect 0 24052 800 24080
rect 0 23996 2044 24052
rect 2100 23996 2110 24052
rect 0 23968 800 23996
rect 5394 23436 5404 23492
rect 5460 23436 6636 23492
rect 6692 23436 6702 23492
rect 35200 23156 36000 23184
rect 25106 23100 25116 23156
rect 25172 23100 36000 23156
rect 35200 23072 36000 23100
rect 5360 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5644 22764
rect 13676 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13960 22764
rect 21992 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22276 22764
rect 30308 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30592 22764
rect 12562 22540 12572 22596
rect 12628 22540 14140 22596
rect 14196 22540 14206 22596
rect 16146 22540 16156 22596
rect 16212 22540 17164 22596
rect 17220 22540 17230 22596
rect 19730 22540 19740 22596
rect 19796 22540 20972 22596
rect 21028 22540 21038 22596
rect 23314 22540 23324 22596
rect 23380 22540 25564 22596
rect 25620 22540 25630 22596
rect 26898 22540 26908 22596
rect 26964 22540 28588 22596
rect 28644 22540 28654 22596
rect 26562 22204 26572 22260
rect 26628 22204 27468 22260
rect 27524 22204 27534 22260
rect 23314 22092 23324 22148
rect 23380 22092 23772 22148
rect 23828 22092 24780 22148
rect 24836 22092 24846 22148
rect 0 22036 800 22064
rect 0 21980 1932 22036
rect 1988 21980 1998 22036
rect 0 21952 800 21980
rect 9518 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9802 21980
rect 17834 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18118 21980
rect 26150 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26434 21980
rect 34466 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34750 21980
rect 8978 21756 8988 21812
rect 9044 21756 11004 21812
rect 11060 21756 11070 21812
rect 12898 21756 12908 21812
rect 12964 21756 17388 21812
rect 17444 21756 17454 21812
rect 19292 21644 29372 21700
rect 29428 21644 29438 21700
rect 4050 21420 4060 21476
rect 4116 21420 6076 21476
rect 6132 21420 6142 21476
rect 19292 21364 19348 21644
rect 35200 21588 36000 21616
rect 25890 21532 25900 21588
rect 25956 21532 26796 21588
rect 26852 21532 26862 21588
rect 31154 21532 31164 21588
rect 31220 21532 36000 21588
rect 35200 21504 36000 21532
rect 19618 21420 19628 21476
rect 19684 21420 20524 21476
rect 20580 21420 20590 21476
rect 25666 21420 25676 21476
rect 25732 21420 31052 21476
rect 31108 21420 31118 21476
rect 4274 21308 4284 21364
rect 4340 21308 5068 21364
rect 5124 21308 5134 21364
rect 16930 21308 16940 21364
rect 16996 21308 17948 21364
rect 18004 21308 19292 21364
rect 19348 21308 19358 21364
rect 24658 21308 24668 21364
rect 24724 21308 25452 21364
rect 25508 21308 25518 21364
rect 27570 21308 27580 21364
rect 27636 21308 33628 21364
rect 33684 21308 33694 21364
rect 5360 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5644 21196
rect 13676 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13960 21196
rect 21992 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22276 21196
rect 30308 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30592 21196
rect 31042 21084 31052 21140
rect 31108 21084 31612 21140
rect 31668 21084 31678 21140
rect 9986 20972 9996 21028
rect 10052 20972 10062 21028
rect 17714 20972 17724 21028
rect 17780 20972 27132 21028
rect 27188 20972 29148 21028
rect 29204 20972 29214 21028
rect 9996 20916 10052 20972
rect 9762 20860 9772 20916
rect 9828 20860 23156 20916
rect 27570 20860 27580 20916
rect 27636 20860 30716 20916
rect 30772 20860 30782 20916
rect 23100 20804 23156 20860
rect 2706 20748 2716 20804
rect 2772 20748 3836 20804
rect 3892 20748 3902 20804
rect 9986 20748 9996 20804
rect 10052 20748 14252 20804
rect 14308 20748 14812 20804
rect 14868 20748 14878 20804
rect 15250 20748 15260 20804
rect 15316 20748 16940 20804
rect 16996 20748 17006 20804
rect 19730 20748 19740 20804
rect 19796 20748 22932 20804
rect 23090 20748 23100 20804
rect 23156 20748 23166 20804
rect 25554 20748 25564 20804
rect 25620 20748 26124 20804
rect 26180 20748 26190 20804
rect 27794 20748 27804 20804
rect 27860 20748 30380 20804
rect 30436 20748 31276 20804
rect 31332 20748 31342 20804
rect 22876 20692 22932 20748
rect 14466 20636 14476 20692
rect 14532 20636 15148 20692
rect 15204 20636 15214 20692
rect 19394 20636 19404 20692
rect 19460 20636 20300 20692
rect 20356 20636 20366 20692
rect 22876 20636 25228 20692
rect 25284 20636 25294 20692
rect 9518 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9802 20412
rect 17834 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18118 20412
rect 25228 20244 25284 20636
rect 26124 20580 26180 20748
rect 26786 20636 26796 20692
rect 26852 20636 29708 20692
rect 29764 20636 29774 20692
rect 26124 20524 29932 20580
rect 29988 20524 30604 20580
rect 30660 20524 30670 20580
rect 26150 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26434 20412
rect 34466 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34750 20412
rect 19842 20188 19852 20244
rect 19908 20188 24668 20244
rect 24724 20188 24734 20244
rect 25228 20188 26628 20244
rect 28466 20188 28476 20244
rect 28532 20188 30716 20244
rect 30772 20188 31836 20244
rect 31892 20188 31902 20244
rect 26572 20132 26628 20188
rect 6514 20076 6524 20132
rect 6580 20076 9772 20132
rect 9828 20076 9838 20132
rect 10546 20076 10556 20132
rect 10612 20076 13244 20132
rect 13300 20076 13310 20132
rect 13458 20076 13468 20132
rect 13524 20076 16156 20132
rect 16212 20076 17724 20132
rect 17780 20076 17790 20132
rect 26534 20076 26572 20132
rect 26628 20076 28924 20132
rect 28980 20076 28990 20132
rect 0 20020 800 20048
rect 13244 20020 13300 20076
rect 35200 20020 36000 20048
rect 0 19964 1932 20020
rect 1988 19964 1998 20020
rect 10434 19964 10444 20020
rect 10500 19964 10892 20020
rect 10948 19964 10958 20020
rect 11218 19964 11228 20020
rect 11284 19964 12012 20020
rect 12068 19964 12078 20020
rect 13244 19964 14252 20020
rect 14308 19964 14318 20020
rect 15026 19964 15036 20020
rect 15092 19964 15372 20020
rect 15428 19964 20076 20020
rect 20132 19964 20142 20020
rect 28466 19964 28476 20020
rect 28532 19964 36000 20020
rect 0 19936 800 19964
rect 35200 19936 36000 19964
rect 12114 19852 12124 19908
rect 12180 19852 14812 19908
rect 14868 19852 14878 19908
rect 23874 19740 23884 19796
rect 23940 19740 25788 19796
rect 25844 19740 25854 19796
rect 5360 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5644 19628
rect 13676 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13960 19628
rect 21992 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22276 19628
rect 30308 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30592 19628
rect 10882 19404 10892 19460
rect 10948 19404 20860 19460
rect 20916 19404 23996 19460
rect 24052 19404 25340 19460
rect 25396 19404 25406 19460
rect 27570 19404 27580 19460
rect 27636 19404 33964 19460
rect 34020 19404 34030 19460
rect 27906 19292 27916 19348
rect 27972 19292 33852 19348
rect 33908 19292 33918 19348
rect 14242 19180 14252 19236
rect 14308 19180 14812 19236
rect 14868 19180 14878 19236
rect 15138 19180 15148 19236
rect 15204 19180 19180 19236
rect 19236 19180 19516 19236
rect 19572 19180 19582 19236
rect 30818 19180 30828 19236
rect 30884 19180 33180 19236
rect 33236 19180 33740 19236
rect 33796 19180 33806 19236
rect 9202 19068 9212 19124
rect 9268 19068 9436 19124
rect 9492 19068 9502 19124
rect 18498 19068 18508 19124
rect 18564 19068 18956 19124
rect 19012 19068 19022 19124
rect 19394 19068 19404 19124
rect 19460 19068 23884 19124
rect 23940 19068 23950 19124
rect 28466 19068 28476 19124
rect 28532 19068 33292 19124
rect 33348 19068 33358 19124
rect 16146 18956 16156 19012
rect 16212 18956 19068 19012
rect 19124 18956 19134 19012
rect 29810 18956 29820 19012
rect 29876 18956 31388 19012
rect 31444 18956 31454 19012
rect 32946 18956 32956 19012
rect 33012 18956 34076 19012
rect 34132 18956 34142 19012
rect 33842 18844 33852 18900
rect 33908 18844 34188 18900
rect 34244 18844 34254 18900
rect 9518 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9802 18844
rect 17834 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18118 18844
rect 26150 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26434 18844
rect 34466 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34750 18844
rect 9202 18732 9212 18788
rect 9268 18732 9278 18788
rect 9212 18676 9268 18732
rect 8754 18620 8764 18676
rect 8820 18620 9660 18676
rect 9716 18620 10892 18676
rect 10948 18620 10958 18676
rect 29362 18620 29372 18676
rect 29428 18620 31164 18676
rect 31220 18620 31230 18676
rect 35200 18452 36000 18480
rect 5730 18396 5740 18452
rect 5796 18396 8428 18452
rect 9090 18396 9100 18452
rect 9156 18396 11676 18452
rect 11732 18396 13692 18452
rect 13748 18396 14476 18452
rect 14532 18396 14542 18452
rect 20514 18396 20524 18452
rect 20580 18396 20860 18452
rect 20916 18396 20926 18452
rect 24434 18396 24444 18452
rect 24500 18396 25228 18452
rect 25284 18396 25294 18452
rect 25554 18396 25564 18452
rect 25620 18396 26236 18452
rect 26292 18396 29036 18452
rect 29092 18396 29102 18452
rect 31826 18396 31836 18452
rect 31892 18396 36000 18452
rect 8372 18284 8428 18396
rect 35200 18368 36000 18396
rect 8484 18284 8494 18340
rect 25778 18284 25788 18340
rect 25844 18284 26460 18340
rect 26516 18284 26526 18340
rect 2706 18172 2716 18228
rect 2772 18172 2782 18228
rect 29250 18172 29260 18228
rect 29316 18172 33068 18228
rect 33124 18172 33134 18228
rect 0 18004 800 18032
rect 2716 18004 2772 18172
rect 5360 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5644 18060
rect 13676 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13960 18060
rect 21992 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22276 18060
rect 30308 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30592 18060
rect 0 17948 2772 18004
rect 0 17920 800 17948
rect 6514 17836 6524 17892
rect 6580 17836 8988 17892
rect 9044 17836 9054 17892
rect 27916 17724 30828 17780
rect 30884 17724 30894 17780
rect 27916 17668 27972 17724
rect 10994 17612 11004 17668
rect 11060 17612 11788 17668
rect 11844 17612 11854 17668
rect 19506 17612 19516 17668
rect 19572 17612 20076 17668
rect 20132 17612 20142 17668
rect 27570 17612 27580 17668
rect 27636 17612 27916 17668
rect 27972 17612 27982 17668
rect 29474 17612 29484 17668
rect 29540 17612 30268 17668
rect 30324 17612 33292 17668
rect 33348 17612 33358 17668
rect 8978 17500 8988 17556
rect 9044 17500 9660 17556
rect 9716 17500 10108 17556
rect 10164 17500 11452 17556
rect 11508 17500 11518 17556
rect 19282 17500 19292 17556
rect 19348 17500 25788 17556
rect 25844 17500 25854 17556
rect 14578 17388 14588 17444
rect 14644 17388 16156 17444
rect 16212 17388 16222 17444
rect 25900 17388 28588 17444
rect 28644 17388 29148 17444
rect 29204 17388 29214 17444
rect 31378 17388 31388 17444
rect 31444 17388 33628 17444
rect 33684 17388 33694 17444
rect 25900 17332 25956 17388
rect 19618 17276 19628 17332
rect 19684 17276 23660 17332
rect 23716 17276 23726 17332
rect 25890 17276 25900 17332
rect 25956 17276 25966 17332
rect 29026 17276 29036 17332
rect 29092 17276 29932 17332
rect 29988 17276 29998 17332
rect 9518 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9802 17276
rect 17834 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18118 17276
rect 25900 17108 25956 17276
rect 26150 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26434 17276
rect 34466 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34750 17276
rect 11442 17052 11452 17108
rect 11508 17052 12348 17108
rect 12404 17052 25956 17108
rect 27682 17052 27692 17108
rect 27748 17052 32060 17108
rect 32116 17052 32126 17108
rect 2716 16940 8652 16996
rect 8708 16940 10668 16996
rect 10724 16940 10734 16996
rect 18834 16940 18844 16996
rect 18900 16940 18910 16996
rect 23650 16940 23660 16996
rect 23716 16940 28700 16996
rect 28756 16940 29260 16996
rect 29316 16940 29326 16996
rect 29586 16940 29596 16996
rect 29652 16940 30604 16996
rect 30660 16940 31724 16996
rect 31780 16940 31790 16996
rect 2716 16884 2772 16940
rect 18844 16884 18900 16940
rect 29596 16884 29652 16940
rect 35200 16884 36000 16912
rect 2706 16828 2716 16884
rect 2772 16828 2782 16884
rect 4946 16828 4956 16884
rect 5012 16828 6972 16884
rect 7028 16828 7038 16884
rect 15586 16828 15596 16884
rect 15652 16828 15662 16884
rect 18610 16828 18620 16884
rect 18676 16828 19740 16884
rect 19796 16828 19806 16884
rect 20066 16828 20076 16884
rect 20132 16828 20636 16884
rect 20692 16828 22988 16884
rect 23044 16828 23054 16884
rect 28466 16828 28476 16884
rect 28532 16828 29652 16884
rect 31602 16828 31612 16884
rect 31668 16828 36000 16884
rect 15596 16660 15652 16828
rect 35200 16800 36000 16828
rect 16034 16716 16044 16772
rect 16100 16716 18844 16772
rect 18900 16716 18910 16772
rect 26674 16716 26684 16772
rect 26740 16716 27356 16772
rect 27412 16716 27422 16772
rect 5506 16604 5516 16660
rect 5572 16604 7980 16660
rect 8036 16604 8046 16660
rect 15596 16604 18956 16660
rect 19012 16604 20188 16660
rect 5360 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5644 16492
rect 13676 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13960 16492
rect 20132 16324 20188 16604
rect 21992 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22276 16492
rect 30308 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30592 16492
rect 20132 16268 22204 16324
rect 22260 16268 22270 16324
rect 23090 16268 23100 16324
rect 23156 16268 26180 16324
rect 30034 16268 30044 16324
rect 30100 16268 33628 16324
rect 33684 16268 33694 16324
rect 1922 16156 1932 16212
rect 1988 16156 1998 16212
rect 0 15988 800 16016
rect 1932 15988 1988 16156
rect 26124 16100 26180 16268
rect 7186 16044 7196 16100
rect 7252 16044 10780 16100
rect 10836 16044 14924 16100
rect 14980 16044 14990 16100
rect 20850 16044 20860 16100
rect 20916 16044 21420 16100
rect 21476 16044 25564 16100
rect 25620 16044 25630 16100
rect 26114 16044 26124 16100
rect 26180 16044 26908 16100
rect 26964 16044 26974 16100
rect 28476 16044 28924 16100
rect 28980 16044 29372 16100
rect 29428 16044 29438 16100
rect 28476 15988 28532 16044
rect 0 15932 1988 15988
rect 7522 15932 7532 15988
rect 7588 15932 11228 15988
rect 11284 15932 11294 15988
rect 12002 15932 12012 15988
rect 12068 15932 18340 15988
rect 0 15904 800 15932
rect 6290 15820 6300 15876
rect 6356 15820 7196 15876
rect 7252 15820 7262 15876
rect 10770 15820 10780 15876
rect 10836 15820 13580 15876
rect 13636 15820 13646 15876
rect 18284 15764 18340 15932
rect 19068 15932 21980 15988
rect 22036 15932 28532 15988
rect 29250 15932 29260 15988
rect 29316 15932 29708 15988
rect 29764 15932 30156 15988
rect 30212 15932 30604 15988
rect 30660 15932 30670 15988
rect 19068 15876 19124 15932
rect 18498 15820 18508 15876
rect 18564 15820 18732 15876
rect 18788 15820 19124 15876
rect 20132 15820 21644 15876
rect 21700 15820 22540 15876
rect 22596 15820 22606 15876
rect 28130 15820 28140 15876
rect 28196 15820 29148 15876
rect 29204 15820 29214 15876
rect 20132 15764 20188 15820
rect 18284 15708 20188 15764
rect 9518 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9802 15708
rect 17834 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18118 15708
rect 26150 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26434 15708
rect 34466 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34750 15708
rect 22978 15596 22988 15652
rect 23044 15596 23548 15652
rect 23604 15596 23614 15652
rect 26852 15596 28700 15652
rect 28756 15596 29932 15652
rect 29988 15596 29998 15652
rect 26852 15540 26908 15596
rect 4620 15484 7308 15540
rect 7364 15484 7374 15540
rect 18386 15484 18396 15540
rect 18452 15484 19404 15540
rect 19460 15484 19852 15540
rect 19908 15484 19918 15540
rect 20132 15484 26908 15540
rect 27458 15484 27468 15540
rect 27524 15484 27804 15540
rect 27860 15484 27870 15540
rect 4620 15316 4676 15484
rect 20132 15428 20188 15484
rect 27468 15428 27524 15484
rect 7074 15372 7084 15428
rect 7140 15372 7644 15428
rect 7700 15372 7710 15428
rect 11106 15372 11116 15428
rect 11172 15372 20188 15428
rect 20626 15372 20636 15428
rect 20692 15372 27524 15428
rect 35200 15316 36000 15344
rect 1698 15260 1708 15316
rect 1764 15260 3836 15316
rect 3892 15260 4620 15316
rect 4676 15260 4686 15316
rect 5842 15260 5852 15316
rect 5908 15260 6412 15316
rect 6468 15260 7308 15316
rect 7364 15260 7374 15316
rect 11442 15260 11452 15316
rect 11508 15260 17724 15316
rect 17780 15260 18732 15316
rect 18788 15260 18798 15316
rect 33506 15260 33516 15316
rect 33572 15260 36000 15316
rect 14018 15148 14028 15204
rect 14084 15148 14812 15204
rect 14868 15148 15596 15204
rect 15652 15148 15662 15204
rect 14028 15092 14084 15148
rect 13346 15036 13356 15092
rect 13412 15036 14084 15092
rect 16044 15092 16100 15260
rect 35200 15232 36000 15260
rect 22418 15148 22428 15204
rect 22484 15148 22652 15204
rect 22708 15148 26684 15204
rect 26740 15148 28924 15204
rect 28980 15148 28990 15204
rect 31602 15148 31612 15204
rect 31668 15148 34188 15204
rect 34244 15148 34254 15204
rect 16044 15036 16156 15092
rect 16212 15036 16222 15092
rect 23650 15036 23660 15092
rect 23716 15036 24220 15092
rect 24276 15036 28700 15092
rect 28756 15036 28766 15092
rect 3938 14924 3948 14980
rect 4004 14924 4284 14980
rect 4340 14924 4350 14980
rect 5360 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5644 14924
rect 13676 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13960 14924
rect 21992 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22276 14924
rect 30308 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30592 14924
rect 6626 14588 6636 14644
rect 6692 14588 8092 14644
rect 8148 14588 10444 14644
rect 10500 14588 11116 14644
rect 11172 14588 11182 14644
rect 28914 14588 28924 14644
rect 28980 14588 29484 14644
rect 29540 14588 29550 14644
rect 2034 14476 2044 14532
rect 2100 14476 2604 14532
rect 2660 14476 3276 14532
rect 3332 14476 3342 14532
rect 4274 14476 4284 14532
rect 4340 14476 6076 14532
rect 6132 14476 6142 14532
rect 22866 14476 22876 14532
rect 22932 14476 23548 14532
rect 23604 14476 23614 14532
rect 2930 14364 2940 14420
rect 2996 14364 3612 14420
rect 3668 14364 4172 14420
rect 4228 14364 6524 14420
rect 6580 14364 6590 14420
rect 23650 14364 23660 14420
rect 23716 14364 24220 14420
rect 24276 14364 24286 14420
rect 26786 14364 26796 14420
rect 26852 14364 31388 14420
rect 31444 14364 31454 14420
rect 4722 14252 4732 14308
rect 4788 14252 5516 14308
rect 5572 14252 5582 14308
rect 7634 14252 7644 14308
rect 7700 14252 9996 14308
rect 10052 14252 20412 14308
rect 20468 14252 21420 14308
rect 21476 14252 21486 14308
rect 22754 14252 22764 14308
rect 22820 14252 23436 14308
rect 23492 14252 27580 14308
rect 27636 14252 27646 14308
rect 9518 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9802 14140
rect 17834 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18118 14140
rect 26150 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26434 14140
rect 34466 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34750 14140
rect 3826 14028 3836 14084
rect 3892 14028 4396 14084
rect 4452 14028 4956 14084
rect 5012 14028 7532 14084
rect 7588 14028 7598 14084
rect 0 13972 800 14000
rect 0 13916 1820 13972
rect 1876 13916 1886 13972
rect 2930 13916 2940 13972
rect 2996 13916 3388 13972
rect 6514 13916 6524 13972
rect 6580 13916 7420 13972
rect 7476 13916 8540 13972
rect 8596 13916 8606 13972
rect 15092 13916 27468 13972
rect 27524 13916 27534 13972
rect 0 13888 800 13916
rect 3332 13804 3388 13916
rect 15092 13860 15148 13916
rect 3444 13804 15148 13860
rect 20626 13804 20636 13860
rect 20692 13804 22204 13860
rect 22260 13804 22270 13860
rect 27794 13804 27804 13860
rect 27860 13804 28588 13860
rect 28644 13804 28654 13860
rect 31892 13804 33684 13860
rect 2482 13692 2492 13748
rect 2548 13692 4172 13748
rect 4228 13692 4238 13748
rect 8306 13692 8316 13748
rect 8372 13692 8382 13748
rect 21074 13692 21084 13748
rect 21140 13692 21756 13748
rect 21812 13692 21822 13748
rect 4610 13580 4620 13636
rect 4676 13580 7084 13636
rect 7140 13580 7150 13636
rect 8316 13524 8372 13692
rect 11442 13580 11452 13636
rect 11508 13580 12348 13636
rect 12404 13580 19964 13636
rect 20020 13580 20030 13636
rect 31826 13580 31836 13636
rect 31892 13580 31948 13804
rect 33628 13748 33684 13804
rect 35200 13748 36000 13776
rect 33058 13692 33068 13748
rect 33124 13692 33134 13748
rect 33628 13692 36000 13748
rect 33068 13524 33124 13692
rect 35200 13664 36000 13692
rect 8316 13468 15596 13524
rect 15652 13468 16492 13524
rect 16548 13468 16558 13524
rect 16930 13468 16940 13524
rect 16996 13468 18620 13524
rect 18676 13468 19516 13524
rect 19572 13468 19582 13524
rect 30706 13468 30716 13524
rect 30772 13468 33124 13524
rect 5360 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5644 13356
rect 13676 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13960 13356
rect 21992 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22276 13356
rect 30308 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30592 13356
rect 23986 13244 23996 13300
rect 24052 13244 29260 13300
rect 29316 13244 29326 13300
rect 3154 13132 3164 13188
rect 3220 13132 11676 13188
rect 11732 13132 11742 13188
rect 13458 13132 13468 13188
rect 13524 13132 20076 13188
rect 20132 13132 20524 13188
rect 20580 13132 20590 13188
rect 29586 13132 29596 13188
rect 29652 13132 33684 13188
rect 12450 13020 12460 13076
rect 12516 13020 14924 13076
rect 14980 13020 15708 13076
rect 15764 13020 21868 13076
rect 21924 13020 21934 13076
rect 33628 12964 33684 13132
rect 5852 12908 6076 12964
rect 6132 12908 6142 12964
rect 15026 12908 15036 12964
rect 15092 12908 15820 12964
rect 15876 12908 15886 12964
rect 19394 12908 19404 12964
rect 19460 12908 22092 12964
rect 22148 12908 23884 12964
rect 23940 12908 23950 12964
rect 29250 12908 29260 12964
rect 29316 12908 31948 12964
rect 33618 12908 33628 12964
rect 33684 12908 33694 12964
rect 5852 12852 5908 12908
rect 31892 12852 31948 12908
rect 5394 12796 5404 12852
rect 5460 12796 5852 12852
rect 5908 12796 5918 12852
rect 14802 12796 14812 12852
rect 14868 12796 16044 12852
rect 16100 12796 16604 12852
rect 16660 12796 16670 12852
rect 24658 12796 24668 12852
rect 24724 12796 27132 12852
rect 27188 12796 27198 12852
rect 31892 12796 34076 12852
rect 34132 12796 34142 12852
rect 8418 12684 8428 12740
rect 8484 12684 12236 12740
rect 12292 12684 12302 12740
rect 13906 12684 13916 12740
rect 13972 12684 14700 12740
rect 14756 12684 14766 12740
rect 19058 12684 19068 12740
rect 19124 12684 19740 12740
rect 19796 12684 19806 12740
rect 21522 12684 21532 12740
rect 21588 12684 24556 12740
rect 24612 12684 24622 12740
rect 6290 12572 6300 12628
rect 6356 12572 6860 12628
rect 6916 12572 6926 12628
rect 19842 12572 19852 12628
rect 19908 12572 20188 12628
rect 20244 12572 20254 12628
rect 23650 12572 23660 12628
rect 23716 12572 23996 12628
rect 24052 12572 24062 12628
rect 9518 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9802 12572
rect 17834 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18118 12572
rect 26150 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26434 12572
rect 34466 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34750 12572
rect 2258 12348 2268 12404
rect 2324 12348 6188 12404
rect 6244 12348 6254 12404
rect 7298 12348 7308 12404
rect 7364 12348 7868 12404
rect 7924 12348 9996 12404
rect 10052 12348 23100 12404
rect 23156 12348 23166 12404
rect 5954 12236 5964 12292
rect 6020 12236 6524 12292
rect 6580 12236 11452 12292
rect 11508 12236 17388 12292
rect 17444 12236 17454 12292
rect 35200 12180 36000 12208
rect 2034 12124 2044 12180
rect 2100 12124 3052 12180
rect 3108 12124 3118 12180
rect 4498 12124 4508 12180
rect 4564 12124 9212 12180
rect 9268 12124 9548 12180
rect 9604 12124 9614 12180
rect 11554 12124 11564 12180
rect 11620 12124 12348 12180
rect 12404 12124 12414 12180
rect 18946 12124 18956 12180
rect 19012 12124 21084 12180
rect 21140 12124 21150 12180
rect 24546 12124 24556 12180
rect 24612 12124 26908 12180
rect 26964 12124 26974 12180
rect 31892 12124 36000 12180
rect 19740 12068 19796 12124
rect 6850 12012 6860 12068
rect 6916 12012 7420 12068
rect 7476 12012 8316 12068
rect 8372 12012 8382 12068
rect 12002 12012 12012 12068
rect 12068 12012 13468 12068
rect 13524 12012 13534 12068
rect 19730 12012 19740 12068
rect 19796 12012 19806 12068
rect 20178 12012 20188 12068
rect 20244 12012 22596 12068
rect 31826 12012 31836 12068
rect 31892 12012 31948 12124
rect 35200 12096 36000 12124
rect 0 11956 800 11984
rect 0 11900 1932 11956
rect 1988 11900 1998 11956
rect 14242 11900 14252 11956
rect 14308 11900 15036 11956
rect 15092 11900 15102 11956
rect 20132 11900 21644 11956
rect 21700 11900 21710 11956
rect 0 11872 800 11900
rect 20132 11844 20188 11900
rect 14466 11788 14476 11844
rect 14532 11788 14924 11844
rect 14980 11788 19964 11844
rect 20020 11788 20188 11844
rect 20402 11788 20412 11844
rect 20468 11788 21532 11844
rect 21588 11788 21598 11844
rect 5360 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5644 11788
rect 13676 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13960 11788
rect 21992 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22276 11788
rect 22540 11732 22596 12012
rect 30308 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30592 11788
rect 12114 11676 12124 11732
rect 12180 11676 12908 11732
rect 12964 11676 12974 11732
rect 22530 11676 22540 11732
rect 22596 11676 22606 11732
rect 22866 11676 22876 11732
rect 22932 11676 26124 11732
rect 26180 11676 26190 11732
rect 28690 11676 28700 11732
rect 28756 11676 29596 11732
rect 29652 11676 29662 11732
rect 22876 11620 22932 11676
rect 18610 11564 18620 11620
rect 18676 11564 21924 11620
rect 22082 11564 22092 11620
rect 22148 11564 22932 11620
rect 29474 11564 29484 11620
rect 29540 11564 31164 11620
rect 31220 11564 31230 11620
rect 21868 11508 21924 11564
rect 11218 11452 11228 11508
rect 11284 11452 20076 11508
rect 20132 11452 20142 11508
rect 21868 11452 25004 11508
rect 25060 11452 25070 11508
rect 29810 11452 29820 11508
rect 29876 11452 30828 11508
rect 30884 11452 30894 11508
rect 3266 11340 3276 11396
rect 3332 11340 3836 11396
rect 3892 11340 3902 11396
rect 19618 11340 19628 11396
rect 19684 11340 20524 11396
rect 20580 11340 20590 11396
rect 21410 11340 21420 11396
rect 21476 11340 23100 11396
rect 23156 11340 23166 11396
rect 26674 11340 26684 11396
rect 26740 11340 27580 11396
rect 27636 11340 27646 11396
rect 11330 11228 11340 11284
rect 11396 11228 14364 11284
rect 14420 11228 14588 11284
rect 14644 11228 14654 11284
rect 14802 11228 14812 11284
rect 14868 11228 16044 11284
rect 16100 11228 16110 11284
rect 19170 11228 19180 11284
rect 19236 11228 21308 11284
rect 21364 11228 21374 11284
rect 22978 11228 22988 11284
rect 23044 11228 23884 11284
rect 23940 11228 24556 11284
rect 24612 11228 24622 11284
rect 14690 11116 14700 11172
rect 14756 11116 15820 11172
rect 15876 11116 15886 11172
rect 16594 11116 16604 11172
rect 16660 11116 17612 11172
rect 17668 11116 17678 11172
rect 21410 11116 21420 11172
rect 21476 11116 25900 11172
rect 25956 11116 25966 11172
rect 31892 11116 34300 11172
rect 34356 11116 34366 11172
rect 9518 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9802 11004
rect 17834 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18118 11004
rect 26150 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26434 11004
rect 28466 10892 28476 10948
rect 28532 10892 31836 10948
rect 31892 10892 31948 11116
rect 34466 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34750 11004
rect 15474 10780 15484 10836
rect 15540 10780 27916 10836
rect 27972 10780 27982 10836
rect 30818 10780 30828 10836
rect 30884 10780 31388 10836
rect 31444 10780 31454 10836
rect 12898 10668 12908 10724
rect 12964 10668 15372 10724
rect 15428 10668 15438 10724
rect 16370 10668 16380 10724
rect 16436 10668 18172 10724
rect 18228 10668 18238 10724
rect 23090 10668 23100 10724
rect 23156 10668 24556 10724
rect 24612 10668 25564 10724
rect 25620 10668 27020 10724
rect 27076 10668 27086 10724
rect 28018 10668 28028 10724
rect 28084 10668 33180 10724
rect 33236 10668 33246 10724
rect 35200 10612 36000 10640
rect 14354 10556 14364 10612
rect 14420 10556 18060 10612
rect 18116 10556 18126 10612
rect 20290 10556 20300 10612
rect 20356 10556 23548 10612
rect 23604 10556 24668 10612
rect 24724 10556 24734 10612
rect 28242 10556 28252 10612
rect 28308 10556 30380 10612
rect 30436 10556 30446 10612
rect 33506 10556 33516 10612
rect 33572 10556 36000 10612
rect 35200 10528 36000 10556
rect 16034 10444 16044 10500
rect 16100 10444 18396 10500
rect 18452 10444 20636 10500
rect 20692 10444 20702 10500
rect 20860 10444 25228 10500
rect 25284 10444 26012 10500
rect 26068 10444 26078 10500
rect 20860 10388 20916 10444
rect 18162 10332 18172 10388
rect 18228 10332 20916 10388
rect 21084 10332 22316 10388
rect 22372 10332 22382 10388
rect 21084 10276 21140 10332
rect 17378 10220 17388 10276
rect 17444 10220 18844 10276
rect 18900 10220 18910 10276
rect 20066 10220 20076 10276
rect 20132 10220 21140 10276
rect 5360 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5644 10220
rect 13676 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13960 10220
rect 21992 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22276 10220
rect 30308 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30592 10220
rect 15362 10108 15372 10164
rect 15428 10108 19180 10164
rect 19236 10108 19246 10164
rect 19954 10108 19964 10164
rect 20020 10108 21308 10164
rect 21364 10108 21374 10164
rect 22530 10108 22540 10164
rect 22596 10108 22876 10164
rect 22932 10108 24332 10164
rect 24388 10108 24398 10164
rect 14802 9996 14812 10052
rect 14868 9996 17724 10052
rect 17780 9996 19068 10052
rect 19124 9996 19134 10052
rect 19282 9996 19292 10052
rect 19348 9996 21756 10052
rect 21812 9996 21822 10052
rect 0 9940 800 9968
rect 0 9884 1932 9940
rect 1988 9884 1998 9940
rect 3266 9884 3276 9940
rect 3332 9884 3836 9940
rect 3892 9884 4732 9940
rect 4788 9884 4798 9940
rect 8306 9884 8316 9940
rect 8372 9884 25564 9940
rect 25620 9884 26460 9940
rect 26516 9884 26526 9940
rect 0 9856 800 9884
rect 6514 9772 6524 9828
rect 6580 9772 7980 9828
rect 8036 9772 8046 9828
rect 12786 9772 12796 9828
rect 12852 9772 14924 9828
rect 14980 9772 18284 9828
rect 18340 9772 18900 9828
rect 19058 9772 19068 9828
rect 19124 9772 20188 9828
rect 20244 9772 20254 9828
rect 20738 9772 20748 9828
rect 20804 9772 23660 9828
rect 23716 9772 23726 9828
rect 26338 9772 26348 9828
rect 26404 9772 26908 9828
rect 26964 9772 26974 9828
rect 18844 9716 18900 9772
rect 2930 9660 2940 9716
rect 2996 9660 4060 9716
rect 4116 9660 4126 9716
rect 14242 9660 14252 9716
rect 14308 9660 16268 9716
rect 16324 9660 16334 9716
rect 16706 9660 16716 9716
rect 16772 9660 17948 9716
rect 18004 9660 18620 9716
rect 18676 9660 18686 9716
rect 18844 9660 22764 9716
rect 22820 9660 22830 9716
rect 23874 9660 23884 9716
rect 23940 9660 25116 9716
rect 25172 9660 25182 9716
rect 26348 9604 26404 9772
rect 2706 9548 2716 9604
rect 2772 9548 6524 9604
rect 6580 9548 6590 9604
rect 14018 9548 14028 9604
rect 14084 9548 15596 9604
rect 15652 9548 15662 9604
rect 17266 9548 17276 9604
rect 17332 9548 19292 9604
rect 19348 9548 19358 9604
rect 21746 9548 21756 9604
rect 21812 9548 26404 9604
rect 32050 9548 32060 9604
rect 32116 9548 33404 9604
rect 33460 9548 33470 9604
rect 19170 9436 19180 9492
rect 19236 9436 23436 9492
rect 23492 9436 23502 9492
rect 9518 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9802 9436
rect 17834 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18118 9436
rect 26150 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26434 9436
rect 34466 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34750 9436
rect 5954 9212 5964 9268
rect 6020 9212 11452 9268
rect 11508 9212 11518 9268
rect 16594 9212 16604 9268
rect 16660 9212 17500 9268
rect 17556 9212 20524 9268
rect 20580 9212 29596 9268
rect 29652 9212 32620 9268
rect 32676 9212 32686 9268
rect 6514 9100 6524 9156
rect 6580 9100 7196 9156
rect 7252 9100 7262 9156
rect 25890 9100 25900 9156
rect 25956 9100 27244 9156
rect 27300 9100 27310 9156
rect 35200 9044 36000 9072
rect 3042 8988 3052 9044
rect 3108 8988 8316 9044
rect 8372 8988 8382 9044
rect 14354 8988 14364 9044
rect 14420 8988 15260 9044
rect 15316 8988 15326 9044
rect 16482 8988 16492 9044
rect 16548 8988 19180 9044
rect 19236 8988 19246 9044
rect 20514 8988 20524 9044
rect 20580 8988 22876 9044
rect 22932 8988 24556 9044
rect 24612 8988 24622 9044
rect 28578 8988 28588 9044
rect 28644 8988 29484 9044
rect 29540 8988 29550 9044
rect 32834 8988 32844 9044
rect 32900 8988 33404 9044
rect 33460 8988 33470 9044
rect 33954 8988 33964 9044
rect 34020 8988 36000 9044
rect 35200 8960 36000 8988
rect 1810 8876 1820 8932
rect 1876 8876 3948 8932
rect 4004 8876 4844 8932
rect 4900 8876 4910 8932
rect 7074 8876 7084 8932
rect 7140 8876 7756 8932
rect 7812 8876 12796 8932
rect 12852 8876 12862 8932
rect 15586 8876 15596 8932
rect 15652 8876 17388 8932
rect 17444 8876 17454 8932
rect 20402 8876 20412 8932
rect 20468 8876 24332 8932
rect 24388 8876 25788 8932
rect 25844 8876 25854 8932
rect 20290 8764 20300 8820
rect 20356 8764 21196 8820
rect 21252 8764 22596 8820
rect 26450 8764 26460 8820
rect 26516 8764 29484 8820
rect 29540 8764 29550 8820
rect 22540 8708 22596 8764
rect 22530 8652 22540 8708
rect 22596 8652 24220 8708
rect 24276 8652 28812 8708
rect 28868 8652 28878 8708
rect 5360 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5644 8652
rect 13676 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13960 8652
rect 21992 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22276 8652
rect 30308 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30592 8652
rect 26562 8428 26572 8484
rect 26628 8428 26908 8484
rect 26964 8428 26974 8484
rect 3490 8316 3500 8372
rect 3556 8316 6076 8372
rect 6132 8316 6142 8372
rect 9202 8316 9212 8372
rect 9268 8316 14028 8372
rect 14084 8316 14094 8372
rect 15092 8316 23380 8372
rect 23538 8316 23548 8372
rect 23604 8316 25788 8372
rect 25844 8316 25854 8372
rect 28466 8316 28476 8372
rect 28532 8316 29260 8372
rect 29316 8316 29326 8372
rect 2370 8204 2380 8260
rect 2436 8204 3836 8260
rect 3892 8204 4620 8260
rect 4676 8204 4686 8260
rect 13794 8204 13804 8260
rect 13860 8204 14476 8260
rect 14532 8204 14542 8260
rect 15092 8148 15148 8316
rect 15362 8204 15372 8260
rect 15428 8204 16716 8260
rect 16772 8204 20300 8260
rect 20356 8204 20366 8260
rect 23324 8148 23380 8316
rect 24658 8204 24668 8260
rect 24724 8204 25900 8260
rect 25956 8204 25966 8260
rect 12450 8092 12460 8148
rect 12516 8092 12796 8148
rect 12852 8092 15148 8148
rect 16940 8092 20076 8148
rect 20132 8092 21308 8148
rect 21364 8092 21374 8148
rect 23324 8092 25788 8148
rect 25844 8092 25854 8148
rect 26012 8092 29820 8148
rect 29876 8092 29886 8148
rect 4946 7980 4956 8036
rect 5012 7980 6636 8036
rect 6692 7980 6702 8036
rect 11218 7980 11228 8036
rect 11284 7980 11294 8036
rect 12898 7980 12908 8036
rect 12964 7980 13916 8036
rect 13972 7980 13982 8036
rect 0 7924 800 7952
rect 11228 7924 11284 7980
rect 16940 7924 16996 8092
rect 19730 7980 19740 8036
rect 19796 7980 20636 8036
rect 20692 7980 20702 8036
rect 0 7868 1932 7924
rect 1988 7868 1998 7924
rect 11228 7868 16996 7924
rect 19506 7868 19516 7924
rect 19572 7868 24780 7924
rect 24836 7868 24846 7924
rect 0 7840 800 7868
rect 9518 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9802 7868
rect 17834 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18118 7868
rect 26012 7812 26068 8092
rect 26226 7980 26236 8036
rect 26292 7980 26460 8036
rect 26516 7980 26526 8036
rect 26150 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26434 7868
rect 34466 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34750 7868
rect 18946 7756 18956 7812
rect 19012 7756 26068 7812
rect 12114 7644 12124 7700
rect 12180 7644 13020 7700
rect 13076 7644 13086 7700
rect 19282 7644 19292 7700
rect 19348 7644 31612 7700
rect 31668 7644 31678 7700
rect 5954 7532 5964 7588
rect 6020 7532 7196 7588
rect 7252 7532 11452 7588
rect 11508 7532 12012 7588
rect 12068 7532 12078 7588
rect 12898 7532 12908 7588
rect 12964 7532 13804 7588
rect 13860 7532 13870 7588
rect 17378 7532 17388 7588
rect 17444 7532 19516 7588
rect 19572 7532 19582 7588
rect 26562 7532 26572 7588
rect 26628 7532 27356 7588
rect 27412 7532 27422 7588
rect 35200 7476 36000 7504
rect 5842 7420 5852 7476
rect 5908 7420 6972 7476
rect 7028 7420 7038 7476
rect 13234 7420 13244 7476
rect 13300 7420 14140 7476
rect 14196 7420 15148 7476
rect 15204 7420 15214 7476
rect 21522 7420 21532 7476
rect 21588 7420 22204 7476
rect 22260 7420 22270 7476
rect 24770 7420 24780 7476
rect 24836 7420 29260 7476
rect 29316 7420 29326 7476
rect 31826 7420 31836 7476
rect 31892 7420 36000 7476
rect 35200 7392 36000 7420
rect 8418 7308 8428 7364
rect 8484 7308 13132 7364
rect 13188 7308 13198 7364
rect 22754 7308 22764 7364
rect 22820 7308 27692 7364
rect 27748 7308 27758 7364
rect 28466 7308 28476 7364
rect 28532 7308 32172 7364
rect 32228 7308 32238 7364
rect 28476 7252 28532 7308
rect 4722 7196 4732 7252
rect 4788 7196 15148 7252
rect 22082 7196 22092 7252
rect 22148 7196 22428 7252
rect 22484 7196 28532 7252
rect 28588 7196 34188 7252
rect 34244 7196 34254 7252
rect 5360 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5644 7084
rect 13676 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13960 7084
rect 2258 6972 2268 7028
rect 2324 6972 5068 7028
rect 5124 6972 5134 7028
rect 15092 6916 15148 7196
rect 28588 7140 28644 7196
rect 25218 7084 25228 7140
rect 25284 7084 26124 7140
rect 26180 7084 28644 7140
rect 21992 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22276 7084
rect 30308 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30592 7084
rect 16156 6972 18956 7028
rect 19012 6972 19740 7028
rect 19796 6972 19806 7028
rect 16156 6916 16212 6972
rect 2482 6860 2492 6916
rect 2548 6860 5628 6916
rect 5684 6860 5694 6916
rect 12562 6860 12572 6916
rect 12628 6860 13468 6916
rect 13524 6860 13534 6916
rect 15092 6860 16212 6916
rect 16370 6860 16380 6916
rect 16436 6860 17388 6916
rect 17444 6860 17454 6916
rect 29026 6860 29036 6916
rect 29092 6860 31948 6916
rect 33506 6860 33516 6916
rect 33572 6860 34076 6916
rect 34132 6860 34142 6916
rect 31892 6804 31948 6860
rect 2930 6748 2940 6804
rect 2996 6748 6300 6804
rect 6356 6748 6366 6804
rect 26786 6748 26796 6804
rect 26852 6748 28252 6804
rect 28308 6748 29596 6804
rect 29652 6748 29662 6804
rect 31892 6748 33852 6804
rect 33908 6748 33918 6804
rect 2146 6636 2156 6692
rect 2212 6636 7756 6692
rect 7812 6636 8316 6692
rect 8372 6636 8382 6692
rect 27122 6636 27132 6692
rect 27188 6636 27468 6692
rect 27524 6636 27534 6692
rect 27906 6636 27916 6692
rect 27972 6636 29932 6692
rect 29988 6636 29998 6692
rect 30146 6636 30156 6692
rect 30212 6636 31164 6692
rect 31220 6636 31230 6692
rect 7410 6524 7420 6580
rect 7476 6524 7980 6580
rect 8036 6524 8540 6580
rect 8596 6524 8606 6580
rect 15474 6524 15484 6580
rect 15540 6524 16604 6580
rect 16660 6524 16670 6580
rect 23202 6524 23212 6580
rect 23268 6524 26572 6580
rect 26628 6524 26638 6580
rect 28578 6524 28588 6580
rect 28644 6524 30268 6580
rect 30324 6524 31052 6580
rect 31108 6524 31118 6580
rect 32050 6524 32060 6580
rect 32116 6524 33516 6580
rect 33572 6524 33582 6580
rect 5170 6412 5180 6468
rect 5236 6412 10668 6468
rect 10724 6412 11116 6468
rect 11172 6412 11182 6468
rect 16930 6412 16940 6468
rect 16996 6412 19516 6468
rect 19572 6412 19582 6468
rect 27682 6412 27692 6468
rect 27748 6412 28364 6468
rect 28420 6412 28430 6468
rect 29586 6412 29596 6468
rect 29652 6412 31164 6468
rect 31220 6412 34300 6468
rect 34356 6412 34366 6468
rect 28690 6300 28700 6356
rect 28756 6300 30604 6356
rect 30660 6300 30670 6356
rect 9518 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9802 6300
rect 17834 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18118 6300
rect 26150 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26434 6300
rect 34466 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34750 6300
rect 9874 6188 9884 6244
rect 9940 6188 15260 6244
rect 15316 6188 15326 6244
rect 5730 6076 5740 6132
rect 5796 6076 6412 6132
rect 6468 6076 9660 6132
rect 9716 6076 9726 6132
rect 12226 6076 12236 6132
rect 12292 6076 12684 6132
rect 12740 6076 12750 6132
rect 14802 6076 14812 6132
rect 14868 6076 16940 6132
rect 16996 6076 17006 6132
rect 17714 6076 17724 6132
rect 17780 6076 18508 6132
rect 18564 6076 18574 6132
rect 31378 6076 31388 6132
rect 31444 6076 31836 6132
rect 31892 6076 32396 6132
rect 32452 6076 33180 6132
rect 33236 6076 33246 6132
rect 6850 5964 6860 6020
rect 6916 5964 10668 6020
rect 10724 5964 10734 6020
rect 13010 5964 13020 6020
rect 13076 5964 14028 6020
rect 14084 5964 14094 6020
rect 15586 5964 15596 6020
rect 15652 5964 16492 6020
rect 16548 5964 16558 6020
rect 18162 5964 18172 6020
rect 18228 5964 18620 6020
rect 18676 5964 19964 6020
rect 20020 5964 20030 6020
rect 26898 5964 26908 6020
rect 26964 5964 28700 6020
rect 28756 5964 28766 6020
rect 0 5908 800 5936
rect 35200 5908 36000 5936
rect 0 5852 2492 5908
rect 2548 5852 2558 5908
rect 6514 5852 6524 5908
rect 6580 5852 11788 5908
rect 11844 5852 11854 5908
rect 13234 5852 13244 5908
rect 13300 5852 13916 5908
rect 13972 5852 13982 5908
rect 16706 5852 16716 5908
rect 16772 5852 20188 5908
rect 20290 5852 20300 5908
rect 20356 5852 24444 5908
rect 24500 5852 24510 5908
rect 29250 5852 29260 5908
rect 29316 5852 29596 5908
rect 29652 5852 29662 5908
rect 34066 5852 34076 5908
rect 34132 5852 36000 5908
rect 0 5824 800 5852
rect 20132 5796 20188 5852
rect 35200 5824 36000 5852
rect 3938 5740 3948 5796
rect 4004 5740 7196 5796
rect 7252 5740 7262 5796
rect 8754 5740 8764 5796
rect 8820 5740 12684 5796
rect 12740 5740 12750 5796
rect 20132 5740 30940 5796
rect 30996 5740 31500 5796
rect 31556 5740 31566 5796
rect 33170 5740 33180 5796
rect 33236 5740 34188 5796
rect 34244 5740 34254 5796
rect 5954 5628 5964 5684
rect 6020 5628 9548 5684
rect 9604 5628 9614 5684
rect 18610 5628 18620 5684
rect 18676 5628 19740 5684
rect 19796 5628 20188 5684
rect 20244 5628 20254 5684
rect 26674 5628 26684 5684
rect 26740 5628 30772 5684
rect 31266 5628 31276 5684
rect 31332 5628 33740 5684
rect 33796 5628 33806 5684
rect 5360 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5644 5516
rect 13676 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13960 5516
rect 21992 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22276 5516
rect 30308 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30592 5516
rect 30716 5460 30772 5628
rect 30716 5404 33628 5460
rect 33684 5404 33694 5460
rect 7746 5292 7756 5348
rect 7812 5292 15148 5348
rect 15204 5292 16044 5348
rect 16100 5292 16604 5348
rect 16660 5292 16670 5348
rect 18162 5292 18172 5348
rect 18228 5292 19180 5348
rect 19236 5292 19246 5348
rect 25778 5292 25788 5348
rect 25844 5292 26796 5348
rect 26852 5292 26862 5348
rect 29474 5292 29484 5348
rect 29540 5292 32060 5348
rect 32116 5292 32126 5348
rect 4162 5180 4172 5236
rect 4228 5180 4732 5236
rect 4788 5180 6748 5236
rect 6804 5180 6814 5236
rect 20402 5180 20412 5236
rect 20468 5180 32844 5236
rect 32900 5180 32910 5236
rect 5618 5068 5628 5124
rect 5684 5068 7420 5124
rect 7476 5068 7486 5124
rect 28354 5068 28364 5124
rect 28420 5068 29988 5124
rect 33282 5068 33292 5124
rect 33348 5068 34188 5124
rect 34244 5068 34254 5124
rect 29932 5012 29988 5068
rect 8530 4956 8540 5012
rect 8596 4956 11564 5012
rect 11620 4956 11630 5012
rect 25890 4956 25900 5012
rect 25956 4956 26908 5012
rect 26964 4956 26974 5012
rect 29922 4956 29932 5012
rect 29988 4956 29998 5012
rect 9996 4900 10052 4956
rect 9986 4844 9996 4900
rect 10052 4844 10062 4900
rect 14018 4844 14028 4900
rect 14084 4844 16156 4900
rect 16212 4844 16222 4900
rect 17612 4844 18956 4900
rect 19012 4844 19022 4900
rect 22642 4844 22652 4900
rect 22708 4844 25116 4900
rect 25172 4844 25182 4900
rect 9518 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9802 4732
rect 17612 4676 17668 4844
rect 17834 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18118 4732
rect 26150 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26434 4732
rect 34466 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34750 4732
rect 10098 4620 10108 4676
rect 10164 4620 13692 4676
rect 13748 4620 17668 4676
rect 9874 4508 9884 4564
rect 9940 4508 10780 4564
rect 10836 4508 10846 4564
rect 19394 4508 19404 4564
rect 19460 4508 22652 4564
rect 22708 4508 22718 4564
rect 10994 4396 11004 4452
rect 11060 4396 12124 4452
rect 12180 4396 13132 4452
rect 13188 4396 13198 4452
rect 18386 4396 18396 4452
rect 18452 4396 20188 4452
rect 20132 4340 20188 4396
rect 35200 4340 36000 4368
rect 9090 4284 9100 4340
rect 9156 4284 11116 4340
rect 11172 4284 11900 4340
rect 11956 4284 11966 4340
rect 20132 4284 21644 4340
rect 21700 4284 21710 4340
rect 26450 4284 26460 4340
rect 26516 4284 28588 4340
rect 28644 4284 28654 4340
rect 32610 4284 32620 4340
rect 32676 4284 34076 4340
rect 34132 4284 34142 4340
rect 34290 4284 34300 4340
rect 34356 4284 36000 4340
rect 35200 4256 36000 4284
rect 5170 4172 5180 4228
rect 5236 4172 11564 4228
rect 11620 4172 11630 4228
rect 28466 4172 28476 4228
rect 28532 4172 33068 4228
rect 33124 4172 33134 4228
rect 1922 4060 1932 4116
rect 1988 4060 1998 4116
rect 0 3892 800 3920
rect 1932 3892 1988 4060
rect 5360 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5644 3948
rect 13676 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13960 3948
rect 21992 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22276 3948
rect 30308 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30592 3948
rect 0 3836 1988 3892
rect 0 3808 800 3836
rect 27570 3724 27580 3780
rect 27636 3724 34076 3780
rect 34132 3724 34142 3780
rect 8978 3612 8988 3668
rect 9044 3612 10332 3668
rect 10388 3612 10398 3668
rect 12562 3612 12572 3668
rect 12628 3612 14140 3668
rect 14196 3612 14206 3668
rect 19730 3612 19740 3668
rect 19796 3612 21868 3668
rect 21924 3612 21934 3668
rect 23314 3612 23324 3668
rect 23380 3612 25564 3668
rect 25620 3612 25630 3668
rect 26898 3612 26908 3668
rect 26964 3612 29372 3668
rect 29428 3612 29438 3668
rect 20066 3500 20076 3556
rect 20132 3500 20748 3556
rect 20804 3500 20814 3556
rect 26002 3500 26012 3556
rect 26068 3500 28588 3556
rect 28644 3500 28654 3556
rect 31714 3500 31724 3556
rect 31780 3500 33292 3556
rect 33348 3500 33358 3556
rect 5394 3388 5404 3444
rect 5460 3388 6636 3444
rect 6692 3388 6702 3444
rect 16146 3388 16156 3444
rect 16212 3388 18508 3444
rect 18564 3388 18574 3444
rect 32498 3388 32508 3444
rect 32564 3388 34188 3444
rect 34244 3388 34254 3444
rect 9518 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9802 3164
rect 17834 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18118 3164
rect 26150 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26434 3164
rect 34466 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34750 3164
rect 35200 2772 36000 2800
rect 34178 2716 34188 2772
rect 34244 2716 36000 2772
rect 35200 2688 36000 2716
rect 0 1876 800 1904
rect 0 1820 3388 1876
rect 3444 1820 3454 1876
rect 0 1792 800 1820
rect 35200 1204 36000 1232
rect 33282 1148 33292 1204
rect 33348 1148 36000 1204
rect 35200 1120 36000 1148
<< via3 >>
rect 5370 22708 5426 22764
rect 5474 22708 5530 22764
rect 5578 22708 5634 22764
rect 13686 22708 13742 22764
rect 13790 22708 13846 22764
rect 13894 22708 13950 22764
rect 22002 22708 22058 22764
rect 22106 22708 22162 22764
rect 22210 22708 22266 22764
rect 30318 22708 30374 22764
rect 30422 22708 30478 22764
rect 30526 22708 30582 22764
rect 9528 21924 9584 21980
rect 9632 21924 9688 21980
rect 9736 21924 9792 21980
rect 17844 21924 17900 21980
rect 17948 21924 18004 21980
rect 18052 21924 18108 21980
rect 26160 21924 26216 21980
rect 26264 21924 26320 21980
rect 26368 21924 26424 21980
rect 34476 21924 34532 21980
rect 34580 21924 34636 21980
rect 34684 21924 34740 21980
rect 5370 21140 5426 21196
rect 5474 21140 5530 21196
rect 5578 21140 5634 21196
rect 13686 21140 13742 21196
rect 13790 21140 13846 21196
rect 13894 21140 13950 21196
rect 22002 21140 22058 21196
rect 22106 21140 22162 21196
rect 22210 21140 22266 21196
rect 30318 21140 30374 21196
rect 30422 21140 30478 21196
rect 30526 21140 30582 21196
rect 9528 20356 9584 20412
rect 9632 20356 9688 20412
rect 9736 20356 9792 20412
rect 17844 20356 17900 20412
rect 17948 20356 18004 20412
rect 18052 20356 18108 20412
rect 26160 20356 26216 20412
rect 26264 20356 26320 20412
rect 26368 20356 26424 20412
rect 34476 20356 34532 20412
rect 34580 20356 34636 20412
rect 34684 20356 34740 20412
rect 5370 19572 5426 19628
rect 5474 19572 5530 19628
rect 5578 19572 5634 19628
rect 13686 19572 13742 19628
rect 13790 19572 13846 19628
rect 13894 19572 13950 19628
rect 22002 19572 22058 19628
rect 22106 19572 22162 19628
rect 22210 19572 22266 19628
rect 30318 19572 30374 19628
rect 30422 19572 30478 19628
rect 30526 19572 30582 19628
rect 9528 18788 9584 18844
rect 9632 18788 9688 18844
rect 9736 18788 9792 18844
rect 17844 18788 17900 18844
rect 17948 18788 18004 18844
rect 18052 18788 18108 18844
rect 26160 18788 26216 18844
rect 26264 18788 26320 18844
rect 26368 18788 26424 18844
rect 34476 18788 34532 18844
rect 34580 18788 34636 18844
rect 34684 18788 34740 18844
rect 5370 18004 5426 18060
rect 5474 18004 5530 18060
rect 5578 18004 5634 18060
rect 13686 18004 13742 18060
rect 13790 18004 13846 18060
rect 13894 18004 13950 18060
rect 22002 18004 22058 18060
rect 22106 18004 22162 18060
rect 22210 18004 22266 18060
rect 30318 18004 30374 18060
rect 30422 18004 30478 18060
rect 30526 18004 30582 18060
rect 9528 17220 9584 17276
rect 9632 17220 9688 17276
rect 9736 17220 9792 17276
rect 17844 17220 17900 17276
rect 17948 17220 18004 17276
rect 18052 17220 18108 17276
rect 26160 17220 26216 17276
rect 26264 17220 26320 17276
rect 26368 17220 26424 17276
rect 34476 17220 34532 17276
rect 34580 17220 34636 17276
rect 34684 17220 34740 17276
rect 5370 16436 5426 16492
rect 5474 16436 5530 16492
rect 5578 16436 5634 16492
rect 13686 16436 13742 16492
rect 13790 16436 13846 16492
rect 13894 16436 13950 16492
rect 22002 16436 22058 16492
rect 22106 16436 22162 16492
rect 22210 16436 22266 16492
rect 30318 16436 30374 16492
rect 30422 16436 30478 16492
rect 30526 16436 30582 16492
rect 9528 15652 9584 15708
rect 9632 15652 9688 15708
rect 9736 15652 9792 15708
rect 17844 15652 17900 15708
rect 17948 15652 18004 15708
rect 18052 15652 18108 15708
rect 26160 15652 26216 15708
rect 26264 15652 26320 15708
rect 26368 15652 26424 15708
rect 34476 15652 34532 15708
rect 34580 15652 34636 15708
rect 34684 15652 34740 15708
rect 5370 14868 5426 14924
rect 5474 14868 5530 14924
rect 5578 14868 5634 14924
rect 13686 14868 13742 14924
rect 13790 14868 13846 14924
rect 13894 14868 13950 14924
rect 22002 14868 22058 14924
rect 22106 14868 22162 14924
rect 22210 14868 22266 14924
rect 30318 14868 30374 14924
rect 30422 14868 30478 14924
rect 30526 14868 30582 14924
rect 9528 14084 9584 14140
rect 9632 14084 9688 14140
rect 9736 14084 9792 14140
rect 17844 14084 17900 14140
rect 17948 14084 18004 14140
rect 18052 14084 18108 14140
rect 26160 14084 26216 14140
rect 26264 14084 26320 14140
rect 26368 14084 26424 14140
rect 34476 14084 34532 14140
rect 34580 14084 34636 14140
rect 34684 14084 34740 14140
rect 5370 13300 5426 13356
rect 5474 13300 5530 13356
rect 5578 13300 5634 13356
rect 13686 13300 13742 13356
rect 13790 13300 13846 13356
rect 13894 13300 13950 13356
rect 22002 13300 22058 13356
rect 22106 13300 22162 13356
rect 22210 13300 22266 13356
rect 30318 13300 30374 13356
rect 30422 13300 30478 13356
rect 30526 13300 30582 13356
rect 20076 13132 20132 13188
rect 9528 12516 9584 12572
rect 9632 12516 9688 12572
rect 9736 12516 9792 12572
rect 17844 12516 17900 12572
rect 17948 12516 18004 12572
rect 18052 12516 18108 12572
rect 26160 12516 26216 12572
rect 26264 12516 26320 12572
rect 26368 12516 26424 12572
rect 34476 12516 34532 12572
rect 34580 12516 34636 12572
rect 34684 12516 34740 12572
rect 19964 11788 20020 11844
rect 5370 11732 5426 11788
rect 5474 11732 5530 11788
rect 5578 11732 5634 11788
rect 13686 11732 13742 11788
rect 13790 11732 13846 11788
rect 13894 11732 13950 11788
rect 22002 11732 22058 11788
rect 22106 11732 22162 11788
rect 22210 11732 22266 11788
rect 30318 11732 30374 11788
rect 30422 11732 30478 11788
rect 30526 11732 30582 11788
rect 9528 10948 9584 11004
rect 9632 10948 9688 11004
rect 9736 10948 9792 11004
rect 17844 10948 17900 11004
rect 17948 10948 18004 11004
rect 18052 10948 18108 11004
rect 26160 10948 26216 11004
rect 26264 10948 26320 11004
rect 26368 10948 26424 11004
rect 34476 10948 34532 11004
rect 34580 10948 34636 11004
rect 34684 10948 34740 11004
rect 20076 10220 20132 10276
rect 5370 10164 5426 10220
rect 5474 10164 5530 10220
rect 5578 10164 5634 10220
rect 13686 10164 13742 10220
rect 13790 10164 13846 10220
rect 13894 10164 13950 10220
rect 22002 10164 22058 10220
rect 22106 10164 22162 10220
rect 22210 10164 22266 10220
rect 30318 10164 30374 10220
rect 30422 10164 30478 10220
rect 30526 10164 30582 10220
rect 19964 10108 20020 10164
rect 19292 9996 19348 10052
rect 19292 9548 19348 9604
rect 9528 9380 9584 9436
rect 9632 9380 9688 9436
rect 9736 9380 9792 9436
rect 17844 9380 17900 9436
rect 17948 9380 18004 9436
rect 18052 9380 18108 9436
rect 26160 9380 26216 9436
rect 26264 9380 26320 9436
rect 26368 9380 26424 9436
rect 34476 9380 34532 9436
rect 34580 9380 34636 9436
rect 34684 9380 34740 9436
rect 5370 8596 5426 8652
rect 5474 8596 5530 8652
rect 5578 8596 5634 8652
rect 13686 8596 13742 8652
rect 13790 8596 13846 8652
rect 13894 8596 13950 8652
rect 22002 8596 22058 8652
rect 22106 8596 22162 8652
rect 22210 8596 22266 8652
rect 30318 8596 30374 8652
rect 30422 8596 30478 8652
rect 30526 8596 30582 8652
rect 9528 7812 9584 7868
rect 9632 7812 9688 7868
rect 9736 7812 9792 7868
rect 17844 7812 17900 7868
rect 17948 7812 18004 7868
rect 18052 7812 18108 7868
rect 26160 7812 26216 7868
rect 26264 7812 26320 7868
rect 26368 7812 26424 7868
rect 34476 7812 34532 7868
rect 34580 7812 34636 7868
rect 34684 7812 34740 7868
rect 5370 7028 5426 7084
rect 5474 7028 5530 7084
rect 5578 7028 5634 7084
rect 13686 7028 13742 7084
rect 13790 7028 13846 7084
rect 13894 7028 13950 7084
rect 22002 7028 22058 7084
rect 22106 7028 22162 7084
rect 22210 7028 22266 7084
rect 30318 7028 30374 7084
rect 30422 7028 30478 7084
rect 30526 7028 30582 7084
rect 9528 6244 9584 6300
rect 9632 6244 9688 6300
rect 9736 6244 9792 6300
rect 17844 6244 17900 6300
rect 17948 6244 18004 6300
rect 18052 6244 18108 6300
rect 26160 6244 26216 6300
rect 26264 6244 26320 6300
rect 26368 6244 26424 6300
rect 34476 6244 34532 6300
rect 34580 6244 34636 6300
rect 34684 6244 34740 6300
rect 5370 5460 5426 5516
rect 5474 5460 5530 5516
rect 5578 5460 5634 5516
rect 13686 5460 13742 5516
rect 13790 5460 13846 5516
rect 13894 5460 13950 5516
rect 22002 5460 22058 5516
rect 22106 5460 22162 5516
rect 22210 5460 22266 5516
rect 30318 5460 30374 5516
rect 30422 5460 30478 5516
rect 30526 5460 30582 5516
rect 9528 4676 9584 4732
rect 9632 4676 9688 4732
rect 9736 4676 9792 4732
rect 17844 4676 17900 4732
rect 17948 4676 18004 4732
rect 18052 4676 18108 4732
rect 26160 4676 26216 4732
rect 26264 4676 26320 4732
rect 26368 4676 26424 4732
rect 34476 4676 34532 4732
rect 34580 4676 34636 4732
rect 34684 4676 34740 4732
rect 5370 3892 5426 3948
rect 5474 3892 5530 3948
rect 5578 3892 5634 3948
rect 13686 3892 13742 3948
rect 13790 3892 13846 3948
rect 13894 3892 13950 3948
rect 22002 3892 22058 3948
rect 22106 3892 22162 3948
rect 22210 3892 22266 3948
rect 30318 3892 30374 3948
rect 30422 3892 30478 3948
rect 30526 3892 30582 3948
rect 9528 3108 9584 3164
rect 9632 3108 9688 3164
rect 9736 3108 9792 3164
rect 17844 3108 17900 3164
rect 17948 3108 18004 3164
rect 18052 3108 18108 3164
rect 26160 3108 26216 3164
rect 26264 3108 26320 3164
rect 26368 3108 26424 3164
rect 34476 3108 34532 3164
rect 34580 3108 34636 3164
rect 34684 3108 34740 3164
<< metal4 >>
rect 5342 22764 5662 22796
rect 5342 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5662 22764
rect 5342 21196 5662 22708
rect 5342 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5662 21196
rect 5342 19628 5662 21140
rect 5342 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5662 19628
rect 5342 18060 5662 19572
rect 5342 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5662 18060
rect 5342 16492 5662 18004
rect 5342 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5662 16492
rect 5342 14924 5662 16436
rect 5342 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5662 14924
rect 5342 13356 5662 14868
rect 5342 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5662 13356
rect 5342 11788 5662 13300
rect 5342 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5662 11788
rect 5342 10220 5662 11732
rect 5342 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5662 10220
rect 5342 8652 5662 10164
rect 5342 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5662 8652
rect 5342 7084 5662 8596
rect 5342 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5662 7084
rect 5342 5516 5662 7028
rect 5342 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5662 5516
rect 5342 3948 5662 5460
rect 5342 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5662 3948
rect 5342 3076 5662 3892
rect 9500 21980 9820 22796
rect 9500 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9820 21980
rect 9500 20412 9820 21924
rect 9500 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9820 20412
rect 9500 18844 9820 20356
rect 9500 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9820 18844
rect 9500 17276 9820 18788
rect 9500 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9820 17276
rect 9500 15708 9820 17220
rect 9500 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9820 15708
rect 9500 14140 9820 15652
rect 9500 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9820 14140
rect 9500 12572 9820 14084
rect 9500 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9820 12572
rect 9500 11004 9820 12516
rect 9500 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9820 11004
rect 9500 9436 9820 10948
rect 9500 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9820 9436
rect 9500 7868 9820 9380
rect 9500 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9820 7868
rect 9500 6300 9820 7812
rect 9500 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9820 6300
rect 9500 4732 9820 6244
rect 9500 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9820 4732
rect 9500 3164 9820 4676
rect 9500 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9820 3164
rect 9500 3076 9820 3108
rect 13658 22764 13978 22796
rect 13658 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13978 22764
rect 13658 21196 13978 22708
rect 13658 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13978 21196
rect 13658 19628 13978 21140
rect 13658 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13978 19628
rect 13658 18060 13978 19572
rect 13658 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13978 18060
rect 13658 16492 13978 18004
rect 13658 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13978 16492
rect 13658 14924 13978 16436
rect 13658 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13978 14924
rect 13658 13356 13978 14868
rect 13658 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13978 13356
rect 13658 11788 13978 13300
rect 13658 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13978 11788
rect 13658 10220 13978 11732
rect 13658 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13978 10220
rect 13658 8652 13978 10164
rect 13658 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13978 8652
rect 13658 7084 13978 8596
rect 13658 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13978 7084
rect 13658 5516 13978 7028
rect 13658 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13978 5516
rect 13658 3948 13978 5460
rect 13658 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13978 3948
rect 13658 3076 13978 3892
rect 17816 21980 18136 22796
rect 17816 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18136 21980
rect 17816 20412 18136 21924
rect 17816 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18136 20412
rect 17816 18844 18136 20356
rect 17816 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18136 18844
rect 17816 17276 18136 18788
rect 17816 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18136 17276
rect 17816 15708 18136 17220
rect 17816 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18136 15708
rect 17816 14140 18136 15652
rect 17816 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18136 14140
rect 17816 12572 18136 14084
rect 21974 22764 22294 22796
rect 21974 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22294 22764
rect 21974 21196 22294 22708
rect 21974 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22294 21196
rect 21974 19628 22294 21140
rect 21974 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22294 19628
rect 21974 18060 22294 19572
rect 21974 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22294 18060
rect 21974 16492 22294 18004
rect 21974 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22294 16492
rect 21974 14924 22294 16436
rect 21974 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22294 14924
rect 21974 13356 22294 14868
rect 21974 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22294 13356
rect 17816 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18136 12572
rect 17816 11004 18136 12516
rect 20076 13188 20132 13198
rect 17816 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18136 11004
rect 17816 9436 18136 10948
rect 19964 11844 20020 11854
rect 19964 10164 20020 11788
rect 20076 10276 20132 13132
rect 20076 10210 20132 10220
rect 21974 11788 22294 13300
rect 21974 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22294 11788
rect 21974 10220 22294 11732
rect 19964 10098 20020 10108
rect 21974 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22294 10220
rect 19292 10052 19348 10062
rect 19292 9604 19348 9996
rect 19292 9538 19348 9548
rect 17816 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18136 9436
rect 17816 7868 18136 9380
rect 17816 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18136 7868
rect 17816 6300 18136 7812
rect 17816 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18136 6300
rect 17816 4732 18136 6244
rect 17816 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18136 4732
rect 17816 3164 18136 4676
rect 17816 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18136 3164
rect 17816 3076 18136 3108
rect 21974 8652 22294 10164
rect 21974 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22294 8652
rect 21974 7084 22294 8596
rect 21974 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22294 7084
rect 21974 5516 22294 7028
rect 21974 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22294 5516
rect 21974 3948 22294 5460
rect 21974 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22294 3948
rect 21974 3076 22294 3892
rect 26132 21980 26452 22796
rect 26132 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26452 21980
rect 26132 20412 26452 21924
rect 26132 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26452 20412
rect 26132 18844 26452 20356
rect 26132 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26452 18844
rect 26132 17276 26452 18788
rect 26132 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26452 17276
rect 26132 15708 26452 17220
rect 26132 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26452 15708
rect 26132 14140 26452 15652
rect 26132 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26452 14140
rect 26132 12572 26452 14084
rect 26132 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26452 12572
rect 26132 11004 26452 12516
rect 26132 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26452 11004
rect 26132 9436 26452 10948
rect 26132 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26452 9436
rect 26132 7868 26452 9380
rect 26132 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26452 7868
rect 26132 6300 26452 7812
rect 26132 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26452 6300
rect 26132 4732 26452 6244
rect 26132 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26452 4732
rect 26132 3164 26452 4676
rect 26132 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26452 3164
rect 26132 3076 26452 3108
rect 30290 22764 30610 22796
rect 30290 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30610 22764
rect 30290 21196 30610 22708
rect 30290 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30610 21196
rect 30290 19628 30610 21140
rect 30290 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30610 19628
rect 30290 18060 30610 19572
rect 30290 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30610 18060
rect 30290 16492 30610 18004
rect 30290 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30610 16492
rect 30290 14924 30610 16436
rect 30290 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30610 14924
rect 30290 13356 30610 14868
rect 30290 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30610 13356
rect 30290 11788 30610 13300
rect 30290 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30610 11788
rect 30290 10220 30610 11732
rect 30290 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30610 10220
rect 30290 8652 30610 10164
rect 30290 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30610 8652
rect 30290 7084 30610 8596
rect 30290 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30610 7084
rect 30290 5516 30610 7028
rect 30290 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30610 5516
rect 30290 3948 30610 5460
rect 30290 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30610 3948
rect 30290 3076 30610 3892
rect 34448 21980 34768 22796
rect 34448 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34768 21980
rect 34448 20412 34768 21924
rect 34448 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34768 20412
rect 34448 18844 34768 20356
rect 34448 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34768 18844
rect 34448 17276 34768 18788
rect 34448 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34768 17276
rect 34448 15708 34768 17220
rect 34448 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34768 15708
rect 34448 14140 34768 15652
rect 34448 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34768 14140
rect 34448 12572 34768 14084
rect 34448 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34768 12572
rect 34448 11004 34768 12516
rect 34448 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34768 11004
rect 34448 9436 34768 10948
rect 34448 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34768 9436
rect 34448 7868 34768 9380
rect 34448 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34768 7868
rect 34448 6300 34768 7812
rect 34448 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34768 6300
rect 34448 4732 34768 6244
rect 34448 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34768 4732
rect 34448 3164 34768 4676
rect 34448 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34768 3164
rect 34448 3076 34768 3108
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _189_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 28224 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _190_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 3136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 4928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _192_
timestamp 1694700623
transform 1 0 29680 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _193_
timestamp 1694700623
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _194_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _195_
timestamp 1694700623
transform 1 0 28896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _196_
timestamp 1694700623
transform 1 0 29904 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _197_
timestamp 1694700623
transform 1 0 30240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _198_
timestamp 1694700623
transform -1 0 28896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _199_
timestamp 1694700623
transform -1 0 28224 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1694700623
transform 1 0 25760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _201_
timestamp 1694700623
transform -1 0 25984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _202_
timestamp 1694700623
transform -1 0 24640 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1694700623
transform 1 0 23296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _204_
timestamp 1694700623
transform -1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _205_
timestamp 1694700623
transform -1 0 25088 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _206_
timestamp 1694700623
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _207_
timestamp 1694700623
transform -1 0 20160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _208_
timestamp 1694700623
transform -1 0 19152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _209_
timestamp 1694700623
transform -1 0 17696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _210_
timestamp 1694700623
transform -1 0 18144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 13104 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _212_
timestamp 1694700623
transform 1 0 11984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _213_
timestamp 1694700623
transform 1 0 9632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1694700623
transform 1 0 10528 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _215_
timestamp 1694700623
transform -1 0 9184 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _216_
timestamp 1694700623
transform -1 0 9184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1694700623
transform 1 0 5488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _218_
timestamp 1694700623
transform -1 0 6608 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _219_
timestamp 1694700623
transform 1 0 12320 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _220_
timestamp 1694700623
transform -1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1694700623
transform 1 0 2464 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _222_
timestamp 1694700623
transform -1 0 3024 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _223_
timestamp 1694700623
transform -1 0 27776 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _224_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _225_
timestamp 1694700623
transform 1 0 19376 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _226_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22736 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _227_
timestamp 1694700623
transform 1 0 18144 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _228_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23856 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _229_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 24192 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _230_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 24192 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _231_
timestamp 1694700623
transform 1 0 18480 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _232_
timestamp 1694700623
transform -1 0 7392 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1694700623
transform -1 0 5152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _234_
timestamp 1694700623
transform -1 0 2464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _235_
timestamp 1694700623
transform -1 0 6496 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _236_
timestamp 1694700623
transform -1 0 2464 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _237_
timestamp 1694700623
transform -1 0 4928 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _238_
timestamp 1694700623
transform -1 0 12320 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _239_
timestamp 1694700623
transform -1 0 5376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _240_
timestamp 1694700623
transform -1 0 5376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _241_
timestamp 1694700623
transform -1 0 19936 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _242_
timestamp 1694700623
transform -1 0 19712 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _243_
timestamp 1694700623
transform 1 0 3136 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _244_
timestamp 1694700623
transform -1 0 12096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _245_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 3584 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _246_
timestamp 1694700623
transform 1 0 25424 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _247_
timestamp 1694700623
transform 1 0 24416 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _248_
timestamp 1694700623
transform 1 0 25088 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _249_
timestamp 1694700623
transform 1 0 18480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _250_
timestamp 1694700623
transform 1 0 18928 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _251_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 26992 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _252_
timestamp 1694700623
transform -1 0 30240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _253_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 28000 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _254_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23968 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _255_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 22736 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _256_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 28112 0 1 9408
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _257_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 25872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _258_
timestamp 1694700623
transform 1 0 27216 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _259_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 26432 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _260_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 28112 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _261_
timestamp 1694700623
transform -1 0 17920 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _262_
timestamp 1694700623
transform -1 0 31360 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _263_
timestamp 1694700623
transform -1 0 28784 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _264_
timestamp 1694700623
transform 1 0 29120 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _265_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 29232 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _266_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 21840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _267_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 19152 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _268_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21056 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _269_
timestamp 1694700623
transform 1 0 26320 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _270_
timestamp 1694700623
transform 1 0 22512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _271_
timestamp 1694700623
transform -1 0 23520 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _272_
timestamp 1694700623
transform 1 0 22176 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _273_
timestamp 1694700623
transform -1 0 26880 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _274_
timestamp 1694700623
transform -1 0 28784 0 -1 12544
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _275_
timestamp 1694700623
transform -1 0 25760 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _276_
timestamp 1694700623
transform -1 0 26432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _277_
timestamp 1694700623
transform 1 0 29008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _278_
timestamp 1694700623
transform 1 0 3136 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _279_
timestamp 1694700623
transform -1 0 22848 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _280_
timestamp 1694700623
transform -1 0 20832 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _281_
timestamp 1694700623
transform 1 0 20384 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _282_
timestamp 1694700623
transform 1 0 27664 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _283_
timestamp 1694700623
transform -1 0 29120 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _284_
timestamp 1694700623
transform 1 0 29008 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _285_
timestamp 1694700623
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _286_
timestamp 1694700623
transform 1 0 29120 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _287_
timestamp 1694700623
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _288_
timestamp 1694700623
transform 1 0 29792 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _289_
timestamp 1694700623
transform 1 0 28896 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _290_
timestamp 1694700623
transform 1 0 32928 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _291_
timestamp 1694700623
transform 1 0 26432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _292_
timestamp 1694700623
transform 1 0 25200 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _293_
timestamp 1694700623
transform -1 0 26880 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _294_
timestamp 1694700623
transform 1 0 27216 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _295_
timestamp 1694700623
transform -1 0 26880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _296_
timestamp 1694700623
transform 1 0 27328 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _297_
timestamp 1694700623
transform -1 0 25984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _298_
timestamp 1694700623
transform 1 0 30912 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _299_
timestamp 1694700623
transform -1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _300_
timestamp 1694700623
transform 1 0 29904 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _301_
timestamp 1694700623
transform -1 0 10528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _302_
timestamp 1694700623
transform -1 0 10080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _303_
timestamp 1694700623
transform -1 0 10192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _304_
timestamp 1694700623
transform -1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _305_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 28896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _306_
timestamp 1694700623
transform 1 0 20048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _307_
timestamp 1694700623
transform -1 0 21504 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _308_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 11424 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _309_
timestamp 1694700623
transform -1 0 24864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _310_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21728 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _311_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 24192 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _312_
timestamp 1694700623
transform -1 0 21056 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _313_
timestamp 1694700623
transform -1 0 18144 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _314_
timestamp 1694700623
transform 1 0 18480 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _315_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 17696 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _316_
timestamp 1694700623
transform 1 0 29008 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 28224 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _318_
timestamp 1694700623
transform -1 0 15008 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _319_
timestamp 1694700623
transform -1 0 15568 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _320_
timestamp 1694700623
transform 1 0 21504 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _321_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 19040 0 1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _322_
timestamp 1694700623
transform 1 0 15232 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_
timestamp 1694700623
transform 1 0 27776 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _324_
timestamp 1694700623
transform 1 0 16128 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _325_
timestamp 1694700623
transform -1 0 16464 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _326_
timestamp 1694700623
transform -1 0 15008 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _327_
timestamp 1694700623
transform -1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1694700623
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _329_
timestamp 1694700623
transform -1 0 17696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _330_
timestamp 1694700623
transform -1 0 14448 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _331_
timestamp 1694700623
transform 1 0 14336 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _332_
timestamp 1694700623
transform 1 0 14336 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _333_
timestamp 1694700623
transform 1 0 21168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _334_
timestamp 1694700623
transform 1 0 15120 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _335_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22176 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _336_
timestamp 1694700623
transform 1 0 23408 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _337_
timestamp 1694700623
transform 1 0 21840 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _338_
timestamp 1694700623
transform 1 0 22736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _339_
timestamp 1694700623
transform -1 0 20496 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _340_
timestamp 1694700623
transform -1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _341_
timestamp 1694700623
transform -1 0 19376 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _342_
timestamp 1694700623
transform -1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _343_
timestamp 1694700623
transform 1 0 19040 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _344_
timestamp 1694700623
transform 1 0 20048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _345_
timestamp 1694700623
transform 1 0 14672 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _346_
timestamp 1694700623
transform -1 0 19600 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _347_
timestamp 1694700623
transform -1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _348_
timestamp 1694700623
transform -1 0 19936 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _349_
timestamp 1694700623
transform 1 0 20160 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _350_
timestamp 1694700623
transform 1 0 19152 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _351_
timestamp 1694700623
transform 1 0 20384 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _352_
timestamp 1694700623
transform 1 0 14672 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _353_
timestamp 1694700623
transform -1 0 14672 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _354_
timestamp 1694700623
transform 1 0 14336 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _355_
timestamp 1694700623
transform -1 0 12320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _356_
timestamp 1694700623
transform -1 0 12096 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _357_
timestamp 1694700623
transform -1 0 11200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _358_
timestamp 1694700623
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _359_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 17024 0 -1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _360_
timestamp 1694700623
transform -1 0 15680 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _361_
timestamp 1694700623
transform -1 0 15008 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _362_
timestamp 1694700623
transform 1 0 11872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _363_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13328 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _364_
timestamp 1694700623
transform 1 0 11872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _365_
timestamp 1694700623
transform 1 0 12432 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _366_
timestamp 1694700623
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _367_
timestamp 1694700623
transform -1 0 13440 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _368_
timestamp 1694700623
transform -1 0 15008 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _369_
timestamp 1694700623
transform -1 0 14560 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _370_
timestamp 1694700623
transform 1 0 15792 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _371_
timestamp 1694700623
transform 1 0 15680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _372_
timestamp 1694700623
transform 1 0 15008 0 1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _373_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 23856 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _374_
timestamp 1694700623
transform -1 0 20944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _375_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21056 0 -1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _376_
timestamp 1694700623
transform -1 0 11424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _377_
timestamp 1694700623
transform 1 0 6608 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _378_
timestamp 1694700623
transform -1 0 6608 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _379_
timestamp 1694700623
transform -1 0 6496 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _380_
timestamp 1694700623
transform -1 0 6160 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _381_
timestamp 1694700623
transform -1 0 6944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _382_
timestamp 1694700623
transform -1 0 6832 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _383_
timestamp 1694700623
transform 1 0 10528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _384_
timestamp 1694700623
transform -1 0 10080 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _385_
timestamp 1694700623
transform -1 0 19936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _386_
timestamp 1694700623
transform 1 0 18928 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1694700623
transform 1 0 17920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _388_
timestamp 1694700623
transform -1 0 12656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _389_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 11088 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _390_
timestamp 1694700623
transform 1 0 11536 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _391_
timestamp 1694700623
transform -1 0 6160 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _392_
timestamp 1694700623
transform -1 0 6496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _393_
timestamp 1694700623
transform 1 0 6272 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _394_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 7840 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _395_
timestamp 1694700623
transform -1 0 20944 0 1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _396_
timestamp 1694700623
transform -1 0 11536 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _397_
timestamp 1694700623
transform 1 0 10416 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1694700623
transform 1 0 2464 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _399_
timestamp 1694700623
transform 1 0 6048 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _400_
timestamp 1694700623
transform 1 0 6384 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _401_
timestamp 1694700623
transform 1 0 7056 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _402_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 4368 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _403_
timestamp 1694700623
transform -1 0 7728 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _404_
timestamp 1694700623
transform 1 0 6720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _405_
timestamp 1694700623
transform 1 0 4032 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _406_
timestamp 1694700623
transform 1 0 3472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _407_
timestamp 1694700623
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _408_
timestamp 1694700623
transform 1 0 3584 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _409_
timestamp 1694700623
transform -1 0 7616 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _410_
timestamp 1694700623
transform 1 0 6160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _411_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 26208 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _412_
timestamp 1694700623
transform 1 0 30576 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _413_
timestamp 1694700623
transform 1 0 22064 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _414_
timestamp 1694700623
transform 1 0 22064 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _415_
timestamp 1694700623
transform 1 0 30576 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _416_
timestamp 1694700623
transform -1 0 34384 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _417_
timestamp 1694700623
transform -1 0 34384 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _418_
timestamp 1694700623
transform -1 0 34384 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _419_
timestamp 1694700623
transform -1 0 32816 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _420_
timestamp 1694700623
transform -1 0 34384 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _421_
timestamp 1694700623
transform -1 0 32704 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _422_
timestamp 1694700623
transform -1 0 30912 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _423_
timestamp 1694700623
transform 1 0 5824 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _424_
timestamp 1694700623
transform 1 0 5488 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _425_
timestamp 1694700623
transform 1 0 28896 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _426_
timestamp 1694700623
transform -1 0 31136 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _427_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15792 0 1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _428_
timestamp 1694700623
transform 1 0 13216 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _429_
timestamp 1694700623
transform 1 0 23856 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _430_
timestamp 1694700623
transform 1 0 22960 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _431_
timestamp 1694700623
transform 1 0 14784 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _432_
timestamp 1694700623
transform 1 0 19936 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _433_
timestamp 1694700623
transform 1 0 14784 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _434_
timestamp 1694700623
transform 1 0 20160 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _435_
timestamp 1694700623
transform 1 0 20944 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _436_
timestamp 1694700623
transform 1 0 13216 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _437_
timestamp 1694700623
transform 1 0 10528 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _438_
timestamp 1694700623
transform 1 0 9968 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _439_
timestamp 1694700623
transform 1 0 8512 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _440_
timestamp 1694700623
transform 1 0 7728 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _441_
timestamp 1694700623
transform 1 0 7952 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _442_
timestamp 1694700623
transform -1 0 16912 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _443_
timestamp 1694700623
transform 1 0 16016 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _444_
timestamp 1694700623
transform 1 0 2800 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _445_
timestamp 1694700623
transform 1 0 1792 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _446_
timestamp 1694700623
transform 1 0 2240 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _447_
timestamp 1694700623
transform 1 0 5376 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _448_
timestamp 1694700623
transform -1 0 22400 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _449_
timestamp 1694700623
transform 1 0 7728 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _450_ pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 12544
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _451_
timestamp 1694700623
transform -1 0 14336 0 -1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _452_
timestamp 1694700623
transform -1 0 5600 0 -1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _453_
timestamp 1694700623
transform 1 0 6272 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 3360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1694700623
transform 1 0 6720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1694700623
transform -1 0 32256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1694700623
transform 1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1694700623
transform -1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1694700623
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1694700623
transform 1 0 20272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1694700623
transform 1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__A2
timestamp 1694700623
transform 1 0 9632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__A2
timestamp 1694700623
transform 1 0 7504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__I
timestamp 1694700623
transform 1 0 4704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__I
timestamp 1694700623
transform 1 0 5600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__I
timestamp 1694700623
transform 1 0 3808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__A2
timestamp 1694700623
transform 1 0 27216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A1
timestamp 1694700623
transform -1 0 25872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__B
timestamp 1694700623
transform 1 0 26992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__277__I
timestamp 1694700623
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A1
timestamp 1694700623
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I
timestamp 1694700623
transform 1 0 27440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1694700623
transform 1 0 23968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A2
timestamp 1694700623
transform -1 0 10976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A1
timestamp 1694700623
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A2
timestamp 1694700623
transform 1 0 10416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__B
timestamp 1694700623
transform 1 0 10864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A1
timestamp 1694700623
transform 1 0 9632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__B
timestamp 1694700623
transform 1 0 12320 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__I
timestamp 1694700623
transform 1 0 12432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__A2
timestamp 1694700623
transform -1 0 20384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1694700623
transform 1 0 23072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A1
timestamp 1694700623
transform 1 0 7728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__A2
timestamp 1694700623
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A1
timestamp 1694700623
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1694700623
transform -1 0 6944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A3
timestamp 1694700623
transform 1 0 7616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__B
timestamp 1694700623
transform 1 0 21392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A1
timestamp 1694700623
transform -1 0 3472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1694700623
transform -1 0 7616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A2
timestamp 1694700623
transform -1 0 7168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A1
timestamp 1694700623
transform 1 0 7840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A2
timestamp 1694700623
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__RN
timestamp 1694700623
transform 1 0 25872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__RN
timestamp 1694700623
transform 1 0 26096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__CLK
timestamp 1694700623
transform 1 0 31360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__RN
timestamp 1694700623
transform 1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout52_I
timestamp 1694700623
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout55_I
timestamp 1694700623
transform 1 0 12320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout56_I
timestamp 1694700623
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout58_I
timestamp 1694700623
transform -1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout76_I
timestamp 1694700623
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout79_I
timestamp 1694700623
transform 1 0 29792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout80_I
timestamp 1694700623
transform 1 0 24080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1694700623
transform -1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1694700623
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1694700623
transform 1 0 1792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1694700623
transform -1 0 33488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1694700623
transform -1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1694700623
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1694700623
transform -1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1694700623
transform 1 0 6048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1694700623
transform -1 0 33376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1694700623
transform 1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1694700623
transform 1 0 31360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1694700623
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1694700623
transform 1 0 23744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1694700623
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1694700623
transform 1 0 28672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1694700623
transform 1 0 7168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1694700623
transform 1 0 4704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1694700623
transform 1 0 4704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout49
timestamp 1694700623
transform -1 0 11872 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout50
timestamp 1694700623
transform -1 0 10528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout51
timestamp 1694700623
transform -1 0 10080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout52
timestamp 1694700623
transform 1 0 18368 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout53
timestamp 1694700623
transform -1 0 19712 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout54
timestamp 1694700623
transform -1 0 18704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout55
timestamp 1694700623
transform -1 0 11648 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout56
timestamp 1694700623
transform -1 0 20384 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout57
timestamp 1694700623
transform -1 0 20608 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout58
timestamp 1694700623
transform -1 0 34384 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout59
timestamp 1694700623
transform 1 0 33488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout60
timestamp 1694700623
transform -1 0 34384 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout61
timestamp 1694700623
transform -1 0 34384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout62
timestamp 1694700623
transform 1 0 33488 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout63
timestamp 1694700623
transform -1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout64
timestamp 1694700623
transform -1 0 33712 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1694700623
transform -1 0 34384 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1694700623
transform -1 0 8848 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout67
timestamp 1694700623
transform 1 0 7840 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout68
timestamp 1694700623
transform -1 0 7952 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout69
timestamp 1694700623
transform -1 0 15680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout70
timestamp 1694700623
transform -1 0 16128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout71
timestamp 1694700623
transform -1 0 14784 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout72
timestamp 1694700623
transform -1 0 8624 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout73
timestamp 1694700623
transform -1 0 16800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout74
timestamp 1694700623
transform -1 0 17024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout75
timestamp 1694700623
transform 1 0 28224 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout76
timestamp 1694700623
transform -1 0 32704 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout77
timestamp 1694700623
transform -1 0 33488 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout78
timestamp 1694700623
transform -1 0 34272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout79
timestamp 1694700623
transform -1 0 29792 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout80
timestamp 1694700623
transform -1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout81
timestamp 1694700623
transform 1 0 31360 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout82
timestamp 1694700623
transform -1 0 31472 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_4 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1792 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_31
timestamp 1694700623
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1694700623
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_36
timestamp 1694700623
transform 1 0 5376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_63
timestamp 1694700623
transform 1 0 8400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_65
timestamp 1694700623
transform 1 0 8624 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_96 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 12096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_130
timestamp 1694700623
transform 1 0 15904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1694700623
transform 1 0 16352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_164
timestamp 1694700623
transform 1 0 19712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1694700623
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1694700623
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1694700623
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1694700623
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1694700623
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1694700623
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1694700623
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_276
timestamp 1694700623
transform 1 0 32256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_279
timestamp 1694700623
transform 1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1694700623
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_98
timestamp 1694700623
transform 1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_102
timestamp 1694700623
transform 1 0 12768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_104
timestamp 1694700623
transform 1 0 12992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1694700623
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1694700623
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_188
timestamp 1694700623
transform 1 0 22400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_192
timestamp 1694700623
transform 1 0 22848 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_200
timestamp 1694700623
transform 1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_204
timestamp 1694700623
transform 1 0 24192 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1694700623
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1694700623
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_256
timestamp 1694700623
transform 1 0 30016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_262
timestamp 1694700623
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_266 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 31136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_276
timestamp 1694700623
transform 1 0 32256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_286
timestamp 1694700623
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_288
timestamp 1694700623
transform 1 0 33600 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_32
timestamp 1694700623
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1694700623
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_37
timestamp 1694700623
transform 1 0 5488 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_46
timestamp 1694700623
transform 1 0 6496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_50
timestamp 1694700623
transform 1 0 6944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_52
timestamp 1694700623
transform 1 0 7168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_93
timestamp 1694700623
transform 1 0 11760 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1694700623
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_111 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13776 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_127
timestamp 1694700623
transform 1 0 15568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_165
timestamp 1694700623
transform 1 0 19824 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1694700623
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1694700623
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1694700623
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_258
timestamp 1694700623
transform 1 0 30240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_260
timestamp 1694700623
transform 1 0 30464 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2
timestamp 1694700623
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_6
timestamp 1694700623
transform 1 0 2016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_50
timestamp 1694700623
transform 1 0 6944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_54
timestamp 1694700623
transform 1 0 7392 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_58
timestamp 1694700623
transform 1 0 7840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_60
timestamp 1694700623
transform 1 0 8064 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_67
timestamp 1694700623
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1694700623
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_78
timestamp 1694700623
transform 1 0 10080 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_142
timestamp 1694700623
transform 1 0 17248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_148
timestamp 1694700623
transform 1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_172 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20608 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_204
timestamp 1694700623
transform 1 0 24192 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1694700623
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_212
timestamp 1694700623
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_216
timestamp 1694700623
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_218
timestamp 1694700623
transform 1 0 25760 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_221
timestamp 1694700623
transform 1 0 26096 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_237
timestamp 1694700623
transform 1 0 27888 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1694700623
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_286
timestamp 1694700623
transform 1 0 33376 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_28
timestamp 1694700623
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1694700623
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1694700623
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_49
timestamp 1694700623
transform 1 0 6832 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_91
timestamp 1694700623
transform 1 0 11536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1694700623
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1694700623
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1694700623
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_123
timestamp 1694700623
transform 1 0 15120 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_127
timestamp 1694700623
transform 1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_144
timestamp 1694700623
transform 1 0 17472 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_152
timestamp 1694700623
transform 1 0 18368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_156
timestamp 1694700623
transform 1 0 18816 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1694700623
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1694700623
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_177
timestamp 1694700623
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_185
timestamp 1694700623
transform 1 0 22064 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_197
timestamp 1694700623
transform 1 0 23408 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_213
timestamp 1694700623
transform 1 0 25200 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_221
timestamp 1694700623
transform 1 0 26096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1694700623
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1694700623
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_54
timestamp 1694700623
transform 1 0 7392 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_72
timestamp 1694700623
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_88
timestamp 1694700623
transform 1 0 11200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_92
timestamp 1694700623
transform 1 0 11648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_98
timestamp 1694700623
transform 1 0 12320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_109
timestamp 1694700623
transform 1 0 13552 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_117
timestamp 1694700623
transform 1 0 14448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_121
timestamp 1694700623
transform 1 0 14896 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_128
timestamp 1694700623
transform 1 0 15680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1694700623
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_148
timestamp 1694700623
transform 1 0 17920 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_164
timestamp 1694700623
transform 1 0 19712 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_172
timestamp 1694700623
transform 1 0 20608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_181
timestamp 1694700623
transform 1 0 21616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_185
timestamp 1694700623
transform 1 0 22064 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_198
timestamp 1694700623
transform 1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1694700623
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1694700623
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1694700623
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_219
timestamp 1694700623
transform 1 0 25872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_223
timestamp 1694700623
transform 1 0 26320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_237
timestamp 1694700623
transform 1 0 27888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_239
timestamp 1694700623
transform 1 0 28112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1694700623
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_284
timestamp 1694700623
transform 1 0 33152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1694700623
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_37
timestamp 1694700623
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_47
timestamp 1694700623
transform 1 0 6608 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_79
timestamp 1694700623
transform 1 0 10192 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_83
timestamp 1694700623
transform 1 0 10640 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_90
timestamp 1694700623
transform 1 0 11424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_98
timestamp 1694700623
transform 1 0 12320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_166
timestamp 1694700623
transform 1 0 19936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_170
timestamp 1694700623
transform 1 0 20384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1694700623
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1694700623
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_227
timestamp 1694700623
transform 1 0 26768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_231
timestamp 1694700623
transform 1 0 27216 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1694700623
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1694700623
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_262
timestamp 1694700623
transform 1 0 30688 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_10
timestamp 1694700623
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_12
timestamp 1694700623
transform 1 0 2688 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_55
timestamp 1694700623
transform 1 0 7504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_59
timestamp 1694700623
transform 1 0 7952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1694700623
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1694700623
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1694700623
transform 1 0 9408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_104
timestamp 1694700623
transform 1 0 12992 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_120
timestamp 1694700623
transform 1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_122
timestamp 1694700623
transform 1 0 15008 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_146
timestamp 1694700623
transform 1 0 17696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_150
timestamp 1694700623
transform 1 0 18144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_152
timestamp 1694700623
transform 1 0 18368 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_162
timestamp 1694700623
transform 1 0 19488 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_195
timestamp 1694700623
transform 1 0 23184 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_199
timestamp 1694700623
transform 1 0 23632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_201
timestamp 1694700623
transform 1 0 23856 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1694700623
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1694700623
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_229
timestamp 1694700623
transform 1 0 26992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_233
timestamp 1694700623
transform 1 0 27440 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_237
timestamp 1694700623
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_239
timestamp 1694700623
transform 1 0 28112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1694700623
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1694700623
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_20
timestamp 1694700623
transform 1 0 3584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_24
timestamp 1694700623
transform 1 0 4032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1694700623
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1694700623
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1694700623
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1694700623
transform 1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_57
timestamp 1694700623
transform 1 0 7728 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1694700623
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1694700623
transform 1 0 13328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_127
timestamp 1694700623
transform 1 0 15568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_131
timestamp 1694700623
transform 1 0 16016 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_138
timestamp 1694700623
transform 1 0 16800 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_156
timestamp 1694700623
transform 1 0 18816 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_164
timestamp 1694700623
transform 1 0 19712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_166
timestamp 1694700623
transform 1 0 19936 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_204
timestamp 1694700623
transform 1 0 24192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_239
timestamp 1694700623
transform 1 0 28112 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1694700623
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_247
timestamp 1694700623
transform 1 0 29008 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_263
timestamp 1694700623
transform 1 0 30800 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_267
timestamp 1694700623
transform 1 0 31248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_28
timestamp 1694700623
transform 1 0 4480 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_60
timestamp 1694700623
transform 1 0 8064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1694700623
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1694700623
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1694700623
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_105
timestamp 1694700623
transform 1 0 13104 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_113
timestamp 1694700623
transform 1 0 14000 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_122
timestamp 1694700623
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1694700623
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1694700623
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_164
timestamp 1694700623
transform 1 0 19712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_166
timestamp 1694700623
transform 1 0 19936 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1694700623
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_214
timestamp 1694700623
transform 1 0 25312 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_223
timestamp 1694700623
transform 1 0 26320 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_231
timestamp 1694700623
transform 1 0 27216 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_266
timestamp 1694700623
transform 1 0 31136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_270
timestamp 1694700623
transform 1 0 31584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1694700623
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1694700623
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1694700623
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1694700623
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1694700623
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1694700623
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1694700623
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1694700623
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1694700623
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_43
timestamp 1694700623
transform 1 0 6160 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_78
timestamp 1694700623
transform 1 0 10080 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_94
timestamp 1694700623
transform 1 0 11872 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1694700623
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1694700623
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1694700623
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_115
timestamp 1694700623
transform 1 0 14224 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1694700623
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_181
timestamp 1694700623
transform 1 0 21616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_204
timestamp 1694700623
transform 1 0 24192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_214
timestamp 1694700623
transform 1 0 25312 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_218
timestamp 1694700623
transform 1 0 25760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1694700623
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1694700623
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1694700623
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1694700623
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_253
timestamp 1694700623
transform 1 0 29680 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_256
timestamp 1694700623
transform 1 0 30016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_260
timestamp 1694700623
transform 1 0 30464 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_56
timestamp 1694700623
transform 1 0 7616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_60
timestamp 1694700623
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_64
timestamp 1694700623
transform 1 0 8512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1694700623
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_78
timestamp 1694700623
transform 1 0 10080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_86
timestamp 1694700623
transform 1 0 10976 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_101
timestamp 1694700623
transform 1 0 12656 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_109
timestamp 1694700623
transform 1 0 13552 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_113
timestamp 1694700623
transform 1 0 14000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_115
timestamp 1694700623
transform 1 0 14224 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_124
timestamp 1694700623
transform 1 0 15232 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_128
timestamp 1694700623
transform 1 0 15680 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_135
timestamp 1694700623
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1694700623
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1694700623
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1694700623
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_152
timestamp 1694700623
transform 1 0 18368 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1694700623
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_245
timestamp 1694700623
transform 1 0 28784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_247
timestamp 1694700623
transform 1 0 29008 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_282
timestamp 1694700623
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_286
timestamp 1694700623
transform 1 0 33376 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1694700623
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_20
timestamp 1694700623
transform 1 0 3584 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1694700623
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1694700623
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1694700623
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_37
timestamp 1694700623
transform 1 0 5488 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_46
timestamp 1694700623
transform 1 0 6496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_50
timestamp 1694700623
transform 1 0 6944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_54
timestamp 1694700623
transform 1 0 7392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_56
timestamp 1694700623
transform 1 0 7616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1694700623
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_113
timestamp 1694700623
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_115
timestamp 1694700623
transform 1 0 14224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_124
timestamp 1694700623
transform 1 0 15232 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_136
timestamp 1694700623
transform 1 0 16576 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_152
timestamp 1694700623
transform 1 0 18368 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_165
timestamp 1694700623
transform 1 0 19824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_192
timestamp 1694700623
transform 1 0 22848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_196
timestamp 1694700623
transform 1 0 23296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_210
timestamp 1694700623
transform 1 0 24864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_220
timestamp 1694700623
transform 1 0 25984 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_236
timestamp 1694700623
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1694700623
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1694700623
transform 1 0 1568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_6
timestamp 1694700623
transform 1 0 2016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_16
timestamp 1694700623
transform 1 0 3136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_43
timestamp 1694700623
transform 1 0 6160 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_48
timestamp 1694700623
transform 1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_52
timestamp 1694700623
transform 1 0 7168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_56
timestamp 1694700623
transform 1 0 7616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_58
timestamp 1694700623
transform 1 0 7840 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_65
timestamp 1694700623
transform 1 0 8624 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1694700623
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1694700623
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1694700623
transform 1 0 10304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1694700623
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_100
timestamp 1694700623
transform 1 0 12544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1694700623
transform 1 0 12992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1694700623
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_158
timestamp 1694700623
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_160
timestamp 1694700623
transform 1 0 19264 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_167
timestamp 1694700623
transform 1 0 20048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_169
timestamp 1694700623
transform 1 0 20272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1694700623
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1694700623
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_228
timestamp 1694700623
transform 1 0 26880 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1694700623
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1694700623
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_8
timestamp 1694700623
transform 1 0 2240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1694700623
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1694700623
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_50
timestamp 1694700623
transform 1 0 6944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_54
timestamp 1694700623
transform 1 0 7392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_81
timestamp 1694700623
transform 1 0 10416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_91
timestamp 1694700623
transform 1 0 11536 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_99
timestamp 1694700623
transform 1 0 12432 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1694700623
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1694700623
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1694700623
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1694700623
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_165
timestamp 1694700623
transform 1 0 19824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_167
timestamp 1694700623
transform 1 0 20048 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1694700623
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1694700623
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_181
timestamp 1694700623
transform 1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_185
timestamp 1694700623
transform 1 0 22064 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_195
timestamp 1694700623
transform 1 0 23184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_235
timestamp 1694700623
transform 1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1694700623
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_263
timestamp 1694700623
transform 1 0 30800 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_267
timestamp 1694700623
transform 1 0 31248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_2
timestamp 1694700623
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_10
timestamp 1694700623
transform 1 0 2464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_14
timestamp 1694700623
transform 1 0 2912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_16
timestamp 1694700623
transform 1 0 3136 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_59
timestamp 1694700623
transform 1 0 7952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1694700623
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1694700623
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1694700623
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_116
timestamp 1694700623
transform 1 0 14336 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1694700623
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1694700623
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1694700623
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1694700623
transform 1 0 18144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1694700623
transform 1 0 18592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_180
timestamp 1694700623
transform 1 0 21504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1694700623
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_190
timestamp 1694700623
transform 1 0 22624 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_201
timestamp 1694700623
transform 1 0 23856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1694700623
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1694700623
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1694700623
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_228
timestamp 1694700623
transform 1 0 26880 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_232
timestamp 1694700623
transform 1 0 27328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_235
timestamp 1694700623
transform 1 0 27664 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_243
timestamp 1694700623
transform 1 0 28560 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_282
timestamp 1694700623
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_290
timestamp 1694700623
transform 1 0 33824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_294
timestamp 1694700623
transform 1 0 34272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_28
timestamp 1694700623
transform 1 0 4480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1694700623
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1694700623
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1694700623
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1694700623
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_48
timestamp 1694700623
transform 1 0 6720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_50
timestamp 1694700623
transform 1 0 6944 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_57
timestamp 1694700623
transform 1 0 7728 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_73
timestamp 1694700623
transform 1 0 9520 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_89
timestamp 1694700623
transform 1 0 11312 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1694700623
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1694700623
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1694700623
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_154
timestamp 1694700623
transform 1 0 18592 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1694700623
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1694700623
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_192
timestamp 1694700623
transform 1 0 22848 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1694700623
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_255
timestamp 1694700623
transform 1 0 29904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_259
timestamp 1694700623
transform 1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_38
timestamp 1694700623
transform 1 0 5600 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_46
timestamp 1694700623
transform 1 0 6496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_56
timestamp 1694700623
transform 1 0 7616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1694700623
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1694700623
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1694700623
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1694700623
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_120
timestamp 1694700623
transform 1 0 14784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1694700623
transform 1 0 15008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1694700623
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1694700623
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1694700623
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1694700623
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1694700623
transform 1 0 18144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_161
timestamp 1694700623
transform 1 0 19376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_165
timestamp 1694700623
transform 1 0 19824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_200
timestamp 1694700623
transform 1 0 23744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1694700623
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_218
timestamp 1694700623
transform 1 0 25760 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_226
timestamp 1694700623
transform 1 0 26656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_230
timestamp 1694700623
transform 1 0 27104 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_237
timestamp 1694700623
transform 1 0 27888 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1694700623
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_286
timestamp 1694700623
transform 1 0 33376 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1694700623
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1694700623
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1694700623
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_53
timestamp 1694700623
transform 1 0 7280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_61
timestamp 1694700623
transform 1 0 8176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_65
timestamp 1694700623
transform 1 0 8624 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_72
timestamp 1694700623
transform 1 0 9408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_76
timestamp 1694700623
transform 1 0 9856 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_96
timestamp 1694700623
transform 1 0 12096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_100
timestamp 1694700623
transform 1 0 12544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1694700623
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1694700623
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_139
timestamp 1694700623
transform 1 0 16912 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_155
timestamp 1694700623
transform 1 0 18704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_157
timestamp 1694700623
transform 1 0 18928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1694700623
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_177
timestamp 1694700623
transform 1 0 21168 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_209
timestamp 1694700623
transform 1 0 24752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_217
timestamp 1694700623
transform 1 0 25648 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_230
timestamp 1694700623
transform 1 0 27104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_240
timestamp 1694700623
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1694700623
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_253
timestamp 1694700623
transform 1 0 29680 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_260
timestamp 1694700623
transform 1 0 30464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_28
timestamp 1694700623
transform 1 0 4480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_36
timestamp 1694700623
transform 1 0 5376 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_47
timestamp 1694700623
transform 1 0 6608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_55
timestamp 1694700623
transform 1 0 7504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_59
timestamp 1694700623
transform 1 0 7952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_61
timestamp 1694700623
transform 1 0 8176 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1694700623
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_76
timestamp 1694700623
transform 1 0 9856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_111
timestamp 1694700623
transform 1 0 13776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_125
timestamp 1694700623
transform 1 0 15344 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_129
timestamp 1694700623
transform 1 0 15792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1694700623
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1694700623
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1694700623
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1694700623
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_155
timestamp 1694700623
transform 1 0 18704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_163
timestamp 1694700623
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_171
timestamp 1694700623
transform 1 0 20496 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_187
timestamp 1694700623
transform 1 0 22288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_195
timestamp 1694700623
transform 1 0 23184 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_199
timestamp 1694700623
transform 1 0 23632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1694700623
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_294
timestamp 1694700623
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1694700623
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_10
timestamp 1694700623
transform 1 0 2464 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_15
timestamp 1694700623
transform 1 0 3024 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1694700623
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_79
timestamp 1694700623
transform 1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_83
timestamp 1694700623
transform 1 0 10640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_87
timestamp 1694700623
transform 1 0 11088 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_91
timestamp 1694700623
transform 1 0 11536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_93
timestamp 1694700623
transform 1 0 11760 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_98
timestamp 1694700623
transform 1 0 12320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1694700623
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1694700623
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1694700623
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1694700623
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_113
timestamp 1694700623
transform 1 0 14000 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1694700623
transform 1 0 20272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1694700623
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1694700623
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_193
timestamp 1694700623
transform 1 0 22960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_201
timestamp 1694700623
transform 1 0 23856 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_212
timestamp 1694700623
transform 1 0 25088 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_287
timestamp 1694700623
transform 1 0 33488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1694700623
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1694700623
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1694700623
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_78
timestamp 1694700623
transform 1 0 10080 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_125
timestamp 1694700623
transform 1 0 15344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1694700623
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1694700623
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1694700623
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1694700623
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1694700623
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_154
timestamp 1694700623
transform 1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_156
timestamp 1694700623
transform 1 0 18816 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_166
timestamp 1694700623
transform 1 0 19936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1694700623
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1694700623
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1694700623
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_286
timestamp 1694700623
transform 1 0 33376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_294
timestamp 1694700623
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_28
timestamp 1694700623
transform 1 0 4480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1694700623
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1694700623
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1694700623
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1694700623
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_82
timestamp 1694700623
transform 1 0 10528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_86
timestamp 1694700623
transform 1 0 10976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1694700623
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1694700623
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1694700623
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_128
timestamp 1694700623
transform 1 0 15680 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1694700623
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1694700623
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1694700623
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_36
timestamp 1694700623
transform 1 0 5376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_40
timestamp 1694700623
transform 1 0 5824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_44
timestamp 1694700623
transform 1 0 6272 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_60
timestamp 1694700623
transform 1 0 8064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_64
timestamp 1694700623
transform 1 0 8512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1694700623
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_88
timestamp 1694700623
transform 1 0 11200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_92
timestamp 1694700623
transform 1 0 11648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_94
timestamp 1694700623
transform 1 0 11872 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_105
timestamp 1694700623
transform 1 0 13104 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_150
timestamp 1694700623
transform 1 0 18144 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_168
timestamp 1694700623
transform 1 0 20160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_174
timestamp 1694700623
transform 1 0 20832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1694700623
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_228
timestamp 1694700623
transform 1 0 26880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_270
timestamp 1694700623
transform 1 0 31584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1694700623
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1694700623
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1694700623
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1694700623
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1694700623
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1694700623
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_4
timestamp 1694700623
transform 1 0 1792 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1694700623
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_33
timestamp 1694700623
transform 1 0 5040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_36
timestamp 1694700623
transform 1 0 5376 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_63
timestamp 1694700623
transform 1 0 8400 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_67
timestamp 1694700623
transform 1 0 8848 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_96
timestamp 1694700623
transform 1 0 12096 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_100
timestamp 1694700623
transform 1 0 12544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_130
timestamp 1694700623
transform 1 0 15904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1694700623
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_164
timestamp 1694700623
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_168
timestamp 1694700623
transform 1 0 20160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_198
timestamp 1694700623
transform 1 0 23520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_202
timestamp 1694700623
transform 1 0 23968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_266
timestamp 1694700623
transform 1 0 31136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_270
timestamp 1694700623
transform 1 0 31584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_274
timestamp 1694700623
transform 1 0 32032 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_290
timestamp 1694700623
transform 1 0 33824 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_294
timestamp 1694700623
transform 1 0 34272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1694700623
transform -1 0 34384 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1694700623
transform -1 0 34384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1694700623
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1694700623
transform -1 0 34384 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1694700623
transform 1 0 33040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 4480 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1694700623
transform -1 0 4816 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1694700623
transform -1 0 28784 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1694700623
transform 1 0 30576 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1694700623
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1694700623
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1694700623
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1694700623
transform 1 0 16800 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1694700623
transform 1 0 12992 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1694700623
transform 1 0 9184 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1694700623
transform 1 0 5488 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1694700623
transform -1 0 4816 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1694700623
transform -1 0 28784 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1694700623
transform -1 0 28784 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1694700623
transform -1 0 31136 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1694700623
transform 1 0 24416 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1694700623
transform -1 0 23520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1694700623
transform -1 0 19712 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1694700623
transform 1 0 12992 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1694700623
transform -1 0 12096 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1694700623
transform 1 0 5488 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1694700623
transform 1 0 31472 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1694700623
transform 1 0 29792 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1694700623
transform 1 0 29792 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1694700623
transform 1 0 31472 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1694700623
transform 1 0 29792 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1694700623
transform 1 0 29792 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1694700623
transform 1 0 25984 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output34
timestamp 1694700623
transform 1 0 26880 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35
timestamp 1694700623
transform 1 0 22960 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1694700623
transform 1 0 29792 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1694700623
transform 1 0 31472 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1694700623
transform -1 0 4480 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1694700623
transform -1 0 4480 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1694700623
transform -1 0 4480 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1694700623
transform -1 0 4480 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1694700623
transform -1 0 4480 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1694700623
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1694700623
transform 1 0 1568 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1694700623
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1694700623
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1694700623
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1694700623
transform 1 0 29792 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_25 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_26
timestamp 1694700623
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_27
timestamp 1694700623
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_28
timestamp 1694700623
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 34608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_29
timestamp 1694700623
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_30
timestamp 1694700623
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 34608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_31
timestamp 1694700623
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_32
timestamp 1694700623
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_33
timestamp 1694700623
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 34608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_34
timestamp 1694700623
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_35
timestamp 1694700623
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_36
timestamp 1694700623
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_37
timestamp 1694700623
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 34608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_38
timestamp 1694700623
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_39
timestamp 1694700623
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_40
timestamp 1694700623
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_41
timestamp 1694700623
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_42
timestamp 1694700623
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 34608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_43
timestamp 1694700623
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_44
timestamp 1694700623
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_45
timestamp 1694700623
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 34608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_46
timestamp 1694700623
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 34608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_47
timestamp 1694700623
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_48
timestamp 1694700623
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_49
timestamp 1694700623
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 34608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_50 pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_51
timestamp 1694700623
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_52
timestamp 1694700623
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_53
timestamp 1694700623
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_54
timestamp 1694700623
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_55
timestamp 1694700623
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_56
timestamp 1694700623
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_57
timestamp 1694700623
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_58
timestamp 1694700623
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_59
timestamp 1694700623
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_60
timestamp 1694700623
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_61
timestamp 1694700623
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_62
timestamp 1694700623
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_63
timestamp 1694700623
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_64
timestamp 1694700623
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_65
timestamp 1694700623
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1694700623
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_67
timestamp 1694700623
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_68
timestamp 1694700623
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_69
timestamp 1694700623
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1694700623
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1694700623
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1694700623
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1694700623
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1694700623
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1694700623
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1694700623
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1694700623
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_78
timestamp 1694700623
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_79
timestamp 1694700623
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_80
timestamp 1694700623
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1694700623
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_82
timestamp 1694700623
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_83
timestamp 1694700623
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_84
timestamp 1694700623
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1694700623
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_86
timestamp 1694700623
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_87
timestamp 1694700623
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_88
timestamp 1694700623
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_89
timestamp 1694700623
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_90
timestamp 1694700623
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_91
timestamp 1694700623
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_92
timestamp 1694700623
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_93
timestamp 1694700623
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_94
timestamp 1694700623
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_95
timestamp 1694700623
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_96
timestamp 1694700623
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_97
timestamp 1694700623
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_98
timestamp 1694700623
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_99
timestamp 1694700623
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_100
timestamp 1694700623
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_101
timestamp 1694700623
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_102
timestamp 1694700623
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_103
timestamp 1694700623
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_104
timestamp 1694700623
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_105
timestamp 1694700623
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_106
timestamp 1694700623
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_107
timestamp 1694700623
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_108
timestamp 1694700623
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_109
timestamp 1694700623
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_110
timestamp 1694700623
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_111
timestamp 1694700623
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_112
timestamp 1694700623
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_113
timestamp 1694700623
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_114
timestamp 1694700623
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_115
timestamp 1694700623
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_116
timestamp 1694700623
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_117
timestamp 1694700623
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_118
timestamp 1694700623
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_119
timestamp 1694700623
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_120
timestamp 1694700623
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_121
timestamp 1694700623
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_122
timestamp 1694700623
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_123
timestamp 1694700623
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_124
timestamp 1694700623
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_125
timestamp 1694700623
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_126
timestamp 1694700623
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_127
timestamp 1694700623
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_128
timestamp 1694700623
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_129
timestamp 1694700623
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_130
timestamp 1694700623
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_131
timestamp 1694700623
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_132
timestamp 1694700623
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_133
timestamp 1694700623
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_134
timestamp 1694700623
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_135
timestamp 1694700623
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_136
timestamp 1694700623
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_137
timestamp 1694700623
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_138
timestamp 1694700623
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_139
timestamp 1694700623
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_140
timestamp 1694700623
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_141
timestamp 1694700623
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_142
timestamp 1694700623
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_143
timestamp 1694700623
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_144
timestamp 1694700623
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_145
timestamp 1694700623
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_146
timestamp 1694700623
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_147
timestamp 1694700623
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_148
timestamp 1694700623
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_149
timestamp 1694700623
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_150
timestamp 1694700623
transform 1 0 5152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_151
timestamp 1694700623
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_152
timestamp 1694700623
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_153
timestamp 1694700623
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_154
timestamp 1694700623
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_155
timestamp 1694700623
transform 1 0 24192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_156
timestamp 1694700623
transform 1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_157
timestamp 1694700623
transform 1 0 31808 0 1 21952
box -86 -86 310 870
<< labels >>
flabel metal3 s 35200 5824 36000 5936 0 FreeSans 448 0 0 0 cal
port 0 nsew signal input
flabel metal3 s 35200 2688 36000 2800 0 FreeSans 448 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 11872 800 11984 0 FreeSans 448 0 0 0 clkc
port 2 nsew signal tristate
flabel metal3 s 0 13888 800 14000 0 FreeSans 448 0 0 0 comp
port 3 nsew signal input
flabel metal2 s 1792 0 1904 800 0 FreeSans 448 90 0 0 ctln[0]
port 4 nsew signal tristate
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 ctln[1]
port 5 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 ctln[2]
port 6 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 ctln[3]
port 7 nsew signal tristate
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 ctln[4]
port 8 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 ctln[5]
port 9 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 ctln[6]
port 10 nsew signal tristate
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 ctln[7]
port 11 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 ctln[8]
port 12 nsew signal tristate
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 ctln[9]
port 13 nsew signal tristate
flabel metal2 s 1792 25200 1904 26000 0 FreeSans 448 90 0 0 ctlp[0]
port 14 nsew signal tristate
flabel metal2 s 34048 25200 34160 26000 0 FreeSans 448 90 0 0 ctlp[1]
port 15 nsew signal tristate
flabel metal2 s 30464 25200 30576 26000 0 FreeSans 448 90 0 0 ctlp[2]
port 16 nsew signal tristate
flabel metal2 s 26880 25200 26992 26000 0 FreeSans 448 90 0 0 ctlp[3]
port 17 nsew signal tristate
flabel metal2 s 23296 25200 23408 26000 0 FreeSans 448 90 0 0 ctlp[4]
port 18 nsew signal tristate
flabel metal2 s 19712 25200 19824 26000 0 FreeSans 448 90 0 0 ctlp[5]
port 19 nsew signal tristate
flabel metal2 s 16128 25200 16240 26000 0 FreeSans 448 90 0 0 ctlp[6]
port 20 nsew signal tristate
flabel metal2 s 12544 25200 12656 26000 0 FreeSans 448 90 0 0 ctlp[7]
port 21 nsew signal tristate
flabel metal2 s 8960 25200 9072 26000 0 FreeSans 448 90 0 0 ctlp[8]
port 22 nsew signal tristate
flabel metal2 s 5376 25200 5488 26000 0 FreeSans 448 90 0 0 ctlp[9]
port 23 nsew signal tristate
flabel metal3 s 35200 4256 36000 4368 0 FreeSans 448 0 0 0 en
port 24 nsew signal input
flabel metal3 s 35200 10528 36000 10640 0 FreeSans 448 0 0 0 result[0]
port 25 nsew signal tristate
flabel metal3 s 35200 12096 36000 12208 0 FreeSans 448 0 0 0 result[1]
port 26 nsew signal tristate
flabel metal3 s 35200 13664 36000 13776 0 FreeSans 448 0 0 0 result[2]
port 27 nsew signal tristate
flabel metal3 s 35200 15232 36000 15344 0 FreeSans 448 0 0 0 result[3]
port 28 nsew signal tristate
flabel metal3 s 35200 16800 36000 16912 0 FreeSans 448 0 0 0 result[4]
port 29 nsew signal tristate
flabel metal3 s 35200 18368 36000 18480 0 FreeSans 448 0 0 0 result[5]
port 30 nsew signal tristate
flabel metal3 s 35200 19936 36000 20048 0 FreeSans 448 0 0 0 result[6]
port 31 nsew signal tristate
flabel metal3 s 35200 21504 36000 21616 0 FreeSans 448 0 0 0 result[7]
port 32 nsew signal tristate
flabel metal3 s 35200 23072 36000 23184 0 FreeSans 448 0 0 0 result[8]
port 33 nsew signal tristate
flabel metal3 s 35200 24640 36000 24752 0 FreeSans 448 0 0 0 result[9]
port 34 nsew signal tristate
flabel metal3 s 35200 1120 36000 1232 0 FreeSans 448 0 0 0 rstn
port 35 nsew signal input
flabel metal3 s 35200 8960 36000 9072 0 FreeSans 448 0 0 0 sample
port 36 nsew signal tristate
flabel metal3 s 0 5824 800 5936 0 FreeSans 448 0 0 0 trim[0]
port 37 nsew signal tristate
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 trim[1]
port 38 nsew signal tristate
flabel metal3 s 0 3808 800 3920 0 FreeSans 448 0 0 0 trim[2]
port 39 nsew signal tristate
flabel metal3 s 0 1792 800 1904 0 FreeSans 448 0 0 0 trim[3]
port 40 nsew signal tristate
flabel metal3 s 0 9856 800 9968 0 FreeSans 448 0 0 0 trim[4]
port 41 nsew signal tristate
flabel metal3 s 0 19936 800 20048 0 FreeSans 448 0 0 0 trimb[0]
port 42 nsew signal tristate
flabel metal3 s 0 17920 800 18032 0 FreeSans 448 0 0 0 trimb[1]
port 43 nsew signal tristate
flabel metal3 s 0 21952 800 22064 0 FreeSans 448 0 0 0 trimb[2]
port 44 nsew signal tristate
flabel metal3 s 0 23968 800 24080 0 FreeSans 448 0 0 0 trimb[3]
port 45 nsew signal tristate
flabel metal3 s 0 15904 800 16016 0 FreeSans 448 0 0 0 trimb[4]
port 46 nsew signal tristate
flabel metal3 s 35200 7392 36000 7504 0 FreeSans 448 0 0 0 valid
port 47 nsew signal tristate
flabel metal4 s 5342 3076 5662 22796 0 FreeSans 1280 90 0 0 vdd
port 48 nsew power bidirectional
flabel metal4 s 13658 3076 13978 22796 0 FreeSans 1280 90 0 0 vdd
port 48 nsew power bidirectional
flabel metal4 s 21974 3076 22294 22796 0 FreeSans 1280 90 0 0 vdd
port 48 nsew power bidirectional
flabel metal4 s 30290 3076 30610 22796 0 FreeSans 1280 90 0 0 vdd
port 48 nsew power bidirectional
flabel metal4 s 9500 3076 9820 22796 0 FreeSans 1280 90 0 0 vss
port 49 nsew ground bidirectional
flabel metal4 s 17816 3076 18136 22796 0 FreeSans 1280 90 0 0 vss
port 49 nsew ground bidirectional
flabel metal4 s 26132 3076 26452 22796 0 FreeSans 1280 90 0 0 vss
port 49 nsew ground bidirectional
flabel metal4 s 34448 3076 34768 22796 0 FreeSans 1280 90 0 0 vss
port 49 nsew ground bidirectional
rlabel metal1 17976 22736 17976 22736 0 vdd
rlabel via1 18056 21952 18056 21952 0 vss
rlabel metal2 26936 4256 26936 4256 0 _000_
rlabel metal3 30688 6664 30688 6664 0 _001_
rlabel metal2 22792 5768 22792 5768 0 _002_
rlabel metal2 22624 7672 22624 7672 0 _003_
rlabel metal2 31192 11480 31192 11480 0 _004_
rlabel metal2 29624 13328 29624 13328 0 _005_
rlabel metal2 33656 16184 33656 16184 0 _006_
rlabel metal2 33656 17920 33656 17920 0 _007_
rlabel metal2 27720 16912 27720 16912 0 _008_
rlabel metal2 33656 21056 33656 21056 0 _009_
rlabel metal2 31864 19992 31864 19992 0 _010_
rlabel metal2 30184 21224 30184 21224 0 _011_
rlabel metal2 6552 20440 6552 20440 0 _012_
rlabel metal2 6552 18536 6552 18536 0 _013_
rlabel metal2 28672 9240 28672 9240 0 _014_
rlabel metal2 28280 10864 28280 10864 0 _015_
rlabel metal2 16352 13048 16352 13048 0 _016_
rlabel metal2 14000 13720 14000 13720 0 _017_
rlabel metal2 24472 14448 24472 14448 0 _018_
rlabel metal2 23016 15568 23016 15568 0 _019_
rlabel metal2 15512 16352 15512 16352 0 _020_
rlabel metal2 20552 16968 20552 16968 0 _021_
rlabel metal2 16072 18928 16072 18928 0 _022_
rlabel metal2 20440 20356 20440 20356 0 _023_
rlabel metal2 21560 21672 21560 21672 0 _024_
rlabel metal2 14392 21280 14392 21280 0 _025_
rlabel metal2 12040 19712 12040 19712 0 _026_
rlabel metal2 10920 18144 10920 18144 0 _027_
rlabel metal3 11648 8344 11648 8344 0 _028_
rlabel metal2 8456 7000 8456 7000 0 _029_
rlabel metal2 8736 5096 8736 5096 0 _030_
rlabel metal2 16184 4592 16184 4592 0 _031_
rlabel metal2 16184 5544 16184 5544 0 _032_
rlabel metal3 4816 8344 4816 8344 0 _033_
rlabel metal2 2520 7168 2520 7168 0 _034_
rlabel metal2 2968 6328 2968 6328 0 _035_
rlabel metal2 5992 4984 5992 4984 0 _036_
rlabel metal3 20916 4312 20916 4312 0 _037_
rlabel metal2 8456 12824 8456 12824 0 _038_
rlabel metal2 2296 12264 2296 12264 0 _039_
rlabel metal2 13608 15568 13608 15568 0 _040_
rlabel metal3 5992 16856 5992 16856 0 _041_
rlabel metal2 6888 11536 6888 11536 0 _042_
rlabel metal3 3164 13944 3164 13944 0 _043_
rlabel metal2 30576 13160 30576 13160 0 _044_
rlabel metal2 30072 14784 30072 14784 0 _045_
rlabel metal2 28168 17248 28168 17248 0 _046_
rlabel metal2 25256 18368 25256 18368 0 _047_
rlabel metal2 24920 19488 24920 19488 0 _048_
rlabel metal2 19320 21000 19320 21000 0 _049_
rlabel metal3 15176 21784 15176 21784 0 _050_
rlabel metal2 10528 21784 10528 21784 0 _051_
rlabel metal3 7084 18424 7084 18424 0 _052_
rlabel metal2 25816 7896 25816 7896 0 _053_
rlabel metal2 2744 9688 2744 9688 0 _054_
rlabel metal2 23128 10528 23128 10528 0 _055_
rlabel metal3 24528 9688 24528 9688 0 _056_
rlabel metal2 20216 12656 20216 12656 0 _057_
rlabel metal3 18872 9744 18872 9744 0 _058_
rlabel metal3 17360 9688 17360 9688 0 _059_
rlabel metal3 25760 12152 25760 12152 0 _060_
rlabel metal2 23576 10976 23576 10976 0 _061_
rlabel metal2 23464 10304 23464 10304 0 _062_
rlabel metal2 6664 7840 6664 7840 0 _063_
rlabel metal2 2296 8008 2296 8008 0 _064_
rlabel metal3 8400 4200 8400 4200 0 _065_
rlabel metal2 19432 6608 19432 6608 0 _066_
rlabel metal2 3192 13048 3192 13048 0 _067_
rlabel metal2 25256 10136 25256 10136 0 _068_
rlabel metal3 23464 11480 23464 11480 0 _069_
rlabel metal2 21392 11144 21392 11144 0 _070_
rlabel metal2 18928 12712 18928 12712 0 _071_
rlabel metal2 25816 10584 25816 10584 0 _072_
rlabel metal2 28392 5768 28392 5768 0 _073_
rlabel metal2 24248 8736 24248 8736 0 _074_
rlabel metal3 25312 8232 25312 8232 0 _075_
rlabel metal2 26880 8680 26880 8680 0 _076_
rlabel metal2 27048 8372 27048 8372 0 _077_
rlabel metal2 26600 7784 26600 7784 0 _078_
rlabel metal2 22848 6664 22848 6664 0 _079_
rlabel metal2 27272 6944 27272 6944 0 _080_
rlabel metal3 27048 7448 27048 7448 0 _081_
rlabel metal3 29456 6552 29456 6552 0 _082_
rlabel metal3 27552 6776 27552 6776 0 _083_
rlabel metal2 29400 5936 29400 5936 0 _084_
rlabel metal2 21112 12488 21112 12488 0 _085_
rlabel metal2 21392 7672 21392 7672 0 _086_
rlabel metal3 21896 7448 21896 7448 0 _087_
rlabel metal3 24920 6552 24920 6552 0 _088_
rlabel metal2 23072 7448 23072 7448 0 _089_
rlabel metal2 26152 11816 26152 11816 0 _090_
rlabel metal2 25592 14280 25592 14280 0 _091_
rlabel metal2 26096 17640 26096 17640 0 _092_
rlabel metal2 25928 17360 25928 17360 0 _093_
rlabel metal2 29456 13944 29456 13944 0 _094_
rlabel metal2 3584 15400 3584 15400 0 _095_
rlabel metal2 20664 14056 20664 14056 0 _096_
rlabel metal2 20552 14952 20552 14952 0 _097_
rlabel metal2 24024 19376 24024 19376 0 _098_
rlabel metal2 29064 14112 29064 14112 0 _099_
rlabel metal2 29176 13216 29176 13216 0 _100_
rlabel metal2 29288 14056 29288 14056 0 _101_
rlabel metal2 29288 16408 29288 16408 0 _102_
rlabel metal2 29176 17136 29176 17136 0 _103_
rlabel metal3 30856 20776 30856 20776 0 _104_
rlabel metal2 26824 21112 26824 21112 0 _105_
rlabel metal2 26712 17528 26712 17528 0 _106_
rlabel metal2 26600 22008 26600 22008 0 _107_
rlabel metal3 28392 21448 28392 21448 0 _108_
rlabel metal2 29848 20888 29848 20888 0 _109_
rlabel metal2 10136 20356 10136 20356 0 _110_
rlabel metal2 9240 17976 9240 17976 0 _111_
rlabel metal2 29624 7728 29624 7728 0 _112_
rlabel metal2 22344 12096 22344 12096 0 _113_
rlabel metal3 21112 10304 21112 10304 0 _114_
rlabel metal2 11536 10808 11536 10808 0 _115_
rlabel metal2 21504 10696 21504 10696 0 _116_
rlabel metal2 22904 11088 22904 11088 0 _117_
rlabel metal2 16072 11368 16072 11368 0 _118_
rlabel metal2 20216 9296 20216 9296 0 _119_
rlabel metal2 17416 11144 17416 11144 0 _120_
rlabel metal2 19040 10584 19040 10584 0 _121_
rlabel metal3 26040 7952 26040 7952 0 _122_
rlabel metal3 28896 8344 28896 8344 0 _123_
rlabel metal2 15848 10864 15848 10864 0 _124_
rlabel metal2 14896 10808 14896 10808 0 _125_
rlabel metal2 21896 13496 21896 13496 0 _126_
rlabel metal2 16632 10864 16632 10864 0 _127_
rlabel metal2 27944 11032 27944 11032 0 _128_
rlabel metal2 16520 10920 16520 10920 0 _129_
rlabel metal2 16184 12600 16184 12600 0 _130_
rlabel metal2 7224 16464 7224 16464 0 _131_
rlabel metal2 14784 18648 14784 18648 0 _132_
rlabel metal3 16520 8904 16520 8904 0 _133_
rlabel metal2 14168 11032 14168 11032 0 _134_
rlabel metal2 14616 12600 14616 12600 0 _135_
rlabel metal3 22120 15848 22120 15848 0 _136_
rlabel metal2 22232 16184 22232 16184 0 _137_
rlabel metal2 22904 14560 22904 14560 0 _138_
rlabel metal2 22904 15792 22904 15792 0 _139_
rlabel metal2 20048 21560 20048 21560 0 _140_
rlabel metal2 19768 17136 19768 17136 0 _141_
rlabel metal2 16072 16800 16072 16800 0 _142_
rlabel metal3 19824 17640 19824 17640 0 _143_
rlabel metal2 15064 20356 15064 20356 0 _144_
rlabel metal2 16184 18704 16184 18704 0 _145_
rlabel metal3 19880 20664 19880 20664 0 _146_
rlabel metal3 20104 21448 20104 21448 0 _147_
rlabel metal3 14840 20664 14840 20664 0 _148_
rlabel metal2 12152 19600 12152 19600 0 _149_
rlabel metal3 11424 17640 11424 17640 0 _150_
rlabel metal3 13440 8008 13440 8008 0 _151_
rlabel metal2 15512 7000 15512 7000 0 _152_
rlabel metal2 15176 7504 15176 7504 0 _153_
rlabel metal3 14168 8232 14168 8232 0 _154_
rlabel metal2 13048 7952 13048 7952 0 _155_
rlabel metal2 12768 6104 12768 6104 0 _156_
rlabel metal3 13608 5880 13608 5880 0 _157_
rlabel metal2 14560 5656 14560 5656 0 _158_
rlabel metal2 15960 6160 15960 6160 0 _159_
rlabel metal2 15288 7112 15288 7112 0 _160_
rlabel metal2 22680 10360 22680 10360 0 _161_
rlabel metal2 20664 9296 20664 9296 0 _162_
rlabel metal2 21336 8456 21336 8456 0 _163_
rlabel metal2 10920 7112 10920 7112 0 _164_
rlabel metal2 6440 8456 6440 8456 0 _165_
rlabel metal2 6048 6888 6048 6888 0 _166_
rlabel metal2 6664 6328 6664 6328 0 _167_
rlabel metal3 10360 4536 10360 4536 0 _168_
rlabel metal2 19600 6888 19600 6888 0 _169_
rlabel metal2 18200 4816 18200 4816 0 _170_
rlabel metal3 11984 12152 11984 12152 0 _171_
rlabel metal2 12040 12656 12040 12656 0 _172_
rlabel metal2 5656 12656 5656 12656 0 _173_
rlabel metal2 8568 14168 8568 14168 0 _174_
rlabel metal2 10360 16072 10360 16072 0 _175_
rlabel metal3 9408 15960 9408 15960 0 _176_
rlabel metal2 11032 15400 11032 15400 0 _177_
rlabel metal2 6216 15540 6216 15540 0 _178_
rlabel metal2 7224 15680 7224 15680 0 _179_
rlabel metal2 7056 15400 7056 15400 0 _180_
rlabel metal3 6888 15288 6888 15288 0 _181_
rlabel metal2 6888 16128 6888 16128 0 _182_
rlabel metal2 7448 16520 7448 16520 0 _183_
rlabel metal2 5544 14392 5544 14392 0 _184_
rlabel metal2 4200 14896 4200 14896 0 _185_
rlabel metal2 5768 14056 5768 14056 0 _186_
rlabel metal2 6216 12152 6216 12152 0 _187_
rlabel metal2 7112 12208 7112 12208 0 _188_
rlabel metal2 34104 5096 34104 5096 0 cal
rlabel metal2 6104 13272 6104 13272 0 cal_count\[0\]
rlabel metal2 6552 15512 6552 15512 0 cal_count\[1\]
rlabel metal3 2800 15288 2800 15288 0 cal_count\[2\]
rlabel metal2 23128 12544 23128 12544 0 cal_count\[3\]
rlabel metal2 30072 5544 30072 5544 0 cal_itt\[0\]
rlabel metal2 31192 6216 31192 6216 0 cal_itt\[1\]
rlabel metal2 26936 6216 26936 6216 0 cal_itt\[2\]
rlabel metal3 24696 8344 24696 8344 0 cal_itt\[3\]
rlabel metal2 20552 9408 20552 9408 0 calibrate
rlabel metal3 33376 3416 33376 3416 0 clk
rlabel metal2 1960 11760 1960 11760 0 clkc
rlabel metal3 1302 13944 1302 13944 0 comp
rlabel metal2 2296 3500 2296 3500 0 ctln[0]
rlabel metal2 27608 4312 27608 4312 0 ctln[1]
rlabel metal2 31528 4872 31528 4872 0 ctln[2]
rlabel metal3 28168 3640 28168 3640 0 ctln[3]
rlabel metal2 23352 2198 23352 2198 0 ctln[4]
rlabel metal2 19768 2198 19768 2198 0 ctln[5]
rlabel metal2 16184 2086 16184 2086 0 ctln[6]
rlabel metal3 13384 3640 13384 3640 0 ctln[7]
rlabel metal3 9688 3640 9688 3640 0 ctln[8]
rlabel metal3 6048 3416 6048 3416 0 ctln[9]
rlabel metal2 2296 23408 2296 23408 0 ctlp[0]
rlabel metal3 30800 19432 30800 19432 0 ctlp[1]
rlabel metal3 29176 20888 29176 20888 0 ctlp[2]
rlabel metal3 27776 22568 27776 22568 0 ctlp[3]
rlabel metal2 23352 23898 23352 23898 0 ctlp[4]
rlabel metal2 19768 23898 19768 23898 0 ctlp[5]
rlabel metal3 16688 22568 16688 22568 0 ctlp[6]
rlabel metal2 12600 23898 12600 23898 0 ctlp[7]
rlabel metal2 9576 23912 9576 23912 0 ctlp[8]
rlabel metal2 5432 24346 5432 24346 0 ctlp[9]
rlabel metal2 34272 5096 34272 5096 0 en
rlabel metal2 11536 13160 11536 13160 0 en_co_clk
rlabel metal2 23464 14000 23464 14000 0 mask\[0\]
rlabel metal2 29512 14280 29512 14280 0 mask\[1\]
rlabel metal3 18816 15848 18816 15848 0 mask\[2\]
rlabel metal2 23688 17192 23688 17192 0 mask\[3\]
rlabel metal2 25816 17920 25816 17920 0 mask\[4\]
rlabel metal2 26096 20552 26096 20552 0 mask\[5\]
rlabel metal2 24696 20776 24696 20776 0 mask\[6\]
rlabel metal2 16968 21056 16968 21056 0 mask\[7\]
rlabel metal2 9968 20776 9968 20776 0 mask\[8\]
rlabel metal3 14112 18424 14112 18424 0 mask\[9\]
rlabel metal2 29064 7112 29064 7112 0 net1
rlabel metal2 26040 3808 26040 3808 0 net10
rlabel metal2 23576 3808 23576 3808 0 net11
rlabel metal3 20440 3528 20440 3528 0 net12
rlabel metal2 17416 3808 17416 3808 0 net13
rlabel metal2 12264 20748 12264 20748 0 net14
rlabel metal2 9352 3696 9352 3696 0 net15
rlabel metal2 6160 18200 6160 18200 0 net16
rlabel metal2 4144 22344 4144 22344 0 net17
rlabel metal2 33152 4424 33152 4424 0 net18
rlabel metal2 30912 4536 30912 4536 0 net19
rlabel metal2 31304 6888 31304 6888 0 net2
rlabel metal2 25928 4704 25928 4704 0 net20
rlabel metal2 23464 4480 23464 4480 0 net21
rlabel metal2 20328 5544 20328 5544 0 net22
rlabel metal3 18144 6104 18144 6104 0 net23
rlabel metal2 12600 22064 12600 22064 0 net24
rlabel metal2 11032 22064 11032 22064 0 net25
rlabel metal2 6216 18424 6216 18424 0 net26
rlabel metal2 31864 10360 31864 10360 0 net27
rlabel metal2 30072 13216 30072 13216 0 net28
rlabel via2 30184 15960 30184 15960 0 net29
rlabel metal3 2968 14504 2968 14504 0 net3
rlabel metal2 30632 17192 30632 17192 0 net30
rlabel metal3 25928 18424 25928 18424 0 net31
rlabel metal3 25872 20776 25872 20776 0 net32
rlabel metal2 25256 21112 25256 21112 0 net33
rlabel metal2 17752 21168 17752 21168 0 net34
rlabel metal3 23128 20832 23128 20832 0 net35
rlabel metal2 10920 18760 10920 18760 0 net36
rlabel metal2 31640 7952 31640 7952 0 net37
rlabel metal2 2968 11424 2968 11424 0 net38
rlabel metal2 2352 9688 2352 9688 0 net39
rlabel metal3 28728 5656 28728 5656 0 net4
rlabel metal2 4760 21168 4760 21168 0 net40
rlabel metal2 5432 21448 5432 21448 0 net41
rlabel metal2 3416 10304 3416 10304 0 net42
rlabel metal3 3304 20776 3304 20776 0 net43
rlabel metal2 2184 14224 2184 14224 0 net44
rlabel metal2 4480 21560 4480 21560 0 net45
rlabel metal3 4704 21336 4704 21336 0 net46
rlabel metal2 4536 16072 4536 16072 0 net47
rlabel metal2 29736 7448 29736 7448 0 net48
rlabel metal2 5208 6384 5208 6384 0 net49
rlabel metal2 33488 3416 33488 3416 0 net5
rlabel metal2 11480 9408 11480 9408 0 net50
rlabel metal2 9576 12208 9576 12208 0 net51
rlabel metal3 18312 4872 18312 4872 0 net52
rlabel metal2 16184 14504 16184 14504 0 net53
rlabel metal2 13496 19376 13496 19376 0 net54
rlabel metal3 2744 16912 2744 16912 0 net55
rlabel metal2 19432 15400 19432 15400 0 net56
rlabel metal2 20216 15568 20216 15568 0 net57
rlabel metal2 29456 4536 29456 4536 0 net58
rlabel metal2 26152 7224 26152 7224 0 net59
rlabel metal2 3304 12040 3304 12040 0 net6
rlabel metal3 32536 17416 32536 17416 0 net60
rlabel metal2 33880 19208 33880 19208 0 net61
rlabel metal3 29120 14392 29120 14392 0 net62
rlabel metal2 23856 21672 23856 21672 0 net63
rlabel metal2 28056 11592 28056 11592 0 net64
rlabel metal2 20440 5544 20440 5544 0 net65
rlabel metal2 2240 5880 2240 5880 0 net66
rlabel metal2 3080 11032 3080 11032 0 net67
rlabel metal3 7280 9800 7280 9800 0 net68
rlabel metal2 15176 5656 15176 5656 0 net69
rlabel metal2 4704 3528 4704 3528 0 net7
rlabel metal2 14056 15232 14056 15232 0 net70
rlabel metal2 10584 19208 10584 19208 0 net71
rlabel metal2 5544 16744 5544 16744 0 net72
rlabel metal2 16296 16408 16296 16408 0 net73
rlabel metal2 15512 5936 15512 5936 0 net74
rlabel metal2 28728 6944 28728 6944 0 net75
rlabel metal2 28504 7392 28504 7392 0 net76
rlabel metal3 33544 18984 33544 18984 0 net77
rlabel metal3 32032 19208 32032 19208 0 net78
rlabel metal2 29288 12824 29288 12824 0 net79
rlabel metal2 28504 4648 28504 4648 0 net8
rlabel metal2 23016 16016 23016 16016 0 net80
rlabel metal2 24192 15176 24192 15176 0 net81
rlabel metal2 31528 5824 31528 5824 0 net82
rlabel metal2 30520 4816 30520 4816 0 net9
rlabel metal2 33544 10304 33544 10304 0 result[0]
rlabel metal3 31892 12040 31892 12040 0 result[1]
rlabel metal3 31892 13608 31892 13608 0 result[2]
rlabel metal3 34426 15288 34426 15288 0 result[3]
rlabel metal3 33474 16856 33474 16856 0 result[4]
rlabel metal2 31864 18368 31864 18368 0 result[5]
rlabel metal2 28504 19936 28504 19936 0 result[6]
rlabel metal2 29400 18480 29400 18480 0 result[7]
rlabel metal2 25144 22008 25144 22008 0 result[8]
rlabel metal2 31080 18144 31080 18144 0 result[9]
rlabel metal3 32536 3528 32536 3528 0 rstn
rlabel metal2 33992 8736 33992 8736 0 sample
rlabel metal3 27160 11368 27160 11368 0 state\[0\]
rlabel metal3 23016 12936 23016 12936 0 state\[1\]
rlabel metal2 18648 13216 18648 13216 0 state\[2\]
rlabel metal3 1638 5880 1638 5880 0 trim[0]
rlabel metal3 1358 7896 1358 7896 0 trim[1]
rlabel metal3 1358 3864 1358 3864 0 trim[2]
rlabel metal3 2086 1848 2086 1848 0 trim[3]
rlabel metal3 1358 9912 1358 9912 0 trim[4]
rlabel metal2 12600 10248 12600 10248 0 trim_mask\[0\]
rlabel metal3 6608 7560 6608 7560 0 trim_mask\[1\]
rlabel metal2 11760 5320 11760 5320 0 trim_mask\[2\]
rlabel metal2 13160 4760 13160 4760 0 trim_mask\[3\]
rlabel metal2 16968 6328 16968 6328 0 trim_mask\[4\]
rlabel metal2 7224 9352 7224 9352 0 trim_val\[0\]
rlabel metal3 6440 7448 6440 7448 0 trim_val\[1\]
rlabel metal2 6104 5880 6104 5880 0 trim_val\[2\]
rlabel metal3 10136 4312 10136 4312 0 trim_val\[3\]
rlabel metal2 20216 6104 20216 6104 0 trim_val\[4\]
rlabel metal3 1358 19992 1358 19992 0 trimb[0]
rlabel metal3 1750 17976 1750 17976 0 trimb[1]
rlabel metal3 1358 22008 1358 22008 0 trimb[2]
rlabel metal3 1414 24024 1414 24024 0 trimb[3]
rlabel metal3 1358 15960 1358 15960 0 trimb[4]
rlabel metal2 31864 7392 31864 7392 0 valid
<< properties >>
string FIXED_BBOX 0 0 36000 26000
<< end >>
