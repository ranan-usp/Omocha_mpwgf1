* NGSPICE file created from buffer.ext - technology: gf180mcuD

.subckt XM2_buffer_inv2 G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 S D 0.090564f
C1 S G 0.138578f
C2 D G 0.001764f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.08816f
C5 S VSUBS 1.2321f
.ends

.subckt XM1_buffer_inv2 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt buffer_inv2 in vdd out vss
XXM2_buffer_inv2_0 in out vdd vss XM2_buffer_inv2
XXM1_buffer_inv2_0 in out vss XM1_buffer_inv2
C0 vdd out 0.086562f
C1 vdd in 0.034991f
C2 out in 0.057341f
C3 out vss 0.51823f
C4 in vss 0.460091f
C5 vdd vss 1.392287f
.ends

.subckt XM1_buffer_inv1 G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt buffer_inv1 in vdd out XM2_buffer_inv1_0/w_n90_n162# vss
XXM1_buffer_inv1_0 in out vss XM1_buffer_inv1
C0 XM2_buffer_inv1_0/w_n90_n162# out 0.007628f
C1 in vdd 0.040357f
C2 in out 0.058676f
C3 vdd out 0.142029f
C4 in XM2_buffer_inv1_0/w_n90_n162# 0.049713f
C5 vdd XM2_buffer_inv1_0/w_n90_n162# 0.009724f
C6 out vss 0.548612f
C7 in vss 0.543919f
C8 vdd vss 0.438255f
C9 XM2_buffer_inv1_0/w_n90_n162# vss 0.176185f
.ends

.subckt buffer middle out in vdd vss
Xbuffer_inv2_0 middle vdd out vss buffer_inv2
Xbuffer_inv1_0 in vdd middle buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vss buffer_inv1
C0 buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# in 0.051621f
C1 middle buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# 0.003733f
C2 vdd out 0.039935f
C3 vdd in 0.054064f
C4 middle vdd 0.190904f
C5 middle out 0.160929f
C6 middle in 0.119536f
C7 buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vdd 0.007171f
C8 middle vss 0.950535f
C9 in vss 0.600677f
C10 vdd vss 1.632177f
C11 buffer_inv1_0/XM2_buffer_inv1_0/w_n90_n162# vss 0.17473f
C12 out vss 0.56762f
.ends

