* NGSPICE file created from dac_in.ext - technology: gf180mcuD

.subckt dac_in inputp inputm vss vdd input_signal[0] input_signal[1] input_signal[2]
+ input_signal[3] input_signal[4] input_signal[5] input_signal[6] input_signal[7]
+ input_signal[8] input_signal[9]
Xphase_inverter_0 input_signal[0] input_signal[1] input_signal[2] input_signal[3]
+ input_signal[4] input_signal[5] input_signal[9] carray_in_1/n0 carray_in_1/n1 carray_in_1/n2
+ carray_in_1/n3 carray_in_1/n4 carray_in_1/n5 carray_in_1/n6 carray_in_1/n7 carray_in_1/n8
+ carray_in_1/n9 carray_in_0/n0 carray_in_0/n1 carray_in_0/n2 carray_in_0/n3 carray_in_0/n4
+ carray_in_0/n5 carray_in_0/n6 carray_in_0/n7 input_signal[7] input_signal[8] carray_in_0/n9
+ input_signal[6] carray_in_0/n8 vdd vss phase_inverter
C0 carray_in_1/n3 carray_in_1/n6 0.339322f
C1 vdd carray_in_0/n0 0.177806f
C2 carray_in_1/n9 carray_in_1/n4 3.741774f
C3 carray_in_1/n5 carray_in_1/n6 29.200403f
C4 vdd carray_in_1/n0 0.193605f
C5 inputp carray_in_0/n7 0.209952p
C6 carray_in_0/n1 carray_in_0/n8 0.333459f
C7 inputp carray_in_0/n3 13.12139f
C8 inputp carray_in_0/n9 0.846091p
C9 carray_in_0/n1 carray_in_1/n1 5.901133f
C10 carray_in_1/n4 carray_in_1/n6 0.617028f
C11 carray_in_1/n8 carray_in_1/n2 0.772498f
C12 carray_in_0/n4 carray_in_0/n7 1.70684f
C13 carray_in_0/n5 carray_in_0/n7 3.37237f
C14 carray_in_1/n8 carray_in_1/n7 50.742203f
C15 carray_in_0/n1 carray_in_0/n6 0.145088f
C16 carray_in_0/n5 carray_in_0/n3 0.350346f
C17 carray_in_0/n4 carray_in_0/n3 26.505903f
C18 carray_in_0/n4 carray_in_0/n9 3.741774f
C19 carray_in_0/n5 carray_in_0/n9 7.400846f
C20 vdd carray_in_0/n9 0.358842f
C21 carray_in_1/n8 carray_in_1/n1 0.333459f
C22 carray_in_0/n8 carray_in_0/n2 0.772498f
C23 carray_in_1/n3 carray_in_1/n2 23.465405f
C24 inputm carray_in_1/n8 0.420079p
C25 carray_in_1/n3 carray_in_1/n7 0.894213f
C26 carray_in_1/n5 carray_in_1/n2 0.210974f
C27 carray_in_0/n6 carray_in_0/n2 0.210444f
C28 carray_in_1/n0 carray_in_1/n1 8.401715f
C29 carray_in_1/n5 carray_in_1/n7 3.37237f
C30 carray_in_1/n9 carray_in_1/n6 14.718489f
C31 carray_in_1/n3 carray_in_1/n1 0.148119f
C32 carray_in_1/n5 carray_in_1/n1 0.145556f
C33 inputm carray_in_1/n0 1.640173f
C34 carray_in_1/n4 carray_in_1/n2 0.215946f
C35 carray_in_1/n9 vdd 0.348295f
C36 carray_in_1/n4 carray_in_1/n7 1.70684f
C37 carray_in_0/n8 carray_in_0/n7 50.742203f
C38 inputm carray_in_1/n3 13.12139f
C39 carray_in_0/n8 carray_in_0/n3 1.46349f
C40 carray_in_0/n8 carray_in_0/n9 87.65757f
C41 inputm carray_in_1/n5 52.485596f
C42 carray_in_1/n4 carray_in_1/n1 0.145617f
C43 carray_in_0/n6 carray_in_0/n7 34.900005f
C44 inputp carray_in_0/n5 52.485596f
C45 inputp carray_in_0/n4 26.242765f
C46 carray_in_0/n6 carray_in_0/n3 0.339322f
C47 carray_in_0/n6 carray_in_0/n9 14.718489f
C48 carray_in_0/n5 carray_in_0/n4 28.094206f
C49 carray_in_0/n1 carray_in_0/n2 15.574605f
C50 inputm carray_in_1/n4 26.242765f
C51 carray_in_0/n1 carray_in_0/n0 8.401715f
C52 carray_in_1/n9 carray_in_1/n2 0.997758f
C53 carray_in_1/n9 carray_in_1/n7 29.520088f
C54 carray_in_1/n9 carray_in_1/n1 0.39415f
C55 carray_in_1/n2 carray_in_1/n6 0.210444f
C56 carray_in_1/n7 carray_in_1/n6 34.900005f
C57 carray_in_0/n1 carray_in_0/n7 0.243006f
C58 carray_in_1/n3 carray_in_1/n8 1.46349f
C59 carray_in_1/n9 inputm 0.846091p
C60 carray_in_0/n1 carray_in_0/n3 0.148119f
C61 carray_in_0/n1 carray_in_0/n9 0.39415f
C62 carray_in_1/n5 carray_in_1/n8 5.6103f
C63 inputp carray_in_0/n8 0.420079p
C64 carray_in_1/n1 carray_in_1/n6 0.145088f
C65 carray_in_0/n8 carray_in_0/n4 2.84594f
C66 carray_in_0/n8 carray_in_0/n5 5.6103f
C67 inputp carray_in_0/n6 0.104976p
C68 carray_in_1/n4 carray_in_1/n8 2.84594f
C69 vdd carray_in_0/n8 0.117452f
C70 inputm carray_in_1/n6 0.104976p
C71 carray_in_0/n7 carray_in_0/n2 0.487626f
C72 carray_in_0/n5 carray_in_0/n6 29.200403f
C73 carray_in_0/n6 carray_in_0/n4 0.617028f
C74 carray_in_0/n3 carray_in_0/n2 23.465405f
C75 carray_in_0/n9 carray_in_0/n2 0.997758f
C76 carray_in_0/n0 carray_in_0/n9 0.82611f
C77 carray_in_1/n3 carray_in_1/n5 0.350346f
C78 carray_in_1/n2 carray_in_1/n7 0.487626f
C79 carray_in_1/n3 carray_in_1/n4 26.505903f
C80 carray_in_1/n4 carray_in_1/n5 28.094206f
C81 carray_in_1/n9 carray_in_1/n8 87.65758f
C82 carray_in_1/n2 carray_in_1/n1 15.574605f
C83 carray_in_0/n3 carray_in_0/n7 0.894213f
C84 carray_in_1/n1 carray_in_1/n7 0.243006f
C85 carray_in_0/n9 carray_in_0/n7 29.520088f
C86 carray_in_0/n1 inputp 3.280347f
C87 carray_in_0/n3 carray_in_0/n9 1.912414f
C88 inputm carray_in_1/n2 6.560692f
C89 carray_in_0/n1 carray_in_0/n5 0.145556f
C90 carray_in_0/n1 carray_in_0/n4 0.145617f
C91 inputm carray_in_1/n7 0.209952p
C92 carray_in_1/n9 carray_in_1/n0 0.82611f
C93 carray_in_0/n8 carray_in_0/n6 11.2197f
C94 carray_in_1/n8 carray_in_1/n6 11.2197f
C95 carray_in_1/n9 carray_in_1/n3 1.912414f
C96 inputm carray_in_1/n1 3.280347f
C97 inputp carray_in_0/n2 6.560692f
C98 inputp carray_in_0/n0 1.640173f
C99 carray_in_1/n9 carray_in_1/n5 7.400846f
C100 carray_in_0/n5 carray_in_0/n2 0.210974f
C101 carray_in_0/n4 carray_in_0/n2 0.215946f
C102 phase_inverter_0/_19_/Z vss 1.174253f
C103 phase_inverter_0/output30/a_224_472# vss 2.386102f
C104 phase_inverter_0/FILLER_0_1_60/a_484_472# vss 0.345058f $ **FLOATING
C105 phase_inverter_0/FILLER_0_1_60/a_36_472# vss 0.404746f
C106 phase_inverter_0/FILLER_0_1_60/a_572_375# vss 0.232991f
C107 phase_inverter_0/FILLER_0_1_60/a_124_375# vss 0.185089f $ **FLOATING
C108 phase_inverter_0/FILLER_0_0_28/a_36_472# vss 0.417394f
C109 phase_inverter_0/FILLER_0_0_28/a_124_375# vss 0.246306f $ **FLOATING
C110 phase_inverter_0/FILLER_0_13_72/a_3172_472# vss 0.345058f $ **FLOATING
C111 phase_inverter_0/FILLER_0_13_72/a_2724_472# vss 0.33241f $ **FLOATING
C112 phase_inverter_0/FILLER_0_13_72/a_2276_472# vss 0.33241f $ **FLOATING
C113 phase_inverter_0/FILLER_0_13_72/a_1828_472# vss 0.33241f $ **FLOATING
C114 phase_inverter_0/FILLER_0_13_72/a_1380_472# vss 0.33241f $ **FLOATING
C115 phase_inverter_0/FILLER_0_13_72/a_932_472# vss 0.33241f $ **FLOATING
C116 phase_inverter_0/FILLER_0_13_72/a_484_472# vss 0.33241f $ **FLOATING
C117 phase_inverter_0/FILLER_0_13_72/a_36_472# vss 0.404746f
C118 phase_inverter_0/FILLER_0_13_72/a_3260_375# vss 0.233093f $ **FLOATING
C119 phase_inverter_0/FILLER_0_13_72/a_2812_375# vss 0.17167f $ **FLOATING
C120 phase_inverter_0/FILLER_0_13_72/a_2364_375# vss 0.17167f $ **FLOATING
C121 phase_inverter_0/FILLER_0_13_72/a_1916_375# vss 0.17167f $ **FLOATING
C122 phase_inverter_0/FILLER_0_13_72/a_1468_375# vss 0.17167f $ **FLOATING
C123 phase_inverter_0/FILLER_0_13_72/a_1020_375# vss 0.17167f $ **FLOATING
C124 phase_inverter_0/FILLER_0_13_72/a_572_375# vss 0.17167f $ **FLOATING
C125 phase_inverter_0/FILLER_0_13_72/a_124_375# vss 0.185915f $ **FLOATING
C126 phase_inverter_0/FILLER_0_2_107/a_1380_472# vss 0.345058f $ **FLOATING
C127 phase_inverter_0/FILLER_0_2_107/a_932_472# vss 0.33241f $ **FLOATING
C128 phase_inverter_0/FILLER_0_2_107/a_484_472# vss 0.33241f $ **FLOATING
C129 phase_inverter_0/FILLER_0_2_107/a_36_472# vss 0.404746f
C130 phase_inverter_0/FILLER_0_2_107/a_1468_375# vss 0.233029f
C131 phase_inverter_0/FILLER_0_2_107/a_1020_375# vss 0.171606f $ **FLOATING
C132 phase_inverter_0/FILLER_0_2_107/a_572_375# vss 0.171606f $ **FLOATING
C133 phase_inverter_0/FILLER_0_2_107/a_124_375# vss 0.185399f $ **FLOATING
C134 phase_inverter_0/FILLER_0_5_104/a_484_472# vss 0.345058f $ **FLOATING
C135 phase_inverter_0/FILLER_0_5_104/a_36_472# vss 0.404746f
C136 phase_inverter_0/FILLER_0_5_104/a_572_375# vss 0.232991f
C137 phase_inverter_0/FILLER_0_5_104/a_124_375# vss 0.185089f $ **FLOATING
C138 phase_inverter_0/FILLER_0_6_37/a_6756_472# vss 0.345058f $ **FLOATING
C139 phase_inverter_0/FILLER_0_6_37/a_6308_472# vss 0.33241f $ **FLOATING
C140 phase_inverter_0/FILLER_0_6_37/a_5860_472# vss 0.33241f $ **FLOATING
C141 phase_inverter_0/FILLER_0_6_37/a_5412_472# vss 0.33241f $ **FLOATING
C142 phase_inverter_0/FILLER_0_6_37/a_4964_472# vss 0.33241f $ **FLOATING
C143 phase_inverter_0/FILLER_0_6_37/a_4516_472# vss 0.33241f $ **FLOATING
C144 phase_inverter_0/FILLER_0_6_37/a_4068_472# vss 0.33241f $ **FLOATING
C145 phase_inverter_0/FILLER_0_6_37/a_3620_472# vss 0.33241f $ **FLOATING
C146 phase_inverter_0/FILLER_0_6_37/a_3172_472# vss 0.33241f $ **FLOATING
C147 phase_inverter_0/FILLER_0_6_37/a_2724_472# vss 0.33241f $ **FLOATING
C148 phase_inverter_0/FILLER_0_6_37/a_2276_472# vss 0.33241f $ **FLOATING
C149 phase_inverter_0/FILLER_0_6_37/a_1828_472# vss 0.33241f $ **FLOATING
C150 phase_inverter_0/FILLER_0_6_37/a_1380_472# vss 0.33241f $ **FLOATING
C151 phase_inverter_0/FILLER_0_6_37/a_932_472# vss 0.33241f $ **FLOATING
C152 phase_inverter_0/FILLER_0_6_37/a_484_472# vss 0.33241f $ **FLOATING
C153 phase_inverter_0/FILLER_0_6_37/a_36_472# vss 0.404746f
C154 phase_inverter_0/FILLER_0_6_37/a_6844_375# vss 0.233068f $ **FLOATING
C155 phase_inverter_0/FILLER_0_6_37/a_6396_375# vss 0.171644f $ **FLOATING
C156 phase_inverter_0/FILLER_0_6_37/a_5948_375# vss 0.171644f $ **FLOATING
C157 phase_inverter_0/FILLER_0_6_37/a_5500_375# vss 0.171644f $ **FLOATING
C158 phase_inverter_0/FILLER_0_6_37/a_5052_375# vss 0.171644f $ **FLOATING
C159 phase_inverter_0/FILLER_0_6_37/a_4604_375# vss 0.171644f $ **FLOATING
C160 phase_inverter_0/FILLER_0_6_37/a_4156_375# vss 0.171644f $ **FLOATING
C161 phase_inverter_0/FILLER_0_6_37/a_3708_375# vss 0.171644f $ **FLOATING
C162 phase_inverter_0/FILLER_0_6_37/a_3260_375# vss 0.171644f $ **FLOATING
C163 phase_inverter_0/FILLER_0_6_37/a_2812_375# vss 0.171644f $ **FLOATING
C164 phase_inverter_0/FILLER_0_6_37/a_2364_375# vss 0.171644f $ **FLOATING
C165 phase_inverter_0/FILLER_0_6_37/a_1916_375# vss 0.171644f $ **FLOATING
C166 phase_inverter_0/FILLER_0_6_37/a_1468_375# vss 0.171644f $ **FLOATING
C167 phase_inverter_0/FILLER_0_6_37/a_1020_375# vss 0.171644f $ **FLOATING
C168 phase_inverter_0/FILLER_0_6_37/a_572_375# vss 0.171644f $ **FLOATING
C169 phase_inverter_0/FILLER_0_6_37/a_124_375# vss 0.185708f $ **FLOATING
C170 input_signal[4] vss 1.095436f
C171 phase_inverter_0/FILLER_0_8_101/a_36_472# vss 0.417394f
C172 phase_inverter_0/FILLER_0_8_101/a_124_375# vss 0.246306f $ **FLOATING
C173 phase_inverter_0/FILLER_0_16_104/a_36_472# vss 0.417394f
C174 phase_inverter_0/FILLER_0_16_104/a_124_375# vss 0.246306f $ **FLOATING
C175 phase_inverter_0/FILLER_0_12_28/a_36_472# vss 0.417394f
C176 phase_inverter_0/FILLER_0_12_28/a_124_375# vss 0.246306f $ **FLOATING
C177 phase_inverter_0/FILLER_0_11_2/a_6756_472# vss 0.345058f $ **FLOATING
C178 phase_inverter_0/FILLER_0_11_2/a_6308_472# vss 0.33241f $ **FLOATING
C179 phase_inverter_0/FILLER_0_11_2/a_5860_472# vss 0.33241f $ **FLOATING
C180 phase_inverter_0/FILLER_0_11_2/a_5412_472# vss 0.33241f $ **FLOATING
C181 phase_inverter_0/FILLER_0_11_2/a_4964_472# vss 0.33241f $ **FLOATING
C182 phase_inverter_0/FILLER_0_11_2/a_4516_472# vss 0.33241f $ **FLOATING
C183 phase_inverter_0/FILLER_0_11_2/a_4068_472# vss 0.33241f $ **FLOATING
C184 phase_inverter_0/FILLER_0_11_2/a_3620_472# vss 0.33241f $ **FLOATING
C185 phase_inverter_0/FILLER_0_11_2/a_3172_472# vss 0.33241f $ **FLOATING
C186 phase_inverter_0/FILLER_0_11_2/a_2724_472# vss 0.33241f $ **FLOATING
C187 phase_inverter_0/FILLER_0_11_2/a_2276_472# vss 0.33241f $ **FLOATING
C188 phase_inverter_0/FILLER_0_11_2/a_1828_472# vss 0.33241f $ **FLOATING
C189 phase_inverter_0/FILLER_0_11_2/a_1380_472# vss 0.33241f $ **FLOATING
C190 phase_inverter_0/FILLER_0_11_2/a_932_472# vss 0.33241f $ **FLOATING
C191 phase_inverter_0/FILLER_0_11_2/a_484_472# vss 0.33241f $ **FLOATING
C192 phase_inverter_0/FILLER_0_11_2/a_36_472# vss 0.404746f
C193 phase_inverter_0/FILLER_0_11_2/a_6844_375# vss 0.233068f $ **FLOATING
C194 phase_inverter_0/FILLER_0_11_2/a_6396_375# vss 0.171644f $ **FLOATING
C195 phase_inverter_0/FILLER_0_11_2/a_5948_375# vss 0.171644f $ **FLOATING
C196 phase_inverter_0/FILLER_0_11_2/a_5500_375# vss 0.171644f $ **FLOATING
C197 phase_inverter_0/FILLER_0_11_2/a_5052_375# vss 0.171644f $ **FLOATING
C198 phase_inverter_0/FILLER_0_11_2/a_4604_375# vss 0.171644f $ **FLOATING
C199 phase_inverter_0/FILLER_0_11_2/a_4156_375# vss 0.171644f $ **FLOATING
C200 phase_inverter_0/FILLER_0_11_2/a_3708_375# vss 0.171644f $ **FLOATING
C201 phase_inverter_0/FILLER_0_11_2/a_3260_375# vss 0.171644f $ **FLOATING
C202 phase_inverter_0/FILLER_0_11_2/a_2812_375# vss 0.171644f $ **FLOATING
C203 phase_inverter_0/FILLER_0_11_2/a_2364_375# vss 0.171644f $ **FLOATING
C204 phase_inverter_0/FILLER_0_11_2/a_1916_375# vss 0.171644f $ **FLOATING
C205 phase_inverter_0/FILLER_0_11_2/a_1468_375# vss 0.171644f $ **FLOATING
C206 phase_inverter_0/FILLER_0_11_2/a_1020_375# vss 0.171644f $ **FLOATING
C207 phase_inverter_0/FILLER_0_11_2/a_572_375# vss 0.171644f $ **FLOATING
C208 phase_inverter_0/FILLER_0_11_2/a_124_375# vss 0.185708f $ **FLOATING
C209 phase_inverter_0/FILLER_0_16_70/a_36_472# vss 0.417394f
C210 phase_inverter_0/FILLER_0_16_70/a_124_375# vss 0.246306f $ **FLOATING
C211 phase_inverter_0/FILLER_0_15_8/a_3172_472# vss 0.345058f $ **FLOATING
C212 phase_inverter_0/FILLER_0_15_8/a_2724_472# vss 0.33241f $ **FLOATING
C213 phase_inverter_0/FILLER_0_15_8/a_2276_472# vss 0.33241f $ **FLOATING
C214 phase_inverter_0/FILLER_0_15_8/a_1828_472# vss 0.33241f $ **FLOATING
C215 phase_inverter_0/FILLER_0_15_8/a_1380_472# vss 0.33241f $ **FLOATING
C216 phase_inverter_0/FILLER_0_15_8/a_932_472# vss 0.33241f $ **FLOATING
C217 phase_inverter_0/FILLER_0_15_8/a_484_472# vss 0.33241f $ **FLOATING
C218 phase_inverter_0/FILLER_0_15_8/a_36_472# vss 0.404746f
C219 phase_inverter_0/FILLER_0_15_8/a_3260_375# vss 0.233093f $ **FLOATING
C220 phase_inverter_0/FILLER_0_15_8/a_2812_375# vss 0.17167f $ **FLOATING
C221 phase_inverter_0/FILLER_0_15_8/a_2364_375# vss 0.17167f $ **FLOATING
C222 phase_inverter_0/FILLER_0_15_8/a_1916_375# vss 0.17167f $ **FLOATING
C223 phase_inverter_0/FILLER_0_15_8/a_1468_375# vss 0.17167f $ **FLOATING
C224 phase_inverter_0/FILLER_0_15_8/a_1020_375# vss 0.17167f $ **FLOATING
C225 phase_inverter_0/FILLER_0_15_8/a_572_375# vss 0.17167f $ **FLOATING
C226 phase_inverter_0/FILLER_0_15_8/a_124_375# vss 0.185915f $ **FLOATING
C227 vdd vss 0.426348p
C228 phase_inverter_0/FILLER_0_0_36/a_3172_472# vss 0.345058f $ **FLOATING
C229 phase_inverter_0/FILLER_0_0_36/a_2724_472# vss 0.33241f $ **FLOATING
C230 phase_inverter_0/FILLER_0_0_36/a_2276_472# vss 0.33241f $ **FLOATING
C231 phase_inverter_0/FILLER_0_0_36/a_1828_472# vss 0.33241f $ **FLOATING
C232 phase_inverter_0/FILLER_0_0_36/a_1380_472# vss 0.33241f $ **FLOATING
C233 phase_inverter_0/FILLER_0_0_36/a_932_472# vss 0.33241f $ **FLOATING
C234 phase_inverter_0/FILLER_0_0_36/a_484_472# vss 0.33241f $ **FLOATING
C235 phase_inverter_0/FILLER_0_0_36/a_36_472# vss 0.409475f
C236 phase_inverter_0/FILLER_0_0_36/a_3260_375# vss 0.233093f $ **FLOATING
C237 phase_inverter_0/FILLER_0_0_36/a_2812_375# vss 0.17167f $ **FLOATING
C238 phase_inverter_0/FILLER_0_0_36/a_2364_375# vss 0.17167f $ **FLOATING
C239 phase_inverter_0/FILLER_0_0_36/a_1916_375# vss 0.17167f $ **FLOATING
C240 phase_inverter_0/FILLER_0_0_36/a_1468_375# vss 0.17167f $ **FLOATING
C241 phase_inverter_0/FILLER_0_0_36/a_1020_375# vss 0.17167f $ **FLOATING
C242 phase_inverter_0/FILLER_0_0_36/a_572_375# vss 0.17167f $ **FLOATING
C243 phase_inverter_0/FILLER_0_0_36/a_124_375# vss 0.185915f $ **FLOATING
C244 phase_inverter_0/_10_/Z vss 1.18279f
C245 phase_inverter_0/_10_/a_36_160# vss 0.386641f $ **FLOATING
C246 phase_inverter_0/FILLER_0_10_107/a_1380_472# vss 0.345058f $ **FLOATING
C247 phase_inverter_0/FILLER_0_10_107/a_932_472# vss 0.33241f $ **FLOATING
C248 phase_inverter_0/FILLER_0_10_107/a_484_472# vss 0.33241f $ **FLOATING
C249 phase_inverter_0/FILLER_0_10_107/a_36_472# vss 0.404746f
C250 phase_inverter_0/FILLER_0_10_107/a_1468_375# vss 0.233029f
C251 phase_inverter_0/FILLER_0_10_107/a_1020_375# vss 0.171606f $ **FLOATING
C252 phase_inverter_0/FILLER_0_10_107/a_572_375# vss 0.171606f $ **FLOATING
C253 phase_inverter_0/FILLER_0_10_107/a_124_375# vss 0.185399f $ **FLOATING
C254 phase_inverter_0/FILLER_0_12_37/a_6756_472# vss 0.345058f $ **FLOATING
C255 phase_inverter_0/FILLER_0_12_37/a_6308_472# vss 0.33241f $ **FLOATING
C256 phase_inverter_0/FILLER_0_12_37/a_5860_472# vss 0.33241f $ **FLOATING
C257 phase_inverter_0/FILLER_0_12_37/a_5412_472# vss 0.33241f $ **FLOATING
C258 phase_inverter_0/FILLER_0_12_37/a_4964_472# vss 0.33241f $ **FLOATING
C259 phase_inverter_0/FILLER_0_12_37/a_4516_472# vss 0.33241f $ **FLOATING
C260 phase_inverter_0/FILLER_0_12_37/a_4068_472# vss 0.33241f $ **FLOATING
C261 phase_inverter_0/FILLER_0_12_37/a_3620_472# vss 0.33241f $ **FLOATING
C262 phase_inverter_0/FILLER_0_12_37/a_3172_472# vss 0.33241f $ **FLOATING
C263 phase_inverter_0/FILLER_0_12_37/a_2724_472# vss 0.33241f $ **FLOATING
C264 phase_inverter_0/FILLER_0_12_37/a_2276_472# vss 0.33241f $ **FLOATING
C265 phase_inverter_0/FILLER_0_12_37/a_1828_472# vss 0.33241f $ **FLOATING
C266 phase_inverter_0/FILLER_0_12_37/a_1380_472# vss 0.33241f $ **FLOATING
C267 phase_inverter_0/FILLER_0_12_37/a_932_472# vss 0.33241f $ **FLOATING
C268 phase_inverter_0/FILLER_0_12_37/a_484_472# vss 0.33241f $ **FLOATING
C269 phase_inverter_0/FILLER_0_12_37/a_36_472# vss 0.404746f
C270 phase_inverter_0/FILLER_0_12_37/a_6844_375# vss 0.233068f $ **FLOATING
C271 phase_inverter_0/FILLER_0_12_37/a_6396_375# vss 0.171644f $ **FLOATING
C272 phase_inverter_0/FILLER_0_12_37/a_5948_375# vss 0.171644f $ **FLOATING
C273 phase_inverter_0/FILLER_0_12_37/a_5500_375# vss 0.171644f $ **FLOATING
C274 phase_inverter_0/FILLER_0_12_37/a_5052_375# vss 0.171644f $ **FLOATING
C275 phase_inverter_0/FILLER_0_12_37/a_4604_375# vss 0.171644f $ **FLOATING
C276 phase_inverter_0/FILLER_0_12_37/a_4156_375# vss 0.171644f $ **FLOATING
C277 phase_inverter_0/FILLER_0_12_37/a_3708_375# vss 0.171644f $ **FLOATING
C278 phase_inverter_0/FILLER_0_12_37/a_3260_375# vss 0.171644f $ **FLOATING
C279 phase_inverter_0/FILLER_0_12_37/a_2812_375# vss 0.171644f $ **FLOATING
C280 phase_inverter_0/FILLER_0_12_37/a_2364_375# vss 0.171644f $ **FLOATING
C281 phase_inverter_0/FILLER_0_12_37/a_1916_375# vss 0.171644f $ **FLOATING
C282 phase_inverter_0/FILLER_0_12_37/a_1468_375# vss 0.171644f $ **FLOATING
C283 phase_inverter_0/FILLER_0_12_37/a_1020_375# vss 0.171644f $ **FLOATING
C284 phase_inverter_0/FILLER_0_12_37/a_572_375# vss 0.171644f $ **FLOATING
C285 phase_inverter_0/FILLER_0_12_37/a_124_375# vss 0.185708f $ **FLOATING
C286 phase_inverter_0/FILLER_0_13_104/a_484_472# vss 0.345058f $ **FLOATING
C287 phase_inverter_0/FILLER_0_13_104/a_36_472# vss 0.404746f
C288 phase_inverter_0/FILLER_0_13_104/a_572_375# vss 0.232991f
C289 phase_inverter_0/FILLER_0_13_104/a_124_375# vss 0.185089f $ **FLOATING
C290 input_signal[6] vss 1.014523f
C291 phase_inverter_0/_11_/Z vss 1.137333f
C292 phase_inverter_0/_11_/a_36_113# vss 0.418095f
C293 phase_inverter_0/FILLER_0_9_66/a_36_472# vss 0.417394f
C294 phase_inverter_0/FILLER_0_9_66/a_124_375# vss 0.246306f $ **FLOATING
C295 phase_inverter_0/FILLER_0_3_12/a_3172_472# vss 0.345058f $ **FLOATING
C296 phase_inverter_0/FILLER_0_3_12/a_2724_472# vss 0.33241f $ **FLOATING
C297 phase_inverter_0/FILLER_0_3_12/a_2276_472# vss 0.33241f $ **FLOATING
C298 phase_inverter_0/FILLER_0_3_12/a_1828_472# vss 0.33241f $ **FLOATING
C299 phase_inverter_0/FILLER_0_3_12/a_1380_472# vss 0.33241f $ **FLOATING
C300 phase_inverter_0/FILLER_0_3_12/a_932_472# vss 0.33241f $ **FLOATING
C301 phase_inverter_0/FILLER_0_3_12/a_484_472# vss 0.33241f $ **FLOATING
C302 phase_inverter_0/FILLER_0_3_12/a_36_472# vss 0.404746f
C303 phase_inverter_0/FILLER_0_3_12/a_3260_375# vss 0.233093f $ **FLOATING
C304 phase_inverter_0/FILLER_0_3_12/a_2812_375# vss 0.17167f $ **FLOATING
C305 phase_inverter_0/FILLER_0_3_12/a_2364_375# vss 0.17167f $ **FLOATING
C306 phase_inverter_0/FILLER_0_3_12/a_1916_375# vss 0.17167f $ **FLOATING
C307 phase_inverter_0/FILLER_0_3_12/a_1468_375# vss 0.17167f $ **FLOATING
C308 phase_inverter_0/FILLER_0_3_12/a_1020_375# vss 0.17167f $ **FLOATING
C309 phase_inverter_0/FILLER_0_3_12/a_572_375# vss 0.17167f $ **FLOATING
C310 phase_inverter_0/FILLER_0_3_12/a_124_375# vss 0.185915f $ **FLOATING
C311 phase_inverter_0/FILLER_0_2_2/a_3172_472# vss 0.345058f $ **FLOATING
C312 phase_inverter_0/FILLER_0_2_2/a_2724_472# vss 0.33241f $ **FLOATING
C313 phase_inverter_0/FILLER_0_2_2/a_2276_472# vss 0.33241f $ **FLOATING
C314 phase_inverter_0/FILLER_0_2_2/a_1828_472# vss 0.33241f $ **FLOATING
C315 phase_inverter_0/FILLER_0_2_2/a_1380_472# vss 0.33241f $ **FLOATING
C316 phase_inverter_0/FILLER_0_2_2/a_932_472# vss 0.33241f $ **FLOATING
C317 phase_inverter_0/FILLER_0_2_2/a_484_472# vss 0.33241f $ **FLOATING
C318 phase_inverter_0/FILLER_0_2_2/a_36_472# vss 0.404746f
C319 phase_inverter_0/FILLER_0_2_2/a_3260_375# vss 0.233093f $ **FLOATING
C320 phase_inverter_0/FILLER_0_2_2/a_2812_375# vss 0.17167f $ **FLOATING
C321 phase_inverter_0/FILLER_0_2_2/a_2364_375# vss 0.17167f $ **FLOATING
C322 phase_inverter_0/FILLER_0_2_2/a_1916_375# vss 0.17167f $ **FLOATING
C323 phase_inverter_0/FILLER_0_2_2/a_1468_375# vss 0.17167f $ **FLOATING
C324 phase_inverter_0/FILLER_0_2_2/a_1020_375# vss 0.17167f $ **FLOATING
C325 phase_inverter_0/FILLER_0_2_2/a_572_375# vss 0.17167f $ **FLOATING
C326 phase_inverter_0/FILLER_0_2_2/a_124_375# vss 0.185915f $ **FLOATING
C327 phase_inverter_0/FILLER_0_13_2/a_6756_472# vss 0.345058f $ **FLOATING
C328 phase_inverter_0/FILLER_0_13_2/a_6308_472# vss 0.33241f $ **FLOATING
C329 phase_inverter_0/FILLER_0_13_2/a_5860_472# vss 0.33241f $ **FLOATING
C330 phase_inverter_0/FILLER_0_13_2/a_5412_472# vss 0.33241f $ **FLOATING
C331 phase_inverter_0/FILLER_0_13_2/a_4964_472# vss 0.33241f $ **FLOATING
C332 phase_inverter_0/FILLER_0_13_2/a_4516_472# vss 0.33241f $ **FLOATING
C333 phase_inverter_0/FILLER_0_13_2/a_4068_472# vss 0.33241f $ **FLOATING
C334 phase_inverter_0/FILLER_0_13_2/a_3620_472# vss 0.33241f $ **FLOATING
C335 phase_inverter_0/FILLER_0_13_2/a_3172_472# vss 0.33241f $ **FLOATING
C336 phase_inverter_0/FILLER_0_13_2/a_2724_472# vss 0.33241f $ **FLOATING
C337 phase_inverter_0/FILLER_0_13_2/a_2276_472# vss 0.33241f $ **FLOATING
C338 phase_inverter_0/FILLER_0_13_2/a_1828_472# vss 0.33241f $ **FLOATING
C339 phase_inverter_0/FILLER_0_13_2/a_1380_472# vss 0.33241f $ **FLOATING
C340 phase_inverter_0/FILLER_0_13_2/a_932_472# vss 0.33241f $ **FLOATING
C341 phase_inverter_0/FILLER_0_13_2/a_484_472# vss 0.33241f $ **FLOATING
C342 phase_inverter_0/FILLER_0_13_2/a_36_472# vss 0.404746f
C343 phase_inverter_0/FILLER_0_13_2/a_6844_375# vss 0.233068f $ **FLOATING
C344 phase_inverter_0/FILLER_0_13_2/a_6396_375# vss 0.171644f $ **FLOATING
C345 phase_inverter_0/FILLER_0_13_2/a_5948_375# vss 0.171644f $ **FLOATING
C346 phase_inverter_0/FILLER_0_13_2/a_5500_375# vss 0.171644f $ **FLOATING
C347 phase_inverter_0/FILLER_0_13_2/a_5052_375# vss 0.171644f $ **FLOATING
C348 phase_inverter_0/FILLER_0_13_2/a_4604_375# vss 0.171644f $ **FLOATING
C349 phase_inverter_0/FILLER_0_13_2/a_4156_375# vss 0.171644f $ **FLOATING
C350 phase_inverter_0/FILLER_0_13_2/a_3708_375# vss 0.171644f $ **FLOATING
C351 phase_inverter_0/FILLER_0_13_2/a_3260_375# vss 0.171644f $ **FLOATING
C352 phase_inverter_0/FILLER_0_13_2/a_2812_375# vss 0.171644f $ **FLOATING
C353 phase_inverter_0/FILLER_0_13_2/a_2364_375# vss 0.171644f $ **FLOATING
C354 phase_inverter_0/FILLER_0_13_2/a_1916_375# vss 0.171644f $ **FLOATING
C355 phase_inverter_0/FILLER_0_13_2/a_1468_375# vss 0.171644f $ **FLOATING
C356 phase_inverter_0/FILLER_0_13_2/a_1020_375# vss 0.171644f $ **FLOATING
C357 phase_inverter_0/FILLER_0_13_2/a_572_375# vss 0.171644f $ **FLOATING
C358 phase_inverter_0/FILLER_0_13_2/a_124_375# vss 0.185708f $ **FLOATING
C359 phase_inverter_0/FILLER_0_0_12/a_1380_472# vss 0.345058f $ **FLOATING
C360 phase_inverter_0/FILLER_0_0_12/a_932_472# vss 0.33241f $ **FLOATING
C361 phase_inverter_0/FILLER_0_0_12/a_484_472# vss 0.33241f $ **FLOATING
C362 phase_inverter_0/FILLER_0_0_12/a_36_472# vss 0.404746f
C363 phase_inverter_0/FILLER_0_0_12/a_1468_375# vss 0.233029f
C364 phase_inverter_0/FILLER_0_0_12/a_1020_375# vss 0.171606f $ **FLOATING
C365 phase_inverter_0/FILLER_0_0_12/a_572_375# vss 0.171606f $ **FLOATING
C366 phase_inverter_0/FILLER_0_0_12/a_124_375# vss 0.185399f $ **FLOATING
C367 phase_inverter_0/FILLER_0_3_44/a_1380_472# vss 0.345058f $ **FLOATING
C368 phase_inverter_0/FILLER_0_3_44/a_932_472# vss 0.33241f $ **FLOATING
C369 phase_inverter_0/FILLER_0_3_44/a_484_472# vss 0.33241f $ **FLOATING
C370 phase_inverter_0/FILLER_0_3_44/a_36_472# vss 0.404746f
C371 phase_inverter_0/FILLER_0_3_44/a_1468_375# vss 0.233029f
C372 phase_inverter_0/FILLER_0_3_44/a_1020_375# vss 0.171606f $ **FLOATING
C373 phase_inverter_0/FILLER_0_3_44/a_572_375# vss 0.171606f $ **FLOATING
C374 phase_inverter_0/FILLER_0_3_44/a_124_375# vss 0.185399f $ **FLOATING
C375 phase_inverter_0/_12_/Z vss 1.135084f
C376 phase_inverter_0/_12_/a_36_113# vss 0.418095f
C377 phase_inverter_0/FILLER_0_15_56/a_484_472# vss 0.345058f $ **FLOATING
C378 phase_inverter_0/FILLER_0_15_56/a_36_472# vss 0.404746f
C379 phase_inverter_0/FILLER_0_15_56/a_572_375# vss 0.232991f
C380 phase_inverter_0/FILLER_0_15_56/a_124_375# vss 0.185089f $ **FLOATING
C381 phase_inverter_0/_13_/Z vss 1.131177f
C382 phase_inverter_0/_13_/a_36_113# vss 0.418095f
C383 phase_inverter_0/FILLER_0_2_101/a_36_472# vss 0.417394f
C384 phase_inverter_0/FILLER_0_2_101/a_124_375# vss 0.246306f $ **FLOATING
C385 phase_inverter_0/FILLER_0_12_12/a_1380_472# vss 0.345058f $ **FLOATING
C386 phase_inverter_0/FILLER_0_12_12/a_932_472# vss 0.33241f $ **FLOATING
C387 phase_inverter_0/FILLER_0_12_12/a_484_472# vss 0.33241f $ **FLOATING
C388 phase_inverter_0/FILLER_0_12_12/a_36_472# vss 0.404746f
C389 phase_inverter_0/FILLER_0_12_12/a_1468_375# vss 0.233029f
C390 phase_inverter_0/FILLER_0_12_12/a_1020_375# vss 0.171606f $ **FLOATING
C391 phase_inverter_0/FILLER_0_12_12/a_572_375# vss 0.171606f $ **FLOATING
C392 phase_inverter_0/FILLER_0_12_12/a_124_375# vss 0.185399f $ **FLOATING
C393 input_signal[8] vss 1.074195f
C394 phase_inverter_0/_14_/Z vss 1.171827f
C395 phase_inverter_0/_14_/a_36_113# vss 0.418095f
C396 phase_inverter_0/FILLER_0_4_2/a_3172_472# vss 0.345058f $ **FLOATING
C397 phase_inverter_0/FILLER_0_4_2/a_2724_472# vss 0.33241f $ **FLOATING
C398 phase_inverter_0/FILLER_0_4_2/a_2276_472# vss 0.33241f $ **FLOATING
C399 phase_inverter_0/FILLER_0_4_2/a_1828_472# vss 0.33241f $ **FLOATING
C400 phase_inverter_0/FILLER_0_4_2/a_1380_472# vss 0.33241f $ **FLOATING
C401 phase_inverter_0/FILLER_0_4_2/a_932_472# vss 0.33241f $ **FLOATING
C402 phase_inverter_0/FILLER_0_4_2/a_484_472# vss 0.33241f $ **FLOATING
C403 phase_inverter_0/FILLER_0_4_2/a_36_472# vss 0.404746f
C404 phase_inverter_0/FILLER_0_4_2/a_3260_375# vss 0.233093f $ **FLOATING
C405 phase_inverter_0/FILLER_0_4_2/a_2812_375# vss 0.17167f $ **FLOATING
C406 phase_inverter_0/FILLER_0_4_2/a_2364_375# vss 0.17167f $ **FLOATING
C407 phase_inverter_0/FILLER_0_4_2/a_1916_375# vss 0.17167f $ **FLOATING
C408 phase_inverter_0/FILLER_0_4_2/a_1468_375# vss 0.17167f $ **FLOATING
C409 phase_inverter_0/FILLER_0_4_2/a_1020_375# vss 0.17167f $ **FLOATING
C410 phase_inverter_0/FILLER_0_4_2/a_572_375# vss 0.17167f $ **FLOATING
C411 phase_inverter_0/FILLER_0_4_2/a_124_375# vss 0.185915f $ **FLOATING
C412 phase_inverter_0/FILLER_0_15_2/a_36_472# vss 0.417394f
C413 phase_inverter_0/FILLER_0_15_2/a_124_375# vss 0.246306f $ **FLOATING
C414 phase_inverter_0/_15_/Z vss 1.167741f
C415 phase_inverter_0/_15_/a_36_113# vss 0.418095f
C416 phase_inverter_0/FILLER_0_6_107/a_36_472# vss 0.417394f
C417 phase_inverter_0/FILLER_0_6_107/a_124_375# vss 0.246306f $ **FLOATING
C418 phase_inverter_0/FILLER_0_9_104/a_484_472# vss 0.345058f $ **FLOATING
C419 phase_inverter_0/FILLER_0_9_104/a_36_472# vss 0.404746f
C420 phase_inverter_0/FILLER_0_9_104/a_572_375# vss 0.232991f
C421 phase_inverter_0/FILLER_0_9_104/a_124_375# vss 0.185089f $ **FLOATING
C422 phase_inverter_0/FILLER_0_9_72/a_3172_472# vss 0.345058f $ **FLOATING
C423 phase_inverter_0/FILLER_0_9_72/a_2724_472# vss 0.33241f $ **FLOATING
C424 phase_inverter_0/FILLER_0_9_72/a_2276_472# vss 0.33241f $ **FLOATING
C425 phase_inverter_0/FILLER_0_9_72/a_1828_472# vss 0.33241f $ **FLOATING
C426 phase_inverter_0/FILLER_0_9_72/a_1380_472# vss 0.33241f $ **FLOATING
C427 phase_inverter_0/FILLER_0_9_72/a_932_472# vss 0.33241f $ **FLOATING
C428 phase_inverter_0/FILLER_0_9_72/a_484_472# vss 0.33241f $ **FLOATING
C429 phase_inverter_0/FILLER_0_9_72/a_36_472# vss 0.404746f
C430 phase_inverter_0/FILLER_0_9_72/a_3260_375# vss 0.233093f $ **FLOATING
C431 phase_inverter_0/FILLER_0_9_72/a_2812_375# vss 0.17167f $ **FLOATING
C432 phase_inverter_0/FILLER_0_9_72/a_2364_375# vss 0.17167f $ **FLOATING
C433 phase_inverter_0/FILLER_0_9_72/a_1916_375# vss 0.17167f $ **FLOATING
C434 phase_inverter_0/FILLER_0_9_72/a_1468_375# vss 0.17167f $ **FLOATING
C435 phase_inverter_0/FILLER_0_9_72/a_1020_375# vss 0.17167f $ **FLOATING
C436 phase_inverter_0/FILLER_0_9_72/a_572_375# vss 0.17167f $ **FLOATING
C437 phase_inverter_0/FILLER_0_9_72/a_124_375# vss 0.185915f $ **FLOATING
C438 phase_inverter_0/FILLER_0_15_64/a_36_472# vss 0.417394f
C439 phase_inverter_0/FILLER_0_15_64/a_124_375# vss 0.246306f $ **FLOATING
C440 phase_inverter_0/_16_/Z vss 1.160526f
C441 phase_inverter_0/_16_/a_36_113# vss 0.418095f
C442 phase_inverter_0/FILLER_0_10_101/a_36_472# vss 0.417394f
C443 phase_inverter_0/FILLER_0_10_101/a_124_375# vss 0.246306f $ **FLOATING
C444 phase_inverter_0/FILLER_0_3_72/a_3172_472# vss 0.345058f $ **FLOATING
C445 phase_inverter_0/FILLER_0_3_72/a_2724_472# vss 0.33241f $ **FLOATING
C446 phase_inverter_0/FILLER_0_3_72/a_2276_472# vss 0.33241f $ **FLOATING
C447 phase_inverter_0/FILLER_0_3_72/a_1828_472# vss 0.33241f $ **FLOATING
C448 phase_inverter_0/FILLER_0_3_72/a_1380_472# vss 0.33241f $ **FLOATING
C449 phase_inverter_0/FILLER_0_3_72/a_932_472# vss 0.33241f $ **FLOATING
C450 phase_inverter_0/FILLER_0_3_72/a_484_472# vss 0.33241f $ **FLOATING
C451 phase_inverter_0/FILLER_0_3_72/a_36_472# vss 0.404746f
C452 phase_inverter_0/FILLER_0_3_72/a_3260_375# vss 0.233093f $ **FLOATING
C453 phase_inverter_0/FILLER_0_3_72/a_2812_375# vss 0.17167f $ **FLOATING
C454 phase_inverter_0/FILLER_0_3_72/a_2364_375# vss 0.17167f $ **FLOATING
C455 phase_inverter_0/FILLER_0_3_72/a_1916_375# vss 0.17167f $ **FLOATING
C456 phase_inverter_0/FILLER_0_3_72/a_1468_375# vss 0.17167f $ **FLOATING
C457 phase_inverter_0/FILLER_0_3_72/a_1020_375# vss 0.17167f $ **FLOATING
C458 phase_inverter_0/FILLER_0_3_72/a_572_375# vss 0.17167f $ **FLOATING
C459 phase_inverter_0/FILLER_0_3_72/a_124_375# vss 0.185915f $ **FLOATING
C460 phase_inverter_0/FILLER_0_8_28/a_36_472# vss 0.417394f
C461 phase_inverter_0/FILLER_0_8_28/a_124_375# vss 0.246306f $ **FLOATING
C462 phase_inverter_0/_17_/a_36_113# vss 0.418095f
C463 phase_inverter_0/FILLER_0_6_2/a_3172_472# vss 0.345058f $ **FLOATING
C464 phase_inverter_0/FILLER_0_6_2/a_2724_472# vss 0.33241f $ **FLOATING
C465 phase_inverter_0/FILLER_0_6_2/a_2276_472# vss 0.33241f $ **FLOATING
C466 phase_inverter_0/FILLER_0_6_2/a_1828_472# vss 0.33241f $ **FLOATING
C467 phase_inverter_0/FILLER_0_6_2/a_1380_472# vss 0.33241f $ **FLOATING
C468 phase_inverter_0/FILLER_0_6_2/a_932_472# vss 0.33241f $ **FLOATING
C469 phase_inverter_0/FILLER_0_6_2/a_484_472# vss 0.33241f $ **FLOATING
C470 phase_inverter_0/FILLER_0_6_2/a_36_472# vss 0.404746f
C471 phase_inverter_0/FILLER_0_6_2/a_3260_375# vss 0.233093f $ **FLOATING
C472 phase_inverter_0/FILLER_0_6_2/a_2812_375# vss 0.17167f $ **FLOATING
C473 phase_inverter_0/FILLER_0_6_2/a_2364_375# vss 0.17167f $ **FLOATING
C474 phase_inverter_0/FILLER_0_6_2/a_1916_375# vss 0.17167f $ **FLOATING
C475 phase_inverter_0/FILLER_0_6_2/a_1468_375# vss 0.17167f $ **FLOATING
C476 phase_inverter_0/FILLER_0_6_2/a_1020_375# vss 0.17167f $ **FLOATING
C477 phase_inverter_0/FILLER_0_6_2/a_572_375# vss 0.17167f $ **FLOATING
C478 phase_inverter_0/FILLER_0_6_2/a_124_375# vss 0.185915f $ **FLOATING
C479 phase_inverter_0/FILLER_0_15_40/a_1380_472# vss 0.345058f $ **FLOATING
C480 phase_inverter_0/FILLER_0_15_40/a_932_472# vss 0.33241f $ **FLOATING
C481 phase_inverter_0/FILLER_0_15_40/a_484_472# vss 0.33241f $ **FLOATING
C482 phase_inverter_0/FILLER_0_15_40/a_36_472# vss 0.404746f
C483 phase_inverter_0/FILLER_0_15_40/a_1468_375# vss 0.233029f
C484 phase_inverter_0/FILLER_0_15_40/a_1020_375# vss 0.171606f $ **FLOATING
C485 phase_inverter_0/FILLER_0_15_40/a_572_375# vss 0.171606f $ **FLOATING
C486 phase_inverter_0/FILLER_0_15_40/a_124_375# vss 0.185399f $ **FLOATING
C487 phase_inverter_0/_18_/a_36_113# vss 0.418095f
C488 phase_inverter_0/FILLER_0_3_60/a_484_472# vss 0.345058f $ **FLOATING
C489 phase_inverter_0/FILLER_0_3_60/a_36_472# vss 0.404746f
C490 phase_inverter_0/FILLER_0_3_60/a_572_375# vss 0.232991f
C491 phase_inverter_0/FILLER_0_3_60/a_124_375# vss 0.185089f $ **FLOATING
C492 phase_inverter_0/FILLER_0_14_107/a_484_472# vss 0.345058f $ **FLOATING
C493 phase_inverter_0/FILLER_0_14_107/a_36_472# vss 0.404746f
C494 phase_inverter_0/FILLER_0_14_107/a_572_375# vss 0.232991f
C495 phase_inverter_0/FILLER_0_14_107/a_124_375# vss 0.185089f $ **FLOATING
C496 phase_inverter_0/FILLER_0_15_72/a_1380_472# vss 0.345058f $ **FLOATING
C497 phase_inverter_0/FILLER_0_15_72/a_932_472# vss 0.33241f $ **FLOATING
C498 phase_inverter_0/FILLER_0_15_72/a_484_472# vss 0.333066f $ **FLOATING
C499 phase_inverter_0/FILLER_0_15_72/a_36_472# vss 0.404746f
C500 phase_inverter_0/FILLER_0_15_72/a_1468_375# vss 0.233029f
C501 phase_inverter_0/FILLER_0_15_72/a_1020_375# vss 0.171606f $ **FLOATING
C502 phase_inverter_0/FILLER_0_15_72/a_572_375# vss 0.171606f $ **FLOATING
C503 phase_inverter_0/FILLER_0_15_72/a_124_375# vss 0.185399f $ **FLOATING
C504 phase_inverter_0/_14_/I vss 1.424187f
C505 phase_inverter_0/FILLER_0_8_37/a_6756_472# vss 0.345058f $ **FLOATING
C506 phase_inverter_0/FILLER_0_8_37/a_6308_472# vss 0.33241f $ **FLOATING
C507 phase_inverter_0/FILLER_0_8_37/a_5860_472# vss 0.33241f $ **FLOATING
C508 phase_inverter_0/FILLER_0_8_37/a_5412_472# vss 0.33241f $ **FLOATING
C509 phase_inverter_0/FILLER_0_8_37/a_4964_472# vss 0.33241f $ **FLOATING
C510 phase_inverter_0/FILLER_0_8_37/a_4516_472# vss 0.33241f $ **FLOATING
C511 phase_inverter_0/FILLER_0_8_37/a_4068_472# vss 0.33241f $ **FLOATING
C512 phase_inverter_0/FILLER_0_8_37/a_3620_472# vss 0.33241f $ **FLOATING
C513 phase_inverter_0/FILLER_0_8_37/a_3172_472# vss 0.33241f $ **FLOATING
C514 phase_inverter_0/FILLER_0_8_37/a_2724_472# vss 0.33241f $ **FLOATING
C515 phase_inverter_0/FILLER_0_8_37/a_2276_472# vss 0.33241f $ **FLOATING
C516 phase_inverter_0/FILLER_0_8_37/a_1828_472# vss 0.33241f $ **FLOATING
C517 phase_inverter_0/FILLER_0_8_37/a_1380_472# vss 0.33241f $ **FLOATING
C518 phase_inverter_0/FILLER_0_8_37/a_932_472# vss 0.33241f $ **FLOATING
C519 phase_inverter_0/FILLER_0_8_37/a_484_472# vss 0.33241f $ **FLOATING
C520 phase_inverter_0/FILLER_0_8_37/a_36_472# vss 0.404746f
C521 phase_inverter_0/FILLER_0_8_37/a_6844_375# vss 0.233068f $ **FLOATING
C522 phase_inverter_0/FILLER_0_8_37/a_6396_375# vss 0.171644f $ **FLOATING
C523 phase_inverter_0/FILLER_0_8_37/a_5948_375# vss 0.171644f $ **FLOATING
C524 phase_inverter_0/FILLER_0_8_37/a_5500_375# vss 0.171644f $ **FLOATING
C525 phase_inverter_0/FILLER_0_8_37/a_5052_375# vss 0.171644f $ **FLOATING
C526 phase_inverter_0/FILLER_0_8_37/a_4604_375# vss 0.171644f $ **FLOATING
C527 phase_inverter_0/FILLER_0_8_37/a_4156_375# vss 0.171644f $ **FLOATING
C528 phase_inverter_0/FILLER_0_8_37/a_3708_375# vss 0.171644f $ **FLOATING
C529 phase_inverter_0/FILLER_0_8_37/a_3260_375# vss 0.171644f $ **FLOATING
C530 phase_inverter_0/FILLER_0_8_37/a_2812_375# vss 0.171644f $ **FLOATING
C531 phase_inverter_0/FILLER_0_8_37/a_2364_375# vss 0.171644f $ **FLOATING
C532 phase_inverter_0/FILLER_0_8_37/a_1916_375# vss 0.171644f $ **FLOATING
C533 phase_inverter_0/FILLER_0_8_37/a_1468_375# vss 0.171644f $ **FLOATING
C534 phase_inverter_0/FILLER_0_8_37/a_1020_375# vss 0.171644f $ **FLOATING
C535 phase_inverter_0/FILLER_0_8_37/a_572_375# vss 0.171644f $ **FLOATING
C536 phase_inverter_0/FILLER_0_8_37/a_124_375# vss 0.185708f $ **FLOATING
C537 phase_inverter_0/_19_/a_36_113# vss 0.418095f
C538 phase_inverter_0/FILLER_0_0_70/a_36_472# vss 0.417394f
C539 phase_inverter_0/FILLER_0_0_70/a_124_375# vss 0.246306f $ **FLOATING
C540 phase_inverter_0/FILLER_0_14_28/a_36_472# vss 0.417394f
C541 phase_inverter_0/FILLER_0_14_28/a_124_375# vss 0.246306f $ **FLOATING
C542 phase_inverter_0/FILLER_0_2_37/a_6756_472# vss 0.345058f $ **FLOATING
C543 phase_inverter_0/FILLER_0_2_37/a_6308_472# vss 0.33241f $ **FLOATING
C544 phase_inverter_0/FILLER_0_2_37/a_5860_472# vss 0.33241f $ **FLOATING
C545 phase_inverter_0/FILLER_0_2_37/a_5412_472# vss 0.33241f $ **FLOATING
C546 phase_inverter_0/FILLER_0_2_37/a_4964_472# vss 0.33241f $ **FLOATING
C547 phase_inverter_0/FILLER_0_2_37/a_4516_472# vss 0.33241f $ **FLOATING
C548 phase_inverter_0/FILLER_0_2_37/a_4068_472# vss 0.33241f $ **FLOATING
C549 phase_inverter_0/FILLER_0_2_37/a_3620_472# vss 0.33241f $ **FLOATING
C550 phase_inverter_0/FILLER_0_2_37/a_3172_472# vss 0.33241f $ **FLOATING
C551 phase_inverter_0/FILLER_0_2_37/a_2724_472# vss 0.33241f $ **FLOATING
C552 phase_inverter_0/FILLER_0_2_37/a_2276_472# vss 0.33241f $ **FLOATING
C553 phase_inverter_0/FILLER_0_2_37/a_1828_472# vss 0.33241f $ **FLOATING
C554 phase_inverter_0/FILLER_0_2_37/a_1380_472# vss 0.33241f $ **FLOATING
C555 phase_inverter_0/FILLER_0_2_37/a_932_472# vss 0.33241f $ **FLOATING
C556 phase_inverter_0/FILLER_0_2_37/a_484_472# vss 0.33241f $ **FLOATING
C557 phase_inverter_0/FILLER_0_2_37/a_36_472# vss 0.404746f
C558 phase_inverter_0/FILLER_0_2_37/a_6844_375# vss 0.233068f $ **FLOATING
C559 phase_inverter_0/FILLER_0_2_37/a_6396_375# vss 0.171644f $ **FLOATING
C560 phase_inverter_0/FILLER_0_2_37/a_5948_375# vss 0.171644f $ **FLOATING
C561 phase_inverter_0/FILLER_0_2_37/a_5500_375# vss 0.171644f $ **FLOATING
C562 phase_inverter_0/FILLER_0_2_37/a_5052_375# vss 0.171644f $ **FLOATING
C563 phase_inverter_0/FILLER_0_2_37/a_4604_375# vss 0.171644f $ **FLOATING
C564 phase_inverter_0/FILLER_0_2_37/a_4156_375# vss 0.171644f $ **FLOATING
C565 phase_inverter_0/FILLER_0_2_37/a_3708_375# vss 0.171644f $ **FLOATING
C566 phase_inverter_0/FILLER_0_2_37/a_3260_375# vss 0.171644f $ **FLOATING
C567 phase_inverter_0/FILLER_0_2_37/a_2812_375# vss 0.171644f $ **FLOATING
C568 phase_inverter_0/FILLER_0_2_37/a_2364_375# vss 0.171644f $ **FLOATING
C569 phase_inverter_0/FILLER_0_2_37/a_1916_375# vss 0.171644f $ **FLOATING
C570 phase_inverter_0/FILLER_0_2_37/a_1468_375# vss 0.171644f $ **FLOATING
C571 phase_inverter_0/FILLER_0_2_37/a_1020_375# vss 0.171644f $ **FLOATING
C572 phase_inverter_0/FILLER_0_2_37/a_572_375# vss 0.171644f $ **FLOATING
C573 phase_inverter_0/FILLER_0_2_37/a_124_375# vss 0.185708f $ **FLOATING
C574 input_signal[9] vss 1.722228f
C575 phase_inverter_0/FILLER_0_3_104/a_484_472# vss 0.345058f $ **FLOATING
C576 phase_inverter_0/FILLER_0_3_104/a_36_472# vss 0.404746f
C577 phase_inverter_0/FILLER_0_3_104/a_572_375# vss 0.232991f
C578 phase_inverter_0/FILLER_0_3_104/a_124_375# vss 0.185089f $ **FLOATING
C579 phase_inverter_0/FILLER_0_6_101/a_36_472# vss 0.417394f
C580 phase_inverter_0/FILLER_0_6_101/a_124_375# vss 0.246306f $ **FLOATING
C581 phase_inverter_0/FILLER_0_14_115/a_36_472# vss 0.417394f
C582 phase_inverter_0/FILLER_0_14_115/a_124_375# vss 0.246306f $ **FLOATING
C583 phase_inverter_0/input9/a_36_113# vss 0.418095f
C584 phase_inverter_0/FILLER_0_8_12/a_1380_472# vss 0.345058f $ **FLOATING
C585 phase_inverter_0/FILLER_0_8_12/a_932_472# vss 0.33241f $ **FLOATING
C586 phase_inverter_0/FILLER_0_8_12/a_484_472# vss 0.33241f $ **FLOATING
C587 phase_inverter_0/FILLER_0_8_12/a_36_472# vss 0.404746f
C588 phase_inverter_0/FILLER_0_8_12/a_1468_375# vss 0.233029f
C589 phase_inverter_0/FILLER_0_8_12/a_1020_375# vss 0.171606f $ **FLOATING
C590 phase_inverter_0/FILLER_0_8_12/a_572_375# vss 0.171606f $ **FLOATING
C591 phase_inverter_0/FILLER_0_8_12/a_124_375# vss 0.185399f $ **FLOATING
C592 phase_inverter_0/FILLER_0_14_37/a_6756_472# vss 0.345058f $ **FLOATING
C593 phase_inverter_0/FILLER_0_14_37/a_6308_472# vss 0.33241f $ **FLOATING
C594 phase_inverter_0/FILLER_0_14_37/a_5860_472# vss 0.33241f $ **FLOATING
C595 phase_inverter_0/FILLER_0_14_37/a_5412_472# vss 0.33241f $ **FLOATING
C596 phase_inverter_0/FILLER_0_14_37/a_4964_472# vss 0.33241f $ **FLOATING
C597 phase_inverter_0/FILLER_0_14_37/a_4516_472# vss 0.33241f $ **FLOATING
C598 phase_inverter_0/FILLER_0_14_37/a_4068_472# vss 0.33241f $ **FLOATING
C599 phase_inverter_0/FILLER_0_14_37/a_3620_472# vss 0.33241f $ **FLOATING
C600 phase_inverter_0/FILLER_0_14_37/a_3172_472# vss 0.33241f $ **FLOATING
C601 phase_inverter_0/FILLER_0_14_37/a_2724_472# vss 0.33241f $ **FLOATING
C602 phase_inverter_0/FILLER_0_14_37/a_2276_472# vss 0.33241f $ **FLOATING
C603 phase_inverter_0/FILLER_0_14_37/a_1828_472# vss 0.33241f $ **FLOATING
C604 phase_inverter_0/FILLER_0_14_37/a_1380_472# vss 0.33241f $ **FLOATING
C605 phase_inverter_0/FILLER_0_14_37/a_932_472# vss 0.33241f $ **FLOATING
C606 phase_inverter_0/FILLER_0_14_37/a_484_472# vss 0.33241f $ **FLOATING
C607 phase_inverter_0/FILLER_0_14_37/a_36_472# vss 0.404746f
C608 phase_inverter_0/FILLER_0_14_37/a_6844_375# vss 0.233068f $ **FLOATING
C609 phase_inverter_0/FILLER_0_14_37/a_6396_375# vss 0.171644f $ **FLOATING
C610 phase_inverter_0/FILLER_0_14_37/a_5948_375# vss 0.171644f $ **FLOATING
C611 phase_inverter_0/FILLER_0_14_37/a_5500_375# vss 0.171644f $ **FLOATING
C612 phase_inverter_0/FILLER_0_14_37/a_5052_375# vss 0.171644f $ **FLOATING
C613 phase_inverter_0/FILLER_0_14_37/a_4604_375# vss 0.171644f $ **FLOATING
C614 phase_inverter_0/FILLER_0_14_37/a_4156_375# vss 0.171644f $ **FLOATING
C615 phase_inverter_0/FILLER_0_14_37/a_3708_375# vss 0.171644f $ **FLOATING
C616 phase_inverter_0/FILLER_0_14_37/a_3260_375# vss 0.171644f $ **FLOATING
C617 phase_inverter_0/FILLER_0_14_37/a_2812_375# vss 0.171644f $ **FLOATING
C618 phase_inverter_0/FILLER_0_14_37/a_2364_375# vss 0.171644f $ **FLOATING
C619 phase_inverter_0/FILLER_0_14_37/a_1916_375# vss 0.171644f $ **FLOATING
C620 phase_inverter_0/FILLER_0_14_37/a_1468_375# vss 0.171644f $ **FLOATING
C621 phase_inverter_0/FILLER_0_14_37/a_1020_375# vss 0.171644f $ **FLOATING
C622 phase_inverter_0/FILLER_0_14_37/a_572_375# vss 0.171644f $ **FLOATING
C623 phase_inverter_0/FILLER_0_14_37/a_124_375# vss 0.185708f $ **FLOATING
C624 phase_inverter_0/input8/a_36_113# vss 0.418095f
C625 phase_inverter_0/FILLER_0_5_12/a_3172_472# vss 0.345058f $ **FLOATING
C626 phase_inverter_0/FILLER_0_5_12/a_2724_472# vss 0.33241f $ **FLOATING
C627 phase_inverter_0/FILLER_0_5_12/a_2276_472# vss 0.33241f $ **FLOATING
C628 phase_inverter_0/FILLER_0_5_12/a_1828_472# vss 0.33241f $ **FLOATING
C629 phase_inverter_0/FILLER_0_5_12/a_1380_472# vss 0.33241f $ **FLOATING
C630 phase_inverter_0/FILLER_0_5_12/a_932_472# vss 0.33241f $ **FLOATING
C631 phase_inverter_0/FILLER_0_5_12/a_484_472# vss 0.33241f $ **FLOATING
C632 phase_inverter_0/FILLER_0_5_12/a_36_472# vss 0.404746f
C633 phase_inverter_0/FILLER_0_5_12/a_3260_375# vss 0.233093f $ **FLOATING
C634 phase_inverter_0/FILLER_0_5_12/a_2812_375# vss 0.17167f $ **FLOATING
C635 phase_inverter_0/FILLER_0_5_12/a_2364_375# vss 0.17167f $ **FLOATING
C636 phase_inverter_0/FILLER_0_5_12/a_1916_375# vss 0.17167f $ **FLOATING
C637 phase_inverter_0/FILLER_0_5_12/a_1468_375# vss 0.17167f $ **FLOATING
C638 phase_inverter_0/FILLER_0_5_12/a_1020_375# vss 0.17167f $ **FLOATING
C639 phase_inverter_0/FILLER_0_5_12/a_572_375# vss 0.17167f $ **FLOATING
C640 phase_inverter_0/FILLER_0_5_12/a_124_375# vss 0.185915f $ **FLOATING
C641 phase_inverter_0/input10/a_36_113# vss 0.418095f
C642 phase_inverter_0/FILLER_0_5_44/a_1380_472# vss 0.345058f $ **FLOATING
C643 phase_inverter_0/FILLER_0_5_44/a_932_472# vss 0.33241f $ **FLOATING
C644 phase_inverter_0/FILLER_0_5_44/a_484_472# vss 0.33241f $ **FLOATING
C645 phase_inverter_0/FILLER_0_5_44/a_36_472# vss 0.404746f
C646 phase_inverter_0/FILLER_0_5_44/a_1468_375# vss 0.233029f
C647 phase_inverter_0/FILLER_0_5_44/a_1020_375# vss 0.171606f $ **FLOATING
C648 phase_inverter_0/FILLER_0_5_44/a_572_375# vss 0.171606f $ **FLOATING
C649 phase_inverter_0/FILLER_0_5_44/a_124_375# vss 0.185399f $ **FLOATING
C650 phase_inverter_0/input7/a_36_113# vss 0.418095f
C651 phase_inverter_0/FILLER_0_0_104/a_36_472# vss 0.417394f
C652 phase_inverter_0/FILLER_0_0_104/a_124_375# vss 0.246306f $ **FLOATING
C653 input_signal[5] vss 1.048828f
C654 phase_inverter_0/input6/a_36_113# vss 0.418095f
C655 phase_inverter_0/FILLER_0_14_101/a_36_472# vss 0.417394f
C656 phase_inverter_0/FILLER_0_14_101/a_124_375# vss 0.246306f $ **FLOATING
C657 phase_inverter_0/FILLER_0_14_12/a_1380_472# vss 0.345058f $ **FLOATING
C658 phase_inverter_0/FILLER_0_14_12/a_932_472# vss 0.33241f $ **FLOATING
C659 phase_inverter_0/FILLER_0_14_12/a_484_472# vss 0.33241f $ **FLOATING
C660 phase_inverter_0/FILLER_0_14_12/a_36_472# vss 0.404746f
C661 phase_inverter_0/FILLER_0_14_12/a_1468_375# vss 0.233029f
C662 phase_inverter_0/FILLER_0_14_12/a_1020_375# vss 0.171606f $ **FLOATING
C663 phase_inverter_0/FILLER_0_14_12/a_572_375# vss 0.171606f $ **FLOATING
C664 phase_inverter_0/FILLER_0_14_12/a_124_375# vss 0.185399f $ **FLOATING
C665 phase_inverter_0/FILLER_0_11_136/a_36_472# vss 0.417394f
C666 phase_inverter_0/FILLER_0_11_136/a_124_375# vss 0.246306f $ **FLOATING
C667 phase_inverter_0/input5/a_36_113# vss 0.418095f
C668 phase_inverter_0/_19_/I vss 1.019585f
C669 input_signal[3] vss 0.969415f
C670 phase_inverter_0/input4/a_36_113# vss 0.418095f
C671 phase_inverter_0/FILLER_0_11_66/a_36_472# vss 0.417394f
C672 phase_inverter_0/FILLER_0_11_66/a_124_375# vss 0.246306f $ **FLOATING
C673 phase_inverter_0/_12_/I vss 1.059653f
C674 phase_inverter_0/input3/a_36_113# vss 0.418095f
C675 phase_inverter_0/_11_/I vss 1.493507f
C676 input_signal[1] vss 1.033314f
C677 phase_inverter_0/input2/a_36_113# vss 0.418095f
C678 phase_inverter_0/FILLER_0_5_72/a_3172_472# vss 0.345058f $ **FLOATING
C679 phase_inverter_0/FILLER_0_5_72/a_2724_472# vss 0.33241f $ **FLOATING
C680 phase_inverter_0/FILLER_0_5_72/a_2276_472# vss 0.33241f $ **FLOATING
C681 phase_inverter_0/FILLER_0_5_72/a_1828_472# vss 0.33241f $ **FLOATING
C682 phase_inverter_0/FILLER_0_5_72/a_1380_472# vss 0.33241f $ **FLOATING
C683 phase_inverter_0/FILLER_0_5_72/a_932_472# vss 0.33241f $ **FLOATING
C684 phase_inverter_0/FILLER_0_5_72/a_484_472# vss 0.33241f $ **FLOATING
C685 phase_inverter_0/FILLER_0_5_72/a_36_472# vss 0.404746f
C686 phase_inverter_0/FILLER_0_5_72/a_3260_375# vss 0.233093f $ **FLOATING
C687 phase_inverter_0/FILLER_0_5_72/a_2812_375# vss 0.17167f $ **FLOATING
C688 phase_inverter_0/FILLER_0_5_72/a_2364_375# vss 0.17167f $ **FLOATING
C689 phase_inverter_0/FILLER_0_5_72/a_1916_375# vss 0.17167f $ **FLOATING
C690 phase_inverter_0/FILLER_0_5_72/a_1468_375# vss 0.17167f $ **FLOATING
C691 phase_inverter_0/FILLER_0_5_72/a_1020_375# vss 0.17167f $ **FLOATING
C692 phase_inverter_0/FILLER_0_5_72/a_572_375# vss 0.17167f $ **FLOATING
C693 phase_inverter_0/FILLER_0_5_72/a_124_375# vss 0.185915f $ **FLOATING
C694 phase_inverter_0/FILLER_0_4_107/a_1380_472# vss 0.345058f $ **FLOATING
C695 phase_inverter_0/FILLER_0_4_107/a_932_472# vss 0.33241f $ **FLOATING
C696 phase_inverter_0/FILLER_0_4_107/a_484_472# vss 0.33241f $ **FLOATING
C697 phase_inverter_0/FILLER_0_4_107/a_36_472# vss 0.404746f
C698 phase_inverter_0/FILLER_0_4_107/a_1468_375# vss 0.233029f
C699 phase_inverter_0/FILLER_0_4_107/a_1020_375# vss 0.171606f $ **FLOATING
C700 phase_inverter_0/FILLER_0_4_107/a_572_375# vss 0.171606f $ **FLOATING
C701 phase_inverter_0/FILLER_0_4_107/a_124_375# vss 0.185399f $ **FLOATING
C702 phase_inverter_0/_10_/I vss 0.979826f
C703 input_signal[0] vss 1.665667f
C704 phase_inverter_0/input1/a_36_113# vss 0.418095f
C705 phase_inverter_0/_03_/ZN vss 1.105776f
C706 phase_inverter_0/FILLER_0_7_104/a_484_472# vss 0.345058f $ **FLOATING
C707 phase_inverter_0/FILLER_0_7_104/a_36_472# vss 0.404746f
C708 phase_inverter_0/FILLER_0_7_104/a_572_375# vss 0.232991f
C709 phase_inverter_0/FILLER_0_7_104/a_124_375# vss 0.185089f $ **FLOATING
C710 phase_inverter_0/FILLER_0_5_60/a_484_472# vss 0.345058f $ **FLOATING
C711 phase_inverter_0/FILLER_0_5_60/a_36_472# vss 0.404746f
C712 phase_inverter_0/FILLER_0_5_60/a_572_375# vss 0.232991f
C713 phase_inverter_0/FILLER_0_5_60/a_124_375# vss 0.185089f $ **FLOATING
C714 phase_inverter_0/FILLER_0_0_142/a_484_472# vss 0.345058f $ **FLOATING
C715 phase_inverter_0/FILLER_0_0_142/a_36_472# vss 0.404746f
C716 phase_inverter_0/FILLER_0_0_142/a_572_375# vss 0.232991f
C717 phase_inverter_0/FILLER_0_0_142/a_124_375# vss 0.185089f $ **FLOATING
C718 phase_inverter_0/_04_/ZN vss 1.111802f
C719 input_signal[7] vss 0.974241f
C720 phase_inverter_0/FILLER_0_16_18/a_1380_472# vss 0.345058f $ **FLOATING
C721 phase_inverter_0/FILLER_0_16_18/a_932_472# vss 0.33241f $ **FLOATING
C722 phase_inverter_0/FILLER_0_16_18/a_484_472# vss 0.33241f $ **FLOATING
C723 phase_inverter_0/FILLER_0_16_18/a_36_472# vss 0.404746f
C724 phase_inverter_0/FILLER_0_16_18/a_1468_375# vss 0.233029f
C725 phase_inverter_0/FILLER_0_16_18/a_1020_375# vss 0.171606f $ **FLOATING
C726 phase_inverter_0/FILLER_0_16_18/a_572_375# vss 0.171606f $ **FLOATING
C727 phase_inverter_0/FILLER_0_16_18/a_124_375# vss 0.185399f $ **FLOATING
C728 phase_inverter_0/net15 vss 1.058175f
C729 phase_inverter_0/_09_/ZN vss 1.363364f
C730 phase_inverter_0/output19/a_224_472# vss 2.38465f
C731 phase_inverter_0/_13_/I vss 1.115417f
C732 phase_inverter_0/FILLER_0_11_72/a_6756_472# vss 0.345058f $ **FLOATING
C733 phase_inverter_0/FILLER_0_11_72/a_6308_472# vss 0.33241f $ **FLOATING
C734 phase_inverter_0/FILLER_0_11_72/a_5860_472# vss 0.33241f $ **FLOATING
C735 phase_inverter_0/FILLER_0_11_72/a_5412_472# vss 0.33241f $ **FLOATING
C736 phase_inverter_0/FILLER_0_11_72/a_4964_472# vss 0.33241f $ **FLOATING
C737 phase_inverter_0/FILLER_0_11_72/a_4516_472# vss 0.33241f $ **FLOATING
C738 phase_inverter_0/FILLER_0_11_72/a_4068_472# vss 0.33241f $ **FLOATING
C739 phase_inverter_0/FILLER_0_11_72/a_3620_472# vss 0.33241f $ **FLOATING
C740 phase_inverter_0/FILLER_0_11_72/a_3172_472# vss 0.33241f $ **FLOATING
C741 phase_inverter_0/FILLER_0_11_72/a_2724_472# vss 0.33241f $ **FLOATING
C742 phase_inverter_0/FILLER_0_11_72/a_2276_472# vss 0.33241f $ **FLOATING
C743 phase_inverter_0/FILLER_0_11_72/a_1828_472# vss 0.33241f $ **FLOATING
C744 phase_inverter_0/FILLER_0_11_72/a_1380_472# vss 0.33241f $ **FLOATING
C745 phase_inverter_0/FILLER_0_11_72/a_932_472# vss 0.33241f $ **FLOATING
C746 phase_inverter_0/FILLER_0_11_72/a_484_472# vss 0.33241f $ **FLOATING
C747 phase_inverter_0/FILLER_0_11_72/a_36_472# vss 0.404746f
C748 phase_inverter_0/FILLER_0_11_72/a_6844_375# vss 0.233068f $ **FLOATING
C749 phase_inverter_0/FILLER_0_11_72/a_6396_375# vss 0.171644f $ **FLOATING
C750 phase_inverter_0/FILLER_0_11_72/a_5948_375# vss 0.171644f $ **FLOATING
C751 phase_inverter_0/FILLER_0_11_72/a_5500_375# vss 0.171644f $ **FLOATING
C752 phase_inverter_0/FILLER_0_11_72/a_5052_375# vss 0.171644f $ **FLOATING
C753 phase_inverter_0/FILLER_0_11_72/a_4604_375# vss 0.171644f $ **FLOATING
C754 phase_inverter_0/FILLER_0_11_72/a_4156_375# vss 0.171644f $ **FLOATING
C755 phase_inverter_0/FILLER_0_11_72/a_3708_375# vss 0.171644f $ **FLOATING
C756 phase_inverter_0/FILLER_0_11_72/a_3260_375# vss 0.171644f $ **FLOATING
C757 phase_inverter_0/FILLER_0_11_72/a_2812_375# vss 0.171644f $ **FLOATING
C758 phase_inverter_0/FILLER_0_11_72/a_2364_375# vss 0.171644f $ **FLOATING
C759 phase_inverter_0/FILLER_0_11_72/a_1916_375# vss 0.171644f $ **FLOATING
C760 phase_inverter_0/FILLER_0_11_72/a_1468_375# vss 0.171644f $ **FLOATING
C761 phase_inverter_0/FILLER_0_11_72/a_1020_375# vss 0.171644f $ **FLOATING
C762 phase_inverter_0/FILLER_0_11_72/a_572_375# vss 0.171644f $ **FLOATING
C763 phase_inverter_0/FILLER_0_11_72/a_124_375# vss 0.185708f $ **FLOATING
C764 phase_inverter_0/FILLER_0_4_37/a_6756_472# vss 0.345058f $ **FLOATING
C765 phase_inverter_0/FILLER_0_4_37/a_6308_472# vss 0.33241f $ **FLOATING
C766 phase_inverter_0/FILLER_0_4_37/a_5860_472# vss 0.33241f $ **FLOATING
C767 phase_inverter_0/FILLER_0_4_37/a_5412_472# vss 0.33241f $ **FLOATING
C768 phase_inverter_0/FILLER_0_4_37/a_4964_472# vss 0.33241f $ **FLOATING
C769 phase_inverter_0/FILLER_0_4_37/a_4516_472# vss 0.33241f $ **FLOATING
C770 phase_inverter_0/FILLER_0_4_37/a_4068_472# vss 0.33241f $ **FLOATING
C771 phase_inverter_0/FILLER_0_4_37/a_3620_472# vss 0.33241f $ **FLOATING
C772 phase_inverter_0/FILLER_0_4_37/a_3172_472# vss 0.33241f $ **FLOATING
C773 phase_inverter_0/FILLER_0_4_37/a_2724_472# vss 0.33241f $ **FLOATING
C774 phase_inverter_0/FILLER_0_4_37/a_2276_472# vss 0.33241f $ **FLOATING
C775 phase_inverter_0/FILLER_0_4_37/a_1828_472# vss 0.33241f $ **FLOATING
C776 phase_inverter_0/FILLER_0_4_37/a_1380_472# vss 0.33241f $ **FLOATING
C777 phase_inverter_0/FILLER_0_4_37/a_932_472# vss 0.33241f $ **FLOATING
C778 phase_inverter_0/FILLER_0_4_37/a_484_472# vss 0.33241f $ **FLOATING
C779 phase_inverter_0/FILLER_0_4_37/a_36_472# vss 0.404746f
C780 phase_inverter_0/FILLER_0_4_37/a_6844_375# vss 0.233068f $ **FLOATING
C781 phase_inverter_0/FILLER_0_4_37/a_6396_375# vss 0.171644f $ **FLOATING
C782 phase_inverter_0/FILLER_0_4_37/a_5948_375# vss 0.171644f $ **FLOATING
C783 phase_inverter_0/FILLER_0_4_37/a_5500_375# vss 0.171644f $ **FLOATING
C784 phase_inverter_0/FILLER_0_4_37/a_5052_375# vss 0.171644f $ **FLOATING
C785 phase_inverter_0/FILLER_0_4_37/a_4604_375# vss 0.171644f $ **FLOATING
C786 phase_inverter_0/FILLER_0_4_37/a_4156_375# vss 0.171644f $ **FLOATING
C787 phase_inverter_0/FILLER_0_4_37/a_3708_375# vss 0.171644f $ **FLOATING
C788 phase_inverter_0/FILLER_0_4_37/a_3260_375# vss 0.171644f $ **FLOATING
C789 phase_inverter_0/FILLER_0_4_37/a_2812_375# vss 0.171644f $ **FLOATING
C790 phase_inverter_0/FILLER_0_4_37/a_2364_375# vss 0.171644f $ **FLOATING
C791 phase_inverter_0/FILLER_0_4_37/a_1916_375# vss 0.171644f $ **FLOATING
C792 phase_inverter_0/FILLER_0_4_37/a_1468_375# vss 0.171644f $ **FLOATING
C793 phase_inverter_0/FILLER_0_4_37/a_1020_375# vss 0.171644f $ **FLOATING
C794 phase_inverter_0/FILLER_0_4_37/a_572_375# vss 0.171644f $ **FLOATING
C795 phase_inverter_0/FILLER_0_4_37/a_124_375# vss 0.185708f $ **FLOATING
C796 phase_inverter_0/_08_/ZN vss 1.295594f
C797 phase_inverter_0/output18/a_224_472# vss 2.39122f
C798 phase_inverter_0/_15_/I vss 1.113137f
C799 phase_inverter_0/_18_/Z vss 1.167483f
C800 phase_inverter_0/output29/a_224_472# vss 2.38465f
C801 phase_inverter_0/FILLER_0_12_107/a_1380_472# vss 0.345058f $ **FLOATING
C802 phase_inverter_0/FILLER_0_12_107/a_932_472# vss 0.33241f $ **FLOATING
C803 phase_inverter_0/FILLER_0_12_107/a_484_472# vss 0.33241f $ **FLOATING
C804 phase_inverter_0/FILLER_0_12_107/a_36_472# vss 0.404746f
C805 phase_inverter_0/FILLER_0_12_107/a_1468_375# vss 0.233029f
C806 phase_inverter_0/FILLER_0_12_107/a_1020_375# vss 0.171606f $ **FLOATING
C807 phase_inverter_0/FILLER_0_12_107/a_572_375# vss 0.171606f $ **FLOATING
C808 phase_inverter_0/FILLER_0_12_107/a_124_375# vss 0.185399f $ **FLOATING
C809 phase_inverter_0/FILLER_0_10_28/a_36_472# vss 0.417394f
C810 phase_inverter_0/FILLER_0_10_28/a_124_375# vss 0.246306f $ **FLOATING
C811 phase_inverter_0/_07_/ZN vss 1.113234f
C812 phase_inverter_0/output17/a_224_472# vss 2.38465f
C813 phase_inverter_0/_16_/I vss 0.912843f
C814 phase_inverter_0/_17_/Z vss 1.120758f
C815 phase_inverter_0/output28/a_224_472# vss 2.38465f
C816 phase_inverter_0/_06_/ZN vss 1.134591f
C817 phase_inverter_0/output16/a_224_472# vss 2.38465f
C818 phase_inverter_0/output27/a_224_472# vss 2.38465f
C819 phase_inverter_0/_17_/I vss 0.917813f
C820 phase_inverter_0/FILLER_0_16_36/a_3172_472# vss 0.345058f $ **FLOATING
C821 phase_inverter_0/FILLER_0_16_36/a_2724_472# vss 0.33241f $ **FLOATING
C822 phase_inverter_0/FILLER_0_16_36/a_2276_472# vss 0.33241f $ **FLOATING
C823 phase_inverter_0/FILLER_0_16_36/a_1828_472# vss 0.33241f $ **FLOATING
C824 phase_inverter_0/FILLER_0_16_36/a_1380_472# vss 0.33241f $ **FLOATING
C825 phase_inverter_0/FILLER_0_16_36/a_932_472# vss 0.33241f $ **FLOATING
C826 phase_inverter_0/FILLER_0_16_36/a_484_472# vss 0.33241f $ **FLOATING
C827 phase_inverter_0/FILLER_0_16_36/a_36_472# vss 0.404746f
C828 phase_inverter_0/FILLER_0_16_36/a_3260_375# vss 0.233093f $ **FLOATING
C829 phase_inverter_0/FILLER_0_16_36/a_2812_375# vss 0.17167f $ **FLOATING
C830 phase_inverter_0/FILLER_0_16_36/a_2364_375# vss 0.17167f $ **FLOATING
C831 phase_inverter_0/FILLER_0_16_36/a_1916_375# vss 0.17167f $ **FLOATING
C832 phase_inverter_0/FILLER_0_16_36/a_1468_375# vss 0.17167f $ **FLOATING
C833 phase_inverter_0/FILLER_0_16_36/a_1020_375# vss 0.17167f $ **FLOATING
C834 phase_inverter_0/FILLER_0_16_36/a_572_375# vss 0.17167f $ **FLOATING
C835 phase_inverter_0/FILLER_0_16_36/a_124_375# vss 0.190644f $ **FLOATING
C836 phase_inverter_0/FILLER_0_10_37/a_6756_472# vss 0.345058f $ **FLOATING
C837 phase_inverter_0/FILLER_0_10_37/a_6308_472# vss 0.33241f $ **FLOATING
C838 phase_inverter_0/FILLER_0_10_37/a_5860_472# vss 0.33241f $ **FLOATING
C839 phase_inverter_0/FILLER_0_10_37/a_5412_472# vss 0.33241f $ **FLOATING
C840 phase_inverter_0/FILLER_0_10_37/a_4964_472# vss 0.33241f $ **FLOATING
C841 phase_inverter_0/FILLER_0_10_37/a_4516_472# vss 0.33241f $ **FLOATING
C842 phase_inverter_0/FILLER_0_10_37/a_4068_472# vss 0.33241f $ **FLOATING
C843 phase_inverter_0/FILLER_0_10_37/a_3620_472# vss 0.33241f $ **FLOATING
C844 phase_inverter_0/FILLER_0_10_37/a_3172_472# vss 0.33241f $ **FLOATING
C845 phase_inverter_0/FILLER_0_10_37/a_2724_472# vss 0.33241f $ **FLOATING
C846 phase_inverter_0/FILLER_0_10_37/a_2276_472# vss 0.33241f $ **FLOATING
C847 phase_inverter_0/FILLER_0_10_37/a_1828_472# vss 0.33241f $ **FLOATING
C848 phase_inverter_0/FILLER_0_10_37/a_1380_472# vss 0.33241f $ **FLOATING
C849 phase_inverter_0/FILLER_0_10_37/a_932_472# vss 0.33241f $ **FLOATING
C850 phase_inverter_0/FILLER_0_10_37/a_484_472# vss 0.33241f $ **FLOATING
C851 phase_inverter_0/FILLER_0_10_37/a_36_472# vss 0.404746f
C852 phase_inverter_0/FILLER_0_10_37/a_6844_375# vss 0.233068f $ **FLOATING
C853 phase_inverter_0/FILLER_0_10_37/a_6396_375# vss 0.171644f $ **FLOATING
C854 phase_inverter_0/FILLER_0_10_37/a_5948_375# vss 0.171644f $ **FLOATING
C855 phase_inverter_0/FILLER_0_10_37/a_5500_375# vss 0.171644f $ **FLOATING
C856 phase_inverter_0/FILLER_0_10_37/a_5052_375# vss 0.171644f $ **FLOATING
C857 phase_inverter_0/FILLER_0_10_37/a_4604_375# vss 0.171644f $ **FLOATING
C858 phase_inverter_0/FILLER_0_10_37/a_4156_375# vss 0.171644f $ **FLOATING
C859 phase_inverter_0/FILLER_0_10_37/a_3708_375# vss 0.171644f $ **FLOATING
C860 phase_inverter_0/FILLER_0_10_37/a_3260_375# vss 0.171644f $ **FLOATING
C861 phase_inverter_0/FILLER_0_10_37/a_2812_375# vss 0.171644f $ **FLOATING
C862 phase_inverter_0/FILLER_0_10_37/a_2364_375# vss 0.171644f $ **FLOATING
C863 phase_inverter_0/FILLER_0_10_37/a_1916_375# vss 0.171644f $ **FLOATING
C864 phase_inverter_0/FILLER_0_10_37/a_1468_375# vss 0.171644f $ **FLOATING
C865 phase_inverter_0/FILLER_0_10_37/a_1020_375# vss 0.171644f $ **FLOATING
C866 phase_inverter_0/FILLER_0_10_37/a_572_375# vss 0.171644f $ **FLOATING
C867 phase_inverter_0/FILLER_0_10_37/a_124_375# vss 0.185708f $ **FLOATING
C868 phase_inverter_0/FILLER_0_7_66/a_36_472# vss 0.417394f
C869 phase_inverter_0/FILLER_0_7_66/a_124_375# vss 0.246306f $ **FLOATING
C870 phase_inverter_0/FILLER_0_4_101/a_36_472# vss 0.417394f
C871 phase_inverter_0/FILLER_0_4_101/a_124_375# vss 0.246306f $ **FLOATING
C872 phase_inverter_0/output15/a_224_472# vss 2.38465f
C873 phase_inverter_0/_18_/I vss 0.865773f
C874 phase_inverter_0/output26/a_224_472# vss 2.38465f
C875 phase_inverter_0/FILLER_0_1_12/a_3172_472# vss 0.345058f $ **FLOATING
C876 phase_inverter_0/FILLER_0_1_12/a_2724_472# vss 0.33241f $ **FLOATING
C877 phase_inverter_0/FILLER_0_1_12/a_2276_472# vss 0.33241f $ **FLOATING
C878 phase_inverter_0/FILLER_0_1_12/a_1828_472# vss 0.33241f $ **FLOATING
C879 phase_inverter_0/FILLER_0_1_12/a_1380_472# vss 0.33241f $ **FLOATING
C880 phase_inverter_0/FILLER_0_1_12/a_932_472# vss 0.33241f $ **FLOATING
C881 phase_inverter_0/FILLER_0_1_12/a_484_472# vss 0.33241f $ **FLOATING
C882 phase_inverter_0/FILLER_0_1_12/a_36_472# vss 0.404746f
C883 phase_inverter_0/FILLER_0_1_12/a_3260_375# vss 0.233093f $ **FLOATING
C884 phase_inverter_0/FILLER_0_1_12/a_2812_375# vss 0.17167f $ **FLOATING
C885 phase_inverter_0/FILLER_0_1_12/a_2364_375# vss 0.17167f $ **FLOATING
C886 phase_inverter_0/FILLER_0_1_12/a_1916_375# vss 0.17167f $ **FLOATING
C887 phase_inverter_0/FILLER_0_1_12/a_1468_375# vss 0.17167f $ **FLOATING
C888 phase_inverter_0/FILLER_0_1_12/a_1020_375# vss 0.17167f $ **FLOATING
C889 phase_inverter_0/FILLER_0_1_12/a_572_375# vss 0.17167f $ **FLOATING
C890 phase_inverter_0/FILLER_0_1_12/a_124_375# vss 0.185915f $ **FLOATING
C891 phase_inverter_0/output14/a_224_472# vss 2.38465f
C892 phase_inverter_0/output25/a_224_472# vss 2.38465f
C893 phase_inverter_0/FILLER_0_1_44/a_1380_472# vss 0.345058f $ **FLOATING
C894 phase_inverter_0/FILLER_0_1_44/a_932_472# vss 0.33241f $ **FLOATING
C895 phase_inverter_0/FILLER_0_1_44/a_484_472# vss 0.33241f $ **FLOATING
C896 phase_inverter_0/FILLER_0_1_44/a_36_472# vss 0.404746f
C897 phase_inverter_0/FILLER_0_1_44/a_1468_375# vss 0.233029f
C898 phase_inverter_0/FILLER_0_1_44/a_1020_375# vss 0.171606f $ **FLOATING
C899 phase_inverter_0/FILLER_0_1_44/a_572_375# vss 0.171606f $ **FLOATING
C900 phase_inverter_0/FILLER_0_1_44/a_124_375# vss 0.185399f $ **FLOATING
C901 phase_inverter_0/FILLER_0_7_2/a_6756_472# vss 0.345058f $ **FLOATING
C902 phase_inverter_0/FILLER_0_7_2/a_6308_472# vss 0.33241f $ **FLOATING
C903 phase_inverter_0/FILLER_0_7_2/a_5860_472# vss 0.33241f $ **FLOATING
C904 phase_inverter_0/FILLER_0_7_2/a_5412_472# vss 0.33241f $ **FLOATING
C905 phase_inverter_0/FILLER_0_7_2/a_4964_472# vss 0.33241f $ **FLOATING
C906 phase_inverter_0/FILLER_0_7_2/a_4516_472# vss 0.33241f $ **FLOATING
C907 phase_inverter_0/FILLER_0_7_2/a_4068_472# vss 0.33241f $ **FLOATING
C908 phase_inverter_0/FILLER_0_7_2/a_3620_472# vss 0.33241f $ **FLOATING
C909 phase_inverter_0/FILLER_0_7_2/a_3172_472# vss 0.33241f $ **FLOATING
C910 phase_inverter_0/FILLER_0_7_2/a_2724_472# vss 0.33241f $ **FLOATING
C911 phase_inverter_0/FILLER_0_7_2/a_2276_472# vss 0.33241f $ **FLOATING
C912 phase_inverter_0/FILLER_0_7_2/a_1828_472# vss 0.33241f $ **FLOATING
C913 phase_inverter_0/FILLER_0_7_2/a_1380_472# vss 0.33241f $ **FLOATING
C914 phase_inverter_0/FILLER_0_7_2/a_932_472# vss 0.33241f $ **FLOATING
C915 phase_inverter_0/FILLER_0_7_2/a_484_472# vss 0.33241f $ **FLOATING
C916 phase_inverter_0/FILLER_0_7_2/a_36_472# vss 0.404746f
C917 phase_inverter_0/FILLER_0_7_2/a_6844_375# vss 0.233068f $ **FLOATING
C918 phase_inverter_0/FILLER_0_7_2/a_6396_375# vss 0.171644f $ **FLOATING
C919 phase_inverter_0/FILLER_0_7_2/a_5948_375# vss 0.171644f $ **FLOATING
C920 phase_inverter_0/FILLER_0_7_2/a_5500_375# vss 0.171644f $ **FLOATING
C921 phase_inverter_0/FILLER_0_7_2/a_5052_375# vss 0.171644f $ **FLOATING
C922 phase_inverter_0/FILLER_0_7_2/a_4604_375# vss 0.171644f $ **FLOATING
C923 phase_inverter_0/FILLER_0_7_2/a_4156_375# vss 0.171644f $ **FLOATING
C924 phase_inverter_0/FILLER_0_7_2/a_3708_375# vss 0.171644f $ **FLOATING
C925 phase_inverter_0/FILLER_0_7_2/a_3260_375# vss 0.171644f $ **FLOATING
C926 phase_inverter_0/FILLER_0_7_2/a_2812_375# vss 0.171644f $ **FLOATING
C927 phase_inverter_0/FILLER_0_7_2/a_2364_375# vss 0.171644f $ **FLOATING
C928 phase_inverter_0/FILLER_0_7_2/a_1916_375# vss 0.171644f $ **FLOATING
C929 phase_inverter_0/FILLER_0_7_2/a_1468_375# vss 0.171644f $ **FLOATING
C930 phase_inverter_0/FILLER_0_7_2/a_1020_375# vss 0.171644f $ **FLOATING
C931 phase_inverter_0/FILLER_0_7_2/a_572_375# vss 0.171644f $ **FLOATING
C932 phase_inverter_0/FILLER_0_7_2/a_124_375# vss 0.185708f $ **FLOATING
C933 phase_inverter_0/output13/a_224_472# vss 2.38465f
C934 phase_inverter_0/FILLER_0_8_107/a_484_472# vss 0.345058f $ **FLOATING
C935 phase_inverter_0/FILLER_0_8_107/a_36_472# vss 0.404746f
C936 phase_inverter_0/FILLER_0_8_107/a_572_375# vss 0.232991f
C937 phase_inverter_0/FILLER_0_8_107/a_124_375# vss 0.185089f $ **FLOATING
C938 phase_inverter_0/output24/a_224_472# vss 2.38465f
C939 phase_inverter_0/FILLER_0_10_12/a_1380_472# vss 0.345058f $ **FLOATING
C940 phase_inverter_0/FILLER_0_10_12/a_932_472# vss 0.33241f $ **FLOATING
C941 phase_inverter_0/FILLER_0_10_12/a_484_472# vss 0.33241f $ **FLOATING
C942 phase_inverter_0/FILLER_0_10_12/a_36_472# vss 0.404746f
C943 phase_inverter_0/FILLER_0_10_12/a_1468_375# vss 0.233029f
C944 phase_inverter_0/FILLER_0_10_12/a_1020_375# vss 0.171606f $ **FLOATING
C945 phase_inverter_0/FILLER_0_10_12/a_572_375# vss 0.171606f $ **FLOATING
C946 phase_inverter_0/FILLER_0_10_12/a_124_375# vss 0.185399f $ **FLOATING
C947 phase_inverter_0/FILLER_0_13_66/a_36_472# vss 0.417394f
C948 phase_inverter_0/FILLER_0_13_66/a_124_375# vss 0.246306f $ **FLOATING
C949 phase_inverter_0/_02_/ZN vss 1.077381f
C950 phase_inverter_0/output12/a_224_472# vss 2.38465f
C951 phase_inverter_0/output23/a_224_472# vss 2.38465f
C952 phase_inverter_0/FILLER_0_12_101/a_36_472# vss 0.417394f
C953 phase_inverter_0/FILLER_0_12_101/a_124_375# vss 0.246306f $ **FLOATING
C954 carray_in_1/n0 vss 19.828964f
C955 phase_inverter_0/_01_/ZN vss 1.235885f
C956 phase_inverter_0/output11/a_224_472# vss 2.38465f
C957 phase_inverter_0/output22/a_224_472# vss 2.38465f
C958 input_signal[2] vss 0.99345f
C959 phase_inverter_0/FILLER_0_7_72/a_3172_472# vss 0.345058f $ **FLOATING
C960 phase_inverter_0/FILLER_0_7_72/a_2724_472# vss 0.33241f $ **FLOATING
C961 phase_inverter_0/FILLER_0_7_72/a_2276_472# vss 0.33241f $ **FLOATING
C962 phase_inverter_0/FILLER_0_7_72/a_1828_472# vss 0.33241f $ **FLOATING
C963 phase_inverter_0/FILLER_0_7_72/a_1380_472# vss 0.33241f $ **FLOATING
C964 phase_inverter_0/FILLER_0_7_72/a_932_472# vss 0.33241f $ **FLOATING
C965 phase_inverter_0/FILLER_0_7_72/a_484_472# vss 0.33241f $ **FLOATING
C966 phase_inverter_0/FILLER_0_7_72/a_36_472# vss 0.404746f
C967 phase_inverter_0/FILLER_0_7_72/a_3260_375# vss 0.233093f $ **FLOATING
C968 phase_inverter_0/FILLER_0_7_72/a_2812_375# vss 0.17167f $ **FLOATING
C969 phase_inverter_0/FILLER_0_7_72/a_2364_375# vss 0.17167f $ **FLOATING
C970 phase_inverter_0/FILLER_0_7_72/a_1916_375# vss 0.17167f $ **FLOATING
C971 phase_inverter_0/FILLER_0_7_72/a_1468_375# vss 0.17167f $ **FLOATING
C972 phase_inverter_0/FILLER_0_7_72/a_1020_375# vss 0.17167f $ **FLOATING
C973 phase_inverter_0/FILLER_0_7_72/a_572_375# vss 0.17167f $ **FLOATING
C974 phase_inverter_0/FILLER_0_7_72/a_124_375# vss 0.185915f $ **FLOATING
C975 phase_inverter_0/FILLER_0_9_2/a_6756_472# vss 0.345058f $ **FLOATING
C976 phase_inverter_0/FILLER_0_9_2/a_6308_472# vss 0.33241f $ **FLOATING
C977 phase_inverter_0/FILLER_0_9_2/a_5860_472# vss 0.33241f $ **FLOATING
C978 phase_inverter_0/FILLER_0_9_2/a_5412_472# vss 0.33241f $ **FLOATING
C979 phase_inverter_0/FILLER_0_9_2/a_4964_472# vss 0.33241f $ **FLOATING
C980 phase_inverter_0/FILLER_0_9_2/a_4516_472# vss 0.33241f $ **FLOATING
C981 phase_inverter_0/FILLER_0_9_2/a_4068_472# vss 0.33241f $ **FLOATING
C982 phase_inverter_0/FILLER_0_9_2/a_3620_472# vss 0.33241f $ **FLOATING
C983 phase_inverter_0/FILLER_0_9_2/a_3172_472# vss 0.33241f $ **FLOATING
C984 phase_inverter_0/FILLER_0_9_2/a_2724_472# vss 0.33241f $ **FLOATING
C985 phase_inverter_0/FILLER_0_9_2/a_2276_472# vss 0.33241f $ **FLOATING
C986 phase_inverter_0/FILLER_0_9_2/a_1828_472# vss 0.33241f $ **FLOATING
C987 phase_inverter_0/FILLER_0_9_2/a_1380_472# vss 0.33241f $ **FLOATING
C988 phase_inverter_0/FILLER_0_9_2/a_932_472# vss 0.33241f $ **FLOATING
C989 phase_inverter_0/FILLER_0_9_2/a_484_472# vss 0.33241f $ **FLOATING
C990 phase_inverter_0/FILLER_0_9_2/a_36_472# vss 0.404746f
C991 phase_inverter_0/FILLER_0_9_2/a_6844_375# vss 0.233068f $ **FLOATING
C992 phase_inverter_0/FILLER_0_9_2/a_6396_375# vss 0.171644f $ **FLOATING
C993 phase_inverter_0/FILLER_0_9_2/a_5948_375# vss 0.171644f $ **FLOATING
C994 phase_inverter_0/FILLER_0_9_2/a_5500_375# vss 0.171644f $ **FLOATING
C995 phase_inverter_0/FILLER_0_9_2/a_5052_375# vss 0.171644f $ **FLOATING
C996 phase_inverter_0/FILLER_0_9_2/a_4604_375# vss 0.171644f $ **FLOATING
C997 phase_inverter_0/FILLER_0_9_2/a_4156_375# vss 0.171644f $ **FLOATING
C998 phase_inverter_0/FILLER_0_9_2/a_3708_375# vss 0.171644f $ **FLOATING
C999 phase_inverter_0/FILLER_0_9_2/a_3260_375# vss 0.171644f $ **FLOATING
C1000 phase_inverter_0/FILLER_0_9_2/a_2812_375# vss 0.171644f $ **FLOATING
C1001 phase_inverter_0/FILLER_0_9_2/a_2364_375# vss 0.171644f $ **FLOATING
C1002 phase_inverter_0/FILLER_0_9_2/a_1916_375# vss 0.171644f $ **FLOATING
C1003 phase_inverter_0/FILLER_0_9_2/a_1468_375# vss 0.171644f $ **FLOATING
C1004 phase_inverter_0/FILLER_0_9_2/a_1020_375# vss 0.171644f $ **FLOATING
C1005 phase_inverter_0/FILLER_0_9_2/a_572_375# vss 0.171644f $ **FLOATING
C1006 phase_inverter_0/FILLER_0_9_2/a_124_375# vss 0.185708f $ **FLOATING
C1007 carray_in_0/n0 vss 18.960093f
C1008 phase_inverter_0/output21/a_224_472# vss 2.390638f
C1009 phase_inverter_0/_00_/ZN vss 1.56724f
C1010 phase_inverter_0/output20/a_224_472# vss 2.386258f
C1011 phase_inverter_0/FILLER_0_1_72/a_1380_472# vss 0.345058f $ **FLOATING
C1012 phase_inverter_0/FILLER_0_1_72/a_932_472# vss 0.33241f $ **FLOATING
C1013 phase_inverter_0/FILLER_0_1_72/a_484_472# vss 0.33241f $ **FLOATING
C1014 phase_inverter_0/FILLER_0_1_72/a_36_472# vss 0.404746f
C1015 phase_inverter_0/FILLER_0_1_72/a_1468_375# vss 0.233029f
C1016 phase_inverter_0/FILLER_0_1_72/a_1020_375# vss 0.171606f $ **FLOATING
C1017 phase_inverter_0/FILLER_0_1_72/a_572_375# vss 0.172262f $ **FLOATING
C1018 phase_inverter_0/FILLER_0_1_72/a_124_375# vss 0.185399f $ **FLOATING
C1019 carray_in_1/n1 vss 26.054531f
C1020 carray_in_1/n4 vss 40.26557f
C1021 carray_in_1/n5 vss 48.29981f
C1022 carray_in_1/n2 vss 31.908575f
C1023 carray_in_1/n3 vss 34.573807f
C1024 carray_in_1/n9 vss 15.677258f
C1025 inputm vss -0.686844p
C1026 carray_in_1/n8 vss 41.236954f
C1027 carray_in_1/n7 vss 56.976776f
C1028 carray_in_1/n6 vss 53.73989f
C1029 carray_in_0/n1 vss 26.210373f
C1030 carray_in_0/n4 vss 40.29222f
C1031 carray_in_0/n5 vss 48.35306f
C1032 carray_in_0/n2 vss 31.825562f
C1033 carray_in_0/n3 vss 34.694798f
C1034 carray_in_0/n9 vss 15.763344f
C1035 inputp vss -0.686844p
C1036 carray_in_0/n8 vss 41.365013f
C1037 carray_in_0/n7 vss 57.173172f
C1038 carray_in_0/n6 vss 53.727947f
.ends

