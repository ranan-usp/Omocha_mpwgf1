module saradc(
	inout vdd,
	inout vss,
	input vinp,
	input vinn,
	input cal,
	input en,
	input clk,
	input rstn,
	output valid,
	output [9:0] result
);
endmodule