* NGSPICE file created from bootstrapped_sw.ext - technology: gf180mcuD

.subckt XM1_bs G D a_811_3903# S a_1507_3903#
X0 D G S a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM4_bs G D S
X0 D G S S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs1_bs G D S a_n2855_n800#
X0 D G S a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668#
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0fF c_width=8u c_length=8u
.ends

.subckt sw_cap_unit in out
Xcap_mim_2p0fF_8JNR63_0 out in cap_mim_2p0fF_8JNR63
.ends

.subckt sw_cap out in
Xsw_cap_unit_0 in out sw_cap_unit
Xsw_cap_unit_1 in out sw_cap_unit
Xsw_cap_unit_2 in out sw_cap_unit
Xsw_cap_unit_3 in out sw_cap_unit
Xsw_cap_unit_4 in out sw_cap_unit
.ends

.subckt XM3_bs G D S
X0 S G D S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs_bs G D S a_846_4542#
X0 S G D a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM1_bs_inv G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2_bs_inv G D S
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt bs_inv in vdd out vss
XXM1_bs_inv_0 in out vss XM1_bs_inv
XXM2_bs_inv_0 in out vdd XM2_bs_inv
.ends

.subckt XM2_bs G D a_811_3460# a_1507_3460# S
X0 S G D a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs2_bs B G D a_n3988_469# S a_n3988_1165#
X0 D G S a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt bootstrapped_sw vbsl vbsh vs vg in vdd vss en enb out
XXM1_bs_0 vg vbsl vss in vss XM1_bs
XXM4_bs_0 enb vg vbsh XM4_bs
XXMs1_bs_0 vdd vs vg vss XMs1_bs
Xsw_cap_0 vbsh vbsl sw_cap
XXM3_bs_0 vg vdd vbsh XM3_bs
XXMs_bs_0 vg out in vss XMs_bs
Xbs_inv_0 en vdd enb vss bs_inv
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 XMs2_bs_0/B enb vss vss vs vss XMs2_bs
.ends

