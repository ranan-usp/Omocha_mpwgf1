magic
tech gf180mcuD
magscale 1 5
timestamp 1702006703
<< obsm1 >>
rect 672 1538 9376 8262
<< obsm2 >>
rect 854 849 9362 9231
<< metal3 >>
rect 9600 9184 10000 9240
rect 0 8960 400 9016
rect 9600 8736 10000 8792
rect 9600 8288 10000 8344
rect 0 8064 400 8120
rect 9600 7840 10000 7896
rect 9600 7392 10000 7448
rect 0 7168 400 7224
rect 9600 6944 10000 7000
rect 9600 6496 10000 6552
rect 0 6272 400 6328
rect 9600 6048 10000 6104
rect 9600 5600 10000 5656
rect 0 5376 400 5432
rect 9600 5152 10000 5208
rect 9600 4704 10000 4760
rect 0 4480 400 4536
rect 9600 4256 10000 4312
rect 9600 3808 10000 3864
rect 0 3584 400 3640
rect 9600 3360 10000 3416
rect 9600 2912 10000 2968
rect 0 2688 400 2744
rect 9600 2464 10000 2520
rect 9600 2016 10000 2072
rect 0 1792 400 1848
rect 9600 1568 10000 1624
rect 9600 1120 10000 1176
rect 0 896 400 952
rect 9600 672 10000 728
<< obsm3 >>
rect 400 9154 9570 9226
rect 400 9046 9600 9154
rect 430 8930 9600 9046
rect 400 8822 9600 8930
rect 400 8706 9570 8822
rect 400 8374 9600 8706
rect 400 8258 9570 8374
rect 400 8150 9600 8258
rect 430 8034 9600 8150
rect 400 7926 9600 8034
rect 400 7810 9570 7926
rect 400 7478 9600 7810
rect 400 7362 9570 7478
rect 400 7254 9600 7362
rect 430 7138 9600 7254
rect 400 7030 9600 7138
rect 400 6914 9570 7030
rect 400 6582 9600 6914
rect 400 6466 9570 6582
rect 400 6358 9600 6466
rect 430 6242 9600 6358
rect 400 6134 9600 6242
rect 400 6018 9570 6134
rect 400 5686 9600 6018
rect 400 5570 9570 5686
rect 400 5462 9600 5570
rect 430 5346 9600 5462
rect 400 5238 9600 5346
rect 400 5122 9570 5238
rect 400 4790 9600 5122
rect 400 4674 9570 4790
rect 400 4566 9600 4674
rect 430 4450 9600 4566
rect 400 4342 9600 4450
rect 400 4226 9570 4342
rect 400 3894 9600 4226
rect 400 3778 9570 3894
rect 400 3670 9600 3778
rect 430 3554 9600 3670
rect 400 3446 9600 3554
rect 400 3330 9570 3446
rect 400 2998 9600 3330
rect 400 2882 9570 2998
rect 400 2774 9600 2882
rect 430 2658 9600 2774
rect 400 2550 9600 2658
rect 400 2434 9570 2550
rect 400 2102 9600 2434
rect 400 1986 9570 2102
rect 400 1878 9600 1986
rect 430 1762 9600 1878
rect 400 1654 9600 1762
rect 400 1538 9570 1654
rect 400 1206 9600 1538
rect 400 1090 9570 1206
rect 400 982 9600 1090
rect 430 866 9600 982
rect 400 758 9600 866
rect 400 686 9570 758
<< metal4 >>
rect 1670 1538 1830 8262
rect 2748 1538 2908 8262
rect 3826 1538 3986 8262
rect 4904 1538 5064 8262
rect 5982 1538 6142 8262
rect 7060 1538 7220 8262
rect 8138 1538 8298 8262
rect 9216 1538 9376 8262
<< labels >>
rlabel metal3 s 0 896 400 952 6 input_signal[0]
port 1 nsew signal input
rlabel metal3 s 0 1792 400 1848 6 input_signal[1]
port 2 nsew signal input
rlabel metal3 s 0 2688 400 2744 6 input_signal[2]
port 3 nsew signal input
rlabel metal3 s 0 3584 400 3640 6 input_signal[3]
port 4 nsew signal input
rlabel metal3 s 0 4480 400 4536 6 input_signal[4]
port 5 nsew signal input
rlabel metal3 s 0 5376 400 5432 6 input_signal[5]
port 6 nsew signal input
rlabel metal3 s 0 6272 400 6328 6 input_signal[6]
port 7 nsew signal input
rlabel metal3 s 0 7168 400 7224 6 input_signal[7]
port 8 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 input_signal[8]
port 9 nsew signal input
rlabel metal3 s 0 8960 400 9016 6 input_signal[9]
port 10 nsew signal input
rlabel metal3 s 9600 672 10000 728 6 output_signal_minus[0]
port 11 nsew signal output
rlabel metal3 s 9600 4704 10000 4760 6 output_signal_minus[1]
port 12 nsew signal output
rlabel metal3 s 9600 4256 10000 4312 6 output_signal_minus[2]
port 13 nsew signal output
rlabel metal3 s 9600 3808 10000 3864 6 output_signal_minus[3]
port 14 nsew signal output
rlabel metal3 s 9600 3360 10000 3416 6 output_signal_minus[4]
port 15 nsew signal output
rlabel metal3 s 9600 2912 10000 2968 6 output_signal_minus[5]
port 16 nsew signal output
rlabel metal3 s 9600 2464 10000 2520 6 output_signal_minus[6]
port 17 nsew signal output
rlabel metal3 s 9600 2016 10000 2072 6 output_signal_minus[7]
port 18 nsew signal output
rlabel metal3 s 9600 1568 10000 1624 6 output_signal_minus[8]
port 19 nsew signal output
rlabel metal3 s 9600 1120 10000 1176 6 output_signal_minus[9]
port 20 nsew signal output
rlabel metal3 s 9600 9184 10000 9240 6 output_signal_plus[0]
port 21 nsew signal output
rlabel metal3 s 9600 5152 10000 5208 6 output_signal_plus[1]
port 22 nsew signal output
rlabel metal3 s 9600 5600 10000 5656 6 output_signal_plus[2]
port 23 nsew signal output
rlabel metal3 s 9600 6048 10000 6104 6 output_signal_plus[3]
port 24 nsew signal output
rlabel metal3 s 9600 6496 10000 6552 6 output_signal_plus[4]
port 25 nsew signal output
rlabel metal3 s 9600 6944 10000 7000 6 output_signal_plus[5]
port 26 nsew signal output
rlabel metal3 s 9600 7392 10000 7448 6 output_signal_plus[6]
port 27 nsew signal output
rlabel metal3 s 9600 7840 10000 7896 6 output_signal_plus[7]
port 28 nsew signal output
rlabel metal3 s 9600 8288 10000 8344 6 output_signal_plus[8]
port 29 nsew signal output
rlabel metal3 s 9600 8736 10000 8792 6 output_signal_plus[9]
port 30 nsew signal output
rlabel metal4 s 1670 1538 1830 8262 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 8262 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 8262 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 8262 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 8262 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 8262 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 8262 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 8262 6 vss
port 32 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 192562
string GDS_FILE /home/oe23ranan/gf_analog/openlane/phase_inverter/runs/23_12_08_12_37/results/signoff/phase_inverter.magic.gds
string GDS_START 65302
<< end >>

