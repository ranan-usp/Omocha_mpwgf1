* NGSPICE file created from dac.ext - technology: gf180mcuD

.subckt XM1_bs G D a_811_3903# S a_1507_3903#
X0 D G S a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM4_bs G D S
X0 D G S S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs1_bs G D S a_n2855_n800#
X0 D G S a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668#
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0fF c_width=8u c_length=8u
.ends

.subckt sw_cap_unit in out
Xcap_mim_2p0fF_8JNR63_0 out in cap_mim_2p0fF_8JNR63
.ends

.subckt sw_cap out in
Xsw_cap_unit_0 in out sw_cap_unit
Xsw_cap_unit_1 in out sw_cap_unit
Xsw_cap_unit_2 in out sw_cap_unit
Xsw_cap_unit_3 in out sw_cap_unit
Xsw_cap_unit_4 in out sw_cap_unit
.ends

.subckt XM3_bs G D S
X0 S G D S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs_bs G D S a_846_4542#
X0 S G D a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XM1_bs_inv G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt XM2_bs_inv G D S
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt bs_inv in vdd out vss
XXM1_bs_inv_0 in out vss XM1_bs_inv
XXM2_bs_inv_0 in out vdd XM2_bs_inv
.ends

.subckt XM2_bs G D a_811_3460# a_1507_3460# S
X0 S G D a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt XMs2_bs G D a_n3988_469# S a_n3988_1165#
X0 D G S a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
.ends

.subckt bootstrapped_sw vbsl vbsh vs vg in vdd vss en enb out
XXM1_bs_0 vg vbsl vss in vss XM1_bs
XXM4_bs_0 enb vg vbsh XM4_bs
XXMs1_bs_0 vdd vs vg vss XMs1_bs
Xsw_cap_0 vbsh vbsl sw_cap
XXM3_bs_0 vg vdd vbsh XM3_bs
XXMs_bs_0 vg out in vss XMs_bs
Xbs_inv_0 en vdd enb vss bs_inv
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 enb vss vss vs vss XMs2_bs
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
.ends

.subckt inv_renketu inv$1_8/I inv$1_1/I inv$1_4/ZN inv$1_1/ZN inv$1_3/I inv$1_5/I
+ inv$1_7/I inv$1_9/ZN inv$1_6/ZN inv$1_3/ZN inv$1_0/ZN inv$1_0/I inv$1_9/I inv$1_2/I
+ inv$1_10/I inv$1_7/ZN inv$1_4/I inv$1_10/ZN vdd inv$1_8/ZN vss inv$1_6/I inv$1_2/ZN
+ inv$1_5/ZN
Xinv$1_10 vss inv$1_10/ZN inv$1_10/I vdd vdd inv$1_10/VPW vss inv$1
Xinv$1_0 vss inv$1_0/ZN inv$1_0/I vdd vdd inv$1_0/VPW vss inv$1
Xinv$1_1 vss inv$1_1/ZN inv$1_1/I vdd vdd inv$1_1/VPW vss inv$1
Xinv$1_2 vss inv$1_2/ZN inv$1_2/I vdd vdd inv$1_2/VPW vss inv$1
Xinv$1_3 vss inv$1_3/ZN inv$1_3/I vdd vdd inv$1_3/VPW vss inv$1
Xinv$1_4 vss inv$1_4/ZN inv$1_4/I vdd vdd inv$1_4/VPW vss inv$1
Xinv$1_5 vss inv$1_5/ZN inv$1_5/I vdd vdd inv$1_5/VPW vss inv$1
Xinv$1_6 vss inv$1_6/ZN inv$1_6/I vdd vdd inv$1_6/VPW vss inv$1
Xinv$1_7 vss inv$1_7/ZN inv$1_7/I vdd vdd inv$1_7/VPW vss inv$1
Xinv$1_8 vss inv$1_8/ZN inv$1_8/I vdd vdd inv$1_8/VPW vss inv$1
Xinv$1_9 vss inv$1_9/ZN inv$1_9/I vdd vdd inv$1_9/VPW vss inv$1
.ends

.subckt dac vdd vss dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10 in out
+ sample
Xbootstrapped_sw_0 bootstrapped_sw_0/vbsl bootstrapped_sw_0/vbsh bootstrapped_sw_0/vs
+ bootstrapped_sw_0/vg in vdd vss sample bootstrapped_sw_0/enb out bootstrapped_sw
Xinv_renketu_0 ctl7 ctl2 carray_0/n3 carray_0/n2 ctl1 ctl4 ctl6 carray_0/n8 carray_0/n5
+ carray_0/n1 carray_0/ndum dum ctl8 ctl10 ctl9 carray_0/n6 ctl3 carray_0/n9 vdd carray_0/n7
+ vss ctl5 carray_0/n0 carray_0/n4 inv_renketu
.ends

