* NGSPICE file created from dac.ext - technology: gf180mcuD

.subckt XM1_bs G D a_811_3903# S a_1507_3903#
X0 D G S a_811_3903# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S G 0.002993f
C1 S D 0.103318f
C2 G D 0.002993f
C3 S a_811_3903# 0.109266f
C4 G a_811_3903# 0.288275f
C5 D a_811_3903# 0.109266f
.ends

.subckt XM4_bs G D S VSUBS
X0 D G S S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D S 0.127372f
C1 S G 0.180042f
C2 D G 0.002993f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.66703f
.ends

.subckt XMs1_bs G D S a_n2855_n800#
X0 D G S a_n2855_n800# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D G 0.002993f
C1 G S 0.002993f
C2 D S 0.103318f
C3 D a_n2855_n800# 0.109266f
C4 S a_n2855_n800# 0.177295f
C5 G a_n2855_n800# 0.288368f
.ends

.subckt cap_mim_2p0fF_8JNR63 m4_n3440_n548# m4_n3800_n668# VSUBS
X0 m4_n3440_n548# m4_n3800_n668# cap_mim_2f0fF c_width=8u c_length=8u
C0 m4_n3800_n668# m4_n3440_n548# 0.646322f
C1 m4_n3440_n548# VSUBS 1.17298f
C2 m4_n3800_n668# VSUBS 1.64833f
.ends

.subckt sw_cap_unit in out VSUBS
Xcap_mim_2p0fF_8JNR63_0 out in VSUBS cap_mim_2p0fF_8JNR63
C0 out VSUBS 1.17298f
C1 in VSUBS 1.64833f
.ends

.subckt sw_cap out in VSUBS
Xsw_cap_unit_0 in out VSUBS sw_cap_unit
Xsw_cap_unit_1 in out VSUBS sw_cap_unit
Xsw_cap_unit_2 in out VSUBS sw_cap_unit
Xsw_cap_unit_3 in out VSUBS sw_cap_unit
Xsw_cap_unit_4 in out VSUBS sw_cap_unit
C0 in out 2.231591f
C1 out VSUBS 6.064711f
C2 in VSUBS 7.39096f
.ends

.subckt XM3_bs G D S VSUBS
X0 S G D S pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D G 0.002993f
C1 S G 0.175929f
C2 S D 0.127372f
C3 D VSUBS 0.094602f
C4 G VSUBS 0.124463f
C5 S VSUBS 1.68221f
.ends

.subckt XMs_bs G D S a_846_4542#
X0 S G D a_846_4542# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 D G 0.002993f
C1 S G 0.002993f
C2 S D 0.103318f
C3 D a_846_4542# 0.387117f
C4 G a_846_4542# 0.288368f
C5 S a_846_4542# 0.109266f
.ends

.subckt XM1_bs_inv G D S
X0 D G S S nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 G D 0.001764f
C1 D S 0.134177f
C2 G S 0.22667f
.ends

.subckt XM2_bs_inv G D S VSUBS
X0 S G D S pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
C0 D G 0.001764f
C1 S G 0.138578f
C2 S D 0.090564f
C3 D VSUBS 0.043675f
C4 G VSUBS 0.08816f
C5 S VSUBS 1.2321f
.ends

.subckt bs_inv in vdd out vss
XXM1_bs_inv_0 in out vss XM1_bs_inv
XXM2_bs_inv_0 in out vdd vss XM2_bs_inv
C0 out in 0.057341f
C1 out vss 0.056311f
C2 in vss 0.019395f
C3 vdd out 0.086562f
C4 vdd in 0.034991f
C5 vdd vss 0.050184f
C6 vss 0 0.154858f
C7 vdd 0 1.342913f
C8 out 0 0.461919f
C9 in 0 0.440696f
.ends

.subckt XM2_bs G D a_811_3460# a_1507_3460# S
X0 S G D a_811_3460# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 G S 0.002993f
C1 G D 0.002993f
C2 D S 0.103318f
C3 D a_811_3460# 0.109266f
C4 G a_811_3460# 0.288275f
C5 S a_811_3460# 0.109266f
.ends

.subckt XMs2_bs G D a_n3988_469# S a_n3988_1165#
X0 D G S a_n3988_469# nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.5u
C0 S G 0.002993f
C1 S D 0.103318f
C2 D G 0.002993f
C3 D a_n3988_469# 0.109266f
C4 S a_n3988_469# 0.109266f
C5 G a_n3988_469# 0.288275f
.ends

.subckt bootstrapped_sw vs vg in vdd vss en enb out vbsh vbsl
XXM1_bs_0 vg vbsl vss in vss XM1_bs
XXM4_bs_0 enb vg vbsh vss XM4_bs
XXMs1_bs_0 vdd vs vg vss XMs1_bs
Xsw_cap_0 vbsh vbsl vss sw_cap
XXM3_bs_0 vg vdd vbsh vss XM3_bs
XXMs_bs_0 vg out in vss XMs_bs
Xbs_inv_0 en vdd enb vss bs_inv
XXM2_bs_0 enb vbsl vss vss vss XM2_bs
XXMs2_bs_0 enb vss vss vs vss XMs2_bs
C0 en enb 0.025502f
C1 vbsh out 0.106418f
C2 vbsh vdd 0.216342f
C3 vbsl out 0.058082f
C4 out vg 0.04429f
C5 vdd vbsl 0.005409f
C6 vbsh enb 0.079647f
C7 vdd vg 0.447811f
C8 vs vbsl 0.001422f
C9 vbsl enb 0.017274f
C10 vs vg 0.01049f
C11 enb vg 0.612108f
C12 vdd out 0.017908f
C13 vbsh in 0.008752f
C14 in vbsl 0.299565f
C15 vdd enb 0.448382f
C16 in vg 0.075595f
C17 vbsh vbsl 0.035648f
C18 vs enb 0.00376f
C19 vbsh vg 0.225467f
C20 vdd en 0.062309f
C21 vbsl vg 0.046114f
C22 vs vss 0.072259f
C23 enb vss 1.595622f
C24 vdd vss 3.10752f
C25 en vss 0.636177f
C26 out vss 1.088543f
C27 vg vss 1.218874f
C28 vbsh vss 9.044386f
C29 vbsl vss 8.368301f
C30 in vss 0.308876f
.ends

.subckt inv$1 VSS ZN I VDD VNW VPW VSUBS
X0 VDD I ZN VNW pfet_06v0 ad=1.2078p pd=4.42u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.2255p pd=1.37u as=0.5084p ps=2.88u w=0.82u l=0.6u
X2 VSS I ZN VSUBS nfet_06v0 ad=0.8118p pd=3.62u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.7564p ps=3.68u w=1.22u l=0.5u
C0 VDD VSS 0.029045f
C1 VDD VNW 0.082022f
C2 VNW VSS 0.006277f
C3 VNW I 0.285482f
C4 VDD I 0.074838f
C5 VSS I 0.091531f
C6 VDD ZN 0.271625f
C7 VNW ZN 0.023676f
C8 VSS ZN 0.180794f
C9 I ZN 0.58604f
C10 VSS VSUBS 0.296769f
C11 ZN VSUBS 0.099188f
C12 VDD VSUBS 0.238483f
C13 I VSUBS 0.610668f
C14 VNW VSUBS 1.31158f
.ends

.subckt inv_renketu inv$1_8/I inv$1_1/I inv$1_4/ZN inv$1_1/ZN inv$1_3/I inv$1_5/I
+ inv$1_7/I inv$1_9/ZN inv$1_6/ZN inv$1_3/ZN inv$1_0/ZN inv$1_0/I inv$1_9/I inv$1_2/I
+ inv$1_10/I inv$1_7/ZN inv$1_4/I inv$1_10/ZN vdd inv$1_8/ZN vss inv$1_6/I inv$1_2/ZN
+ inv$1_5/ZN
Xinv$1_10 vss inv$1_10/ZN inv$1_10/I vdd vdd inv$1_10/VPW vss inv$1
Xinv$1_0 vss inv$1_0/ZN inv$1_0/I vdd vdd inv$1_0/VPW vss inv$1
Xinv$1_1 vss inv$1_1/ZN inv$1_1/I vdd vdd inv$1_1/VPW vss inv$1
Xinv$1_2 vss inv$1_2/ZN inv$1_2/I vdd vdd inv$1_2/VPW vss inv$1
Xinv$1_3 vss inv$1_3/ZN inv$1_3/I vdd vdd inv$1_3/VPW vss inv$1
Xinv$1_4 vss inv$1_4/ZN inv$1_4/I vdd vdd inv$1_4/VPW vss inv$1
Xinv$1_5 vss inv$1_5/ZN inv$1_5/I vdd vdd inv$1_5/VPW vss inv$1
Xinv$1_6 vss inv$1_6/ZN inv$1_6/I vdd vdd inv$1_6/VPW vss inv$1
Xinv$1_7 vss inv$1_7/ZN inv$1_7/I vdd vdd inv$1_7/VPW vss inv$1
Xinv$1_8 vss inv$1_8/ZN inv$1_8/I vdd vdd inv$1_8/VPW vss inv$1
Xinv$1_9 vss inv$1_9/ZN inv$1_9/I vdd vdd inv$1_9/VPW vss inv$1
C0 vss inv$1_5/I 0.166388f
C1 vdd inv$1_1/I 0.019437f
C2 inv$1_4/I inv$1_5/ZN 0.028928f
C3 inv$1_10/ZN inv$1_10/I 0.029333f
C4 vss inv$1_10/I 0.166388f
C5 inv$1_8/ZN inv$1_9/I 0.002086f
C6 inv$1_10/ZN vdd 0.159176f
C7 vdd vss 0.009518f
C8 inv$1_2/ZN inv$1_10/I 0.028928f
C9 inv$1_6/I inv$1_6/ZN 0.029333f
C10 inv$1_0/I vss 0.170492f
C11 inv$1_2/ZN vdd 0.174722f
C12 vss inv$1_8/I 0.166388f
C13 inv$1_10/ZN inv$1_9/ZN 0.080571f
C14 vss inv$1_9/ZN 0.003326f
C15 inv$1_4/I inv$1_4/ZN 0.029333f
C16 vss inv$1_7/ZN 0.003326f
C17 inv$1_3/ZN inv$1_3/I 0.029333f
C18 inv$1_4/ZN inv$1_5/ZN 0.080571f
C19 inv$1_6/ZN inv$1_7/I 0.002086f
C20 inv$1_6/ZN inv$1_5/ZN 0.080571f
C21 inv$1_1/ZN inv$1_1/I 0.029333f
C22 inv$1_0/ZN vdd 0.184001f
C23 inv$1_0/I inv$1_0/ZN 0.029333f
C24 vss inv$1_8/ZN 0.003326f
C25 inv$1_10/ZN inv$1_2/I 0.002086f
C26 inv$1_2/I vss 0.164788f
C27 inv$1_2/ZN inv$1_2/I 0.029333f
C28 inv$1_1/ZN vss 0.003326f
C29 vdd inv$1_5/I 0.019437f
C30 inv$1_6/I vss 0.166388f
C31 inv$1_1/I inv$1_4/I 0.084161f
C32 vdd inv$1_10/I 0.019437f
C33 inv$1_3/ZN inv$1_1/I 0.002086f
C34 inv$1_0/I vdd 0.026972f
C35 vdd inv$1_8/I 0.019437f
C36 inv$1_4/I vss 0.166388f
C37 inv$1_9/ZN inv$1_10/I 0.002086f
C38 vdd inv$1_9/ZN 0.159176f
C39 vss inv$1_7/I 0.166388f
C40 inv$1_9/ZN inv$1_8/I 0.028928f
C41 vdd inv$1_7/ZN 0.159176f
C42 inv$1_3/ZN vss 0.003326f
C43 vss inv$1_5/ZN 0.003326f
C44 inv$1_7/ZN inv$1_8/I 0.002086f
C45 inv$1_3/I inv$1_1/I 0.084161f
C46 inv$1_1/I inv$1_4/ZN 0.028928f
C47 inv$1_2/I inv$1_10/I 0.084161f
C48 vdd inv$1_8/ZN 0.159176f
C49 inv$1_2/I vdd 0.035575f
C50 inv$1_3/I vss 0.166388f
C51 inv$1_8/ZN inv$1_8/I 0.029333f
C52 inv$1_8/ZN inv$1_9/ZN 0.080571f
C53 inv$1_4/ZN vss 0.003326f
C54 inv$1_6/I inv$1_5/I 0.084161f
C55 inv$1_3/ZN inv$1_0/ZN 0.080571f
C56 inv$1_7/ZN inv$1_8/ZN 0.080571f
C57 inv$1_1/ZN vdd 0.159176f
C58 vss inv$1_6/ZN 0.003326f
C59 inv$1_4/I inv$1_5/I 0.084161f
C60 inv$1_0/ZN inv$1_3/I 0.002086f
C61 vdd inv$1_6/I 0.019437f
C62 inv$1_5/I inv$1_5/ZN 0.029333f
C63 inv$1_6/I inv$1_7/ZN 0.028928f
C64 inv$1_10/ZN inv$1_9/I 0.028928f
C65 vss inv$1_9/I 0.166388f
C66 vdd inv$1_4/I 0.019437f
C67 vdd inv$1_7/I 0.019437f
C68 inv$1_8/I inv$1_7/I 0.084161f
C69 inv$1_3/ZN vdd 0.159176f
C70 vdd inv$1_5/ZN 0.159176f
C71 inv$1_0/I inv$1_3/ZN 0.028928f
C72 inv$1_4/ZN inv$1_5/I 0.002086f
C73 inv$1_1/I vss 0.166388f
C74 inv$1_7/ZN inv$1_7/I 0.029333f
C75 inv$1_6/ZN inv$1_5/I 0.028928f
C76 inv$1_3/I vdd 0.019437f
C77 inv$1_0/I inv$1_3/I 0.08416f
C78 inv$1_10/ZN vss 0.003326f
C79 inv$1_10/ZN inv$1_2/ZN 0.080571f
C80 inv$1_2/ZN vss 0.005014f
C81 inv$1_8/ZN inv$1_7/I 0.028928f
C82 vdd inv$1_4/ZN 0.159176f
C83 vdd inv$1_6/ZN 0.159176f
C84 inv$1_1/ZN inv$1_4/I 0.002086f
C85 inv$1_1/ZN inv$1_3/ZN 0.080571f
C86 inv$1_7/ZN inv$1_6/ZN 0.080571f
C87 inv$1_0/ZN vss 0.005399f
C88 inv$1_6/I inv$1_7/I 0.084161f
C89 inv$1_9/I inv$1_10/I 0.084161f
C90 inv$1_1/ZN inv$1_3/I 0.028928f
C91 inv$1_6/I inv$1_5/ZN 0.002086f
C92 vdd inv$1_9/I 0.019437f
C93 inv$1_9/I inv$1_8/I 0.084161f
C94 inv$1_1/ZN inv$1_4/ZN 0.080571f
C95 inv$1_9/ZN inv$1_9/I 0.029333f
C96 inv$1_9/ZN 0 0.131999f
C97 inv$1_9/I 0 0.64919f
C98 inv$1_8/ZN 0 0.131999f
C99 inv$1_8/I 0 0.64919f
C100 inv$1_7/ZN 0 0.131999f
C101 inv$1_7/I 0 0.64919f
C102 inv$1_6/ZN 0 0.131999f
C103 inv$1_6/I 0 0.64919f
C104 inv$1_5/ZN 0 0.131999f
C105 inv$1_5/I 0 0.64919f
C106 inv$1_4/ZN 0 0.131999f
C107 inv$1_4/I 0 0.64919f
C108 inv$1_3/ZN 0 0.131999f
C109 inv$1_3/I 0 0.64919f
C110 vss 0 3.02573f
C111 inv$1_2/ZN 0 0.206166f
C112 vdd 0 16.013325f
C113 inv$1_2/I 0 0.750024f
C114 inv$1_1/ZN 0 0.131999f
C115 inv$1_1/I 0 0.64919f
C116 inv$1_0/ZN 0 0.209411f
C117 inv$1_0/I 0 0.731246f
C118 inv$1_10/ZN 0 0.131999f
C119 inv$1_10/I 0 0.64919f
.ends

.subckt dac vdd vss dum ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 ctl8 ctl9 ctl10 in out
+ sample
Xbootstrapped_sw_0 bootstrapped_sw_0/vs bootstrapped_sw_0/vg in vdd vss sample bootstrapped_sw_0/enb
+ out bootstrapped_sw_0/vbsh bootstrapped_sw_0/vbsl bootstrapped_sw
Xinv_renketu_0 ctl7 ctl2 carray_0/n3 carray_0/n2 ctl1 ctl4 ctl6 carray_0/n8 carray_0/n5
+ carray_0/n1 carray_0/ndum dum ctl8 ctl10 ctl9 carray_0/n6 ctl3 carray_0/n9 vdd carray_0/n7
+ vss ctl5 carray_0/n0 carray_0/n4 inv_renketu
C0 carray_0/n1 carray_0/n5 0.142354f
C1 carray_0/n8 carray_0/n9 87.43916f
C2 carray_0/n2 vdd 0.002151f
C3 out carray_0/n4 26.32268f
C4 carray_0/n3 carray_0/n4 26.229404f
C5 vdd carray_0/n5 0.002151f
C6 carray_0/n2 carray_0/ndum 0.041162f
C7 carray_0/n7 carray_0/n4 1.70387f
C8 carray_0/n5 carray_0/ndum 0.025424f
C9 carray_0/n8 carray_0/n0 0.097254f
C10 carray_0/n8 carray_0/n6 11.2161f
C11 ctl2 ctl1 0.104537f
C12 sample carray_0/ndum 0.045492f
C13 carray_0/n9 carray_0/n0 0.521489f
C14 carray_0/n2 carray_0/n5 0.208112f
C15 carray_0/n6 carray_0/n9 14.716781f
C16 carray_0/n1 carray_0/n4 0.142475f
C17 carray_0/n8 out 0.420152p
C18 carray_0/n3 carray_0/n8 1.46111f
C19 carray_0/n6 carray_0/n0 0.025424f
C20 carray_0/n9 out 0.846161p
C21 carray_0/n8 carray_0/n7 50.514606f
C22 carray_0/n3 carray_0/n9 1.911225f
C23 vdd carray_0/n4 0.002151f
C24 carray_0/n7 carray_0/n9 29.51607f
C25 carray_0/n4 carray_0/ndum 0.025424f
C26 ctl4 ctl3 0.104537f
C27 carray_0/n2 carray_0/n4 0.213209f
C28 out carray_0/n0 1.750611f
C29 carray_0/n3 carray_0/n0 0.051666f
C30 carray_0/n6 out 0.105055p
C31 carray_0/n3 carray_0/n6 0.336612f
C32 carray_0/n5 carray_0/n4 27.828503f
C33 carray_0/n7 carray_0/n0 0.06073f
C34 carray_0/n6 carray_0/n7 34.66261f
C35 carray_0/n8 carray_0/n1 0.28587f
C36 carray_0/n1 carray_0/n9 0.350042f
C37 bootstrapped_sw_0/vbsh out 0.137967f
C38 carray_0/n8 vdd 0.002151f
C39 carray_0/n3 out 13.201303f
C40 ctl6 ctl7 0.104537f
C41 ctl10 ctl9 0.104537f
C42 vdd carray_0/n9 0.002151f
C43 carray_0/n8 carray_0/ndum 0.097254f
C44 ctl6 ctl5 0.104537f
C45 carray_0/n7 out 0.210032p
C46 ctl4 ctl5 0.104537f
C47 carray_0/n3 carray_0/n7 0.891504f
C48 carray_0/n1 carray_0/n0 8.476913f
C49 carray_0/n1 carray_0/n6 0.142211f
C50 carray_0/n9 carray_0/ndum 0.127951f
C51 carray_0/n8 carray_0/n2 0.770227f
C52 carray_0/n8 carray_0/n5 5.60732f
C53 carray_0/n2 carray_0/n9 0.996681f
C54 vdd carray_0/n0 0.002151f
C55 vdd carray_0/n6 0.002151f
C56 out bootstrapped_sw_0/vbsl 0.061234f
C57 carray_0/n5 carray_0/n9 7.39935f
C58 carray_0/n6 carray_0/ndum 0.025424f
C59 carray_0/n1 out 3.367623f
C60 carray_0/n3 carray_0/n1 0.145048f
C61 carray_0/n2 carray_0/n0 0.099314f
C62 carray_0/n2 carray_0/n6 0.20799f
C63 ctl9 ctl8 0.104537f
C64 carray_0/n1 carray_0/n7 0.212822f
C65 carray_0/n5 carray_0/n0 0.025424f
C66 carray_0/n5 carray_0/n6 28.925903f
C67 carray_0/n3 vdd 0.002151f
C68 vdd carray_0/n7 0.002151f
C69 out carray_0/ndum 1.640173f
C70 carray_0/n3 carray_0/ndum 0.025424f
C71 ctl3 ctl2 0.104537f
C72 carray_0/n8 carray_0/n4 2.84323f
C73 carray_0/n7 carray_0/ndum 0.06073f
C74 carray_0/n2 out 6.640605f
C75 ctl1 dum 0.104537f
C76 carray_0/n3 carray_0/n2 23.177216f
C77 carray_0/n9 carray_0/n4 3.740571f
C78 carray_0/n5 out 52.565495f
C79 carray_0/n2 carray_0/n7 0.485355f
C80 carray_0/n3 carray_0/n5 0.346757f
C81 carray_0/n5 carray_0/n7 3.36878f
C82 carray_0/n1 vdd 0.002151f
C83 carray_0/n4 carray_0/n0 0.040502f
C84 carray_0/n6 carray_0/n4 0.614078f
C85 carray_0/n1 carray_0/ndum 8.4982f
C86 ctl7 ctl8 0.104537f
C87 carray_0/n1 carray_0/n2 16.941956f
C88 vdd carray_0/ndum 0.004405f
C89 ctl8 vss 0.916847f
C90 ctl7 vss 0.916847f
C91 ctl6 vss 0.916847f
C92 ctl5 vss 0.916847f
C93 ctl4 vss 0.916847f
C94 ctl3 vss 0.916847f
C95 ctl1 vss 0.916847f
C96 carray_0/n0 vss 17.398035f
C97 vdd vss 19.487324f
C98 ctl10 vss 1.146163f
C99 ctl2 vss 0.916847f
C100 carray_0/ndum vss 14.881927f
C101 dum vss 1.125528f
C102 ctl9 vss 0.916847f
C103 carray_0/n4 vss 39.983227f
C104 carray_0/n5 vss 47.48966f
C105 carray_0/n9 vss 14.559587f
C106 out vss -0.683569p
C107 carray_0/n8 vss 40.389835f
C108 carray_0/n7 vss 57.16868f
C109 carray_0/n6 vss 53.444874f
C110 carray_0/n2 vss 30.239845f
C111 carray_0/n1 vss 16.427063f
C112 carray_0/n3 vss 33.722244f
C113 bootstrapped_sw_0/vs vss 0.065021f
C114 bootstrapped_sw_0/enb vss 1.52928f
C115 sample vss 20.507322f
C116 bootstrapped_sw_0/vg vss 1.162193f
C117 bootstrapped_sw_0/vbsh vss 9.037161f
C118 bootstrapped_sw_0/vbsl vss 8.446682f
C119 in vss 0.297821f
.ends

